
module ctrl ( clk, rst_n, s_p_flag_in, mux_flag, rotation, demux_flag );
  output [2:0] rotation;
  input clk, rst_n, s_p_flag_in;
  output mux_flag, demux_flag;
  wire   n11, n12, n13, N17, N18, N19, n3, n2, n7, n9, n10;
  wire   [2:0] core_tick;

  DFFRHQX4 rotation_reg_2_ ( .D(core_tick[2]), .CK(clk), .RN(rst_n), .Q(n11)
         );
  DFFRHQX4 rotation_reg_1_ ( .D(core_tick[1]), .CK(clk), .RN(rst_n), .Q(n12)
         );
  DFFRHQX4 rotation_reg_0_ ( .D(core_tick[0]), .CK(clk), .RN(rst_n), .Q(n13)
         );
  DFFRHQX1 core_tick_reg_2_ ( .D(N19), .CK(clk), .RN(rst_n), .Q(core_tick[2])
         );
  DFFRHQX1 core_tick_reg_1_ ( .D(N18), .CK(clk), .RN(rst_n), .Q(core_tick[1])
         );
  DFFRHQX1 core_tick_reg_0_ ( .D(N17), .CK(clk), .RN(rst_n), .Q(core_tick[0])
         );
  DFFRX1 demux_flag_reg ( .D(n10), .CK(clk), .RN(rst_n), .Q(demux_flag) );
  DFFRHQX4 mux_flag_reg ( .D(core_tick[2]), .CK(clk), .RN(rst_n), .Q(mux_flag)
         );
  INVX4 U3 ( .A(n11), .Y(n2) );
  BUFX12 U4 ( .A(n12), .Y(rotation[1]) );
  INVX8 U5 ( .A(n2), .Y(rotation[2]) );
  INVX4 U6 ( .A(n13), .Y(n7) );
  INVX8 U7 ( .A(n7), .Y(rotation[0]) );
  INVX1 U8 ( .A(core_tick[2]), .Y(n10) );
  AOI2BB1X1 U9 ( .A0N(n9), .A1N(core_tick[1]), .B0(core_tick[0]), .Y(N17) );
  OR2X2 U10 ( .A(s_p_flag_in), .B(core_tick[2]), .Y(n9) );
  XOR2X1 U11 ( .A(core_tick[1]), .B(core_tick[0]), .Y(N18) );
  XOR2X1 U12 ( .A(n10), .B(n3), .Y(N19) );
  NAND2X1 U13 ( .A(core_tick[1]), .B(core_tick[0]), .Y(n3) );
endmodule


module s_p ( clk, rst_n, data_in_1, data_out_1, s_p_flag_out );
  input [33:0] data_in_1;
  output [135:0] data_out_1;
  input clk, rst_n;
  output s_p_flag_out;
  wire   N13, N14, N15, N171, n550, n551, n552, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n980, n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n978, n979, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046;
  wire   [3:0] counter;
  wire   [33:0] R15;
  wire   [33:0] R11;
  wire   [33:0] R7;
  wire   [33:0] R3;
  wire   [33:0] R12;
  wire   [33:0] R8;
  wire   [33:0] R4;
  wire   [33:0] R0;
  wire   [33:0] R13;
  wire   [33:0] R9;
  wire   [33:0] R5;
  wire   [33:0] R1;
  wire   [33:0] R14;
  wire   [33:0] R10;
  wire   [33:0] R6;
  wire   [33:0] R2;

  DFFHQX4 data_out_1_reg_135_ ( .D(n832), .CK(clk), .Q(data_out_1[135]) );
  DFFHQX4 data_out_1_reg_118_ ( .D(n849), .CK(clk), .Q(data_out_1[118]) );
  EDFFX1 R15_reg_33_ ( .D(data_in_1[33]), .E(n1032), .CK(clk), .Q(R15[33]) );
  EDFFX1 R15_reg_32_ ( .D(data_in_1[32]), .E(n1032), .CK(clk), .Q(R15[32]) );
  EDFFX1 R15_reg_31_ ( .D(data_in_1[31]), .E(n1032), .CK(clk), .Q(R15[31]) );
  EDFFX1 R15_reg_30_ ( .D(data_in_1[30]), .E(n1032), .CK(clk), .Q(R15[30]) );
  EDFFX1 R15_reg_29_ ( .D(data_in_1[29]), .E(n1032), .CK(clk), .Q(R15[29]) );
  EDFFX1 R15_reg_28_ ( .D(data_in_1[28]), .E(n1032), .CK(clk), .Q(R15[28]) );
  EDFFX1 R15_reg_27_ ( .D(data_in_1[27]), .E(n1032), .CK(clk), .Q(R15[27]) );
  EDFFX1 R15_reg_26_ ( .D(data_in_1[26]), .E(n1032), .CK(clk), .Q(R15[26]) );
  EDFFX1 R15_reg_25_ ( .D(data_in_1[25]), .E(n1032), .CK(clk), .Q(R15[25]) );
  EDFFX1 R15_reg_24_ ( .D(data_in_1[24]), .E(n1029), .CK(clk), .Q(R15[24]) );
  EDFFX1 R15_reg_23_ ( .D(data_in_1[23]), .E(n1029), .CK(clk), .Q(R15[23]) );
  EDFFX1 R15_reg_22_ ( .D(data_in_1[22]), .E(n1032), .CK(clk), .Q(R15[22]) );
  EDFFX1 R15_reg_21_ ( .D(data_in_1[21]), .E(n1032), .CK(clk), .Q(R15[21]) );
  EDFFX1 R15_reg_20_ ( .D(data_in_1[20]), .E(n1031), .CK(clk), .Q(R15[20]) );
  EDFFX1 R15_reg_19_ ( .D(data_in_1[19]), .E(n1030), .CK(clk), .Q(R15[19]) );
  EDFFX1 R15_reg_18_ ( .D(data_in_1[18]), .E(n1029), .CK(clk), .Q(R15[18]) );
  EDFFX1 R15_reg_17_ ( .D(data_in_1[17]), .E(n1031), .CK(clk), .Q(R15[17]) );
  EDFFX1 R15_reg_16_ ( .D(data_in_1[16]), .E(n1032), .CK(clk), .Q(R15[16]) );
  EDFFX1 R15_reg_15_ ( .D(data_in_1[15]), .E(n1031), .CK(clk), .Q(R15[15]) );
  EDFFX1 R15_reg_14_ ( .D(data_in_1[14]), .E(n1031), .CK(clk), .Q(R15[14]) );
  EDFFX1 R15_reg_13_ ( .D(data_in_1[13]), .E(n1030), .CK(clk), .Q(R15[13]) );
  EDFFX1 R15_reg_12_ ( .D(data_in_1[12]), .E(n1029), .CK(clk), .Q(R15[12]) );
  EDFFX1 R15_reg_11_ ( .D(data_in_1[11]), .E(n1030), .CK(clk), .Q(R15[11]) );
  EDFFX1 R15_reg_10_ ( .D(data_in_1[10]), .E(n1032), .CK(clk), .Q(R15[10]) );
  EDFFX1 R15_reg_9_ ( .D(data_in_1[9]), .E(n1030), .CK(clk), .Q(R15[9]) );
  EDFFX1 R15_reg_8_ ( .D(data_in_1[8]), .E(n1031), .CK(clk), .Q(R15[8]) );
  EDFFX1 R15_reg_7_ ( .D(data_in_1[7]), .E(n1030), .CK(clk), .Q(R15[7]) );
  EDFFX1 R15_reg_6_ ( .D(data_in_1[6]), .E(n1029), .CK(clk), .Q(R15[6]) );
  EDFFX1 R15_reg_5_ ( .D(data_in_1[5]), .E(n1032), .CK(clk), .Q(R15[5]) );
  EDFFX1 R15_reg_4_ ( .D(data_in_1[4]), .E(n1032), .CK(clk), .Q(R15[4]) );
  EDFFX1 R15_reg_3_ ( .D(data_in_1[3]), .E(n1030), .CK(clk), .Q(R15[3]) );
  EDFFX1 R15_reg_2_ ( .D(data_in_1[2]), .E(n1029), .CK(clk), .Q(R15[2]) );
  EDFFX1 R15_reg_1_ ( .D(data_in_1[1]), .E(n1029), .CK(clk), .Q(R15[1]) );
  EDFFX1 R15_reg_0_ ( .D(data_in_1[0]), .E(n1032), .CK(clk), .Q(R15[0]) );
  EDFFX1 R3_reg_33_ ( .D(data_in_1[33]), .E(n984), .CK(clk), .Q(R3[33]) );
  EDFFX1 R3_reg_32_ ( .D(data_in_1[32]), .E(n984), .CK(clk), .Q(R3[32]) );
  EDFFX1 R3_reg_31_ ( .D(data_in_1[31]), .E(n984), .CK(clk), .Q(R3[31]) );
  EDFFX1 R3_reg_30_ ( .D(data_in_1[30]), .E(n984), .CK(clk), .Q(R3[30]) );
  EDFFX1 R3_reg_29_ ( .D(data_in_1[29]), .E(n984), .CK(clk), .Q(R3[29]) );
  EDFFX1 R3_reg_28_ ( .D(data_in_1[28]), .E(n984), .CK(clk), .Q(R3[28]) );
  EDFFX1 R3_reg_27_ ( .D(data_in_1[27]), .E(n984), .CK(clk), .Q(R3[27]) );
  EDFFX1 R3_reg_26_ ( .D(data_in_1[26]), .E(n984), .CK(clk), .Q(R3[26]) );
  EDFFX1 R3_reg_25_ ( .D(data_in_1[25]), .E(n984), .CK(clk), .Q(R3[25]) );
  EDFFX1 R3_reg_24_ ( .D(data_in_1[24]), .E(n984), .CK(clk), .Q(R3[24]) );
  EDFFX1 R3_reg_23_ ( .D(data_in_1[23]), .E(n984), .CK(clk), .Q(R3[23]) );
  EDFFX1 R3_reg_22_ ( .D(data_in_1[22]), .E(n984), .CK(clk), .Q(R3[22]) );
  EDFFX1 R3_reg_21_ ( .D(data_in_1[21]), .E(n985), .CK(clk), .Q(R3[21]) );
  EDFFX1 R3_reg_20_ ( .D(data_in_1[20]), .E(n985), .CK(clk), .Q(R3[20]) );
  EDFFX1 R3_reg_19_ ( .D(data_in_1[19]), .E(n985), .CK(clk), .Q(R3[19]) );
  EDFFX1 R3_reg_18_ ( .D(data_in_1[18]), .E(n985), .CK(clk), .Q(R3[18]) );
  EDFFX1 R3_reg_17_ ( .D(data_in_1[17]), .E(n985), .CK(clk), .Q(R3[17]) );
  EDFFX1 R3_reg_16_ ( .D(data_in_1[16]), .E(n985), .CK(clk), .Q(R3[16]) );
  EDFFX1 R3_reg_15_ ( .D(data_in_1[15]), .E(n985), .CK(clk), .Q(R3[15]) );
  EDFFX1 R3_reg_14_ ( .D(data_in_1[14]), .E(n985), .CK(clk), .Q(R3[14]) );
  EDFFX1 R3_reg_13_ ( .D(data_in_1[13]), .E(n985), .CK(clk), .Q(R3[13]) );
  EDFFX1 R3_reg_12_ ( .D(data_in_1[12]), .E(n985), .CK(clk), .Q(R3[12]) );
  EDFFX1 R3_reg_11_ ( .D(data_in_1[11]), .E(n985), .CK(clk), .Q(R3[11]) );
  EDFFX1 R3_reg_10_ ( .D(data_in_1[10]), .E(n985), .CK(clk), .Q(R3[10]) );
  EDFFX1 R3_reg_9_ ( .D(data_in_1[9]), .E(n984), .CK(clk), .Q(R3[9]) );
  EDFFX1 R3_reg_8_ ( .D(data_in_1[8]), .E(n985), .CK(clk), .Q(R3[8]) );
  EDFFX1 R3_reg_7_ ( .D(data_in_1[7]), .E(n984), .CK(clk), .Q(R3[7]) );
  EDFFX1 R3_reg_6_ ( .D(data_in_1[6]), .E(n985), .CK(clk), .Q(R3[6]) );
  EDFFX1 R3_reg_5_ ( .D(data_in_1[5]), .E(n984), .CK(clk), .Q(R3[5]) );
  EDFFX1 R3_reg_4_ ( .D(data_in_1[4]), .E(n985), .CK(clk), .Q(R3[4]) );
  EDFFX1 R3_reg_3_ ( .D(data_in_1[3]), .E(n984), .CK(clk), .Q(R3[3]) );
  EDFFX1 R3_reg_2_ ( .D(data_in_1[2]), .E(n985), .CK(clk), .Q(R3[2]) );
  EDFFX1 R3_reg_1_ ( .D(data_in_1[1]), .E(n984), .CK(clk), .Q(R3[1]) );
  EDFFX1 R3_reg_0_ ( .D(data_in_1[0]), .E(n985), .CK(clk), .Q(R3[0]) );
  EDFFX1 R7_reg_33_ ( .D(data_in_1[33]), .E(n992), .CK(clk), .Q(R7[33]) );
  EDFFX1 R7_reg_32_ ( .D(data_in_1[32]), .E(n993), .CK(clk), .Q(R7[32]) );
  EDFFX1 R7_reg_31_ ( .D(data_in_1[31]), .E(n992), .CK(clk), .Q(R7[31]) );
  EDFFX1 R7_reg_30_ ( .D(data_in_1[30]), .E(n993), .CK(clk), .Q(R7[30]) );
  EDFFX1 R7_reg_29_ ( .D(data_in_1[29]), .E(n992), .CK(clk), .Q(R7[29]) );
  EDFFX1 R7_reg_28_ ( .D(data_in_1[28]), .E(n993), .CK(clk), .Q(R7[28]) );
  EDFFX1 R7_reg_27_ ( .D(data_in_1[27]), .E(n992), .CK(clk), .Q(R7[27]) );
  EDFFX1 R7_reg_26_ ( .D(data_in_1[26]), .E(n993), .CK(clk), .Q(R7[26]) );
  EDFFX1 R7_reg_25_ ( .D(data_in_1[25]), .E(n992), .CK(clk), .Q(R7[25]) );
  EDFFX1 R7_reg_24_ ( .D(data_in_1[24]), .E(n993), .CK(clk), .Q(R7[24]) );
  EDFFX1 R7_reg_23_ ( .D(data_in_1[23]), .E(n993), .CK(clk), .Q(R7[23]) );
  EDFFX1 R7_reg_22_ ( .D(data_in_1[22]), .E(n993), .CK(clk), .Q(R7[22]) );
  EDFFX1 R7_reg_21_ ( .D(data_in_1[21]), .E(n993), .CK(clk), .Q(R7[21]) );
  EDFFX1 R7_reg_20_ ( .D(data_in_1[20]), .E(n993), .CK(clk), .Q(R7[20]) );
  EDFFX1 R7_reg_19_ ( .D(data_in_1[19]), .E(n993), .CK(clk), .Q(R7[19]) );
  EDFFX1 R7_reg_18_ ( .D(data_in_1[18]), .E(n993), .CK(clk), .Q(R7[18]) );
  EDFFX1 R7_reg_17_ ( .D(data_in_1[17]), .E(n993), .CK(clk), .Q(R7[17]) );
  EDFFX1 R7_reg_16_ ( .D(data_in_1[16]), .E(n993), .CK(clk), .Q(R7[16]) );
  EDFFX1 R7_reg_15_ ( .D(data_in_1[15]), .E(n993), .CK(clk), .Q(R7[15]) );
  EDFFX1 R7_reg_14_ ( .D(data_in_1[14]), .E(n993), .CK(clk), .Q(R7[14]) );
  EDFFX1 R7_reg_13_ ( .D(data_in_1[13]), .E(n993), .CK(clk), .Q(R7[13]) );
  EDFFX1 R7_reg_12_ ( .D(data_in_1[12]), .E(n993), .CK(clk), .Q(R7[12]) );
  EDFFX1 R7_reg_11_ ( .D(data_in_1[11]), .E(n992), .CK(clk), .Q(R7[11]) );
  EDFFX1 R7_reg_10_ ( .D(data_in_1[10]), .E(n992), .CK(clk), .Q(R7[10]) );
  EDFFX1 R7_reg_9_ ( .D(data_in_1[9]), .E(n992), .CK(clk), .Q(R7[9]) );
  EDFFX1 R7_reg_8_ ( .D(data_in_1[8]), .E(n992), .CK(clk), .Q(R7[8]) );
  EDFFX1 R7_reg_7_ ( .D(data_in_1[7]), .E(n992), .CK(clk), .Q(R7[7]) );
  EDFFX1 R7_reg_6_ ( .D(data_in_1[6]), .E(n992), .CK(clk), .Q(R7[6]) );
  EDFFX1 R7_reg_5_ ( .D(data_in_1[5]), .E(n992), .CK(clk), .Q(R7[5]) );
  EDFFX1 R7_reg_4_ ( .D(data_in_1[4]), .E(n992), .CK(clk), .Q(R7[4]) );
  EDFFX1 R7_reg_3_ ( .D(data_in_1[3]), .E(n992), .CK(clk), .Q(R7[3]) );
  EDFFX1 R7_reg_2_ ( .D(data_in_1[2]), .E(n992), .CK(clk), .Q(R7[2]) );
  EDFFX1 R7_reg_1_ ( .D(data_in_1[1]), .E(n992), .CK(clk), .Q(R7[1]) );
  EDFFX1 R7_reg_0_ ( .D(data_in_1[0]), .E(n992), .CK(clk), .Q(R7[0]) );
  EDFFX1 R11_reg_33_ ( .D(data_in_1[33]), .E(n1000), .CK(clk), .Q(R11[33]) );
  EDFFX1 R11_reg_32_ ( .D(data_in_1[32]), .E(n1000), .CK(clk), .Q(R11[32]) );
  EDFFX1 R11_reg_31_ ( .D(data_in_1[31]), .E(n1000), .CK(clk), .Q(R11[31]) );
  EDFFX1 R11_reg_30_ ( .D(data_in_1[30]), .E(n1000), .CK(clk), .Q(R11[30]) );
  EDFFX1 R11_reg_29_ ( .D(data_in_1[29]), .E(n1000), .CK(clk), .Q(R11[29]) );
  EDFFX1 R11_reg_28_ ( .D(data_in_1[28]), .E(n1000), .CK(clk), .Q(R11[28]) );
  EDFFX1 R11_reg_27_ ( .D(data_in_1[27]), .E(n1000), .CK(clk), .Q(R11[27]) );
  EDFFX1 R11_reg_26_ ( .D(data_in_1[26]), .E(n1000), .CK(clk), .Q(R11[26]) );
  EDFFX1 R11_reg_25_ ( .D(data_in_1[25]), .E(n1000), .CK(clk), .Q(R11[25]) );
  EDFFX1 R11_reg_24_ ( .D(data_in_1[24]), .E(n1000), .CK(clk), .Q(R11[24]) );
  EDFFX1 R11_reg_23_ ( .D(data_in_1[23]), .E(n1000), .CK(clk), .Q(R11[23]) );
  EDFFX1 R11_reg_22_ ( .D(data_in_1[22]), .E(n1000), .CK(clk), .Q(R11[22]) );
  EDFFX1 R11_reg_21_ ( .D(data_in_1[21]), .E(n1001), .CK(clk), .Q(R11[21]) );
  EDFFX1 R11_reg_20_ ( .D(data_in_1[20]), .E(n1001), .CK(clk), .Q(R11[20]) );
  EDFFX1 R11_reg_19_ ( .D(data_in_1[19]), .E(n1001), .CK(clk), .Q(R11[19]) );
  EDFFX1 R11_reg_18_ ( .D(data_in_1[18]), .E(n1001), .CK(clk), .Q(R11[18]) );
  EDFFX1 R11_reg_17_ ( .D(data_in_1[17]), .E(n1001), .CK(clk), .Q(R11[17]) );
  EDFFX1 R11_reg_16_ ( .D(data_in_1[16]), .E(n1001), .CK(clk), .Q(R11[16]) );
  EDFFX1 R11_reg_15_ ( .D(data_in_1[15]), .E(n1001), .CK(clk), .Q(R11[15]) );
  EDFFX1 R11_reg_14_ ( .D(data_in_1[14]), .E(n1001), .CK(clk), .Q(R11[14]) );
  EDFFX1 R11_reg_13_ ( .D(data_in_1[13]), .E(n1001), .CK(clk), .Q(R11[13]) );
  EDFFX1 R11_reg_12_ ( .D(data_in_1[12]), .E(n1001), .CK(clk), .Q(R11[12]) );
  EDFFX1 R11_reg_11_ ( .D(data_in_1[11]), .E(n1001), .CK(clk), .Q(R11[11]) );
  EDFFX1 R11_reg_10_ ( .D(data_in_1[10]), .E(n1001), .CK(clk), .Q(R11[10]) );
  EDFFX1 R11_reg_9_ ( .D(data_in_1[9]), .E(n1000), .CK(clk), .Q(R11[9]) );
  EDFFX1 R11_reg_8_ ( .D(data_in_1[8]), .E(n1001), .CK(clk), .Q(R11[8]) );
  EDFFX1 R11_reg_7_ ( .D(data_in_1[7]), .E(n1000), .CK(clk), .Q(R11[7]) );
  EDFFX1 R11_reg_6_ ( .D(data_in_1[6]), .E(n1001), .CK(clk), .Q(R11[6]) );
  EDFFX1 R11_reg_5_ ( .D(data_in_1[5]), .E(n1000), .CK(clk), .Q(R11[5]) );
  EDFFX1 R11_reg_4_ ( .D(data_in_1[4]), .E(n1001), .CK(clk), .Q(R11[4]) );
  EDFFX1 R11_reg_3_ ( .D(data_in_1[3]), .E(n1000), .CK(clk), .Q(R11[3]) );
  EDFFX1 R11_reg_2_ ( .D(data_in_1[2]), .E(n1001), .CK(clk), .Q(R11[2]) );
  EDFFX1 R11_reg_1_ ( .D(data_in_1[1]), .E(n1000), .CK(clk), .Q(R11[1]) );
  EDFFX1 R11_reg_0_ ( .D(data_in_1[0]), .E(n1001), .CK(clk), .Q(R11[0]) );
  DFFRHQX1 s_p_flag_out_reg ( .D(n1003), .CK(clk), .RN(rst_n), .Q(s_p_flag_out) );
  EDFFX1 R13_reg_33_ ( .D(data_in_1[33]), .E(n1008), .CK(clk), .Q(R13[33]) );
  EDFFX1 R13_reg_32_ ( .D(data_in_1[32]), .E(n1008), .CK(clk), .Q(R13[32]) );
  EDFFX1 R13_reg_31_ ( .D(data_in_1[31]), .E(n1008), .CK(clk), .Q(R13[31]) );
  EDFFX1 R13_reg_30_ ( .D(data_in_1[30]), .E(n1008), .CK(clk), .Q(R13[30]) );
  EDFFX1 R13_reg_29_ ( .D(data_in_1[29]), .E(n1008), .CK(clk), .Q(R13[29]) );
  EDFFX1 R13_reg_28_ ( .D(data_in_1[28]), .E(n1008), .CK(clk), .Q(R13[28]) );
  EDFFX1 R13_reg_27_ ( .D(data_in_1[27]), .E(n1008), .CK(clk), .Q(R13[27]) );
  EDFFX1 R13_reg_26_ ( .D(data_in_1[26]), .E(n1006), .CK(clk), .Q(R13[26]) );
  EDFFX1 R13_reg_25_ ( .D(data_in_1[25]), .E(n1008), .CK(clk), .Q(R13[25]) );
  EDFFX1 R13_reg_24_ ( .D(data_in_1[24]), .E(n1007), .CK(clk), .Q(R13[24]) );
  EDFFX1 R13_reg_23_ ( .D(data_in_1[23]), .E(n1007), .CK(clk), .Q(R13[23]) );
  EDFFX1 R13_reg_22_ ( .D(data_in_1[22]), .E(n1008), .CK(clk), .Q(R13[22]) );
  EDFFX1 R13_reg_21_ ( .D(data_in_1[21]), .E(n1005), .CK(clk), .Q(R13[21]) );
  EDFFX1 R13_reg_20_ ( .D(data_in_1[20]), .E(n1006), .CK(clk), .Q(R13[20]) );
  EDFFX1 R13_reg_19_ ( .D(data_in_1[19]), .E(n1007), .CK(clk), .Q(R13[19]) );
  EDFFX1 R13_reg_18_ ( .D(data_in_1[18]), .E(n1008), .CK(clk), .Q(R13[18]) );
  EDFFX1 R13_reg_17_ ( .D(data_in_1[17]), .E(n1006), .CK(clk), .Q(R13[17]) );
  EDFFX1 R13_reg_16_ ( .D(data_in_1[16]), .E(n1005), .CK(clk), .Q(R13[16]) );
  EDFFX1 R13_reg_15_ ( .D(data_in_1[15]), .E(n1007), .CK(clk), .Q(R13[15]) );
  EDFFX1 R13_reg_14_ ( .D(data_in_1[14]), .E(n1008), .CK(clk), .Q(R13[14]) );
  EDFFX1 R13_reg_13_ ( .D(data_in_1[13]), .E(n1006), .CK(clk), .Q(R13[13]) );
  EDFFX1 R13_reg_12_ ( .D(data_in_1[12]), .E(n1005), .CK(clk), .Q(R13[12]) );
  EDFFX1 R13_reg_11_ ( .D(data_in_1[11]), .E(n1007), .CK(clk), .Q(R13[11]) );
  EDFFX1 R13_reg_10_ ( .D(data_in_1[10]), .E(n1008), .CK(clk), .Q(R13[10]) );
  EDFFX1 R13_reg_9_ ( .D(data_in_1[9]), .E(n1006), .CK(clk), .Q(R13[9]) );
  EDFFX1 R13_reg_8_ ( .D(data_in_1[8]), .E(n1005), .CK(clk), .Q(R13[8]) );
  EDFFX1 R13_reg_7_ ( .D(data_in_1[7]), .E(n1007), .CK(clk), .Q(R13[7]) );
  EDFFX1 R13_reg_6_ ( .D(data_in_1[6]), .E(n1008), .CK(clk), .Q(R13[6]) );
  EDFFX1 R13_reg_5_ ( .D(data_in_1[5]), .E(n1005), .CK(clk), .Q(R13[5]) );
  EDFFX1 R13_reg_4_ ( .D(data_in_1[4]), .E(n1007), .CK(clk), .Q(R13[4]) );
  EDFFX1 R13_reg_3_ ( .D(data_in_1[3]), .E(n1007), .CK(clk), .Q(R13[3]) );
  EDFFX1 R13_reg_2_ ( .D(data_in_1[2]), .E(n1008), .CK(clk), .Q(R13[2]) );
  EDFFX1 R13_reg_1_ ( .D(data_in_1[1]), .E(n1006), .CK(clk), .Q(R13[1]) );
  EDFFX1 R13_reg_0_ ( .D(data_in_1[0]), .E(n1005), .CK(clk), .Q(R13[0]) );
  EDFFX1 R1_reg_33_ ( .D(data_in_1[33]), .E(n978), .CK(clk), .Q(R1[33]) );
  EDFFX1 R1_reg_32_ ( .D(data_in_1[32]), .E(n978), .CK(clk), .Q(R1[32]) );
  EDFFX1 R1_reg_31_ ( .D(data_in_1[31]), .E(n978), .CK(clk), .Q(R1[31]) );
  EDFFX1 R1_reg_30_ ( .D(data_in_1[30]), .E(n978), .CK(clk), .Q(R1[30]) );
  EDFFX1 R1_reg_29_ ( .D(data_in_1[29]), .E(n978), .CK(clk), .Q(R1[29]) );
  EDFFX1 R1_reg_28_ ( .D(data_in_1[28]), .E(n978), .CK(clk), .Q(R1[28]) );
  EDFFX1 R1_reg_27_ ( .D(data_in_1[27]), .E(n978), .CK(clk), .Q(R1[27]) );
  EDFFX1 R1_reg_26_ ( .D(data_in_1[26]), .E(n978), .CK(clk), .Q(R1[26]) );
  EDFFX1 R1_reg_25_ ( .D(data_in_1[25]), .E(n978), .CK(clk), .Q(R1[25]) );
  EDFFX1 R1_reg_24_ ( .D(data_in_1[24]), .E(n978), .CK(clk), .Q(R1[24]) );
  EDFFX1 R1_reg_23_ ( .D(data_in_1[23]), .E(n978), .CK(clk), .Q(R1[23]) );
  EDFFX1 R1_reg_22_ ( .D(data_in_1[22]), .E(n978), .CK(clk), .Q(R1[22]) );
  EDFFX1 R1_reg_21_ ( .D(data_in_1[21]), .E(n979), .CK(clk), .Q(R1[21]) );
  EDFFX1 R1_reg_20_ ( .D(data_in_1[20]), .E(n979), .CK(clk), .Q(R1[20]) );
  EDFFX1 R1_reg_19_ ( .D(data_in_1[19]), .E(n979), .CK(clk), .Q(R1[19]) );
  EDFFX1 R1_reg_18_ ( .D(data_in_1[18]), .E(n979), .CK(clk), .Q(R1[18]) );
  EDFFX1 R1_reg_17_ ( .D(data_in_1[17]), .E(n979), .CK(clk), .Q(R1[17]) );
  EDFFX1 R1_reg_16_ ( .D(data_in_1[16]), .E(n979), .CK(clk), .Q(R1[16]) );
  EDFFX1 R1_reg_15_ ( .D(data_in_1[15]), .E(n979), .CK(clk), .Q(R1[15]) );
  EDFFX1 R1_reg_14_ ( .D(data_in_1[14]), .E(n979), .CK(clk), .Q(R1[14]) );
  EDFFX1 R1_reg_13_ ( .D(data_in_1[13]), .E(n979), .CK(clk), .Q(R1[13]) );
  EDFFX1 R1_reg_12_ ( .D(data_in_1[12]), .E(n979), .CK(clk), .Q(R1[12]) );
  EDFFX1 R1_reg_11_ ( .D(data_in_1[11]), .E(n979), .CK(clk), .Q(R1[11]) );
  EDFFX1 R1_reg_10_ ( .D(data_in_1[10]), .E(n979), .CK(clk), .Q(R1[10]) );
  EDFFX1 R1_reg_9_ ( .D(data_in_1[9]), .E(n978), .CK(clk), .Q(R1[9]) );
  EDFFX1 R1_reg_8_ ( .D(data_in_1[8]), .E(n979), .CK(clk), .Q(R1[8]) );
  EDFFX1 R1_reg_7_ ( .D(data_in_1[7]), .E(n978), .CK(clk), .Q(R1[7]) );
  EDFFX1 R1_reg_6_ ( .D(data_in_1[6]), .E(n979), .CK(clk), .Q(R1[6]) );
  EDFFX1 R1_reg_5_ ( .D(data_in_1[5]), .E(n978), .CK(clk), .Q(R1[5]) );
  EDFFX1 R1_reg_4_ ( .D(data_in_1[4]), .E(n979), .CK(clk), .Q(R1[4]) );
  EDFFX1 R1_reg_3_ ( .D(data_in_1[3]), .E(n978), .CK(clk), .Q(R1[3]) );
  EDFFX1 R1_reg_2_ ( .D(data_in_1[2]), .E(n979), .CK(clk), .Q(R1[2]) );
  EDFFX1 R1_reg_1_ ( .D(data_in_1[1]), .E(n978), .CK(clk), .Q(R1[1]) );
  EDFFX1 R1_reg_0_ ( .D(data_in_1[0]), .E(n979), .CK(clk), .Q(R1[0]) );
  EDFFX1 R5_reg_33_ ( .D(data_in_1[33]), .E(n988), .CK(clk), .Q(R5[33]) );
  EDFFX1 R5_reg_32_ ( .D(data_in_1[32]), .E(n988), .CK(clk), .Q(R5[32]) );
  EDFFX1 R5_reg_31_ ( .D(data_in_1[31]), .E(n988), .CK(clk), .Q(R5[31]) );
  EDFFX1 R5_reg_30_ ( .D(data_in_1[30]), .E(n988), .CK(clk), .Q(R5[30]) );
  EDFFX1 R5_reg_29_ ( .D(data_in_1[29]), .E(n988), .CK(clk), .Q(R5[29]) );
  EDFFX1 R5_reg_28_ ( .D(data_in_1[28]), .E(n988), .CK(clk), .Q(R5[28]) );
  EDFFX1 R5_reg_27_ ( .D(data_in_1[27]), .E(n988), .CK(clk), .Q(R5[27]) );
  EDFFX1 R5_reg_26_ ( .D(data_in_1[26]), .E(n988), .CK(clk), .Q(R5[26]) );
  EDFFX1 R5_reg_25_ ( .D(data_in_1[25]), .E(n988), .CK(clk), .Q(R5[25]) );
  EDFFX1 R5_reg_24_ ( .D(data_in_1[24]), .E(n988), .CK(clk), .Q(R5[24]) );
  EDFFX1 R5_reg_23_ ( .D(data_in_1[23]), .E(n988), .CK(clk), .Q(R5[23]) );
  EDFFX1 R5_reg_22_ ( .D(data_in_1[22]), .E(n988), .CK(clk), .Q(R5[22]) );
  EDFFX1 R5_reg_21_ ( .D(data_in_1[21]), .E(n989), .CK(clk), .Q(R5[21]) );
  EDFFX1 R5_reg_20_ ( .D(data_in_1[20]), .E(n989), .CK(clk), .Q(R5[20]) );
  EDFFX1 R5_reg_19_ ( .D(data_in_1[19]), .E(n989), .CK(clk), .Q(R5[19]) );
  EDFFX1 R5_reg_18_ ( .D(data_in_1[18]), .E(n989), .CK(clk), .Q(R5[18]) );
  EDFFX1 R5_reg_17_ ( .D(data_in_1[17]), .E(n989), .CK(clk), .Q(R5[17]) );
  EDFFX1 R5_reg_16_ ( .D(data_in_1[16]), .E(n989), .CK(clk), .Q(R5[16]) );
  EDFFX1 R5_reg_15_ ( .D(data_in_1[15]), .E(n989), .CK(clk), .Q(R5[15]) );
  EDFFX1 R5_reg_14_ ( .D(data_in_1[14]), .E(n989), .CK(clk), .Q(R5[14]) );
  EDFFX1 R5_reg_13_ ( .D(data_in_1[13]), .E(n989), .CK(clk), .Q(R5[13]) );
  EDFFX1 R5_reg_12_ ( .D(data_in_1[12]), .E(n989), .CK(clk), .Q(R5[12]) );
  EDFFX1 R5_reg_11_ ( .D(data_in_1[11]), .E(n989), .CK(clk), .Q(R5[11]) );
  EDFFX1 R5_reg_10_ ( .D(data_in_1[10]), .E(n989), .CK(clk), .Q(R5[10]) );
  EDFFX1 R5_reg_9_ ( .D(data_in_1[9]), .E(n988), .CK(clk), .Q(R5[9]) );
  EDFFX1 R5_reg_8_ ( .D(data_in_1[8]), .E(n989), .CK(clk), .Q(R5[8]) );
  EDFFX1 R5_reg_7_ ( .D(data_in_1[7]), .E(n988), .CK(clk), .Q(R5[7]) );
  EDFFX1 R5_reg_6_ ( .D(data_in_1[6]), .E(n989), .CK(clk), .Q(R5[6]) );
  EDFFX1 R5_reg_5_ ( .D(data_in_1[5]), .E(n988), .CK(clk), .Q(R5[5]) );
  EDFFX1 R5_reg_4_ ( .D(data_in_1[4]), .E(n989), .CK(clk), .Q(R5[4]) );
  EDFFX1 R5_reg_3_ ( .D(data_in_1[3]), .E(n988), .CK(clk), .Q(R5[3]) );
  EDFFX1 R5_reg_2_ ( .D(data_in_1[2]), .E(n989), .CK(clk), .Q(R5[2]) );
  EDFFX1 R5_reg_1_ ( .D(data_in_1[1]), .E(n988), .CK(clk), .Q(R5[1]) );
  EDFFX1 R5_reg_0_ ( .D(data_in_1[0]), .E(n989), .CK(clk), .Q(R5[0]) );
  EDFFX1 R9_reg_33_ ( .D(data_in_1[33]), .E(n996), .CK(clk), .Q(R9[33]) );
  EDFFX1 R9_reg_32_ ( .D(data_in_1[32]), .E(n996), .CK(clk), .Q(R9[32]) );
  EDFFX1 R9_reg_31_ ( .D(data_in_1[31]), .E(n996), .CK(clk), .Q(R9[31]) );
  EDFFX1 R9_reg_30_ ( .D(data_in_1[30]), .E(n996), .CK(clk), .Q(R9[30]) );
  EDFFX1 R9_reg_29_ ( .D(data_in_1[29]), .E(n996), .CK(clk), .Q(R9[29]) );
  EDFFX1 R9_reg_28_ ( .D(data_in_1[28]), .E(n996), .CK(clk), .Q(R9[28]) );
  EDFFX1 R9_reg_27_ ( .D(data_in_1[27]), .E(n996), .CK(clk), .Q(R9[27]) );
  EDFFX1 R9_reg_26_ ( .D(data_in_1[26]), .E(n996), .CK(clk), .Q(R9[26]) );
  EDFFX1 R9_reg_25_ ( .D(data_in_1[25]), .E(n996), .CK(clk), .Q(R9[25]) );
  EDFFX1 R9_reg_24_ ( .D(data_in_1[24]), .E(n996), .CK(clk), .Q(R9[24]) );
  EDFFX1 R9_reg_23_ ( .D(data_in_1[23]), .E(n996), .CK(clk), .Q(R9[23]) );
  EDFFX1 R9_reg_22_ ( .D(data_in_1[22]), .E(n996), .CK(clk), .Q(R9[22]) );
  EDFFX1 R9_reg_21_ ( .D(data_in_1[21]), .E(n997), .CK(clk), .Q(R9[21]) );
  EDFFX1 R9_reg_20_ ( .D(data_in_1[20]), .E(n997), .CK(clk), .Q(R9[20]) );
  EDFFX1 R9_reg_19_ ( .D(data_in_1[19]), .E(n997), .CK(clk), .Q(R9[19]) );
  EDFFX1 R9_reg_18_ ( .D(data_in_1[18]), .E(n997), .CK(clk), .Q(R9[18]) );
  EDFFX1 R9_reg_17_ ( .D(data_in_1[17]), .E(n997), .CK(clk), .Q(R9[17]) );
  EDFFX1 R9_reg_16_ ( .D(data_in_1[16]), .E(n997), .CK(clk), .Q(R9[16]) );
  EDFFX1 R9_reg_15_ ( .D(data_in_1[15]), .E(n997), .CK(clk), .Q(R9[15]) );
  EDFFX1 R9_reg_14_ ( .D(data_in_1[14]), .E(n997), .CK(clk), .Q(R9[14]) );
  EDFFX1 R9_reg_13_ ( .D(data_in_1[13]), .E(n997), .CK(clk), .Q(R9[13]) );
  EDFFX1 R9_reg_12_ ( .D(data_in_1[12]), .E(n997), .CK(clk), .Q(R9[12]) );
  EDFFX1 R9_reg_11_ ( .D(data_in_1[11]), .E(n997), .CK(clk), .Q(R9[11]) );
  EDFFX1 R9_reg_10_ ( .D(data_in_1[10]), .E(n997), .CK(clk), .Q(R9[10]) );
  EDFFX1 R9_reg_9_ ( .D(data_in_1[9]), .E(n996), .CK(clk), .Q(R9[9]) );
  EDFFX1 R9_reg_8_ ( .D(data_in_1[8]), .E(n997), .CK(clk), .Q(R9[8]) );
  EDFFX1 R9_reg_7_ ( .D(data_in_1[7]), .E(n996), .CK(clk), .Q(R9[7]) );
  EDFFX1 R9_reg_6_ ( .D(data_in_1[6]), .E(n997), .CK(clk), .Q(R9[6]) );
  EDFFX1 R9_reg_5_ ( .D(data_in_1[5]), .E(n996), .CK(clk), .Q(R9[5]) );
  EDFFX1 R9_reg_4_ ( .D(data_in_1[4]), .E(n997), .CK(clk), .Q(R9[4]) );
  EDFFX1 R9_reg_3_ ( .D(data_in_1[3]), .E(n996), .CK(clk), .Q(R9[3]) );
  EDFFX1 R9_reg_2_ ( .D(data_in_1[2]), .E(n997), .CK(clk), .Q(R9[2]) );
  EDFFX1 R9_reg_1_ ( .D(data_in_1[1]), .E(n996), .CK(clk), .Q(R9[1]) );
  EDFFX1 R9_reg_0_ ( .D(data_in_1[0]), .E(n997), .CK(clk), .Q(R9[0]) );
  EDFFX1 R14_reg_33_ ( .D(data_in_1[33]), .E(n1010), .CK(clk), .Q(R14[33]) );
  EDFFX1 R14_reg_32_ ( .D(data_in_1[32]), .E(n1011), .CK(clk), .Q(R14[32]) );
  EDFFX1 R14_reg_31_ ( .D(data_in_1[31]), .E(n1013), .CK(clk), .Q(R14[31]) );
  EDFFX1 R14_reg_30_ ( .D(data_in_1[30]), .E(n1012), .CK(clk), .Q(R14[30]) );
  EDFFX1 R14_reg_29_ ( .D(data_in_1[29]), .E(n1012), .CK(clk), .Q(R14[29]) );
  EDFFX1 R14_reg_28_ ( .D(data_in_1[28]), .E(n1011), .CK(clk), .Q(R14[28]) );
  EDFFX1 R14_reg_27_ ( .D(data_in_1[27]), .E(n1013), .CK(clk), .Q(R14[27]) );
  EDFFX1 R14_reg_26_ ( .D(data_in_1[26]), .E(n1012), .CK(clk), .Q(R14[26]) );
  EDFFX1 R14_reg_25_ ( .D(data_in_1[25]), .E(n1010), .CK(clk), .Q(R14[25]) );
  EDFFX1 R14_reg_24_ ( .D(data_in_1[24]), .E(n1013), .CK(clk), .Q(R14[24]) );
  EDFFX1 R14_reg_23_ ( .D(data_in_1[23]), .E(n1011), .CK(clk), .Q(R14[23]) );
  EDFFX1 R14_reg_22_ ( .D(data_in_1[22]), .E(n1011), .CK(clk), .Q(R14[22]) );
  EDFFX1 R14_reg_21_ ( .D(data_in_1[21]), .E(n1012), .CK(clk), .Q(R14[21]) );
  EDFFX1 R14_reg_20_ ( .D(data_in_1[20]), .E(n1013), .CK(clk), .Q(R14[20]) );
  EDFFX1 R14_reg_19_ ( .D(data_in_1[19]), .E(n1010), .CK(clk), .Q(R14[19]) );
  EDFFX1 R14_reg_18_ ( .D(data_in_1[18]), .E(n1010), .CK(clk), .Q(R14[18]) );
  EDFFX1 R14_reg_17_ ( .D(data_in_1[17]), .E(n1010), .CK(clk), .Q(R14[17]) );
  EDFFX1 R14_reg_16_ ( .D(data_in_1[16]), .E(n1010), .CK(clk), .Q(R14[16]) );
  EDFFX1 R14_reg_15_ ( .D(data_in_1[15]), .E(n1010), .CK(clk), .Q(R14[15]) );
  EDFFX1 R14_reg_14_ ( .D(data_in_1[14]), .E(n1010), .CK(clk), .Q(R14[14]) );
  EDFFX1 R14_reg_13_ ( .D(data_in_1[13]), .E(n1010), .CK(clk), .Q(R14[13]) );
  EDFFX1 R14_reg_12_ ( .D(data_in_1[12]), .E(n1010), .CK(clk), .Q(R14[12]) );
  EDFFX1 R14_reg_11_ ( .D(data_in_1[11]), .E(n1010), .CK(clk), .Q(R14[11]) );
  EDFFX1 R14_reg_10_ ( .D(data_in_1[10]), .E(n1010), .CK(clk), .Q(R14[10]) );
  EDFFX1 R14_reg_9_ ( .D(data_in_1[9]), .E(n1010), .CK(clk), .Q(R14[9]) );
  EDFFX1 R14_reg_8_ ( .D(data_in_1[8]), .E(n1010), .CK(clk), .Q(R14[8]) );
  EDFFX1 R14_reg_7_ ( .D(data_in_1[7]), .E(n1010), .CK(clk), .Q(R14[7]) );
  EDFFX1 R14_reg_6_ ( .D(data_in_1[6]), .E(n1010), .CK(clk), .Q(R14[6]) );
  EDFFX1 R14_reg_5_ ( .D(data_in_1[5]), .E(n1010), .CK(clk), .Q(R14[5]) );
  EDFFX1 R14_reg_4_ ( .D(data_in_1[4]), .E(n1010), .CK(clk), .Q(R14[4]) );
  EDFFX1 R14_reg_3_ ( .D(data_in_1[3]), .E(n1010), .CK(clk), .Q(R14[3]) );
  EDFFX1 R14_reg_2_ ( .D(data_in_1[2]), .E(n1010), .CK(clk), .Q(R14[2]) );
  EDFFX1 R14_reg_1_ ( .D(data_in_1[1]), .E(n1010), .CK(clk), .Q(R14[1]) );
  EDFFX1 R14_reg_0_ ( .D(data_in_1[0]), .E(n1010), .CK(clk), .Q(R14[0]) );
  EDFFX1 R2_reg_33_ ( .D(data_in_1[33]), .E(n981), .CK(clk), .Q(R2[33]) );
  EDFFX1 R2_reg_32_ ( .D(data_in_1[32]), .E(n981), .CK(clk), .Q(R2[32]) );
  EDFFX1 R2_reg_31_ ( .D(data_in_1[31]), .E(n981), .CK(clk), .Q(R2[31]) );
  EDFFX1 R2_reg_30_ ( .D(data_in_1[30]), .E(n981), .CK(clk), .Q(R2[30]) );
  EDFFX1 R2_reg_29_ ( .D(data_in_1[29]), .E(n981), .CK(clk), .Q(R2[29]) );
  EDFFX1 R2_reg_28_ ( .D(data_in_1[28]), .E(n981), .CK(clk), .Q(R2[28]) );
  EDFFX1 R2_reg_27_ ( .D(data_in_1[27]), .E(n981), .CK(clk), .Q(R2[27]) );
  EDFFX1 R2_reg_26_ ( .D(data_in_1[26]), .E(n981), .CK(clk), .Q(R2[26]) );
  EDFFX1 R2_reg_25_ ( .D(data_in_1[25]), .E(n981), .CK(clk), .Q(R2[25]) );
  EDFFX1 R2_reg_24_ ( .D(data_in_1[24]), .E(n981), .CK(clk), .Q(R2[24]) );
  EDFFX1 R2_reg_23_ ( .D(data_in_1[23]), .E(n981), .CK(clk), .Q(R2[23]) );
  EDFFX1 R2_reg_22_ ( .D(data_in_1[22]), .E(n981), .CK(clk), .Q(R2[22]) );
  EDFFX1 R2_reg_21_ ( .D(data_in_1[21]), .E(n982), .CK(clk), .Q(R2[21]) );
  EDFFX1 R2_reg_20_ ( .D(data_in_1[20]), .E(n982), .CK(clk), .Q(R2[20]) );
  EDFFX1 R2_reg_19_ ( .D(data_in_1[19]), .E(n982), .CK(clk), .Q(R2[19]) );
  EDFFX1 R2_reg_18_ ( .D(data_in_1[18]), .E(n982), .CK(clk), .Q(R2[18]) );
  EDFFX1 R2_reg_17_ ( .D(data_in_1[17]), .E(n982), .CK(clk), .Q(R2[17]) );
  EDFFX1 R2_reg_16_ ( .D(data_in_1[16]), .E(n982), .CK(clk), .Q(R2[16]) );
  EDFFX1 R2_reg_15_ ( .D(data_in_1[15]), .E(n982), .CK(clk), .Q(R2[15]) );
  EDFFX1 R2_reg_14_ ( .D(data_in_1[14]), .E(n982), .CK(clk), .Q(R2[14]) );
  EDFFX1 R2_reg_13_ ( .D(data_in_1[13]), .E(n982), .CK(clk), .Q(R2[13]) );
  EDFFX1 R2_reg_12_ ( .D(data_in_1[12]), .E(n982), .CK(clk), .Q(R2[12]) );
  EDFFX1 R2_reg_11_ ( .D(data_in_1[11]), .E(n982), .CK(clk), .Q(R2[11]) );
  EDFFX1 R2_reg_10_ ( .D(data_in_1[10]), .E(n982), .CK(clk), .Q(R2[10]) );
  EDFFX1 R2_reg_9_ ( .D(data_in_1[9]), .E(n980), .CK(clk), .Q(R2[9]) );
  EDFFX1 R2_reg_8_ ( .D(data_in_1[8]), .E(n980), .CK(clk), .Q(R2[8]) );
  EDFFX1 R2_reg_7_ ( .D(data_in_1[7]), .E(n980), .CK(clk), .Q(R2[7]) );
  EDFFX1 R2_reg_6_ ( .D(data_in_1[6]), .E(n980), .CK(clk), .Q(R2[6]) );
  EDFFX1 R2_reg_5_ ( .D(data_in_1[5]), .E(n980), .CK(clk), .Q(R2[5]) );
  EDFFX1 R2_reg_4_ ( .D(data_in_1[4]), .E(n980), .CK(clk), .Q(R2[4]) );
  EDFFX1 R2_reg_3_ ( .D(data_in_1[3]), .E(n981), .CK(clk), .Q(R2[3]) );
  EDFFX1 R2_reg_2_ ( .D(data_in_1[2]), .E(n982), .CK(clk), .Q(R2[2]) );
  EDFFX1 R2_reg_1_ ( .D(data_in_1[1]), .E(n981), .CK(clk), .Q(R2[1]) );
  EDFFX1 R2_reg_0_ ( .D(data_in_1[0]), .E(n982), .CK(clk), .Q(R2[0]) );
  EDFFX1 R6_reg_33_ ( .D(data_in_1[33]), .E(n990), .CK(clk), .Q(R6[33]) );
  EDFFX1 R6_reg_32_ ( .D(data_in_1[32]), .E(n990), .CK(clk), .Q(R6[32]) );
  EDFFX1 R6_reg_31_ ( .D(data_in_1[31]), .E(n990), .CK(clk), .Q(R6[31]) );
  EDFFX1 R6_reg_30_ ( .D(data_in_1[30]), .E(n990), .CK(clk), .Q(R6[30]) );
  EDFFX1 R6_reg_29_ ( .D(data_in_1[29]), .E(n990), .CK(clk), .Q(R6[29]) );
  EDFFX1 R6_reg_28_ ( .D(data_in_1[28]), .E(n990), .CK(clk), .Q(R6[28]) );
  EDFFX1 R6_reg_27_ ( .D(data_in_1[27]), .E(n990), .CK(clk), .Q(R6[27]) );
  EDFFX1 R6_reg_26_ ( .D(data_in_1[26]), .E(n990), .CK(clk), .Q(R6[26]) );
  EDFFX1 R6_reg_25_ ( .D(data_in_1[25]), .E(n990), .CK(clk), .Q(R6[25]) );
  EDFFX1 R6_reg_24_ ( .D(data_in_1[24]), .E(n990), .CK(clk), .Q(R6[24]) );
  EDFFX1 R6_reg_23_ ( .D(data_in_1[23]), .E(n990), .CK(clk), .Q(R6[23]) );
  EDFFX1 R6_reg_22_ ( .D(data_in_1[22]), .E(n990), .CK(clk), .Q(R6[22]) );
  EDFFX1 R6_reg_21_ ( .D(data_in_1[21]), .E(n991), .CK(clk), .Q(R6[21]) );
  EDFFX1 R6_reg_20_ ( .D(data_in_1[20]), .E(n991), .CK(clk), .Q(R6[20]) );
  EDFFX1 R6_reg_19_ ( .D(data_in_1[19]), .E(n991), .CK(clk), .Q(R6[19]) );
  EDFFX1 R6_reg_18_ ( .D(data_in_1[18]), .E(n991), .CK(clk), .Q(R6[18]) );
  EDFFX1 R6_reg_17_ ( .D(data_in_1[17]), .E(n991), .CK(clk), .Q(R6[17]) );
  EDFFX1 R6_reg_16_ ( .D(data_in_1[16]), .E(n991), .CK(clk), .Q(R6[16]) );
  EDFFX1 R6_reg_15_ ( .D(data_in_1[15]), .E(n991), .CK(clk), .Q(R6[15]) );
  EDFFX1 R6_reg_14_ ( .D(data_in_1[14]), .E(n991), .CK(clk), .Q(R6[14]) );
  EDFFX1 R6_reg_13_ ( .D(data_in_1[13]), .E(n991), .CK(clk), .Q(R6[13]) );
  EDFFX1 R6_reg_12_ ( .D(data_in_1[12]), .E(n991), .CK(clk), .Q(R6[12]) );
  EDFFX1 R6_reg_11_ ( .D(data_in_1[11]), .E(n991), .CK(clk), .Q(R6[11]) );
  EDFFX1 R6_reg_10_ ( .D(data_in_1[10]), .E(n991), .CK(clk), .Q(R6[10]) );
  EDFFX1 R6_reg_9_ ( .D(data_in_1[9]), .E(n990), .CK(clk), .Q(R6[9]) );
  EDFFX1 R6_reg_8_ ( .D(data_in_1[8]), .E(n991), .CK(clk), .Q(R6[8]) );
  EDFFX1 R6_reg_7_ ( .D(data_in_1[7]), .E(n990), .CK(clk), .Q(R6[7]) );
  EDFFX1 R6_reg_6_ ( .D(data_in_1[6]), .E(n991), .CK(clk), .Q(R6[6]) );
  EDFFX1 R6_reg_5_ ( .D(data_in_1[5]), .E(n990), .CK(clk), .Q(R6[5]) );
  EDFFX1 R6_reg_4_ ( .D(data_in_1[4]), .E(n991), .CK(clk), .Q(R6[4]) );
  EDFFX1 R6_reg_3_ ( .D(data_in_1[3]), .E(n990), .CK(clk), .Q(R6[3]) );
  EDFFX1 R6_reg_2_ ( .D(data_in_1[2]), .E(n991), .CK(clk), .Q(R6[2]) );
  EDFFX1 R6_reg_1_ ( .D(data_in_1[1]), .E(n990), .CK(clk), .Q(R6[1]) );
  EDFFX1 R6_reg_0_ ( .D(data_in_1[0]), .E(n991), .CK(clk), .Q(R6[0]) );
  EDFFX1 R10_reg_33_ ( .D(data_in_1[33]), .E(n998), .CK(clk), .Q(R10[33]) );
  EDFFX1 R10_reg_32_ ( .D(data_in_1[32]), .E(n998), .CK(clk), .Q(R10[32]) );
  EDFFX1 R10_reg_31_ ( .D(data_in_1[31]), .E(n998), .CK(clk), .Q(R10[31]) );
  EDFFX1 R10_reg_30_ ( .D(data_in_1[30]), .E(n998), .CK(clk), .Q(R10[30]) );
  EDFFX1 R10_reg_29_ ( .D(data_in_1[29]), .E(n998), .CK(clk), .Q(R10[29]) );
  EDFFX1 R10_reg_28_ ( .D(data_in_1[28]), .E(n998), .CK(clk), .Q(R10[28]) );
  EDFFX1 R10_reg_27_ ( .D(data_in_1[27]), .E(n998), .CK(clk), .Q(R10[27]) );
  EDFFX1 R10_reg_26_ ( .D(data_in_1[26]), .E(n998), .CK(clk), .Q(R10[26]) );
  EDFFX1 R10_reg_25_ ( .D(data_in_1[25]), .E(n998), .CK(clk), .Q(R10[25]) );
  EDFFX1 R10_reg_24_ ( .D(data_in_1[24]), .E(n998), .CK(clk), .Q(R10[24]) );
  EDFFX1 R10_reg_23_ ( .D(data_in_1[23]), .E(n998), .CK(clk), .Q(R10[23]) );
  EDFFX1 R10_reg_22_ ( .D(data_in_1[22]), .E(n998), .CK(clk), .Q(R10[22]) );
  EDFFX1 R10_reg_21_ ( .D(data_in_1[21]), .E(n999), .CK(clk), .Q(R10[21]) );
  EDFFX1 R10_reg_20_ ( .D(data_in_1[20]), .E(n999), .CK(clk), .Q(R10[20]) );
  EDFFX1 R10_reg_19_ ( .D(data_in_1[19]), .E(n999), .CK(clk), .Q(R10[19]) );
  EDFFX1 R10_reg_18_ ( .D(data_in_1[18]), .E(n999), .CK(clk), .Q(R10[18]) );
  EDFFX1 R10_reg_17_ ( .D(data_in_1[17]), .E(n999), .CK(clk), .Q(R10[17]) );
  EDFFX1 R10_reg_16_ ( .D(data_in_1[16]), .E(n999), .CK(clk), .Q(R10[16]) );
  EDFFX1 R10_reg_15_ ( .D(data_in_1[15]), .E(n999), .CK(clk), .Q(R10[15]) );
  EDFFX1 R10_reg_14_ ( .D(data_in_1[14]), .E(n999), .CK(clk), .Q(R10[14]) );
  EDFFX1 R10_reg_13_ ( .D(data_in_1[13]), .E(n999), .CK(clk), .Q(R10[13]) );
  EDFFX1 R10_reg_12_ ( .D(data_in_1[12]), .E(n999), .CK(clk), .Q(R10[12]) );
  EDFFX1 R10_reg_11_ ( .D(data_in_1[11]), .E(n999), .CK(clk), .Q(R10[11]) );
  EDFFX1 R10_reg_10_ ( .D(data_in_1[10]), .E(n999), .CK(clk), .Q(R10[10]) );
  EDFFX1 R10_reg_9_ ( .D(data_in_1[9]), .E(n998), .CK(clk), .Q(R10[9]) );
  EDFFX1 R10_reg_8_ ( .D(data_in_1[8]), .E(n999), .CK(clk), .Q(R10[8]) );
  EDFFX1 R10_reg_7_ ( .D(data_in_1[7]), .E(n998), .CK(clk), .Q(R10[7]) );
  EDFFX1 R10_reg_6_ ( .D(data_in_1[6]), .E(n999), .CK(clk), .Q(R10[6]) );
  EDFFX1 R10_reg_5_ ( .D(data_in_1[5]), .E(n998), .CK(clk), .Q(R10[5]) );
  EDFFX1 R10_reg_4_ ( .D(data_in_1[4]), .E(n999), .CK(clk), .Q(R10[4]) );
  EDFFX1 R10_reg_3_ ( .D(data_in_1[3]), .E(n998), .CK(clk), .Q(R10[3]) );
  EDFFX1 R10_reg_2_ ( .D(data_in_1[2]), .E(n999), .CK(clk), .Q(R10[2]) );
  EDFFX1 R10_reg_1_ ( .D(data_in_1[1]), .E(n998), .CK(clk), .Q(R10[1]) );
  EDFFX1 R10_reg_0_ ( .D(data_in_1[0]), .E(n999), .CK(clk), .Q(R10[0]) );
  EDFFX1 R0_reg_33_ ( .D(data_in_1[33]), .E(n1042), .CK(clk), .Q(R0[33]) );
  EDFFX1 R0_reg_32_ ( .D(data_in_1[32]), .E(n1042), .CK(clk), .Q(R0[32]) );
  EDFFX1 R0_reg_31_ ( .D(data_in_1[31]), .E(n1042), .CK(clk), .Q(R0[31]) );
  EDFFX1 R0_reg_30_ ( .D(data_in_1[30]), .E(n1042), .CK(clk), .Q(R0[30]) );
  EDFFX1 R0_reg_29_ ( .D(data_in_1[29]), .E(n1042), .CK(clk), .Q(R0[29]) );
  EDFFX1 R0_reg_28_ ( .D(data_in_1[28]), .E(n1042), .CK(clk), .Q(R0[28]) );
  EDFFX1 R0_reg_27_ ( .D(data_in_1[27]), .E(n1042), .CK(clk), .Q(R0[27]) );
  EDFFX1 R0_reg_26_ ( .D(data_in_1[26]), .E(n1042), .CK(clk), .Q(R0[26]) );
  EDFFX1 R0_reg_25_ ( .D(data_in_1[25]), .E(n1042), .CK(clk), .Q(R0[25]) );
  EDFFX1 R0_reg_24_ ( .D(data_in_1[24]), .E(n1042), .CK(clk), .Q(R0[24]) );
  EDFFX1 R0_reg_23_ ( .D(data_in_1[23]), .E(n1040), .CK(clk), .Q(R0[23]) );
  EDFFX1 R0_reg_22_ ( .D(data_in_1[22]), .E(n1036), .CK(clk), .Q(R0[22]) );
  EDFFX1 R0_reg_21_ ( .D(data_in_1[21]), .E(n1039), .CK(clk), .Q(R0[21]) );
  EDFFX1 R0_reg_20_ ( .D(data_in_1[20]), .E(n1033), .CK(clk), .Q(R0[20]) );
  EDFFX1 R0_reg_19_ ( .D(data_in_1[19]), .E(n1034), .CK(clk), .Q(R0[19]) );
  EDFFX1 R0_reg_18_ ( .D(data_in_1[18]), .E(n1035), .CK(clk), .Q(R0[18]) );
  EDFFX1 R0_reg_17_ ( .D(data_in_1[17]), .E(n1037), .CK(clk), .Q(R0[17]) );
  EDFFX1 R0_reg_16_ ( .D(data_in_1[16]), .E(n1038), .CK(clk), .Q(R0[16]) );
  EDFFX1 R0_reg_15_ ( .D(data_in_1[15]), .E(n1041), .CK(clk), .Q(R0[15]) );
  EDFFX1 R0_reg_14_ ( .D(data_in_1[14]), .E(n1040), .CK(clk), .Q(R0[14]) );
  EDFFX1 R0_reg_13_ ( .D(data_in_1[13]), .E(n1036), .CK(clk), .Q(R0[13]) );
  EDFFX1 R0_reg_12_ ( .D(data_in_1[12]), .E(n1039), .CK(clk), .Q(R0[12]) );
  EDFFX1 R0_reg_11_ ( .D(data_in_1[11]), .E(n1033), .CK(clk), .Q(R0[11]) );
  EDFFX1 R0_reg_10_ ( .D(data_in_1[10]), .E(n1034), .CK(clk), .Q(R0[10]) );
  EDFFX1 R0_reg_9_ ( .D(data_in_1[9]), .E(n1035), .CK(clk), .Q(R0[9]) );
  EDFFX1 R0_reg_8_ ( .D(data_in_1[8]), .E(n1037), .CK(clk), .Q(R0[8]) );
  EDFFX1 R0_reg_7_ ( .D(data_in_1[7]), .E(n1038), .CK(clk), .Q(R0[7]) );
  EDFFX1 R0_reg_6_ ( .D(data_in_1[6]), .E(n1041), .CK(clk), .Q(R0[6]) );
  EDFFX1 R0_reg_5_ ( .D(data_in_1[5]), .E(n1040), .CK(clk), .Q(R0[5]) );
  EDFFX1 R0_reg_4_ ( .D(data_in_1[4]), .E(n1036), .CK(clk), .Q(R0[4]) );
  EDFFX1 R0_reg_3_ ( .D(data_in_1[3]), .E(n1039), .CK(clk), .Q(R0[3]) );
  EDFFX1 R0_reg_2_ ( .D(data_in_1[2]), .E(n1040), .CK(clk), .Q(R0[2]) );
  EDFFX1 R0_reg_1_ ( .D(data_in_1[1]), .E(n1036), .CK(clk), .Q(R0[1]) );
  EDFFX1 R0_reg_0_ ( .D(data_in_1[0]), .E(n1039), .CK(clk), .Q(R0[0]) );
  EDFFX1 R4_reg_33_ ( .D(data_in_1[33]), .E(n986), .CK(clk), .Q(R4[33]) );
  EDFFX1 R4_reg_32_ ( .D(data_in_1[32]), .E(n986), .CK(clk), .Q(R4[32]) );
  EDFFX1 R4_reg_31_ ( .D(data_in_1[31]), .E(n986), .CK(clk), .Q(R4[31]) );
  EDFFX1 R4_reg_30_ ( .D(data_in_1[30]), .E(n986), .CK(clk), .Q(R4[30]) );
  EDFFX1 R4_reg_29_ ( .D(data_in_1[29]), .E(n986), .CK(clk), .Q(R4[29]) );
  EDFFX1 R4_reg_28_ ( .D(data_in_1[28]), .E(n986), .CK(clk), .Q(R4[28]) );
  EDFFX1 R4_reg_27_ ( .D(data_in_1[27]), .E(n986), .CK(clk), .Q(R4[27]) );
  EDFFX1 R4_reg_26_ ( .D(data_in_1[26]), .E(n986), .CK(clk), .Q(R4[26]) );
  EDFFX1 R4_reg_25_ ( .D(data_in_1[25]), .E(n986), .CK(clk), .Q(R4[25]) );
  EDFFX1 R4_reg_24_ ( .D(data_in_1[24]), .E(n986), .CK(clk), .Q(R4[24]) );
  EDFFX1 R4_reg_23_ ( .D(data_in_1[23]), .E(n986), .CK(clk), .Q(R4[23]) );
  EDFFX1 R4_reg_22_ ( .D(data_in_1[22]), .E(n986), .CK(clk), .Q(R4[22]) );
  EDFFX1 R4_reg_21_ ( .D(data_in_1[21]), .E(n987), .CK(clk), .Q(R4[21]) );
  EDFFX1 R4_reg_20_ ( .D(data_in_1[20]), .E(n987), .CK(clk), .Q(R4[20]) );
  EDFFX1 R4_reg_19_ ( .D(data_in_1[19]), .E(n987), .CK(clk), .Q(R4[19]) );
  EDFFX1 R4_reg_18_ ( .D(data_in_1[18]), .E(n987), .CK(clk), .Q(R4[18]) );
  EDFFX1 R4_reg_17_ ( .D(data_in_1[17]), .E(n987), .CK(clk), .Q(R4[17]) );
  EDFFX1 R4_reg_16_ ( .D(data_in_1[16]), .E(n987), .CK(clk), .Q(R4[16]) );
  EDFFX1 R4_reg_15_ ( .D(data_in_1[15]), .E(n987), .CK(clk), .Q(R4[15]) );
  EDFFX1 R4_reg_14_ ( .D(data_in_1[14]), .E(n987), .CK(clk), .Q(R4[14]) );
  EDFFX1 R4_reg_13_ ( .D(data_in_1[13]), .E(n987), .CK(clk), .Q(R4[13]) );
  EDFFX1 R4_reg_12_ ( .D(data_in_1[12]), .E(n987), .CK(clk), .Q(R4[12]) );
  EDFFX1 R4_reg_11_ ( .D(data_in_1[11]), .E(n987), .CK(clk), .Q(R4[11]) );
  EDFFX1 R4_reg_10_ ( .D(data_in_1[10]), .E(n987), .CK(clk), .Q(R4[10]) );
  EDFFX1 R4_reg_9_ ( .D(data_in_1[9]), .E(n986), .CK(clk), .Q(R4[9]) );
  EDFFX1 R4_reg_8_ ( .D(data_in_1[8]), .E(n987), .CK(clk), .Q(R4[8]) );
  EDFFX1 R4_reg_7_ ( .D(data_in_1[7]), .E(n986), .CK(clk), .Q(R4[7]) );
  EDFFX1 R4_reg_6_ ( .D(data_in_1[6]), .E(n987), .CK(clk), .Q(R4[6]) );
  EDFFX1 R4_reg_5_ ( .D(data_in_1[5]), .E(n986), .CK(clk), .Q(R4[5]) );
  EDFFX1 R4_reg_4_ ( .D(data_in_1[4]), .E(n987), .CK(clk), .Q(R4[4]) );
  EDFFX1 R4_reg_3_ ( .D(data_in_1[3]), .E(n986), .CK(clk), .Q(R4[3]) );
  EDFFX1 R4_reg_2_ ( .D(data_in_1[2]), .E(n987), .CK(clk), .Q(R4[2]) );
  EDFFX1 R4_reg_1_ ( .D(data_in_1[1]), .E(n986), .CK(clk), .Q(R4[1]) );
  EDFFX1 R4_reg_0_ ( .D(data_in_1[0]), .E(n987), .CK(clk), .Q(R4[0]) );
  EDFFX1 R8_reg_33_ ( .D(data_in_1[33]), .E(n994), .CK(clk), .Q(R8[33]) );
  EDFFX1 R8_reg_32_ ( .D(data_in_1[32]), .E(n994), .CK(clk), .Q(R8[32]) );
  EDFFX1 R8_reg_31_ ( .D(data_in_1[31]), .E(n994), .CK(clk), .Q(R8[31]) );
  EDFFX1 R8_reg_30_ ( .D(data_in_1[30]), .E(n994), .CK(clk), .Q(R8[30]) );
  EDFFX1 R8_reg_29_ ( .D(data_in_1[29]), .E(n994), .CK(clk), .Q(R8[29]) );
  EDFFX1 R8_reg_28_ ( .D(data_in_1[28]), .E(n994), .CK(clk), .Q(R8[28]) );
  EDFFX1 R8_reg_27_ ( .D(data_in_1[27]), .E(n994), .CK(clk), .Q(R8[27]) );
  EDFFX1 R8_reg_26_ ( .D(data_in_1[26]), .E(n994), .CK(clk), .Q(R8[26]) );
  EDFFX1 R8_reg_25_ ( .D(data_in_1[25]), .E(n994), .CK(clk), .Q(R8[25]) );
  EDFFX1 R8_reg_24_ ( .D(data_in_1[24]), .E(n994), .CK(clk), .Q(R8[24]) );
  EDFFX1 R8_reg_23_ ( .D(data_in_1[23]), .E(n994), .CK(clk), .Q(R8[23]) );
  EDFFX1 R8_reg_22_ ( .D(data_in_1[22]), .E(n994), .CK(clk), .Q(R8[22]) );
  EDFFX1 R8_reg_21_ ( .D(data_in_1[21]), .E(n995), .CK(clk), .Q(R8[21]) );
  EDFFX1 R8_reg_20_ ( .D(data_in_1[20]), .E(n995), .CK(clk), .Q(R8[20]) );
  EDFFX1 R8_reg_19_ ( .D(data_in_1[19]), .E(n995), .CK(clk), .Q(R8[19]) );
  EDFFX1 R8_reg_18_ ( .D(data_in_1[18]), .E(n995), .CK(clk), .Q(R8[18]) );
  EDFFX1 R8_reg_17_ ( .D(data_in_1[17]), .E(n995), .CK(clk), .Q(R8[17]) );
  EDFFX1 R8_reg_16_ ( .D(data_in_1[16]), .E(n995), .CK(clk), .Q(R8[16]) );
  EDFFX1 R8_reg_15_ ( .D(data_in_1[15]), .E(n995), .CK(clk), .Q(R8[15]) );
  EDFFX1 R8_reg_14_ ( .D(data_in_1[14]), .E(n995), .CK(clk), .Q(R8[14]) );
  EDFFX1 R8_reg_13_ ( .D(data_in_1[13]), .E(n995), .CK(clk), .Q(R8[13]) );
  EDFFX1 R8_reg_12_ ( .D(data_in_1[12]), .E(n995), .CK(clk), .Q(R8[12]) );
  EDFFX1 R8_reg_11_ ( .D(data_in_1[11]), .E(n995), .CK(clk), .Q(R8[11]) );
  EDFFX1 R8_reg_10_ ( .D(data_in_1[10]), .E(n995), .CK(clk), .Q(R8[10]) );
  EDFFX1 R8_reg_9_ ( .D(data_in_1[9]), .E(n994), .CK(clk), .Q(R8[9]) );
  EDFFX1 R8_reg_8_ ( .D(data_in_1[8]), .E(n995), .CK(clk), .Q(R8[8]) );
  EDFFX1 R8_reg_7_ ( .D(data_in_1[7]), .E(n994), .CK(clk), .Q(R8[7]) );
  EDFFX1 R8_reg_6_ ( .D(data_in_1[6]), .E(n995), .CK(clk), .Q(R8[6]) );
  EDFFX1 R8_reg_5_ ( .D(data_in_1[5]), .E(n994), .CK(clk), .Q(R8[5]) );
  EDFFX1 R8_reg_4_ ( .D(data_in_1[4]), .E(n995), .CK(clk), .Q(R8[4]) );
  EDFFX1 R8_reg_3_ ( .D(data_in_1[3]), .E(n994), .CK(clk), .Q(R8[3]) );
  EDFFX1 R8_reg_2_ ( .D(data_in_1[2]), .E(n995), .CK(clk), .Q(R8[2]) );
  EDFFX1 R8_reg_1_ ( .D(data_in_1[1]), .E(n994), .CK(clk), .Q(R8[1]) );
  EDFFX1 R8_reg_0_ ( .D(data_in_1[0]), .E(n995), .CK(clk), .Q(R8[0]) );
  EDFFX1 R12_reg_33_ ( .D(data_in_1[33]), .E(n1003), .CK(clk), .Q(R12[33]) );
  EDFFX1 R12_reg_32_ ( .D(data_in_1[32]), .E(n1003), .CK(clk), .Q(R12[32]) );
  EDFFX1 R12_reg_31_ ( .D(data_in_1[31]), .E(n1003), .CK(clk), .Q(R12[31]) );
  EDFFX1 R12_reg_30_ ( .D(data_in_1[30]), .E(n1003), .CK(clk), .Q(R12[30]) );
  EDFFX1 R12_reg_29_ ( .D(data_in_1[29]), .E(n1003), .CK(clk), .Q(R12[29]) );
  EDFFX1 R12_reg_28_ ( .D(data_in_1[28]), .E(n1003), .CK(clk), .Q(R12[28]) );
  EDFFX1 R12_reg_27_ ( .D(data_in_1[27]), .E(n1003), .CK(clk), .Q(R12[27]) );
  EDFFX1 R12_reg_26_ ( .D(data_in_1[26]), .E(n1003), .CK(clk), .Q(R12[26]) );
  EDFFX1 R12_reg_25_ ( .D(data_in_1[25]), .E(n1003), .CK(clk), .Q(R12[25]) );
  EDFFX1 R12_reg_24_ ( .D(data_in_1[24]), .E(n1003), .CK(clk), .Q(R12[24]) );
  EDFFX1 R12_reg_23_ ( .D(data_in_1[23]), .E(n1002), .CK(clk), .Q(R12[23]) );
  EDFFX1 R12_reg_22_ ( .D(data_in_1[22]), .E(n1002), .CK(clk), .Q(R12[22]) );
  EDFFX1 R12_reg_21_ ( .D(data_in_1[21]), .E(n1002), .CK(clk), .Q(R12[21]) );
  EDFFX1 R12_reg_20_ ( .D(data_in_1[20]), .E(n1002), .CK(clk), .Q(R12[20]) );
  EDFFX1 R12_reg_19_ ( .D(data_in_1[19]), .E(n1002), .CK(clk), .Q(R12[19]) );
  EDFFX1 R12_reg_18_ ( .D(data_in_1[18]), .E(n1002), .CK(clk), .Q(R12[18]) );
  EDFFX1 R12_reg_17_ ( .D(data_in_1[17]), .E(n1002), .CK(clk), .Q(R12[17]) );
  EDFFX1 R12_reg_16_ ( .D(data_in_1[16]), .E(n1002), .CK(clk), .Q(R12[16]) );
  EDFFX1 R12_reg_15_ ( .D(data_in_1[15]), .E(n1002), .CK(clk), .Q(R12[15]) );
  EDFFX1 R12_reg_14_ ( .D(data_in_1[14]), .E(n1002), .CK(clk), .Q(R12[14]) );
  EDFFX1 R12_reg_13_ ( .D(data_in_1[13]), .E(n1002), .CK(clk), .Q(R12[13]) );
  EDFFX1 R12_reg_12_ ( .D(data_in_1[12]), .E(n1002), .CK(clk), .Q(R12[12]) );
  EDFFX1 R12_reg_11_ ( .D(data_in_1[11]), .E(n970), .CK(clk), .Q(R12[11]) );
  EDFFX1 R12_reg_10_ ( .D(data_in_1[10]), .E(n970), .CK(clk), .Q(R12[10]) );
  EDFFX1 R12_reg_9_ ( .D(data_in_1[9]), .E(n970), .CK(clk), .Q(R12[9]) );
  EDFFX1 R12_reg_8_ ( .D(data_in_1[8]), .E(n970), .CK(clk), .Q(R12[8]) );
  EDFFX1 R12_reg_7_ ( .D(data_in_1[7]), .E(n970), .CK(clk), .Q(R12[7]) );
  EDFFX1 R12_reg_6_ ( .D(data_in_1[6]), .E(n970), .CK(clk), .Q(R12[6]) );
  EDFFX1 R12_reg_5_ ( .D(data_in_1[5]), .E(n970), .CK(clk), .Q(R12[5]) );
  EDFFX1 R12_reg_4_ ( .D(data_in_1[4]), .E(n1002), .CK(clk), .Q(R12[4]) );
  EDFFX1 R12_reg_3_ ( .D(data_in_1[3]), .E(n1003), .CK(clk), .Q(R12[3]) );
  EDFFX1 R12_reg_2_ ( .D(data_in_1[2]), .E(n1002), .CK(clk), .Q(R12[2]) );
  EDFFX1 R12_reg_1_ ( .D(data_in_1[1]), .E(n1003), .CK(clk), .Q(R12[1]) );
  EDFFX1 R12_reg_0_ ( .D(data_in_1[0]), .E(n1003), .CK(clk), .Q(R12[0]) );
  DFFHQX1 data_out_1_reg_51_ ( .D(n916), .CK(clk), .Q(data_out_1[51]) );
  DFFHQX1 data_out_1_reg_34_ ( .D(n933), .CK(clk), .Q(data_out_1[34]) );
  DFFHQX1 data_out_1_reg_85_ ( .D(n882), .CK(clk), .Q(data_out_1[85]) );
  DFFHQX1 data_out_1_reg_68_ ( .D(n899), .CK(clk), .Q(data_out_1[68]) );
  DFFHQX1 data_out_1_reg_119_ ( .D(n848), .CK(clk), .Q(data_out_1[119]) );
  DFFHQX1 data_out_1_reg_102_ ( .D(n865), .CK(clk), .Q(data_out_1[102]) );
  DFFHQX1 data_out_1_reg_66_ ( .D(n901), .CK(clk), .Q(data_out_1[66]) );
  DFFHQX1 data_out_1_reg_65_ ( .D(n902), .CK(clk), .Q(data_out_1[65]) );
  DFFHQX1 data_out_1_reg_64_ ( .D(n903), .CK(clk), .Q(data_out_1[64]) );
  DFFHQX1 data_out_1_reg_63_ ( .D(n904), .CK(clk), .Q(data_out_1[63]) );
  DFFHQX1 data_out_1_reg_62_ ( .D(n905), .CK(clk), .Q(data_out_1[62]) );
  DFFHQX1 data_out_1_reg_61_ ( .D(n906), .CK(clk), .Q(data_out_1[61]) );
  DFFHQX1 data_out_1_reg_60_ ( .D(n907), .CK(clk), .Q(data_out_1[60]) );
  DFFHQX1 data_out_1_reg_59_ ( .D(n908), .CK(clk), .Q(data_out_1[59]) );
  DFFHQX1 data_out_1_reg_58_ ( .D(n909), .CK(clk), .Q(data_out_1[58]) );
  DFFHQX1 data_out_1_reg_57_ ( .D(n910), .CK(clk), .Q(data_out_1[57]) );
  DFFHQX1 data_out_1_reg_56_ ( .D(n911), .CK(clk), .Q(data_out_1[56]) );
  DFFHQX1 data_out_1_reg_55_ ( .D(n912), .CK(clk), .Q(data_out_1[55]) );
  DFFHQX1 data_out_1_reg_54_ ( .D(n913), .CK(clk), .Q(data_out_1[54]) );
  DFFHQX1 data_out_1_reg_53_ ( .D(n914), .CK(clk), .Q(data_out_1[53]) );
  DFFHQX1 data_out_1_reg_52_ ( .D(n915), .CK(clk), .Q(data_out_1[52]) );
  DFFHQX1 data_out_1_reg_49_ ( .D(n918), .CK(clk), .Q(data_out_1[49]) );
  DFFHQX1 data_out_1_reg_48_ ( .D(n919), .CK(clk), .Q(data_out_1[48]) );
  DFFHQX1 data_out_1_reg_47_ ( .D(n920), .CK(clk), .Q(data_out_1[47]) );
  DFFHQX1 data_out_1_reg_46_ ( .D(n921), .CK(clk), .Q(data_out_1[46]) );
  DFFHQX1 data_out_1_reg_45_ ( .D(n922), .CK(clk), .Q(data_out_1[45]) );
  DFFHQX1 data_out_1_reg_44_ ( .D(n923), .CK(clk), .Q(data_out_1[44]) );
  DFFHQX1 data_out_1_reg_43_ ( .D(n924), .CK(clk), .Q(data_out_1[43]) );
  DFFHQX1 data_out_1_reg_42_ ( .D(n925), .CK(clk), .Q(data_out_1[42]) );
  DFFHQX1 data_out_1_reg_41_ ( .D(n926), .CK(clk), .Q(data_out_1[41]) );
  DFFHQX1 data_out_1_reg_40_ ( .D(n927), .CK(clk), .Q(data_out_1[40]) );
  DFFHQX1 data_out_1_reg_39_ ( .D(n928), .CK(clk), .Q(data_out_1[39]) );
  DFFHQX1 data_out_1_reg_38_ ( .D(n929), .CK(clk), .Q(data_out_1[38]) );
  DFFHQX1 data_out_1_reg_37_ ( .D(n930), .CK(clk), .Q(data_out_1[37]) );
  DFFHQX1 data_out_1_reg_36_ ( .D(n931), .CK(clk), .Q(data_out_1[36]) );
  DFFHQX1 data_out_1_reg_35_ ( .D(n932), .CK(clk), .Q(data_out_1[35]) );
  DFFHQX1 data_out_1_reg_100_ ( .D(n867), .CK(clk), .Q(data_out_1[100]) );
  DFFHQX1 data_out_1_reg_99_ ( .D(n868), .CK(clk), .Q(data_out_1[99]) );
  DFFHQX1 data_out_1_reg_98_ ( .D(n869), .CK(clk), .Q(data_out_1[98]) );
  DFFHQX1 data_out_1_reg_97_ ( .D(n870), .CK(clk), .Q(data_out_1[97]) );
  DFFHQX1 data_out_1_reg_96_ ( .D(n871), .CK(clk), .Q(data_out_1[96]) );
  DFFHQX1 data_out_1_reg_95_ ( .D(n872), .CK(clk), .Q(data_out_1[95]) );
  DFFHQX1 data_out_1_reg_94_ ( .D(n873), .CK(clk), .Q(data_out_1[94]) );
  DFFHQX1 data_out_1_reg_93_ ( .D(n874), .CK(clk), .Q(data_out_1[93]) );
  DFFHQX1 data_out_1_reg_92_ ( .D(n875), .CK(clk), .Q(data_out_1[92]) );
  DFFHQX1 data_out_1_reg_91_ ( .D(n876), .CK(clk), .Q(data_out_1[91]) );
  DFFHQX1 data_out_1_reg_90_ ( .D(n877), .CK(clk), .Q(data_out_1[90]) );
  DFFHQX1 data_out_1_reg_89_ ( .D(n878), .CK(clk), .Q(data_out_1[89]) );
  DFFHQX1 data_out_1_reg_88_ ( .D(n879), .CK(clk), .Q(data_out_1[88]) );
  DFFHQX1 data_out_1_reg_87_ ( .D(n880), .CK(clk), .Q(data_out_1[87]) );
  DFFHQX1 data_out_1_reg_86_ ( .D(n881), .CK(clk), .Q(data_out_1[86]) );
  DFFHQX1 data_out_1_reg_83_ ( .D(n884), .CK(clk), .Q(data_out_1[83]) );
  DFFHQX1 data_out_1_reg_82_ ( .D(n885), .CK(clk), .Q(data_out_1[82]) );
  DFFHQX1 data_out_1_reg_81_ ( .D(n886), .CK(clk), .Q(data_out_1[81]) );
  DFFHQX1 data_out_1_reg_80_ ( .D(n887), .CK(clk), .Q(data_out_1[80]) );
  DFFHQX1 data_out_1_reg_79_ ( .D(n888), .CK(clk), .Q(data_out_1[79]) );
  DFFHQX1 data_out_1_reg_78_ ( .D(n889), .CK(clk), .Q(data_out_1[78]) );
  DFFHQX1 data_out_1_reg_77_ ( .D(n890), .CK(clk), .Q(data_out_1[77]) );
  DFFHQX1 data_out_1_reg_76_ ( .D(n891), .CK(clk), .Q(data_out_1[76]) );
  DFFHQX1 data_out_1_reg_75_ ( .D(n892), .CK(clk), .Q(data_out_1[75]) );
  DFFHQX1 data_out_1_reg_74_ ( .D(n893), .CK(clk), .Q(data_out_1[74]) );
  DFFHQX1 data_out_1_reg_73_ ( .D(n894), .CK(clk), .Q(data_out_1[73]) );
  DFFHQX1 data_out_1_reg_72_ ( .D(n895), .CK(clk), .Q(data_out_1[72]) );
  DFFHQX1 data_out_1_reg_71_ ( .D(n896), .CK(clk), .Q(data_out_1[71]) );
  DFFHQX1 data_out_1_reg_70_ ( .D(n897), .CK(clk), .Q(data_out_1[70]) );
  DFFHQX1 data_out_1_reg_69_ ( .D(n898), .CK(clk), .Q(data_out_1[69]) );
  DFFHQX1 data_out_1_reg_134_ ( .D(n833), .CK(clk), .Q(data_out_1[134]) );
  DFFHQX1 data_out_1_reg_133_ ( .D(n834), .CK(clk), .Q(data_out_1[133]) );
  DFFHQX1 data_out_1_reg_132_ ( .D(n835), .CK(clk), .Q(data_out_1[132]) );
  DFFHQX1 data_out_1_reg_131_ ( .D(n836), .CK(clk), .Q(data_out_1[131]) );
  DFFHQX1 data_out_1_reg_130_ ( .D(n837), .CK(clk), .Q(data_out_1[130]) );
  DFFHQX1 data_out_1_reg_129_ ( .D(n838), .CK(clk), .Q(data_out_1[129]) );
  DFFHQX1 data_out_1_reg_128_ ( .D(n839), .CK(clk), .Q(data_out_1[128]) );
  DFFHQX1 data_out_1_reg_127_ ( .D(n840), .CK(clk), .Q(data_out_1[127]) );
  DFFHQX1 data_out_1_reg_126_ ( .D(n841), .CK(clk), .Q(data_out_1[126]) );
  DFFHQX1 data_out_1_reg_125_ ( .D(n842), .CK(clk), .Q(data_out_1[125]) );
  DFFHQX1 data_out_1_reg_124_ ( .D(n843), .CK(clk), .Q(data_out_1[124]) );
  DFFHQX1 data_out_1_reg_123_ ( .D(n844), .CK(clk), .Q(data_out_1[123]) );
  DFFHQX1 data_out_1_reg_122_ ( .D(n845), .CK(clk), .Q(data_out_1[122]) );
  DFFHQX1 data_out_1_reg_121_ ( .D(n846), .CK(clk), .Q(data_out_1[121]) );
  DFFHQX1 data_out_1_reg_120_ ( .D(n847), .CK(clk), .Q(data_out_1[120]) );
  DFFHQX1 data_out_1_reg_117_ ( .D(n850), .CK(clk), .Q(data_out_1[117]) );
  DFFHQX1 data_out_1_reg_116_ ( .D(n851), .CK(clk), .Q(data_out_1[116]) );
  DFFHQX1 data_out_1_reg_115_ ( .D(n852), .CK(clk), .Q(data_out_1[115]) );
  DFFHQX1 data_out_1_reg_114_ ( .D(n853), .CK(clk), .Q(data_out_1[114]) );
  DFFHQX1 data_out_1_reg_113_ ( .D(n854), .CK(clk), .Q(data_out_1[113]) );
  DFFHQX1 data_out_1_reg_112_ ( .D(n855), .CK(clk), .Q(data_out_1[112]) );
  DFFHQX1 data_out_1_reg_111_ ( .D(n856), .CK(clk), .Q(data_out_1[111]) );
  DFFHQX1 data_out_1_reg_110_ ( .D(n857), .CK(clk), .Q(data_out_1[110]) );
  DFFHQX1 data_out_1_reg_109_ ( .D(n858), .CK(clk), .Q(data_out_1[109]) );
  DFFHQX1 data_out_1_reg_108_ ( .D(n859), .CK(clk), .Q(data_out_1[108]) );
  DFFHQX1 data_out_1_reg_107_ ( .D(n860), .CK(clk), .Q(data_out_1[107]) );
  DFFHQX1 data_out_1_reg_106_ ( .D(n861), .CK(clk), .Q(data_out_1[106]) );
  DFFHQX1 data_out_1_reg_105_ ( .D(n862), .CK(clk), .Q(data_out_1[105]) );
  DFFHQX1 data_out_1_reg_104_ ( .D(n863), .CK(clk), .Q(data_out_1[104]) );
  DFFHQX1 data_out_1_reg_103_ ( .D(n864), .CK(clk), .Q(data_out_1[103]) );
  DFFHQX1 data_out_1_reg_33_ ( .D(n934), .CK(clk), .Q(data_out_1[33]) );
  DFFHQX1 data_out_1_reg_16_ ( .D(n951), .CK(clk), .Q(data_out_1[16]) );
  DFFHQX1 data_out_1_reg_32_ ( .D(n935), .CK(clk), .Q(data_out_1[32]) );
  DFFHQX1 data_out_1_reg_15_ ( .D(n952), .CK(clk), .Q(data_out_1[15]) );
  DFFRHQX1 counter_reg_3_ ( .D(N15), .CK(clk), .RN(rst_n), .Q(counter[3]) );
  DFFRHQX1 counter_reg_1_ ( .D(N13), .CK(clk), .RN(rst_n), .Q(counter[1]) );
  JKFFRXL counter_reg_0_ ( .J(1'b1), .K(1'b1), .CK(clk), .RN(rst_n), .Q(
        counter[0]), .QN(n550) );
  DFFHQX1 data_out_1_reg_31_ ( .D(n936), .CK(clk), .Q(data_out_1[31]) );
  DFFHQX1 data_out_1_reg_30_ ( .D(n937), .CK(clk), .Q(data_out_1[30]) );
  DFFHQX1 data_out_1_reg_29_ ( .D(n938), .CK(clk), .Q(data_out_1[29]) );
  DFFHQX1 data_out_1_reg_28_ ( .D(n939), .CK(clk), .Q(data_out_1[28]) );
  DFFHQX1 data_out_1_reg_27_ ( .D(n940), .CK(clk), .Q(data_out_1[27]) );
  DFFHQX1 data_out_1_reg_26_ ( .D(n941), .CK(clk), .Q(data_out_1[26]) );
  DFFHQX1 data_out_1_reg_25_ ( .D(n942), .CK(clk), .Q(data_out_1[25]) );
  DFFHQX1 data_out_1_reg_14_ ( .D(n953), .CK(clk), .Q(data_out_1[14]) );
  DFFHQX1 data_out_1_reg_13_ ( .D(n954), .CK(clk), .Q(data_out_1[13]) );
  DFFHQX1 data_out_1_reg_12_ ( .D(n955), .CK(clk), .Q(data_out_1[12]) );
  DFFHQX1 data_out_1_reg_11_ ( .D(n956), .CK(clk), .Q(data_out_1[11]) );
  DFFHQX1 data_out_1_reg_10_ ( .D(n957), .CK(clk), .Q(data_out_1[10]) );
  DFFHQX1 data_out_1_reg_24_ ( .D(n943), .CK(clk), .Q(data_out_1[24]) );
  DFFHQX1 data_out_1_reg_22_ ( .D(n945), .CK(clk), .Q(data_out_1[22]) );
  DFFHQX1 data_out_1_reg_21_ ( .D(n946), .CK(clk), .Q(data_out_1[21]) );
  DFFHQX1 data_out_1_reg_20_ ( .D(n947), .CK(clk), .Q(data_out_1[20]) );
  DFFHQX1 data_out_1_reg_19_ ( .D(n948), .CK(clk), .Q(data_out_1[19]) );
  DFFHQX1 data_out_1_reg_18_ ( .D(n949), .CK(clk), .Q(data_out_1[18]) );
  DFFHQX1 data_out_1_reg_17_ ( .D(n950), .CK(clk), .Q(data_out_1[17]) );
  DFFHQX1 data_out_1_reg_9_ ( .D(n958), .CK(clk), .Q(data_out_1[9]) );
  DFFHQX1 data_out_1_reg_7_ ( .D(n960), .CK(clk), .Q(data_out_1[7]) );
  DFFHQX1 data_out_1_reg_6_ ( .D(n961), .CK(clk), .Q(data_out_1[6]) );
  DFFHQX1 data_out_1_reg_4_ ( .D(n963), .CK(clk), .Q(data_out_1[4]) );
  DFFHQX1 data_out_1_reg_3_ ( .D(n964), .CK(clk), .Q(data_out_1[3]) );
  DFFHQX1 data_out_1_reg_2_ ( .D(n965), .CK(clk), .Q(data_out_1[2]) );
  DFFHQX1 data_out_1_reg_1_ ( .D(n966), .CK(clk), .Q(data_out_1[1]) );
  DFFHQX1 data_out_1_reg_0_ ( .D(n967), .CK(clk), .Q(data_out_1[0]) );
  DFFHQX1 data_out_1_reg_5_ ( .D(n962), .CK(clk), .Q(data_out_1[5]) );
  DFFHQXL data_out_1_reg_23_ ( .D(n944), .CK(clk), .Q(data_out_1[23]) );
  DFFHQX1 data_out_1_reg_8_ ( .D(n959), .CK(clk), .Q(data_out_1[8]) );
  DFFRHQX1 counter_reg_2_ ( .D(N14), .CK(clk), .RN(rst_n), .Q(counter[2]) );
  DFFHQX1 data_out_1_reg_67_ ( .D(n900), .CK(clk), .Q(data_out_1[67]) );
  DFFHQX2 data_out_1_reg_50_ ( .D(n917), .CK(clk), .Q(data_out_1[50]) );
  DFFHQX2 data_out_1_reg_101_ ( .D(n866), .CK(clk), .Q(data_out_1[101]) );
  DFFHQX2 data_out_1_reg_84_ ( .D(n883), .CK(clk), .Q(data_out_1[84]) );
  INVX1 U4 ( .A(counter[3]), .Y(n1046) );
  INVX1 U5 ( .A(counter[2]), .Y(n1045) );
  OR3XL U6 ( .A(n1045), .B(n826), .C(n1046), .Y(n1) );
  OR2X2 U7 ( .A(n829), .B(n826), .Y(n2) );
  OR2X2 U8 ( .A(n828), .B(n827), .Y(n3) );
  OR2X2 U9 ( .A(n824), .B(n827), .Y(n4) );
  OR2X2 U10 ( .A(n825), .B(n827), .Y(n5) );
  OR2X2 U11 ( .A(n826), .B(n827), .Y(n6) );
  OR2X2 U12 ( .A(n825), .B(n830), .Y(n7) );
  OR2X2 U13 ( .A(n826), .B(n830), .Y(n8) );
  OR2X2 U14 ( .A(n828), .B(n829), .Y(n9) );
  OR2X2 U15 ( .A(n824), .B(n829), .Y(n10) );
  OR2X2 U16 ( .A(n825), .B(n829), .Y(n11) );
  NOR2X1 U17 ( .A(n830), .B(n828), .Y(N171) );
  INVX2 U18 ( .A(n1024), .Y(n1020) );
  INVXL U19 ( .A(n1027), .Y(n1025) );
  INVXL U20 ( .A(n1027), .Y(n1026) );
  NOR2XL U21 ( .A(n824), .B(n830), .Y(n980) );
  AOI22XL U22 ( .A0(R3[0]), .A1(n1042), .B0(data_out_1[0]), .B1(n1015), .Y(
        n822) );
  AOI22XL U23 ( .A0(R3[1]), .A1(n1042), .B0(data_out_1[1]), .B1(n1015), .Y(
        n820) );
  AOI22XL U24 ( .A0(R3[2]), .A1(n1042), .B0(data_out_1[2]), .B1(n1015), .Y(
        n818) );
  AOI22XL U25 ( .A0(R3[3]), .A1(n1042), .B0(data_out_1[3]), .B1(n1015), .Y(
        n816) );
  AOI22XL U26 ( .A0(R3[5]), .A1(n1042), .B0(data_out_1[5]), .B1(n1015), .Y(
        n812) );
  AOI22XL U27 ( .A0(R3[7]), .A1(n1041), .B0(data_out_1[7]), .B1(n1020), .Y(
        n808) );
  AOI22XL U28 ( .A0(R3[8]), .A1(n1041), .B0(data_out_1[8]), .B1(n1020), .Y(
        n806) );
  AOI22XL U29 ( .A0(R3[17]), .A1(n1041), .B0(data_out_1[17]), .B1(n1015), .Y(
        n788) );
  AOI22XL U30 ( .A0(R3[18]), .A1(n1041), .B0(data_out_1[18]), .B1(n1015), .Y(
        n786) );
  AOI22XL U31 ( .A0(R3[23]), .A1(n1040), .B0(data_out_1[23]), .B1(n1015), .Y(
        n776) );
  AOI22XL U32 ( .A0(R15[30]), .A1(n1041), .B0(data_out_1[132]), .B1(n1020), 
        .Y(n558) );
  AOI22XL U33 ( .A0(R15[31]), .A1(n1038), .B0(data_out_1[133]), .B1(n1021), 
        .Y(n556) );
  AOI22XL U34 ( .A0(R15[32]), .A1(n1037), .B0(data_out_1[134]), .B1(n1020), 
        .Y(n554) );
  NAND2XL U35 ( .A(counter[3]), .B(n1045), .Y(n827) );
  NAND2XL U36 ( .A(counter[2]), .B(n1046), .Y(n829) );
  OAI22XL U37 ( .A0(n831), .A1(n1045), .B0(counter[2]), .B1(n826), .Y(N14) );
  INVX1 U38 ( .A(n1024), .Y(n1022) );
  INVX1 U39 ( .A(n1026), .Y(n1023) );
  INVX1 U40 ( .A(n1024), .Y(n1021) );
  INVX1 U41 ( .A(n1026), .Y(n1017) );
  INVX1 U42 ( .A(n1025), .Y(n1018) );
  INVX1 U43 ( .A(n1025), .Y(n1019) );
  INVX1 U44 ( .A(n12), .Y(n1015) );
  INVX1 U45 ( .A(n1026), .Y(n1016) );
  INVX1 U46 ( .A(n1027), .Y(n1024) );
  INVX1 U47 ( .A(n12), .Y(n1027) );
  CLKINVX3 U48 ( .A(n1), .Y(n1028) );
  OR4X2 U49 ( .A(n968), .B(n969), .C(n1028), .D(N171), .Y(n12) );
  CLKINVX3 U50 ( .A(n1009), .Y(n1006) );
  CLKINVX3 U51 ( .A(n1009), .Y(n1005) );
  CLKINVX3 U52 ( .A(n1009), .Y(n1007) );
  INVX1 U53 ( .A(n1043), .Y(n1033) );
  INVX1 U54 ( .A(n1043), .Y(n1036) );
  INVX1 U55 ( .A(n1043), .Y(n1035) );
  INVX1 U56 ( .A(n1043), .Y(n1034) );
  INVX1 U57 ( .A(n1043), .Y(n1038) );
  INVX1 U58 ( .A(n1043), .Y(n1037) );
  INVX1 U59 ( .A(n1043), .Y(n1041) );
  INVX1 U60 ( .A(n1043), .Y(n1040) );
  INVX1 U61 ( .A(n1043), .Y(n1039) );
  CLKINVX3 U62 ( .A(n1), .Y(n1032) );
  CLKINVX3 U63 ( .A(n1), .Y(n1029) );
  CLKINVX3 U64 ( .A(n1), .Y(n1031) );
  CLKINVX3 U65 ( .A(n1), .Y(n1030) );
  CLKINVX3 U66 ( .A(n1009), .Y(n1008) );
  INVX1 U67 ( .A(n1043), .Y(n1042) );
  CLKINVX3 U68 ( .A(n1014), .Y(n1011) );
  CLKINVX3 U69 ( .A(n1014), .Y(n1010) );
  CLKINVX3 U70 ( .A(n1014), .Y(n1013) );
  CLKINVX3 U71 ( .A(n1014), .Y(n1012) );
  INVX1 U72 ( .A(n1004), .Y(n1002) );
  INVX1 U73 ( .A(n6), .Y(n1001) );
  INVX1 U74 ( .A(n4), .Y(n999) );
  INVX1 U75 ( .A(n5), .Y(n997) );
  INVX1 U76 ( .A(n3), .Y(n995) );
  INVX1 U77 ( .A(n2), .Y(n992) );
  INVX1 U78 ( .A(n2), .Y(n993) );
  INVX1 U79 ( .A(n10), .Y(n991) );
  INVX1 U80 ( .A(n11), .Y(n989) );
  INVX1 U81 ( .A(n9), .Y(n987) );
  INVX1 U82 ( .A(n8), .Y(n985) );
  INVX1 U83 ( .A(n983), .Y(n982) );
  INVX1 U84 ( .A(n7), .Y(n979) );
  INVX1 U85 ( .A(n1004), .Y(n1003) );
  INVX1 U86 ( .A(n6), .Y(n1000) );
  INVX1 U87 ( .A(n4), .Y(n998) );
  INVX1 U88 ( .A(n5), .Y(n996) );
  INVX1 U89 ( .A(n3), .Y(n994) );
  INVX1 U90 ( .A(n10), .Y(n990) );
  INVX1 U91 ( .A(n11), .Y(n988) );
  INVX1 U92 ( .A(n9), .Y(n986) );
  INVX1 U93 ( .A(n8), .Y(n984) );
  INVX1 U94 ( .A(n983), .Y(n981) );
  INVX1 U95 ( .A(n980), .Y(n983) );
  INVX1 U96 ( .A(n7), .Y(n978) );
  INVX1 U97 ( .A(n968), .Y(n1014) );
  INVX1 U98 ( .A(n969), .Y(n1009) );
  INVX1 U99 ( .A(N171), .Y(n1043) );
  INVX1 U100 ( .A(n970), .Y(n1004) );
  NOR3X1 U101 ( .A(n1046), .B(n1045), .C(n825), .Y(n969) );
  NOR3X1 U102 ( .A(n1046), .B(n1045), .C(n824), .Y(n968) );
  NAND2X1 U103 ( .A(n1045), .B(n1046), .Y(n830) );
  NOR3X1 U104 ( .A(n1046), .B(n1045), .C(n828), .Y(n970) );
  OAI211X1 U105 ( .A0(n831), .A1(n1046), .B0(n827), .C0(n2), .Y(N15) );
  NAND2X1 U106 ( .A(n824), .B(n825), .Y(N13) );
  NAND2X1 U107 ( .A(counter[0]), .B(n1044), .Y(n825) );
  NAND2X1 U108 ( .A(counter[1]), .B(counter[0]), .Y(n826) );
  NAND2X1 U109 ( .A(n618), .B(n619), .Y(n865) );
  AOI222X1 U110 ( .A0(R12[0]), .A1(n1008), .B0(R14[0]), .B1(n1031), .C0(R13[0]), .C1(n1010), .Y(n619) );
  AOI22X1 U111 ( .A0(R15[0]), .A1(n1034), .B0(data_out_1[102]), .B1(n1021), 
        .Y(n618) );
  NAND2X1 U112 ( .A(n616), .B(n617), .Y(n864) );
  AOI222X1 U113 ( .A0(R12[1]), .A1(n1006), .B0(R14[1]), .B1(n1030), .C0(R13[1]), .C1(n1010), .Y(n617) );
  AOI22X1 U114 ( .A0(R15[1]), .A1(n1034), .B0(data_out_1[103]), .B1(n1021), 
        .Y(n616) );
  NAND2X1 U115 ( .A(n614), .B(n615), .Y(n863) );
  AOI222X1 U116 ( .A0(R12[2]), .A1(n1007), .B0(R14[2]), .B1(n1029), .C0(R13[2]), .C1(n1010), .Y(n615) );
  AOI22X1 U117 ( .A0(R15[2]), .A1(n1034), .B0(data_out_1[104]), .B1(n1021), 
        .Y(n614) );
  NAND2X1 U118 ( .A(n612), .B(n613), .Y(n862) );
  AOI222X1 U119 ( .A0(R12[3]), .A1(n1005), .B0(R14[3]), .B1(n1030), .C0(R13[3]), .C1(n1010), .Y(n613) );
  AOI22X1 U120 ( .A0(R15[3]), .A1(n1034), .B0(data_out_1[105]), .B1(n1021), 
        .Y(n612) );
  NAND2X1 U121 ( .A(n610), .B(n611), .Y(n861) );
  AOI222X1 U122 ( .A0(R12[4]), .A1(n1008), .B0(R14[4]), .B1(n1030), .C0(R13[4]), .C1(n1010), .Y(n611) );
  AOI22X1 U123 ( .A0(R15[4]), .A1(n1034), .B0(data_out_1[106]), .B1(n1021), 
        .Y(n610) );
  NAND2X1 U124 ( .A(n608), .B(n609), .Y(n860) );
  AOI222X1 U125 ( .A0(R12[5]), .A1(n1006), .B0(R14[5]), .B1(n1031), .C0(R13[5]), .C1(n1010), .Y(n609) );
  AOI22X1 U126 ( .A0(R15[5]), .A1(n1034), .B0(data_out_1[107]), .B1(n1021), 
        .Y(n608) );
  NAND2X1 U127 ( .A(n606), .B(n607), .Y(n859) );
  AOI222X1 U128 ( .A0(R12[6]), .A1(n1007), .B0(R14[6]), .B1(n1031), .C0(R13[6]), .C1(n1010), .Y(n607) );
  AOI22X1 U129 ( .A0(R15[6]), .A1(n1034), .B0(data_out_1[108]), .B1(n1022), 
        .Y(n606) );
  NAND2X1 U130 ( .A(n604), .B(n605), .Y(n858) );
  AOI222X1 U131 ( .A0(R12[7]), .A1(n1005), .B0(R14[7]), .B1(n1029), .C0(R13[7]), .C1(n1010), .Y(n605) );
  AOI22X1 U132 ( .A0(R15[7]), .A1(n1034), .B0(data_out_1[109]), .B1(n1022), 
        .Y(n604) );
  NAND2X1 U133 ( .A(n602), .B(n603), .Y(n857) );
  AOI222X1 U134 ( .A0(R12[8]), .A1(n1008), .B0(R14[8]), .B1(n1030), .C0(R13[8]), .C1(n1010), .Y(n603) );
  AOI22X1 U135 ( .A0(R15[8]), .A1(n1033), .B0(data_out_1[110]), .B1(n1022), 
        .Y(n602) );
  NAND2X1 U136 ( .A(n600), .B(n601), .Y(n856) );
  AOI222X1 U137 ( .A0(R12[9]), .A1(n1006), .B0(R14[9]), .B1(n1030), .C0(R13[9]), .C1(n1010), .Y(n601) );
  AOI22X1 U138 ( .A0(R15[9]), .A1(n1033), .B0(data_out_1[111]), .B1(n1022), 
        .Y(n600) );
  NAND2X1 U139 ( .A(n598), .B(n599), .Y(n855) );
  AOI222X1 U140 ( .A0(R12[10]), .A1(n1007), .B0(R14[10]), .B1(n1031), .C0(
        R13[10]), .C1(n1010), .Y(n599) );
  AOI22X1 U141 ( .A0(R15[10]), .A1(n1033), .B0(data_out_1[112]), .B1(n1022), 
        .Y(n598) );
  NAND2X1 U142 ( .A(n596), .B(n597), .Y(n854) );
  AOI222X1 U143 ( .A0(R12[11]), .A1(n1005), .B0(R14[11]), .B1(n1030), .C0(
        R13[11]), .C1(n1010), .Y(n597) );
  AOI22X1 U144 ( .A0(R15[11]), .A1(n1033), .B0(data_out_1[113]), .B1(n1022), 
        .Y(n596) );
  NAND2X1 U145 ( .A(n594), .B(n595), .Y(n853) );
  AOI222X1 U146 ( .A0(R12[12]), .A1(n1008), .B0(R14[12]), .B1(n1029), .C0(
        R13[12]), .C1(n1010), .Y(n595) );
  AOI22X1 U147 ( .A0(R15[12]), .A1(n1033), .B0(data_out_1[114]), .B1(n1022), 
        .Y(n594) );
  NAND2X1 U148 ( .A(n592), .B(n593), .Y(n852) );
  AOI222X1 U149 ( .A0(R12[13]), .A1(n1006), .B0(R14[13]), .B1(n1030), .C0(
        R13[13]), .C1(n1010), .Y(n593) );
  AOI22X1 U150 ( .A0(R15[13]), .A1(n1033), .B0(data_out_1[115]), .B1(n1022), 
        .Y(n592) );
  NAND2X1 U151 ( .A(n590), .B(n591), .Y(n851) );
  AOI222X1 U152 ( .A0(R12[14]), .A1(n1007), .B0(R14[14]), .B1(n1030), .C0(
        R13[14]), .C1(n1010), .Y(n591) );
  AOI22X1 U153 ( .A0(R15[14]), .A1(n1033), .B0(data_out_1[116]), .B1(n1022), 
        .Y(n590) );
  NAND2X1 U154 ( .A(n588), .B(n589), .Y(n850) );
  AOI222X1 U155 ( .A0(R12[15]), .A1(n1005), .B0(R14[15]), .B1(n1032), .C0(
        R13[15]), .C1(n1010), .Y(n589) );
  AOI22X1 U156 ( .A0(R15[15]), .A1(n1033), .B0(data_out_1[117]), .B1(n1022), 
        .Y(n588) );
  NAND2X1 U157 ( .A(n586), .B(n587), .Y(n849) );
  AOI222X1 U158 ( .A0(R12[16]), .A1(n1008), .B0(R14[16]), .B1(n1028), .C0(
        R13[16]), .C1(n968), .Y(n587) );
  AOI22XL U159 ( .A0(R15[16]), .A1(n1033), .B0(data_out_1[118]), .B1(n1022), 
        .Y(n586) );
  NAND2X1 U160 ( .A(n584), .B(n585), .Y(n848) );
  AOI222X1 U161 ( .A0(R12[17]), .A1(n1006), .B0(R14[17]), .B1(n1028), .C0(
        R13[17]), .C1(n1012), .Y(n585) );
  AOI22X1 U162 ( .A0(R15[17]), .A1(n1033), .B0(data_out_1[119]), .B1(n1022), 
        .Y(n584) );
  NAND2X1 U163 ( .A(n582), .B(n583), .Y(n847) );
  AOI222X1 U164 ( .A0(R12[18]), .A1(n1005), .B0(R14[18]), .B1(n1028), .C0(
        R13[18]), .C1(n1012), .Y(n583) );
  AOI22X1 U165 ( .A0(R15[18]), .A1(n1033), .B0(data_out_1[120]), .B1(n1023), 
        .Y(n582) );
  NAND2X1 U166 ( .A(n580), .B(n581), .Y(n846) );
  AOI222X1 U167 ( .A0(R12[19]), .A1(n1007), .B0(R14[19]), .B1(n1028), .C0(
        R13[19]), .C1(n1011), .Y(n581) );
  AOI22X1 U168 ( .A0(R15[19]), .A1(n1033), .B0(data_out_1[121]), .B1(n1023), 
        .Y(n580) );
  NAND2X1 U169 ( .A(n578), .B(n579), .Y(n845) );
  AOI222X1 U170 ( .A0(R12[20]), .A1(n969), .B0(R14[20]), .B1(n1028), .C0(
        R13[20]), .C1(n1012), .Y(n579) );
  AOI22X1 U171 ( .A0(R15[20]), .A1(n1033), .B0(data_out_1[122]), .B1(n1023), 
        .Y(n578) );
  NAND2X1 U172 ( .A(n576), .B(n577), .Y(n844) );
  AOI222X1 U173 ( .A0(R12[21]), .A1(n969), .B0(R14[21]), .B1(n1028), .C0(
        R13[21]), .C1(n1011), .Y(n577) );
  AOI22X1 U174 ( .A0(R15[21]), .A1(n1035), .B0(data_out_1[123]), .B1(n1023), 
        .Y(n576) );
  NAND2X1 U175 ( .A(n574), .B(n575), .Y(n843) );
  AOI222X1 U176 ( .A0(R12[22]), .A1(n969), .B0(R14[22]), .B1(n1028), .C0(
        R13[22]), .C1(n1010), .Y(n575) );
  AOI22X1 U177 ( .A0(R15[22]), .A1(n1033), .B0(data_out_1[124]), .B1(n1023), 
        .Y(n574) );
  NAND2X1 U178 ( .A(n572), .B(n573), .Y(n842) );
  AOI222X1 U179 ( .A0(R12[23]), .A1(n969), .B0(R14[23]), .B1(n1028), .C0(
        R13[23]), .C1(n968), .Y(n573) );
  AOI22X1 U180 ( .A0(R15[23]), .A1(n1034), .B0(data_out_1[125]), .B1(n1023), 
        .Y(n572) );
  NAND2X1 U181 ( .A(n570), .B(n571), .Y(n841) );
  AOI222X1 U182 ( .A0(R12[24]), .A1(n1006), .B0(R14[24]), .B1(n1028), .C0(
        R13[24]), .C1(n1013), .Y(n571) );
  AOI22X1 U183 ( .A0(R15[24]), .A1(n1041), .B0(data_out_1[126]), .B1(n1023), 
        .Y(n570) );
  NAND2X1 U184 ( .A(n568), .B(n569), .Y(n840) );
  AOI222X1 U185 ( .A0(R12[25]), .A1(n1008), .B0(R14[25]), .B1(n1028), .C0(
        R13[25]), .C1(n1011), .Y(n569) );
  AOI22X1 U186 ( .A0(R15[25]), .A1(n1038), .B0(data_out_1[127]), .B1(n1023), 
        .Y(n568) );
  NAND2X1 U187 ( .A(n566), .B(n567), .Y(n839) );
  AOI222X1 U188 ( .A0(R12[26]), .A1(n1007), .B0(R14[26]), .B1(n1028), .C0(
        R13[26]), .C1(n1013), .Y(n567) );
  AOI22X1 U189 ( .A0(R15[26]), .A1(n1037), .B0(data_out_1[128]), .B1(n1023), 
        .Y(n566) );
  NAND2X1 U190 ( .A(n564), .B(n565), .Y(n838) );
  AOI222X1 U191 ( .A0(R12[27]), .A1(n1008), .B0(R14[27]), .B1(n1028), .C0(
        R13[27]), .C1(n1012), .Y(n565) );
  AOI22X1 U192 ( .A0(R15[27]), .A1(n1035), .B0(data_out_1[129]), .B1(n1023), 
        .Y(n564) );
  NAND2X1 U193 ( .A(n562), .B(n563), .Y(n837) );
  AOI222X1 U194 ( .A0(R12[28]), .A1(n1006), .B0(R14[28]), .B1(n1028), .C0(
        R13[28]), .C1(n1012), .Y(n563) );
  AOI22X1 U195 ( .A0(R15[28]), .A1(n1033), .B0(data_out_1[130]), .B1(n1023), 
        .Y(n562) );
  NAND2X1 U196 ( .A(n560), .B(n561), .Y(n836) );
  AOI222X1 U197 ( .A0(R12[29]), .A1(n1005), .B0(R14[29]), .B1(n1028), .C0(
        R13[29]), .C1(n1013), .Y(n561) );
  AOI22X1 U198 ( .A0(R15[29]), .A1(n1034), .B0(data_out_1[131]), .B1(n1023), 
        .Y(n560) );
  NAND2X1 U199 ( .A(n686), .B(n687), .Y(n899) );
  AOI222X1 U200 ( .A0(R8[0]), .A1(n1005), .B0(R10[0]), .B1(n1030), .C0(R9[0]), 
        .C1(n1011), .Y(n687) );
  AOI22X1 U201 ( .A0(R11[0]), .A1(n1037), .B0(data_out_1[68]), .B1(n1019), .Y(
        n686) );
  NAND2X1 U202 ( .A(n684), .B(n685), .Y(n898) );
  AOI222X1 U203 ( .A0(R8[1]), .A1(n1005), .B0(R10[1]), .B1(n1030), .C0(R9[1]), 
        .C1(n1013), .Y(n685) );
  AOI22X1 U204 ( .A0(R11[1]), .A1(n1037), .B0(data_out_1[69]), .B1(n1019), .Y(
        n684) );
  NAND2X1 U205 ( .A(n682), .B(n683), .Y(n897) );
  AOI222X1 U206 ( .A0(R8[2]), .A1(n1005), .B0(R10[2]), .B1(n1030), .C0(R9[2]), 
        .C1(n1012), .Y(n683) );
  AOI22X1 U207 ( .A0(R11[2]), .A1(n1037), .B0(data_out_1[70]), .B1(n1019), .Y(
        n682) );
  NAND2X1 U208 ( .A(n680), .B(n681), .Y(n896) );
  AOI222X1 U209 ( .A0(R8[3]), .A1(n1005), .B0(R10[3]), .B1(n1030), .C0(R9[3]), 
        .C1(n1011), .Y(n681) );
  AOI22X1 U210 ( .A0(R11[3]), .A1(n1036), .B0(data_out_1[71]), .B1(n1019), .Y(
        n680) );
  NAND2X1 U211 ( .A(n678), .B(n679), .Y(n895) );
  AOI222X1 U212 ( .A0(R8[4]), .A1(n1005), .B0(R10[4]), .B1(n1030), .C0(R9[4]), 
        .C1(n1013), .Y(n679) );
  AOI22X1 U213 ( .A0(R11[4]), .A1(n1036), .B0(data_out_1[72]), .B1(n1020), .Y(
        n678) );
  NAND2X1 U214 ( .A(n676), .B(n677), .Y(n894) );
  AOI222X1 U215 ( .A0(R8[5]), .A1(n1005), .B0(R10[5]), .B1(n1030), .C0(R9[5]), 
        .C1(n1012), .Y(n677) );
  AOI22X1 U216 ( .A0(R11[5]), .A1(n1036), .B0(data_out_1[73]), .B1(n1020), .Y(
        n676) );
  NAND2X1 U217 ( .A(n674), .B(n675), .Y(n893) );
  AOI222X1 U218 ( .A0(R8[6]), .A1(n1005), .B0(R10[6]), .B1(n1030), .C0(R9[6]), 
        .C1(n1011), .Y(n675) );
  AOI22X1 U219 ( .A0(R11[6]), .A1(n1036), .B0(data_out_1[74]), .B1(n1020), .Y(
        n674) );
  NAND2X1 U220 ( .A(n672), .B(n673), .Y(n892) );
  AOI222X1 U221 ( .A0(R8[7]), .A1(n1005), .B0(R10[7]), .B1(n1030), .C0(R9[7]), 
        .C1(n1013), .Y(n673) );
  AOI22X1 U222 ( .A0(R11[7]), .A1(n1036), .B0(data_out_1[75]), .B1(n1020), .Y(
        n672) );
  NAND2X1 U223 ( .A(n670), .B(n671), .Y(n891) );
  AOI222X1 U224 ( .A0(R8[8]), .A1(n1005), .B0(R10[8]), .B1(n1030), .C0(R9[8]), 
        .C1(n1012), .Y(n671) );
  AOI22X1 U225 ( .A0(R11[8]), .A1(n1036), .B0(data_out_1[76]), .B1(n1020), .Y(
        n670) );
  NAND2X1 U226 ( .A(n668), .B(n669), .Y(n890) );
  AOI222X1 U227 ( .A0(R8[9]), .A1(n1005), .B0(R10[9]), .B1(n1030), .C0(R9[9]), 
        .C1(n1011), .Y(n669) );
  AOI22X1 U228 ( .A0(R11[9]), .A1(n1036), .B0(data_out_1[77]), .B1(n1020), .Y(
        n668) );
  NAND2X1 U229 ( .A(n666), .B(n667), .Y(n889) );
  AOI222X1 U230 ( .A0(R8[10]), .A1(n1005), .B0(R10[10]), .B1(n1030), .C0(
        R9[10]), .C1(n1013), .Y(n667) );
  AOI22X1 U231 ( .A0(R11[10]), .A1(n1036), .B0(data_out_1[78]), .B1(n1020), 
        .Y(n666) );
  NAND2X1 U232 ( .A(n664), .B(n665), .Y(n888) );
  AOI222X1 U233 ( .A0(R8[11]), .A1(n1005), .B0(R10[11]), .B1(n1030), .C0(
        R9[11]), .C1(n1012), .Y(n665) );
  AOI22X1 U234 ( .A0(R11[11]), .A1(n1036), .B0(data_out_1[79]), .B1(n1020), 
        .Y(n664) );
  NAND2X1 U235 ( .A(n662), .B(n663), .Y(n887) );
  AOI222X1 U236 ( .A0(R8[12]), .A1(n1005), .B0(R10[12]), .B1(n1030), .C0(
        R9[12]), .C1(n1011), .Y(n663) );
  AOI22X1 U237 ( .A0(R11[12]), .A1(n1036), .B0(data_out_1[80]), .B1(n1020), 
        .Y(n662) );
  NAND2X1 U238 ( .A(n660), .B(n661), .Y(n886) );
  AOI222X1 U239 ( .A0(R8[13]), .A1(n1005), .B0(R10[13]), .B1(n1030), .C0(
        R9[13]), .C1(n1013), .Y(n661) );
  AOI22X1 U240 ( .A0(R11[13]), .A1(n1036), .B0(data_out_1[81]), .B1(n1020), 
        .Y(n660) );
  NAND2X1 U241 ( .A(n658), .B(n659), .Y(n885) );
  AOI222X1 U242 ( .A0(R8[14]), .A1(n1005), .B0(R10[14]), .B1(n1029), .C0(
        R9[14]), .C1(n1011), .Y(n659) );
  AOI22X1 U243 ( .A0(R11[14]), .A1(n1036), .B0(data_out_1[82]), .B1(n1020), 
        .Y(n658) );
  NAND2X1 U244 ( .A(n656), .B(n657), .Y(n884) );
  AOI222X1 U245 ( .A0(R8[15]), .A1(n1005), .B0(R10[15]), .B1(n1029), .C0(
        R9[15]), .C1(n1011), .Y(n657) );
  AOI22X1 U246 ( .A0(R11[15]), .A1(n1036), .B0(data_out_1[83]), .B1(n1020), 
        .Y(n656) );
  NAND2X1 U247 ( .A(n654), .B(n655), .Y(n883) );
  AOI222X1 U248 ( .A0(R8[16]), .A1(n1006), .B0(R10[16]), .B1(n1029), .C0(
        R9[16]), .C1(n1011), .Y(n655) );
  AOI22XL U249 ( .A0(R11[16]), .A1(n1035), .B0(data_out_1[84]), .B1(n1020), 
        .Y(n654) );
  NAND2X1 U250 ( .A(n652), .B(n653), .Y(n882) );
  AOI222X1 U251 ( .A0(R8[17]), .A1(n1007), .B0(R10[17]), .B1(n1029), .C0(
        R9[17]), .C1(n1011), .Y(n653) );
  AOI22X1 U252 ( .A0(R11[17]), .A1(n1035), .B0(data_out_1[85]), .B1(n1020), 
        .Y(n652) );
  NAND2X1 U253 ( .A(n650), .B(n651), .Y(n881) );
  AOI222X1 U254 ( .A0(R8[18]), .A1(n1005), .B0(R10[18]), .B1(n1029), .C0(
        R9[18]), .C1(n1011), .Y(n651) );
  AOI22X1 U255 ( .A0(R11[18]), .A1(n1035), .B0(data_out_1[86]), .B1(n1020), 
        .Y(n650) );
  NAND2X1 U256 ( .A(n648), .B(n649), .Y(n880) );
  AOI222X1 U257 ( .A0(R8[19]), .A1(n1006), .B0(R10[19]), .B1(n1029), .C0(
        R9[19]), .C1(n1011), .Y(n649) );
  AOI22X1 U258 ( .A0(R11[19]), .A1(n1035), .B0(data_out_1[87]), .B1(n1020), 
        .Y(n648) );
  NAND2X1 U259 ( .A(n646), .B(n647), .Y(n879) );
  AOI222X1 U260 ( .A0(R8[20]), .A1(n1007), .B0(R10[20]), .B1(n1029), .C0(
        R9[20]), .C1(n1011), .Y(n647) );
  AOI22X1 U261 ( .A0(R11[20]), .A1(n1035), .B0(data_out_1[88]), .B1(n1020), 
        .Y(n646) );
  NAND2X1 U262 ( .A(n644), .B(n645), .Y(n878) );
  AOI222X1 U263 ( .A0(R8[21]), .A1(n1008), .B0(R10[21]), .B1(n1029), .C0(
        R9[21]), .C1(n1011), .Y(n645) );
  AOI22X1 U264 ( .A0(R11[21]), .A1(n1035), .B0(data_out_1[89]), .B1(n1020), 
        .Y(n644) );
  NAND2X1 U265 ( .A(n642), .B(n643), .Y(n877) );
  AOI222X1 U266 ( .A0(R8[22]), .A1(n1005), .B0(R10[22]), .B1(n1029), .C0(
        R9[22]), .C1(n1011), .Y(n643) );
  AOI22X1 U267 ( .A0(R11[22]), .A1(n1035), .B0(data_out_1[90]), .B1(n1018), 
        .Y(n642) );
  NAND2X1 U268 ( .A(n640), .B(n641), .Y(n876) );
  AOI222X1 U269 ( .A0(R8[23]), .A1(n1006), .B0(R10[23]), .B1(n1029), .C0(
        R9[23]), .C1(n1011), .Y(n641) );
  AOI22X1 U270 ( .A0(R11[23]), .A1(n1035), .B0(data_out_1[91]), .B1(n1020), 
        .Y(n640) );
  NAND2X1 U271 ( .A(n638), .B(n639), .Y(n875) );
  AOI222X1 U272 ( .A0(R8[24]), .A1(n1007), .B0(R10[24]), .B1(n1029), .C0(
        R9[24]), .C1(n1011), .Y(n639) );
  AOI22X1 U273 ( .A0(R11[24]), .A1(n1035), .B0(data_out_1[92]), .B1(n1020), 
        .Y(n638) );
  NAND2X1 U274 ( .A(n636), .B(n637), .Y(n874) );
  AOI222X1 U275 ( .A0(R8[25]), .A1(n1008), .B0(R10[25]), .B1(n1029), .C0(
        R9[25]), .C1(n1011), .Y(n637) );
  AOI22X1 U276 ( .A0(R11[25]), .A1(n1035), .B0(data_out_1[93]), .B1(n1019), 
        .Y(n636) );
  NAND2X1 U277 ( .A(n634), .B(n635), .Y(n873) );
  AOI222X1 U278 ( .A0(R8[26]), .A1(n1005), .B0(R10[26]), .B1(n1029), .C0(
        R9[26]), .C1(n1011), .Y(n635) );
  AOI22X1 U279 ( .A0(R11[26]), .A1(n1035), .B0(data_out_1[94]), .B1(n1020), 
        .Y(n634) );
  NAND2X1 U280 ( .A(n632), .B(n633), .Y(n872) );
  AOI222X1 U281 ( .A0(R8[27]), .A1(n1006), .B0(R10[27]), .B1(n1029), .C0(
        R9[27]), .C1(n1011), .Y(n633) );
  AOI22X1 U282 ( .A0(R11[27]), .A1(n1035), .B0(data_out_1[95]), .B1(n1020), 
        .Y(n632) );
  NAND2X1 U283 ( .A(n630), .B(n631), .Y(n871) );
  AOI222X1 U284 ( .A0(R8[28]), .A1(n1007), .B0(R10[28]), .B1(n1029), .C0(
        R9[28]), .C1(n1011), .Y(n631) );
  AOI22X1 U285 ( .A0(R11[28]), .A1(n1035), .B0(data_out_1[96]), .B1(n1021), 
        .Y(n630) );
  NAND2X1 U286 ( .A(n628), .B(n629), .Y(n870) );
  AOI222X1 U287 ( .A0(R8[29]), .A1(n1008), .B0(R10[29]), .B1(n1029), .C0(
        R9[29]), .C1(n1011), .Y(n629) );
  AOI22X1 U288 ( .A0(R11[29]), .A1(n1034), .B0(data_out_1[97]), .B1(n1021), 
        .Y(n628) );
  NAND2X1 U289 ( .A(n626), .B(n627), .Y(n869) );
  AOI222X1 U290 ( .A0(R8[30]), .A1(n1005), .B0(R10[30]), .B1(n1029), .C0(
        R9[30]), .C1(n1011), .Y(n627) );
  AOI22X1 U291 ( .A0(R11[30]), .A1(n1034), .B0(data_out_1[98]), .B1(n1021), 
        .Y(n626) );
  NAND2X1 U292 ( .A(n624), .B(n625), .Y(n868) );
  AOI222X1 U293 ( .A0(R8[31]), .A1(n1006), .B0(R10[31]), .B1(n1029), .C0(
        R9[31]), .C1(n1011), .Y(n625) );
  AOI22X1 U294 ( .A0(R11[31]), .A1(n1034), .B0(data_out_1[99]), .B1(n1021), 
        .Y(n624) );
  NAND2X1 U295 ( .A(n622), .B(n623), .Y(n867) );
  AOI222X1 U296 ( .A0(R8[32]), .A1(n1006), .B0(R10[32]), .B1(n1031), .C0(
        R9[32]), .C1(n1010), .Y(n623) );
  AOI22X1 U297 ( .A0(R11[32]), .A1(n1034), .B0(data_out_1[100]), .B1(n1021), 
        .Y(n622) );
  NAND2X1 U298 ( .A(n620), .B(n621), .Y(n866) );
  AOI222X1 U299 ( .A0(R8[33]), .A1(n1006), .B0(R10[33]), .B1(n1029), .C0(
        R9[33]), .C1(n1010), .Y(n621) );
  AOI22XL U300 ( .A0(R11[33]), .A1(n1034), .B0(data_out_1[101]), .B1(n1021), 
        .Y(n620) );
  NAND2X1 U301 ( .A(n754), .B(n755), .Y(n933) );
  AOI222X1 U302 ( .A0(R4[0]), .A1(n1008), .B0(R6[0]), .B1(n1030), .C0(R5[0]), 
        .C1(n1012), .Y(n755) );
  AOI22X1 U303 ( .A0(R7[0]), .A1(n1039), .B0(data_out_1[34]), .B1(n1016), .Y(
        n754) );
  NAND2X1 U304 ( .A(n752), .B(n753), .Y(n932) );
  AOI222X1 U305 ( .A0(R4[1]), .A1(n1005), .B0(R6[1]), .B1(n1031), .C0(R5[1]), 
        .C1(n1012), .Y(n753) );
  AOI22X1 U306 ( .A0(R7[1]), .A1(n1039), .B0(data_out_1[35]), .B1(n1016), .Y(
        n752) );
  NAND2X1 U307 ( .A(n750), .B(n751), .Y(n931) );
  AOI222X1 U308 ( .A0(R4[2]), .A1(n1007), .B0(R6[2]), .B1(n1031), .C0(R5[2]), 
        .C1(n1012), .Y(n751) );
  AOI22X1 U309 ( .A0(R7[2]), .A1(n1039), .B0(data_out_1[36]), .B1(n1017), .Y(
        n750) );
  NAND2X1 U310 ( .A(n748), .B(n749), .Y(n930) );
  AOI222X1 U311 ( .A0(R4[3]), .A1(n1008), .B0(R6[3]), .B1(n1031), .C0(R5[3]), 
        .C1(n1012), .Y(n749) );
  AOI22X1 U312 ( .A0(R7[3]), .A1(n1039), .B0(data_out_1[37]), .B1(n1017), .Y(
        n748) );
  NAND2X1 U313 ( .A(n746), .B(n747), .Y(n929) );
  AOI222X1 U314 ( .A0(R4[4]), .A1(n1005), .B0(R6[4]), .B1(n1032), .C0(R5[4]), 
        .C1(n1012), .Y(n747) );
  AOI22X1 U315 ( .A0(R7[4]), .A1(n1039), .B0(data_out_1[38]), .B1(n1017), .Y(
        n746) );
  NAND2X1 U316 ( .A(n744), .B(n745), .Y(n928) );
  AOI222X1 U317 ( .A0(R4[5]), .A1(n1007), .B0(R6[5]), .B1(n1032), .C0(R5[5]), 
        .C1(n1012), .Y(n745) );
  AOI22X1 U318 ( .A0(R7[5]), .A1(n1039), .B0(data_out_1[39]), .B1(n1017), .Y(
        n744) );
  NAND2X1 U319 ( .A(n742), .B(n743), .Y(n927) );
  AOI222X1 U320 ( .A0(R4[6]), .A1(n1006), .B0(R6[6]), .B1(n1029), .C0(R5[6]), 
        .C1(n1012), .Y(n743) );
  AOI22X1 U321 ( .A0(R7[6]), .A1(n1039), .B0(data_out_1[40]), .B1(n1017), .Y(
        n742) );
  NAND2X1 U322 ( .A(n740), .B(n741), .Y(n926) );
  AOI222X1 U323 ( .A0(R4[7]), .A1(n1007), .B0(R6[7]), .B1(n1029), .C0(R5[7]), 
        .C1(n1012), .Y(n741) );
  AOI22X1 U324 ( .A0(R7[7]), .A1(n1039), .B0(data_out_1[41]), .B1(n1017), .Y(
        n740) );
  NAND2X1 U325 ( .A(n738), .B(n739), .Y(n925) );
  AOI222X1 U326 ( .A0(R4[8]), .A1(n1008), .B0(R6[8]), .B1(n1032), .C0(R5[8]), 
        .C1(n1012), .Y(n739) );
  AOI22X1 U327 ( .A0(R7[8]), .A1(n1039), .B0(data_out_1[42]), .B1(n1017), .Y(
        n738) );
  NAND2X1 U328 ( .A(n736), .B(n737), .Y(n924) );
  AOI222X1 U329 ( .A0(R4[9]), .A1(n1005), .B0(R6[9]), .B1(n1032), .C0(R5[9]), 
        .C1(n1012), .Y(n737) );
  AOI22X1 U330 ( .A0(R7[9]), .A1(n1039), .B0(data_out_1[43]), .B1(n1017), .Y(
        n736) );
  NAND2X1 U331 ( .A(n734), .B(n735), .Y(n923) );
  AOI222X1 U332 ( .A0(R4[10]), .A1(n1007), .B0(R6[10]), .B1(n1030), .C0(R5[10]), .C1(n1012), .Y(n735) );
  AOI22X1 U333 ( .A0(R7[10]), .A1(n1039), .B0(data_out_1[44]), .B1(n1017), .Y(
        n734) );
  NAND2X1 U334 ( .A(n732), .B(n733), .Y(n922) );
  AOI222X1 U335 ( .A0(R4[11]), .A1(n1006), .B0(R6[11]), .B1(n1031), .C0(R5[11]), .C1(n1012), .Y(n733) );
  AOI22X1 U336 ( .A0(R7[11]), .A1(n1039), .B0(data_out_1[45]), .B1(n1017), .Y(
        n732) );
  NAND2X1 U337 ( .A(n730), .B(n731), .Y(n921) );
  AOI222X1 U338 ( .A0(R4[12]), .A1(n1008), .B0(R6[12]), .B1(n1032), .C0(R5[12]), .C1(n1012), .Y(n731) );
  AOI22X1 U339 ( .A0(R7[12]), .A1(n1038), .B0(data_out_1[46]), .B1(n1017), .Y(
        n730) );
  NAND2X1 U340 ( .A(n728), .B(n729), .Y(n920) );
  AOI222X1 U341 ( .A0(R4[13]), .A1(n1008), .B0(R6[13]), .B1(n1031), .C0(R5[13]), .C1(n1012), .Y(n729) );
  AOI22X1 U342 ( .A0(R7[13]), .A1(n1038), .B0(data_out_1[47]), .B1(n1017), .Y(
        n728) );
  NAND2X1 U343 ( .A(n726), .B(n727), .Y(n919) );
  AOI222X1 U344 ( .A0(R4[14]), .A1(n1006), .B0(R6[14]), .B1(n1031), .C0(R5[14]), .C1(n1012), .Y(n727) );
  AOI22X1 U345 ( .A0(R7[14]), .A1(n1038), .B0(data_out_1[48]), .B1(n1018), .Y(
        n726) );
  NAND2X1 U346 ( .A(n724), .B(n725), .Y(n918) );
  AOI222X1 U347 ( .A0(R4[15]), .A1(n1006), .B0(R6[15]), .B1(n1031), .C0(R5[15]), .C1(n1013), .Y(n725) );
  AOI22X1 U348 ( .A0(R7[15]), .A1(n1038), .B0(data_out_1[49]), .B1(n1018), .Y(
        n724) );
  NAND2X1 U349 ( .A(n722), .B(n723), .Y(n917) );
  AOI222X1 U350 ( .A0(R4[16]), .A1(n1006), .B0(R6[16]), .B1(n1031), .C0(R5[16]), .C1(n1013), .Y(n723) );
  AOI22XL U351 ( .A0(R7[16]), .A1(n1038), .B0(data_out_1[50]), .B1(n1018), .Y(
        n722) );
  NAND2X1 U352 ( .A(n720), .B(n721), .Y(n916) );
  AOI222X1 U353 ( .A0(R4[17]), .A1(n1006), .B0(R6[17]), .B1(n1031), .C0(R5[17]), .C1(n1011), .Y(n721) );
  AOI22X1 U354 ( .A0(R7[17]), .A1(n1038), .B0(data_out_1[51]), .B1(n1018), .Y(
        n720) );
  NAND2X1 U355 ( .A(n718), .B(n719), .Y(n915) );
  AOI222X1 U356 ( .A0(R4[18]), .A1(n1006), .B0(R6[18]), .B1(n1031), .C0(R5[18]), .C1(n1013), .Y(n719) );
  AOI22X1 U357 ( .A0(R7[18]), .A1(n1038), .B0(data_out_1[52]), .B1(n1018), .Y(
        n718) );
  NAND2X1 U358 ( .A(n716), .B(n717), .Y(n914) );
  AOI222X1 U359 ( .A0(R4[19]), .A1(n1006), .B0(R6[19]), .B1(n1031), .C0(R5[19]), .C1(n1012), .Y(n717) );
  AOI22X1 U360 ( .A0(R7[19]), .A1(n1038), .B0(data_out_1[53]), .B1(n1018), .Y(
        n716) );
  NAND2X1 U361 ( .A(n714), .B(n715), .Y(n913) );
  AOI222X1 U362 ( .A0(R4[20]), .A1(n1006), .B0(R6[20]), .B1(n1031), .C0(R5[20]), .C1(n1013), .Y(n715) );
  AOI22X1 U363 ( .A0(R7[20]), .A1(n1038), .B0(data_out_1[54]), .B1(n1018), .Y(
        n714) );
  NAND2X1 U364 ( .A(n712), .B(n713), .Y(n912) );
  AOI222X1 U365 ( .A0(R4[21]), .A1(n1006), .B0(R6[21]), .B1(n1031), .C0(R5[21]), .C1(n1011), .Y(n713) );
  AOI22X1 U366 ( .A0(R7[21]), .A1(n1038), .B0(data_out_1[55]), .B1(n1018), .Y(
        n712) );
  NAND2X1 U367 ( .A(n710), .B(n711), .Y(n911) );
  AOI222X1 U368 ( .A0(R4[22]), .A1(n1006), .B0(R6[22]), .B1(n1031), .C0(R5[22]), .C1(n1012), .Y(n711) );
  AOI22X1 U369 ( .A0(R7[22]), .A1(n1038), .B0(data_out_1[56]), .B1(n1018), .Y(
        n710) );
  NAND2X1 U370 ( .A(n708), .B(n709), .Y(n910) );
  AOI222X1 U371 ( .A0(R4[23]), .A1(n1006), .B0(R6[23]), .B1(n1031), .C0(R5[23]), .C1(n1012), .Y(n709) );
  AOI22X1 U372 ( .A0(R7[23]), .A1(n1038), .B0(data_out_1[57]), .B1(n1018), .Y(
        n708) );
  NAND2X1 U373 ( .A(n706), .B(n707), .Y(n909) );
  AOI222X1 U374 ( .A0(R4[24]), .A1(n1006), .B0(R6[24]), .B1(n1031), .C0(R5[24]), .C1(n1013), .Y(n707) );
  AOI22X1 U375 ( .A0(R7[24]), .A1(n1037), .B0(data_out_1[58]), .B1(n1018), .Y(
        n706) );
  NAND2X1 U376 ( .A(n704), .B(n705), .Y(n908) );
  AOI222X1 U377 ( .A0(R4[25]), .A1(n1006), .B0(R6[25]), .B1(n1031), .C0(R5[25]), .C1(n1011), .Y(n705) );
  AOI22X1 U378 ( .A0(R7[25]), .A1(n1037), .B0(data_out_1[59]), .B1(n1018), .Y(
        n704) );
  NAND2X1 U379 ( .A(n702), .B(n703), .Y(n907) );
  AOI222X1 U380 ( .A0(R4[26]), .A1(n1006), .B0(R6[26]), .B1(n1031), .C0(R5[26]), .C1(n1011), .Y(n703) );
  AOI22X1 U381 ( .A0(R7[26]), .A1(n1037), .B0(data_out_1[60]), .B1(n1019), .Y(
        n702) );
  NAND2X1 U382 ( .A(n700), .B(n701), .Y(n906) );
  AOI222X1 U383 ( .A0(R4[27]), .A1(n1006), .B0(R6[27]), .B1(n1031), .C0(R5[27]), .C1(n1012), .Y(n701) );
  AOI22X1 U384 ( .A0(R7[27]), .A1(n1037), .B0(data_out_1[61]), .B1(n1019), .Y(
        n700) );
  NAND2X1 U385 ( .A(n698), .B(n699), .Y(n905) );
  AOI222X1 U386 ( .A0(R4[28]), .A1(n1006), .B0(R6[28]), .B1(n1031), .C0(R5[28]), .C1(n1013), .Y(n699) );
  AOI22X1 U387 ( .A0(R7[28]), .A1(n1037), .B0(data_out_1[62]), .B1(n1019), .Y(
        n698) );
  NAND2X1 U388 ( .A(n696), .B(n697), .Y(n904) );
  AOI222X1 U389 ( .A0(R4[29]), .A1(n1006), .B0(R6[29]), .B1(n1031), .C0(R5[29]), .C1(n1011), .Y(n697) );
  AOI22X1 U390 ( .A0(R7[29]), .A1(n1037), .B0(data_out_1[63]), .B1(n1019), .Y(
        n696) );
  NAND2X1 U391 ( .A(n694), .B(n695), .Y(n903) );
  AOI222X1 U392 ( .A0(R4[30]), .A1(n1006), .B0(R6[30]), .B1(n1030), .C0(R5[30]), .C1(n1013), .Y(n695) );
  AOI22X1 U393 ( .A0(R7[30]), .A1(n1037), .B0(data_out_1[64]), .B1(n1019), .Y(
        n694) );
  NAND2X1 U394 ( .A(n692), .B(n693), .Y(n902) );
  AOI222X1 U395 ( .A0(R4[31]), .A1(n1005), .B0(R6[31]), .B1(n1030), .C0(R5[31]), .C1(n1012), .Y(n693) );
  AOI22X1 U396 ( .A0(R7[31]), .A1(n1037), .B0(data_out_1[65]), .B1(n1019), .Y(
        n692) );
  NAND2X1 U397 ( .A(n690), .B(n691), .Y(n901) );
  AOI222X1 U398 ( .A0(R4[32]), .A1(n1005), .B0(R6[32]), .B1(n1030), .C0(R5[32]), .C1(n1011), .Y(n691) );
  AOI22X1 U399 ( .A0(R7[32]), .A1(n1037), .B0(data_out_1[66]), .B1(n1019), .Y(
        n690) );
  NAND2X1 U400 ( .A(n688), .B(n689), .Y(n900) );
  AOI222X1 U401 ( .A0(R4[33]), .A1(n1005), .B0(R6[33]), .B1(n1030), .C0(R5[33]), .C1(n1011), .Y(n689) );
  AOI22XL U402 ( .A0(R7[33]), .A1(n1037), .B0(data_out_1[67]), .B1(n1019), .Y(
        n688) );
  NAND2X1 U403 ( .A(n822), .B(n823), .Y(n967) );
  AOI222X1 U404 ( .A0(R0[0]), .A1(n1008), .B0(R2[0]), .B1(n1032), .C0(R1[0]), 
        .C1(n1012), .Y(n823) );
  NAND2X1 U405 ( .A(n820), .B(n821), .Y(n966) );
  AOI222X1 U406 ( .A0(R0[1]), .A1(n1008), .B0(R2[1]), .B1(n1032), .C0(R1[1]), 
        .C1(n1012), .Y(n821) );
  NAND2X1 U407 ( .A(n818), .B(n819), .Y(n965) );
  AOI222X1 U408 ( .A0(R0[2]), .A1(n1008), .B0(R2[2]), .B1(n1032), .C0(R1[2]), 
        .C1(n1013), .Y(n819) );
  NAND2X1 U409 ( .A(n816), .B(n817), .Y(n964) );
  AOI222X1 U410 ( .A0(R0[3]), .A1(n1008), .B0(R2[3]), .B1(n1032), .C0(R1[3]), 
        .C1(n1011), .Y(n817) );
  NAND2X1 U411 ( .A(n814), .B(n815), .Y(n963) );
  AOI222X1 U412 ( .A0(R0[4]), .A1(n1008), .B0(R2[4]), .B1(n1032), .C0(R1[4]), 
        .C1(n1013), .Y(n815) );
  AOI22X1 U413 ( .A0(R3[4]), .A1(n1042), .B0(data_out_1[4]), .B1(n1022), .Y(
        n814) );
  NAND2X1 U414 ( .A(n812), .B(n813), .Y(n962) );
  AOI222X1 U415 ( .A0(R0[5]), .A1(n1008), .B0(R2[5]), .B1(n1032), .C0(R1[5]), 
        .C1(n1011), .Y(n813) );
  NAND2X1 U416 ( .A(n810), .B(n811), .Y(n961) );
  AOI222X1 U417 ( .A0(R0[6]), .A1(n1008), .B0(R2[6]), .B1(n1032), .C0(R1[6]), 
        .C1(n1011), .Y(n811) );
  AOI22X1 U418 ( .A0(R3[6]), .A1(n1042), .B0(data_out_1[6]), .B1(n1017), .Y(
        n810) );
  NAND2X1 U419 ( .A(n808), .B(n809), .Y(n960) );
  AOI222X1 U420 ( .A0(R0[7]), .A1(n1008), .B0(R2[7]), .B1(n1032), .C0(R1[7]), 
        .C1(n1013), .Y(n809) );
  NAND2X1 U421 ( .A(n806), .B(n807), .Y(n959) );
  AOI222X1 U422 ( .A0(R0[8]), .A1(n1008), .B0(R2[8]), .B1(n1032), .C0(R1[8]), 
        .C1(n1012), .Y(n807) );
  NAND2X1 U423 ( .A(n804), .B(n805), .Y(n958) );
  AOI222X1 U424 ( .A0(R0[9]), .A1(n1008), .B0(R2[9]), .B1(n1032), .C0(R1[9]), 
        .C1(n1010), .Y(n805) );
  AOI22X1 U425 ( .A0(R3[9]), .A1(n1041), .B0(data_out_1[9]), .B1(n1023), .Y(
        n804) );
  NAND2X1 U426 ( .A(n802), .B(n803), .Y(n957) );
  AOI222X1 U427 ( .A0(R0[10]), .A1(n1008), .B0(R2[10]), .B1(n1032), .C0(R1[10]), .C1(n1011), .Y(n803) );
  AOI22X1 U428 ( .A0(R3[10]), .A1(n1041), .B0(data_out_1[10]), .B1(n1020), .Y(
        n802) );
  NAND2X1 U429 ( .A(n800), .B(n801), .Y(n956) );
  AOI222X1 U430 ( .A0(R0[11]), .A1(n1008), .B0(R2[11]), .B1(n1031), .C0(R1[11]), .C1(n1013), .Y(n801) );
  AOI22X1 U431 ( .A0(R3[11]), .A1(n1041), .B0(data_out_1[11]), .B1(n1016), .Y(
        n800) );
  NAND2X1 U432 ( .A(n798), .B(n799), .Y(n955) );
  AOI222X1 U433 ( .A0(R0[12]), .A1(n1007), .B0(R2[12]), .B1(n1031), .C0(R1[12]), .C1(n1013), .Y(n799) );
  AOI22X1 U434 ( .A0(R3[12]), .A1(n1041), .B0(data_out_1[12]), .B1(n1015), .Y(
        n798) );
  NAND2X1 U435 ( .A(n796), .B(n797), .Y(n954) );
  AOI222X1 U436 ( .A0(R0[13]), .A1(n1007), .B0(R2[13]), .B1(n1029), .C0(R1[13]), .C1(n1013), .Y(n797) );
  AOI22X1 U437 ( .A0(R3[13]), .A1(n1041), .B0(data_out_1[13]), .B1(n1015), .Y(
        n796) );
  NAND2X1 U438 ( .A(n794), .B(n795), .Y(n953) );
  AOI222X1 U439 ( .A0(R0[14]), .A1(n1007), .B0(R2[14]), .B1(n1032), .C0(R1[14]), .C1(n1013), .Y(n795) );
  AOI22X1 U440 ( .A0(R3[14]), .A1(n1041), .B0(data_out_1[14]), .B1(n1015), .Y(
        n794) );
  NAND2X1 U441 ( .A(n792), .B(n793), .Y(n952) );
  AOI222X1 U442 ( .A0(R0[15]), .A1(n1007), .B0(R2[15]), .B1(n1030), .C0(R1[15]), .C1(n1013), .Y(n793) );
  AOI22X1 U443 ( .A0(R3[15]), .A1(n1041), .B0(data_out_1[15]), .B1(n1015), .Y(
        n792) );
  NAND2X1 U444 ( .A(n790), .B(n791), .Y(n951) );
  AOI222X1 U445 ( .A0(R0[16]), .A1(n1007), .B0(R2[16]), .B1(n1031), .C0(R1[16]), .C1(n1013), .Y(n791) );
  AOI22X1 U446 ( .A0(R3[16]), .A1(n1041), .B0(data_out_1[16]), .B1(n1015), .Y(
        n790) );
  NAND2X1 U447 ( .A(n788), .B(n789), .Y(n950) );
  AOI222X1 U448 ( .A0(R0[17]), .A1(n1007), .B0(R2[17]), .B1(n1029), .C0(R1[17]), .C1(n1013), .Y(n789) );
  NAND2X1 U449 ( .A(n786), .B(n787), .Y(n949) );
  AOI222X1 U450 ( .A0(R0[18]), .A1(n1007), .B0(R2[18]), .B1(n1029), .C0(R1[18]), .C1(n1013), .Y(n787) );
  NAND2X1 U451 ( .A(n784), .B(n785), .Y(n948) );
  AOI222X1 U452 ( .A0(R0[19]), .A1(n1007), .B0(R2[19]), .B1(n1029), .C0(R1[19]), .C1(n1013), .Y(n785) );
  AOI22X1 U453 ( .A0(R3[19]), .A1(n1041), .B0(data_out_1[19]), .B1(n1015), .Y(
        n784) );
  NAND2X1 U454 ( .A(n782), .B(n783), .Y(n947) );
  AOI222X1 U455 ( .A0(R0[20]), .A1(n1007), .B0(R2[20]), .B1(n1032), .C0(R1[20]), .C1(n1013), .Y(n783) );
  AOI22X1 U456 ( .A0(R3[20]), .A1(n1040), .B0(data_out_1[20]), .B1(n1015), .Y(
        n782) );
  NAND2X1 U457 ( .A(n780), .B(n781), .Y(n946) );
  AOI222X1 U458 ( .A0(R0[21]), .A1(n1007), .B0(R2[21]), .B1(n1030), .C0(R1[21]), .C1(n1013), .Y(n781) );
  AOI22X1 U459 ( .A0(R3[21]), .A1(n1040), .B0(data_out_1[21]), .B1(n1015), .Y(
        n780) );
  NAND2X1 U460 ( .A(n778), .B(n779), .Y(n945) );
  AOI222X1 U461 ( .A0(R0[22]), .A1(n1007), .B0(R2[22]), .B1(n1031), .C0(R1[22]), .C1(n1013), .Y(n779) );
  AOI22X1 U462 ( .A0(R3[22]), .A1(n1040), .B0(data_out_1[22]), .B1(n1015), .Y(
        n778) );
  NAND2X1 U463 ( .A(n776), .B(n777), .Y(n944) );
  AOI222X1 U464 ( .A0(R0[23]), .A1(n1007), .B0(R2[23]), .B1(n1031), .C0(R1[23]), .C1(n1013), .Y(n777) );
  NAND2X1 U465 ( .A(n774), .B(n775), .Y(n943) );
  AOI222X1 U466 ( .A0(R0[24]), .A1(n1007), .B0(R2[24]), .B1(n1029), .C0(R1[24]), .C1(n1013), .Y(n775) );
  AOI22X1 U467 ( .A0(R3[24]), .A1(n1040), .B0(data_out_1[24]), .B1(n1016), .Y(
        n774) );
  NAND2X1 U468 ( .A(n772), .B(n773), .Y(n942) );
  AOI222X1 U469 ( .A0(R0[25]), .A1(n1007), .B0(R2[25]), .B1(n1032), .C0(R1[25]), .C1(n1013), .Y(n773) );
  AOI22X1 U470 ( .A0(R3[25]), .A1(n1040), .B0(data_out_1[25]), .B1(n1016), .Y(
        n772) );
  NAND2X1 U471 ( .A(n770), .B(n771), .Y(n941) );
  AOI222X1 U472 ( .A0(R0[26]), .A1(n1007), .B0(R2[26]), .B1(n1030), .C0(R1[26]), .C1(n1013), .Y(n771) );
  AOI22X1 U473 ( .A0(R3[26]), .A1(n1040), .B0(data_out_1[26]), .B1(n1016), .Y(
        n770) );
  NAND2X1 U474 ( .A(n768), .B(n769), .Y(n940) );
  AOI222X1 U475 ( .A0(R0[27]), .A1(n1007), .B0(R2[27]), .B1(n1031), .C0(R1[27]), .C1(n1013), .Y(n769) );
  AOI22X1 U476 ( .A0(R3[27]), .A1(n1040), .B0(data_out_1[27]), .B1(n1016), .Y(
        n768) );
  NAND2X1 U477 ( .A(n766), .B(n767), .Y(n939) );
  AOI222X1 U478 ( .A0(R0[28]), .A1(n1007), .B0(R2[28]), .B1(n1029), .C0(R1[28]), .C1(n1013), .Y(n767) );
  AOI22X1 U479 ( .A0(R3[28]), .A1(n1040), .B0(data_out_1[28]), .B1(n1016), .Y(
        n766) );
  NAND2X1 U480 ( .A(n764), .B(n765), .Y(n938) );
  AOI222X1 U481 ( .A0(R0[29]), .A1(n1007), .B0(R2[29]), .B1(n1032), .C0(R1[29]), .C1(n1012), .Y(n765) );
  AOI22X1 U482 ( .A0(R3[29]), .A1(n1040), .B0(data_out_1[29]), .B1(n1016), .Y(
        n764) );
  NAND2X1 U483 ( .A(n762), .B(n763), .Y(n937) );
  AOI222X1 U484 ( .A0(R0[30]), .A1(n1005), .B0(R2[30]), .B1(n1029), .C0(R1[30]), .C1(n1012), .Y(n763) );
  AOI22X1 U485 ( .A0(R3[30]), .A1(n1040), .B0(data_out_1[30]), .B1(n1016), .Y(
        n762) );
  NAND2X1 U486 ( .A(n760), .B(n761), .Y(n936) );
  AOI222X1 U487 ( .A0(R0[31]), .A1(n1007), .B0(R2[31]), .B1(n1032), .C0(R1[31]), .C1(n1012), .Y(n761) );
  AOI22X1 U488 ( .A0(R3[31]), .A1(n1040), .B0(data_out_1[31]), .B1(n1016), .Y(
        n760) );
  NAND2X1 U489 ( .A(n758), .B(n759), .Y(n935) );
  AOI222X1 U490 ( .A0(R0[32]), .A1(n1006), .B0(R2[32]), .B1(n1029), .C0(R1[32]), .C1(n1012), .Y(n759) );
  AOI22X1 U491 ( .A0(R3[32]), .A1(n1040), .B0(data_out_1[32]), .B1(n1016), .Y(
        n758) );
  NAND2X1 U492 ( .A(n756), .B(n757), .Y(n934) );
  AOI222X1 U493 ( .A0(R0[33]), .A1(n1005), .B0(R2[33]), .B1(n1030), .C0(R1[33]), .C1(n1012), .Y(n757) );
  AOI22X1 U494 ( .A0(R3[33]), .A1(n1039), .B0(data_out_1[33]), .B1(n1016), .Y(
        n756) );
  NAND2X1 U495 ( .A(counter[1]), .B(n550), .Y(n824) );
  NAND2X1 U496 ( .A(n550), .B(n1044), .Y(n828) );
  INVX1 U497 ( .A(counter[1]), .Y(n1044) );
  NAND2X1 U498 ( .A(n558), .B(n559), .Y(n835) );
  AOI222X1 U499 ( .A0(R12[30]), .A1(n1008), .B0(R14[30]), .B1(n1028), .C0(
        R13[30]), .C1(n1013), .Y(n559) );
  NAND2X1 U500 ( .A(n556), .B(n557), .Y(n834) );
  AOI222X1 U501 ( .A0(R12[31]), .A1(n1005), .B0(R14[31]), .B1(n1028), .C0(
        R13[31]), .C1(n1011), .Y(n557) );
  NAND2X1 U502 ( .A(n554), .B(n555), .Y(n833) );
  AOI222X1 U503 ( .A0(R12[32]), .A1(n1006), .B0(R14[32]), .B1(n1028), .C0(
        R13[32]), .C1(n1013), .Y(n555) );
  NAND2X1 U504 ( .A(n551), .B(n552), .Y(n832) );
  AOI222X1 U505 ( .A0(R12[33]), .A1(n1006), .B0(R14[33]), .B1(n1031), .C0(
        R13[33]), .C1(n1012), .Y(n552) );
  AOI22XL U506 ( .A0(R15[33]), .A1(n1038), .B0(data_out_1[135]), .B1(n1015), 
        .Y(n551) );
  NOR2X1 U507 ( .A(n550), .B(n1044), .Y(n831) );
endmodule


module mux ( mux_flag, clk, rst_n, data_in_1, data_in_2, data_out, 
        data_in_3_33_, data_in_3_32_, data_in_3_31_, data_in_3_30_, 
        data_in_3_29_, data_in_3_28_, data_in_3_27_, data_in_3_26_, 
        data_in_3_25_, data_in_3_24_, data_in_3_23_, data_in_3_22_, 
        data_in_3_21_, data_in_3_20_, data_in_3_19_, data_in_3_18_, 
        data_in_3_17_, data_in_3_16_, data_in_3_15_, data_in_3_14_, 
        data_in_3_13_, data_in_3_12_, data_in_3_11_, data_in_3_10_, 
        data_in_3_9_, data_in_3_8_, data_in_3_7_, data_in_3_6_, data_in_3_5_, 
        data_in_3_4_, data_in_3_3_, data_in_3_2_, data_in_3_1_, data_in_3_0_
 );
  input [135:0] data_in_1;
  input [135:0] data_in_2;
  output [135:0] data_out;
  input mux_flag, clk, rst_n, data_in_3_33_, data_in_3_32_, data_in_3_31_,
         data_in_3_30_, data_in_3_29_, data_in_3_28_, data_in_3_27_,
         data_in_3_26_, data_in_3_25_, data_in_3_24_, data_in_3_23_,
         data_in_3_22_, data_in_3_21_, data_in_3_20_, data_in_3_19_,
         data_in_3_18_, data_in_3_17_, data_in_3_16_, data_in_3_15_,
         data_in_3_14_, data_in_3_13_, data_in_3_12_, data_in_3_11_,
         data_in_3_10_, data_in_3_9_, data_in_3_8_, data_in_3_7_, data_in_3_6_,
         data_in_3_5_, data_in_3_4_, data_in_3_3_, data_in_3_2_, data_in_3_1_,
         data_in_3_0_;
  wire   n561, n562, n563, N6, N7, N8, n140, n141, n281, n282, n285, n1, n2,
         n4, n5, n6, n7, n8, n9, n10, n11, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n48, n49, n50, n51, n174, n175, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n283,
         n284, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n559, n560;
  wire   [3:1] counter;
  wire   [33:0] R4;
  wire   [33:0] R3;
  wire   [32:0] R2;
  wire   [33:0] R1;

  JKFFRX4 counter_reg_0_ ( .J(1'b1), .K(1'b1), .CK(clk), .RN(rst_n), .Q(n31), 
        .QN(n140) );
  DFFRHQX4 counter_reg_1_ ( .D(N6), .CK(clk), .RN(rst_n), .Q(counter[1]) );
  DFFRHQX4 counter_reg_2_ ( .D(N7), .CK(clk), .RN(rst_n), .Q(counter[2]) );
  DFFRHQX4 counter_reg_3_ ( .D(N8), .CK(clk), .RN(rst_n), .Q(counter[3]) );
  TLATXL R4_reg_33_ ( .G(n199), .D(data_in_3_33_), .Q(R4[33]) );
  TLATXL R3_reg_33_ ( .G(n1), .D(data_in_3_33_), .Q(R3[33]) );
  TLATXL R2_reg_33_ ( .G(n200), .D(data_in_3_33_), .Q(n11) );
  TLATXL R1_reg_33_ ( .G(n285), .D(data_in_3_33_), .Q(R1[33]) );
  TLATXL R3_reg_16_ ( .G(n1), .D(data_in_3_16_), .QN(n10) );
  TLATXL R4_reg_16_ ( .G(n199), .D(data_in_3_16_), .QN(n9) );
  TLATXL R2_reg_32_ ( .G(n200), .D(data_in_3_32_), .Q(R2[32]) );
  TLATXL R2_reg_31_ ( .G(n200), .D(data_in_3_31_), .Q(R2[31]) );
  TLATXL R2_reg_30_ ( .G(n200), .D(data_in_3_30_), .Q(R2[30]) );
  TLATXL R2_reg_29_ ( .G(n200), .D(data_in_3_29_), .Q(R2[29]) );
  TLATXL R2_reg_28_ ( .G(n200), .D(data_in_3_28_), .Q(R2[28]) );
  TLATXL R2_reg_27_ ( .G(n200), .D(data_in_3_27_), .Q(R2[27]) );
  TLATXL R2_reg_26_ ( .G(n200), .D(data_in_3_26_), .Q(R2[26]) );
  TLATXL R2_reg_25_ ( .G(n200), .D(data_in_3_25_), .Q(R2[25]) );
  TLATXL R2_reg_24_ ( .G(n200), .D(data_in_3_24_), .Q(R2[24]) );
  TLATXL R3_reg_9_ ( .G(n1), .D(data_in_3_9_), .Q(R3[9]) );
  TLATXL R3_reg_8_ ( .G(n1), .D(data_in_3_8_), .Q(R3[8]) );
  TLATXL R3_reg_7_ ( .G(n1), .D(data_in_3_7_), .Q(R3[7]) );
  TLATXL R3_reg_6_ ( .G(n1), .D(data_in_3_6_), .Q(R3[6]) );
  TLATXL R3_reg_5_ ( .G(n1), .D(data_in_3_5_), .Q(R3[5]) );
  TLATXL R3_reg_4_ ( .G(n1), .D(data_in_3_4_), .Q(R3[4]) );
  TLATXL R3_reg_3_ ( .G(n1), .D(data_in_3_3_), .Q(R3[3]) );
  TLATX1 R3_reg_2_ ( .G(n1), .D(data_in_3_2_), .Q(R3[2]) );
  TLATX1 R3_reg_1_ ( .G(n1), .D(data_in_3_1_), .Q(R3[1]) );
  TLATXL R4_reg_9_ ( .G(n199), .D(data_in_3_9_), .Q(R4[9]) );
  TLATXL R4_reg_8_ ( .G(n199), .D(data_in_3_8_), .Q(R4[8]) );
  TLATXL R4_reg_7_ ( .G(n199), .D(data_in_3_7_), .Q(R4[7]) );
  TLATXL R4_reg_6_ ( .G(n199), .D(data_in_3_6_), .Q(R4[6]) );
  TLATXL R4_reg_5_ ( .G(n199), .D(data_in_3_5_), .Q(R4[5]) );
  TLATXL R4_reg_4_ ( .G(n199), .D(data_in_3_4_), .Q(R4[4]) );
  TLATXL R4_reg_3_ ( .G(n199), .D(data_in_3_3_), .Q(R4[3]) );
  TLATX1 R4_reg_2_ ( .G(n199), .D(data_in_3_2_), .Q(R4[2]) );
  TLATX1 R4_reg_1_ ( .G(n199), .D(data_in_3_1_), .Q(R4[1]) );
  TLATXL R1_reg_5_ ( .G(n285), .D(data_in_3_5_), .Q(R1[5]) );
  TLATXL R2_reg_23_ ( .G(n200), .D(data_in_3_23_), .Q(R2[23]) );
  TLATXL R2_reg_22_ ( .G(n200), .D(data_in_3_22_), .Q(R2[22]) );
  TLATXL R2_reg_21_ ( .G(n200), .D(data_in_3_21_), .Q(R2[21]) );
  TLATX1 R2_reg_20_ ( .G(n200), .D(data_in_3_20_), .Q(R2[20]) );
  TLATX1 R2_reg_19_ ( .G(n200), .D(data_in_3_19_), .Q(R2[19]) );
  TLATXL R2_reg_16_ ( .G(n200), .D(data_in_3_16_), .Q(R2[16]) );
  TLATXL R2_reg_15_ ( .G(n200), .D(data_in_3_15_), .Q(R2[15]) );
  TLATXL R2_reg_14_ ( .G(n200), .D(data_in_3_14_), .Q(R2[14]) );
  TLATXL R2_reg_13_ ( .G(n200), .D(data_in_3_13_), .Q(R2[13]) );
  TLATXL R2_reg_12_ ( .G(n200), .D(data_in_3_12_), .Q(R2[12]) );
  TLATXL R2_reg_11_ ( .G(n200), .D(data_in_3_11_), .Q(R2[11]) );
  TLATXL R2_reg_10_ ( .G(n200), .D(data_in_3_10_), .Q(R2[10]) );
  TLATXL R2_reg_9_ ( .G(n200), .D(data_in_3_9_), .Q(R2[9]) );
  TLATXL R2_reg_8_ ( .G(n200), .D(data_in_3_8_), .Q(R2[8]) );
  TLATXL R2_reg_7_ ( .G(n200), .D(data_in_3_7_), .Q(R2[7]) );
  TLATXL R2_reg_6_ ( .G(n200), .D(data_in_3_6_), .Q(R2[6]) );
  TLATXL R2_reg_5_ ( .G(n200), .D(data_in_3_5_), .Q(R2[5]) );
  TLATXL R2_reg_4_ ( .G(n200), .D(data_in_3_4_), .Q(R2[4]) );
  TLATXL R2_reg_3_ ( .G(n200), .D(data_in_3_3_), .Q(R2[3]) );
  TLATX1 R2_reg_2_ ( .G(n200), .D(data_in_3_2_), .Q(R2[2]) );
  TLATX1 R2_reg_1_ ( .G(n200), .D(data_in_3_1_), .Q(R2[1]) );
  TLATXL R3_reg_32_ ( .G(n1), .D(data_in_3_32_), .Q(R3[32]) );
  TLATXL R3_reg_31_ ( .G(n1), .D(data_in_3_31_), .Q(R3[31]) );
  TLATXL R3_reg_30_ ( .G(n1), .D(data_in_3_30_), .Q(R3[30]) );
  TLATXL R3_reg_29_ ( .G(n1), .D(data_in_3_29_), .Q(R3[29]) );
  TLATXL R3_reg_28_ ( .G(n1), .D(data_in_3_28_), .Q(R3[28]) );
  TLATXL R3_reg_27_ ( .G(n1), .D(data_in_3_27_), .Q(R3[27]) );
  TLATXL R3_reg_26_ ( .G(n1), .D(data_in_3_26_), .Q(R3[26]) );
  TLATXL R3_reg_25_ ( .G(n1), .D(data_in_3_25_), .Q(R3[25]) );
  TLATXL R3_reg_24_ ( .G(n1), .D(data_in_3_24_), .Q(R3[24]) );
  TLATXL R3_reg_23_ ( .G(n1), .D(data_in_3_23_), .Q(R3[23]) );
  TLATXL R3_reg_22_ ( .G(n1), .D(data_in_3_22_), .Q(R3[22]) );
  TLATXL R3_reg_21_ ( .G(n1), .D(data_in_3_21_), .Q(R3[21]) );
  TLATX1 R3_reg_20_ ( .G(n1), .D(data_in_3_20_), .Q(R3[20]) );
  TLATX1 R3_reg_19_ ( .G(n1), .D(data_in_3_19_), .Q(R3[19]) );
  TLATXL R3_reg_15_ ( .G(n1), .D(data_in_3_15_), .Q(R3[15]) );
  TLATXL R3_reg_14_ ( .G(n1), .D(data_in_3_14_), .Q(R3[14]) );
  TLATXL R3_reg_13_ ( .G(n1), .D(data_in_3_13_), .Q(R3[13]) );
  TLATXL R3_reg_12_ ( .G(n1), .D(data_in_3_12_), .Q(R3[12]) );
  TLATXL R3_reg_11_ ( .G(n1), .D(data_in_3_11_), .Q(R3[11]) );
  TLATXL R3_reg_10_ ( .G(n1), .D(data_in_3_10_), .Q(R3[10]) );
  TLATXL R4_reg_32_ ( .G(n199), .D(data_in_3_32_), .Q(R4[32]) );
  TLATXL R4_reg_31_ ( .G(n199), .D(data_in_3_31_), .Q(R4[31]) );
  TLATXL R4_reg_30_ ( .G(n199), .D(data_in_3_30_), .Q(R4[30]) );
  TLATXL R4_reg_29_ ( .G(n199), .D(data_in_3_29_), .Q(R4[29]) );
  TLATXL R4_reg_28_ ( .G(n199), .D(data_in_3_28_), .Q(R4[28]) );
  TLATXL R4_reg_27_ ( .G(n199), .D(data_in_3_27_), .Q(R4[27]) );
  TLATXL R4_reg_26_ ( .G(n199), .D(data_in_3_26_), .Q(R4[26]) );
  TLATXL R4_reg_25_ ( .G(n199), .D(data_in_3_25_), .Q(R4[25]) );
  TLATXL R4_reg_24_ ( .G(n199), .D(data_in_3_24_), .Q(R4[24]) );
  TLATXL R4_reg_23_ ( .G(n199), .D(data_in_3_23_), .Q(R4[23]) );
  TLATXL R4_reg_22_ ( .G(n199), .D(data_in_3_22_), .Q(R4[22]) );
  TLATXL R4_reg_21_ ( .G(n199), .D(data_in_3_21_), .Q(R4[21]) );
  TLATX1 R4_reg_20_ ( .G(n199), .D(data_in_3_20_), .Q(R4[20]) );
  TLATX1 R4_reg_19_ ( .G(n199), .D(data_in_3_19_), .Q(R4[19]) );
  TLATXL R4_reg_15_ ( .G(n199), .D(data_in_3_15_), .Q(R4[15]) );
  TLATXL R4_reg_14_ ( .G(n199), .D(data_in_3_14_), .Q(R4[14]) );
  TLATXL R4_reg_13_ ( .G(n199), .D(data_in_3_13_), .Q(R4[13]) );
  TLATXL R4_reg_12_ ( .G(n199), .D(data_in_3_12_), .Q(R4[12]) );
  TLATXL R4_reg_11_ ( .G(n199), .D(data_in_3_11_), .Q(R4[11]) );
  TLATXL R4_reg_10_ ( .G(n199), .D(data_in_3_10_), .Q(R4[10]) );
  TLATXL R1_reg_32_ ( .G(n197), .D(data_in_3_32_), .Q(R1[32]) );
  TLATXL R1_reg_31_ ( .G(n285), .D(data_in_3_31_), .Q(R1[31]) );
  TLATXL R1_reg_30_ ( .G(n197), .D(data_in_3_30_), .Q(R1[30]) );
  TLATXL R1_reg_29_ ( .G(n285), .D(data_in_3_29_), .Q(R1[29]) );
  TLATXL R1_reg_28_ ( .G(n285), .D(data_in_3_28_), .Q(R1[28]) );
  TLATXL R1_reg_27_ ( .G(n285), .D(data_in_3_27_), .Q(R1[27]) );
  TLATXL R1_reg_26_ ( .G(n285), .D(data_in_3_26_), .Q(R1[26]) );
  TLATXL R1_reg_25_ ( .G(n285), .D(data_in_3_25_), .Q(R1[25]) );
  TLATXL R1_reg_24_ ( .G(n285), .D(data_in_3_24_), .Q(R1[24]) );
  TLATXL R1_reg_23_ ( .G(n197), .D(data_in_3_23_), .Q(R1[23]) );
  TLATXL R1_reg_22_ ( .G(n197), .D(data_in_3_22_), .Q(R1[22]) );
  TLATXL R1_reg_21_ ( .G(n197), .D(data_in_3_21_), .Q(R1[21]) );
  TLATX1 R1_reg_20_ ( .G(n197), .D(data_in_3_20_), .Q(R1[20]) );
  TLATX1 R1_reg_19_ ( .G(n197), .D(data_in_3_19_), .Q(R1[19]) );
  TLATX1 R1_reg_18_ ( .G(n197), .D(data_in_3_18_), .Q(R1[18]) );
  TLATXL R1_reg_16_ ( .G(n197), .D(data_in_3_16_), .Q(R1[16]) );
  TLATXL R1_reg_15_ ( .G(n197), .D(data_in_3_15_), .Q(R1[15]) );
  TLATXL R1_reg_14_ ( .G(n197), .D(data_in_3_14_), .Q(R1[14]) );
  TLATXL R1_reg_13_ ( .G(n197), .D(data_in_3_13_), .Q(R1[13]) );
  TLATXL R1_reg_12_ ( .G(n197), .D(data_in_3_12_), .Q(R1[12]) );
  TLATXL R1_reg_11_ ( .G(n285), .D(data_in_3_11_), .Q(R1[11]) );
  TLATXL R1_reg_10_ ( .G(n285), .D(data_in_3_10_), .Q(R1[10]) );
  TLATXL R1_reg_9_ ( .G(n285), .D(data_in_3_9_), .Q(R1[9]) );
  TLATXL R1_reg_8_ ( .G(n285), .D(data_in_3_8_), .Q(R1[8]) );
  TLATXL R1_reg_7_ ( .G(n285), .D(data_in_3_7_), .Q(R1[7]) );
  TLATXL R1_reg_6_ ( .G(n285), .D(data_in_3_6_), .Q(R1[6]) );
  TLATXL R1_reg_4_ ( .G(n285), .D(data_in_3_4_), .Q(R1[4]) );
  TLATXL R1_reg_3_ ( .G(n285), .D(data_in_3_3_), .Q(R1[3]) );
  TLATX1 R1_reg_2_ ( .G(n285), .D(data_in_3_2_), .Q(R1[2]) );
  TLATX1 R1_reg_1_ ( .G(n285), .D(data_in_3_1_), .Q(R1[1]) );
  TLATXL R3_reg_18_ ( .G(n1), .D(data_in_3_18_), .Q(R3[18]) );
  TLATXL R2_reg_18_ ( .G(n200), .D(data_in_3_18_), .Q(R2[18]) );
  TLATXL R4_reg_18_ ( .G(n199), .D(data_in_3_18_), .Q(R4[18]) );
  TLATXL R1_reg_0_ ( .G(n285), .D(data_in_3_0_), .Q(R1[0]) );
  TLATXL R2_reg_17_ ( .G(n200), .D(data_in_3_17_), .Q(R2[17]) );
  TLATXL R2_reg_0_ ( .G(n200), .D(data_in_3_0_), .Q(R2[0]) );
  TLATXL R3_reg_17_ ( .G(n1), .D(data_in_3_17_), .Q(R3[17]) );
  TLATXL R3_reg_0_ ( .G(n1), .D(data_in_3_0_), .Q(R3[0]) );
  TLATXL R4_reg_17_ ( .G(n199), .D(data_in_3_17_), .Q(R4[17]) );
  TLATXL R4_reg_0_ ( .G(n199), .D(data_in_3_0_), .Q(R4[0]) );
  TLATXL R1_reg_17_ ( .G(n197), .D(data_in_3_17_), .Q(R1[17]) );
  AOI22X2 U4 ( .A0(data_in_1[17]), .A1(n185), .B0(R1[17]), .B1(n193), .Y(n230)
         );
  BUFX16 U5 ( .A(counter[3]), .Y(n174) );
  NAND2BX2 U6 ( .AN(n555), .B(R4[33]), .Y(n32) );
  NAND3X1 U7 ( .A(n555), .B(n19), .C(data_in_1[135]), .Y(n554) );
  CLKINVX3 U8 ( .A(data_in_2[101]), .Y(n452) );
  MXI2X4 U9 ( .A(n7), .B(R3[33]), .S0(n556), .Y(n15) );
  NOR4BX4 U10 ( .AN(n26), .B(n559), .C(n560), .D(n23), .Y(n285) );
  CLKINVX3 U11 ( .A(n4), .Y(n200) );
  NOR2X4 U12 ( .A(n24), .B(n141), .Y(n1) );
  CLKINVX3 U13 ( .A(n5), .Y(n199) );
  CLKINVX4 U14 ( .A(n549), .Y(n188) );
  INVX20 U15 ( .A(n211), .Y(n549) );
  INVX4 U16 ( .A(n188), .Y(n183) );
  INVX4 U17 ( .A(n196), .Y(n194) );
  INVX4 U18 ( .A(n196), .Y(n192) );
  INVX4 U19 ( .A(n182), .Y(n180) );
  INVX12 U20 ( .A(n246), .Y(n181) );
  OAI2BB1X1 U21 ( .A0N(data_in_2[20]), .A1N(n181), .B0(n233), .Y(data_out[20])
         );
  INVX4 U22 ( .A(n19), .Y(n2) );
  CLKINVX4 U23 ( .A(n34), .Y(n19) );
  OR2X2 U24 ( .A(n21), .B(n20), .Y(n201) );
  OR2XL U25 ( .A(n452), .B(n179), .Y(n29) );
  BUFX16 U26 ( .A(mux_flag), .Y(n179) );
  NAND2X2 U27 ( .A(data_in_1[118]), .B(n179), .Y(n500) );
  INVX4 U28 ( .A(n27), .Y(n28) );
  NAND2X2 U29 ( .A(data_in_2[50]), .B(n34), .Y(n27) );
  INVX8 U30 ( .A(n179), .Y(n34) );
  CLKINVXL U31 ( .A(n246), .Y(n216) );
  INVX16 U32 ( .A(n50), .Y(n246) );
  BUFX8 U33 ( .A(n563), .Y(data_out[1]) );
  OAI2BB1X1 U34 ( .A0N(data_in_2[1]), .A1N(n181), .B0(n203), .Y(n563) );
  CLKINVX8 U35 ( .A(n550), .Y(n196) );
  CLKINVX8 U36 ( .A(n196), .Y(n195) );
  INVX8 U37 ( .A(n196), .Y(n193) );
  INVX4 U38 ( .A(n196), .Y(n190) );
  AOI22XL U39 ( .A0(data_in_1[29]), .A1(n184), .B0(R1[29]), .B1(n192), .Y(n249) );
  AOI22XL U40 ( .A0(data_in_1[30]), .A1(n185), .B0(R1[30]), .B1(n194), .Y(n250) );
  AOI22X2 U41 ( .A0(data_in_1[18]), .A1(n549), .B0(R1[18]), .B1(n550), .Y(n231) );
  OAI2BB1X2 U42 ( .A0N(data_in_2[25]), .A1N(n181), .B0(n241), .Y(data_out[25])
         );
  INVX4 U43 ( .A(n189), .Y(n184) );
  INVX8 U44 ( .A(n189), .Y(n186) );
  INVX4 U45 ( .A(n196), .Y(n191) );
  OR3XL U46 ( .A(n26), .B(n33), .C(n17), .Y(n141) );
  BUFX3 U47 ( .A(n23), .Y(n24) );
  CLKINVX8 U48 ( .A(n549), .Y(n189) );
  OR3XL U49 ( .A(n282), .B(n559), .C(n560), .Y(n4) );
  OR2XL U50 ( .A(n504), .B(n141), .Y(n5) );
  OR2XL U51 ( .A(n179), .B(n30), .Y(n6) );
  AND2X1 U52 ( .A(data_in_1[101]), .B(n179), .Y(n7) );
  AND2X2 U53 ( .A(data_in_1[50]), .B(n179), .Y(n8) );
  OAI2BB1X2 U54 ( .A0N(data_in_2[9]), .A1N(n221), .B0(n220), .Y(data_out[9])
         );
  OAI2BB1X2 U55 ( .A0N(data_in_2[13]), .A1N(n235), .B0(n226), .Y(data_out[13])
         );
  BUFX3 U56 ( .A(n562), .Y(data_out[31]) );
  OR2X4 U57 ( .A(n179), .B(n501), .Y(n13) );
  NAND2X4 U58 ( .A(n13), .B(n500), .Y(n502) );
  INVX1 U59 ( .A(data_in_2[118]), .Y(n501) );
  NAND3X4 U60 ( .A(n14), .B(n32), .C(n554), .Y(n561) );
  OR2X4 U61 ( .A(n556), .B(n6), .Y(n14) );
  NAND2X2 U62 ( .A(n556), .B(n11), .Y(n48) );
  NAND2X4 U63 ( .A(n15), .B(n49), .Y(data_out[101]) );
  NAND3X4 U64 ( .A(n48), .B(n352), .C(n353), .Y(data_out[67]) );
  OAI2BB1X4 U65 ( .A0N(R2[16]), .A1N(n16), .B0(n51), .Y(data_out[50]) );
  CLKINVX1 U66 ( .A(n351), .Y(n16) );
  OAI2BB1X4 U67 ( .A0N(data_in_2[27]), .A1N(n245), .B0(n244), .Y(data_out[27])
         );
  OAI21X4 U68 ( .A0(n20), .A1(n21), .B0(n502), .Y(n503) );
  DLY1X1 U69 ( .A(n174), .Y(n17) );
  BUFX12 U70 ( .A(counter[2]), .Y(n18) );
  INVXL U71 ( .A(n504), .Y(n23) );
  NOR2X4 U72 ( .A(n403), .B(n9), .Y(n505) );
  XOR2XL U73 ( .A(n26), .B(n23), .Y(N6) );
  AOI22X2 U74 ( .A0(data_in_1[20]), .A1(n549), .B0(R1[20]), .B1(n195), .Y(n233) );
  CLKBUFX8 U75 ( .A(counter[1]), .Y(n175) );
  CLKINVX8 U76 ( .A(n504), .Y(n20) );
  INVX8 U77 ( .A(n31), .Y(n504) );
  NAND2X4 U78 ( .A(n499), .B(n175), .Y(n21) );
  OAI2BB1X2 U79 ( .A0N(data_in_2[29]), .A1N(n221), .B0(n249), .Y(data_out[29])
         );
  AND2X2 U80 ( .A(data_in_1[67]), .B(n179), .Y(n22) );
  NAND3X2 U81 ( .A(n351), .B(n2), .C(data_in_2[67]), .Y(n353) );
  AOI22X1 U82 ( .A0(data_in_1[3]), .A1(n186), .B0(R1[3]), .B1(n195), .Y(n206)
         );
  NAND2X2 U83 ( .A(data_in_1[84]), .B(n179), .Y(n401) );
  OAI2BB1X2 U84 ( .A0N(data_in_2[30]), .A1N(n205), .B0(n250), .Y(data_out[30])
         );
  OAI2BB1X2 U85 ( .A0N(data_in_2[12]), .A1N(n245), .B0(n225), .Y(data_out[12])
         );
  OAI2BB1X4 U86 ( .A0N(data_in_2[7]), .A1N(n181), .B0(n217), .Y(data_out[7])
         );
  OAI2BB1X2 U87 ( .A0N(data_in_2[11]), .A1N(n224), .B0(n223), .Y(data_out[11])
         );
  NOR2BX1 U88 ( .AN(n201), .B(n19), .Y(n50) );
  NAND2X2 U89 ( .A(n351), .B(n22), .Y(n352) );
  INVX1 U90 ( .A(data_in_2[135]), .Y(n30) );
  OAI2BB1X2 U91 ( .A0N(data_in_2[10]), .A1N(n224), .B0(n222), .Y(data_out[10])
         );
  BUFX20 U92 ( .A(n561), .Y(data_out[135]) );
  OR2X4 U93 ( .A(n556), .B(n29), .Y(n49) );
  DLY1X1 U94 ( .A(n175), .Y(n26) );
  NAND2X2 U95 ( .A(n351), .B(n28), .Y(n304) );
  INVX8 U96 ( .A(n189), .Y(n185) );
  INVX1 U97 ( .A(n559), .Y(n33) );
  NOR2X4 U98 ( .A(n403), .B(n10), .Y(n405) );
  OAI21X4 U99 ( .A0(n21), .A1(n20), .B0(n402), .Y(n404) );
  AOI22X4 U100 ( .A0(data_in_1[0]), .A1(n186), .B0(R1[0]), .B1(n193), .Y(n202)
         );
  NAND2X2 U101 ( .A(n351), .B(n8), .Y(n303) );
  AND2X4 U102 ( .A(n303), .B(n304), .Y(n51) );
  OAI2BB1X4 U103 ( .A0N(data_in_2[23]), .A1N(n181), .B0(n238), .Y(data_out[23]) );
  INVX12 U104 ( .A(n188), .Y(n187) );
  INVX12 U105 ( .A(n201), .Y(n550) );
  NOR3BX4 U106 ( .AN(counter[1]), .B(n18), .C(n174), .Y(n35) );
  CLKINVX8 U107 ( .A(n140), .Y(n36) );
  INVXL U108 ( .A(n235), .Y(n182) );
  NAND2XL U109 ( .A(n19), .B(n201), .Y(n211) );
  AOI22XL U110 ( .A0(data_in_1[28]), .A1(n187), .B0(R1[28]), .B1(n190), .Y(
        n247) );
  AOI22XL U111 ( .A0(data_in_1[31]), .A1(n185), .B0(R1[31]), .B1(n195), .Y(
        n251) );
  INVX1 U112 ( .A(n198), .Y(n197) );
  INVX1 U113 ( .A(n285), .Y(n198) );
  XOR2X1 U114 ( .A(n559), .B(n282), .Y(N7) );
  XOR2X1 U115 ( .A(n17), .B(n281), .Y(N8) );
  NOR2X1 U116 ( .A(n559), .B(n282), .Y(n281) );
  INVXL U117 ( .A(n17), .Y(n560) );
  INVXL U118 ( .A(n246), .Y(n207) );
  OAI2BB1X4 U119 ( .A0N(data_in_2[84]), .A1N(n34), .B0(n401), .Y(n402) );
  INVXL U120 ( .A(n246), .Y(n209) );
  AOI22XL U121 ( .A0(data_in_1[4]), .A1(n183), .B0(R1[4]), .B1(n194), .Y(n208)
         );
  INVXL U122 ( .A(n246), .Y(n235) );
  AOI22XL U123 ( .A0(data_in_1[21]), .A1(n187), .B0(R1[21]), .B1(n192), .Y(
        n234) );
  INVXL U124 ( .A(n246), .Y(n248) );
  INVXL U125 ( .A(n246), .Y(n240) );
  AOI22XL U126 ( .A0(data_in_1[24]), .A1(n186), .B0(R1[24]), .B1(n190), .Y(
        n239) );
  AOI22X1 U127 ( .A0(data_in_1[1]), .A1(n185), .B0(R1[1]), .B1(n195), .Y(n203)
         );
  INVXL U128 ( .A(n246), .Y(n237) );
  AOI22XL U129 ( .A0(data_in_1[22]), .A1(n184), .B0(R1[22]), .B1(n194), .Y(
        n236) );
  AOI22XL U130 ( .A0(data_in_1[6]), .A1(n184), .B0(R1[6]), .B1(n191), .Y(n215)
         );
  INVXL U131 ( .A(n246), .Y(n205) );
  AOI22X2 U132 ( .A0(data_in_1[2]), .A1(n185), .B0(R1[2]), .B1(n194), .Y(n204)
         );
  AOI22XL U133 ( .A0(data_in_1[7]), .A1(n183), .B0(R1[7]), .B1(n190), .Y(n217)
         );
  INVXL U134 ( .A(n246), .Y(n221) );
  AOI22XL U135 ( .A0(data_in_1[9]), .A1(n185), .B0(R1[9]), .B1(n550), .Y(n220)
         );
  INVXL U136 ( .A(n246), .Y(n243) );
  AOI22XL U137 ( .A0(data_in_1[26]), .A1(n187), .B0(R1[26]), .B1(n192), .Y(
        n242) );
  INVXL U138 ( .A(n246), .Y(n219) );
  AOI22XL U139 ( .A0(data_in_1[8]), .A1(n183), .B0(R1[8]), .B1(n193), .Y(n218)
         );
  INVXL U140 ( .A(n246), .Y(n245) );
  AOI22XL U141 ( .A0(data_in_1[27]), .A1(n187), .B0(R1[27]), .B1(n192), .Y(
        n244) );
  AOI22XL U142 ( .A0(data_in_1[13]), .A1(n186), .B0(R1[13]), .B1(n193), .Y(
        n226) );
  AOI22XL U143 ( .A0(data_in_1[25]), .A1(n185), .B0(R1[25]), .B1(n193), .Y(
        n241) );
  AOI22XL U144 ( .A0(data_in_1[10]), .A1(n187), .B0(R1[10]), .B1(n190), .Y(
        n222) );
  OAI2BB1X1 U145 ( .A0N(data_in_2[15]), .A1N(n216), .B0(n228), .Y(data_out[15]) );
  AOI22XL U146 ( .A0(data_in_1[15]), .A1(n186), .B0(R1[15]), .B1(n194), .Y(
        n228) );
  AOI22XL U147 ( .A0(data_in_1[12]), .A1(n187), .B0(R1[12]), .B1(n191), .Y(
        n225) );
  OAI2BB1X1 U148 ( .A0N(data_in_2[32]), .A1N(n209), .B0(n252), .Y(data_out[32]) );
  AOI22XL U149 ( .A0(data_in_1[32]), .A1(n184), .B0(R1[32]), .B1(n190), .Y(
        n252) );
  OAI2BB1X1 U150 ( .A0N(data_in_2[31]), .A1N(n243), .B0(n251), .Y(n562) );
  OAI2BB1X1 U151 ( .A0N(data_in_2[14]), .A1N(n181), .B0(n227), .Y(data_out[14]) );
  AOI22XL U152 ( .A0(data_in_1[14]), .A1(n549), .B0(R1[14]), .B1(n195), .Y(
        n227) );
  AOI22XL U153 ( .A0(data_in_1[23]), .A1(n184), .B0(R1[23]), .B1(n192), .Y(
        n238) );
  INVXL U154 ( .A(n246), .Y(n224) );
  AOI22XL U155 ( .A0(data_in_1[11]), .A1(n185), .B0(R1[11]), .B1(n190), .Y(
        n223) );
  OAI22XL U156 ( .A0(n246), .A1(n212), .B0(n188), .B1(n210), .Y(n214) );
  OAI2BB1X1 U157 ( .A0N(data_in_2[33]), .A1N(n248), .B0(n253), .Y(data_out[33]) );
  AOI22XL U158 ( .A0(data_in_1[33]), .A1(n183), .B0(R1[33]), .B1(n550), .Y(
        n253) );
  OAI2BB1X1 U159 ( .A0N(data_in_2[16]), .A1N(n219), .B0(n229), .Y(data_out[16]) );
  AOI22XL U160 ( .A0(data_in_1[16]), .A1(n549), .B0(R1[16]), .B1(n191), .Y(
        n229) );
  INVX1 U161 ( .A(data_in_2[5]), .Y(n212) );
  INVX1 U162 ( .A(data_in_1[5]), .Y(n210) );
  INVXL U163 ( .A(n18), .Y(n559) );
  OAI2BB1X1 U164 ( .A0N(data_in_2[51]), .A1N(n248), .B0(n305), .Y(data_out[51]) );
  AOI22XL U165 ( .A0(data_in_1[51]), .A1(n183), .B0(R2[17]), .B1(n194), .Y(
        n305) );
  OAI2BB1X1 U166 ( .A0N(data_in_2[119]), .A1N(n240), .B0(n506), .Y(
        data_out[119]) );
  AOI22XL U167 ( .A0(data_in_1[119]), .A1(n187), .B0(R4[17]), .B1(n190), .Y(
        n506) );
  OAI2BB1X1 U168 ( .A0N(data_in_2[102]), .A1N(n181), .B0(n453), .Y(
        data_out[102]) );
  AOI22XL U169 ( .A0(data_in_1[102]), .A1(n187), .B0(R4[0]), .B1(n193), .Y(
        n453) );
  NAND3X1 U170 ( .A(n308), .B(n307), .C(n306), .Y(data_out[52]) );
  NAND2X1 U171 ( .A(data_in_1[52]), .B(n185), .Y(n307) );
  NAND2X1 U172 ( .A(data_in_2[52]), .B(n216), .Y(n308) );
  NAND2X1 U173 ( .A(R2[18]), .B(n550), .Y(n306) );
  NAND3X1 U174 ( .A(n509), .B(n508), .C(n507), .Y(data_out[120]) );
  NAND2X1 U175 ( .A(data_in_1[120]), .B(n187), .Y(n508) );
  NAND2X1 U176 ( .A(data_in_2[120]), .B(n180), .Y(n509) );
  NAND2X1 U177 ( .A(R4[18]), .B(n194), .Y(n507) );
  NAND3X1 U178 ( .A(n456), .B(n455), .C(n454), .Y(data_out[103]) );
  NAND2X1 U179 ( .A(data_in_1[103]), .B(n183), .Y(n455) );
  NAND2X1 U180 ( .A(data_in_2[103]), .B(n180), .Y(n456) );
  NAND2X1 U181 ( .A(R4[1]), .B(n550), .Y(n454) );
  NAND3X1 U182 ( .A(n311), .B(n310), .C(n309), .Y(data_out[53]) );
  NAND2X1 U183 ( .A(data_in_1[53]), .B(n549), .Y(n310) );
  NAND2X1 U184 ( .A(data_in_2[53]), .B(n209), .Y(n311) );
  NAND2X1 U185 ( .A(R2[19]), .B(n192), .Y(n309) );
  NAND3X1 U186 ( .A(n512), .B(n511), .C(n510), .Y(data_out[121]) );
  NAND2X1 U187 ( .A(data_in_1[121]), .B(n187), .Y(n511) );
  NAND2X1 U188 ( .A(data_in_2[121]), .B(n180), .Y(n512) );
  NAND2X1 U189 ( .A(R4[19]), .B(n191), .Y(n510) );
  NAND3X1 U190 ( .A(n459), .B(n458), .C(n457), .Y(data_out[104]) );
  NAND2X1 U191 ( .A(data_in_1[104]), .B(n187), .Y(n458) );
  NAND2X1 U192 ( .A(data_in_2[104]), .B(n180), .Y(n459) );
  NAND2X1 U193 ( .A(R4[2]), .B(n193), .Y(n457) );
  NAND3X1 U194 ( .A(n314), .B(n313), .C(n312), .Y(data_out[54]) );
  NAND2X1 U195 ( .A(data_in_1[54]), .B(n187), .Y(n313) );
  NAND2X1 U196 ( .A(data_in_2[54]), .B(n221), .Y(n314) );
  NAND2X1 U197 ( .A(R2[20]), .B(n191), .Y(n312) );
  NAND3X1 U198 ( .A(n263), .B(n262), .C(n261), .Y(data_out[37]) );
  NAND2X1 U199 ( .A(data_in_1[37]), .B(n183), .Y(n262) );
  NAND2X1 U200 ( .A(R2[3]), .B(n191), .Y(n261) );
  NAND2X1 U201 ( .A(data_in_2[37]), .B(n219), .Y(n263) );
  NAND3X1 U202 ( .A(n415), .B(n414), .C(n413), .Y(data_out[88]) );
  NAND2X1 U203 ( .A(data_in_1[88]), .B(n549), .Y(n414) );
  NAND2X1 U204 ( .A(data_in_2[88]), .B(n237), .Y(n415) );
  NAND2X1 U205 ( .A(R3[20]), .B(n193), .Y(n413) );
  NAND3X1 U206 ( .A(n364), .B(n363), .C(n362), .Y(data_out[71]) );
  NAND2X1 U207 ( .A(data_in_1[71]), .B(n187), .Y(n363) );
  NAND2X1 U208 ( .A(data_in_2[71]), .B(n240), .Y(n364) );
  NAND2X1 U209 ( .A(R3[3]), .B(n192), .Y(n362) );
  NAND3X1 U210 ( .A(n515), .B(n514), .C(n513), .Y(data_out[122]) );
  NAND2X1 U211 ( .A(data_in_1[122]), .B(n187), .Y(n514) );
  NAND2X1 U212 ( .A(data_in_2[122]), .B(n180), .Y(n515) );
  NAND2X1 U213 ( .A(R4[20]), .B(n193), .Y(n513) );
  NAND3X1 U214 ( .A(n462), .B(n461), .C(n460), .Y(data_out[105]) );
  NAND2X1 U215 ( .A(data_in_1[105]), .B(n186), .Y(n461) );
  NAND2X1 U216 ( .A(data_in_2[105]), .B(n180), .Y(n462) );
  NAND2X1 U217 ( .A(R4[3]), .B(n190), .Y(n460) );
  NAND3X1 U218 ( .A(n418), .B(n417), .C(n416), .Y(data_out[89]) );
  NAND2X1 U219 ( .A(data_in_1[89]), .B(n187), .Y(n417) );
  NAND2X1 U220 ( .A(data_in_2[89]), .B(n245), .Y(n418) );
  NAND2X1 U221 ( .A(R3[21]), .B(n191), .Y(n416) );
  NAND3X1 U222 ( .A(n367), .B(n366), .C(n365), .Y(data_out[72]) );
  NAND2X1 U223 ( .A(data_in_1[72]), .B(n184), .Y(n366) );
  NAND2X1 U224 ( .A(data_in_2[72]), .B(n180), .Y(n367) );
  NAND2X1 U225 ( .A(R3[4]), .B(n550), .Y(n365) );
  NAND3X1 U226 ( .A(n518), .B(n517), .C(n516), .Y(data_out[123]) );
  NAND2X1 U227 ( .A(data_in_1[123]), .B(n184), .Y(n517) );
  NAND2X1 U228 ( .A(data_in_2[123]), .B(n180), .Y(n518) );
  NAND2X1 U229 ( .A(R4[21]), .B(n190), .Y(n516) );
  NAND3X1 U230 ( .A(n465), .B(n464), .C(n463), .Y(data_out[106]) );
  NAND2X1 U231 ( .A(data_in_1[106]), .B(n185), .Y(n464) );
  NAND2X1 U232 ( .A(data_in_2[106]), .B(n180), .Y(n465) );
  NAND2X1 U233 ( .A(R4[4]), .B(n193), .Y(n463) );
  NAND3X1 U234 ( .A(n269), .B(n268), .C(n267), .Y(data_out[39]) );
  NAND2X1 U235 ( .A(data_in_1[39]), .B(n549), .Y(n268) );
  NAND2X1 U236 ( .A(R2[5]), .B(n193), .Y(n267) );
  NAND2X1 U237 ( .A(data_in_2[39]), .B(n180), .Y(n269) );
  NAND3X1 U238 ( .A(n421), .B(n420), .C(n419), .Y(data_out[90]) );
  NAND2X1 U239 ( .A(data_in_1[90]), .B(n184), .Y(n420) );
  NAND2X1 U240 ( .A(data_in_2[90]), .B(n224), .Y(n421) );
  NAND2X1 U241 ( .A(R3[22]), .B(n192), .Y(n419) );
  NAND3X1 U242 ( .A(n370), .B(n369), .C(n368), .Y(data_out[73]) );
  NAND2X1 U243 ( .A(data_in_1[73]), .B(n183), .Y(n369) );
  NAND2X1 U244 ( .A(data_in_2[73]), .B(n245), .Y(n370) );
  NAND2X1 U245 ( .A(R3[5]), .B(n192), .Y(n368) );
  NAND3X1 U246 ( .A(n521), .B(n520), .C(n519), .Y(data_out[124]) );
  NAND2X1 U247 ( .A(data_in_1[124]), .B(n183), .Y(n520) );
  NAND2XL U248 ( .A(R4[22]), .B(n193), .Y(n519) );
  NAND2X1 U249 ( .A(data_in_2[124]), .B(n180), .Y(n521) );
  NAND3X1 U250 ( .A(n468), .B(n467), .C(n466), .Y(data_out[107]) );
  NAND2X1 U251 ( .A(data_in_1[107]), .B(n187), .Y(n467) );
  NAND2X1 U252 ( .A(data_in_2[107]), .B(n180), .Y(n468) );
  NAND2X1 U253 ( .A(R4[5]), .B(n550), .Y(n466) );
  NAND3X1 U254 ( .A(n323), .B(n322), .C(n321), .Y(data_out[57]) );
  NAND2X1 U255 ( .A(data_in_1[57]), .B(n187), .Y(n322) );
  NAND2X1 U256 ( .A(data_in_2[57]), .B(n205), .Y(n323) );
  NAND2X1 U257 ( .A(R2[23]), .B(n190), .Y(n321) );
  NAND3X1 U258 ( .A(n272), .B(n271), .C(n270), .Y(data_out[40]) );
  NAND2X1 U259 ( .A(data_in_1[40]), .B(n185), .Y(n271) );
  NAND2X1 U260 ( .A(R2[6]), .B(n193), .Y(n270) );
  NAND2X1 U261 ( .A(data_in_2[40]), .B(n180), .Y(n272) );
  NAND3X1 U262 ( .A(n424), .B(n423), .C(n422), .Y(data_out[91]) );
  NAND2X1 U263 ( .A(data_in_1[91]), .B(n183), .Y(n423) );
  NAND2X1 U264 ( .A(data_in_2[91]), .B(n180), .Y(n424) );
  NAND2X1 U265 ( .A(R3[23]), .B(n192), .Y(n422) );
  NAND3X1 U266 ( .A(n373), .B(n372), .C(n371), .Y(data_out[74]) );
  NAND2X1 U267 ( .A(data_in_1[74]), .B(n187), .Y(n372) );
  NAND2X1 U268 ( .A(data_in_2[74]), .B(n180), .Y(n373) );
  NAND2X1 U269 ( .A(R3[6]), .B(n195), .Y(n371) );
  NAND3X1 U270 ( .A(n524), .B(n523), .C(n522), .Y(data_out[125]) );
  NAND2X1 U271 ( .A(data_in_1[125]), .B(n549), .Y(n523) );
  NAND2X1 U272 ( .A(data_in_2[125]), .B(n180), .Y(n524) );
  NAND2X1 U273 ( .A(R4[23]), .B(n193), .Y(n522) );
  NAND3X1 U274 ( .A(n471), .B(n470), .C(n469), .Y(data_out[108]) );
  NAND2X1 U275 ( .A(data_in_1[108]), .B(n187), .Y(n470) );
  NAND2X1 U276 ( .A(data_in_2[108]), .B(n180), .Y(n471) );
  NAND2X1 U277 ( .A(R4[6]), .B(n192), .Y(n469) );
  NAND3X1 U278 ( .A(n326), .B(n325), .C(n324), .Y(data_out[58]) );
  NAND2X1 U279 ( .A(data_in_1[58]), .B(n549), .Y(n325) );
  NAND2X1 U280 ( .A(data_in_2[58]), .B(n224), .Y(n326) );
  NAND2X1 U281 ( .A(R2[24]), .B(n190), .Y(n324) );
  NAND3X1 U282 ( .A(n275), .B(n274), .C(n273), .Y(data_out[41]) );
  NAND2X1 U283 ( .A(data_in_1[41]), .B(n186), .Y(n274) );
  NAND2X1 U284 ( .A(R2[7]), .B(n191), .Y(n273) );
  NAND2X1 U285 ( .A(data_in_2[41]), .B(n180), .Y(n275) );
  NAND3X1 U286 ( .A(n427), .B(n426), .C(n425), .Y(data_out[92]) );
  NAND2X1 U287 ( .A(data_in_1[92]), .B(n549), .Y(n426) );
  NAND2X1 U288 ( .A(data_in_2[92]), .B(n180), .Y(n427) );
  NAND2X1 U289 ( .A(R3[24]), .B(n191), .Y(n425) );
  NAND3X1 U290 ( .A(n376), .B(n375), .C(n374), .Y(data_out[75]) );
  NAND2X1 U291 ( .A(data_in_1[75]), .B(n185), .Y(n375) );
  NAND2X1 U292 ( .A(data_in_2[75]), .B(n180), .Y(n376) );
  NAND2X1 U293 ( .A(R3[7]), .B(n192), .Y(n374) );
  NAND3X1 U294 ( .A(n527), .B(n526), .C(n525), .Y(data_out[126]) );
  NAND2X1 U295 ( .A(data_in_1[126]), .B(n187), .Y(n526) );
  NAND2XL U296 ( .A(R4[24]), .B(n195), .Y(n525) );
  NAND2X1 U297 ( .A(data_in_2[126]), .B(n180), .Y(n527) );
  NAND3X1 U298 ( .A(n474), .B(n473), .C(n472), .Y(data_out[109]) );
  NAND2X1 U299 ( .A(data_in_1[109]), .B(n187), .Y(n473) );
  NAND2X1 U300 ( .A(data_in_2[109]), .B(n180), .Y(n474) );
  NAND2X1 U301 ( .A(R4[7]), .B(n194), .Y(n472) );
  NAND3X1 U302 ( .A(n329), .B(n328), .C(n327), .Y(data_out[59]) );
  NAND2X1 U303 ( .A(data_in_1[59]), .B(n187), .Y(n328) );
  NAND2X1 U304 ( .A(data_in_2[59]), .B(n245), .Y(n329) );
  NAND2X1 U305 ( .A(R2[25]), .B(n195), .Y(n327) );
  NAND3X1 U306 ( .A(n278), .B(n277), .C(n276), .Y(data_out[42]) );
  NAND2X1 U307 ( .A(R2[8]), .B(n192), .Y(n276) );
  NAND2X1 U308 ( .A(data_in_1[42]), .B(n184), .Y(n277) );
  NAND2X1 U309 ( .A(data_in_2[42]), .B(n207), .Y(n278) );
  NAND3X1 U310 ( .A(n430), .B(n429), .C(n428), .Y(data_out[93]) );
  NAND2X1 U311 ( .A(data_in_1[93]), .B(n185), .Y(n429) );
  NAND2X1 U312 ( .A(data_in_2[93]), .B(n180), .Y(n430) );
  NAND2X1 U313 ( .A(R3[25]), .B(n190), .Y(n428) );
  NAND3X1 U314 ( .A(n379), .B(n378), .C(n377), .Y(data_out[76]) );
  NAND2X1 U315 ( .A(data_in_1[76]), .B(n187), .Y(n378) );
  NAND2X1 U316 ( .A(data_in_2[76]), .B(n243), .Y(n379) );
  NAND2X1 U317 ( .A(R3[8]), .B(n193), .Y(n377) );
  NAND3X1 U318 ( .A(n530), .B(n529), .C(n528), .Y(data_out[127]) );
  NAND2X1 U319 ( .A(data_in_1[127]), .B(n187), .Y(n529) );
  NAND2XL U320 ( .A(R4[25]), .B(n193), .Y(n528) );
  NAND2X1 U321 ( .A(data_in_2[127]), .B(n180), .Y(n530) );
  NAND3X1 U322 ( .A(n477), .B(n476), .C(n475), .Y(data_out[110]) );
  NAND2X1 U323 ( .A(data_in_1[110]), .B(n184), .Y(n476) );
  NAND2X1 U324 ( .A(data_in_2[110]), .B(n180), .Y(n477) );
  NAND2X1 U325 ( .A(R4[8]), .B(n191), .Y(n475) );
  NAND3X1 U326 ( .A(n332), .B(n331), .C(n330), .Y(data_out[60]) );
  NAND2X1 U327 ( .A(data_in_1[60]), .B(n187), .Y(n331) );
  NAND2X1 U328 ( .A(data_in_2[60]), .B(n235), .Y(n332) );
  NAND2X1 U329 ( .A(R2[26]), .B(n194), .Y(n330) );
  NAND3X1 U330 ( .A(n283), .B(n280), .C(n279), .Y(data_out[43]) );
  NAND2X1 U331 ( .A(R2[9]), .B(n195), .Y(n279) );
  NAND2X1 U332 ( .A(data_in_1[43]), .B(n183), .Y(n280) );
  NAND2X1 U333 ( .A(data_in_2[43]), .B(n180), .Y(n283) );
  NAND3X1 U334 ( .A(n433), .B(n432), .C(n431), .Y(data_out[94]) );
  NAND2X1 U335 ( .A(data_in_1[94]), .B(n185), .Y(n432) );
  NAND2X1 U336 ( .A(data_in_2[94]), .B(n180), .Y(n433) );
  NAND2X1 U337 ( .A(R3[26]), .B(n192), .Y(n431) );
  NAND3X1 U338 ( .A(n382), .B(n381), .C(n380), .Y(data_out[77]) );
  NAND2X1 U339 ( .A(data_in_1[77]), .B(n186), .Y(n381) );
  NAND2X1 U340 ( .A(data_in_2[77]), .B(n219), .Y(n382) );
  NAND2X1 U341 ( .A(R3[9]), .B(n195), .Y(n380) );
  NAND3X1 U342 ( .A(n533), .B(n532), .C(n531), .Y(data_out[128]) );
  NAND2X1 U343 ( .A(data_in_1[128]), .B(n187), .Y(n532) );
  NAND2XL U344 ( .A(R4[26]), .B(n195), .Y(n531) );
  NAND2X1 U345 ( .A(data_in_2[128]), .B(n180), .Y(n533) );
  NAND3X1 U346 ( .A(n480), .B(n479), .C(n478), .Y(data_out[111]) );
  NAND2X1 U347 ( .A(data_in_1[111]), .B(n183), .Y(n479) );
  NAND2X1 U348 ( .A(data_in_2[111]), .B(n180), .Y(n480) );
  NAND2X1 U349 ( .A(R4[9]), .B(n194), .Y(n478) );
  NAND3X1 U350 ( .A(n335), .B(n334), .C(n333), .Y(data_out[61]) );
  NAND2X1 U351 ( .A(data_in_1[61]), .B(n184), .Y(n334) );
  NAND2X1 U352 ( .A(data_in_2[61]), .B(n219), .Y(n335) );
  NAND2X1 U353 ( .A(R2[27]), .B(n550), .Y(n333) );
  NAND3X1 U354 ( .A(n287), .B(n286), .C(n284), .Y(data_out[44]) );
  NAND2X1 U355 ( .A(R2[10]), .B(n192), .Y(n284) );
  NAND2X1 U356 ( .A(data_in_1[44]), .B(n549), .Y(n286) );
  NAND2X1 U357 ( .A(data_in_2[44]), .B(n248), .Y(n287) );
  NAND3X1 U358 ( .A(n436), .B(n435), .C(n434), .Y(data_out[95]) );
  NAND2X1 U359 ( .A(data_in_1[95]), .B(n187), .Y(n435) );
  NAND2X1 U360 ( .A(data_in_2[95]), .B(n180), .Y(n436) );
  NAND2X1 U361 ( .A(R3[27]), .B(n550), .Y(n434) );
  NAND3X1 U362 ( .A(n385), .B(n384), .C(n383), .Y(data_out[78]) );
  NAND2X1 U363 ( .A(data_in_1[78]), .B(n185), .Y(n384) );
  NAND2X1 U364 ( .A(data_in_2[78]), .B(n248), .Y(n385) );
  NAND2X1 U365 ( .A(R3[10]), .B(n190), .Y(n383) );
  NAND3X1 U366 ( .A(n536), .B(n535), .C(n534), .Y(data_out[129]) );
  NAND2X1 U367 ( .A(data_in_1[129]), .B(n186), .Y(n535) );
  NAND2XL U368 ( .A(R4[27]), .B(n191), .Y(n534) );
  NAND2X1 U369 ( .A(data_in_2[129]), .B(n180), .Y(n536) );
  NAND3X1 U370 ( .A(n483), .B(n482), .C(n481), .Y(data_out[112]) );
  NAND2X1 U371 ( .A(data_in_1[112]), .B(n549), .Y(n482) );
  NAND2X1 U372 ( .A(data_in_2[112]), .B(n180), .Y(n483) );
  NAND2X1 U373 ( .A(R4[10]), .B(n195), .Y(n481) );
  NAND3X1 U374 ( .A(n338), .B(n337), .C(n336), .Y(data_out[62]) );
  NAND2X1 U375 ( .A(data_in_1[62]), .B(n186), .Y(n337) );
  NAND2X1 U376 ( .A(data_in_2[62]), .B(n240), .Y(n338) );
  NAND2X1 U377 ( .A(R2[28]), .B(n190), .Y(n336) );
  NAND3X1 U378 ( .A(n290), .B(n289), .C(n288), .Y(data_out[45]) );
  NAND2X1 U379 ( .A(R2[11]), .B(n190), .Y(n288) );
  NAND2X1 U380 ( .A(data_in_1[45]), .B(n186), .Y(n289) );
  NAND2X1 U381 ( .A(data_in_2[45]), .B(n180), .Y(n290) );
  NAND3X1 U382 ( .A(n439), .B(n438), .C(n437), .Y(data_out[96]) );
  NAND2X1 U383 ( .A(data_in_1[96]), .B(n186), .Y(n438) );
  NAND2X1 U384 ( .A(data_in_2[96]), .B(n180), .Y(n439) );
  NAND2X1 U385 ( .A(R3[28]), .B(n193), .Y(n437) );
  NAND3X1 U386 ( .A(n388), .B(n387), .C(n386), .Y(data_out[79]) );
  NAND2X1 U387 ( .A(data_in_1[79]), .B(n549), .Y(n387) );
  NAND2X1 U388 ( .A(data_in_2[79]), .B(n237), .Y(n388) );
  NAND2X1 U389 ( .A(R3[11]), .B(n193), .Y(n386) );
  NAND3X1 U390 ( .A(n539), .B(n538), .C(n537), .Y(data_out[130]) );
  NAND2X1 U391 ( .A(data_in_1[130]), .B(n185), .Y(n538) );
  NAND2XL U392 ( .A(R4[28]), .B(n194), .Y(n537) );
  NAND2X1 U393 ( .A(data_in_2[130]), .B(n180), .Y(n539) );
  NAND3X1 U394 ( .A(n486), .B(n485), .C(n484), .Y(data_out[113]) );
  NAND2X1 U395 ( .A(data_in_1[113]), .B(n187), .Y(n485) );
  NAND2X1 U396 ( .A(data_in_2[113]), .B(n180), .Y(n486) );
  NAND2X1 U397 ( .A(R4[11]), .B(n193), .Y(n484) );
  NAND3X1 U398 ( .A(n341), .B(n340), .C(n339), .Y(data_out[63]) );
  NAND2X1 U399 ( .A(data_in_1[63]), .B(n185), .Y(n340) );
  NAND2X1 U400 ( .A(data_in_2[63]), .B(n180), .Y(n341) );
  NAND2X1 U401 ( .A(R2[29]), .B(n193), .Y(n339) );
  NAND3X1 U402 ( .A(n293), .B(n292), .C(n291), .Y(data_out[46]) );
  NAND2X1 U403 ( .A(data_in_1[46]), .B(n187), .Y(n292) );
  NAND2X1 U404 ( .A(data_in_2[46]), .B(n180), .Y(n293) );
  NAND2X1 U405 ( .A(R2[12]), .B(n194), .Y(n291) );
  NAND3X1 U406 ( .A(n442), .B(n441), .C(n440), .Y(data_out[97]) );
  NAND2X1 U407 ( .A(data_in_1[97]), .B(n185), .Y(n441) );
  NAND2X1 U408 ( .A(data_in_2[97]), .B(n180), .Y(n442) );
  NAND2X1 U409 ( .A(R3[29]), .B(n195), .Y(n440) );
  NAND3X1 U410 ( .A(n391), .B(n390), .C(n389), .Y(data_out[80]) );
  NAND2X1 U411 ( .A(data_in_1[80]), .B(n187), .Y(n390) );
  NAND2X1 U412 ( .A(data_in_2[80]), .B(n245), .Y(n391) );
  NAND2X1 U413 ( .A(R3[12]), .B(n191), .Y(n389) );
  NAND3X1 U414 ( .A(n542), .B(n541), .C(n540), .Y(data_out[131]) );
  NAND2X1 U415 ( .A(data_in_1[131]), .B(n549), .Y(n541) );
  NAND2XL U416 ( .A(R4[29]), .B(n192), .Y(n540) );
  NAND2X1 U417 ( .A(data_in_2[131]), .B(n180), .Y(n542) );
  NAND3X1 U418 ( .A(n489), .B(n488), .C(n487), .Y(data_out[114]) );
  NAND2X1 U419 ( .A(data_in_1[114]), .B(n186), .Y(n488) );
  NAND2X1 U420 ( .A(data_in_2[114]), .B(n180), .Y(n489) );
  NAND2X1 U421 ( .A(R4[12]), .B(n195), .Y(n487) );
  NAND3X1 U422 ( .A(n344), .B(n343), .C(n342), .Y(data_out[64]) );
  NAND2X1 U423 ( .A(data_in_1[64]), .B(n186), .Y(n343) );
  NAND2X1 U424 ( .A(data_in_2[64]), .B(n243), .Y(n344) );
  NAND2X1 U425 ( .A(R2[30]), .B(n191), .Y(n342) );
  NAND3X1 U426 ( .A(n296), .B(n295), .C(n294), .Y(data_out[47]) );
  NAND2X1 U427 ( .A(data_in_1[47]), .B(n187), .Y(n295) );
  NAND2X1 U428 ( .A(data_in_2[47]), .B(n219), .Y(n296) );
  NAND2X1 U429 ( .A(R2[13]), .B(n192), .Y(n294) );
  NAND3X1 U430 ( .A(n445), .B(n444), .C(n443), .Y(data_out[98]) );
  NAND2X1 U431 ( .A(data_in_1[98]), .B(n186), .Y(n444) );
  NAND2X1 U432 ( .A(data_in_2[98]), .B(n180), .Y(n445) );
  NAND2X1 U433 ( .A(R3[30]), .B(n194), .Y(n443) );
  NAND3X1 U434 ( .A(n394), .B(n393), .C(n392), .Y(data_out[81]) );
  NAND2X1 U435 ( .A(data_in_1[81]), .B(n187), .Y(n393) );
  NAND2X1 U436 ( .A(data_in_2[81]), .B(n224), .Y(n394) );
  NAND2X1 U437 ( .A(R3[13]), .B(n192), .Y(n392) );
  NAND3X1 U438 ( .A(n545), .B(n544), .C(n543), .Y(data_out[132]) );
  NAND2X1 U439 ( .A(data_in_1[132]), .B(n187), .Y(n544) );
  NAND2XL U440 ( .A(R4[30]), .B(n550), .Y(n543) );
  NAND2X1 U441 ( .A(data_in_2[132]), .B(n180), .Y(n545) );
  NAND3X1 U442 ( .A(n492), .B(n491), .C(n490), .Y(data_out[115]) );
  NAND2X1 U443 ( .A(data_in_1[115]), .B(n185), .Y(n491) );
  NAND2X1 U444 ( .A(data_in_2[115]), .B(n180), .Y(n492) );
  NAND2X1 U445 ( .A(R4[13]), .B(n190), .Y(n490) );
  NAND3X1 U446 ( .A(n347), .B(n346), .C(n345), .Y(data_out[65]) );
  NAND2X1 U447 ( .A(data_in_1[65]), .B(n187), .Y(n346) );
  NAND2X1 U448 ( .A(data_in_2[65]), .B(n180), .Y(n347) );
  NAND2X1 U449 ( .A(R2[31]), .B(n192), .Y(n345) );
  NAND3X1 U450 ( .A(n299), .B(n298), .C(n297), .Y(data_out[48]) );
  NAND2X1 U451 ( .A(data_in_1[48]), .B(n186), .Y(n298) );
  NAND2X1 U452 ( .A(data_in_2[48]), .B(n248), .Y(n299) );
  NAND2X1 U453 ( .A(R2[14]), .B(n550), .Y(n297) );
  NAND3X1 U454 ( .A(n448), .B(n447), .C(n446), .Y(data_out[99]) );
  NAND2X1 U455 ( .A(data_in_1[99]), .B(n187), .Y(n447) );
  NAND2X1 U456 ( .A(data_in_2[99]), .B(n180), .Y(n448) );
  NAND2X1 U457 ( .A(R3[31]), .B(n195), .Y(n446) );
  NAND3X1 U458 ( .A(n397), .B(n396), .C(n395), .Y(data_out[82]) );
  NAND2X1 U459 ( .A(data_in_1[82]), .B(n184), .Y(n396) );
  NAND2X1 U460 ( .A(data_in_2[82]), .B(n216), .Y(n397) );
  NAND2X1 U461 ( .A(R3[14]), .B(n193), .Y(n395) );
  NAND3X1 U462 ( .A(n548), .B(n547), .C(n546), .Y(data_out[133]) );
  NAND2X1 U463 ( .A(data_in_1[133]), .B(n185), .Y(n547) );
  NAND2XL U464 ( .A(R4[31]), .B(n192), .Y(n546) );
  NAND2X1 U465 ( .A(data_in_2[133]), .B(n180), .Y(n548) );
  NAND3X1 U466 ( .A(n495), .B(n494), .C(n493), .Y(data_out[116]) );
  NAND2X1 U467 ( .A(data_in_1[116]), .B(n186), .Y(n494) );
  NAND2X1 U468 ( .A(data_in_2[116]), .B(n180), .Y(n495) );
  NAND2X1 U469 ( .A(R4[14]), .B(n190), .Y(n493) );
  NAND3X1 U470 ( .A(n350), .B(n349), .C(n348), .Y(data_out[66]) );
  NAND2X1 U471 ( .A(data_in_1[66]), .B(n187), .Y(n349) );
  NAND2X1 U472 ( .A(data_in_2[66]), .B(n180), .Y(n350) );
  NAND2X1 U473 ( .A(R2[32]), .B(n195), .Y(n348) );
  NAND3X1 U474 ( .A(n302), .B(n301), .C(n300), .Y(data_out[49]) );
  NAND2X1 U475 ( .A(data_in_1[49]), .B(n185), .Y(n301) );
  NAND2X1 U476 ( .A(data_in_2[49]), .B(n243), .Y(n302) );
  NAND2X1 U477 ( .A(R2[15]), .B(n194), .Y(n300) );
  NAND3X1 U478 ( .A(n451), .B(n450), .C(n449), .Y(data_out[100]) );
  NAND2X1 U479 ( .A(data_in_1[100]), .B(n187), .Y(n450) );
  NAND2X1 U480 ( .A(data_in_2[100]), .B(n180), .Y(n451) );
  NAND2X1 U481 ( .A(R3[32]), .B(n550), .Y(n449) );
  NAND3X1 U482 ( .A(n400), .B(n399), .C(n398), .Y(data_out[83]) );
  NAND2X1 U483 ( .A(data_in_1[83]), .B(n183), .Y(n399) );
  NAND2X1 U484 ( .A(data_in_2[83]), .B(n221), .Y(n400) );
  NAND2X1 U485 ( .A(R3[15]), .B(n190), .Y(n398) );
  NAND3X1 U486 ( .A(n553), .B(n552), .C(n551), .Y(data_out[134]) );
  NAND2X1 U487 ( .A(data_in_1[134]), .B(n549), .Y(n552) );
  NAND2X1 U488 ( .A(data_in_2[134]), .B(n248), .Y(n553) );
  NAND2X1 U489 ( .A(R4[32]), .B(n550), .Y(n551) );
  NAND3X1 U490 ( .A(n498), .B(n497), .C(n496), .Y(data_out[117]) );
  NAND2X1 U491 ( .A(data_in_1[117]), .B(n185), .Y(n497) );
  NAND2X1 U492 ( .A(data_in_2[117]), .B(n180), .Y(n498) );
  NAND2X1 U493 ( .A(R4[15]), .B(n192), .Y(n496) );
  NAND3X1 U494 ( .A(n320), .B(n319), .C(n318), .Y(data_out[56]) );
  NAND2X1 U495 ( .A(data_in_1[56]), .B(n187), .Y(n319) );
  NAND2X1 U496 ( .A(data_in_2[56]), .B(n207), .Y(n320) );
  NAND2X1 U497 ( .A(R2[22]), .B(n190), .Y(n318) );
  NAND3X1 U498 ( .A(n317), .B(n316), .C(n315), .Y(data_out[55]) );
  NAND2X1 U499 ( .A(data_in_1[55]), .B(n187), .Y(n316) );
  NAND2X1 U500 ( .A(data_in_2[55]), .B(n237), .Y(n317) );
  NAND2X1 U501 ( .A(R2[21]), .B(n195), .Y(n315) );
  NAND3X1 U502 ( .A(n257), .B(n256), .C(n255), .Y(data_out[35]) );
  NAND2X1 U503 ( .A(R2[1]), .B(n191), .Y(n255) );
  NAND2X1 U504 ( .A(data_in_1[35]), .B(n184), .Y(n256) );
  NAND2X1 U505 ( .A(data_in_2[35]), .B(n180), .Y(n257) );
  NAND3X1 U506 ( .A(n260), .B(n259), .C(n258), .Y(data_out[36]) );
  NAND2X1 U507 ( .A(data_in_1[36]), .B(n186), .Y(n259) );
  NAND2X1 U508 ( .A(R2[2]), .B(n195), .Y(n258) );
  NAND2X1 U509 ( .A(data_in_2[36]), .B(n237), .Y(n260) );
  NAND3X1 U510 ( .A(n266), .B(n265), .C(n264), .Y(data_out[38]) );
  NAND2X1 U511 ( .A(data_in_1[38]), .B(n186), .Y(n265) );
  NAND2X1 U512 ( .A(R2[4]), .B(n194), .Y(n264) );
  NAND2X1 U513 ( .A(data_in_2[38]), .B(n180), .Y(n266) );
  NAND3X1 U514 ( .A(n409), .B(n408), .C(n407), .Y(data_out[86]) );
  NAND2X1 U515 ( .A(data_in_1[86]), .B(n184), .Y(n408) );
  NAND2X1 U516 ( .A(data_in_2[86]), .B(n243), .Y(n409) );
  NAND2X1 U517 ( .A(R3[18]), .B(n191), .Y(n407) );
  NAND3X1 U518 ( .A(n412), .B(n411), .C(n410), .Y(data_out[87]) );
  NAND2X1 U519 ( .A(data_in_1[87]), .B(n184), .Y(n411) );
  NAND2X1 U520 ( .A(data_in_2[87]), .B(n235), .Y(n412) );
  NAND2X1 U521 ( .A(R3[19]), .B(n195), .Y(n410) );
  NAND3X1 U522 ( .A(n358), .B(n357), .C(n356), .Y(data_out[69]) );
  NAND2X1 U523 ( .A(data_in_1[69]), .B(n184), .Y(n357) );
  NAND2X1 U524 ( .A(data_in_2[69]), .B(n180), .Y(n358) );
  NAND2X1 U525 ( .A(R3[1]), .B(n194), .Y(n356) );
  NAND3X1 U526 ( .A(n361), .B(n360), .C(n359), .Y(data_out[70]) );
  NAND2X1 U527 ( .A(data_in_1[70]), .B(n183), .Y(n360) );
  NAND2X1 U528 ( .A(data_in_2[70]), .B(n248), .Y(n361) );
  NAND2X1 U529 ( .A(R3[2]), .B(n195), .Y(n359) );
  OAI2BB1X1 U530 ( .A0N(data_in_2[34]), .A1N(n216), .B0(n254), .Y(data_out[34]) );
  AOI22XL U531 ( .A0(data_in_1[34]), .A1(n186), .B0(R2[0]), .B1(n195), .Y(n254) );
  OAI2BB1X1 U532 ( .A0N(data_in_2[85]), .A1N(n209), .B0(n406), .Y(data_out[85]) );
  AOI22XL U533 ( .A0(data_in_1[85]), .A1(n185), .B0(R3[17]), .B1(n192), .Y(
        n406) );
  OAI2BB1X1 U534 ( .A0N(data_in_2[68]), .A1N(n181), .B0(n355), .Y(data_out[68]) );
  AOI22XL U535 ( .A0(data_in_1[68]), .A1(n549), .B0(R3[0]), .B1(n550), .Y(n355) );
  NAND2X4 U536 ( .A(n175), .B(n499), .Y(n403) );
  INVX8 U537 ( .A(n555), .Y(n556) );
  NAND2XL U538 ( .A(n26), .B(n24), .Y(n282) );
  OAI2BB1X4 U539 ( .A0N(data_in_2[0]), .A1N(n181), .B0(n202), .Y(data_out[0])
         );
  OAI2BB1X4 U540 ( .A0N(data_in_2[2]), .A1N(n205), .B0(n204), .Y(data_out[2])
         );
  OAI2BB1X4 U541 ( .A0N(data_in_2[3]), .A1N(n207), .B0(n206), .Y(data_out[3])
         );
  OAI2BB1X4 U542 ( .A0N(data_in_2[4]), .A1N(n209), .B0(n208), .Y(data_out[4])
         );
  NAND2X4 U543 ( .A(R1[5]), .B(n550), .Y(n213) );
  NAND2BX4 U544 ( .AN(n214), .B(n213), .Y(data_out[5]) );
  OAI2BB1X4 U545 ( .A0N(data_in_2[6]), .A1N(n216), .B0(n215), .Y(data_out[6])
         );
  OAI2BB1X4 U546 ( .A0N(data_in_2[8]), .A1N(n219), .B0(n218), .Y(data_out[8])
         );
  OAI2BB1X4 U547 ( .A0N(data_in_2[17]), .A1N(n181), .B0(n230), .Y(data_out[17]) );
  OAI2BB1X4 U548 ( .A0N(data_in_2[18]), .A1N(n205), .B0(n231), .Y(data_out[18]) );
  AOI22X4 U549 ( .A0(data_in_1[19]), .A1(n187), .B0(R1[19]), .B1(n191), .Y(
        n232) );
  OAI2BB1X4 U550 ( .A0N(data_in_2[19]), .A1N(n181), .B0(n232), .Y(data_out[19]) );
  OAI2BB1X4 U551 ( .A0N(data_in_2[21]), .A1N(n235), .B0(n234), .Y(data_out[21]) );
  OAI2BB1X4 U552 ( .A0N(data_in_2[22]), .A1N(n237), .B0(n236), .Y(data_out[22]) );
  OAI2BB1X4 U553 ( .A0N(data_in_2[24]), .A1N(n240), .B0(n239), .Y(data_out[24]) );
  OAI2BB1X4 U554 ( .A0N(data_in_2[26]), .A1N(n243), .B0(n242), .Y(data_out[26]) );
  OAI2BB1X4 U555 ( .A0N(data_in_2[28]), .A1N(n248), .B0(n247), .Y(data_out[28]) );
  NOR3BX4 U556 ( .AN(counter[1]), .B(n18), .C(n174), .Y(n354) );
  NAND2BX4 U557 ( .AN(n36), .B(n354), .Y(n351) );
  NAND2BX4 U558 ( .AN(n36), .B(n35), .Y(n555) );
  OAI2BB1X4 U559 ( .A0N(n504), .A1N(n405), .B0(n404), .Y(data_out[84]) );
  NOR2X4 U560 ( .A(n18), .B(n174), .Y(n499) );
  OAI2BB1X4 U561 ( .A0N(n504), .A1N(n505), .B0(n503), .Y(data_out[118]) );
endmodule


module multi16_0_DW01_add_5 ( A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, 
        A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, 
        A_4_, B_23_, B_22_, B_21_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, 
        B_14_, B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, 
        SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, 
        SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, 
        SUM_7_ );
  input A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_,
         A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, B_23_, B_22_,
         B_21_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_,
         B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_;
  output SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_,
         SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_,
         SUM_8_, SUM_7_;
  wire   n1, n2, n3, n4;
  wire   [23:7] carry;

  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry[7]), .CO(carry[8]), .S(SUM_7_)
         );
  ADDFX2 U1_21 ( .A(A_21_), .B(B_21_), .CI(carry[21]), .CO(carry[22]), .S(
        SUM_21_) );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry[20]), .CO(carry[21]), .S(
        SUM_20_) );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry[19]), .CO(carry[20]), .S(
        SUM_19_) );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry[18]), .CO(carry[19]), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry[17]), .CO(carry[18]), .S(
        SUM_17_) );
  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry[16]), .CO(carry[17]), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry[15]), .CO(carry[16]), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry[14]), .CO(carry[15]), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry[13]), .CO(carry[14]), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry[12]), .CO(carry[13]), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry[11]), .CO(carry[12]), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry[10]), .CO(carry[11]), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry[9]), .CO(carry[10]), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry[8]), .CO(carry[9]), .S(SUM_8_)
         );
  ADDFX2 U1_22 ( .A(A_22_), .B(B_22_), .CI(carry[22]), .CO(carry[23]), .S(
        SUM_22_) );
  AND2X2 U1 ( .A(A_4_), .B(B_4_), .Y(n1) );
  XOR2X1 U2 ( .A(B_23_), .B(carry[23]), .Y(SUM_23_) );
  OAI2BB1X1 U3 ( .A0N(n2), .A1N(A_6_), .B0(n3), .Y(carry[7]) );
  OAI21XL U4 ( .A0(A_6_), .A1(n2), .B0(B_6_), .Y(n3) );
  OAI2BB1X1 U5 ( .A0N(n1), .A1N(A_5_), .B0(n4), .Y(n2) );
  OAI21XL U6 ( .A0(A_5_), .A1(n1), .B0(B_5_), .Y(n4) );
endmodule


module multi16_0_DW01_add_3 ( A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, 
        A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, 
        B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, 
        B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, SUM_22_, SUM_21_, SUM_20_, 
        SUM_19_, SUM_18_, SUM_17_, SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, 
        SUM_11_, SUM_10_, SUM_9_, SUM_8_, SUM_7_ );
  input A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_,
         A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, B_20_, B_19_,
         B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, B_10_, B_9_,
         B_8_, B_7_, B_6_, B_5_;
  output SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_,
         SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_,
         SUM_7_;
  wire   carry_21_, carry_20_, carry_19_, carry_18_, carry_17_, carry_16_,
         carry_15_, carry_14_, carry_13_, carry_12_, carry_11_, carry_10_,
         carry_9_, carry_8_, carry_7_, n1;

  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry_16_), .CO(carry_17_), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry_15_), .CO(carry_16_), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry_14_), .CO(carry_15_), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry_13_), .CO(carry_14_), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry_12_), .CO(carry_13_), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry_11_), .CO(carry_12_), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry_10_), .CO(carry_11_), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry_9_), .CO(carry_10_), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry_8_), .CO(carry_9_), .S(SUM_8_)
         );
  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry_7_), .CO(carry_8_), .S(SUM_7_)
         );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry_20_), .CO(carry_21_), .S(
        SUM_20_) );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry_19_), .CO(carry_20_), .S(
        SUM_19_) );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry_18_), .CO(carry_19_), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry_17_), .CO(carry_18_), .S(
        SUM_17_) );
  ADDFX2 U1_21 ( .A(A_21_), .B(B_21_), .CI(carry_21_), .CO(SUM_22_), .S(
        SUM_21_) );
  OAI2BB1X1 U1 ( .A0N(A_6_), .A1N(B_6_), .B0(n1), .Y(carry_7_) );
  OAI211X1 U2 ( .A0(B_6_), .A1(A_6_), .B0(A_5_), .C0(B_5_), .Y(n1) );
endmodule


module multi16_0_DW01_add_0 ( A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, 
        A_16_, A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, 
        A_6_, A_5_, A_4_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, 
        B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, 
        SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, 
        SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, 
        SUM_7_ );
  input A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_,
         A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, B_20_,
         B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, B_10_,
         B_9_, B_8_, B_7_, B_6_, B_5_, B_4_;
  output SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_,
         SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_,
         SUM_8_, SUM_7_;
  wire   n1, n2, n3, n4, n5, n6;
  wire   [21:7] carry;

  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry[7]), .CO(carry[8]), .S(SUM_7_)
         );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry[18]), .CO(carry[19]), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry[17]), .CO(carry[18]), .S(
        SUM_17_) );
  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry[16]), .CO(carry[17]), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry[15]), .CO(carry[16]), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry[14]), .CO(carry[15]), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry[13]), .CO(carry[14]), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry[12]), .CO(carry[13]), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry[11]), .CO(carry[12]), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry[10]), .CO(carry[11]), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry[9]), .CO(carry[10]), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry[8]), .CO(carry[9]), .S(SUM_8_)
         );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry[19]), .CO(carry[20]), .S(
        SUM_19_) );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry[20]), .CO(carry[21]), .S(
        SUM_20_) );
  AND2X2 U1 ( .A(A_22_), .B(n2), .Y(n1) );
  AND2X2 U2 ( .A(A_21_), .B(carry[21]), .Y(n2) );
  AND2X2 U3 ( .A(A_4_), .B(B_4_), .Y(n3) );
  XOR2X1 U4 ( .A(A_23_), .B(n1), .Y(SUM_23_) );
  XOR2X1 U5 ( .A(A_21_), .B(carry[21]), .Y(SUM_21_) );
  XOR2X1 U6 ( .A(A_22_), .B(n2), .Y(SUM_22_) );
  OAI2BB1X1 U7 ( .A0N(n4), .A1N(A_6_), .B0(n5), .Y(carry[7]) );
  OAI21XL U8 ( .A0(A_6_), .A1(n4), .B0(B_6_), .Y(n5) );
  OAI2BB1X1 U9 ( .A0N(n3), .A1N(A_5_), .B0(n6), .Y(n4) );
  OAI21XL U10 ( .A0(A_5_), .A1(n3), .B0(B_5_), .Y(n6) );
endmodule


module multi16_0 ( in_17bit, in_8bit, out );
  input [16:0] in_17bit;
  input [7:0] in_8bit;
  output [16:0] out;
  wire   n225, n226, n227, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23,
         N24, N25, N26, N27, N28, N29, N108, N109, N110, N111, N112, N113,
         N114, N115, N116, N117, N118, N119, N120, N121, N122, N123, N205,
         N206, N207, N208, N209, N210, N211, N212, N213, N214, N215, N216,
         N217, N218, N219, N220, N221, N347, N348, N349, N350, N351, N352,
         N353, N354, N355, N356, N357, N358, N359, N360, N361, N362, N363,
         N446, N447, N448, N449, N450, N451, N452, N453, N454, N455, N456,
         N457, N458, N459, N460, N461, N462, N463, N479, N480, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         add_2_root_r115_carry_10_, add_2_root_r115_carry_11_,
         add_2_root_r115_carry_12_, add_2_root_r115_carry_13_,
         add_2_root_r115_carry_14_, add_2_root_r115_carry_15_,
         add_2_root_r115_carry_16_, add_2_root_r115_carry_17_,
         add_2_root_r115_carry_18_, add_2_root_r115_carry_19_,
         add_2_root_r115_carry_5_, add_2_root_r115_carry_6_,
         add_2_root_r115_carry_7_, add_2_root_r115_carry_8_,
         add_2_root_r115_carry_9_, add_2_root_r115_SUM_3_,
         add_2_root_r115_SUM_4_, add_2_root_r115_SUM_5_,
         add_2_root_r115_SUM_6_, add_2_root_r115_SUM_7_,
         add_2_root_r115_SUM_8_, add_2_root_r115_SUM_9_,
         add_2_root_r115_SUM_10_, add_2_root_r115_SUM_11_,
         add_2_root_r115_SUM_12_, add_2_root_r115_SUM_13_,
         add_2_root_r115_SUM_14_, add_2_root_r115_SUM_15_,
         add_2_root_r115_SUM_16_, add_2_root_r115_SUM_17_,
         add_2_root_r115_SUM_18_, add_2_root_r115_SUM_19_,
         add_2_root_r115_SUM_20_, add_1_root_r115_carry_10_,
         add_1_root_r115_carry_11_, add_1_root_r115_carry_12_,
         add_1_root_r115_carry_13_, add_1_root_r115_carry_14_,
         add_1_root_r115_carry_15_, add_1_root_r115_carry_16_,
         add_1_root_r115_carry_17_, add_1_root_r115_carry_18_,
         add_1_root_r115_carry_19_, add_1_root_r115_carry_20_,
         add_1_root_r115_carry_21_, add_1_root_r115_carry_22_,
         add_1_root_r115_carry_7_, add_1_root_r115_carry_8_,
         add_1_root_r115_carry_9_, add_1_root_r115_SUM_7_,
         add_1_root_r115_SUM_8_, add_1_root_r115_SUM_9_,
         add_1_root_r115_SUM_10_, add_1_root_r115_SUM_11_,
         add_1_root_r115_SUM_12_, add_1_root_r115_SUM_13_,
         add_1_root_r115_SUM_14_, add_1_root_r115_SUM_15_,
         add_1_root_r115_SUM_16_, add_1_root_r115_SUM_17_,
         add_1_root_r115_SUM_18_, add_1_root_r115_SUM_19_,
         add_1_root_r115_SUM_20_, add_1_root_r115_SUM_21_,
         add_1_root_r115_SUM_22_, add_1_root_r115_SUM_23_,
         add_1_root_r112_carry_10_, add_1_root_r112_carry_11_,
         add_1_root_r112_carry_12_, add_1_root_r112_carry_13_,
         add_1_root_r112_carry_14_, add_1_root_r112_carry_15_,
         add_1_root_r112_carry_16_, add_1_root_r112_carry_17_,
         add_1_root_r112_carry_18_, add_1_root_r112_carry_19_,
         add_1_root_r112_carry_20_, add_1_root_r112_carry_5_,
         add_1_root_r112_carry_6_, add_1_root_r112_carry_7_,
         add_1_root_r112_carry_8_, add_1_root_r112_carry_9_,
         add_1_root_r112_SUM_1_, add_1_root_r112_SUM_2_,
         add_1_root_r112_SUM_3_, add_1_root_r112_SUM_4_,
         add_1_root_r112_SUM_5_, add_1_root_r112_SUM_6_,
         add_1_root_r112_SUM_7_, add_1_root_r112_SUM_8_,
         add_1_root_r112_SUM_9_, add_1_root_r112_SUM_10_,
         add_1_root_r112_SUM_11_, add_1_root_r112_SUM_12_,
         add_1_root_r112_SUM_13_, add_1_root_r112_SUM_14_,
         add_1_root_r112_SUM_15_, add_1_root_r112_SUM_16_,
         add_1_root_r112_SUM_17_, add_1_root_r112_SUM_18_,
         add_1_root_r112_SUM_19_, add_1_root_r112_SUM_20_,
         add_1_root_r112_SUM_21_, add_2_root_r119_carry_10_,
         add_2_root_r119_carry_11_, add_2_root_r119_carry_12_,
         add_2_root_r119_carry_13_, add_2_root_r119_carry_14_,
         add_2_root_r119_carry_15_, add_2_root_r119_carry_16_,
         add_2_root_r119_carry_17_, add_2_root_r119_carry_18_,
         add_2_root_r119_carry_19_, add_2_root_r119_carry_20_,
         add_2_root_r119_carry_21_, add_2_root_r119_carry_7_,
         add_2_root_r119_carry_8_, add_2_root_r119_carry_9_,
         add_2_root_r119_SUM_5_, add_2_root_r119_SUM_6_,
         add_2_root_r119_SUM_7_, add_2_root_r119_SUM_8_,
         add_2_root_r119_SUM_9_, add_2_root_r119_SUM_10_,
         add_2_root_r119_SUM_11_, add_2_root_r119_SUM_12_,
         add_2_root_r119_SUM_13_, add_2_root_r119_SUM_14_,
         add_2_root_r119_SUM_15_, add_2_root_r119_SUM_16_,
         add_2_root_r119_SUM_17_, add_2_root_r119_SUM_18_,
         add_2_root_r119_SUM_19_, add_2_root_r119_SUM_20_,
         add_2_root_r119_SUM_21_, add_2_root_r119_SUM_22_,
         add_1_root_r119_SUM_6_, add_1_root_r119_SUM_7_,
         add_1_root_r119_SUM_8_, add_1_root_r119_SUM_9_,
         add_1_root_r119_SUM_10_, add_1_root_r119_SUM_11_,
         add_1_root_r119_SUM_12_, add_1_root_r119_SUM_13_,
         add_1_root_r119_SUM_14_, add_1_root_r119_SUM_15_,
         add_1_root_r119_SUM_16_, add_1_root_r119_SUM_17_,
         add_1_root_r119_SUM_18_, add_1_root_r119_SUM_19_,
         add_1_root_r119_SUM_20_, add_1_root_r119_SUM_21_,
         add_1_root_r119_SUM_22_, add_1_root_r119_SUM_23_,
         add_1_root_r119_A_3_, add_1_root_r119_A_4_, add_1_root_r119_A_5_,
         add_1_root_r119_A_6_, add_1_root_r119_A_7_, add_1_root_r119_A_8_,
         add_1_root_r119_A_9_, add_1_root_r119_A_10_, add_1_root_r119_A_11_,
         add_1_root_r119_A_12_, add_1_root_r119_A_13_, add_1_root_r119_A_14_,
         add_1_root_r119_A_15_, add_1_root_r119_A_16_, add_1_root_r119_A_17_,
         add_1_root_r119_A_18_, add_1_root_r119_A_19_,
         add_3_root_r119_carry_10_, add_3_root_r119_carry_11_,
         add_3_root_r119_carry_12_, add_3_root_r119_carry_13_,
         add_3_root_r119_carry_14_, add_3_root_r119_carry_15_,
         add_3_root_r119_carry_16_, add_3_root_r119_carry_17_,
         add_3_root_r119_carry_18_, add_3_root_r119_carry_3_,
         add_3_root_r119_carry_4_, add_3_root_r119_carry_5_,
         add_3_root_r119_carry_6_, add_3_root_r119_carry_7_,
         add_3_root_r119_carry_8_, add_3_root_r119_carry_9_, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n15, n16, n17, n19, n21, n22,
         n23, n24, n25, n26, n27, n28, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205;
  wire   [16:0] in_17bit_b;
  wire   [23:8] neg_mul;
  wire   [15:13] sub_add_75_b0_carry;
  wire   [16:2] sub_add_54_b0_carry;
  wire   [22:7] add_1_root_r119_carry;

  multi16_0_DW01_add_5 add_0_root_r119 ( .A_22_(add_2_root_r119_SUM_22_), 
        .A_21_(add_2_root_r119_SUM_21_), .A_20_(add_2_root_r119_SUM_20_), 
        .A_19_(add_2_root_r119_SUM_19_), .A_18_(add_2_root_r119_SUM_18_), 
        .A_17_(add_2_root_r119_SUM_17_), .A_16_(add_2_root_r119_SUM_16_), 
        .A_15_(add_2_root_r119_SUM_15_), .A_14_(add_2_root_r119_SUM_14_), 
        .A_13_(add_2_root_r119_SUM_13_), .A_12_(add_2_root_r119_SUM_12_), 
        .A_11_(add_2_root_r119_SUM_11_), .A_10_(add_2_root_r119_SUM_10_), 
        .A_9_(add_2_root_r119_SUM_9_), .A_8_(add_2_root_r119_SUM_8_), .A_7_(
        add_2_root_r119_SUM_7_), .A_6_(add_2_root_r119_SUM_6_), .A_5_(
        add_2_root_r119_SUM_5_), .A_4_(in_17bit_b[0]), .B_23_(
        add_1_root_r119_SUM_23_), .B_22_(add_1_root_r119_SUM_22_), .B_21_(
        add_1_root_r119_SUM_21_), .B_20_(add_1_root_r119_SUM_20_), .B_19_(
        add_1_root_r119_SUM_19_), .B_18_(add_1_root_r119_SUM_18_), .B_17_(
        add_1_root_r119_SUM_17_), .B_16_(add_1_root_r119_SUM_16_), .B_15_(
        add_1_root_r119_SUM_15_), .B_14_(add_1_root_r119_SUM_14_), .B_13_(
        add_1_root_r119_SUM_13_), .B_12_(add_1_root_r119_SUM_12_), .B_11_(
        add_1_root_r119_SUM_11_), .B_10_(add_1_root_r119_SUM_10_), .B_9_(
        add_1_root_r119_SUM_9_), .B_8_(add_1_root_r119_SUM_8_), .B_7_(
        add_1_root_r119_SUM_7_), .B_6_(add_1_root_r119_SUM_6_), .B_5_(
        add_1_root_r119_A_5_), .B_4_(add_1_root_r119_A_4_), .SUM_23_(N363), 
        .SUM_22_(N362), .SUM_21_(N361), .SUM_20_(N360), .SUM_19_(N359), 
        .SUM_18_(N358), .SUM_17_(N357), .SUM_16_(N356), .SUM_15_(N355), 
        .SUM_14_(N354), .SUM_13_(N353), .SUM_12_(N352), .SUM_11_(N351), 
        .SUM_10_(N350), .SUM_9_(N349), .SUM_8_(N348), .SUM_7_(N347) );
  multi16_0_DW01_add_3 add_0_root_r112 ( .A_21_(in_17bit_b[16]), .A_20_(
        in_17bit_b[15]), .A_19_(in_17bit_b[14]), .A_18_(in_17bit_b[13]), 
        .A_17_(in_17bit_b[12]), .A_16_(in_17bit_b[11]), .A_15_(in_17bit_b[10]), 
        .A_14_(in_17bit_b[9]), .A_13_(in_17bit_b[8]), .A_12_(in_17bit_b[7]), 
        .A_11_(in_17bit_b[6]), .A_10_(in_17bit_b[5]), .A_9_(in_17bit_b[4]), 
        .A_8_(in_17bit_b[3]), .A_7_(in_17bit_b[2]), .A_6_(in_17bit_b[1]), 
        .A_5_(in_17bit_b[0]), .B_21_(add_1_root_r112_SUM_21_), .B_20_(
        add_1_root_r112_SUM_20_), .B_19_(add_1_root_r112_SUM_19_), .B_18_(
        add_1_root_r112_SUM_18_), .B_17_(add_1_root_r112_SUM_17_), .B_16_(
        add_1_root_r112_SUM_16_), .B_15_(add_1_root_r112_SUM_15_), .B_14_(
        add_1_root_r112_SUM_14_), .B_13_(add_1_root_r112_SUM_13_), .B_12_(
        add_1_root_r112_SUM_12_), .B_11_(add_1_root_r112_SUM_11_), .B_10_(
        add_1_root_r112_SUM_10_), .B_9_(add_1_root_r112_SUM_9_), .B_8_(
        add_1_root_r112_SUM_8_), .B_7_(add_1_root_r112_SUM_7_), .B_6_(
        add_1_root_r112_SUM_6_), .B_5_(add_1_root_r112_SUM_5_), .SUM_22_(N123), 
        .SUM_21_(N122), .SUM_20_(N121), .SUM_19_(N120), .SUM_18_(N119), 
        .SUM_17_(N118), .SUM_16_(N117), .SUM_15_(N116), .SUM_14_(N115), 
        .SUM_13_(N114), .SUM_12_(N113), .SUM_11_(N112), .SUM_10_(N111), 
        .SUM_9_(N110), .SUM_8_(N109), .SUM_7_(N108) );
  multi16_0_DW01_add_0 add_0_root_r115 ( .A_23_(add_1_root_r115_SUM_23_), 
        .A_22_(add_1_root_r115_SUM_22_), .A_21_(add_1_root_r115_SUM_21_), 
        .A_20_(add_1_root_r115_SUM_20_), .A_19_(add_1_root_r115_SUM_19_), 
        .A_18_(add_1_root_r115_SUM_18_), .A_17_(add_1_root_r115_SUM_17_), 
        .A_16_(add_1_root_r115_SUM_16_), .A_15_(add_1_root_r115_SUM_15_), 
        .A_14_(add_1_root_r115_SUM_14_), .A_13_(add_1_root_r115_SUM_13_), 
        .A_12_(add_1_root_r115_SUM_12_), .A_11_(add_1_root_r115_SUM_11_), 
        .A_10_(add_1_root_r115_SUM_10_), .A_9_(add_1_root_r115_SUM_9_), .A_8_(
        add_1_root_r115_SUM_8_), .A_7_(add_1_root_r115_SUM_7_), .A_6_(
        add_2_root_r115_SUM_3_), .A_5_(in_17bit_b[1]), .A_4_(in_17bit_b[0]), 
        .B_20_(add_2_root_r115_SUM_20_), .B_19_(add_2_root_r115_SUM_19_), 
        .B_18_(add_2_root_r115_SUM_18_), .B_17_(add_2_root_r115_SUM_17_), 
        .B_16_(add_2_root_r115_SUM_16_), .B_15_(add_2_root_r115_SUM_15_), 
        .B_14_(add_2_root_r115_SUM_14_), .B_13_(add_2_root_r115_SUM_13_), 
        .B_12_(add_2_root_r115_SUM_12_), .B_11_(add_2_root_r115_SUM_11_), 
        .B_10_(add_2_root_r115_SUM_10_), .B_9_(add_2_root_r115_SUM_9_), .B_8_(
        add_2_root_r115_SUM_8_), .B_7_(add_2_root_r115_SUM_7_), .B_6_(
        add_2_root_r115_SUM_6_), .B_5_(add_2_root_r115_SUM_5_), .B_4_(
        add_2_root_r115_SUM_4_), .SUM_23_(N221), .SUM_22_(N220), .SUM_21_(N219), .SUM_20_(N218), .SUM_19_(N217), .SUM_18_(N216), .SUM_17_(N215), .SUM_16_(
        N214), .SUM_15_(N213), .SUM_14_(N212), .SUM_13_(N211), .SUM_12_(N210), 
        .SUM_11_(N209), .SUM_10_(N208), .SUM_9_(N207), .SUM_8_(N206), .SUM_7_(
        N205) );
  TLATX1 neg_mul_reg_19_ ( .G(N446), .D(N459), .QN(n5) );
  TLATX1 neg_mul_reg_18_ ( .G(N446), .D(N458), .QN(n4) );
  TLATX1 neg_mul_reg_17_ ( .G(N446), .D(N457), .Q(neg_mul[17]), .QN(n12) );
  TLATX1 neg_mul_reg_16_ ( .G(N446), .D(N456), .QN(n3) );
  TLATX1 neg_mul_reg_11_ ( .G(N446), .D(N451), .QN(n2) );
  TLATX1 neg_mul_reg_23_ ( .G(N446), .D(N463), .Q(neg_mul[23]), .QN(n1) );
  TLATX1 neg_mul_reg_22_ ( .G(N446), .D(N462), .Q(neg_mul[22]), .QN(n6) );
  TLATX1 neg_mul_reg_21_ ( .G(N446), .D(N461), .Q(neg_mul[21]), .QN(n7) );
  TLATX1 neg_mul_reg_20_ ( .G(N446), .D(N460), .QN(n8) );
  TLATX1 neg_mul_reg_8_ ( .G(N446), .D(N448), .Q(neg_mul[8]) );
  TLATX1 neg_mul_reg_9_ ( .G(N446), .D(N449), .Q(neg_mul[9]), .QN(n11) );
  TLATX1 neg_mul_reg_15_ ( .G(N446), .D(N455), .Q(neg_mul[15]) );
  TLATX1 neg_mul_reg_14_ ( .G(N446), .D(N454), .Q(neg_mul[14]), .QN(n10) );
  TLATX1 neg_mul_reg_13_ ( .G(N446), .D(N453), .Q(neg_mul[13]), .QN(n9) );
  TLATX1 neg_mul_reg_12_ ( .G(N446), .D(N452), .Q(neg_mul[12]) );
  TLATX1 neg_mul_reg_10_ ( .G(N446), .D(N450), .Q(neg_mul[10]) );
  TLATX1 neg_mul_reg_7_ ( .G(N446), .D(N447), .Q(out[0]) );
  BUFX16 U2 ( .A(n226), .Y(out[4]) );
  BUFX8 U3 ( .A(in_17bit[16]), .Y(n21) );
  CLKINVX3 U4 ( .A(n102), .Y(in_17bit_b[16]) );
  MXI2X4 U5 ( .A(n8), .B(n26), .S0(n185), .Y(out[13]) );
  NOR2X2 U6 ( .A(n41), .B(n79), .Y(n81) );
  INVX1 U7 ( .A(n58), .Y(n19) );
  INVX1 U8 ( .A(n88), .Y(n17) );
  INVX1 U9 ( .A(n174), .Y(n16) );
  XNOR2X2 U10 ( .A(n183), .B(n5), .Y(out[12]) );
  MX2X1 U11 ( .A(neg_mul[21]), .B(N479), .S0(n185), .Y(out[14]) );
  AOI22X1 U12 ( .A0(N27), .A1(n42), .B0(in_17bit[14]), .B1(n44), .Y(n113) );
  XNOR2X1 U13 ( .A(neg_mul[23]), .B(n28), .Y(n13) );
  CLKINVX3 U14 ( .A(n15), .Y(n42) );
  BUFX12 U15 ( .A(n225), .Y(out[5]) );
  BUFX8 U16 ( .A(n227), .Y(out[2]) );
  OAI21X4 U17 ( .A0(n41), .A1(n50), .B0(n49), .Y(n51) );
  INVXL U18 ( .A(n21), .Y(n15) );
  AND2X1 U19 ( .A(n40), .B(n16), .Y(n175) );
  NOR2X2 U20 ( .A(n21), .B(n97), .Y(n99) );
  AND2X2 U21 ( .A(n40), .B(n17), .Y(n90) );
  INVX8 U22 ( .A(n40), .Y(n41) );
  AND2X4 U23 ( .A(n40), .B(n19), .Y(n60) );
  XOR2X4 U24 ( .A(n180), .B(neg_mul[17]), .Y(out[10]) );
  INVXL U25 ( .A(in_8bit[0]), .Y(n38) );
  INVX4 U26 ( .A(n184), .Y(n185) );
  XNOR2X2 U27 ( .A(n21), .B(in_8bit[7]), .Y(n184) );
  XNOR2X2 U28 ( .A(n22), .B(in_8bit[7]), .Y(n181) );
  AOI211X2 U29 ( .A0(n21), .A1(n61), .B0(n60), .C0(n59), .Y(n227) );
  NOR2X4 U30 ( .A(n23), .B(n179), .Y(n180) );
  NOR2X4 U31 ( .A(n24), .B(n181), .Y(n182) );
  INVX8 U32 ( .A(in_17bit[16]), .Y(n40) );
  INVXL U33 ( .A(n42), .Y(n43) );
  INVXL U34 ( .A(n42), .Y(n44) );
  INVX8 U35 ( .A(n40), .Y(n22) );
  NOR2X4 U36 ( .A(n27), .B(n177), .Y(n178) );
  XNOR2X4 U37 ( .A(n41), .B(in_8bit[7]), .Y(n177) );
  OAI21X4 U38 ( .A0(n21), .A1(n68), .B0(n67), .Y(n69) );
  NOR2X2 U39 ( .A(n184), .B(n25), .Y(n183) );
  AOI211X4 U40 ( .A0(n41), .A1(n176), .B0(n175), .C0(n27), .Y(out[8]) );
  XNOR2X4 U41 ( .A(n22), .B(in_8bit[7]), .Y(n71) );
  XNOR2X2 U42 ( .A(n22), .B(in_8bit[7]), .Y(n179) );
  NOR2X4 U43 ( .A(n72), .B(n71), .Y(n73) );
  AOI21X4 U44 ( .A0(n41), .A1(n70), .B0(n69), .Y(out[3]) );
  INVX1 U45 ( .A(n152), .Y(in_17bit_b[1]) );
  INVX1 U46 ( .A(n113), .Y(in_17bit_b[14]) );
  INVX1 U47 ( .A(n116), .Y(in_17bit_b[13]) );
  INVX1 U48 ( .A(n149), .Y(in_17bit_b[2]) );
  INVX1 U49 ( .A(n140), .Y(in_17bit_b[5]) );
  INVX1 U50 ( .A(n137), .Y(in_17bit_b[6]) );
  INVX1 U51 ( .A(n134), .Y(in_17bit_b[7]) );
  INVX1 U52 ( .A(n131), .Y(in_17bit_b[8]) );
  INVX1 U53 ( .A(n128), .Y(in_17bit_b[9]) );
  INVX1 U54 ( .A(n125), .Y(in_17bit_b[10]) );
  INVX1 U55 ( .A(n122), .Y(in_17bit_b[11]) );
  INVX1 U56 ( .A(n119), .Y(in_17bit_b[12]) );
  INVX1 U57 ( .A(n143), .Y(in_17bit_b[4]) );
  INVX1 U58 ( .A(n146), .Y(in_17bit_b[3]) );
  AOI21X4 U59 ( .A0(n22), .A1(n52), .B0(n51), .Y(out[1]) );
  INVX1 U60 ( .A(n38), .Y(n37) );
  ADDFX2 U61 ( .A(in_17bit_b[16]), .B(in_17bit_b[12]), .CI(
        add_1_root_r112_carry_16_), .CO(add_1_root_r112_carry_17_), .S(
        add_1_root_r112_SUM_16_) );
  ADDFX2 U62 ( .A(add_1_root_r119_A_19_), .B(in_17bit_b[13]), .CI(
        add_1_root_r119_carry[19]), .CO(add_1_root_r119_carry[20]), .S(
        add_1_root_r119_SUM_19_) );
  ADDFX2 U63 ( .A(in_17bit_b[16]), .B(in_17bit_b[15]), .CI(
        add_3_root_r119_carry_17_), .CO(add_3_root_r119_carry_18_), .S(
        add_1_root_r119_A_17_) );
  ADDFX2 U64 ( .A(in_17bit_b[16]), .B(in_17bit_b[14]), .CI(
        add_2_root_r115_carry_17_), .CO(add_2_root_r115_carry_18_), .S(
        add_2_root_r115_SUM_17_) );
  ADDFX2 U65 ( .A(in_17bit_b[16]), .B(in_17bit_b[14]), .CI(
        add_1_root_r115_carry_20_), .CO(add_1_root_r115_carry_21_), .S(
        add_1_root_r115_SUM_20_) );
  ADDFX2 U66 ( .A(in_17bit_b[16]), .B(in_17bit_b[15]), .CI(
        add_2_root_r119_carry_20_), .CO(add_2_root_r119_carry_21_), .S(
        add_2_root_r119_SUM_20_) );
  ADDFX2 U67 ( .A(in_17bit_b[3]), .B(in_17bit_b[1]), .CI(
        add_1_root_r115_carry_7_), .CO(add_2_root_r115_carry_5_), .S(
        add_2_root_r115_SUM_4_) );
  ADDFX2 U68 ( .A(in_17bit_b[4]), .B(in_17bit_b[2]), .CI(
        add_2_root_r115_carry_5_), .CO(add_2_root_r115_carry_6_), .S(
        add_2_root_r115_SUM_5_) );
  ADDFX2 U69 ( .A(in_17bit_b[5]), .B(in_17bit_b[1]), .CI(
        add_1_root_r112_carry_5_), .CO(add_1_root_r112_carry_6_), .S(
        add_1_root_r112_SUM_5_) );
  ADDFX2 U70 ( .A(in_17bit_b[6]), .B(in_17bit_b[5]), .CI(
        add_3_root_r119_carry_7_), .CO(add_3_root_r119_carry_8_), .S(
        add_1_root_r119_A_7_) );
  ADDFX2 U71 ( .A(in_17bit_b[6]), .B(in_17bit_b[2]), .CI(
        add_1_root_r112_carry_6_), .CO(add_1_root_r112_carry_7_), .S(
        add_1_root_r112_SUM_6_) );
  ADDFX2 U72 ( .A(in_17bit_b[3]), .B(in_17bit_b[1]), .CI(
        add_1_root_r115_carry_7_), .CO(add_1_root_r115_carry_8_), .S(
        add_1_root_r115_SUM_7_) );
  ADDFX2 U73 ( .A(in_17bit_b[7]), .B(in_17bit_b[6]), .CI(
        add_3_root_r119_carry_8_), .CO(add_3_root_r119_carry_9_), .S(
        add_1_root_r119_A_8_) );
  ADDFX2 U74 ( .A(add_1_root_r119_A_7_), .B(in_17bit_b[1]), .CI(
        add_1_root_r119_carry[7]), .CO(add_1_root_r119_carry[8]), .S(
        add_1_root_r119_SUM_7_) );
  ADDFX2 U75 ( .A(in_17bit_b[2]), .B(in_17bit_b[1]), .CI(
        add_3_root_r119_carry_3_), .CO(add_2_root_r119_carry_7_), .S(
        add_2_root_r119_SUM_6_) );
  ADDFX2 U76 ( .A(in_17bit_b[4]), .B(in_17bit_b[2]), .CI(
        add_1_root_r115_carry_8_), .CO(add_1_root_r115_carry_9_), .S(
        add_1_root_r115_SUM_8_) );
  ADDFX2 U77 ( .A(in_17bit_b[8]), .B(in_17bit_b[7]), .CI(
        add_3_root_r119_carry_9_), .CO(add_3_root_r119_carry_10_), .S(
        add_1_root_r119_A_9_) );
  ADDFX2 U78 ( .A(add_1_root_r119_A_8_), .B(in_17bit_b[2]), .CI(
        add_1_root_r119_carry[8]), .CO(add_1_root_r119_carry[9]), .S(
        add_1_root_r119_SUM_8_) );
  ADDFX2 U79 ( .A(in_17bit_b[9]), .B(in_17bit_b[8]), .CI(
        add_3_root_r119_carry_10_), .CO(add_3_root_r119_carry_11_), .S(
        add_1_root_r119_A_10_) );
  ADDFX2 U80 ( .A(in_17bit_b[3]), .B(in_17bit_b[2]), .CI(
        add_2_root_r119_carry_7_), .CO(add_2_root_r119_carry_8_), .S(
        add_2_root_r119_SUM_7_) );
  ADDFX2 U81 ( .A(in_17bit_b[6]), .B(in_17bit_b[4]), .CI(
        add_2_root_r115_carry_7_), .CO(add_2_root_r115_carry_8_), .S(
        add_2_root_r115_SUM_7_) );
  ADDFX2 U82 ( .A(in_17bit_b[8]), .B(in_17bit_b[4]), .CI(
        add_1_root_r112_carry_8_), .CO(add_1_root_r112_carry_9_), .S(
        add_1_root_r112_SUM_8_) );
  ADDFX2 U83 ( .A(in_17bit_b[7]), .B(in_17bit_b[5]), .CI(
        add_2_root_r115_carry_8_), .CO(add_2_root_r115_carry_9_), .S(
        add_2_root_r115_SUM_8_) );
  ADDFX2 U84 ( .A(in_17bit_b[9]), .B(in_17bit_b[5]), .CI(
        add_1_root_r112_carry_9_), .CO(add_1_root_r112_carry_10_), .S(
        add_1_root_r112_SUM_9_) );
  ADDFX2 U85 ( .A(in_17bit_b[6]), .B(in_17bit_b[4]), .CI(
        add_1_root_r115_carry_10_), .CO(add_1_root_r115_carry_11_), .S(
        add_1_root_r115_SUM_10_) );
  ADDFX2 U86 ( .A(in_17bit_b[10]), .B(in_17bit_b[9]), .CI(
        add_3_root_r119_carry_11_), .CO(add_3_root_r119_carry_12_), .S(
        add_1_root_r119_A_11_) );
  ADDFX2 U87 ( .A(in_17bit_b[10]), .B(in_17bit_b[6]), .CI(
        add_1_root_r112_carry_10_), .CO(add_1_root_r112_carry_11_), .S(
        add_1_root_r112_SUM_10_) );
  ADDFX2 U88 ( .A(in_17bit_b[7]), .B(in_17bit_b[5]), .CI(
        add_1_root_r115_carry_11_), .CO(add_1_root_r115_carry_12_), .S(
        add_1_root_r115_SUM_11_) );
  ADDFX2 U89 ( .A(in_17bit_b[11]), .B(in_17bit_b[10]), .CI(
        add_3_root_r119_carry_12_), .CO(add_3_root_r119_carry_13_), .S(
        add_1_root_r119_A_12_) );
  ADDFX2 U90 ( .A(add_1_root_r119_A_11_), .B(in_17bit_b[5]), .CI(
        add_1_root_r119_carry[11]), .CO(add_1_root_r119_carry[12]), .S(
        add_1_root_r119_SUM_11_) );
  ADDFX2 U91 ( .A(in_17bit_b[6]), .B(in_17bit_b[5]), .CI(
        add_2_root_r119_carry_10_), .CO(add_2_root_r119_carry_11_), .S(
        add_2_root_r119_SUM_10_) );
  ADDFX2 U92 ( .A(in_17bit_b[9]), .B(in_17bit_b[7]), .CI(
        add_2_root_r115_carry_10_), .CO(add_2_root_r115_carry_11_), .S(
        add_2_root_r115_SUM_10_) );
  ADDFX2 U93 ( .A(in_17bit_b[11]), .B(in_17bit_b[7]), .CI(
        add_1_root_r112_carry_11_), .CO(add_1_root_r112_carry_12_), .S(
        add_1_root_r112_SUM_11_) );
  ADDFX2 U94 ( .A(in_17bit_b[8]), .B(in_17bit_b[6]), .CI(
        add_1_root_r115_carry_12_), .CO(add_1_root_r115_carry_13_), .S(
        add_1_root_r115_SUM_12_) );
  ADDFX2 U95 ( .A(in_17bit_b[12]), .B(in_17bit_b[11]), .CI(
        add_3_root_r119_carry_13_), .CO(add_3_root_r119_carry_14_), .S(
        add_1_root_r119_A_13_) );
  ADDFX2 U96 ( .A(add_1_root_r119_A_12_), .B(in_17bit_b[6]), .CI(
        add_1_root_r119_carry[12]), .CO(add_1_root_r119_carry[13]), .S(
        add_1_root_r119_SUM_12_) );
  ADDFX2 U97 ( .A(in_17bit_b[7]), .B(in_17bit_b[6]), .CI(
        add_2_root_r119_carry_11_), .CO(add_2_root_r119_carry_12_), .S(
        add_2_root_r119_SUM_11_) );
  ADDFX2 U98 ( .A(in_17bit_b[10]), .B(in_17bit_b[8]), .CI(
        add_2_root_r115_carry_11_), .CO(add_2_root_r115_carry_12_), .S(
        add_2_root_r115_SUM_11_) );
  ADDFX2 U99 ( .A(in_17bit_b[12]), .B(in_17bit_b[8]), .CI(
        add_1_root_r112_carry_12_), .CO(add_1_root_r112_carry_13_), .S(
        add_1_root_r112_SUM_12_) );
  ADDFX2 U100 ( .A(in_17bit_b[9]), .B(in_17bit_b[7]), .CI(
        add_1_root_r115_carry_13_), .CO(add_1_root_r115_carry_14_), .S(
        add_1_root_r115_SUM_13_) );
  ADDFX2 U101 ( .A(in_17bit_b[13]), .B(in_17bit_b[12]), .CI(
        add_3_root_r119_carry_14_), .CO(add_3_root_r119_carry_15_), .S(
        add_1_root_r119_A_14_) );
  ADDFX2 U102 ( .A(add_1_root_r119_A_13_), .B(in_17bit_b[7]), .CI(
        add_1_root_r119_carry[13]), .CO(add_1_root_r119_carry[14]), .S(
        add_1_root_r119_SUM_13_) );
  ADDFX2 U103 ( .A(in_17bit_b[8]), .B(in_17bit_b[7]), .CI(
        add_2_root_r119_carry_12_), .CO(add_2_root_r119_carry_13_), .S(
        add_2_root_r119_SUM_12_) );
  ADDFX2 U104 ( .A(in_17bit_b[11]), .B(in_17bit_b[9]), .CI(
        add_2_root_r115_carry_12_), .CO(add_2_root_r115_carry_13_), .S(
        add_2_root_r115_SUM_12_) );
  ADDFX2 U105 ( .A(in_17bit_b[14]), .B(in_17bit_b[13]), .CI(
        add_3_root_r119_carry_15_), .CO(add_3_root_r119_carry_16_), .S(
        add_1_root_r119_A_15_) );
  ADDFX2 U106 ( .A(add_1_root_r119_A_14_), .B(in_17bit_b[8]), .CI(
        add_1_root_r119_carry[14]), .CO(add_1_root_r119_carry[15]), .S(
        add_1_root_r119_SUM_14_) );
  ADDFX2 U107 ( .A(in_17bit_b[9]), .B(in_17bit_b[8]), .CI(
        add_2_root_r119_carry_13_), .CO(add_2_root_r119_carry_14_), .S(
        add_2_root_r119_SUM_13_) );
  ADDFX2 U108 ( .A(in_17bit_b[12]), .B(in_17bit_b[10]), .CI(
        add_2_root_r115_carry_13_), .CO(add_2_root_r115_carry_14_), .S(
        add_2_root_r115_SUM_13_) );
  ADDFX2 U109 ( .A(in_17bit_b[14]), .B(in_17bit_b[10]), .CI(
        add_1_root_r112_carry_14_), .CO(add_1_root_r112_carry_15_), .S(
        add_1_root_r112_SUM_14_) );
  ADDFX2 U110 ( .A(in_17bit_b[11]), .B(in_17bit_b[9]), .CI(
        add_1_root_r115_carry_15_), .CO(add_1_root_r115_carry_16_), .S(
        add_1_root_r115_SUM_15_) );
  ADDFX2 U111 ( .A(add_1_root_r119_A_15_), .B(in_17bit_b[9]), .CI(
        add_1_root_r119_carry[15]), .CO(add_1_root_r119_carry[16]), .S(
        add_1_root_r119_SUM_15_) );
  ADDFX2 U112 ( .A(in_17bit_b[10]), .B(in_17bit_b[9]), .CI(
        add_2_root_r119_carry_14_), .CO(add_2_root_r119_carry_15_), .S(
        add_2_root_r119_SUM_14_) );
  ADDFX2 U113 ( .A(in_17bit_b[13]), .B(in_17bit_b[11]), .CI(
        add_2_root_r115_carry_14_), .CO(add_2_root_r115_carry_15_), .S(
        add_2_root_r115_SUM_14_) );
  ADDFX2 U114 ( .A(in_17bit_b[15]), .B(in_17bit_b[11]), .CI(
        add_1_root_r112_carry_15_), .CO(add_1_root_r112_carry_16_), .S(
        add_1_root_r112_SUM_15_) );
  ADDFX2 U115 ( .A(in_17bit_b[12]), .B(in_17bit_b[10]), .CI(
        add_1_root_r115_carry_16_), .CO(add_1_root_r115_carry_17_), .S(
        add_1_root_r115_SUM_16_) );
  ADDFX2 U116 ( .A(add_1_root_r119_A_16_), .B(in_17bit_b[10]), .CI(
        add_1_root_r119_carry[16]), .CO(add_1_root_r119_carry[17]), .S(
        add_1_root_r119_SUM_16_) );
  ADDFX2 U117 ( .A(in_17bit_b[11]), .B(in_17bit_b[10]), .CI(
        add_2_root_r119_carry_15_), .CO(add_2_root_r119_carry_16_), .S(
        add_2_root_r119_SUM_15_) );
  ADDFX2 U118 ( .A(in_17bit_b[14]), .B(in_17bit_b[12]), .CI(
        add_2_root_r115_carry_15_), .CO(add_2_root_r115_carry_16_), .S(
        add_2_root_r115_SUM_15_) );
  ADDFX2 U119 ( .A(in_17bit_b[13]), .B(in_17bit_b[11]), .CI(
        add_1_root_r115_carry_17_), .CO(add_1_root_r115_carry_18_), .S(
        add_1_root_r115_SUM_17_) );
  ADDFX2 U120 ( .A(add_1_root_r119_A_17_), .B(in_17bit_b[11]), .CI(
        add_1_root_r119_carry[17]), .CO(add_1_root_r119_carry[18]), .S(
        add_1_root_r119_SUM_17_) );
  ADDFX2 U121 ( .A(in_17bit_b[12]), .B(in_17bit_b[11]), .CI(
        add_2_root_r119_carry_16_), .CO(add_2_root_r119_carry_17_), .S(
        add_2_root_r119_SUM_16_) );
  ADDFX2 U122 ( .A(in_17bit_b[15]), .B(in_17bit_b[13]), .CI(
        add_2_root_r115_carry_16_), .CO(add_2_root_r115_carry_17_), .S(
        add_2_root_r115_SUM_16_) );
  ADDFX2 U123 ( .A(in_17bit_b[14]), .B(in_17bit_b[12]), .CI(
        add_1_root_r115_carry_18_), .CO(add_1_root_r115_carry_19_), .S(
        add_1_root_r115_SUM_18_) );
  ADDFX2 U124 ( .A(add_1_root_r119_A_18_), .B(in_17bit_b[12]), .CI(
        add_1_root_r119_carry[18]), .CO(add_1_root_r119_carry[19]), .S(
        add_1_root_r119_SUM_18_) );
  ADDFX2 U125 ( .A(in_17bit_b[15]), .B(in_17bit_b[13]), .CI(
        add_1_root_r115_carry_19_), .CO(add_1_root_r115_carry_20_), .S(
        add_1_root_r115_SUM_19_) );
  ADDFX2 U126 ( .A(in_17bit_b[7]), .B(in_17bit_b[3]), .CI(
        add_1_root_r112_carry_7_), .CO(add_1_root_r112_carry_8_), .S(
        add_1_root_r112_SUM_7_) );
  ADDFX2 U127 ( .A(in_17bit_b[5]), .B(in_17bit_b[3]), .CI(
        add_1_root_r115_carry_9_), .CO(add_1_root_r115_carry_10_), .S(
        add_1_root_r115_SUM_9_) );
  ADDFX2 U128 ( .A(add_1_root_r119_A_9_), .B(in_17bit_b[3]), .CI(
        add_1_root_r119_carry[9]), .CO(add_1_root_r119_carry[10]), .S(
        add_1_root_r119_SUM_9_) );
  ADDFX2 U129 ( .A(in_17bit_b[4]), .B(in_17bit_b[3]), .CI(
        add_2_root_r119_carry_8_), .CO(add_2_root_r119_carry_9_), .S(
        add_2_root_r119_SUM_8_) );
  ADDFX2 U130 ( .A(add_1_root_r119_A_10_), .B(in_17bit_b[4]), .CI(
        add_1_root_r119_carry[10]), .CO(add_1_root_r119_carry[11]), .S(
        add_1_root_r119_SUM_10_) );
  ADDFX2 U131 ( .A(in_17bit_b[5]), .B(in_17bit_b[4]), .CI(
        add_2_root_r119_carry_9_), .CO(add_2_root_r119_carry_10_), .S(
        add_2_root_r119_SUM_9_) );
  ADDFX2 U132 ( .A(in_17bit_b[8]), .B(in_17bit_b[6]), .CI(
        add_2_root_r115_carry_9_), .CO(add_2_root_r115_carry_10_), .S(
        add_2_root_r115_SUM_9_) );
  ADDFX2 U133 ( .A(in_17bit_b[13]), .B(in_17bit_b[9]), .CI(
        add_1_root_r112_carry_13_), .CO(add_1_root_r112_carry_14_), .S(
        add_1_root_r112_SUM_13_) );
  ADDFX2 U134 ( .A(in_17bit_b[10]), .B(in_17bit_b[8]), .CI(
        add_1_root_r115_carry_14_), .CO(add_1_root_r115_carry_15_), .S(
        add_1_root_r115_SUM_14_) );
  ADDFX2 U135 ( .A(in_17bit_b[13]), .B(in_17bit_b[12]), .CI(
        add_2_root_r119_carry_17_), .CO(add_2_root_r119_carry_18_), .S(
        add_2_root_r119_SUM_17_) );
  ADDFX2 U136 ( .A(in_17bit_b[15]), .B(in_17bit_b[14]), .CI(
        add_3_root_r119_carry_16_), .CO(add_3_root_r119_carry_17_), .S(
        add_1_root_r119_A_16_) );
  ADDFX2 U137 ( .A(in_17bit_b[3]), .B(in_17bit_b[2]), .CI(
        add_3_root_r119_carry_4_), .CO(add_3_root_r119_carry_5_), .S(
        add_1_root_r119_A_4_) );
  ADDFX2 U138 ( .A(in_17bit_b[2]), .B(in_17bit_b[1]), .CI(
        add_3_root_r119_carry_3_), .CO(add_3_root_r119_carry_4_), .S(
        add_1_root_r119_A_3_) );
  ADDFX2 U139 ( .A(in_17bit_b[4]), .B(in_17bit_b[3]), .CI(
        add_3_root_r119_carry_5_), .CO(add_3_root_r119_carry_6_), .S(
        add_1_root_r119_A_5_) );
  ADDFX2 U140 ( .A(in_17bit_b[5]), .B(in_17bit_b[4]), .CI(
        add_3_root_r119_carry_6_), .CO(add_3_root_r119_carry_7_), .S(
        add_1_root_r119_A_6_) );
  ADDFX2 U141 ( .A(in_17bit_b[14]), .B(in_17bit_b[13]), .CI(
        add_2_root_r119_carry_18_), .CO(add_2_root_r119_carry_19_), .S(
        add_2_root_r119_SUM_18_) );
  ADDFX2 U142 ( .A(in_17bit_b[5]), .B(in_17bit_b[3]), .CI(
        add_2_root_r115_carry_6_), .CO(add_2_root_r115_carry_7_), .S(
        add_2_root_r115_SUM_6_) );
  ADDFX2 U143 ( .A(in_17bit_b[15]), .B(in_17bit_b[14]), .CI(
        add_2_root_r119_carry_19_), .CO(add_2_root_r119_carry_20_), .S(
        add_2_root_r119_SUM_19_) );
  INVX1 U144 ( .A(in_8bit[2]), .Y(n39) );
  NOR3X1 U145 ( .A(n39), .B(n205), .C(n38), .Y(n157) );
  CLKINVX3 U146 ( .A(n155), .Y(in_17bit_b[0]) );
  INVX1 U147 ( .A(n103), .Y(n202) );
  OAI21XL U148 ( .A0(n103), .A1(n102), .B0(n104), .Y(N463) );
  AOI22X1 U149 ( .A0(N221), .A1(n35), .B0(N363), .B1(n34), .Y(n104) );
  NAND2XL U150 ( .A(N29), .B(n42), .Y(n102) );
  CLKINVX3 U151 ( .A(n110), .Y(in_17bit_b[15]) );
  BUFX3 U152 ( .A(in_8bit[1]), .Y(n36) );
  MXI2XL U153 ( .A(n1), .B(n13), .S0(n185), .Y(out[16]) );
  AOI32X1 U154 ( .A0(n157), .A1(n203), .A2(in_8bit[5]), .B0(n158), .B1(n159), 
        .Y(n103) );
  INVX1 U155 ( .A(n160), .Y(n203) );
  INVXL U156 ( .A(in_8bit[3]), .Y(n205) );
  NAND3BXL U157 ( .AN(in_8bit[5]), .B(n39), .C(in_8bit[3]), .Y(n166) );
  NOR4BX1 U158 ( .AN(n165), .B(n38), .C(n36), .D(in_8bit[2]), .Y(n159) );
  NOR2XL U159 ( .A(in_8bit[6]), .B(in_8bit[3]), .Y(n165) );
  AOI22XL U160 ( .A0(in_17bit[0]), .A1(n42), .B0(in_17bit[0]), .B1(n44), .Y(
        n155) );
  NAND3X1 U161 ( .A(in_8bit[2]), .B(n205), .C(in_8bit[5]), .Y(n167) );
  AOI22XL U162 ( .A0(N26), .A1(n42), .B0(in_17bit[13]), .B1(n43), .Y(n116) );
  AOI22XL U163 ( .A0(N14), .A1(n42), .B0(in_17bit[1]), .B1(n44), .Y(n152) );
  AOI22XL U164 ( .A0(N15), .A1(n42), .B0(in_17bit[2]), .B1(n43), .Y(n149) );
  AOI22XL U165 ( .A0(N16), .A1(n42), .B0(in_17bit[3]), .B1(n15), .Y(n146) );
  AOI22XL U166 ( .A0(N18), .A1(n42), .B0(in_17bit[5]), .B1(n44), .Y(n140) );
  AOI22XL U167 ( .A0(N19), .A1(n42), .B0(in_17bit[6]), .B1(n15), .Y(n137) );
  AOI22XL U168 ( .A0(N20), .A1(n42), .B0(in_17bit[7]), .B1(n15), .Y(n134) );
  AOI22XL U169 ( .A0(N21), .A1(n42), .B0(in_17bit[8]), .B1(n44), .Y(n131) );
  AOI22XL U170 ( .A0(N22), .A1(n42), .B0(in_17bit[9]), .B1(n43), .Y(n128) );
  AOI22XL U171 ( .A0(N23), .A1(n42), .B0(in_17bit[10]), .B1(n43), .Y(n125) );
  AOI22XL U172 ( .A0(N24), .A1(n42), .B0(in_17bit[11]), .B1(n15), .Y(n122) );
  AOI22XL U173 ( .A0(N25), .A1(n42), .B0(in_17bit[12]), .B1(n44), .Y(n119) );
  AOI22XL U174 ( .A0(N28), .A1(n42), .B0(in_17bit[15]), .B1(n43), .Y(n110) );
  INVX1 U175 ( .A(n67), .Y(n72) );
  AND2X2 U176 ( .A(n27), .B(n3), .Y(n23) );
  AND2X2 U177 ( .A(n23), .B(n12), .Y(n24) );
  BUFX3 U178 ( .A(n106), .Y(n34) );
  OAI32X1 U179 ( .A0(n167), .A1(n37), .A2(n160), .B0(n166), .B1(n168), .Y(n106) );
  BUFX3 U180 ( .A(n105), .Y(n35) );
  OAI32X1 U181 ( .A0(n160), .A1(n37), .A2(n166), .B0(n167), .B1(n168), .Y(n105) );
  INVX1 U182 ( .A(n49), .Y(n53) );
  NAND2X1 U183 ( .A(n72), .B(n2), .Y(n74) );
  INVX1 U184 ( .A(n83), .Y(n80) );
  INVX1 U185 ( .A(n92), .Y(n89) );
  INVX1 U186 ( .A(n101), .Y(n98) );
  AND2X2 U187 ( .A(n24), .B(n4), .Y(n25) );
  INVX1 U188 ( .A(in_17bit[0]), .Y(n186) );
  INVX1 U189 ( .A(in_17bit[1]), .Y(n187) );
  INVX1 U190 ( .A(in_17bit[2]), .Y(n188) );
  INVX1 U191 ( .A(in_17bit[3]), .Y(n189) );
  INVX1 U192 ( .A(in_17bit[6]), .Y(n192) );
  INVX1 U193 ( .A(in_17bit[7]), .Y(n193) );
  INVX1 U194 ( .A(in_17bit[8]), .Y(n194) );
  INVX1 U195 ( .A(in_17bit[9]), .Y(n195) );
  INVX1 U196 ( .A(in_17bit[10]), .Y(n196) );
  INVX1 U197 ( .A(in_17bit[11]), .Y(n197) );
  INVX1 U198 ( .A(in_17bit[12]), .Y(n198) );
  INVX1 U199 ( .A(in_17bit[13]), .Y(n199) );
  INVX1 U200 ( .A(in_17bit[14]), .Y(n200) );
  INVX1 U201 ( .A(in_17bit[15]), .Y(n201) );
  INVX1 U202 ( .A(in_17bit[5]), .Y(n191) );
  INVX1 U203 ( .A(in_17bit[4]), .Y(n190) );
  NAND2X1 U204 ( .A(n153), .B(n154), .Y(N447) );
  AOI22X1 U205 ( .A0(N108), .A1(n109), .B0(N205), .B1(n35), .Y(n154) );
  AOI22X1 U206 ( .A0(N347), .A1(n34), .B0(n202), .B1(in_17bit_b[0]), .Y(n153)
         );
  NAND2X1 U207 ( .A(n150), .B(n151), .Y(N448) );
  AOI22X1 U208 ( .A0(N109), .A1(n109), .B0(N206), .B1(n35), .Y(n151) );
  AOI22X1 U209 ( .A0(N348), .A1(n34), .B0(n202), .B1(in_17bit_b[1]), .Y(n150)
         );
  NAND2X1 U210 ( .A(n147), .B(n148), .Y(N449) );
  AOI22X1 U211 ( .A0(N110), .A1(n109), .B0(N207), .B1(n35), .Y(n148) );
  AOI22X1 U212 ( .A0(N349), .A1(n34), .B0(n202), .B1(in_17bit_b[2]), .Y(n147)
         );
  NAND2X1 U213 ( .A(n144), .B(n145), .Y(N450) );
  AOI22X1 U214 ( .A0(N111), .A1(n109), .B0(N208), .B1(n35), .Y(n145) );
  AOI22X1 U215 ( .A0(N350), .A1(n34), .B0(n202), .B1(in_17bit_b[3]), .Y(n144)
         );
  NAND2X1 U216 ( .A(n141), .B(n142), .Y(N451) );
  AOI22X1 U217 ( .A0(N112), .A1(n109), .B0(N209), .B1(n35), .Y(n142) );
  AOI22X1 U218 ( .A0(N351), .A1(n34), .B0(n202), .B1(in_17bit_b[4]), .Y(n141)
         );
  NAND2X1 U219 ( .A(n138), .B(n139), .Y(N452) );
  AOI22X1 U220 ( .A0(N113), .A1(n109), .B0(N210), .B1(n35), .Y(n139) );
  AOI22X1 U221 ( .A0(N352), .A1(n34), .B0(n202), .B1(in_17bit_b[5]), .Y(n138)
         );
  NAND2X1 U222 ( .A(n135), .B(n136), .Y(N453) );
  AOI22X1 U223 ( .A0(N114), .A1(n109), .B0(N211), .B1(n35), .Y(n136) );
  AOI22X1 U224 ( .A0(N353), .A1(n34), .B0(n202), .B1(in_17bit_b[6]), .Y(n135)
         );
  NAND2X1 U225 ( .A(n132), .B(n133), .Y(N454) );
  AOI22X1 U226 ( .A0(N115), .A1(n109), .B0(N212), .B1(n35), .Y(n133) );
  AOI22X1 U227 ( .A0(N354), .A1(n34), .B0(n202), .B1(in_17bit_b[7]), .Y(n132)
         );
  NAND2X1 U228 ( .A(n129), .B(n130), .Y(N455) );
  AOI22X1 U229 ( .A0(N116), .A1(n109), .B0(N213), .B1(n35), .Y(n130) );
  AOI22X1 U230 ( .A0(N355), .A1(n34), .B0(n202), .B1(in_17bit_b[8]), .Y(n129)
         );
  NAND2X1 U231 ( .A(n126), .B(n127), .Y(N456) );
  AOI22X1 U232 ( .A0(N117), .A1(n109), .B0(N214), .B1(n35), .Y(n127) );
  AOI22X1 U233 ( .A0(N356), .A1(n34), .B0(n202), .B1(in_17bit_b[9]), .Y(n126)
         );
  NAND2X1 U234 ( .A(n123), .B(n124), .Y(N457) );
  AOI22X1 U235 ( .A0(N118), .A1(n109), .B0(N215), .B1(n35), .Y(n124) );
  AOI22X1 U236 ( .A0(N357), .A1(n34), .B0(n202), .B1(in_17bit_b[10]), .Y(n123)
         );
  NAND2X1 U237 ( .A(n120), .B(n121), .Y(N458) );
  AOI22X1 U238 ( .A0(N119), .A1(n109), .B0(N216), .B1(n35), .Y(n121) );
  AOI22X1 U239 ( .A0(N358), .A1(n34), .B0(n202), .B1(in_17bit_b[11]), .Y(n120)
         );
  NAND2X1 U240 ( .A(n117), .B(n118), .Y(N459) );
  AOI22X1 U241 ( .A0(N120), .A1(n109), .B0(N217), .B1(n35), .Y(n118) );
  AOI22X1 U242 ( .A0(N359), .A1(n34), .B0(n202), .B1(in_17bit_b[12]), .Y(n117)
         );
  NAND2X1 U243 ( .A(n114), .B(n115), .Y(N460) );
  AOI22X1 U244 ( .A0(N121), .A1(n109), .B0(N218), .B1(n35), .Y(n115) );
  AOI22X1 U245 ( .A0(N360), .A1(n34), .B0(n202), .B1(in_17bit_b[13]), .Y(n114)
         );
  NAND2X1 U246 ( .A(n111), .B(n112), .Y(N461) );
  AOI22X1 U247 ( .A0(N122), .A1(n109), .B0(N219), .B1(n35), .Y(n112) );
  AOI22X1 U248 ( .A0(N361), .A1(n34), .B0(n202), .B1(in_17bit_b[14]), .Y(n111)
         );
  NAND2X1 U249 ( .A(n107), .B(n108), .Y(N462) );
  AOI22X1 U250 ( .A0(N123), .A1(n109), .B0(N220), .B1(n35), .Y(n108) );
  AOI22X1 U251 ( .A0(N362), .A1(n34), .B0(n202), .B1(in_17bit_b[15]), .Y(n107)
         );
  OAI21XL U252 ( .A0(in_8bit[7]), .A1(n171), .B0(n170), .Y(n176) );
  NAND2BX1 U253 ( .AN(neg_mul[15]), .B(in_8bit[7]), .Y(n170) );
  XNOR2X1 U254 ( .A(n8), .B(sub_add_75_b0_carry[13]), .Y(n26) );
  OAI21XL U255 ( .A0(in_8bit[7]), .A1(n46), .B0(n45), .Y(n52) );
  NAND2BX1 U256 ( .AN(neg_mul[8]), .B(in_8bit[7]), .Y(n45) );
  OAI21XL U257 ( .A0(in_8bit[7]), .A1(n64), .B0(n63), .Y(n70) );
  NAND2BX1 U258 ( .AN(neg_mul[10]), .B(in_8bit[7]), .Y(n63) );
  OAI21XL U259 ( .A0(in_8bit[7]), .A1(n76), .B0(n75), .Y(n82) );
  NAND2BX1 U260 ( .AN(neg_mul[12]), .B(in_8bit[7]), .Y(n75) );
  OAI21XL U261 ( .A0(in_8bit[7]), .A1(n85), .B0(n84), .Y(n91) );
  NAND2BX1 U262 ( .AN(neg_mul[13]), .B(in_8bit[7]), .Y(n84) );
  INVX1 U263 ( .A(n62), .Y(n59) );
  OAI21XL U264 ( .A0(in_8bit[7]), .A1(n55), .B0(n54), .Y(n61) );
  OAI21XL U265 ( .A0(in_8bit[7]), .A1(n94), .B0(n93), .Y(n100) );
  NAND2BX1 U266 ( .AN(neg_mul[14]), .B(in_8bit[7]), .Y(n93) );
  MX2X1 U267 ( .A(neg_mul[22]), .B(N480), .S0(n185), .Y(out[15]) );
  NAND4BBX1 U268 ( .AN(n34), .BN(n35), .C(n156), .D(n103), .Y(N446) );
  AOI2BB1X1 U269 ( .A0N(n161), .A1N(n162), .B0(n109), .Y(n156) );
  OR4X2 U270 ( .A(in_8bit[4]), .B(in_8bit[5]), .C(in_8bit[6]), .D(in_8bit[7]), 
        .Y(n161) );
  OR4XL U271 ( .A(n36), .B(n37), .C(in_8bit[2]), .D(in_8bit[3]), .Y(n162) );
  NOR3X1 U272 ( .A(in_8bit[4]), .B(in_8bit[5]), .C(n204), .Y(n158) );
  NAND4X1 U273 ( .A(in_8bit[6]), .B(in_8bit[4]), .C(n36), .D(n204), .Y(n160)
         );
  NOR2BX1 U274 ( .AN(n98), .B(neg_mul[15]), .Y(n27) );
  NAND4X1 U275 ( .A(n36), .B(in_8bit[7]), .C(n169), .D(n38), .Y(n168) );
  NOR2X1 U276 ( .A(in_8bit[6]), .B(in_8bit[4]), .Y(n169) );
  NAND2X1 U277 ( .A(n53), .B(n11), .Y(n62) );
  NAND2X1 U278 ( .A(out[0]), .B(neg_mul[8]), .Y(n46) );
  NAND2X1 U279 ( .A(neg_mul[10]), .B(n62), .Y(n64) );
  NAND2X1 U280 ( .A(neg_mul[12]), .B(n74), .Y(n76) );
  NAND2X1 U281 ( .A(neg_mul[14]), .B(n92), .Y(n94) );
  NAND2BX1 U282 ( .AN(n53), .B(neg_mul[9]), .Y(n55) );
  AOI21X1 U283 ( .A0(n173), .A1(in_8bit[7]), .B0(n172), .Y(n174) );
  INVX1 U284 ( .A(n171), .Y(n173) );
  NOR2X1 U285 ( .A(in_8bit[7]), .B(neg_mul[15]), .Y(n172) );
  AOI21X1 U286 ( .A0(n87), .A1(in_8bit[7]), .B0(n86), .Y(n88) );
  INVX1 U287 ( .A(n85), .Y(n87) );
  NOR2X1 U288 ( .A(in_8bit[7]), .B(neg_mul[13]), .Y(n86) );
  NAND2X1 U289 ( .A(n163), .B(n164), .Y(n109) );
  NAND4X1 U290 ( .A(n158), .B(n157), .C(in_8bit[6]), .D(n36), .Y(n164) );
  NAND4X1 U291 ( .A(n159), .B(in_8bit[5]), .C(in_8bit[4]), .D(n204), .Y(n163)
         );
  NAND2X1 U292 ( .A(neg_mul[15]), .B(n101), .Y(n171) );
  NAND2X1 U293 ( .A(neg_mul[13]), .B(n83), .Y(n85) );
  OR2X2 U294 ( .A(n62), .B(neg_mul[10]), .Y(n67) );
  OR2X2 U295 ( .A(n74), .B(neg_mul[12]), .Y(n83) );
  NAND2X1 U296 ( .A(n80), .B(n9), .Y(n92) );
  NAND2X1 U297 ( .A(n89), .B(n10), .Y(n101) );
  NOR2X1 U298 ( .A(n48), .B(n47), .Y(n50) );
  NOR2X1 U299 ( .A(in_8bit[7]), .B(neg_mul[8]), .Y(n47) );
  NOR2X1 U300 ( .A(n204), .B(n46), .Y(n48) );
  NOR2X1 U301 ( .A(n66), .B(n65), .Y(n68) );
  NOR2X1 U302 ( .A(in_8bit[7]), .B(neg_mul[10]), .Y(n65) );
  NOR2X1 U303 ( .A(n204), .B(n64), .Y(n66) );
  NOR2X1 U304 ( .A(n78), .B(n77), .Y(n79) );
  NOR2X1 U305 ( .A(in_8bit[7]), .B(neg_mul[12]), .Y(n77) );
  NOR2X1 U306 ( .A(n204), .B(n76), .Y(n78) );
  NOR2X1 U307 ( .A(n96), .B(n95), .Y(n97) );
  NOR2X1 U308 ( .A(in_8bit[7]), .B(neg_mul[14]), .Y(n95) );
  NOR2X1 U309 ( .A(n204), .B(n94), .Y(n96) );
  AOI21X1 U310 ( .A0(n57), .A1(in_8bit[7]), .B0(n56), .Y(n58) );
  INVX1 U311 ( .A(n55), .Y(n57) );
  NOR2X1 U312 ( .A(in_8bit[7]), .B(neg_mul[9]), .Y(n56) );
  OR2X2 U313 ( .A(out[0]), .B(neg_mul[8]), .Y(n49) );
  NAND2X1 U314 ( .A(sub_add_75_b0_carry[15]), .B(n6), .Y(n28) );
  NAND2BX1 U315 ( .AN(neg_mul[9]), .B(in_8bit[7]), .Y(n54) );
  INVX1 U316 ( .A(in_8bit[7]), .Y(n204) );
  AOI211X4 U317 ( .A0(n22), .A1(n91), .B0(n90), .C0(n89), .Y(out[6]) );
  AOI211X4 U318 ( .A0(n41), .A1(n100), .B0(n99), .C0(n98), .Y(out[7]) );
  AOI22XL U319 ( .A0(N17), .A1(n42), .B0(in_17bit[4]), .B1(n43), .Y(n143) );
  AOI211X4 U320 ( .A0(n22), .A1(n82), .B0(n81), .C0(n80), .Y(n225) );
  XNOR2X4 U321 ( .A(n73), .B(n2), .Y(n226) );
  XNOR2X4 U322 ( .A(n178), .B(n3), .Y(out[9]) );
  XNOR2X4 U323 ( .A(n182), .B(n4), .Y(out[11]) );
  AND2X1 U324 ( .A(add_1_root_r112_carry_20_), .B(in_17bit_b[16]), .Y(
        add_1_root_r112_SUM_21_) );
  XOR2X1 U325 ( .A(in_17bit_b[16]), .B(add_1_root_r112_carry_20_), .Y(
        add_1_root_r112_SUM_20_) );
  AND2X1 U326 ( .A(add_1_root_r112_carry_19_), .B(in_17bit_b[15]), .Y(
        add_1_root_r112_carry_20_) );
  XOR2X1 U327 ( .A(in_17bit_b[15]), .B(add_1_root_r112_carry_19_), .Y(
        add_1_root_r112_SUM_19_) );
  AND2X1 U328 ( .A(add_1_root_r112_carry_18_), .B(in_17bit_b[14]), .Y(
        add_1_root_r112_carry_19_) );
  XOR2X1 U329 ( .A(in_17bit_b[14]), .B(add_1_root_r112_carry_18_), .Y(
        add_1_root_r112_SUM_18_) );
  AND2X1 U330 ( .A(add_1_root_r112_carry_17_), .B(in_17bit_b[13]), .Y(
        add_1_root_r112_carry_18_) );
  XOR2X1 U331 ( .A(in_17bit_b[13]), .B(add_1_root_r112_carry_17_), .Y(
        add_1_root_r112_SUM_17_) );
  AND2X1 U332 ( .A(add_2_root_r119_carry_21_), .B(in_17bit_b[16]), .Y(
        add_2_root_r119_SUM_22_) );
  XOR2X1 U333 ( .A(in_17bit_b[16]), .B(add_2_root_r119_carry_21_), .Y(
        add_2_root_r119_SUM_21_) );
  XOR2X1 U334 ( .A(in_17bit_b[0]), .B(in_17bit_b[1]), .Y(
        add_2_root_r119_SUM_5_) );
  AND2X1 U335 ( .A(add_1_root_r119_carry[22]), .B(in_17bit_b[16]), .Y(
        add_1_root_r119_SUM_23_) );
  XOR2X1 U336 ( .A(in_17bit_b[16]), .B(add_1_root_r119_carry[22]), .Y(
        add_1_root_r119_SUM_22_) );
  AND2X1 U337 ( .A(add_1_root_r119_carry[21]), .B(in_17bit_b[15]), .Y(
        add_1_root_r119_carry[22]) );
  XOR2X1 U338 ( .A(in_17bit_b[15]), .B(add_1_root_r119_carry[21]), .Y(
        add_1_root_r119_SUM_21_) );
  AND2X1 U339 ( .A(add_1_root_r119_carry[20]), .B(in_17bit_b[14]), .Y(
        add_1_root_r119_carry[21]) );
  XOR2X1 U340 ( .A(in_17bit_b[14]), .B(add_1_root_r119_carry[20]), .Y(
        add_1_root_r119_SUM_20_) );
  AND2X1 U341 ( .A(add_1_root_r119_A_6_), .B(in_17bit_b[0]), .Y(
        add_1_root_r119_carry[7]) );
  XOR2X1 U342 ( .A(in_17bit_b[0]), .B(add_1_root_r119_A_6_), .Y(
        add_1_root_r119_SUM_6_) );
  AND2X1 U343 ( .A(add_3_root_r119_carry_18_), .B(in_17bit_b[16]), .Y(
        add_1_root_r119_A_19_) );
  XOR2X1 U344 ( .A(in_17bit_b[16]), .B(add_3_root_r119_carry_18_), .Y(
        add_1_root_r119_A_18_) );
  AND2X1 U345 ( .A(in_17bit_b[1]), .B(in_17bit_b[0]), .Y(
        add_3_root_r119_carry_3_) );
  AND2X1 U346 ( .A(add_2_root_r115_carry_19_), .B(in_17bit_b[16]), .Y(
        add_2_root_r115_SUM_20_) );
  XOR2X1 U347 ( .A(in_17bit_b[16]), .B(add_2_root_r115_carry_19_), .Y(
        add_2_root_r115_SUM_19_) );
  AND2X1 U348 ( .A(add_2_root_r115_carry_18_), .B(in_17bit_b[15]), .Y(
        add_2_root_r115_carry_19_) );
  XOR2X1 U349 ( .A(in_17bit_b[15]), .B(add_2_root_r115_carry_18_), .Y(
        add_2_root_r115_SUM_18_) );
  XOR2X1 U350 ( .A(in_17bit_b[0]), .B(in_17bit_b[2]), .Y(
        add_2_root_r115_SUM_3_) );
  AND2X1 U351 ( .A(add_1_root_r115_carry_22_), .B(in_17bit_b[16]), .Y(
        add_1_root_r115_SUM_23_) );
  XOR2X1 U352 ( .A(in_17bit_b[16]), .B(add_1_root_r115_carry_22_), .Y(
        add_1_root_r115_SUM_22_) );
  AND2X1 U353 ( .A(add_1_root_r115_carry_21_), .B(in_17bit_b[15]), .Y(
        add_1_root_r115_carry_22_) );
  XOR2X1 U354 ( .A(in_17bit_b[15]), .B(add_1_root_r115_carry_21_), .Y(
        add_1_root_r115_SUM_21_) );
  AND2X1 U355 ( .A(in_17bit_b[2]), .B(in_17bit_b[0]), .Y(
        add_1_root_r115_carry_7_) );
  XOR2X1 U356 ( .A(n15), .B(sub_add_54_b0_carry[16]), .Y(N29) );
  AND2X1 U357 ( .A(sub_add_54_b0_carry[15]), .B(n201), .Y(
        sub_add_54_b0_carry[16]) );
  XOR2X1 U358 ( .A(n201), .B(sub_add_54_b0_carry[15]), .Y(N28) );
  AND2X1 U359 ( .A(sub_add_54_b0_carry[14]), .B(n200), .Y(
        sub_add_54_b0_carry[15]) );
  XOR2X1 U360 ( .A(n200), .B(sub_add_54_b0_carry[14]), .Y(N27) );
  AND2X1 U361 ( .A(sub_add_54_b0_carry[13]), .B(n199), .Y(
        sub_add_54_b0_carry[14]) );
  XOR2X1 U362 ( .A(n199), .B(sub_add_54_b0_carry[13]), .Y(N26) );
  AND2X1 U363 ( .A(sub_add_54_b0_carry[12]), .B(n198), .Y(
        sub_add_54_b0_carry[13]) );
  XOR2X1 U364 ( .A(n198), .B(sub_add_54_b0_carry[12]), .Y(N25) );
  AND2X1 U365 ( .A(sub_add_54_b0_carry[11]), .B(n197), .Y(
        sub_add_54_b0_carry[12]) );
  XOR2X1 U366 ( .A(n197), .B(sub_add_54_b0_carry[11]), .Y(N24) );
  AND2X1 U367 ( .A(sub_add_54_b0_carry[10]), .B(n196), .Y(
        sub_add_54_b0_carry[11]) );
  XOR2X1 U368 ( .A(n196), .B(sub_add_54_b0_carry[10]), .Y(N23) );
  AND2X1 U369 ( .A(sub_add_54_b0_carry[9]), .B(n195), .Y(
        sub_add_54_b0_carry[10]) );
  XOR2X1 U370 ( .A(n195), .B(sub_add_54_b0_carry[9]), .Y(N22) );
  AND2X1 U371 ( .A(sub_add_54_b0_carry[8]), .B(n194), .Y(
        sub_add_54_b0_carry[9]) );
  XOR2X1 U372 ( .A(n194), .B(sub_add_54_b0_carry[8]), .Y(N21) );
  AND2X1 U373 ( .A(sub_add_54_b0_carry[7]), .B(n193), .Y(
        sub_add_54_b0_carry[8]) );
  XOR2X1 U374 ( .A(n193), .B(sub_add_54_b0_carry[7]), .Y(N20) );
  AND2X1 U375 ( .A(sub_add_54_b0_carry[6]), .B(n192), .Y(
        sub_add_54_b0_carry[7]) );
  XOR2X1 U376 ( .A(n192), .B(sub_add_54_b0_carry[6]), .Y(N19) );
  AND2X1 U377 ( .A(sub_add_54_b0_carry[5]), .B(n191), .Y(
        sub_add_54_b0_carry[6]) );
  XOR2X1 U378 ( .A(n191), .B(sub_add_54_b0_carry[5]), .Y(N18) );
  AND2X1 U379 ( .A(sub_add_54_b0_carry[4]), .B(n190), .Y(
        sub_add_54_b0_carry[5]) );
  XOR2X1 U380 ( .A(n190), .B(sub_add_54_b0_carry[4]), .Y(N17) );
  AND2X1 U381 ( .A(sub_add_54_b0_carry[3]), .B(n189), .Y(
        sub_add_54_b0_carry[4]) );
  XOR2X1 U382 ( .A(n189), .B(sub_add_54_b0_carry[3]), .Y(N16) );
  AND2X1 U383 ( .A(sub_add_54_b0_carry[2]), .B(n188), .Y(
        sub_add_54_b0_carry[3]) );
  XOR2X1 U384 ( .A(n188), .B(sub_add_54_b0_carry[2]), .Y(N15) );
  AND2X1 U385 ( .A(n186), .B(n187), .Y(sub_add_54_b0_carry[2]) );
  XOR2X1 U386 ( .A(n187), .B(n186), .Y(N14) );
  XOR2X1 U387 ( .A(n6), .B(sub_add_75_b0_carry[15]), .Y(N480) );
  AND2X1 U388 ( .A(sub_add_75_b0_carry[14]), .B(n7), .Y(
        sub_add_75_b0_carry[15]) );
  XOR2X1 U389 ( .A(n7), .B(sub_add_75_b0_carry[14]), .Y(N479) );
  AND2X1 U390 ( .A(sub_add_75_b0_carry[13]), .B(n8), .Y(
        sub_add_75_b0_carry[14]) );
  AND2X1 U391 ( .A(n25), .B(n5), .Y(sub_add_75_b0_carry[13]) );
  AND2X1 U392 ( .A(in_17bit_b[0]), .B(in_17bit_b[4]), .Y(
        add_1_root_r112_carry_5_) );
endmodule


module multi16_11_DW01_add_0 ( A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, 
        A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, 
        A_4_, B_23_, B_22_, B_21_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, 
        B_14_, B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, 
        SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, 
        SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, 
        SUM_7_ );
  input A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_,
         A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, B_23_, B_22_,
         B_21_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_,
         B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_;
  output SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_,
         SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_,
         SUM_8_, SUM_7_;
  wire   n1, n2, n3, n4;
  wire   [23:7] carry;

  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry[7]), .CO(carry[8]), .S(SUM_7_)
         );
  ADDFX2 U1_21 ( .A(A_21_), .B(B_21_), .CI(carry[21]), .CO(carry[22]), .S(
        SUM_21_) );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry[20]), .CO(carry[21]), .S(
        SUM_20_) );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry[19]), .CO(carry[20]), .S(
        SUM_19_) );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry[18]), .CO(carry[19]), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry[17]), .CO(carry[18]), .S(
        SUM_17_) );
  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry[16]), .CO(carry[17]), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry[15]), .CO(carry[16]), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry[14]), .CO(carry[15]), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry[13]), .CO(carry[14]), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry[12]), .CO(carry[13]), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry[11]), .CO(carry[12]), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry[10]), .CO(carry[11]), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry[9]), .CO(carry[10]), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry[8]), .CO(carry[9]), .S(SUM_8_)
         );
  ADDFX2 U1_22 ( .A(A_22_), .B(B_22_), .CI(carry[22]), .CO(carry[23]), .S(
        SUM_22_) );
  AND2X2 U1 ( .A(A_4_), .B(B_4_), .Y(n1) );
  XOR2X1 U2 ( .A(B_23_), .B(carry[23]), .Y(SUM_23_) );
  OAI2BB1X1 U3 ( .A0N(n2), .A1N(A_6_), .B0(n3), .Y(carry[7]) );
  OAI21XL U4 ( .A0(A_6_), .A1(n2), .B0(B_6_), .Y(n3) );
  OAI2BB1X1 U5 ( .A0N(n1), .A1N(A_5_), .B0(n4), .Y(n2) );
  OAI21XL U6 ( .A0(A_5_), .A1(n1), .B0(B_5_), .Y(n4) );
endmodule


module multi16_11_DW01_add_4 ( A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, 
        A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, 
        B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, 
        B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, SUM_22_, SUM_21_, SUM_20_, 
        SUM_19_, SUM_18_, SUM_17_, SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, 
        SUM_11_, SUM_10_, SUM_9_, SUM_8_, SUM_7_ );
  input A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_,
         A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, B_20_, B_19_,
         B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, B_10_, B_9_,
         B_8_, B_7_, B_6_, B_5_;
  output SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_,
         SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_,
         SUM_7_;
  wire   carry_21_, carry_20_, carry_19_, carry_18_, carry_17_, carry_16_,
         carry_15_, carry_14_, carry_13_, carry_12_, carry_11_, carry_10_,
         carry_9_, carry_8_, carry_7_, n1;

  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry_16_), .CO(carry_17_), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry_15_), .CO(carry_16_), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry_14_), .CO(carry_15_), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry_13_), .CO(carry_14_), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry_12_), .CO(carry_13_), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry_11_), .CO(carry_12_), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry_10_), .CO(carry_11_), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry_9_), .CO(carry_10_), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry_8_), .CO(carry_9_), .S(SUM_8_)
         );
  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry_7_), .CO(carry_8_), .S(SUM_7_)
         );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry_20_), .CO(carry_21_), .S(
        SUM_20_) );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry_19_), .CO(carry_20_), .S(
        SUM_19_) );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry_18_), .CO(carry_19_), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry_17_), .CO(carry_18_), .S(
        SUM_17_) );
  ADDFX2 U1_21 ( .A(A_21_), .B(B_21_), .CI(carry_21_), .CO(SUM_22_), .S(
        SUM_21_) );
  OAI2BB1X1 U1 ( .A0N(A_6_), .A1N(B_6_), .B0(n1), .Y(carry_7_) );
  OAI211X1 U2 ( .A0(B_6_), .A1(A_6_), .B0(A_5_), .C0(B_5_), .Y(n1) );
endmodule


module multi16_11_DW01_add_6 ( A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, 
        A_16_, A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, 
        A_6_, A_5_, A_4_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, 
        B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, 
        SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, 
        SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, 
        SUM_7_ );
  input A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_,
         A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, B_20_,
         B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, B_10_,
         B_9_, B_8_, B_7_, B_6_, B_5_, B_4_;
  output SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_,
         SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_,
         SUM_8_, SUM_7_;
  wire   n1, n2, n3, n4, n5, n6;
  wire   [21:7] carry;

  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry[7]), .CO(carry[8]), .S(SUM_7_)
         );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry[18]), .CO(carry[19]), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry[17]), .CO(carry[18]), .S(
        SUM_17_) );
  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry[16]), .CO(carry[17]), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry[15]), .CO(carry[16]), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry[14]), .CO(carry[15]), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry[13]), .CO(carry[14]), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry[12]), .CO(carry[13]), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry[11]), .CO(carry[12]), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry[10]), .CO(carry[11]), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry[9]), .CO(carry[10]), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry[8]), .CO(carry[9]), .S(SUM_8_)
         );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry[19]), .CO(carry[20]), .S(
        SUM_19_) );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry[20]), .CO(carry[21]), .S(
        SUM_20_) );
  AND2X2 U1 ( .A(A_22_), .B(n2), .Y(n1) );
  AND2X2 U2 ( .A(A_21_), .B(carry[21]), .Y(n2) );
  AND2X2 U3 ( .A(A_4_), .B(B_4_), .Y(n3) );
  XOR2X1 U4 ( .A(A_23_), .B(n1), .Y(SUM_23_) );
  XOR2X1 U5 ( .A(A_21_), .B(carry[21]), .Y(SUM_21_) );
  XOR2X1 U6 ( .A(A_22_), .B(n2), .Y(SUM_22_) );
  OAI2BB1X1 U7 ( .A0N(n4), .A1N(A_6_), .B0(n5), .Y(carry[7]) );
  OAI21XL U8 ( .A0(A_6_), .A1(n4), .B0(B_6_), .Y(n5) );
  OAI2BB1X1 U9 ( .A0N(n3), .A1N(A_5_), .B0(n6), .Y(n4) );
  OAI21XL U10 ( .A0(A_5_), .A1(n3), .B0(B_5_), .Y(n6) );
endmodule


module multi16_11 ( in_17bit, in_8bit, out );
  input [16:0] in_17bit;
  input [7:0] in_8bit;
  output [16:0] out;
  wire   n289, n290, n291, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23,
         N24, N25, N26, N27, N28, N29, N108, N109, N110, N111, N112, N113,
         N114, N115, N116, N117, N118, N119, N120, N121, N122, N123, N205,
         N206, N207, N208, N209, N210, N211, N212, N213, N214, N215, N216,
         N217, N218, N219, N220, N221, N347, N348, N349, N350, N351, N352,
         N353, N354, N355, N356, N357, N358, N359, N360, N361, N362, N363,
         N446, N447, N448, N449, N450, N451, N452, N453, N454, N455, N456,
         N457, N458, N459, N460, N461, N462, N463, N479, N480, N481,
         add_2_root_r119_carry_10_, add_2_root_r119_carry_11_,
         add_2_root_r119_carry_12_, add_2_root_r119_carry_13_,
         add_2_root_r119_carry_14_, add_2_root_r119_carry_15_,
         add_2_root_r119_carry_16_, add_2_root_r119_carry_17_,
         add_2_root_r119_carry_18_, add_2_root_r119_carry_19_,
         add_2_root_r119_carry_20_, add_2_root_r119_carry_21_,
         add_2_root_r119_carry_6_, add_2_root_r119_carry_7_,
         add_2_root_r119_carry_8_, add_2_root_r119_carry_9_,
         add_2_root_r119_SUM_6_, add_2_root_r119_SUM_7_,
         add_2_root_r119_SUM_8_, add_2_root_r119_SUM_9_,
         add_2_root_r119_SUM_10_, add_2_root_r119_SUM_11_,
         add_2_root_r119_SUM_12_, add_2_root_r119_SUM_13_,
         add_2_root_r119_SUM_14_, add_2_root_r119_SUM_15_,
         add_2_root_r119_SUM_16_, add_2_root_r119_SUM_17_,
         add_2_root_r119_SUM_18_, add_2_root_r119_SUM_19_,
         add_2_root_r119_SUM_20_, add_2_root_r119_SUM_21_,
         add_2_root_r119_SUM_22_, add_1_root_r119_SUM_6_,
         add_1_root_r119_SUM_7_, add_1_root_r119_SUM_8_,
         add_1_root_r119_SUM_9_, add_1_root_r119_SUM_10_,
         add_1_root_r119_SUM_11_, add_1_root_r119_SUM_12_,
         add_1_root_r119_SUM_13_, add_1_root_r119_SUM_14_,
         add_1_root_r119_SUM_15_, add_1_root_r119_SUM_16_,
         add_1_root_r119_SUM_17_, add_1_root_r119_SUM_18_,
         add_1_root_r119_SUM_19_, add_1_root_r119_SUM_20_,
         add_1_root_r119_SUM_21_, add_1_root_r119_SUM_22_,
         add_1_root_r119_SUM_23_, add_1_root_r119_A_2_, add_1_root_r119_A_3_,
         add_1_root_r119_A_4_, add_1_root_r119_A_5_, add_1_root_r119_A_6_,
         add_1_root_r119_A_7_, add_1_root_r119_A_8_, add_1_root_r119_A_9_,
         add_1_root_r119_A_10_, add_1_root_r119_A_11_, add_1_root_r119_A_12_,
         add_1_root_r119_A_13_, add_1_root_r119_A_14_, add_1_root_r119_A_15_,
         add_1_root_r119_A_16_, add_1_root_r119_A_17_, add_1_root_r119_A_18_,
         add_1_root_r119_A_19_, add_3_root_r119_carry_10_,
         add_3_root_r119_carry_11_, add_3_root_r119_carry_12_,
         add_3_root_r119_carry_13_, add_3_root_r119_carry_14_,
         add_3_root_r119_carry_15_, add_3_root_r119_carry_16_,
         add_3_root_r119_carry_17_, add_3_root_r119_carry_18_,
         add_3_root_r119_carry_4_, add_3_root_r119_carry_5_,
         add_3_root_r119_carry_6_, add_3_root_r119_carry_7_,
         add_3_root_r119_carry_8_, add_3_root_r119_carry_9_,
         add_1_root_r112_carry_10_, add_1_root_r112_carry_11_,
         add_1_root_r112_carry_12_, add_1_root_r112_carry_13_,
         add_1_root_r112_carry_14_, add_1_root_r112_carry_15_,
         add_1_root_r112_carry_16_, add_1_root_r112_carry_17_,
         add_1_root_r112_carry_18_, add_1_root_r112_carry_19_,
         add_1_root_r112_carry_20_, add_1_root_r112_carry_5_,
         add_1_root_r112_carry_6_, add_1_root_r112_carry_7_,
         add_1_root_r112_carry_8_, add_1_root_r112_carry_9_,
         add_1_root_r112_SUM_1_, add_1_root_r112_SUM_2_,
         add_1_root_r112_SUM_3_, add_1_root_r112_SUM_4_,
         add_1_root_r112_SUM_5_, add_1_root_r112_SUM_6_,
         add_1_root_r112_SUM_7_, add_1_root_r112_SUM_8_,
         add_1_root_r112_SUM_9_, add_1_root_r112_SUM_10_,
         add_1_root_r112_SUM_11_, add_1_root_r112_SUM_12_,
         add_1_root_r112_SUM_13_, add_1_root_r112_SUM_14_,
         add_1_root_r112_SUM_15_, add_1_root_r112_SUM_16_,
         add_1_root_r112_SUM_17_, add_1_root_r112_SUM_18_,
         add_1_root_r112_SUM_19_, add_1_root_r112_SUM_20_,
         add_1_root_r112_SUM_21_, add_2_root_r115_carry_10_,
         add_2_root_r115_carry_11_, add_2_root_r115_carry_12_,
         add_2_root_r115_carry_13_, add_2_root_r115_carry_14_,
         add_2_root_r115_carry_15_, add_2_root_r115_carry_16_,
         add_2_root_r115_carry_17_, add_2_root_r115_carry_18_,
         add_2_root_r115_carry_19_, add_2_root_r115_carry_5_,
         add_2_root_r115_carry_6_, add_2_root_r115_carry_7_,
         add_2_root_r115_carry_8_, add_2_root_r115_carry_9_,
         add_2_root_r115_SUM_3_, add_2_root_r115_SUM_4_,
         add_2_root_r115_SUM_5_, add_2_root_r115_SUM_6_,
         add_2_root_r115_SUM_7_, add_2_root_r115_SUM_8_,
         add_2_root_r115_SUM_9_, add_2_root_r115_SUM_10_,
         add_2_root_r115_SUM_11_, add_2_root_r115_SUM_12_,
         add_2_root_r115_SUM_13_, add_2_root_r115_SUM_14_,
         add_2_root_r115_SUM_15_, add_2_root_r115_SUM_16_,
         add_2_root_r115_SUM_17_, add_2_root_r115_SUM_18_,
         add_2_root_r115_SUM_19_, add_2_root_r115_SUM_20_,
         add_1_root_r115_carry_10_, add_1_root_r115_carry_11_,
         add_1_root_r115_carry_12_, add_1_root_r115_carry_13_,
         add_1_root_r115_carry_14_, add_1_root_r115_carry_15_,
         add_1_root_r115_carry_16_, add_1_root_r115_carry_17_,
         add_1_root_r115_carry_18_, add_1_root_r115_carry_19_,
         add_1_root_r115_carry_20_, add_1_root_r115_carry_21_,
         add_1_root_r115_carry_22_, add_1_root_r115_carry_7_,
         add_1_root_r115_carry_8_, add_1_root_r115_carry_9_,
         add_1_root_r115_SUM_7_, add_1_root_r115_SUM_8_,
         add_1_root_r115_SUM_9_, add_1_root_r115_SUM_10_,
         add_1_root_r115_SUM_11_, add_1_root_r115_SUM_12_,
         add_1_root_r115_SUM_13_, add_1_root_r115_SUM_14_,
         add_1_root_r115_SUM_15_, add_1_root_r115_SUM_16_,
         add_1_root_r115_SUM_17_, add_1_root_r115_SUM_18_,
         add_1_root_r115_SUM_19_, add_1_root_r115_SUM_20_,
         add_1_root_r115_SUM_21_, add_1_root_r115_SUM_22_,
         add_1_root_r115_SUM_23_, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n20, n21, n22, n23, n24, n25, n26, n28,
         n29, n30, n31, n32, n33, n34, n35, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n158, n160, n163, n164, n168, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288;
  wire   [16:0] in_17bit_b;
  wire   [23:8] neg_mul;
  wire   [16:13] sub_add_75_b0_carry;
  wire   [16:2] sub_add_54_b0_carry;
  wire   [22:7] add_1_root_r119_carry;

  multi16_11_DW01_add_0 add_0_root_r119 ( .A_22_(add_2_root_r119_SUM_22_), 
        .A_21_(add_2_root_r119_SUM_21_), .A_20_(add_2_root_r119_SUM_20_), 
        .A_19_(add_2_root_r119_SUM_19_), .A_18_(add_2_root_r119_SUM_18_), 
        .A_17_(add_2_root_r119_SUM_17_), .A_16_(add_2_root_r119_SUM_16_), 
        .A_15_(add_2_root_r119_SUM_15_), .A_14_(add_2_root_r119_SUM_14_), 
        .A_13_(add_2_root_r119_SUM_13_), .A_12_(add_2_root_r119_SUM_12_), 
        .A_11_(add_2_root_r119_SUM_11_), .A_10_(add_2_root_r119_SUM_10_), 
        .A_9_(add_2_root_r119_SUM_9_), .A_8_(add_2_root_r119_SUM_8_), .A_7_(
        add_2_root_r119_SUM_7_), .A_6_(add_2_root_r119_SUM_6_), .A_5_(
        add_1_root_r119_A_2_), .A_4_(in_17bit_b[0]), .B_23_(
        add_1_root_r119_SUM_23_), .B_22_(add_1_root_r119_SUM_22_), .B_21_(
        add_1_root_r119_SUM_21_), .B_20_(add_1_root_r119_SUM_20_), .B_19_(
        add_1_root_r119_SUM_19_), .B_18_(add_1_root_r119_SUM_18_), .B_17_(
        add_1_root_r119_SUM_17_), .B_16_(add_1_root_r119_SUM_16_), .B_15_(
        add_1_root_r119_SUM_15_), .B_14_(add_1_root_r119_SUM_14_), .B_13_(
        add_1_root_r119_SUM_13_), .B_12_(add_1_root_r119_SUM_12_), .B_11_(
        add_1_root_r119_SUM_11_), .B_10_(add_1_root_r119_SUM_10_), .B_9_(
        add_1_root_r119_SUM_9_), .B_8_(add_1_root_r119_SUM_8_), .B_7_(
        add_1_root_r119_SUM_7_), .B_6_(add_1_root_r119_SUM_6_), .B_5_(
        add_1_root_r119_A_5_), .B_4_(add_1_root_r119_A_4_), .SUM_23_(N363), 
        .SUM_22_(N362), .SUM_21_(N361), .SUM_20_(N360), .SUM_19_(N359), 
        .SUM_18_(N358), .SUM_17_(N357), .SUM_16_(N356), .SUM_15_(N355), 
        .SUM_14_(N354), .SUM_13_(N353), .SUM_12_(N352), .SUM_11_(N351), 
        .SUM_10_(N350), .SUM_9_(N349), .SUM_8_(N348), .SUM_7_(N347) );
  multi16_11_DW01_add_4 add_0_root_r112 ( .A_21_(in_17bit_b[16]), .A_20_(
        in_17bit_b[15]), .A_19_(in_17bit_b[14]), .A_18_(in_17bit_b[13]), 
        .A_17_(in_17bit_b[12]), .A_16_(in_17bit_b[11]), .A_15_(in_17bit_b[10]), 
        .A_14_(in_17bit_b[9]), .A_13_(in_17bit_b[8]), .A_12_(in_17bit_b[7]), 
        .A_11_(in_17bit_b[6]), .A_10_(in_17bit_b[5]), .A_9_(in_17bit_b[4]), 
        .A_8_(in_17bit_b[3]), .A_7_(in_17bit_b[2]), .A_6_(n205), .A_5_(
        in_17bit_b[0]), .B_21_(add_1_root_r112_SUM_21_), .B_20_(
        add_1_root_r112_SUM_20_), .B_19_(add_1_root_r112_SUM_19_), .B_18_(
        add_1_root_r112_SUM_18_), .B_17_(add_1_root_r112_SUM_17_), .B_16_(
        add_1_root_r112_SUM_16_), .B_15_(add_1_root_r112_SUM_15_), .B_14_(
        add_1_root_r112_SUM_14_), .B_13_(add_1_root_r112_SUM_13_), .B_12_(
        add_1_root_r112_SUM_12_), .B_11_(add_1_root_r112_SUM_11_), .B_10_(
        add_1_root_r112_SUM_10_), .B_9_(add_1_root_r112_SUM_9_), .B_8_(
        add_1_root_r112_SUM_8_), .B_7_(add_1_root_r112_SUM_7_), .B_6_(
        add_1_root_r112_SUM_6_), .B_5_(add_1_root_r112_SUM_5_), .SUM_22_(N123), 
        .SUM_21_(N122), .SUM_20_(N121), .SUM_19_(N120), .SUM_18_(N119), 
        .SUM_17_(N118), .SUM_16_(N117), .SUM_15_(N116), .SUM_14_(N115), 
        .SUM_13_(N114), .SUM_12_(N113), .SUM_11_(N112), .SUM_10_(N111), 
        .SUM_9_(N110), .SUM_8_(N109), .SUM_7_(N108) );
  multi16_11_DW01_add_6 add_0_root_r115 ( .A_23_(add_1_root_r115_SUM_23_), 
        .A_22_(add_1_root_r115_SUM_22_), .A_21_(add_1_root_r115_SUM_21_), 
        .A_20_(add_1_root_r115_SUM_20_), .A_19_(add_1_root_r115_SUM_19_), 
        .A_18_(add_1_root_r115_SUM_18_), .A_17_(add_1_root_r115_SUM_17_), 
        .A_16_(add_1_root_r115_SUM_16_), .A_15_(add_1_root_r115_SUM_15_), 
        .A_14_(add_1_root_r115_SUM_14_), .A_13_(add_1_root_r115_SUM_13_), 
        .A_12_(add_1_root_r115_SUM_12_), .A_11_(add_1_root_r115_SUM_11_), 
        .A_10_(add_1_root_r115_SUM_10_), .A_9_(add_1_root_r115_SUM_9_), .A_8_(
        add_1_root_r115_SUM_8_), .A_7_(add_1_root_r115_SUM_7_), .A_6_(
        add_2_root_r115_SUM_3_), .A_5_(n205), .A_4_(in_17bit_b[0]), .B_20_(
        add_2_root_r115_SUM_20_), .B_19_(add_2_root_r115_SUM_19_), .B_18_(
        add_2_root_r115_SUM_18_), .B_17_(add_2_root_r115_SUM_17_), .B_16_(
        add_2_root_r115_SUM_16_), .B_15_(add_2_root_r115_SUM_15_), .B_14_(
        add_2_root_r115_SUM_14_), .B_13_(add_2_root_r115_SUM_13_), .B_12_(
        add_2_root_r115_SUM_12_), .B_11_(add_2_root_r115_SUM_11_), .B_10_(
        add_2_root_r115_SUM_10_), .B_9_(add_2_root_r115_SUM_9_), .B_8_(
        add_2_root_r115_SUM_8_), .B_7_(add_2_root_r115_SUM_7_), .B_6_(
        add_2_root_r115_SUM_6_), .B_5_(add_2_root_r115_SUM_5_), .B_4_(
        add_2_root_r115_SUM_4_), .SUM_23_(N221), .SUM_22_(N220), .SUM_21_(N219), .SUM_20_(N218), .SUM_19_(N217), .SUM_18_(N216), .SUM_17_(N215), .SUM_16_(
        N214), .SUM_15_(N213), .SUM_14_(N212), .SUM_13_(N211), .SUM_12_(N210), 
        .SUM_11_(N209), .SUM_10_(N208), .SUM_9_(N207), .SUM_8_(N206), .SUM_7_(
        N205) );
  TLATX1 neg_mul_reg_19_ ( .G(N446), .D(N459), .QN(n4) );
  TLATX1 neg_mul_reg_18_ ( .G(N446), .D(N458), .QN(n2) );
  TLATX1 neg_mul_reg_17_ ( .G(N446), .D(N457), .Q(neg_mul[17]), .QN(n1) );
  TLATX1 neg_mul_reg_16_ ( .G(N446), .D(N456), .QN(n3) );
  TLATX1 neg_mul_reg_23_ ( .G(N446), .D(N463), .Q(neg_mul[23]), .QN(n17) );
  TLATX1 neg_mul_reg_22_ ( .G(N446), .D(N462), .Q(neg_mul[22]), .QN(n10) );
  TLATX1 neg_mul_reg_21_ ( .G(N446), .D(N461), .Q(neg_mul[21]), .QN(n9) );
  TLATX1 neg_mul_reg_20_ ( .G(N446), .D(N460), .QN(n15) );
  TLATX1 neg_mul_reg_11_ ( .G(N446), .D(N451), .Q(neg_mul[11]), .QN(n11) );
  TLATX1 neg_mul_reg_12_ ( .G(N446), .D(N452), .Q(neg_mul[12]), .QN(n12) );
  TLATX1 neg_mul_reg_9_ ( .G(N446), .D(N449), .Q(neg_mul[9]), .QN(n5) );
  TLATX1 neg_mul_reg_15_ ( .G(N446), .D(N455), .Q(neg_mul[15]), .QN(n13) );
  TLATX1 neg_mul_reg_14_ ( .G(N446), .D(N454), .Q(neg_mul[14]), .QN(n7) );
  TLATX1 neg_mul_reg_13_ ( .G(N446), .D(N453), .Q(neg_mul[13]), .QN(n8) );
  TLATX1 neg_mul_reg_10_ ( .G(N446), .D(N450), .Q(neg_mul[10]), .QN(n6) );
  TLATX1 neg_mul_reg_8_ ( .G(N446), .D(N448), .Q(neg_mul[8]), .QN(n16) );
  TLATX1 neg_mul_reg_7_ ( .G(N446), .D(N447), .Q(out[0]) );
  BUFX16 U2 ( .A(n20), .Y(n37) );
  BUFX16 U3 ( .A(n24), .Y(n22) );
  CLKINVX3 U4 ( .A(n288), .Y(in_17bit_b[16]) );
  CLKINVX8 U5 ( .A(n47), .Y(n46) );
  BUFX20 U6 ( .A(n24), .Y(n21) );
  NOR2X1 U7 ( .A(n82), .B(n20), .Y(n84) );
  INVX8 U8 ( .A(n47), .Y(n20) );
  INVX8 U9 ( .A(in_17bit[16]), .Y(n47) );
  OAI21X1 U10 ( .A0(n23), .A1(n65), .B0(n64), .Y(n69) );
  NAND2X2 U11 ( .A(n23), .B(n6), .Y(n64) );
  MX2X2 U12 ( .A(neg_mul[21]), .B(N479), .S0(n177), .Y(out[14]) );
  MXI2X2 U13 ( .A(n15), .B(n34), .S0(n177), .Y(out[13]) );
  INVX8 U14 ( .A(n176), .Y(n177) );
  BUFX8 U15 ( .A(n290), .Y(out[5]) );
  AOI2BB2X2 U16 ( .B0(n52), .B1(n23), .A0N(n22), .A1N(neg_mul[8]), .Y(n53) );
  AOI2BB2X1 U17 ( .B0(n89), .B1(n21), .A0N(n21), .A1N(neg_mul[13]), .Y(n90) );
  AOI2BB2X2 U18 ( .B0(n58), .B1(n23), .A0N(n22), .A1N(neg_mul[9]), .Y(n59) );
  NAND4BXL U19 ( .AN(n22), .B(in_8bit[4]), .C(n40), .D(in_8bit[6]), .Y(n186)
         );
  INVX1 U20 ( .A(n186), .Y(n182) );
  BUFX12 U21 ( .A(n24), .Y(n23) );
  AND4X1 U22 ( .A(n40), .B(n22), .C(n226), .D(n41), .Y(n14) );
  AOI22X1 U23 ( .A0(N27), .A1(n25), .B0(in_17bit[14]), .B1(n49), .Y(n277) );
  NOR2X1 U24 ( .A(n20), .B(n74), .Y(n76) );
  CLKBUFX8 U25 ( .A(n291), .Y(out[4]) );
  NAND2X1 U26 ( .A(n21), .B(n7), .Y(n95) );
  BUFX16 U27 ( .A(in_8bit[7]), .Y(n24) );
  NOR2XL U28 ( .A(n20), .B(n168), .Y(n170) );
  NOR2X2 U29 ( .A(n46), .B(n59), .Y(n61) );
  OAI21X2 U30 ( .A0(n46), .A1(n67), .B0(n70), .Y(n68) );
  OR4XL U31 ( .A(in_8bit[4]), .B(in_8bit[5]), .C(in_8bit[6]), .D(n22), .Y(n231) );
  AOI211X2 U32 ( .A0(n37), .A1(n77), .B0(n76), .C0(n75), .Y(n291) );
  AOI211X2 U33 ( .A0(n85), .A1(n37), .B0(n84), .C0(n83), .Y(n290) );
  XOR2X4 U34 ( .A(n173), .B(neg_mul[17]), .Y(out[10]) );
  NOR2X1 U35 ( .A(n20), .B(n98), .Y(n100) );
  AOI2BB2X2 U36 ( .B0(n97), .B1(n23), .A0N(n23), .A1N(neg_mul[14]), .Y(n98) );
  OAI21X2 U37 ( .A0(n21), .A1(n51), .B0(n50), .Y(n55) );
  AOI2BB2X4 U38 ( .B0(n66), .B1(n23), .A0N(n23), .A1N(neg_mul[10]), .Y(n67) );
  NOR2X4 U39 ( .A(n46), .B(n53), .Y(n54) );
  XNOR2X2 U40 ( .A(n20), .B(n21), .Y(n176) );
  NOR2X2 U41 ( .A(n176), .B(n33), .Y(n175) );
  AOI211X2 U42 ( .A0(n20), .A1(n55), .B0(n54), .C0(n35), .Y(out[1]) );
  INVX1 U43 ( .A(n48), .Y(n25) );
  INVXL U44 ( .A(n37), .Y(n48) );
  OAI21X1 U45 ( .A0(n22), .A1(n57), .B0(n56), .Y(n62) );
  NAND2X2 U46 ( .A(n21), .B(n5), .Y(n56) );
  NAND2X2 U47 ( .A(n21), .B(n16), .Y(n50) );
  NOR2X4 U48 ( .A(n29), .B(n174), .Y(n172) );
  AOI211X2 U49 ( .A0(n20), .A1(n62), .B0(n61), .C0(n60), .Y(out[2]) );
  NOR2X4 U50 ( .A(n32), .B(n174), .Y(n28) );
  XNOR2X4 U51 ( .A(n46), .B(n21), .Y(n174) );
  AOI21X4 U52 ( .A0(n37), .A1(n69), .B0(n68), .Y(out[3]) );
  AOI2BB2X1 U53 ( .B0(n81), .B1(n23), .A0N(n21), .A1N(neg_mul[12]), .Y(n82) );
  INVX4 U54 ( .A(n289), .Y(n26) );
  CLKINVX8 U55 ( .A(n26), .Y(out[7]) );
  INVX1 U56 ( .A(n277), .Y(in_17bit_b[14]) );
  INVX1 U57 ( .A(n274), .Y(in_17bit_b[13]) );
  INVX1 U58 ( .A(n241), .Y(in_17bit_b[2]) );
  INVX1 U59 ( .A(n250), .Y(in_17bit_b[5]) );
  INVX1 U60 ( .A(n253), .Y(in_17bit_b[6]) );
  INVX1 U61 ( .A(n256), .Y(in_17bit_b[7]) );
  INVX1 U62 ( .A(n259), .Y(in_17bit_b[8]) );
  INVX1 U63 ( .A(n262), .Y(in_17bit_b[9]) );
  INVX1 U64 ( .A(n265), .Y(in_17bit_b[10]) );
  INVX1 U65 ( .A(n268), .Y(in_17bit_b[11]) );
  INVX1 U66 ( .A(n271), .Y(in_17bit_b[12]) );
  INVX1 U67 ( .A(n247), .Y(in_17bit_b[4]) );
  INVX1 U68 ( .A(n244), .Y(in_17bit_b[3]) );
  XNOR2X4 U69 ( .A(n28), .B(n2), .Y(out[11]) );
  INVX1 U70 ( .A(n45), .Y(n44) );
  NOR3X1 U71 ( .A(n45), .B(n43), .C(n41), .Y(n233) );
  NOR4BX1 U72 ( .AN(n229), .B(n41), .C(n40), .D(n44), .Y(n232) );
  NOR2X1 U73 ( .A(in_8bit[6]), .B(in_8bit[3]), .Y(n229) );
  NAND3X1 U74 ( .A(n44), .B(n43), .C(in_8bit[5]), .Y(n227) );
  ADDFX2 U75 ( .A(in_17bit_b[16]), .B(in_17bit_b[12]), .CI(
        add_1_root_r112_carry_16_), .CO(add_1_root_r112_carry_17_), .S(
        add_1_root_r112_SUM_16_) );
  ADDFX2 U76 ( .A(add_1_root_r119_A_19_), .B(in_17bit_b[13]), .CI(
        add_1_root_r119_carry[19]), .CO(add_1_root_r119_carry[20]), .S(
        add_1_root_r119_SUM_19_) );
  ADDFX2 U77 ( .A(in_17bit_b[16]), .B(in_17bit_b[15]), .CI(
        add_3_root_r119_carry_17_), .CO(add_3_root_r119_carry_18_), .S(
        add_1_root_r119_A_17_) );
  ADDFX2 U78 ( .A(in_17bit_b[16]), .B(in_17bit_b[14]), .CI(
        add_2_root_r115_carry_17_), .CO(add_2_root_r115_carry_18_), .S(
        add_2_root_r115_SUM_17_) );
  ADDFX2 U79 ( .A(in_17bit_b[16]), .B(in_17bit_b[14]), .CI(
        add_1_root_r115_carry_20_), .CO(add_1_root_r115_carry_21_), .S(
        add_1_root_r115_SUM_20_) );
  ADDFX2 U80 ( .A(in_17bit_b[16]), .B(in_17bit_b[15]), .CI(
        add_2_root_r119_carry_20_), .CO(add_2_root_r119_carry_21_), .S(
        add_2_root_r119_SUM_20_) );
  ADDFX2 U81 ( .A(in_17bit_b[3]), .B(n205), .CI(add_1_root_r115_carry_7_), 
        .CO(add_2_root_r115_carry_5_), .S(add_2_root_r115_SUM_4_) );
  ADDFX2 U82 ( .A(in_17bit_b[4]), .B(in_17bit_b[2]), .CI(
        add_2_root_r115_carry_5_), .CO(add_2_root_r115_carry_6_), .S(
        add_2_root_r115_SUM_5_) );
  ADDFX2 U83 ( .A(in_17bit_b[5]), .B(n205), .CI(add_1_root_r112_carry_5_), 
        .CO(add_1_root_r112_carry_6_), .S(add_1_root_r112_SUM_5_) );
  ADDFX2 U84 ( .A(in_17bit_b[6]), .B(in_17bit_b[5]), .CI(
        add_3_root_r119_carry_7_), .CO(add_3_root_r119_carry_8_), .S(
        add_1_root_r119_A_7_) );
  ADDFX2 U85 ( .A(in_17bit_b[6]), .B(in_17bit_b[2]), .CI(
        add_1_root_r112_carry_6_), .CO(add_1_root_r112_carry_7_), .S(
        add_1_root_r112_SUM_6_) );
  ADDFX2 U86 ( .A(in_17bit_b[3]), .B(n205), .CI(add_1_root_r115_carry_7_), 
        .CO(add_1_root_r115_carry_8_), .S(add_1_root_r115_SUM_7_) );
  ADDFX2 U87 ( .A(in_17bit_b[7]), .B(in_17bit_b[6]), .CI(
        add_3_root_r119_carry_8_), .CO(add_3_root_r119_carry_9_), .S(
        add_1_root_r119_A_8_) );
  ADDFX2 U88 ( .A(add_1_root_r119_A_7_), .B(n205), .CI(
        add_1_root_r119_carry[7]), .CO(add_1_root_r119_carry[8]), .S(
        add_1_root_r119_SUM_7_) );
  ADDFX2 U89 ( .A(in_17bit_b[2]), .B(n205), .CI(add_2_root_r119_carry_6_), 
        .CO(add_2_root_r119_carry_7_), .S(add_2_root_r119_SUM_6_) );
  ADDFX2 U90 ( .A(in_17bit_b[4]), .B(in_17bit_b[2]), .CI(
        add_1_root_r115_carry_8_), .CO(add_1_root_r115_carry_9_), .S(
        add_1_root_r115_SUM_8_) );
  ADDFX2 U91 ( .A(in_17bit_b[8]), .B(in_17bit_b[7]), .CI(
        add_3_root_r119_carry_9_), .CO(add_3_root_r119_carry_10_), .S(
        add_1_root_r119_A_9_) );
  ADDFX2 U92 ( .A(add_1_root_r119_A_8_), .B(in_17bit_b[2]), .CI(
        add_1_root_r119_carry[8]), .CO(add_1_root_r119_carry[9]), .S(
        add_1_root_r119_SUM_8_) );
  ADDFX2 U93 ( .A(in_17bit_b[3]), .B(in_17bit_b[2]), .CI(
        add_2_root_r119_carry_7_), .CO(add_2_root_r119_carry_8_), .S(
        add_2_root_r119_SUM_7_) );
  ADDFX2 U94 ( .A(in_17bit_b[6]), .B(in_17bit_b[4]), .CI(
        add_2_root_r115_carry_7_), .CO(add_2_root_r115_carry_8_), .S(
        add_2_root_r115_SUM_7_) );
  ADDFX2 U95 ( .A(in_17bit_b[9]), .B(in_17bit_b[8]), .CI(
        add_3_root_r119_carry_10_), .CO(add_3_root_r119_carry_11_), .S(
        add_1_root_r119_A_10_) );
  ADDFX2 U96 ( .A(in_17bit_b[9]), .B(in_17bit_b[5]), .CI(
        add_1_root_r112_carry_9_), .CO(add_1_root_r112_carry_10_), .S(
        add_1_root_r112_SUM_9_) );
  ADDFX2 U97 ( .A(in_17bit_b[6]), .B(in_17bit_b[4]), .CI(
        add_1_root_r115_carry_10_), .CO(add_1_root_r115_carry_11_), .S(
        add_1_root_r115_SUM_10_) );
  ADDFX2 U98 ( .A(add_1_root_r119_A_9_), .B(in_17bit_b[3]), .CI(
        add_1_root_r119_carry[9]), .CO(add_1_root_r119_carry[10]), .S(
        add_1_root_r119_SUM_9_) );
  ADDFX2 U99 ( .A(in_17bit_b[7]), .B(in_17bit_b[5]), .CI(
        add_2_root_r115_carry_8_), .CO(add_2_root_r115_carry_9_), .S(
        add_2_root_r115_SUM_8_) );
  ADDFX2 U100 ( .A(in_17bit_b[10]), .B(in_17bit_b[9]), .CI(
        add_3_root_r119_carry_11_), .CO(add_3_root_r119_carry_12_), .S(
        add_1_root_r119_A_11_) );
  ADDFX2 U101 ( .A(in_17bit_b[5]), .B(in_17bit_b[4]), .CI(
        add_2_root_r119_carry_9_), .CO(add_2_root_r119_carry_10_), .S(
        add_2_root_r119_SUM_9_) );
  ADDFX2 U102 ( .A(in_17bit_b[8]), .B(in_17bit_b[6]), .CI(
        add_2_root_r115_carry_9_), .CO(add_2_root_r115_carry_10_), .S(
        add_2_root_r115_SUM_9_) );
  ADDFX2 U103 ( .A(in_17bit_b[10]), .B(in_17bit_b[6]), .CI(
        add_1_root_r112_carry_10_), .CO(add_1_root_r112_carry_11_), .S(
        add_1_root_r112_SUM_10_) );
  ADDFX2 U104 ( .A(in_17bit_b[11]), .B(in_17bit_b[10]), .CI(
        add_3_root_r119_carry_12_), .CO(add_3_root_r119_carry_13_), .S(
        add_1_root_r119_A_12_) );
  ADDFX2 U105 ( .A(add_1_root_r119_A_11_), .B(in_17bit_b[5]), .CI(
        add_1_root_r119_carry[11]), .CO(add_1_root_r119_carry[12]), .S(
        add_1_root_r119_SUM_11_) );
  ADDFX2 U106 ( .A(in_17bit_b[6]), .B(in_17bit_b[5]), .CI(
        add_2_root_r119_carry_10_), .CO(add_2_root_r119_carry_11_), .S(
        add_2_root_r119_SUM_10_) );
  ADDFX2 U107 ( .A(in_17bit_b[9]), .B(in_17bit_b[7]), .CI(
        add_2_root_r115_carry_10_), .CO(add_2_root_r115_carry_11_), .S(
        add_2_root_r115_SUM_10_) );
  ADDFX2 U108 ( .A(in_17bit_b[11]), .B(in_17bit_b[7]), .CI(
        add_1_root_r112_carry_11_), .CO(add_1_root_r112_carry_12_), .S(
        add_1_root_r112_SUM_11_) );
  ADDFX2 U109 ( .A(in_17bit_b[8]), .B(in_17bit_b[6]), .CI(
        add_1_root_r115_carry_12_), .CO(add_1_root_r115_carry_13_), .S(
        add_1_root_r115_SUM_12_) );
  ADDFX2 U110 ( .A(in_17bit_b[12]), .B(in_17bit_b[11]), .CI(
        add_3_root_r119_carry_13_), .CO(add_3_root_r119_carry_14_), .S(
        add_1_root_r119_A_13_) );
  ADDFX2 U111 ( .A(add_1_root_r119_A_12_), .B(in_17bit_b[6]), .CI(
        add_1_root_r119_carry[12]), .CO(add_1_root_r119_carry[13]), .S(
        add_1_root_r119_SUM_12_) );
  ADDFX2 U112 ( .A(in_17bit_b[7]), .B(in_17bit_b[6]), .CI(
        add_2_root_r119_carry_11_), .CO(add_2_root_r119_carry_12_), .S(
        add_2_root_r119_SUM_11_) );
  ADDFX2 U113 ( .A(in_17bit_b[10]), .B(in_17bit_b[8]), .CI(
        add_2_root_r115_carry_11_), .CO(add_2_root_r115_carry_12_), .S(
        add_2_root_r115_SUM_11_) );
  ADDFX2 U114 ( .A(in_17bit_b[12]), .B(in_17bit_b[8]), .CI(
        add_1_root_r112_carry_12_), .CO(add_1_root_r112_carry_13_), .S(
        add_1_root_r112_SUM_12_) );
  ADDFX2 U115 ( .A(in_17bit_b[9]), .B(in_17bit_b[7]), .CI(
        add_1_root_r115_carry_13_), .CO(add_1_root_r115_carry_14_), .S(
        add_1_root_r115_SUM_13_) );
  ADDFX2 U116 ( .A(in_17bit_b[13]), .B(in_17bit_b[12]), .CI(
        add_3_root_r119_carry_14_), .CO(add_3_root_r119_carry_15_), .S(
        add_1_root_r119_A_14_) );
  ADDFX2 U117 ( .A(add_1_root_r119_A_13_), .B(in_17bit_b[7]), .CI(
        add_1_root_r119_carry[13]), .CO(add_1_root_r119_carry[14]), .S(
        add_1_root_r119_SUM_13_) );
  ADDFX2 U118 ( .A(in_17bit_b[8]), .B(in_17bit_b[7]), .CI(
        add_2_root_r119_carry_12_), .CO(add_2_root_r119_carry_13_), .S(
        add_2_root_r119_SUM_12_) );
  ADDFX2 U119 ( .A(in_17bit_b[11]), .B(in_17bit_b[9]), .CI(
        add_2_root_r115_carry_12_), .CO(add_2_root_r115_carry_13_), .S(
        add_2_root_r115_SUM_12_) );
  ADDFX2 U120 ( .A(in_17bit_b[13]), .B(in_17bit_b[9]), .CI(
        add_1_root_r112_carry_13_), .CO(add_1_root_r112_carry_14_), .S(
        add_1_root_r112_SUM_13_) );
  ADDFX2 U121 ( .A(in_17bit_b[14]), .B(in_17bit_b[13]), .CI(
        add_3_root_r119_carry_15_), .CO(add_3_root_r119_carry_16_), .S(
        add_1_root_r119_A_15_) );
  ADDFX2 U122 ( .A(add_1_root_r119_A_14_), .B(in_17bit_b[8]), .CI(
        add_1_root_r119_carry[14]), .CO(add_1_root_r119_carry[15]), .S(
        add_1_root_r119_SUM_14_) );
  ADDFX2 U123 ( .A(in_17bit_b[3]), .B(in_17bit_b[2]), .CI(
        add_3_root_r119_carry_4_), .CO(add_3_root_r119_carry_5_), .S(
        add_1_root_r119_A_4_) );
  ADDFX2 U124 ( .A(in_17bit_b[2]), .B(n205), .CI(add_2_root_r119_carry_6_), 
        .CO(add_3_root_r119_carry_4_), .S(add_1_root_r119_A_3_) );
  ADDFX2 U125 ( .A(in_17bit_b[9]), .B(in_17bit_b[8]), .CI(
        add_2_root_r119_carry_13_), .CO(add_2_root_r119_carry_14_), .S(
        add_2_root_r119_SUM_13_) );
  ADDFX2 U126 ( .A(in_17bit_b[14]), .B(in_17bit_b[10]), .CI(
        add_1_root_r112_carry_14_), .CO(add_1_root_r112_carry_15_), .S(
        add_1_root_r112_SUM_14_) );
  ADDFX2 U127 ( .A(in_17bit_b[11]), .B(in_17bit_b[9]), .CI(
        add_1_root_r115_carry_15_), .CO(add_1_root_r115_carry_16_), .S(
        add_1_root_r115_SUM_15_) );
  ADDFX2 U128 ( .A(add_1_root_r119_A_15_), .B(in_17bit_b[9]), .CI(
        add_1_root_r119_carry[15]), .CO(add_1_root_r119_carry[16]), .S(
        add_1_root_r119_SUM_15_) );
  ADDFX2 U129 ( .A(in_17bit_b[10]), .B(in_17bit_b[9]), .CI(
        add_2_root_r119_carry_14_), .CO(add_2_root_r119_carry_15_), .S(
        add_2_root_r119_SUM_14_) );
  ADDFX2 U130 ( .A(in_17bit_b[13]), .B(in_17bit_b[11]), .CI(
        add_2_root_r115_carry_14_), .CO(add_2_root_r115_carry_15_), .S(
        add_2_root_r115_SUM_14_) );
  ADDFX2 U131 ( .A(in_17bit_b[15]), .B(in_17bit_b[11]), .CI(
        add_1_root_r112_carry_15_), .CO(add_1_root_r112_carry_16_), .S(
        add_1_root_r112_SUM_15_) );
  ADDFX2 U132 ( .A(in_17bit_b[12]), .B(in_17bit_b[10]), .CI(
        add_1_root_r115_carry_16_), .CO(add_1_root_r115_carry_17_), .S(
        add_1_root_r115_SUM_16_) );
  ADDFX2 U133 ( .A(add_1_root_r119_A_16_), .B(in_17bit_b[10]), .CI(
        add_1_root_r119_carry[16]), .CO(add_1_root_r119_carry[17]), .S(
        add_1_root_r119_SUM_16_) );
  ADDFX2 U134 ( .A(in_17bit_b[11]), .B(in_17bit_b[10]), .CI(
        add_2_root_r119_carry_15_), .CO(add_2_root_r119_carry_16_), .S(
        add_2_root_r119_SUM_15_) );
  ADDFX2 U135 ( .A(in_17bit_b[14]), .B(in_17bit_b[12]), .CI(
        add_2_root_r115_carry_15_), .CO(add_2_root_r115_carry_16_), .S(
        add_2_root_r115_SUM_15_) );
  ADDFX2 U136 ( .A(in_17bit_b[13]), .B(in_17bit_b[11]), .CI(
        add_1_root_r115_carry_17_), .CO(add_1_root_r115_carry_18_), .S(
        add_1_root_r115_SUM_17_) );
  ADDFX2 U137 ( .A(add_1_root_r119_A_17_), .B(in_17bit_b[11]), .CI(
        add_1_root_r119_carry[17]), .CO(add_1_root_r119_carry[18]), .S(
        add_1_root_r119_SUM_17_) );
  ADDFX2 U138 ( .A(in_17bit_b[12]), .B(in_17bit_b[11]), .CI(
        add_2_root_r119_carry_16_), .CO(add_2_root_r119_carry_17_), .S(
        add_2_root_r119_SUM_16_) );
  ADDFX2 U139 ( .A(in_17bit_b[15]), .B(in_17bit_b[13]), .CI(
        add_2_root_r115_carry_16_), .CO(add_2_root_r115_carry_17_), .S(
        add_2_root_r115_SUM_16_) );
  ADDFX2 U140 ( .A(in_17bit_b[14]), .B(in_17bit_b[12]), .CI(
        add_1_root_r115_carry_18_), .CO(add_1_root_r115_carry_19_), .S(
        add_1_root_r115_SUM_18_) );
  ADDFX2 U141 ( .A(add_1_root_r119_A_18_), .B(in_17bit_b[12]), .CI(
        add_1_root_r119_carry[18]), .CO(add_1_root_r119_carry[19]), .S(
        add_1_root_r119_SUM_18_) );
  ADDFX2 U142 ( .A(in_17bit_b[13]), .B(in_17bit_b[12]), .CI(
        add_2_root_r119_carry_17_), .CO(add_2_root_r119_carry_18_), .S(
        add_2_root_r119_SUM_17_) );
  ADDFX2 U143 ( .A(in_17bit_b[15]), .B(in_17bit_b[13]), .CI(
        add_1_root_r115_carry_19_), .CO(add_1_root_r115_carry_20_), .S(
        add_1_root_r115_SUM_19_) );
  ADDFX2 U144 ( .A(in_17bit_b[14]), .B(in_17bit_b[13]), .CI(
        add_2_root_r119_carry_18_), .CO(add_2_root_r119_carry_19_), .S(
        add_2_root_r119_SUM_18_) );
  ADDFX2 U145 ( .A(in_17bit_b[5]), .B(in_17bit_b[3]), .CI(
        add_2_root_r115_carry_6_), .CO(add_2_root_r115_carry_7_), .S(
        add_2_root_r115_SUM_6_) );
  ADDFX2 U146 ( .A(in_17bit_b[7]), .B(in_17bit_b[3]), .CI(
        add_1_root_r112_carry_7_), .CO(add_1_root_r112_carry_8_), .S(
        add_1_root_r112_SUM_7_) );
  ADDFX2 U147 ( .A(in_17bit_b[8]), .B(in_17bit_b[4]), .CI(
        add_1_root_r112_carry_8_), .CO(add_1_root_r112_carry_9_), .S(
        add_1_root_r112_SUM_8_) );
  ADDFX2 U148 ( .A(in_17bit_b[5]), .B(in_17bit_b[3]), .CI(
        add_1_root_r115_carry_9_), .CO(add_1_root_r115_carry_10_), .S(
        add_1_root_r115_SUM_9_) );
  ADDFX2 U149 ( .A(in_17bit_b[4]), .B(in_17bit_b[3]), .CI(
        add_2_root_r119_carry_8_), .CO(add_2_root_r119_carry_9_), .S(
        add_2_root_r119_SUM_8_) );
  ADDFX2 U150 ( .A(add_1_root_r119_A_10_), .B(in_17bit_b[4]), .CI(
        add_1_root_r119_carry[10]), .CO(add_1_root_r119_carry[11]), .S(
        add_1_root_r119_SUM_10_) );
  ADDFX2 U151 ( .A(in_17bit_b[7]), .B(in_17bit_b[5]), .CI(
        add_1_root_r115_carry_11_), .CO(add_1_root_r115_carry_12_), .S(
        add_1_root_r115_SUM_11_) );
  ADDFX2 U152 ( .A(in_17bit_b[10]), .B(in_17bit_b[8]), .CI(
        add_1_root_r115_carry_14_), .CO(add_1_root_r115_carry_15_), .S(
        add_1_root_r115_SUM_14_) );
  ADDFX2 U153 ( .A(in_17bit_b[12]), .B(in_17bit_b[10]), .CI(
        add_2_root_r115_carry_13_), .CO(add_2_root_r115_carry_14_), .S(
        add_2_root_r115_SUM_13_) );
  ADDFX2 U154 ( .A(in_17bit_b[15]), .B(in_17bit_b[14]), .CI(
        add_3_root_r119_carry_16_), .CO(add_3_root_r119_carry_17_), .S(
        add_1_root_r119_A_16_) );
  ADDFX2 U155 ( .A(in_17bit_b[5]), .B(in_17bit_b[4]), .CI(
        add_3_root_r119_carry_6_), .CO(add_3_root_r119_carry_7_), .S(
        add_1_root_r119_A_6_) );
  ADDFX2 U156 ( .A(in_17bit_b[4]), .B(in_17bit_b[3]), .CI(
        add_3_root_r119_carry_5_), .CO(add_3_root_r119_carry_6_), .S(
        add_1_root_r119_A_5_) );
  ADDFX2 U157 ( .A(in_17bit_b[15]), .B(in_17bit_b[14]), .CI(
        add_2_root_r119_carry_19_), .CO(add_2_root_r119_carry_20_), .S(
        add_2_root_r119_SUM_19_) );
  INVX1 U158 ( .A(n228), .Y(n185) );
  NAND3BX1 U159 ( .AN(in_8bit[5]), .B(n45), .C(in_8bit[3]), .Y(n228) );
  INVX1 U160 ( .A(n25), .Y(n49) );
  INVX1 U161 ( .A(in_8bit[6]), .Y(n42) );
  CLKINVX3 U162 ( .A(n235), .Y(in_17bit_b[0]) );
  INVX1 U163 ( .A(n206), .Y(n287) );
  NAND2XL U164 ( .A(N29), .B(n25), .Y(n288) );
  OAI21XL U165 ( .A0(n287), .A1(n288), .B0(n286), .Y(N463) );
  AOI22X1 U166 ( .A0(N221), .A1(n39), .B0(N363), .B1(n38), .Y(n286) );
  INVX1 U167 ( .A(n158), .Y(n99) );
  CLKINVX3 U168 ( .A(n280), .Y(in_17bit_b[15]) );
  INVX1 U169 ( .A(n94), .Y(n91) );
  INVX1 U170 ( .A(n78), .Y(n75) );
  INVX1 U171 ( .A(n86), .Y(n83) );
  NAND2X1 U172 ( .A(n237), .B(n236), .Y(N447) );
  AOI22X1 U173 ( .A0(N108), .A1(n281), .B0(N205), .B1(n39), .Y(n236) );
  AOI22X1 U174 ( .A0(N347), .A1(n38), .B0(n206), .B1(in_17bit_b[0]), .Y(n237)
         );
  NAND2X1 U175 ( .A(n240), .B(n239), .Y(N448) );
  AOI22X1 U176 ( .A0(N109), .A1(n281), .B0(N206), .B1(n39), .Y(n239) );
  AOI22X1 U177 ( .A0(N348), .A1(n38), .B0(n206), .B1(n205), .Y(n240) );
  INVX1 U178 ( .A(n238), .Y(n205) );
  NAND2X1 U179 ( .A(n243), .B(n242), .Y(N449) );
  AOI22X1 U180 ( .A0(N110), .A1(n281), .B0(N207), .B1(n39), .Y(n242) );
  AOI22X1 U181 ( .A0(N349), .A1(n38), .B0(n206), .B1(in_17bit_b[2]), .Y(n243)
         );
  NAND2X1 U182 ( .A(n246), .B(n245), .Y(N450) );
  AOI22X1 U183 ( .A0(N111), .A1(n281), .B0(N208), .B1(n39), .Y(n245) );
  AOI22X1 U184 ( .A0(N350), .A1(n38), .B0(n206), .B1(in_17bit_b[3]), .Y(n246)
         );
  NAND2X1 U185 ( .A(n249), .B(n248), .Y(N451) );
  AOI22X1 U186 ( .A0(N112), .A1(n281), .B0(N209), .B1(n39), .Y(n248) );
  AOI22X1 U187 ( .A0(N351), .A1(n38), .B0(n206), .B1(in_17bit_b[4]), .Y(n249)
         );
  NAND2X1 U188 ( .A(n252), .B(n251), .Y(N452) );
  AOI22X1 U189 ( .A0(N113), .A1(n281), .B0(N210), .B1(n39), .Y(n251) );
  AOI22X1 U190 ( .A0(N352), .A1(n38), .B0(n206), .B1(in_17bit_b[5]), .Y(n252)
         );
  NAND2X1 U191 ( .A(n255), .B(n254), .Y(N453) );
  AOI22X1 U192 ( .A0(N114), .A1(n281), .B0(N211), .B1(n39), .Y(n254) );
  AOI22X1 U193 ( .A0(N353), .A1(n38), .B0(n206), .B1(in_17bit_b[6]), .Y(n255)
         );
  NAND2X1 U194 ( .A(n258), .B(n257), .Y(N454) );
  AOI22X1 U195 ( .A0(N115), .A1(n281), .B0(N212), .B1(n39), .Y(n257) );
  AOI22X1 U196 ( .A0(N354), .A1(n38), .B0(n206), .B1(in_17bit_b[7]), .Y(n258)
         );
  NAND2X1 U197 ( .A(n261), .B(n260), .Y(N455) );
  AOI22X1 U198 ( .A0(N116), .A1(n281), .B0(N213), .B1(n39), .Y(n260) );
  AOI22X1 U199 ( .A0(N355), .A1(n38), .B0(n206), .B1(in_17bit_b[8]), .Y(n261)
         );
  NAND2X1 U200 ( .A(n264), .B(n263), .Y(N456) );
  AOI22X1 U201 ( .A0(N117), .A1(n281), .B0(N214), .B1(n39), .Y(n263) );
  AOI22X1 U202 ( .A0(N356), .A1(n38), .B0(n206), .B1(in_17bit_b[9]), .Y(n264)
         );
  NAND2X1 U203 ( .A(n267), .B(n266), .Y(N457) );
  AOI22X1 U204 ( .A0(N118), .A1(n281), .B0(N215), .B1(n39), .Y(n266) );
  AOI22X1 U205 ( .A0(N357), .A1(n38), .B0(n206), .B1(in_17bit_b[10]), .Y(n267)
         );
  NAND2X1 U206 ( .A(n270), .B(n269), .Y(N458) );
  AOI22X1 U207 ( .A0(N119), .A1(n281), .B0(N216), .B1(n39), .Y(n269) );
  AOI22X1 U208 ( .A0(N358), .A1(n38), .B0(n206), .B1(in_17bit_b[11]), .Y(n270)
         );
  NAND2X1 U209 ( .A(n273), .B(n272), .Y(N459) );
  AOI22X1 U210 ( .A0(N120), .A1(n281), .B0(N217), .B1(n39), .Y(n272) );
  AOI22X1 U211 ( .A0(N359), .A1(n38), .B0(n206), .B1(in_17bit_b[12]), .Y(n273)
         );
  NAND2X1 U212 ( .A(n276), .B(n275), .Y(N460) );
  AOI22X1 U213 ( .A0(N121), .A1(n281), .B0(N218), .B1(n39), .Y(n275) );
  AOI22X1 U214 ( .A0(N360), .A1(n38), .B0(n206), .B1(in_17bit_b[13]), .Y(n276)
         );
  NAND2X1 U215 ( .A(n279), .B(n278), .Y(N461) );
  AOI22X1 U216 ( .A0(N122), .A1(n281), .B0(N219), .B1(n39), .Y(n278) );
  AOI22X1 U217 ( .A0(N361), .A1(n38), .B0(n206), .B1(in_17bit_b[14]), .Y(n279)
         );
  NAND2X1 U218 ( .A(n283), .B(n282), .Y(N462) );
  AOI22X1 U219 ( .A0(N123), .A1(n281), .B0(N220), .B1(n39), .Y(n282) );
  AOI22X1 U220 ( .A0(N362), .A1(n38), .B0(n206), .B1(in_17bit_b[15]), .Y(n283)
         );
  CLKBUFXL U221 ( .A(in_8bit[1]), .Y(n40) );
  INVX1 U222 ( .A(in_8bit[0]), .Y(n41) );
  INVX1 U223 ( .A(in_8bit[3]), .Y(n43) );
  OAI21XL U224 ( .A0(n22), .A1(n96), .B0(n95), .Y(n101) );
  OAI21XL U225 ( .A0(n23), .A1(n88), .B0(n87), .Y(n93) );
  NOR2XL U226 ( .A(n90), .B(n20), .Y(n92) );
  NAND2XL U227 ( .A(n21), .B(n13), .Y(n160) );
  INVX1 U228 ( .A(n63), .Y(n60) );
  AOI22XL U229 ( .A0(N26), .A1(n25), .B0(in_17bit[13]), .B1(n49), .Y(n274) );
  AOI22XL U230 ( .A0(N18), .A1(n25), .B0(in_17bit[5]), .B1(n49), .Y(n250) );
  AOI22XL U231 ( .A0(N19), .A1(n25), .B0(in_17bit[6]), .B1(n49), .Y(n253) );
  AOI22XL U232 ( .A0(N20), .A1(n25), .B0(in_17bit[7]), .B1(n49), .Y(n256) );
  AOI22XL U233 ( .A0(N21), .A1(n25), .B0(in_17bit[8]), .B1(n49), .Y(n259) );
  AOI22XL U234 ( .A0(N22), .A1(n25), .B0(in_17bit[9]), .B1(n48), .Y(n262) );
  AOI22XL U235 ( .A0(N23), .A1(n25), .B0(in_17bit[10]), .B1(n48), .Y(n265) );
  AOI22XL U236 ( .A0(N24), .A1(n25), .B0(in_17bit[11]), .B1(n49), .Y(n268) );
  AOI22XL U237 ( .A0(N25), .A1(n25), .B0(in_17bit[12]), .B1(n49), .Y(n271) );
  AOI22XL U238 ( .A0(N28), .A1(n25), .B0(in_17bit[15]), .B1(n49), .Y(n280) );
  AOI22XL U239 ( .A0(N16), .A1(n25), .B0(in_17bit[3]), .B1(n49), .Y(n244) );
  NAND2BX1 U240 ( .AN(n63), .B(n6), .Y(n70) );
  AND2X2 U241 ( .A(n99), .B(n13), .Y(n29) );
  NAND2X1 U242 ( .A(n35), .B(n5), .Y(n63) );
  BUFX3 U243 ( .A(n284), .Y(n38) );
  OAI2BB1X1 U244 ( .A0N(n185), .A1N(n14), .B0(n183), .Y(n284) );
  NAND2BX1 U245 ( .AN(n227), .B(n31), .Y(n183) );
  BUFX3 U246 ( .A(n285), .Y(n39) );
  OAI2BB1X1 U247 ( .A0N(n31), .A1N(n185), .B0(n184), .Y(n285) );
  NAND2BX1 U248 ( .AN(n227), .B(n14), .Y(n184) );
  AND2X2 U249 ( .A(n29), .B(n3), .Y(n30) );
  NAND2X1 U250 ( .A(n181), .B(n180), .Y(n281) );
  NAND3X1 U251 ( .A(n232), .B(in_8bit[5]), .C(n179), .Y(n180) );
  NAND4BXL U252 ( .AN(n42), .B(n233), .C(n188), .D(n40), .Y(n181) );
  OAI2BB1X1 U253 ( .A0N(n232), .A1N(n188), .B0(n187), .Y(n206) );
  NAND3BX1 U254 ( .AN(n186), .B(n233), .C(in_8bit[5]), .Y(n187) );
  AND2X2 U255 ( .A(n182), .B(n41), .Y(n31) );
  NAND2X1 U256 ( .A(n83), .B(n8), .Y(n94) );
  NAND2X1 U257 ( .A(n91), .B(n7), .Y(n158) );
  NAND2X1 U258 ( .A(n75), .B(n12), .Y(n86) );
  NAND2BX1 U259 ( .AN(n70), .B(n11), .Y(n78) );
  AND2X2 U260 ( .A(n30), .B(n1), .Y(n32) );
  AND2X2 U261 ( .A(n32), .B(n2), .Y(n33) );
  INVX1 U262 ( .A(in_17bit[3]), .Y(n192) );
  INVX1 U263 ( .A(in_17bit[5]), .Y(n194) );
  INVX1 U264 ( .A(in_17bit[6]), .Y(n195) );
  INVX1 U265 ( .A(in_17bit[7]), .Y(n196) );
  INVX1 U266 ( .A(in_17bit[8]), .Y(n197) );
  INVX1 U267 ( .A(in_17bit[9]), .Y(n198) );
  INVX1 U268 ( .A(in_17bit[10]), .Y(n199) );
  INVX1 U269 ( .A(in_17bit[11]), .Y(n200) );
  INVX1 U270 ( .A(in_17bit[12]), .Y(n201) );
  INVX1 U271 ( .A(in_17bit[13]), .Y(n202) );
  INVX1 U272 ( .A(in_17bit[14]), .Y(n203) );
  INVX1 U273 ( .A(in_17bit[15]), .Y(n204) );
  INVX1 U274 ( .A(in_17bit[1]), .Y(n190) );
  INVX1 U275 ( .A(in_17bit[2]), .Y(n191) );
  INVX1 U276 ( .A(in_17bit[4]), .Y(n193) );
  INVX1 U277 ( .A(in_17bit[0]), .Y(n189) );
  INVX1 U278 ( .A(n72), .Y(n73) );
  INVX1 U279 ( .A(n80), .Y(n81) );
  XNOR2X1 U280 ( .A(n15), .B(sub_add_75_b0_carry[13]), .Y(n34) );
  INVX1 U281 ( .A(n65), .Y(n66) );
  INVX1 U282 ( .A(n88), .Y(n89) );
  INVX1 U283 ( .A(n57), .Y(n58) );
  INVX1 U284 ( .A(n96), .Y(n97) );
  AOI2BB2X1 U285 ( .B0(n164), .B1(n23), .A0N(n22), .A1N(neg_mul[15]), .Y(n168)
         );
  INVX1 U286 ( .A(n163), .Y(n164) );
  INVX1 U287 ( .A(n51), .Y(n52) );
  MX2X1 U288 ( .A(neg_mul[22]), .B(N480), .S0(n177), .Y(out[15]) );
  MX2X1 U289 ( .A(neg_mul[23]), .B(N481), .S0(n177), .Y(out[16]) );
  NAND4BBX1 U290 ( .AN(n38), .BN(n39), .C(n234), .D(n287), .Y(N446) );
  AOI2BB1X1 U291 ( .A0N(n231), .A1N(n230), .B0(n281), .Y(n234) );
  OR4X2 U292 ( .A(n40), .B(in_8bit[0]), .C(n44), .D(in_8bit[3]), .Y(n230) );
  INVX1 U293 ( .A(in_8bit[4]), .Y(n178) );
  NOR3BXL U294 ( .AN(n22), .B(in_8bit[5]), .C(in_8bit[4]), .Y(n188) );
  NOR2X1 U295 ( .A(out[0]), .B(neg_mul[8]), .Y(n35) );
  NOR2X1 U296 ( .A(in_8bit[6]), .B(in_8bit[4]), .Y(n226) );
  NAND2X1 U297 ( .A(out[0]), .B(neg_mul[8]), .Y(n51) );
  NAND2BX1 U298 ( .AN(n35), .B(neg_mul[9]), .Y(n57) );
  NAND2X1 U299 ( .A(neg_mul[10]), .B(n63), .Y(n65) );
  NAND2X1 U300 ( .A(neg_mul[14]), .B(n94), .Y(n96) );
  NAND2X1 U301 ( .A(neg_mul[11]), .B(n70), .Y(n72) );
  NAND2X1 U302 ( .A(neg_mul[13]), .B(n86), .Y(n88) );
  NAND2X1 U303 ( .A(neg_mul[15]), .B(n158), .Y(n163) );
  NAND2X1 U304 ( .A(neg_mul[12]), .B(n78), .Y(n80) );
  INVXL U305 ( .A(in_8bit[2]), .Y(n45) );
  AOI211X4 U306 ( .A0(n37), .A1(n93), .B0(n92), .C0(n91), .Y(out[6]) );
  AOI211X4 U307 ( .A0(n37), .A1(n171), .B0(n170), .C0(n29), .Y(out[8]) );
  OAI21XL U308 ( .A0(n22), .A1(n72), .B0(n71), .Y(n77) );
  OAI21XL U309 ( .A0(n22), .A1(n80), .B0(n79), .Y(n85) );
  OAI21XL U310 ( .A0(n22), .A1(n163), .B0(n160), .Y(n171) );
  AOI2BB2X1 U311 ( .B0(n73), .B1(n23), .A0N(n21), .A1N(neg_mul[11]), .Y(n74)
         );
  NOR2XL U312 ( .A(n22), .B(n178), .Y(n179) );
  NAND2XL U313 ( .A(n21), .B(n11), .Y(n71) );
  NAND2XL U314 ( .A(n21), .B(n12), .Y(n79) );
  NAND2X1 U315 ( .A(n23), .B(n8), .Y(n87) );
  NOR2X2 U316 ( .A(n30), .B(n174), .Y(n173) );
  AOI22XL U317 ( .A0(N17), .A1(n25), .B0(in_17bit[4]), .B1(n49), .Y(n247) );
  AOI22XL U318 ( .A0(in_17bit[0]), .A1(n25), .B0(in_17bit[0]), .B1(n48), .Y(
        n235) );
  AOI22XL U319 ( .A0(N15), .A1(n25), .B0(in_17bit[2]), .B1(n49), .Y(n241) );
  AOI22XL U320 ( .A0(N14), .A1(n25), .B0(in_17bit[1]), .B1(n49), .Y(n238) );
  AOI211X2 U321 ( .A0(n37), .A1(n101), .B0(n100), .C0(n99), .Y(n289) );
  XNOR2X4 U322 ( .A(n172), .B(n3), .Y(out[9]) );
  XNOR2X4 U323 ( .A(n175), .B(n4), .Y(out[12]) );
  AND2X1 U324 ( .A(add_1_root_r112_carry_20_), .B(in_17bit_b[16]), .Y(
        add_1_root_r112_SUM_21_) );
  XOR2X1 U325 ( .A(in_17bit_b[16]), .B(add_1_root_r112_carry_20_), .Y(
        add_1_root_r112_SUM_20_) );
  AND2X1 U326 ( .A(add_1_root_r112_carry_19_), .B(in_17bit_b[15]), .Y(
        add_1_root_r112_carry_20_) );
  XOR2X1 U327 ( .A(in_17bit_b[15]), .B(add_1_root_r112_carry_19_), .Y(
        add_1_root_r112_SUM_19_) );
  AND2X1 U328 ( .A(add_1_root_r112_carry_18_), .B(in_17bit_b[14]), .Y(
        add_1_root_r112_carry_19_) );
  XOR2X1 U329 ( .A(in_17bit_b[14]), .B(add_1_root_r112_carry_18_), .Y(
        add_1_root_r112_SUM_18_) );
  AND2X1 U330 ( .A(add_1_root_r112_carry_17_), .B(in_17bit_b[13]), .Y(
        add_1_root_r112_carry_18_) );
  XOR2X1 U331 ( .A(in_17bit_b[13]), .B(add_1_root_r112_carry_17_), .Y(
        add_1_root_r112_SUM_17_) );
  AND2X1 U332 ( .A(add_2_root_r119_carry_21_), .B(in_17bit_b[16]), .Y(
        add_2_root_r119_SUM_22_) );
  XOR2X1 U333 ( .A(in_17bit_b[16]), .B(add_2_root_r119_carry_21_), .Y(
        add_2_root_r119_SUM_21_) );
  AND2X1 U334 ( .A(n205), .B(in_17bit_b[0]), .Y(add_2_root_r119_carry_6_) );
  AND2X1 U335 ( .A(add_1_root_r119_carry[22]), .B(in_17bit_b[16]), .Y(
        add_1_root_r119_SUM_23_) );
  XOR2X1 U336 ( .A(in_17bit_b[16]), .B(add_1_root_r119_carry[22]), .Y(
        add_1_root_r119_SUM_22_) );
  AND2X1 U337 ( .A(add_1_root_r119_carry[21]), .B(in_17bit_b[15]), .Y(
        add_1_root_r119_carry[22]) );
  XOR2X1 U338 ( .A(in_17bit_b[15]), .B(add_1_root_r119_carry[21]), .Y(
        add_1_root_r119_SUM_21_) );
  AND2X1 U339 ( .A(add_1_root_r119_carry[20]), .B(in_17bit_b[14]), .Y(
        add_1_root_r119_carry[21]) );
  XOR2X1 U340 ( .A(in_17bit_b[14]), .B(add_1_root_r119_carry[20]), .Y(
        add_1_root_r119_SUM_20_) );
  AND2X1 U341 ( .A(add_1_root_r119_A_6_), .B(in_17bit_b[0]), .Y(
        add_1_root_r119_carry[7]) );
  XOR2X1 U342 ( .A(in_17bit_b[0]), .B(add_1_root_r119_A_6_), .Y(
        add_1_root_r119_SUM_6_) );
  AND2X1 U343 ( .A(add_3_root_r119_carry_18_), .B(in_17bit_b[16]), .Y(
        add_1_root_r119_A_19_) );
  XOR2X1 U344 ( .A(in_17bit_b[16]), .B(add_3_root_r119_carry_18_), .Y(
        add_1_root_r119_A_18_) );
  XOR2X1 U345 ( .A(in_17bit_b[0]), .B(n205), .Y(add_1_root_r119_A_2_) );
  AND2X1 U346 ( .A(add_2_root_r115_carry_19_), .B(in_17bit_b[16]), .Y(
        add_2_root_r115_SUM_20_) );
  XOR2X1 U347 ( .A(in_17bit_b[16]), .B(add_2_root_r115_carry_19_), .Y(
        add_2_root_r115_SUM_19_) );
  AND2X1 U348 ( .A(add_2_root_r115_carry_18_), .B(in_17bit_b[15]), .Y(
        add_2_root_r115_carry_19_) );
  XOR2X1 U349 ( .A(in_17bit_b[15]), .B(add_2_root_r115_carry_18_), .Y(
        add_2_root_r115_SUM_18_) );
  XOR2X1 U350 ( .A(in_17bit_b[0]), .B(in_17bit_b[2]), .Y(
        add_2_root_r115_SUM_3_) );
  AND2X1 U351 ( .A(add_1_root_r115_carry_22_), .B(in_17bit_b[16]), .Y(
        add_1_root_r115_SUM_23_) );
  XOR2X1 U352 ( .A(in_17bit_b[16]), .B(add_1_root_r115_carry_22_), .Y(
        add_1_root_r115_SUM_22_) );
  AND2X1 U353 ( .A(add_1_root_r115_carry_21_), .B(in_17bit_b[15]), .Y(
        add_1_root_r115_carry_22_) );
  XOR2X1 U354 ( .A(in_17bit_b[15]), .B(add_1_root_r115_carry_21_), .Y(
        add_1_root_r115_SUM_21_) );
  AND2X1 U355 ( .A(in_17bit_b[2]), .B(in_17bit_b[0]), .Y(
        add_1_root_r115_carry_7_) );
  XOR2X1 U356 ( .A(n49), .B(sub_add_54_b0_carry[16]), .Y(N29) );
  AND2X1 U357 ( .A(sub_add_54_b0_carry[15]), .B(n204), .Y(
        sub_add_54_b0_carry[16]) );
  XOR2X1 U358 ( .A(n204), .B(sub_add_54_b0_carry[15]), .Y(N28) );
  AND2X1 U359 ( .A(sub_add_54_b0_carry[14]), .B(n203), .Y(
        sub_add_54_b0_carry[15]) );
  XOR2X1 U360 ( .A(n203), .B(sub_add_54_b0_carry[14]), .Y(N27) );
  AND2X1 U361 ( .A(sub_add_54_b0_carry[13]), .B(n202), .Y(
        sub_add_54_b0_carry[14]) );
  XOR2X1 U362 ( .A(n202), .B(sub_add_54_b0_carry[13]), .Y(N26) );
  AND2X1 U363 ( .A(sub_add_54_b0_carry[12]), .B(n201), .Y(
        sub_add_54_b0_carry[13]) );
  XOR2X1 U364 ( .A(n201), .B(sub_add_54_b0_carry[12]), .Y(N25) );
  AND2X1 U365 ( .A(sub_add_54_b0_carry[11]), .B(n200), .Y(
        sub_add_54_b0_carry[12]) );
  XOR2X1 U366 ( .A(n200), .B(sub_add_54_b0_carry[11]), .Y(N24) );
  AND2X1 U367 ( .A(sub_add_54_b0_carry[10]), .B(n199), .Y(
        sub_add_54_b0_carry[11]) );
  XOR2X1 U368 ( .A(n199), .B(sub_add_54_b0_carry[10]), .Y(N23) );
  AND2X1 U369 ( .A(sub_add_54_b0_carry[9]), .B(n198), .Y(
        sub_add_54_b0_carry[10]) );
  XOR2X1 U370 ( .A(n198), .B(sub_add_54_b0_carry[9]), .Y(N22) );
  AND2X1 U371 ( .A(sub_add_54_b0_carry[8]), .B(n197), .Y(
        sub_add_54_b0_carry[9]) );
  XOR2X1 U372 ( .A(n197), .B(sub_add_54_b0_carry[8]), .Y(N21) );
  AND2X1 U373 ( .A(sub_add_54_b0_carry[7]), .B(n196), .Y(
        sub_add_54_b0_carry[8]) );
  XOR2X1 U374 ( .A(n196), .B(sub_add_54_b0_carry[7]), .Y(N20) );
  AND2X1 U375 ( .A(sub_add_54_b0_carry[6]), .B(n195), .Y(
        sub_add_54_b0_carry[7]) );
  XOR2X1 U376 ( .A(n195), .B(sub_add_54_b0_carry[6]), .Y(N19) );
  AND2X1 U377 ( .A(sub_add_54_b0_carry[5]), .B(n194), .Y(
        sub_add_54_b0_carry[6]) );
  XOR2X1 U378 ( .A(n194), .B(sub_add_54_b0_carry[5]), .Y(N18) );
  AND2X1 U379 ( .A(sub_add_54_b0_carry[4]), .B(n193), .Y(
        sub_add_54_b0_carry[5]) );
  XOR2X1 U380 ( .A(n193), .B(sub_add_54_b0_carry[4]), .Y(N17) );
  AND2X1 U381 ( .A(sub_add_54_b0_carry[3]), .B(n192), .Y(
        sub_add_54_b0_carry[4]) );
  XOR2X1 U382 ( .A(n192), .B(sub_add_54_b0_carry[3]), .Y(N16) );
  AND2X1 U383 ( .A(sub_add_54_b0_carry[2]), .B(n191), .Y(
        sub_add_54_b0_carry[3]) );
  XOR2X1 U384 ( .A(n191), .B(sub_add_54_b0_carry[2]), .Y(N15) );
  AND2X1 U385 ( .A(n189), .B(n190), .Y(sub_add_54_b0_carry[2]) );
  XOR2X1 U386 ( .A(n190), .B(n189), .Y(N14) );
  XOR2X1 U387 ( .A(n17), .B(sub_add_75_b0_carry[16]), .Y(N481) );
  AND2X1 U388 ( .A(sub_add_75_b0_carry[15]), .B(n10), .Y(
        sub_add_75_b0_carry[16]) );
  XOR2X1 U389 ( .A(n10), .B(sub_add_75_b0_carry[15]), .Y(N480) );
  AND2X1 U390 ( .A(sub_add_75_b0_carry[14]), .B(n9), .Y(
        sub_add_75_b0_carry[15]) );
  XOR2X1 U391 ( .A(n9), .B(sub_add_75_b0_carry[14]), .Y(N479) );
  AND2X1 U392 ( .A(sub_add_75_b0_carry[13]), .B(n15), .Y(
        sub_add_75_b0_carry[14]) );
  AND2X1 U393 ( .A(n33), .B(n4), .Y(sub_add_75_b0_carry[13]) );
  AND2X1 U394 ( .A(in_17bit_b[0]), .B(in_17bit_b[4]), .Y(
        add_1_root_r112_carry_5_) );
endmodule


module multi16_10_DW01_add_0 ( A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, 
        A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, 
        A_4_, B_23_, B_22_, B_21_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, 
        B_14_, B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, 
        SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, 
        SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, 
        SUM_7_ );
  input A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_,
         A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, B_23_, B_22_,
         B_21_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_,
         B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_;
  output SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_,
         SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_,
         SUM_8_, SUM_7_;
  wire   n1, n2, n3, n4;
  wire   [23:7] carry;

  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry[7]), .CO(carry[8]), .S(SUM_7_)
         );
  ADDFX2 U1_21 ( .A(A_21_), .B(B_21_), .CI(carry[21]), .CO(carry[22]), .S(
        SUM_21_) );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry[20]), .CO(carry[21]), .S(
        SUM_20_) );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry[19]), .CO(carry[20]), .S(
        SUM_19_) );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry[18]), .CO(carry[19]), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry[17]), .CO(carry[18]), .S(
        SUM_17_) );
  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry[16]), .CO(carry[17]), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry[15]), .CO(carry[16]), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry[14]), .CO(carry[15]), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry[13]), .CO(carry[14]), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry[12]), .CO(carry[13]), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry[11]), .CO(carry[12]), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry[10]), .CO(carry[11]), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry[9]), .CO(carry[10]), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry[8]), .CO(carry[9]), .S(SUM_8_)
         );
  ADDFX2 U1_22 ( .A(A_22_), .B(B_22_), .CI(carry[22]), .CO(carry[23]), .S(
        SUM_22_) );
  AND2X2 U1 ( .A(A_4_), .B(B_4_), .Y(n1) );
  XOR2X1 U2 ( .A(B_23_), .B(carry[23]), .Y(SUM_23_) );
  OAI2BB1X1 U3 ( .A0N(n2), .A1N(A_6_), .B0(n3), .Y(carry[7]) );
  OAI21XL U4 ( .A0(A_6_), .A1(n2), .B0(B_6_), .Y(n3) );
  OAI2BB1X1 U5 ( .A0N(n1), .A1N(A_5_), .B0(n4), .Y(n2) );
  OAI21XL U6 ( .A0(A_5_), .A1(n1), .B0(B_5_), .Y(n4) );
endmodule


module multi16_10_DW01_add_4 ( A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, 
        A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, 
        B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, 
        B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, SUM_22_, SUM_21_, SUM_20_, 
        SUM_19_, SUM_18_, SUM_17_, SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, 
        SUM_11_, SUM_10_, SUM_9_, SUM_8_, SUM_7_ );
  input A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_,
         A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, B_20_, B_19_,
         B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, B_10_, B_9_,
         B_8_, B_7_, B_6_, B_5_;
  output SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_,
         SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_,
         SUM_7_;
  wire   carry_21_, carry_20_, carry_19_, carry_18_, carry_17_, carry_16_,
         carry_15_, carry_14_, carry_13_, carry_12_, carry_11_, carry_10_,
         carry_9_, carry_8_, carry_7_, n1;

  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry_16_), .CO(carry_17_), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry_15_), .CO(carry_16_), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry_14_), .CO(carry_15_), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry_13_), .CO(carry_14_), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry_12_), .CO(carry_13_), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry_11_), .CO(carry_12_), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry_10_), .CO(carry_11_), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry_9_), .CO(carry_10_), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry_8_), .CO(carry_9_), .S(SUM_8_)
         );
  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry_7_), .CO(carry_8_), .S(SUM_7_)
         );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry_20_), .CO(carry_21_), .S(
        SUM_20_) );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry_19_), .CO(carry_20_), .S(
        SUM_19_) );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry_18_), .CO(carry_19_), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry_17_), .CO(carry_18_), .S(
        SUM_17_) );
  ADDFX2 U1_21 ( .A(A_21_), .B(B_21_), .CI(carry_21_), .CO(SUM_22_), .S(
        SUM_21_) );
  OAI2BB1X1 U1 ( .A0N(A_6_), .A1N(B_6_), .B0(n1), .Y(carry_7_) );
  OAI211X1 U2 ( .A0(B_6_), .A1(A_6_), .B0(A_5_), .C0(B_5_), .Y(n1) );
endmodule


module multi16_10_DW01_add_6 ( A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, 
        A_16_, A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, 
        A_6_, A_5_, A_4_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, 
        B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, 
        SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, 
        SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, 
        SUM_7_ );
  input A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_,
         A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, B_20_,
         B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, B_10_,
         B_9_, B_8_, B_7_, B_6_, B_5_, B_4_;
  output SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_,
         SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_,
         SUM_8_, SUM_7_;
  wire   n1, n2, n3, n4, n5, n6;
  wire   [21:7] carry;

  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry[7]), .CO(carry[8]), .S(SUM_7_)
         );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry[18]), .CO(carry[19]), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry[17]), .CO(carry[18]), .S(
        SUM_17_) );
  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry[16]), .CO(carry[17]), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry[15]), .CO(carry[16]), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry[14]), .CO(carry[15]), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry[13]), .CO(carry[14]), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry[12]), .CO(carry[13]), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry[11]), .CO(carry[12]), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry[10]), .CO(carry[11]), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry[9]), .CO(carry[10]), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry[8]), .CO(carry[9]), .S(SUM_8_)
         );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry[19]), .CO(carry[20]), .S(
        SUM_19_) );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry[20]), .CO(carry[21]), .S(
        SUM_20_) );
  AND2X2 U1 ( .A(A_22_), .B(n2), .Y(n1) );
  AND2X2 U2 ( .A(A_21_), .B(carry[21]), .Y(n2) );
  AND2X2 U3 ( .A(A_4_), .B(B_4_), .Y(n3) );
  XOR2X1 U4 ( .A(A_23_), .B(n1), .Y(SUM_23_) );
  XOR2X1 U5 ( .A(A_21_), .B(carry[21]), .Y(SUM_21_) );
  XOR2X1 U6 ( .A(A_22_), .B(n2), .Y(SUM_22_) );
  OAI2BB1X1 U7 ( .A0N(n4), .A1N(A_6_), .B0(n5), .Y(carry[7]) );
  OAI21XL U8 ( .A0(A_6_), .A1(n4), .B0(B_6_), .Y(n5) );
  OAI2BB1X1 U9 ( .A0N(n3), .A1N(A_5_), .B0(n6), .Y(n4) );
  OAI21XL U10 ( .A0(A_5_), .A1(n3), .B0(B_5_), .Y(n6) );
endmodule


module multi16_10 ( in_17bit, in_8bit, out );
  input [16:0] in_17bit;
  input [7:0] in_8bit;
  output [16:0] out;
  wire   N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27,
         N28, N29, N108, N109, N110, N111, N112, N113, N114, N115, N116, N117,
         N118, N119, N120, N121, N122, N123, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220,
         N221, N347, N348, N349, N350, N351, N352, N353, N354, N355, N356,
         N357, N358, N359, N360, N361, N362, N363, N446, N447, N448, N449,
         N450, N451, N452, N453, N454, N455, N456, N457, N458, N459, N460,
         N461, N462, N463, N479, N480, N481, add_2_root_r119_carry_10_,
         add_2_root_r119_carry_11_, add_2_root_r119_carry_12_,
         add_2_root_r119_carry_13_, add_2_root_r119_carry_14_,
         add_2_root_r119_carry_15_, add_2_root_r119_carry_16_,
         add_2_root_r119_carry_17_, add_2_root_r119_carry_18_,
         add_2_root_r119_carry_19_, add_2_root_r119_carry_20_,
         add_2_root_r119_carry_21_, add_2_root_r119_carry_7_,
         add_2_root_r119_carry_8_, add_2_root_r119_carry_9_,
         add_2_root_r119_SUM_6_, add_2_root_r119_SUM_7_,
         add_2_root_r119_SUM_8_, add_2_root_r119_SUM_9_,
         add_2_root_r119_SUM_10_, add_2_root_r119_SUM_11_,
         add_2_root_r119_SUM_12_, add_2_root_r119_SUM_13_,
         add_2_root_r119_SUM_14_, add_2_root_r119_SUM_15_,
         add_2_root_r119_SUM_16_, add_2_root_r119_SUM_17_,
         add_2_root_r119_SUM_18_, add_2_root_r119_SUM_19_,
         add_2_root_r119_SUM_20_, add_2_root_r119_SUM_21_,
         add_2_root_r119_SUM_22_, add_1_root_r119_SUM_6_,
         add_1_root_r119_SUM_7_, add_1_root_r119_SUM_8_,
         add_1_root_r119_SUM_9_, add_1_root_r119_SUM_10_,
         add_1_root_r119_SUM_11_, add_1_root_r119_SUM_12_,
         add_1_root_r119_SUM_13_, add_1_root_r119_SUM_14_,
         add_1_root_r119_SUM_15_, add_1_root_r119_SUM_16_,
         add_1_root_r119_SUM_17_, add_1_root_r119_SUM_18_,
         add_1_root_r119_SUM_19_, add_1_root_r119_SUM_20_,
         add_1_root_r119_SUM_21_, add_1_root_r119_SUM_22_,
         add_1_root_r119_SUM_23_, add_1_root_r119_A_2_, add_1_root_r119_A_3_,
         add_1_root_r119_A_4_, add_1_root_r119_A_5_, add_1_root_r119_A_6_,
         add_1_root_r119_A_7_, add_1_root_r119_A_8_, add_1_root_r119_A_9_,
         add_1_root_r119_A_10_, add_1_root_r119_A_11_, add_1_root_r119_A_12_,
         add_1_root_r119_A_13_, add_1_root_r119_A_14_, add_1_root_r119_A_15_,
         add_1_root_r119_A_16_, add_1_root_r119_A_17_, add_1_root_r119_A_18_,
         add_1_root_r119_A_19_, add_3_root_r119_carry_10_,
         add_3_root_r119_carry_11_, add_3_root_r119_carry_12_,
         add_3_root_r119_carry_13_, add_3_root_r119_carry_14_,
         add_3_root_r119_carry_15_, add_3_root_r119_carry_16_,
         add_3_root_r119_carry_17_, add_3_root_r119_carry_18_,
         add_3_root_r119_carry_3_, add_3_root_r119_carry_4_,
         add_3_root_r119_carry_5_, add_3_root_r119_carry_6_,
         add_3_root_r119_carry_7_, add_3_root_r119_carry_8_,
         add_3_root_r119_carry_9_, add_1_root_r112_carry_10_,
         add_1_root_r112_carry_11_, add_1_root_r112_carry_12_,
         add_1_root_r112_carry_13_, add_1_root_r112_carry_14_,
         add_1_root_r112_carry_15_, add_1_root_r112_carry_16_,
         add_1_root_r112_carry_17_, add_1_root_r112_carry_18_,
         add_1_root_r112_carry_19_, add_1_root_r112_carry_20_,
         add_1_root_r112_carry_5_, add_1_root_r112_carry_6_,
         add_1_root_r112_carry_7_, add_1_root_r112_carry_8_,
         add_1_root_r112_carry_9_, add_1_root_r112_SUM_1_,
         add_1_root_r112_SUM_2_, add_1_root_r112_SUM_3_,
         add_1_root_r112_SUM_4_, add_1_root_r112_SUM_5_,
         add_1_root_r112_SUM_6_, add_1_root_r112_SUM_7_,
         add_1_root_r112_SUM_8_, add_1_root_r112_SUM_9_,
         add_1_root_r112_SUM_10_, add_1_root_r112_SUM_11_,
         add_1_root_r112_SUM_12_, add_1_root_r112_SUM_13_,
         add_1_root_r112_SUM_14_, add_1_root_r112_SUM_15_,
         add_1_root_r112_SUM_16_, add_1_root_r112_SUM_17_,
         add_1_root_r112_SUM_18_, add_1_root_r112_SUM_19_,
         add_1_root_r112_SUM_20_, add_1_root_r112_SUM_21_,
         add_2_root_r115_carry_10_, add_2_root_r115_carry_11_,
         add_2_root_r115_carry_12_, add_2_root_r115_carry_13_,
         add_2_root_r115_carry_14_, add_2_root_r115_carry_15_,
         add_2_root_r115_carry_16_, add_2_root_r115_carry_17_,
         add_2_root_r115_carry_18_, add_2_root_r115_carry_19_,
         add_2_root_r115_carry_4_, add_2_root_r115_carry_5_,
         add_2_root_r115_carry_6_, add_2_root_r115_carry_7_,
         add_2_root_r115_carry_8_, add_2_root_r115_carry_9_,
         add_2_root_r115_SUM_4_, add_2_root_r115_SUM_5_,
         add_2_root_r115_SUM_6_, add_2_root_r115_SUM_7_,
         add_2_root_r115_SUM_8_, add_2_root_r115_SUM_9_,
         add_2_root_r115_SUM_10_, add_2_root_r115_SUM_11_,
         add_2_root_r115_SUM_12_, add_2_root_r115_SUM_13_,
         add_2_root_r115_SUM_14_, add_2_root_r115_SUM_15_,
         add_2_root_r115_SUM_16_, add_2_root_r115_SUM_17_,
         add_2_root_r115_SUM_18_, add_2_root_r115_SUM_19_,
         add_2_root_r115_SUM_20_, add_1_root_r115_carry_10_,
         add_1_root_r115_carry_11_, add_1_root_r115_carry_12_,
         add_1_root_r115_carry_13_, add_1_root_r115_carry_14_,
         add_1_root_r115_carry_15_, add_1_root_r115_carry_16_,
         add_1_root_r115_carry_17_, add_1_root_r115_carry_18_,
         add_1_root_r115_carry_19_, add_1_root_r115_carry_20_,
         add_1_root_r115_carry_21_, add_1_root_r115_carry_22_,
         add_1_root_r115_carry_8_, add_1_root_r115_carry_9_,
         add_1_root_r115_SUM_6_, add_1_root_r115_SUM_7_,
         add_1_root_r115_SUM_8_, add_1_root_r115_SUM_9_,
         add_1_root_r115_SUM_10_, add_1_root_r115_SUM_11_,
         add_1_root_r115_SUM_12_, add_1_root_r115_SUM_13_,
         add_1_root_r115_SUM_14_, add_1_root_r115_SUM_15_,
         add_1_root_r115_SUM_16_, add_1_root_r115_SUM_17_,
         add_1_root_r115_SUM_18_, add_1_root_r115_SUM_19_,
         add_1_root_r115_SUM_20_, add_1_root_r115_SUM_21_,
         add_1_root_r115_SUM_22_, add_1_root_r115_SUM_23_, n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n158, n160, n161,
         n162, n163, n164, n168, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274;
  wire   [16:0] in_17bit_b;
  wire   [23:8] neg_mul;
  wire   [16:13] sub_add_75_b0_carry;
  wire   [16:2] sub_add_54_b0_carry;
  wire   [22:7] add_1_root_r119_carry;

  multi16_10_DW01_add_0 add_0_root_r119 ( .A_22_(add_2_root_r119_SUM_22_), 
        .A_21_(add_2_root_r119_SUM_21_), .A_20_(add_2_root_r119_SUM_20_), 
        .A_19_(add_2_root_r119_SUM_19_), .A_18_(add_2_root_r119_SUM_18_), 
        .A_17_(add_2_root_r119_SUM_17_), .A_16_(add_2_root_r119_SUM_16_), 
        .A_15_(add_2_root_r119_SUM_15_), .A_14_(add_2_root_r119_SUM_14_), 
        .A_13_(add_2_root_r119_SUM_13_), .A_12_(add_2_root_r119_SUM_12_), 
        .A_11_(add_2_root_r119_SUM_11_), .A_10_(add_2_root_r119_SUM_10_), 
        .A_9_(add_2_root_r119_SUM_9_), .A_8_(add_2_root_r119_SUM_8_), .A_7_(
        add_2_root_r119_SUM_7_), .A_6_(add_2_root_r119_SUM_6_), .A_5_(
        add_1_root_r119_A_2_), .A_4_(in_17bit_b[0]), .B_23_(
        add_1_root_r119_SUM_23_), .B_22_(add_1_root_r119_SUM_22_), .B_21_(
        add_1_root_r119_SUM_21_), .B_20_(add_1_root_r119_SUM_20_), .B_19_(
        add_1_root_r119_SUM_19_), .B_18_(add_1_root_r119_SUM_18_), .B_17_(
        add_1_root_r119_SUM_17_), .B_16_(add_1_root_r119_SUM_16_), .B_15_(
        add_1_root_r119_SUM_15_), .B_14_(add_1_root_r119_SUM_14_), .B_13_(
        add_1_root_r119_SUM_13_), .B_12_(add_1_root_r119_SUM_12_), .B_11_(
        add_1_root_r119_SUM_11_), .B_10_(add_1_root_r119_SUM_10_), .B_9_(
        add_1_root_r119_SUM_9_), .B_8_(add_1_root_r119_SUM_8_), .B_7_(
        add_1_root_r119_SUM_7_), .B_6_(add_1_root_r119_SUM_6_), .B_5_(
        add_1_root_r119_A_5_), .B_4_(add_1_root_r119_A_4_), .SUM_23_(N363), 
        .SUM_22_(N362), .SUM_21_(N361), .SUM_20_(N360), .SUM_19_(N359), 
        .SUM_18_(N358), .SUM_17_(N357), .SUM_16_(N356), .SUM_15_(N355), 
        .SUM_14_(N354), .SUM_13_(N353), .SUM_12_(N352), .SUM_11_(N351), 
        .SUM_10_(N350), .SUM_9_(N349), .SUM_8_(N348), .SUM_7_(N347) );
  multi16_10_DW01_add_4 add_0_root_r112 ( .A_21_(in_17bit_b[16]), .A_20_(
        in_17bit_b[15]), .A_19_(in_17bit_b[14]), .A_18_(in_17bit_b[13]), 
        .A_17_(in_17bit_b[12]), .A_16_(in_17bit_b[11]), .A_15_(in_17bit_b[10]), 
        .A_14_(in_17bit_b[9]), .A_13_(in_17bit_b[8]), .A_12_(in_17bit_b[7]), 
        .A_11_(in_17bit_b[6]), .A_10_(in_17bit_b[5]), .A_9_(in_17bit_b[4]), 
        .A_8_(in_17bit_b[3]), .A_7_(in_17bit_b[2]), .A_6_(in_17bit_b[1]), 
        .A_5_(in_17bit_b[0]), .B_21_(add_1_root_r112_SUM_21_), .B_20_(
        add_1_root_r112_SUM_20_), .B_19_(add_1_root_r112_SUM_19_), .B_18_(
        add_1_root_r112_SUM_18_), .B_17_(add_1_root_r112_SUM_17_), .B_16_(
        add_1_root_r112_SUM_16_), .B_15_(add_1_root_r112_SUM_15_), .B_14_(
        add_1_root_r112_SUM_14_), .B_13_(add_1_root_r112_SUM_13_), .B_12_(
        add_1_root_r112_SUM_12_), .B_11_(add_1_root_r112_SUM_11_), .B_10_(
        add_1_root_r112_SUM_10_), .B_9_(add_1_root_r112_SUM_9_), .B_8_(
        add_1_root_r112_SUM_8_), .B_7_(add_1_root_r112_SUM_7_), .B_6_(
        add_1_root_r112_SUM_6_), .B_5_(add_1_root_r112_SUM_5_), .SUM_22_(N123), 
        .SUM_21_(N122), .SUM_20_(N121), .SUM_19_(N120), .SUM_18_(N119), 
        .SUM_17_(N118), .SUM_16_(N117), .SUM_15_(N116), .SUM_14_(N115), 
        .SUM_13_(N114), .SUM_12_(N113), .SUM_11_(N112), .SUM_10_(N111), 
        .SUM_9_(N110), .SUM_8_(N109), .SUM_7_(N108) );
  multi16_10_DW01_add_6 add_0_root_r115 ( .A_23_(add_1_root_r115_SUM_23_), 
        .A_22_(add_1_root_r115_SUM_22_), .A_21_(add_1_root_r115_SUM_21_), 
        .A_20_(add_1_root_r115_SUM_20_), .A_19_(add_1_root_r115_SUM_19_), 
        .A_18_(add_1_root_r115_SUM_18_), .A_17_(add_1_root_r115_SUM_17_), 
        .A_16_(add_1_root_r115_SUM_16_), .A_15_(add_1_root_r115_SUM_15_), 
        .A_14_(add_1_root_r115_SUM_14_), .A_13_(add_1_root_r115_SUM_13_), 
        .A_12_(add_1_root_r115_SUM_12_), .A_11_(add_1_root_r115_SUM_11_), 
        .A_10_(add_1_root_r115_SUM_10_), .A_9_(add_1_root_r115_SUM_9_), .A_8_(
        add_1_root_r115_SUM_8_), .A_7_(add_1_root_r115_SUM_7_), .A_6_(
        add_1_root_r115_SUM_6_), .A_5_(in_17bit_b[1]), .A_4_(in_17bit_b[0]), 
        .B_20_(add_2_root_r115_SUM_20_), .B_19_(add_2_root_r115_SUM_19_), 
        .B_18_(add_2_root_r115_SUM_18_), .B_17_(add_2_root_r115_SUM_17_), 
        .B_16_(add_2_root_r115_SUM_16_), .B_15_(add_2_root_r115_SUM_15_), 
        .B_14_(add_2_root_r115_SUM_14_), .B_13_(add_2_root_r115_SUM_13_), 
        .B_12_(add_2_root_r115_SUM_12_), .B_11_(add_2_root_r115_SUM_11_), 
        .B_10_(add_2_root_r115_SUM_10_), .B_9_(add_2_root_r115_SUM_9_), .B_8_(
        add_2_root_r115_SUM_8_), .B_7_(add_2_root_r115_SUM_7_), .B_6_(
        add_2_root_r115_SUM_6_), .B_5_(add_2_root_r115_SUM_5_), .B_4_(
        add_2_root_r115_SUM_4_), .SUM_23_(N221), .SUM_22_(N220), .SUM_21_(N219), .SUM_20_(N218), .SUM_19_(N217), .SUM_18_(N216), .SUM_17_(N215), .SUM_16_(
        N214), .SUM_15_(N213), .SUM_14_(N212), .SUM_13_(N211), .SUM_12_(N210), 
        .SUM_11_(N209), .SUM_10_(N208), .SUM_9_(N207), .SUM_8_(N206), .SUM_7_(
        N205) );
  TLATX1 neg_mul_reg_19_ ( .G(N446), .D(N459), .Q(n1), .QN(n15) );
  TLATX1 neg_mul_reg_18_ ( .G(N446), .D(N458), .QN(n6) );
  TLATX1 neg_mul_reg_17_ ( .G(N446), .D(N457), .QN(n5) );
  TLATX1 neg_mul_reg_16_ ( .G(N446), .D(N456), .QN(n4) );
  TLATX1 neg_mul_reg_15_ ( .G(N446), .D(N455), .QN(n3) );
  TLATX1 neg_mul_reg_11_ ( .G(N446), .D(N451), .Q(neg_mul[11]), .QN(n2) );
  TLATX1 neg_mul_reg_23_ ( .G(N446), .D(N463), .Q(neg_mul[23]), .QN(n17) );
  TLATX1 neg_mul_reg_22_ ( .G(N446), .D(N462), .Q(neg_mul[22]), .QN(n12) );
  TLATX1 neg_mul_reg_21_ ( .G(N446), .D(N461), .Q(neg_mul[21]), .QN(n13) );
  TLATX1 neg_mul_reg_20_ ( .G(N446), .D(N460), .QN(n16) );
  TLATX1 neg_mul_reg_12_ ( .G(N446), .D(N452), .Q(neg_mul[12]), .QN(n8) );
  TLATX1 neg_mul_reg_9_ ( .G(N446), .D(N449), .Q(neg_mul[9]), .QN(n10) );
  TLATX1 neg_mul_reg_14_ ( .G(N446), .D(N454), .Q(neg_mul[14]), .QN(n11) );
  TLATX1 neg_mul_reg_13_ ( .G(N446), .D(N453), .Q(neg_mul[13]), .QN(n9) );
  TLATX1 neg_mul_reg_10_ ( .G(N446), .D(N450), .Q(neg_mul[10]), .QN(n7) );
  TLATX1 neg_mul_reg_8_ ( .G(N446), .D(N448), .Q(neg_mul[8]), .QN(n14) );
  TLATX1 neg_mul_reg_7_ ( .G(N446), .D(N447), .Q(out[0]) );
  CLKINVX3 U2 ( .A(n274), .Y(in_17bit_b[16]) );
  NOR2X2 U3 ( .A(n20), .B(n86), .Y(n88) );
  MXI2X2 U4 ( .A(n16), .B(n32), .S0(n162), .Y(out[13]) );
  OAI21X1 U5 ( .A0(n19), .A1(n58), .B0(n57), .Y(n62) );
  OAI21X1 U6 ( .A0(n19), .A1(n50), .B0(n49), .Y(n55) );
  BUFX12 U7 ( .A(in_8bit[7]), .Y(n19) );
  AOI2BB2X1 U8 ( .B0(n85), .B1(n19), .A0N(n19), .A1N(neg_mul[13]), .Y(n86) );
  NAND2X2 U9 ( .A(n19), .B(n14), .Y(n49) );
  AOI2BB2X1 U10 ( .B0(n93), .B1(n37), .A0N(n18), .A1N(neg_mul[14]), .Y(n94) );
  NOR2X2 U11 ( .A(n161), .B(n31), .Y(n22) );
  NAND2X1 U12 ( .A(n37), .B(n8), .Y(n75) );
  OAI21XL U13 ( .A0(n18), .A1(n65), .B0(n64), .Y(n70) );
  NAND2X1 U14 ( .A(n37), .B(n11), .Y(n91) );
  OAI21XL U15 ( .A0(n19), .A1(n84), .B0(n83), .Y(n89) );
  NAND2X1 U16 ( .A(n18), .B(n9), .Y(n83) );
  INVX4 U17 ( .A(n161), .Y(n162) );
  INVX1 U18 ( .A(n175), .Y(n171) );
  AOI22X1 U19 ( .A0(N27), .A1(n44), .B0(in_17bit[14]), .B1(n21), .Y(n263) );
  INVX1 U20 ( .A(n21), .Y(n44) );
  NOR2X2 U21 ( .A(n20), .B(n94), .Y(n95) );
  CLKINVX8 U22 ( .A(n45), .Y(n20) );
  AOI2BB2X2 U23 ( .B0(n77), .B1(n37), .A0N(n37), .A1N(neg_mul[12]), .Y(n78) );
  AOI2BB2X2 U24 ( .B0(n66), .B1(n37), .A0N(n37), .A1N(neg_mul[10]), .Y(n68) );
  AOI2BB2X2 U25 ( .B0(n59), .B1(n37), .A0N(n37), .A1N(neg_mul[9]), .Y(n60) );
  NOR2X2 U26 ( .A(n46), .B(n78), .Y(n80) );
  XOR2X4 U27 ( .A(n73), .B(neg_mul[11]), .Y(out[4]) );
  BUFX16 U28 ( .A(in_8bit[7]), .Y(n18) );
  NOR2X4 U29 ( .A(n27), .B(n99), .Y(n100) );
  INVXL U30 ( .A(n20), .Y(n21) );
  INVX8 U31 ( .A(in_8bit[7]), .Y(n38) );
  INVX8 U32 ( .A(n38), .Y(n37) );
  INVX8 U33 ( .A(in_17bit[16]), .Y(n45) );
  INVXL U34 ( .A(n44), .Y(n48) );
  NAND2X2 U35 ( .A(n18), .B(n7), .Y(n64) );
  XNOR2X2 U36 ( .A(n20), .B(n19), .Y(n99) );
  XNOR2X4 U37 ( .A(n46), .B(n19), .Y(n97) );
  NOR2X4 U38 ( .A(n161), .B(n29), .Y(n160) );
  NOR2X4 U39 ( .A(n28), .B(n101), .Y(n158) );
  XNOR2X2 U40 ( .A(n46), .B(n19), .Y(n101) );
  XNOR2X4 U41 ( .A(n46), .B(n19), .Y(n161) );
  AOI211X4 U42 ( .A0(n20), .A1(n89), .B0(n88), .C0(n87), .Y(out[6]) );
  INVX8 U43 ( .A(n45), .Y(n46) );
  AOI22XL U44 ( .A0(N18), .A1(n44), .B0(in_17bit[5]), .B1(n21), .Y(n236) );
  NOR2X4 U45 ( .A(n26), .B(n97), .Y(n98) );
  AOI2BB2X4 U46 ( .B0(n51), .B1(n18), .A0N(n18), .A1N(neg_mul[8]), .Y(n53) );
  INVX8 U47 ( .A(n45), .Y(n47) );
  AOI211X4 U48 ( .A0(n46), .A1(n96), .B0(n95), .C0(n26), .Y(out[7]) );
  XNOR2X4 U49 ( .A(n47), .B(n19), .Y(n71) );
  NOR2X4 U50 ( .A(n72), .B(n71), .Y(n73) );
  OAI21XL U51 ( .A0(n18), .A1(n92), .B0(n91), .Y(n96) );
  MX2X1 U52 ( .A(neg_mul[21]), .B(N479), .S0(n162), .Y(out[14]) );
  INVX1 U53 ( .A(n224), .Y(in_17bit_b[1]) );
  INVX1 U54 ( .A(n263), .Y(in_17bit_b[14]) );
  INVX1 U55 ( .A(n260), .Y(in_17bit_b[13]) );
  INVX1 U56 ( .A(n227), .Y(in_17bit_b[2]) );
  INVX1 U57 ( .A(n245), .Y(in_17bit_b[8]) );
  INVX1 U58 ( .A(n239), .Y(in_17bit_b[6]) );
  INVX1 U59 ( .A(n242), .Y(in_17bit_b[7]) );
  INVX1 U60 ( .A(n248), .Y(in_17bit_b[9]) );
  INVX1 U61 ( .A(n251), .Y(in_17bit_b[10]) );
  INVX1 U62 ( .A(n254), .Y(in_17bit_b[11]) );
  INVX1 U63 ( .A(n257), .Y(in_17bit_b[12]) );
  INVX1 U64 ( .A(n233), .Y(in_17bit_b[4]) );
  INVX1 U65 ( .A(n236), .Y(in_17bit_b[5]) );
  INVX1 U66 ( .A(n230), .Y(in_17bit_b[3]) );
  NAND2X2 U67 ( .A(n37), .B(n10), .Y(n57) );
  OAI21X4 U68 ( .A0(n47), .A1(n60), .B0(n63), .Y(n61) );
  XOR2X4 U69 ( .A(n22), .B(n1), .Y(out[12]) );
  AOI21X1 U70 ( .A0(n23), .A1(n24), .B0(n267), .Y(n220) );
  NOR4XL U71 ( .A(in_8bit[4]), .B(in_8bit[5]), .C(in_8bit[6]), .D(n19), .Y(n23) );
  NOR4X1 U72 ( .A(n36), .B(in_8bit[0]), .C(n42), .D(in_8bit[3]), .Y(n24) );
  AND4X1 U73 ( .A(n36), .B(n19), .C(n214), .D(n39), .Y(n25) );
  INVX1 U74 ( .A(n43), .Y(n42) );
  NOR3X1 U75 ( .A(n43), .B(n41), .C(n39), .Y(n219) );
  NOR4BX1 U76 ( .AN(n217), .B(n39), .C(n36), .D(n42), .Y(n218) );
  NOR2X1 U77 ( .A(in_8bit[6]), .B(in_8bit[3]), .Y(n217) );
  NAND3X1 U78 ( .A(n42), .B(n41), .C(in_8bit[5]), .Y(n215) );
  ADDFX2 U79 ( .A(in_17bit_b[16]), .B(in_17bit_b[12]), .CI(
        add_1_root_r112_carry_16_), .CO(add_1_root_r112_carry_17_), .S(
        add_1_root_r112_SUM_16_) );
  ADDFX2 U80 ( .A(add_1_root_r119_A_19_), .B(in_17bit_b[13]), .CI(
        add_1_root_r119_carry[19]), .CO(add_1_root_r119_carry[20]), .S(
        add_1_root_r119_SUM_19_) );
  ADDFX2 U81 ( .A(in_17bit_b[16]), .B(in_17bit_b[15]), .CI(
        add_3_root_r119_carry_17_), .CO(add_3_root_r119_carry_18_), .S(
        add_1_root_r119_A_17_) );
  ADDFX2 U82 ( .A(in_17bit_b[16]), .B(in_17bit_b[14]), .CI(
        add_2_root_r115_carry_17_), .CO(add_2_root_r115_carry_18_), .S(
        add_2_root_r115_SUM_17_) );
  ADDFX2 U83 ( .A(in_17bit_b[16]), .B(in_17bit_b[14]), .CI(
        add_1_root_r115_carry_20_), .CO(add_1_root_r115_carry_21_), .S(
        add_1_root_r115_SUM_20_) );
  ADDFX2 U84 ( .A(in_17bit_b[16]), .B(in_17bit_b[15]), .CI(
        add_2_root_r119_carry_20_), .CO(add_2_root_r119_carry_21_), .S(
        add_2_root_r119_SUM_20_) );
  ADDFX2 U85 ( .A(in_17bit_b[3]), .B(in_17bit_b[1]), .CI(
        add_2_root_r115_carry_4_), .CO(add_2_root_r115_carry_5_), .S(
        add_2_root_r115_SUM_4_) );
  ADDFX2 U86 ( .A(in_17bit_b[4]), .B(in_17bit_b[2]), .CI(
        add_2_root_r115_carry_5_), .CO(add_2_root_r115_carry_6_), .S(
        add_2_root_r115_SUM_5_) );
  ADDFX2 U87 ( .A(in_17bit_b[5]), .B(in_17bit_b[1]), .CI(
        add_1_root_r112_carry_5_), .CO(add_1_root_r112_carry_6_), .S(
        add_1_root_r112_SUM_5_) );
  ADDFX2 U88 ( .A(in_17bit_b[6]), .B(in_17bit_b[5]), .CI(
        add_3_root_r119_carry_7_), .CO(add_3_root_r119_carry_8_), .S(
        add_1_root_r119_A_7_) );
  ADDFX2 U89 ( .A(in_17bit_b[6]), .B(in_17bit_b[2]), .CI(
        add_1_root_r112_carry_6_), .CO(add_1_root_r112_carry_7_), .S(
        add_1_root_r112_SUM_6_) );
  ADDFX2 U90 ( .A(in_17bit_b[3]), .B(in_17bit_b[1]), .CI(
        add_2_root_r115_carry_4_), .CO(add_1_root_r115_carry_8_), .S(
        add_1_root_r115_SUM_7_) );
  ADDFX2 U91 ( .A(in_17bit_b[7]), .B(in_17bit_b[6]), .CI(
        add_3_root_r119_carry_8_), .CO(add_3_root_r119_carry_9_), .S(
        add_1_root_r119_A_8_) );
  ADDFX2 U92 ( .A(add_1_root_r119_A_7_), .B(in_17bit_b[1]), .CI(
        add_1_root_r119_carry[7]), .CO(add_1_root_r119_carry[8]), .S(
        add_1_root_r119_SUM_7_) );
  ADDFX2 U93 ( .A(in_17bit_b[2]), .B(in_17bit_b[1]), .CI(
        add_3_root_r119_carry_3_), .CO(add_2_root_r119_carry_7_), .S(
        add_2_root_r119_SUM_6_) );
  ADDFX2 U94 ( .A(in_17bit_b[4]), .B(in_17bit_b[2]), .CI(
        add_1_root_r115_carry_8_), .CO(add_1_root_r115_carry_9_), .S(
        add_1_root_r115_SUM_8_) );
  ADDFX2 U95 ( .A(in_17bit_b[8]), .B(in_17bit_b[7]), .CI(
        add_3_root_r119_carry_9_), .CO(add_3_root_r119_carry_10_), .S(
        add_1_root_r119_A_9_) );
  ADDFX2 U96 ( .A(add_1_root_r119_A_8_), .B(in_17bit_b[2]), .CI(
        add_1_root_r119_carry[8]), .CO(add_1_root_r119_carry[9]), .S(
        add_1_root_r119_SUM_8_) );
  ADDFX2 U97 ( .A(in_17bit_b[3]), .B(in_17bit_b[2]), .CI(
        add_2_root_r119_carry_7_), .CO(add_2_root_r119_carry_8_), .S(
        add_2_root_r119_SUM_7_) );
  ADDFX2 U98 ( .A(in_17bit_b[6]), .B(in_17bit_b[4]), .CI(
        add_2_root_r115_carry_7_), .CO(add_2_root_r115_carry_8_), .S(
        add_2_root_r115_SUM_7_) );
  ADDFX2 U99 ( .A(in_17bit_b[9]), .B(in_17bit_b[8]), .CI(
        add_3_root_r119_carry_10_), .CO(add_3_root_r119_carry_11_), .S(
        add_1_root_r119_A_10_) );
  ADDFX2 U100 ( .A(in_17bit_b[7]), .B(in_17bit_b[5]), .CI(
        add_2_root_r115_carry_8_), .CO(add_2_root_r115_carry_9_), .S(
        add_2_root_r115_SUM_8_) );
  ADDFX2 U101 ( .A(in_17bit_b[9]), .B(in_17bit_b[5]), .CI(
        add_1_root_r112_carry_9_), .CO(add_1_root_r112_carry_10_), .S(
        add_1_root_r112_SUM_9_) );
  ADDFX2 U102 ( .A(in_17bit_b[6]), .B(in_17bit_b[4]), .CI(
        add_1_root_r115_carry_10_), .CO(add_1_root_r115_carry_11_), .S(
        add_1_root_r115_SUM_10_) );
  ADDFX2 U103 ( .A(in_17bit_b[10]), .B(in_17bit_b[9]), .CI(
        add_3_root_r119_carry_11_), .CO(add_3_root_r119_carry_12_), .S(
        add_1_root_r119_A_11_) );
  ADDFX2 U104 ( .A(add_1_root_r119_A_10_), .B(in_17bit_b[4]), .CI(
        add_1_root_r119_carry[10]), .CO(add_1_root_r119_carry[11]), .S(
        add_1_root_r119_SUM_10_) );
  ADDFX2 U105 ( .A(in_17bit_b[8]), .B(in_17bit_b[4]), .CI(
        add_1_root_r112_carry_8_), .CO(add_1_root_r112_carry_9_), .S(
        add_1_root_r112_SUM_8_) );
  ADDFX2 U106 ( .A(in_17bit_b[5]), .B(in_17bit_b[4]), .CI(
        add_2_root_r119_carry_9_), .CO(add_2_root_r119_carry_10_), .S(
        add_2_root_r119_SUM_9_) );
  ADDFX2 U107 ( .A(in_17bit_b[8]), .B(in_17bit_b[6]), .CI(
        add_2_root_r115_carry_9_), .CO(add_2_root_r115_carry_10_), .S(
        add_2_root_r115_SUM_9_) );
  ADDFX2 U108 ( .A(in_17bit_b[10]), .B(in_17bit_b[6]), .CI(
        add_1_root_r112_carry_10_), .CO(add_1_root_r112_carry_11_), .S(
        add_1_root_r112_SUM_10_) );
  ADDFX2 U109 ( .A(in_17bit_b[7]), .B(in_17bit_b[5]), .CI(
        add_1_root_r115_carry_11_), .CO(add_1_root_r115_carry_12_), .S(
        add_1_root_r115_SUM_11_) );
  ADDFX2 U110 ( .A(in_17bit_b[11]), .B(in_17bit_b[10]), .CI(
        add_3_root_r119_carry_12_), .CO(add_3_root_r119_carry_13_), .S(
        add_1_root_r119_A_12_) );
  ADDFX2 U111 ( .A(add_1_root_r119_A_11_), .B(in_17bit_b[5]), .CI(
        add_1_root_r119_carry[11]), .CO(add_1_root_r119_carry[12]), .S(
        add_1_root_r119_SUM_11_) );
  ADDFX2 U112 ( .A(in_17bit_b[6]), .B(in_17bit_b[5]), .CI(
        add_2_root_r119_carry_10_), .CO(add_2_root_r119_carry_11_), .S(
        add_2_root_r119_SUM_10_) );
  ADDFX2 U113 ( .A(in_17bit_b[9]), .B(in_17bit_b[7]), .CI(
        add_2_root_r115_carry_10_), .CO(add_2_root_r115_carry_11_), .S(
        add_2_root_r115_SUM_10_) );
  ADDFX2 U114 ( .A(in_17bit_b[11]), .B(in_17bit_b[7]), .CI(
        add_1_root_r112_carry_11_), .CO(add_1_root_r112_carry_12_), .S(
        add_1_root_r112_SUM_11_) );
  ADDFX2 U115 ( .A(in_17bit_b[8]), .B(in_17bit_b[6]), .CI(
        add_1_root_r115_carry_12_), .CO(add_1_root_r115_carry_13_), .S(
        add_1_root_r115_SUM_12_) );
  ADDFX2 U116 ( .A(in_17bit_b[12]), .B(in_17bit_b[11]), .CI(
        add_3_root_r119_carry_13_), .CO(add_3_root_r119_carry_14_), .S(
        add_1_root_r119_A_13_) );
  ADDFX2 U117 ( .A(add_1_root_r119_A_12_), .B(in_17bit_b[6]), .CI(
        add_1_root_r119_carry[12]), .CO(add_1_root_r119_carry[13]), .S(
        add_1_root_r119_SUM_12_) );
  ADDFX2 U118 ( .A(in_17bit_b[7]), .B(in_17bit_b[6]), .CI(
        add_2_root_r119_carry_11_), .CO(add_2_root_r119_carry_12_), .S(
        add_2_root_r119_SUM_11_) );
  ADDFX2 U119 ( .A(in_17bit_b[10]), .B(in_17bit_b[8]), .CI(
        add_2_root_r115_carry_11_), .CO(add_2_root_r115_carry_12_), .S(
        add_2_root_r115_SUM_11_) );
  ADDFX2 U120 ( .A(in_17bit_b[12]), .B(in_17bit_b[8]), .CI(
        add_1_root_r112_carry_12_), .CO(add_1_root_r112_carry_13_), .S(
        add_1_root_r112_SUM_12_) );
  ADDFX2 U121 ( .A(in_17bit_b[9]), .B(in_17bit_b[7]), .CI(
        add_1_root_r115_carry_13_), .CO(add_1_root_r115_carry_14_), .S(
        add_1_root_r115_SUM_13_) );
  ADDFX2 U122 ( .A(in_17bit_b[13]), .B(in_17bit_b[12]), .CI(
        add_3_root_r119_carry_14_), .CO(add_3_root_r119_carry_15_), .S(
        add_1_root_r119_A_14_) );
  ADDFX2 U123 ( .A(in_17bit_b[8]), .B(in_17bit_b[7]), .CI(
        add_2_root_r119_carry_12_), .CO(add_2_root_r119_carry_13_), .S(
        add_2_root_r119_SUM_12_) );
  ADDFX2 U124 ( .A(in_17bit_b[11]), .B(in_17bit_b[9]), .CI(
        add_2_root_r115_carry_12_), .CO(add_2_root_r115_carry_13_), .S(
        add_2_root_r115_SUM_12_) );
  ADDFX2 U125 ( .A(in_17bit_b[13]), .B(in_17bit_b[9]), .CI(
        add_1_root_r112_carry_13_), .CO(add_1_root_r112_carry_14_), .S(
        add_1_root_r112_SUM_13_) );
  ADDFX2 U126 ( .A(in_17bit_b[10]), .B(in_17bit_b[8]), .CI(
        add_1_root_r115_carry_14_), .CO(add_1_root_r115_carry_15_), .S(
        add_1_root_r115_SUM_14_) );
  ADDFX2 U127 ( .A(in_17bit_b[14]), .B(in_17bit_b[13]), .CI(
        add_3_root_r119_carry_15_), .CO(add_3_root_r119_carry_16_), .S(
        add_1_root_r119_A_15_) );
  ADDFX2 U128 ( .A(add_1_root_r119_A_14_), .B(in_17bit_b[8]), .CI(
        add_1_root_r119_carry[14]), .CO(add_1_root_r119_carry[15]), .S(
        add_1_root_r119_SUM_14_) );
  ADDFX2 U129 ( .A(in_17bit_b[9]), .B(in_17bit_b[8]), .CI(
        add_2_root_r119_carry_13_), .CO(add_2_root_r119_carry_14_), .S(
        add_2_root_r119_SUM_13_) );
  ADDFX2 U130 ( .A(in_17bit_b[12]), .B(in_17bit_b[10]), .CI(
        add_2_root_r115_carry_13_), .CO(add_2_root_r115_carry_14_), .S(
        add_2_root_r115_SUM_13_) );
  ADDFX2 U131 ( .A(in_17bit_b[14]), .B(in_17bit_b[10]), .CI(
        add_1_root_r112_carry_14_), .CO(add_1_root_r112_carry_15_), .S(
        add_1_root_r112_SUM_14_) );
  ADDFX2 U132 ( .A(in_17bit_b[11]), .B(in_17bit_b[9]), .CI(
        add_1_root_r115_carry_15_), .CO(add_1_root_r115_carry_16_), .S(
        add_1_root_r115_SUM_15_) );
  ADDFX2 U133 ( .A(add_1_root_r119_A_15_), .B(in_17bit_b[9]), .CI(
        add_1_root_r119_carry[15]), .CO(add_1_root_r119_carry[16]), .S(
        add_1_root_r119_SUM_15_) );
  ADDFX2 U134 ( .A(in_17bit_b[3]), .B(in_17bit_b[2]), .CI(
        add_3_root_r119_carry_4_), .CO(add_3_root_r119_carry_5_), .S(
        add_1_root_r119_A_4_) );
  ADDFX2 U135 ( .A(in_17bit_b[2]), .B(in_17bit_b[1]), .CI(
        add_3_root_r119_carry_3_), .CO(add_3_root_r119_carry_4_), .S(
        add_1_root_r119_A_3_) );
  ADDFX2 U136 ( .A(in_17bit_b[10]), .B(in_17bit_b[9]), .CI(
        add_2_root_r119_carry_14_), .CO(add_2_root_r119_carry_15_), .S(
        add_2_root_r119_SUM_14_) );
  ADDFX2 U137 ( .A(in_17bit_b[13]), .B(in_17bit_b[11]), .CI(
        add_2_root_r115_carry_14_), .CO(add_2_root_r115_carry_15_), .S(
        add_2_root_r115_SUM_14_) );
  ADDFX2 U138 ( .A(in_17bit_b[15]), .B(in_17bit_b[11]), .CI(
        add_1_root_r112_carry_15_), .CO(add_1_root_r112_carry_16_), .S(
        add_1_root_r112_SUM_15_) );
  ADDFX2 U139 ( .A(in_17bit_b[12]), .B(in_17bit_b[10]), .CI(
        add_1_root_r115_carry_16_), .CO(add_1_root_r115_carry_17_), .S(
        add_1_root_r115_SUM_16_) );
  ADDFX2 U140 ( .A(add_1_root_r119_A_16_), .B(in_17bit_b[10]), .CI(
        add_1_root_r119_carry[16]), .CO(add_1_root_r119_carry[17]), .S(
        add_1_root_r119_SUM_16_) );
  ADDFX2 U141 ( .A(in_17bit_b[11]), .B(in_17bit_b[10]), .CI(
        add_2_root_r119_carry_15_), .CO(add_2_root_r119_carry_16_), .S(
        add_2_root_r119_SUM_15_) );
  ADDFX2 U142 ( .A(in_17bit_b[14]), .B(in_17bit_b[12]), .CI(
        add_2_root_r115_carry_15_), .CO(add_2_root_r115_carry_16_), .S(
        add_2_root_r115_SUM_15_) );
  ADDFX2 U143 ( .A(in_17bit_b[13]), .B(in_17bit_b[11]), .CI(
        add_1_root_r115_carry_17_), .CO(add_1_root_r115_carry_18_), .S(
        add_1_root_r115_SUM_17_) );
  ADDFX2 U144 ( .A(add_1_root_r119_A_17_), .B(in_17bit_b[11]), .CI(
        add_1_root_r119_carry[17]), .CO(add_1_root_r119_carry[18]), .S(
        add_1_root_r119_SUM_17_) );
  ADDFX2 U145 ( .A(in_17bit_b[12]), .B(in_17bit_b[11]), .CI(
        add_2_root_r119_carry_16_), .CO(add_2_root_r119_carry_17_), .S(
        add_2_root_r119_SUM_16_) );
  ADDFX2 U146 ( .A(in_17bit_b[15]), .B(in_17bit_b[13]), .CI(
        add_2_root_r115_carry_16_), .CO(add_2_root_r115_carry_17_), .S(
        add_2_root_r115_SUM_16_) );
  ADDFX2 U147 ( .A(in_17bit_b[14]), .B(in_17bit_b[12]), .CI(
        add_1_root_r115_carry_18_), .CO(add_1_root_r115_carry_19_), .S(
        add_1_root_r115_SUM_18_) );
  ADDFX2 U148 ( .A(add_1_root_r119_A_18_), .B(in_17bit_b[12]), .CI(
        add_1_root_r119_carry[18]), .CO(add_1_root_r119_carry[19]), .S(
        add_1_root_r119_SUM_18_) );
  ADDFX2 U149 ( .A(in_17bit_b[13]), .B(in_17bit_b[12]), .CI(
        add_2_root_r119_carry_17_), .CO(add_2_root_r119_carry_18_), .S(
        add_2_root_r119_SUM_17_) );
  ADDFX2 U150 ( .A(in_17bit_b[14]), .B(in_17bit_b[13]), .CI(
        add_2_root_r119_carry_18_), .CO(add_2_root_r119_carry_19_), .S(
        add_2_root_r119_SUM_18_) );
  ADDFX2 U151 ( .A(in_17bit_b[5]), .B(in_17bit_b[3]), .CI(
        add_2_root_r115_carry_6_), .CO(add_2_root_r115_carry_7_), .S(
        add_2_root_r115_SUM_6_) );
  ADDFX2 U152 ( .A(in_17bit_b[7]), .B(in_17bit_b[3]), .CI(
        add_1_root_r112_carry_7_), .CO(add_1_root_r112_carry_8_), .S(
        add_1_root_r112_SUM_7_) );
  ADDFX2 U153 ( .A(in_17bit_b[5]), .B(in_17bit_b[3]), .CI(
        add_1_root_r115_carry_9_), .CO(add_1_root_r115_carry_10_), .S(
        add_1_root_r115_SUM_9_) );
  ADDFX2 U154 ( .A(in_17bit_b[4]), .B(in_17bit_b[3]), .CI(
        add_2_root_r119_carry_8_), .CO(add_2_root_r119_carry_9_), .S(
        add_2_root_r119_SUM_8_) );
  ADDFX2 U155 ( .A(add_1_root_r119_A_13_), .B(in_17bit_b[7]), .CI(
        add_1_root_r119_carry[13]), .CO(add_1_root_r119_carry[14]), .S(
        add_1_root_r119_SUM_13_) );
  ADDFX2 U156 ( .A(in_17bit_b[15]), .B(in_17bit_b[14]), .CI(
        add_3_root_r119_carry_16_), .CO(add_3_root_r119_carry_17_), .S(
        add_1_root_r119_A_16_) );
  ADDFX2 U157 ( .A(in_17bit_b[4]), .B(in_17bit_b[3]), .CI(
        add_3_root_r119_carry_5_), .CO(add_3_root_r119_carry_6_), .S(
        add_1_root_r119_A_5_) );
  ADDFX2 U158 ( .A(in_17bit_b[15]), .B(in_17bit_b[13]), .CI(
        add_1_root_r115_carry_19_), .CO(add_1_root_r115_carry_20_), .S(
        add_1_root_r115_SUM_19_) );
  ADDFX2 U159 ( .A(in_17bit_b[5]), .B(in_17bit_b[4]), .CI(
        add_3_root_r119_carry_6_), .CO(add_3_root_r119_carry_7_), .S(
        add_1_root_r119_A_6_) );
  ADDFX2 U160 ( .A(add_1_root_r119_A_9_), .B(in_17bit_b[3]), .CI(
        add_1_root_r119_carry[9]), .CO(add_1_root_r119_carry[10]), .S(
        add_1_root_r119_SUM_9_) );
  ADDFX2 U161 ( .A(in_17bit_b[15]), .B(in_17bit_b[14]), .CI(
        add_2_root_r119_carry_19_), .CO(add_2_root_r119_carry_20_), .S(
        add_2_root_r119_SUM_19_) );
  INVX1 U162 ( .A(n216), .Y(n174) );
  NAND3BX1 U163 ( .AN(in_8bit[5]), .B(n43), .C(in_8bit[3]), .Y(n216) );
  INVX1 U164 ( .A(in_8bit[6]), .Y(n40) );
  CLKINVX3 U165 ( .A(n221), .Y(in_17bit_b[0]) );
  INVX1 U166 ( .A(n194), .Y(n273) );
  NAND2XL U167 ( .A(N29), .B(n44), .Y(n274) );
  INVX1 U168 ( .A(n67), .Y(n72) );
  OAI21XL U169 ( .A0(n273), .A1(n274), .B0(n272), .Y(N463) );
  AOI22X1 U170 ( .A0(N221), .A1(n35), .B0(N363), .B1(n34), .Y(n272) );
  INVX1 U171 ( .A(n90), .Y(n87) );
  CLKINVX3 U172 ( .A(n266), .Y(in_17bit_b[15]) );
  INVX1 U173 ( .A(n82), .Y(n79) );
  NAND2X1 U174 ( .A(n223), .B(n222), .Y(N447) );
  AOI22X1 U175 ( .A0(N108), .A1(n267), .B0(N205), .B1(n35), .Y(n222) );
  AOI22X1 U176 ( .A0(N347), .A1(n34), .B0(n194), .B1(in_17bit_b[0]), .Y(n223)
         );
  NAND2X1 U177 ( .A(n226), .B(n225), .Y(N448) );
  AOI22X1 U178 ( .A0(N109), .A1(n267), .B0(N206), .B1(n35), .Y(n225) );
  AOI22X1 U179 ( .A0(N348), .A1(n34), .B0(n194), .B1(in_17bit_b[1]), .Y(n226)
         );
  NAND2X1 U180 ( .A(n229), .B(n228), .Y(N449) );
  AOI22X1 U181 ( .A0(N110), .A1(n267), .B0(N207), .B1(n35), .Y(n228) );
  AOI22X1 U182 ( .A0(N349), .A1(n34), .B0(n194), .B1(in_17bit_b[2]), .Y(n229)
         );
  NAND2X1 U183 ( .A(n232), .B(n231), .Y(N450) );
  AOI22X1 U184 ( .A0(N111), .A1(n267), .B0(N208), .B1(n35), .Y(n231) );
  AOI22X1 U185 ( .A0(N350), .A1(n34), .B0(n194), .B1(in_17bit_b[3]), .Y(n232)
         );
  NAND2X1 U186 ( .A(n235), .B(n234), .Y(N451) );
  AOI22X1 U187 ( .A0(N112), .A1(n267), .B0(N209), .B1(n35), .Y(n234) );
  AOI22X1 U188 ( .A0(N351), .A1(n34), .B0(n194), .B1(in_17bit_b[4]), .Y(n235)
         );
  NAND2X1 U189 ( .A(n238), .B(n237), .Y(N452) );
  AOI22X1 U190 ( .A0(N113), .A1(n267), .B0(N210), .B1(n35), .Y(n237) );
  AOI22X1 U191 ( .A0(N352), .A1(n34), .B0(n194), .B1(in_17bit_b[5]), .Y(n238)
         );
  NAND2X1 U192 ( .A(n241), .B(n240), .Y(N453) );
  AOI22X1 U193 ( .A0(N114), .A1(n267), .B0(N211), .B1(n35), .Y(n240) );
  AOI22X1 U194 ( .A0(N353), .A1(n34), .B0(n194), .B1(in_17bit_b[6]), .Y(n241)
         );
  NAND2X1 U195 ( .A(n244), .B(n243), .Y(N454) );
  AOI22X1 U196 ( .A0(N115), .A1(n267), .B0(N212), .B1(n35), .Y(n243) );
  AOI22X1 U197 ( .A0(N354), .A1(n34), .B0(n194), .B1(in_17bit_b[7]), .Y(n244)
         );
  NAND2X1 U198 ( .A(n247), .B(n246), .Y(N455) );
  AOI22X1 U199 ( .A0(N116), .A1(n267), .B0(N213), .B1(n35), .Y(n246) );
  AOI22X1 U200 ( .A0(N355), .A1(n34), .B0(n194), .B1(in_17bit_b[8]), .Y(n247)
         );
  NAND2X1 U201 ( .A(n250), .B(n249), .Y(N456) );
  AOI22X1 U202 ( .A0(N117), .A1(n267), .B0(N214), .B1(n35), .Y(n249) );
  AOI22X1 U203 ( .A0(N356), .A1(n34), .B0(n194), .B1(in_17bit_b[9]), .Y(n250)
         );
  NAND2X1 U204 ( .A(n253), .B(n252), .Y(N457) );
  AOI22X1 U205 ( .A0(N118), .A1(n267), .B0(N215), .B1(n35), .Y(n252) );
  AOI22X1 U206 ( .A0(N357), .A1(n34), .B0(n194), .B1(in_17bit_b[10]), .Y(n253)
         );
  NAND2X1 U207 ( .A(n256), .B(n255), .Y(N458) );
  AOI22X1 U208 ( .A0(N119), .A1(n267), .B0(N216), .B1(n35), .Y(n255) );
  AOI22X1 U209 ( .A0(N358), .A1(n34), .B0(n194), .B1(in_17bit_b[11]), .Y(n256)
         );
  NAND2X1 U210 ( .A(n259), .B(n258), .Y(N459) );
  AOI22X1 U211 ( .A0(N120), .A1(n267), .B0(N217), .B1(n35), .Y(n258) );
  AOI22X1 U212 ( .A0(N359), .A1(n34), .B0(n194), .B1(in_17bit_b[12]), .Y(n259)
         );
  NAND2X1 U213 ( .A(n262), .B(n261), .Y(N460) );
  AOI22X1 U214 ( .A0(N121), .A1(n267), .B0(N218), .B1(n35), .Y(n261) );
  AOI22X1 U215 ( .A0(N360), .A1(n34), .B0(n194), .B1(in_17bit_b[13]), .Y(n262)
         );
  NAND2X1 U216 ( .A(n265), .B(n264), .Y(N461) );
  AOI22X1 U217 ( .A0(N122), .A1(n267), .B0(N219), .B1(n35), .Y(n264) );
  AOI22X1 U218 ( .A0(N361), .A1(n34), .B0(n194), .B1(in_17bit_b[14]), .Y(n265)
         );
  NAND2X1 U219 ( .A(n269), .B(n268), .Y(N462) );
  AOI22X1 U220 ( .A0(N123), .A1(n267), .B0(N220), .B1(n35), .Y(n268) );
  AOI22X1 U221 ( .A0(N362), .A1(n34), .B0(n194), .B1(in_17bit_b[15]), .Y(n269)
         );
  CLKBUFXL U222 ( .A(in_8bit[1]), .Y(n36) );
  INVX1 U223 ( .A(in_8bit[0]), .Y(n39) );
  INVX1 U224 ( .A(in_8bit[3]), .Y(n41) );
  OAI21XL U225 ( .A0(n18), .A1(n76), .B0(n75), .Y(n81) );
  AOI22XL U226 ( .A0(in_17bit[0]), .A1(n44), .B0(in_17bit[0]), .B1(n48), .Y(
        n221) );
  AOI22XL U227 ( .A0(N26), .A1(n44), .B0(in_17bit[13]), .B1(n21), .Y(n260) );
  AOI22XL U228 ( .A0(N28), .A1(n44), .B0(in_17bit[15]), .B1(n48), .Y(n266) );
  AOI22XL U229 ( .A0(N14), .A1(n44), .B0(in_17bit[1]), .B1(n48), .Y(n224) );
  AOI22XL U230 ( .A0(N15), .A1(n44), .B0(in_17bit[2]), .B1(n48), .Y(n227) );
  AOI22XL U231 ( .A0(N16), .A1(n44), .B0(in_17bit[3]), .B1(n48), .Y(n230) );
  AOI22XL U232 ( .A0(N17), .A1(n44), .B0(in_17bit[4]), .B1(n21), .Y(n233) );
  AOI22XL U233 ( .A0(N20), .A1(n44), .B0(in_17bit[7]), .B1(n48), .Y(n242) );
  AOI22XL U234 ( .A0(N21), .A1(n44), .B0(in_17bit[8]), .B1(n48), .Y(n245) );
  AOI22XL U235 ( .A0(N22), .A1(n44), .B0(in_17bit[9]), .B1(n21), .Y(n248) );
  AOI22XL U236 ( .A0(N23), .A1(n44), .B0(in_17bit[10]), .B1(n21), .Y(n251) );
  AOI22XL U237 ( .A0(N24), .A1(n44), .B0(in_17bit[11]), .B1(n48), .Y(n254) );
  AOI22XL U238 ( .A0(N25), .A1(n44), .B0(in_17bit[12]), .B1(n48), .Y(n257) );
  AOI22XL U239 ( .A0(N19), .A1(n44), .B0(in_17bit[6]), .B1(n21), .Y(n239) );
  AND2X2 U240 ( .A(n87), .B(n11), .Y(n26) );
  NAND2X1 U241 ( .A(n56), .B(n10), .Y(n63) );
  AND2X2 U242 ( .A(n26), .B(n3), .Y(n27) );
  AND2X2 U243 ( .A(n27), .B(n4), .Y(n28) );
  AND2X2 U244 ( .A(n28), .B(n5), .Y(n29) );
  BUFX3 U245 ( .A(n270), .Y(n34) );
  OAI2BB1X1 U246 ( .A0N(n174), .A1N(n25), .B0(n172), .Y(n270) );
  NAND2BX1 U247 ( .AN(n215), .B(n30), .Y(n172) );
  BUFX3 U248 ( .A(n271), .Y(n35) );
  OAI2BB1X1 U249 ( .A0N(n30), .A1N(n174), .B0(n173), .Y(n271) );
  NAND2BX1 U250 ( .AN(n215), .B(n25), .Y(n173) );
  NAND2X1 U251 ( .A(n170), .B(n168), .Y(n267) );
  NAND3X1 U252 ( .A(n218), .B(in_8bit[5]), .C(n164), .Y(n168) );
  NAND4BXL U253 ( .AN(n40), .B(n219), .C(n177), .D(n36), .Y(n170) );
  NAND2BX1 U254 ( .AN(n63), .B(n7), .Y(n67) );
  INVX1 U255 ( .A(n52), .Y(n56) );
  NAND2X1 U256 ( .A(n72), .B(n2), .Y(n74) );
  NAND2X1 U257 ( .A(n79), .B(n9), .Y(n90) );
  OAI2BB1X1 U258 ( .A0N(n218), .A1N(n177), .B0(n176), .Y(n194) );
  NAND3BX1 U259 ( .AN(n175), .B(n219), .C(in_8bit[5]), .Y(n176) );
  NAND2BX1 U260 ( .AN(n74), .B(n8), .Y(n82) );
  AND2X2 U261 ( .A(n171), .B(n39), .Y(n30) );
  AND2X2 U262 ( .A(n29), .B(n6), .Y(n31) );
  INVX1 U263 ( .A(in_17bit[0]), .Y(n178) );
  INVX1 U264 ( .A(in_17bit[1]), .Y(n179) );
  INVX1 U265 ( .A(in_17bit[2]), .Y(n180) );
  INVX1 U266 ( .A(in_17bit[3]), .Y(n181) );
  INVX1 U267 ( .A(in_17bit[6]), .Y(n184) );
  INVX1 U268 ( .A(in_17bit[7]), .Y(n185) );
  INVX1 U269 ( .A(in_17bit[8]), .Y(n186) );
  INVX1 U270 ( .A(in_17bit[9]), .Y(n187) );
  INVX1 U271 ( .A(in_17bit[10]), .Y(n188) );
  INVX1 U272 ( .A(in_17bit[11]), .Y(n189) );
  INVX1 U273 ( .A(in_17bit[12]), .Y(n190) );
  INVX1 U274 ( .A(in_17bit[13]), .Y(n191) );
  INVX1 U275 ( .A(in_17bit[14]), .Y(n192) );
  INVX1 U276 ( .A(in_17bit[15]), .Y(n193) );
  INVX1 U277 ( .A(in_17bit[5]), .Y(n183) );
  INVX1 U278 ( .A(in_17bit[4]), .Y(n182) );
  XNOR2X1 U279 ( .A(n16), .B(sub_add_75_b0_carry[13]), .Y(n32) );
  INVX1 U280 ( .A(n76), .Y(n77) );
  INVX1 U281 ( .A(n50), .Y(n51) );
  INVX1 U282 ( .A(n84), .Y(n85) );
  INVX1 U283 ( .A(n65), .Y(n66) );
  INVX1 U284 ( .A(n58), .Y(n59) );
  INVX1 U285 ( .A(n92), .Y(n93) );
  MX2X1 U286 ( .A(neg_mul[22]), .B(N480), .S0(n162), .Y(out[15]) );
  MX2X1 U287 ( .A(neg_mul[23]), .B(N481), .S0(n162), .Y(out[16]) );
  NAND4BBX1 U288 ( .AN(n34), .BN(n35), .C(n220), .D(n273), .Y(N446) );
  NOR3BXL U289 ( .AN(n19), .B(in_8bit[5]), .C(in_8bit[4]), .Y(n177) );
  NAND4BXL U290 ( .AN(n19), .B(in_8bit[4]), .C(n36), .D(in_8bit[6]), .Y(n175)
         );
  NAND2BX1 U291 ( .AN(n56), .B(neg_mul[9]), .Y(n58) );
  NAND2X1 U292 ( .A(neg_mul[10]), .B(n63), .Y(n65) );
  NAND2X1 U293 ( .A(out[0]), .B(neg_mul[8]), .Y(n50) );
  NOR2X1 U294 ( .A(in_8bit[6]), .B(in_8bit[4]), .Y(n214) );
  NAND2X1 U295 ( .A(neg_mul[12]), .B(n74), .Y(n76) );
  NAND2X1 U296 ( .A(neg_mul[14]), .B(n90), .Y(n92) );
  NAND2X1 U297 ( .A(neg_mul[13]), .B(n82), .Y(n84) );
  NOR2XL U298 ( .A(n19), .B(n163), .Y(n164) );
  INVX1 U299 ( .A(in_8bit[4]), .Y(n163) );
  OR2X2 U300 ( .A(out[0]), .B(neg_mul[8]), .Y(n52) );
  AOI211X4 U301 ( .A0(n20), .A1(n81), .B0(n80), .C0(n79), .Y(out[5]) );
  INVXL U302 ( .A(in_8bit[2]), .Y(n43) );
  OAI21X4 U303 ( .A0(n53), .A1(n47), .B0(n52), .Y(n54) );
  AOI21X4 U304 ( .A0(n46), .A1(n55), .B0(n54), .Y(out[1]) );
  AOI21X4 U305 ( .A0(n20), .A1(n62), .B0(n61), .Y(out[2]) );
  OAI21X4 U306 ( .A0(n47), .A1(n68), .B0(n67), .Y(n69) );
  AOI21X4 U307 ( .A0(n70), .A1(n46), .B0(n69), .Y(out[3]) );
  XNOR2X4 U308 ( .A(n98), .B(n3), .Y(out[8]) );
  XNOR2X4 U309 ( .A(n100), .B(n4), .Y(out[9]) );
  XNOR2X4 U310 ( .A(n158), .B(n5), .Y(out[10]) );
  XNOR2X4 U311 ( .A(n160), .B(n6), .Y(out[11]) );
  AND2X1 U312 ( .A(add_1_root_r112_carry_20_), .B(in_17bit_b[16]), .Y(
        add_1_root_r112_SUM_21_) );
  XOR2X1 U313 ( .A(in_17bit_b[16]), .B(add_1_root_r112_carry_20_), .Y(
        add_1_root_r112_SUM_20_) );
  AND2X1 U314 ( .A(add_1_root_r112_carry_19_), .B(in_17bit_b[15]), .Y(
        add_1_root_r112_carry_20_) );
  XOR2X1 U315 ( .A(in_17bit_b[15]), .B(add_1_root_r112_carry_19_), .Y(
        add_1_root_r112_SUM_19_) );
  AND2X1 U316 ( .A(add_1_root_r112_carry_18_), .B(in_17bit_b[14]), .Y(
        add_1_root_r112_carry_19_) );
  XOR2X1 U317 ( .A(in_17bit_b[14]), .B(add_1_root_r112_carry_18_), .Y(
        add_1_root_r112_SUM_18_) );
  AND2X1 U318 ( .A(add_1_root_r112_carry_17_), .B(in_17bit_b[13]), .Y(
        add_1_root_r112_carry_18_) );
  XOR2X1 U319 ( .A(in_17bit_b[13]), .B(add_1_root_r112_carry_17_), .Y(
        add_1_root_r112_SUM_17_) );
  AND2X1 U320 ( .A(add_2_root_r119_carry_21_), .B(in_17bit_b[16]), .Y(
        add_2_root_r119_SUM_22_) );
  XOR2X1 U321 ( .A(in_17bit_b[16]), .B(add_2_root_r119_carry_21_), .Y(
        add_2_root_r119_SUM_21_) );
  AND2X1 U322 ( .A(add_1_root_r119_carry[22]), .B(in_17bit_b[16]), .Y(
        add_1_root_r119_SUM_23_) );
  XOR2X1 U323 ( .A(in_17bit_b[16]), .B(add_1_root_r119_carry[22]), .Y(
        add_1_root_r119_SUM_22_) );
  AND2X1 U324 ( .A(add_1_root_r119_carry[21]), .B(in_17bit_b[15]), .Y(
        add_1_root_r119_carry[22]) );
  XOR2X1 U325 ( .A(in_17bit_b[15]), .B(add_1_root_r119_carry[21]), .Y(
        add_1_root_r119_SUM_21_) );
  AND2X1 U326 ( .A(add_1_root_r119_carry[20]), .B(in_17bit_b[14]), .Y(
        add_1_root_r119_carry[21]) );
  XOR2X1 U327 ( .A(in_17bit_b[14]), .B(add_1_root_r119_carry[20]), .Y(
        add_1_root_r119_SUM_20_) );
  AND2X1 U328 ( .A(add_1_root_r119_A_6_), .B(in_17bit_b[0]), .Y(
        add_1_root_r119_carry[7]) );
  XOR2X1 U329 ( .A(in_17bit_b[0]), .B(add_1_root_r119_A_6_), .Y(
        add_1_root_r119_SUM_6_) );
  AND2X1 U330 ( .A(add_3_root_r119_carry_18_), .B(in_17bit_b[16]), .Y(
        add_1_root_r119_A_19_) );
  XOR2X1 U331 ( .A(in_17bit_b[16]), .B(add_3_root_r119_carry_18_), .Y(
        add_1_root_r119_A_18_) );
  AND2X1 U332 ( .A(in_17bit_b[1]), .B(in_17bit_b[0]), .Y(
        add_3_root_r119_carry_3_) );
  XOR2X1 U333 ( .A(in_17bit_b[0]), .B(in_17bit_b[1]), .Y(add_1_root_r119_A_2_)
         );
  AND2X1 U334 ( .A(add_2_root_r115_carry_19_), .B(in_17bit_b[16]), .Y(
        add_2_root_r115_SUM_20_) );
  XOR2X1 U335 ( .A(in_17bit_b[16]), .B(add_2_root_r115_carry_19_), .Y(
        add_2_root_r115_SUM_19_) );
  AND2X1 U336 ( .A(add_2_root_r115_carry_18_), .B(in_17bit_b[15]), .Y(
        add_2_root_r115_carry_19_) );
  XOR2X1 U337 ( .A(in_17bit_b[15]), .B(add_2_root_r115_carry_18_), .Y(
        add_2_root_r115_SUM_18_) );
  AND2X1 U338 ( .A(in_17bit_b[2]), .B(in_17bit_b[0]), .Y(
        add_2_root_r115_carry_4_) );
  AND2X1 U339 ( .A(add_1_root_r115_carry_22_), .B(in_17bit_b[16]), .Y(
        add_1_root_r115_SUM_23_) );
  XOR2X1 U340 ( .A(in_17bit_b[16]), .B(add_1_root_r115_carry_22_), .Y(
        add_1_root_r115_SUM_22_) );
  AND2X1 U341 ( .A(add_1_root_r115_carry_21_), .B(in_17bit_b[15]), .Y(
        add_1_root_r115_carry_22_) );
  XOR2X1 U342 ( .A(in_17bit_b[15]), .B(add_1_root_r115_carry_21_), .Y(
        add_1_root_r115_SUM_21_) );
  XOR2X1 U343 ( .A(in_17bit_b[0]), .B(in_17bit_b[2]), .Y(
        add_1_root_r115_SUM_6_) );
  XOR2X1 U344 ( .A(n21), .B(sub_add_54_b0_carry[16]), .Y(N29) );
  AND2X1 U345 ( .A(sub_add_54_b0_carry[15]), .B(n193), .Y(
        sub_add_54_b0_carry[16]) );
  XOR2X1 U346 ( .A(n193), .B(sub_add_54_b0_carry[15]), .Y(N28) );
  AND2X1 U347 ( .A(sub_add_54_b0_carry[14]), .B(n192), .Y(
        sub_add_54_b0_carry[15]) );
  XOR2X1 U348 ( .A(n192), .B(sub_add_54_b0_carry[14]), .Y(N27) );
  AND2X1 U349 ( .A(sub_add_54_b0_carry[13]), .B(n191), .Y(
        sub_add_54_b0_carry[14]) );
  XOR2X1 U350 ( .A(n191), .B(sub_add_54_b0_carry[13]), .Y(N26) );
  AND2X1 U351 ( .A(sub_add_54_b0_carry[12]), .B(n190), .Y(
        sub_add_54_b0_carry[13]) );
  XOR2X1 U352 ( .A(n190), .B(sub_add_54_b0_carry[12]), .Y(N25) );
  AND2X1 U353 ( .A(sub_add_54_b0_carry[11]), .B(n189), .Y(
        sub_add_54_b0_carry[12]) );
  XOR2X1 U354 ( .A(n189), .B(sub_add_54_b0_carry[11]), .Y(N24) );
  AND2X1 U355 ( .A(sub_add_54_b0_carry[10]), .B(n188), .Y(
        sub_add_54_b0_carry[11]) );
  XOR2X1 U356 ( .A(n188), .B(sub_add_54_b0_carry[10]), .Y(N23) );
  AND2X1 U357 ( .A(sub_add_54_b0_carry[9]), .B(n187), .Y(
        sub_add_54_b0_carry[10]) );
  XOR2X1 U358 ( .A(n187), .B(sub_add_54_b0_carry[9]), .Y(N22) );
  AND2X1 U359 ( .A(sub_add_54_b0_carry[8]), .B(n186), .Y(
        sub_add_54_b0_carry[9]) );
  XOR2X1 U360 ( .A(n186), .B(sub_add_54_b0_carry[8]), .Y(N21) );
  AND2X1 U361 ( .A(sub_add_54_b0_carry[7]), .B(n185), .Y(
        sub_add_54_b0_carry[8]) );
  XOR2X1 U362 ( .A(n185), .B(sub_add_54_b0_carry[7]), .Y(N20) );
  AND2X1 U363 ( .A(sub_add_54_b0_carry[6]), .B(n184), .Y(
        sub_add_54_b0_carry[7]) );
  XOR2X1 U364 ( .A(n184), .B(sub_add_54_b0_carry[6]), .Y(N19) );
  AND2X1 U365 ( .A(sub_add_54_b0_carry[5]), .B(n183), .Y(
        sub_add_54_b0_carry[6]) );
  XOR2X1 U366 ( .A(n183), .B(sub_add_54_b0_carry[5]), .Y(N18) );
  AND2X1 U367 ( .A(sub_add_54_b0_carry[4]), .B(n182), .Y(
        sub_add_54_b0_carry[5]) );
  XOR2X1 U368 ( .A(n182), .B(sub_add_54_b0_carry[4]), .Y(N17) );
  AND2X1 U369 ( .A(sub_add_54_b0_carry[3]), .B(n181), .Y(
        sub_add_54_b0_carry[4]) );
  XOR2X1 U370 ( .A(n181), .B(sub_add_54_b0_carry[3]), .Y(N16) );
  AND2X1 U371 ( .A(sub_add_54_b0_carry[2]), .B(n180), .Y(
        sub_add_54_b0_carry[3]) );
  XOR2X1 U372 ( .A(n180), .B(sub_add_54_b0_carry[2]), .Y(N15) );
  AND2X1 U373 ( .A(n178), .B(n179), .Y(sub_add_54_b0_carry[2]) );
  XOR2X1 U374 ( .A(n179), .B(n178), .Y(N14) );
  XOR2X1 U375 ( .A(n17), .B(sub_add_75_b0_carry[16]), .Y(N481) );
  AND2X1 U376 ( .A(sub_add_75_b0_carry[15]), .B(n12), .Y(
        sub_add_75_b0_carry[16]) );
  XOR2X1 U377 ( .A(n12), .B(sub_add_75_b0_carry[15]), .Y(N480) );
  AND2X1 U378 ( .A(sub_add_75_b0_carry[14]), .B(n13), .Y(
        sub_add_75_b0_carry[15]) );
  XOR2X1 U379 ( .A(n13), .B(sub_add_75_b0_carry[14]), .Y(N479) );
  AND2X1 U380 ( .A(sub_add_75_b0_carry[13]), .B(n16), .Y(
        sub_add_75_b0_carry[14]) );
  AND2X1 U381 ( .A(n31), .B(n15), .Y(sub_add_75_b0_carry[13]) );
  AND2X1 U382 ( .A(in_17bit_b[0]), .B(in_17bit_b[4]), .Y(
        add_1_root_r112_carry_5_) );
endmodule


module multi16_9_DW01_add_0 ( A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, 
        A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, 
        A_4_, B_23_, B_22_, B_21_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, 
        B_14_, B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, 
        SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, 
        SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, 
        SUM_7_ );
  input A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_,
         A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, B_23_, B_22_,
         B_21_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_,
         B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_;
  output SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_,
         SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_,
         SUM_8_, SUM_7_;
  wire   n1, n2, n3, n4;
  wire   [23:7] carry;

  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry[7]), .CO(carry[8]), .S(SUM_7_)
         );
  ADDFX2 U1_21 ( .A(A_21_), .B(B_21_), .CI(carry[21]), .CO(carry[22]), .S(
        SUM_21_) );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry[20]), .CO(carry[21]), .S(
        SUM_20_) );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry[19]), .CO(carry[20]), .S(
        SUM_19_) );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry[18]), .CO(carry[19]), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry[17]), .CO(carry[18]), .S(
        SUM_17_) );
  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry[16]), .CO(carry[17]), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry[15]), .CO(carry[16]), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry[14]), .CO(carry[15]), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry[13]), .CO(carry[14]), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry[12]), .CO(carry[13]), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry[11]), .CO(carry[12]), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry[10]), .CO(carry[11]), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry[9]), .CO(carry[10]), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry[8]), .CO(carry[9]), .S(SUM_8_)
         );
  ADDFX2 U1_22 ( .A(A_22_), .B(B_22_), .CI(carry[22]), .CO(carry[23]), .S(
        SUM_22_) );
  AND2X2 U1 ( .A(A_4_), .B(B_4_), .Y(n1) );
  XOR2X1 U2 ( .A(B_23_), .B(carry[23]), .Y(SUM_23_) );
  OAI2BB1X1 U3 ( .A0N(n2), .A1N(A_6_), .B0(n3), .Y(carry[7]) );
  OAI21XL U4 ( .A0(A_6_), .A1(n2), .B0(B_6_), .Y(n3) );
  OAI2BB1X1 U5 ( .A0N(n1), .A1N(A_5_), .B0(n4), .Y(n2) );
  OAI21XL U6 ( .A0(A_5_), .A1(n1), .B0(B_5_), .Y(n4) );
endmodule


module multi16_9_DW01_add_4 ( A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, 
        A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, 
        B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, 
        B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, SUM_22_, SUM_21_, SUM_20_, 
        SUM_19_, SUM_18_, SUM_17_, SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, 
        SUM_11_, SUM_10_, SUM_9_, SUM_8_, SUM_7_ );
  input A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_,
         A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, B_20_, B_19_,
         B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, B_10_, B_9_,
         B_8_, B_7_, B_6_, B_5_;
  output SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_,
         SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_,
         SUM_7_;
  wire   carry_21_, carry_20_, carry_19_, carry_18_, carry_17_, carry_16_,
         carry_15_, carry_14_, carry_13_, carry_12_, carry_11_, carry_10_,
         carry_9_, carry_8_, carry_7_, n1;

  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry_16_), .CO(carry_17_), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry_15_), .CO(carry_16_), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry_14_), .CO(carry_15_), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry_13_), .CO(carry_14_), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry_12_), .CO(carry_13_), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry_11_), .CO(carry_12_), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry_10_), .CO(carry_11_), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry_9_), .CO(carry_10_), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry_8_), .CO(carry_9_), .S(SUM_8_)
         );
  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry_7_), .CO(carry_8_), .S(SUM_7_)
         );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry_20_), .CO(carry_21_), .S(
        SUM_20_) );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry_19_), .CO(carry_20_), .S(
        SUM_19_) );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry_18_), .CO(carry_19_), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry_17_), .CO(carry_18_), .S(
        SUM_17_) );
  ADDFX2 U1_21 ( .A(A_21_), .B(B_21_), .CI(carry_21_), .CO(SUM_22_), .S(
        SUM_21_) );
  OAI2BB1X1 U1 ( .A0N(A_6_), .A1N(B_6_), .B0(n1), .Y(carry_7_) );
  OAI211X1 U2 ( .A0(B_6_), .A1(A_6_), .B0(A_5_), .C0(B_5_), .Y(n1) );
endmodule


module multi16_9_DW01_add_6 ( A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, 
        A_16_, A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, 
        A_6_, A_5_, A_4_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, 
        B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, 
        SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, 
        SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, 
        SUM_7_ );
  input A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_,
         A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, B_20_,
         B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, B_10_,
         B_9_, B_8_, B_7_, B_6_, B_5_, B_4_;
  output SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_,
         SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_,
         SUM_8_, SUM_7_;
  wire   n1, n2, n3, n4, n5, n6;
  wire   [21:7] carry;

  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry[7]), .CO(carry[8]), .S(SUM_7_)
         );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry[18]), .CO(carry[19]), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry[17]), .CO(carry[18]), .S(
        SUM_17_) );
  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry[16]), .CO(carry[17]), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry[15]), .CO(carry[16]), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry[14]), .CO(carry[15]), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry[13]), .CO(carry[14]), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry[12]), .CO(carry[13]), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry[11]), .CO(carry[12]), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry[10]), .CO(carry[11]), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry[9]), .CO(carry[10]), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry[8]), .CO(carry[9]), .S(SUM_8_)
         );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry[19]), .CO(carry[20]), .S(
        SUM_19_) );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry[20]), .CO(carry[21]), .S(
        SUM_20_) );
  AND2X2 U1 ( .A(A_22_), .B(n2), .Y(n1) );
  AND2X2 U2 ( .A(A_21_), .B(carry[21]), .Y(n2) );
  AND2X2 U3 ( .A(A_4_), .B(B_4_), .Y(n3) );
  XOR2X1 U4 ( .A(A_23_), .B(n1), .Y(SUM_23_) );
  XOR2X1 U5 ( .A(A_21_), .B(carry[21]), .Y(SUM_21_) );
  XOR2X1 U6 ( .A(A_22_), .B(n2), .Y(SUM_22_) );
  OAI2BB1X1 U7 ( .A0N(n4), .A1N(A_6_), .B0(n5), .Y(carry[7]) );
  OAI21XL U8 ( .A0(A_6_), .A1(n4), .B0(B_6_), .Y(n5) );
  OAI2BB1X1 U9 ( .A0N(n3), .A1N(A_5_), .B0(n6), .Y(n4) );
  OAI21XL U10 ( .A0(A_5_), .A1(n3), .B0(B_5_), .Y(n6) );
endmodule


module multi16_9 ( in_17bit, in_8bit, out );
  input [16:0] in_17bit;
  input [7:0] in_8bit;
  output [16:0] out;
  wire   n289, n290, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24,
         N25, N26, N27, N28, N29, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, N205, N206,
         N207, N208, N209, N210, N211, N212, N213, N214, N215, N216, N217,
         N218, N219, N220, N221, N347, N348, N349, N350, N351, N352, N353,
         N354, N355, N356, N357, N358, N359, N360, N361, N362, N363, N446,
         N447, N448, N449, N450, N451, N452, N453, N454, N455, N456, N457,
         N458, N459, N460, N461, N462, N463, N479, N480,
         add_2_root_r119_carry_10_, add_2_root_r119_carry_11_,
         add_2_root_r119_carry_12_, add_2_root_r119_carry_13_,
         add_2_root_r119_carry_14_, add_2_root_r119_carry_15_,
         add_2_root_r119_carry_16_, add_2_root_r119_carry_17_,
         add_2_root_r119_carry_18_, add_2_root_r119_carry_19_,
         add_2_root_r119_carry_20_, add_2_root_r119_carry_21_,
         add_2_root_r119_carry_7_, add_2_root_r119_carry_8_,
         add_2_root_r119_carry_9_, add_2_root_r119_SUM_6_,
         add_2_root_r119_SUM_7_, add_2_root_r119_SUM_8_,
         add_2_root_r119_SUM_9_, add_2_root_r119_SUM_10_,
         add_2_root_r119_SUM_11_, add_2_root_r119_SUM_12_,
         add_2_root_r119_SUM_13_, add_2_root_r119_SUM_14_,
         add_2_root_r119_SUM_15_, add_2_root_r119_SUM_16_,
         add_2_root_r119_SUM_17_, add_2_root_r119_SUM_18_,
         add_2_root_r119_SUM_19_, add_2_root_r119_SUM_20_,
         add_2_root_r119_SUM_21_, add_2_root_r119_SUM_22_,
         add_1_root_r119_SUM_6_, add_1_root_r119_SUM_7_,
         add_1_root_r119_SUM_8_, add_1_root_r119_SUM_9_,
         add_1_root_r119_SUM_10_, add_1_root_r119_SUM_11_,
         add_1_root_r119_SUM_12_, add_1_root_r119_SUM_13_,
         add_1_root_r119_SUM_14_, add_1_root_r119_SUM_15_,
         add_1_root_r119_SUM_16_, add_1_root_r119_SUM_17_,
         add_1_root_r119_SUM_18_, add_1_root_r119_SUM_19_,
         add_1_root_r119_SUM_20_, add_1_root_r119_SUM_21_,
         add_1_root_r119_SUM_22_, add_1_root_r119_SUM_23_,
         add_1_root_r119_A_2_, add_1_root_r119_A_3_, add_1_root_r119_A_4_,
         add_1_root_r119_A_5_, add_1_root_r119_A_6_, add_1_root_r119_A_7_,
         add_1_root_r119_A_8_, add_1_root_r119_A_9_, add_1_root_r119_A_10_,
         add_1_root_r119_A_11_, add_1_root_r119_A_12_, add_1_root_r119_A_13_,
         add_1_root_r119_A_14_, add_1_root_r119_A_15_, add_1_root_r119_A_16_,
         add_1_root_r119_A_17_, add_1_root_r119_A_18_, add_1_root_r119_A_19_,
         add_3_root_r119_carry_10_, add_3_root_r119_carry_11_,
         add_3_root_r119_carry_12_, add_3_root_r119_carry_13_,
         add_3_root_r119_carry_14_, add_3_root_r119_carry_15_,
         add_3_root_r119_carry_16_, add_3_root_r119_carry_17_,
         add_3_root_r119_carry_18_, add_3_root_r119_carry_3_,
         add_3_root_r119_carry_4_, add_3_root_r119_carry_5_,
         add_3_root_r119_carry_6_, add_3_root_r119_carry_7_,
         add_3_root_r119_carry_8_, add_3_root_r119_carry_9_,
         add_1_root_r112_carry_10_, add_1_root_r112_carry_11_,
         add_1_root_r112_carry_12_, add_1_root_r112_carry_13_,
         add_1_root_r112_carry_14_, add_1_root_r112_carry_15_,
         add_1_root_r112_carry_16_, add_1_root_r112_carry_17_,
         add_1_root_r112_carry_18_, add_1_root_r112_carry_19_,
         add_1_root_r112_carry_20_, add_1_root_r112_carry_5_,
         add_1_root_r112_carry_6_, add_1_root_r112_carry_7_,
         add_1_root_r112_carry_8_, add_1_root_r112_carry_9_,
         add_1_root_r112_SUM_1_, add_1_root_r112_SUM_2_,
         add_1_root_r112_SUM_3_, add_1_root_r112_SUM_4_,
         add_1_root_r112_SUM_5_, add_1_root_r112_SUM_6_,
         add_1_root_r112_SUM_7_, add_1_root_r112_SUM_8_,
         add_1_root_r112_SUM_9_, add_1_root_r112_SUM_10_,
         add_1_root_r112_SUM_11_, add_1_root_r112_SUM_12_,
         add_1_root_r112_SUM_13_, add_1_root_r112_SUM_14_,
         add_1_root_r112_SUM_15_, add_1_root_r112_SUM_16_,
         add_1_root_r112_SUM_17_, add_1_root_r112_SUM_18_,
         add_1_root_r112_SUM_19_, add_1_root_r112_SUM_20_,
         add_1_root_r112_SUM_21_, add_2_root_r115_carry_10_,
         add_2_root_r115_carry_11_, add_2_root_r115_carry_12_,
         add_2_root_r115_carry_13_, add_2_root_r115_carry_14_,
         add_2_root_r115_carry_15_, add_2_root_r115_carry_16_,
         add_2_root_r115_carry_17_, add_2_root_r115_carry_18_,
         add_2_root_r115_carry_19_, add_2_root_r115_carry_5_,
         add_2_root_r115_carry_6_, add_2_root_r115_carry_7_,
         add_2_root_r115_carry_8_, add_2_root_r115_carry_9_,
         add_2_root_r115_SUM_4_, add_2_root_r115_SUM_5_,
         add_2_root_r115_SUM_6_, add_2_root_r115_SUM_7_,
         add_2_root_r115_SUM_8_, add_2_root_r115_SUM_9_,
         add_2_root_r115_SUM_10_, add_2_root_r115_SUM_11_,
         add_2_root_r115_SUM_12_, add_2_root_r115_SUM_13_,
         add_2_root_r115_SUM_14_, add_2_root_r115_SUM_15_,
         add_2_root_r115_SUM_16_, add_2_root_r115_SUM_17_,
         add_2_root_r115_SUM_18_, add_2_root_r115_SUM_19_,
         add_2_root_r115_SUM_20_, add_1_root_r115_carry_10_,
         add_1_root_r115_carry_11_, add_1_root_r115_carry_12_,
         add_1_root_r115_carry_13_, add_1_root_r115_carry_14_,
         add_1_root_r115_carry_15_, add_1_root_r115_carry_16_,
         add_1_root_r115_carry_17_, add_1_root_r115_carry_18_,
         add_1_root_r115_carry_19_, add_1_root_r115_carry_20_,
         add_1_root_r115_carry_21_, add_1_root_r115_carry_22_,
         add_1_root_r115_carry_7_, add_1_root_r115_carry_8_,
         add_1_root_r115_carry_9_, add_1_root_r115_SUM_6_,
         add_1_root_r115_SUM_7_, add_1_root_r115_SUM_8_,
         add_1_root_r115_SUM_9_, add_1_root_r115_SUM_10_,
         add_1_root_r115_SUM_11_, add_1_root_r115_SUM_12_,
         add_1_root_r115_SUM_13_, add_1_root_r115_SUM_14_,
         add_1_root_r115_SUM_15_, add_1_root_r115_SUM_16_,
         add_1_root_r115_SUM_17_, add_1_root_r115_SUM_18_,
         add_1_root_r115_SUM_19_, add_1_root_r115_SUM_20_,
         add_1_root_r115_SUM_21_, add_1_root_r115_SUM_22_,
         add_1_root_r115_SUM_23_, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n17, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288;
  wire   [16:0] in_17bit_b;
  wire   [23:8] neg_mul;
  wire   [15:13] sub_add_75_b0_carry;
  wire   [16:2] sub_add_54_b0_carry;
  wire   [22:7] add_1_root_r119_carry;

  multi16_9_DW01_add_0 add_0_root_r119 ( .A_22_(add_2_root_r119_SUM_22_), 
        .A_21_(add_2_root_r119_SUM_21_), .A_20_(add_2_root_r119_SUM_20_), 
        .A_19_(add_2_root_r119_SUM_19_), .A_18_(add_2_root_r119_SUM_18_), 
        .A_17_(add_2_root_r119_SUM_17_), .A_16_(add_2_root_r119_SUM_16_), 
        .A_15_(add_2_root_r119_SUM_15_), .A_14_(add_2_root_r119_SUM_14_), 
        .A_13_(add_2_root_r119_SUM_13_), .A_12_(add_2_root_r119_SUM_12_), 
        .A_11_(add_2_root_r119_SUM_11_), .A_10_(add_2_root_r119_SUM_10_), 
        .A_9_(add_2_root_r119_SUM_9_), .A_8_(add_2_root_r119_SUM_8_), .A_7_(
        add_2_root_r119_SUM_7_), .A_6_(add_2_root_r119_SUM_6_), .A_5_(
        add_1_root_r119_A_2_), .A_4_(in_17bit_b[0]), .B_23_(
        add_1_root_r119_SUM_23_), .B_22_(add_1_root_r119_SUM_22_), .B_21_(
        add_1_root_r119_SUM_21_), .B_20_(add_1_root_r119_SUM_20_), .B_19_(
        add_1_root_r119_SUM_19_), .B_18_(add_1_root_r119_SUM_18_), .B_17_(
        add_1_root_r119_SUM_17_), .B_16_(add_1_root_r119_SUM_16_), .B_15_(
        add_1_root_r119_SUM_15_), .B_14_(add_1_root_r119_SUM_14_), .B_13_(
        add_1_root_r119_SUM_13_), .B_12_(add_1_root_r119_SUM_12_), .B_11_(
        add_1_root_r119_SUM_11_), .B_10_(add_1_root_r119_SUM_10_), .B_9_(
        add_1_root_r119_SUM_9_), .B_8_(add_1_root_r119_SUM_8_), .B_7_(
        add_1_root_r119_SUM_7_), .B_6_(add_1_root_r119_SUM_6_), .B_5_(
        add_1_root_r119_A_5_), .B_4_(add_1_root_r119_A_4_), .SUM_23_(N363), 
        .SUM_22_(N362), .SUM_21_(N361), .SUM_20_(N360), .SUM_19_(N359), 
        .SUM_18_(N358), .SUM_17_(N357), .SUM_16_(N356), .SUM_15_(N355), 
        .SUM_14_(N354), .SUM_13_(N353), .SUM_12_(N352), .SUM_11_(N351), 
        .SUM_10_(N350), .SUM_9_(N349), .SUM_8_(N348), .SUM_7_(N347) );
  multi16_9_DW01_add_4 add_0_root_r112 ( .A_21_(in_17bit_b[16]), .A_20_(
        in_17bit_b[15]), .A_19_(in_17bit_b[14]), .A_18_(in_17bit_b[13]), 
        .A_17_(in_17bit_b[12]), .A_16_(in_17bit_b[11]), .A_15_(in_17bit_b[10]), 
        .A_14_(in_17bit_b[9]), .A_13_(in_17bit_b[8]), .A_12_(in_17bit_b[7]), 
        .A_11_(in_17bit_b[6]), .A_10_(in_17bit_b[5]), .A_9_(in_17bit_b[4]), 
        .A_8_(in_17bit_b[3]), .A_7_(in_17bit_b[2]), .A_6_(in_17bit_b[1]), 
        .A_5_(in_17bit_b[0]), .B_21_(add_1_root_r112_SUM_21_), .B_20_(
        add_1_root_r112_SUM_20_), .B_19_(add_1_root_r112_SUM_19_), .B_18_(
        add_1_root_r112_SUM_18_), .B_17_(add_1_root_r112_SUM_17_), .B_16_(
        add_1_root_r112_SUM_16_), .B_15_(add_1_root_r112_SUM_15_), .B_14_(
        add_1_root_r112_SUM_14_), .B_13_(add_1_root_r112_SUM_13_), .B_12_(
        add_1_root_r112_SUM_12_), .B_11_(add_1_root_r112_SUM_11_), .B_10_(
        add_1_root_r112_SUM_10_), .B_9_(add_1_root_r112_SUM_9_), .B_8_(
        add_1_root_r112_SUM_8_), .B_7_(add_1_root_r112_SUM_7_), .B_6_(
        add_1_root_r112_SUM_6_), .B_5_(add_1_root_r112_SUM_5_), .SUM_22_(N123), 
        .SUM_21_(N122), .SUM_20_(N121), .SUM_19_(N120), .SUM_18_(N119), 
        .SUM_17_(N118), .SUM_16_(N117), .SUM_15_(N116), .SUM_14_(N115), 
        .SUM_13_(N114), .SUM_12_(N113), .SUM_11_(N112), .SUM_10_(N111), 
        .SUM_9_(N110), .SUM_8_(N109), .SUM_7_(N108) );
  multi16_9_DW01_add_6 add_0_root_r115 ( .A_23_(add_1_root_r115_SUM_23_), 
        .A_22_(add_1_root_r115_SUM_22_), .A_21_(add_1_root_r115_SUM_21_), 
        .A_20_(add_1_root_r115_SUM_20_), .A_19_(add_1_root_r115_SUM_19_), 
        .A_18_(add_1_root_r115_SUM_18_), .A_17_(add_1_root_r115_SUM_17_), 
        .A_16_(add_1_root_r115_SUM_16_), .A_15_(add_1_root_r115_SUM_15_), 
        .A_14_(add_1_root_r115_SUM_14_), .A_13_(add_1_root_r115_SUM_13_), 
        .A_12_(add_1_root_r115_SUM_12_), .A_11_(add_1_root_r115_SUM_11_), 
        .A_10_(add_1_root_r115_SUM_10_), .A_9_(add_1_root_r115_SUM_9_), .A_8_(
        add_1_root_r115_SUM_8_), .A_7_(add_1_root_r115_SUM_7_), .A_6_(
        add_1_root_r115_SUM_6_), .A_5_(in_17bit_b[1]), .A_4_(in_17bit_b[0]), 
        .B_20_(add_2_root_r115_SUM_20_), .B_19_(add_2_root_r115_SUM_19_), 
        .B_18_(add_2_root_r115_SUM_18_), .B_17_(add_2_root_r115_SUM_17_), 
        .B_16_(add_2_root_r115_SUM_16_), .B_15_(add_2_root_r115_SUM_15_), 
        .B_14_(add_2_root_r115_SUM_14_), .B_13_(add_2_root_r115_SUM_13_), 
        .B_12_(add_2_root_r115_SUM_12_), .B_11_(add_2_root_r115_SUM_11_), 
        .B_10_(add_2_root_r115_SUM_10_), .B_9_(add_2_root_r115_SUM_9_), .B_8_(
        add_2_root_r115_SUM_8_), .B_7_(add_2_root_r115_SUM_7_), .B_6_(
        add_2_root_r115_SUM_6_), .B_5_(add_2_root_r115_SUM_5_), .B_4_(
        add_2_root_r115_SUM_4_), .SUM_23_(N221), .SUM_22_(N220), .SUM_21_(N219), .SUM_20_(N218), .SUM_19_(N217), .SUM_18_(N216), .SUM_17_(N215), .SUM_16_(
        N214), .SUM_15_(N213), .SUM_14_(N212), .SUM_13_(N211), .SUM_12_(N210), 
        .SUM_11_(N209), .SUM_10_(N208), .SUM_9_(N207), .SUM_8_(N206), .SUM_7_(
        N205) );
  TLATX1 neg_mul_reg_19_ ( .G(N446), .D(N459), .QN(n8) );
  TLATX1 neg_mul_reg_18_ ( .G(N446), .D(N458), .QN(n7) );
  TLATX1 neg_mul_reg_17_ ( .G(N446), .D(N457), .Q(neg_mul[17]), .QN(n5) );
  TLATX1 neg_mul_reg_16_ ( .G(N446), .D(N456), .Q(neg_mul[16]), .QN(n4) );
  TLATX1 neg_mul_reg_11_ ( .G(N446), .D(N451), .Q(neg_mul[11]), .QN(n3) );
  TLATX1 neg_mul_reg_23_ ( .G(N446), .D(N463), .Q(neg_mul[23]), .QN(n6) );
  TLATX1 neg_mul_reg_22_ ( .G(N446), .D(N462), .Q(neg_mul[22]), .QN(n9) );
  TLATX1 neg_mul_reg_21_ ( .G(N446), .D(N461), .Q(neg_mul[21]), .QN(n10) );
  TLATX1 neg_mul_reg_20_ ( .G(N446), .D(N460), .QN(n11) );
  TLATX1 neg_mul_reg_8_ ( .G(N446), .D(N448), .Q(neg_mul[8]) );
  TLATX1 neg_mul_reg_9_ ( .G(N446), .D(N449), .Q(neg_mul[9]), .QN(n14) );
  TLATX1 neg_mul_reg_15_ ( .G(N446), .D(N455), .Q(neg_mul[15]) );
  TLATX1 neg_mul_reg_14_ ( .G(N446), .D(N454), .Q(neg_mul[14]), .QN(n13) );
  TLATX1 neg_mul_reg_13_ ( .G(N446), .D(N453), .Q(neg_mul[13]), .QN(n12) );
  TLATX1 neg_mul_reg_12_ ( .G(N446), .D(N452), .Q(neg_mul[12]) );
  TLATX1 neg_mul_reg_10_ ( .G(N446), .D(N450), .Q(neg_mul[10]) );
  TLATX1 neg_mul_reg_7_ ( .G(N446), .D(N447), .Q(out[0]) );
  XOR2X4 U2 ( .A(n180), .B(n1), .Y(out[11]) );
  CLKINVX20 U3 ( .A(n7), .Y(n1) );
  BUFX20 U4 ( .A(n43), .Y(n23) );
  NOR2X2 U5 ( .A(n23), .B(n88), .Y(n90) );
  CLKINVX1 U6 ( .A(n22), .Y(n45) );
  CLKINVX3 U7 ( .A(n288), .Y(in_17bit_b[16]) );
  NOR2BX4 U8 ( .AN(n2), .B(n71), .Y(n73) );
  CLKINVX20 U9 ( .A(n72), .Y(n2) );
  INVX8 U10 ( .A(in_17bit[16]), .Y(n46) );
  AOI211X4 U11 ( .A0(n42), .A1(n176), .B0(n175), .C0(n29), .Y(out[8]) );
  INVX1 U12 ( .A(n25), .Y(n19) );
  NOR2X1 U13 ( .A(n97), .B(n44), .Y(n99) );
  AOI22X1 U14 ( .A0(N27), .A1(n22), .B0(in_17bit[14]), .B1(n45), .Y(n277) );
  XNOR2X1 U15 ( .A(neg_mul[23]), .B(n30), .Y(n15) );
  DLY1X1 U16 ( .A(n23), .Y(n22) );
  INVX12 U17 ( .A(n177), .Y(n181) );
  OAI21X4 U18 ( .A0(n52), .A1(n43), .B0(n51), .Y(n53) );
  XOR2X4 U19 ( .A(n73), .B(neg_mul[11]), .Y(out[4]) );
  CLKINVX8 U20 ( .A(n46), .Y(n43) );
  OAI2BB1X2 U21 ( .A0N(n21), .A1N(n46), .B0(n68), .Y(n69) );
  NOR2X4 U22 ( .A(n23), .B(n79), .Y(n81) );
  XNOR2X4 U23 ( .A(n42), .B(in_8bit[7]), .Y(n179) );
  XNOR2X4 U24 ( .A(n42), .B(in_8bit[7]), .Y(n177) );
  BUFX8 U25 ( .A(n289), .Y(out[7]) );
  AOI211X2 U26 ( .A0(n42), .A1(n100), .B0(n99), .C0(n98), .Y(n289) );
  XOR2X4 U27 ( .A(n178), .B(neg_mul[16]), .Y(out[9]) );
  XNOR2X4 U28 ( .A(n17), .B(neg_mul[17]), .Y(out[10]) );
  NAND2X4 U29 ( .A(n19), .B(n20), .Y(n17) );
  NOR2X1 U30 ( .A(n42), .B(n174), .Y(n175) );
  INVX4 U31 ( .A(n46), .Y(n44) );
  NOR2X4 U32 ( .A(n26), .B(n179), .Y(n180) );
  BUFX8 U33 ( .A(n290), .Y(out[6]) );
  AOI211X2 U34 ( .A0(n23), .A1(n91), .B0(n90), .C0(n89), .Y(n290) );
  AOI211X2 U35 ( .A0(n42), .A1(n82), .B0(n81), .C0(n80), .Y(out[5]) );
  INVX20 U36 ( .A(n46), .Y(n42) );
  XOR2X2 U37 ( .A(n42), .B(in_8bit[7]), .Y(n20) );
  NOR2X4 U38 ( .A(n29), .B(n177), .Y(n178) );
  OR2X2 U39 ( .A(n67), .B(n66), .Y(n21) );
  MX2X2 U40 ( .A(neg_mul[21]), .B(N479), .S0(n181), .Y(out[14]) );
  INVX1 U41 ( .A(n238), .Y(in_17bit_b[1]) );
  INVX1 U42 ( .A(n277), .Y(in_17bit_b[14]) );
  INVX1 U43 ( .A(n274), .Y(in_17bit_b[13]) );
  INVX1 U44 ( .A(n241), .Y(in_17bit_b[2]) );
  INVX1 U45 ( .A(n250), .Y(in_17bit_b[5]) );
  INVX1 U46 ( .A(n253), .Y(in_17bit_b[6]) );
  INVX1 U47 ( .A(n256), .Y(in_17bit_b[7]) );
  INVX1 U48 ( .A(n262), .Y(in_17bit_b[9]) );
  INVX1 U49 ( .A(n265), .Y(in_17bit_b[10]) );
  INVX1 U50 ( .A(n268), .Y(in_17bit_b[11]) );
  INVX1 U51 ( .A(n271), .Y(in_17bit_b[12]) );
  INVX1 U52 ( .A(n259), .Y(in_17bit_b[8]) );
  INVX1 U53 ( .A(n247), .Y(in_17bit_b[4]) );
  INVX1 U54 ( .A(n244), .Y(in_17bit_b[3]) );
  XOR2X4 U55 ( .A(n24), .B(n8), .Y(out[12]) );
  OR2X4 U56 ( .A(n179), .B(n27), .Y(n24) );
  ADDFX2 U57 ( .A(in_17bit_b[16]), .B(in_17bit_b[12]), .CI(
        add_1_root_r112_carry_16_), .CO(add_1_root_r112_carry_17_), .S(
        add_1_root_r112_SUM_16_) );
  ADDFX2 U58 ( .A(add_1_root_r119_A_19_), .B(in_17bit_b[13]), .CI(
        add_1_root_r119_carry[19]), .CO(add_1_root_r119_carry[20]), .S(
        add_1_root_r119_SUM_19_) );
  ADDFX2 U59 ( .A(in_17bit_b[16]), .B(in_17bit_b[15]), .CI(
        add_3_root_r119_carry_17_), .CO(add_3_root_r119_carry_18_), .S(
        add_1_root_r119_A_17_) );
  ADDFX2 U60 ( .A(in_17bit_b[16]), .B(in_17bit_b[14]), .CI(
        add_2_root_r115_carry_17_), .CO(add_2_root_r115_carry_18_), .S(
        add_2_root_r115_SUM_17_) );
  ADDFX2 U61 ( .A(in_17bit_b[16]), .B(in_17bit_b[14]), .CI(
        add_1_root_r115_carry_20_), .CO(add_1_root_r115_carry_21_), .S(
        add_1_root_r115_SUM_20_) );
  ADDFX2 U62 ( .A(in_17bit_b[16]), .B(in_17bit_b[15]), .CI(
        add_2_root_r119_carry_20_), .CO(add_2_root_r119_carry_21_), .S(
        add_2_root_r119_SUM_20_) );
  ADDFX2 U63 ( .A(in_17bit_b[3]), .B(in_17bit_b[1]), .CI(
        add_1_root_r115_carry_7_), .CO(add_2_root_r115_carry_5_), .S(
        add_2_root_r115_SUM_4_) );
  ADDFX2 U64 ( .A(in_17bit_b[4]), .B(in_17bit_b[2]), .CI(
        add_2_root_r115_carry_5_), .CO(add_2_root_r115_carry_6_), .S(
        add_2_root_r115_SUM_5_) );
  ADDFX2 U65 ( .A(in_17bit_b[5]), .B(in_17bit_b[1]), .CI(
        add_1_root_r112_carry_5_), .CO(add_1_root_r112_carry_6_), .S(
        add_1_root_r112_SUM_5_) );
  ADDFX2 U66 ( .A(in_17bit_b[6]), .B(in_17bit_b[5]), .CI(
        add_3_root_r119_carry_7_), .CO(add_3_root_r119_carry_8_), .S(
        add_1_root_r119_A_7_) );
  ADDFX2 U67 ( .A(in_17bit_b[6]), .B(in_17bit_b[2]), .CI(
        add_1_root_r112_carry_6_), .CO(add_1_root_r112_carry_7_), .S(
        add_1_root_r112_SUM_6_) );
  ADDFX2 U68 ( .A(in_17bit_b[3]), .B(in_17bit_b[1]), .CI(
        add_1_root_r115_carry_7_), .CO(add_1_root_r115_carry_8_), .S(
        add_1_root_r115_SUM_7_) );
  ADDFX2 U69 ( .A(in_17bit_b[7]), .B(in_17bit_b[6]), .CI(
        add_3_root_r119_carry_8_), .CO(add_3_root_r119_carry_9_), .S(
        add_1_root_r119_A_8_) );
  ADDFX2 U70 ( .A(add_1_root_r119_A_7_), .B(in_17bit_b[1]), .CI(
        add_1_root_r119_carry[7]), .CO(add_1_root_r119_carry[8]), .S(
        add_1_root_r119_SUM_7_) );
  ADDFX2 U71 ( .A(in_17bit_b[2]), .B(in_17bit_b[1]), .CI(
        add_3_root_r119_carry_3_), .CO(add_2_root_r119_carry_7_), .S(
        add_2_root_r119_SUM_6_) );
  ADDFX2 U72 ( .A(in_17bit_b[4]), .B(in_17bit_b[2]), .CI(
        add_1_root_r115_carry_8_), .CO(add_1_root_r115_carry_9_), .S(
        add_1_root_r115_SUM_8_) );
  ADDFX2 U73 ( .A(in_17bit_b[8]), .B(in_17bit_b[7]), .CI(
        add_3_root_r119_carry_9_), .CO(add_3_root_r119_carry_10_), .S(
        add_1_root_r119_A_9_) );
  ADDFX2 U74 ( .A(add_1_root_r119_A_8_), .B(in_17bit_b[2]), .CI(
        add_1_root_r119_carry[8]), .CO(add_1_root_r119_carry[9]), .S(
        add_1_root_r119_SUM_8_) );
  ADDFX2 U75 ( .A(in_17bit_b[3]), .B(in_17bit_b[2]), .CI(
        add_2_root_r119_carry_7_), .CO(add_2_root_r119_carry_8_), .S(
        add_2_root_r119_SUM_7_) );
  ADDFX2 U76 ( .A(in_17bit_b[6]), .B(in_17bit_b[4]), .CI(
        add_2_root_r115_carry_7_), .CO(add_2_root_r115_carry_8_), .S(
        add_2_root_r115_SUM_7_) );
  ADDFX2 U77 ( .A(in_17bit_b[8]), .B(in_17bit_b[4]), .CI(
        add_1_root_r112_carry_8_), .CO(add_1_root_r112_carry_9_), .S(
        add_1_root_r112_SUM_8_) );
  ADDFX2 U78 ( .A(in_17bit_b[9]), .B(in_17bit_b[8]), .CI(
        add_3_root_r119_carry_10_), .CO(add_3_root_r119_carry_11_), .S(
        add_1_root_r119_A_10_) );
  ADDFX2 U79 ( .A(in_17bit_b[7]), .B(in_17bit_b[5]), .CI(
        add_2_root_r115_carry_8_), .CO(add_2_root_r115_carry_9_), .S(
        add_2_root_r115_SUM_8_) );
  ADDFX2 U80 ( .A(in_17bit_b[10]), .B(in_17bit_b[9]), .CI(
        add_3_root_r119_carry_11_), .CO(add_3_root_r119_carry_12_), .S(
        add_1_root_r119_A_11_) );
  ADDFX2 U81 ( .A(add_1_root_r119_A_10_), .B(in_17bit_b[4]), .CI(
        add_1_root_r119_carry[10]), .CO(add_1_root_r119_carry[11]), .S(
        add_1_root_r119_SUM_10_) );
  ADDFX2 U82 ( .A(in_17bit_b[9]), .B(in_17bit_b[5]), .CI(
        add_1_root_r112_carry_9_), .CO(add_1_root_r112_carry_10_), .S(
        add_1_root_r112_SUM_9_) );
  ADDFX2 U83 ( .A(in_17bit_b[8]), .B(in_17bit_b[6]), .CI(
        add_2_root_r115_carry_9_), .CO(add_2_root_r115_carry_10_), .S(
        add_2_root_r115_SUM_9_) );
  ADDFX2 U84 ( .A(in_17bit_b[10]), .B(in_17bit_b[6]), .CI(
        add_1_root_r112_carry_10_), .CO(add_1_root_r112_carry_11_), .S(
        add_1_root_r112_SUM_10_) );
  ADDFX2 U85 ( .A(in_17bit_b[7]), .B(in_17bit_b[5]), .CI(
        add_1_root_r115_carry_11_), .CO(add_1_root_r115_carry_12_), .S(
        add_1_root_r115_SUM_11_) );
  ADDFX2 U86 ( .A(in_17bit_b[11]), .B(in_17bit_b[10]), .CI(
        add_3_root_r119_carry_12_), .CO(add_3_root_r119_carry_13_), .S(
        add_1_root_r119_A_12_) );
  ADDFX2 U87 ( .A(add_1_root_r119_A_11_), .B(in_17bit_b[5]), .CI(
        add_1_root_r119_carry[11]), .CO(add_1_root_r119_carry[12]), .S(
        add_1_root_r119_SUM_11_) );
  ADDFX2 U88 ( .A(in_17bit_b[6]), .B(in_17bit_b[5]), .CI(
        add_2_root_r119_carry_10_), .CO(add_2_root_r119_carry_11_), .S(
        add_2_root_r119_SUM_10_) );
  ADDFX2 U89 ( .A(in_17bit_b[9]), .B(in_17bit_b[7]), .CI(
        add_2_root_r115_carry_10_), .CO(add_2_root_r115_carry_11_), .S(
        add_2_root_r115_SUM_10_) );
  ADDFX2 U90 ( .A(in_17bit_b[11]), .B(in_17bit_b[7]), .CI(
        add_1_root_r112_carry_11_), .CO(add_1_root_r112_carry_12_), .S(
        add_1_root_r112_SUM_11_) );
  ADDFX2 U91 ( .A(in_17bit_b[8]), .B(in_17bit_b[6]), .CI(
        add_1_root_r115_carry_12_), .CO(add_1_root_r115_carry_13_), .S(
        add_1_root_r115_SUM_12_) );
  ADDFX2 U92 ( .A(in_17bit_b[12]), .B(in_17bit_b[11]), .CI(
        add_3_root_r119_carry_13_), .CO(add_3_root_r119_carry_14_), .S(
        add_1_root_r119_A_13_) );
  ADDFX2 U93 ( .A(add_1_root_r119_A_12_), .B(in_17bit_b[6]), .CI(
        add_1_root_r119_carry[12]), .CO(add_1_root_r119_carry[13]), .S(
        add_1_root_r119_SUM_12_) );
  ADDFX2 U94 ( .A(in_17bit_b[7]), .B(in_17bit_b[6]), .CI(
        add_2_root_r119_carry_11_), .CO(add_2_root_r119_carry_12_), .S(
        add_2_root_r119_SUM_11_) );
  ADDFX2 U95 ( .A(in_17bit_b[10]), .B(in_17bit_b[8]), .CI(
        add_2_root_r115_carry_11_), .CO(add_2_root_r115_carry_12_), .S(
        add_2_root_r115_SUM_11_) );
  ADDFX2 U96 ( .A(in_17bit_b[12]), .B(in_17bit_b[8]), .CI(
        add_1_root_r112_carry_12_), .CO(add_1_root_r112_carry_13_), .S(
        add_1_root_r112_SUM_12_) );
  ADDFX2 U97 ( .A(in_17bit_b[9]), .B(in_17bit_b[7]), .CI(
        add_1_root_r115_carry_13_), .CO(add_1_root_r115_carry_14_), .S(
        add_1_root_r115_SUM_13_) );
  ADDFX2 U98 ( .A(in_17bit_b[13]), .B(in_17bit_b[12]), .CI(
        add_3_root_r119_carry_14_), .CO(add_3_root_r119_carry_15_), .S(
        add_1_root_r119_A_14_) );
  ADDFX2 U99 ( .A(add_1_root_r119_A_13_), .B(in_17bit_b[7]), .CI(
        add_1_root_r119_carry[13]), .CO(add_1_root_r119_carry[14]), .S(
        add_1_root_r119_SUM_13_) );
  ADDFX2 U100 ( .A(in_17bit_b[8]), .B(in_17bit_b[7]), .CI(
        add_2_root_r119_carry_12_), .CO(add_2_root_r119_carry_13_), .S(
        add_2_root_r119_SUM_12_) );
  ADDFX2 U101 ( .A(in_17bit_b[11]), .B(in_17bit_b[9]), .CI(
        add_2_root_r115_carry_12_), .CO(add_2_root_r115_carry_13_), .S(
        add_2_root_r115_SUM_12_) );
  ADDFX2 U102 ( .A(in_17bit_b[13]), .B(in_17bit_b[9]), .CI(
        add_1_root_r112_carry_13_), .CO(add_1_root_r112_carry_14_), .S(
        add_1_root_r112_SUM_13_) );
  ADDFX2 U103 ( .A(in_17bit_b[10]), .B(in_17bit_b[8]), .CI(
        add_1_root_r115_carry_14_), .CO(add_1_root_r115_carry_15_), .S(
        add_1_root_r115_SUM_14_) );
  ADDFX2 U104 ( .A(in_17bit_b[14]), .B(in_17bit_b[13]), .CI(
        add_3_root_r119_carry_15_), .CO(add_3_root_r119_carry_16_), .S(
        add_1_root_r119_A_15_) );
  ADDFX2 U105 ( .A(add_1_root_r119_A_14_), .B(in_17bit_b[8]), .CI(
        add_1_root_r119_carry[14]), .CO(add_1_root_r119_carry[15]), .S(
        add_1_root_r119_SUM_14_) );
  ADDFX2 U106 ( .A(in_17bit_b[9]), .B(in_17bit_b[8]), .CI(
        add_2_root_r119_carry_13_), .CO(add_2_root_r119_carry_14_), .S(
        add_2_root_r119_SUM_13_) );
  ADDFX2 U107 ( .A(in_17bit_b[12]), .B(in_17bit_b[10]), .CI(
        add_2_root_r115_carry_13_), .CO(add_2_root_r115_carry_14_), .S(
        add_2_root_r115_SUM_13_) );
  ADDFX2 U108 ( .A(in_17bit_b[14]), .B(in_17bit_b[10]), .CI(
        add_1_root_r112_carry_14_), .CO(add_1_root_r112_carry_15_), .S(
        add_1_root_r112_SUM_14_) );
  ADDFX2 U109 ( .A(in_17bit_b[11]), .B(in_17bit_b[9]), .CI(
        add_1_root_r115_carry_15_), .CO(add_1_root_r115_carry_16_), .S(
        add_1_root_r115_SUM_15_) );
  ADDFX2 U110 ( .A(add_1_root_r119_A_15_), .B(in_17bit_b[9]), .CI(
        add_1_root_r119_carry[15]), .CO(add_1_root_r119_carry[16]), .S(
        add_1_root_r119_SUM_15_) );
  ADDFX2 U111 ( .A(in_17bit_b[3]), .B(in_17bit_b[2]), .CI(
        add_3_root_r119_carry_4_), .CO(add_3_root_r119_carry_5_), .S(
        add_1_root_r119_A_4_) );
  ADDFX2 U112 ( .A(in_17bit_b[2]), .B(in_17bit_b[1]), .CI(
        add_3_root_r119_carry_3_), .CO(add_3_root_r119_carry_4_), .S(
        add_1_root_r119_A_3_) );
  ADDFX2 U113 ( .A(in_17bit_b[10]), .B(in_17bit_b[9]), .CI(
        add_2_root_r119_carry_14_), .CO(add_2_root_r119_carry_15_), .S(
        add_2_root_r119_SUM_14_) );
  ADDFX2 U114 ( .A(in_17bit_b[13]), .B(in_17bit_b[11]), .CI(
        add_2_root_r115_carry_14_), .CO(add_2_root_r115_carry_15_), .S(
        add_2_root_r115_SUM_14_) );
  ADDFX2 U115 ( .A(in_17bit_b[15]), .B(in_17bit_b[11]), .CI(
        add_1_root_r112_carry_15_), .CO(add_1_root_r112_carry_16_), .S(
        add_1_root_r112_SUM_15_) );
  ADDFX2 U116 ( .A(add_1_root_r119_A_16_), .B(in_17bit_b[10]), .CI(
        add_1_root_r119_carry[16]), .CO(add_1_root_r119_carry[17]), .S(
        add_1_root_r119_SUM_16_) );
  ADDFX2 U117 ( .A(in_17bit_b[11]), .B(in_17bit_b[10]), .CI(
        add_2_root_r119_carry_15_), .CO(add_2_root_r119_carry_16_), .S(
        add_2_root_r119_SUM_15_) );
  ADDFX2 U118 ( .A(in_17bit_b[14]), .B(in_17bit_b[12]), .CI(
        add_2_root_r115_carry_15_), .CO(add_2_root_r115_carry_16_), .S(
        add_2_root_r115_SUM_15_) );
  ADDFX2 U119 ( .A(in_17bit_b[13]), .B(in_17bit_b[11]), .CI(
        add_1_root_r115_carry_17_), .CO(add_1_root_r115_carry_18_), .S(
        add_1_root_r115_SUM_17_) );
  ADDFX2 U120 ( .A(add_1_root_r119_A_17_), .B(in_17bit_b[11]), .CI(
        add_1_root_r119_carry[17]), .CO(add_1_root_r119_carry[18]), .S(
        add_1_root_r119_SUM_17_) );
  ADDFX2 U121 ( .A(in_17bit_b[12]), .B(in_17bit_b[11]), .CI(
        add_2_root_r119_carry_16_), .CO(add_2_root_r119_carry_17_), .S(
        add_2_root_r119_SUM_16_) );
  ADDFX2 U122 ( .A(in_17bit_b[15]), .B(in_17bit_b[13]), .CI(
        add_2_root_r115_carry_16_), .CO(add_2_root_r115_carry_17_), .S(
        add_2_root_r115_SUM_16_) );
  ADDFX2 U123 ( .A(add_1_root_r119_A_18_), .B(in_17bit_b[12]), .CI(
        add_1_root_r119_carry[18]), .CO(add_1_root_r119_carry[19]), .S(
        add_1_root_r119_SUM_18_) );
  ADDFX2 U124 ( .A(in_17bit_b[13]), .B(in_17bit_b[12]), .CI(
        add_2_root_r119_carry_17_), .CO(add_2_root_r119_carry_18_), .S(
        add_2_root_r119_SUM_17_) );
  ADDFX2 U125 ( .A(in_17bit_b[5]), .B(in_17bit_b[3]), .CI(
        add_2_root_r115_carry_6_), .CO(add_2_root_r115_carry_7_), .S(
        add_2_root_r115_SUM_6_) );
  ADDFX2 U126 ( .A(in_17bit_b[7]), .B(in_17bit_b[3]), .CI(
        add_1_root_r112_carry_7_), .CO(add_1_root_r112_carry_8_), .S(
        add_1_root_r112_SUM_7_) );
  ADDFX2 U127 ( .A(add_1_root_r119_A_9_), .B(in_17bit_b[3]), .CI(
        add_1_root_r119_carry[9]), .CO(add_1_root_r119_carry[10]), .S(
        add_1_root_r119_SUM_9_) );
  ADDFX2 U128 ( .A(in_17bit_b[14]), .B(in_17bit_b[13]), .CI(
        add_2_root_r119_carry_18_), .CO(add_2_root_r119_carry_19_), .S(
        add_2_root_r119_SUM_18_) );
  ADDFX2 U129 ( .A(in_17bit_b[5]), .B(in_17bit_b[3]), .CI(
        add_1_root_r115_carry_9_), .CO(add_1_root_r115_carry_10_), .S(
        add_1_root_r115_SUM_9_) );
  ADDFX2 U130 ( .A(in_17bit_b[4]), .B(in_17bit_b[3]), .CI(
        add_2_root_r119_carry_8_), .CO(add_2_root_r119_carry_9_), .S(
        add_2_root_r119_SUM_8_) );
  ADDFX2 U131 ( .A(in_17bit_b[6]), .B(in_17bit_b[4]), .CI(
        add_1_root_r115_carry_10_), .CO(add_1_root_r115_carry_11_), .S(
        add_1_root_r115_SUM_10_) );
  ADDFX2 U132 ( .A(in_17bit_b[5]), .B(in_17bit_b[4]), .CI(
        add_2_root_r119_carry_9_), .CO(add_2_root_r119_carry_10_), .S(
        add_2_root_r119_SUM_9_) );
  ADDFX2 U133 ( .A(in_17bit_b[12]), .B(in_17bit_b[10]), .CI(
        add_1_root_r115_carry_16_), .CO(add_1_root_r115_carry_17_), .S(
        add_1_root_r115_SUM_16_) );
  ADDFX2 U134 ( .A(in_17bit_b[15]), .B(in_17bit_b[14]), .CI(
        add_3_root_r119_carry_16_), .CO(add_3_root_r119_carry_17_), .S(
        add_1_root_r119_A_16_) );
  ADDFX2 U135 ( .A(in_17bit_b[14]), .B(in_17bit_b[12]), .CI(
        add_1_root_r115_carry_18_), .CO(add_1_root_r115_carry_19_), .S(
        add_1_root_r115_SUM_18_) );
  ADDFX2 U136 ( .A(in_17bit_b[4]), .B(in_17bit_b[3]), .CI(
        add_3_root_r119_carry_5_), .CO(add_3_root_r119_carry_6_), .S(
        add_1_root_r119_A_5_) );
  ADDFX2 U137 ( .A(in_17bit_b[5]), .B(in_17bit_b[4]), .CI(
        add_3_root_r119_carry_6_), .CO(add_3_root_r119_carry_7_), .S(
        add_1_root_r119_A_6_) );
  ADDFX2 U138 ( .A(in_17bit_b[15]), .B(in_17bit_b[13]), .CI(
        add_1_root_r115_carry_19_), .CO(add_1_root_r115_carry_20_), .S(
        add_1_root_r115_SUM_19_) );
  ADDFX2 U139 ( .A(in_17bit_b[15]), .B(in_17bit_b[14]), .CI(
        add_2_root_r119_carry_19_), .CO(add_2_root_r119_carry_20_), .S(
        add_2_root_r119_SUM_19_) );
  INVX1 U140 ( .A(in_8bit[2]), .Y(n41) );
  INVX1 U141 ( .A(in_8bit[0]), .Y(n40) );
  NOR3X1 U142 ( .A(n41), .B(n201), .C(n40), .Y(n233) );
  CLKINVX3 U143 ( .A(n235), .Y(in_17bit_b[0]) );
  INVX1 U144 ( .A(n287), .Y(n198) );
  OAI21XL U145 ( .A0(n287), .A1(n288), .B0(n286), .Y(N463) );
  AOI22X1 U146 ( .A0(N221), .A1(n37), .B0(N363), .B1(n36), .Y(n286) );
  NAND2XL U147 ( .A(N29), .B(n22), .Y(n288) );
  CLKINVX3 U148 ( .A(n280), .Y(in_17bit_b[15]) );
  BUFX3 U149 ( .A(in_8bit[6]), .Y(n39) );
  BUFX3 U150 ( .A(in_8bit[1]), .Y(n38) );
  MXI2XL U151 ( .A(n6), .B(n15), .S0(n181), .Y(out[16]) );
  AOI32X1 U152 ( .A0(n233), .A1(n199), .A2(in_8bit[5]), .B0(n232), .B1(n231), 
        .Y(n287) );
  INVX1 U153 ( .A(n230), .Y(n199) );
  INVXL U154 ( .A(in_8bit[3]), .Y(n201) );
  NAND3BXL U155 ( .AN(in_8bit[5]), .B(n41), .C(in_8bit[3]), .Y(n224) );
  AOI22X1 U156 ( .A0(in_17bit[0]), .A1(n22), .B0(in_17bit[0]), .B1(n45), .Y(
        n235) );
  NOR4BX1 U157 ( .AN(n225), .B(n40), .C(n38), .D(in_8bit[2]), .Y(n231) );
  NOR2XL U158 ( .A(n39), .B(in_8bit[3]), .Y(n225) );
  AOI22X1 U159 ( .A0(N14), .A1(n22), .B0(in_17bit[1]), .B1(n45), .Y(n238) );
  AOI22X1 U160 ( .A0(N15), .A1(n22), .B0(in_17bit[2]), .B1(n45), .Y(n241) );
  AOI22X1 U161 ( .A0(N16), .A1(n22), .B0(in_17bit[3]), .B1(n45), .Y(n244) );
  AOI22X1 U162 ( .A0(N17), .A1(n22), .B0(in_17bit[4]), .B1(n45), .Y(n247) );
  AOI22X1 U163 ( .A0(N21), .A1(n22), .B0(in_17bit[8]), .B1(n45), .Y(n259) );
  NAND3X1 U164 ( .A(in_8bit[2]), .B(n201), .C(in_8bit[5]), .Y(n223) );
  AOI22XL U165 ( .A0(N26), .A1(n22), .B0(in_17bit[13]), .B1(n45), .Y(n274) );
  AOI22XL U166 ( .A0(N28), .A1(n22), .B0(in_17bit[15]), .B1(n45), .Y(n280) );
  AOI22XL U167 ( .A0(N18), .A1(n22), .B0(in_17bit[5]), .B1(n45), .Y(n250) );
  AOI22XL U168 ( .A0(N19), .A1(n22), .B0(in_17bit[6]), .B1(n45), .Y(n253) );
  AOI22XL U169 ( .A0(N20), .A1(n22), .B0(in_17bit[7]), .B1(n45), .Y(n256) );
  AOI22XL U170 ( .A0(N22), .A1(n22), .B0(in_17bit[9]), .B1(n45), .Y(n262) );
  AOI22XL U171 ( .A0(N23), .A1(n22), .B0(in_17bit[10]), .B1(n45), .Y(n265) );
  AOI22XL U172 ( .A0(N24), .A1(n22), .B0(in_17bit[11]), .B1(n45), .Y(n268) );
  AOI22XL U173 ( .A0(N25), .A1(n22), .B0(in_17bit[12]), .B1(n45), .Y(n271) );
  INVX1 U174 ( .A(n68), .Y(n72) );
  AND2X2 U175 ( .A(n29), .B(n4), .Y(n25) );
  AND2X2 U176 ( .A(n25), .B(n5), .Y(n26) );
  INVX1 U177 ( .A(n83), .Y(n80) );
  INVX1 U178 ( .A(n92), .Y(n89) );
  INVX1 U179 ( .A(n101), .Y(n98) );
  BUFX3 U180 ( .A(n284), .Y(n36) );
  OAI32X1 U181 ( .A0(n223), .A1(in_8bit[0]), .A2(n230), .B0(n224), .B1(n222), 
        .Y(n284) );
  BUFX3 U182 ( .A(n285), .Y(n37) );
  OAI32X1 U183 ( .A0(n230), .A1(in_8bit[0]), .A2(n224), .B0(n223), .B1(n222), 
        .Y(n285) );
  INVX1 U184 ( .A(n51), .Y(n55) );
  NAND2X1 U185 ( .A(n72), .B(n3), .Y(n74) );
  AND2X2 U186 ( .A(n26), .B(n7), .Y(n27) );
  INVX1 U187 ( .A(in_17bit[3]), .Y(n185) );
  INVX1 U188 ( .A(in_17bit[5]), .Y(n187) );
  INVX1 U189 ( .A(in_17bit[6]), .Y(n188) );
  INVX1 U190 ( .A(in_17bit[7]), .Y(n189) );
  INVX1 U191 ( .A(in_17bit[8]), .Y(n190) );
  INVX1 U192 ( .A(in_17bit[9]), .Y(n191) );
  INVX1 U193 ( .A(in_17bit[10]), .Y(n192) );
  INVX1 U194 ( .A(in_17bit[11]), .Y(n193) );
  INVX1 U195 ( .A(in_17bit[12]), .Y(n194) );
  INVX1 U196 ( .A(in_17bit[13]), .Y(n195) );
  INVX1 U197 ( .A(in_17bit[14]), .Y(n196) );
  INVX1 U198 ( .A(in_17bit[15]), .Y(n197) );
  INVX1 U199 ( .A(in_17bit[1]), .Y(n183) );
  INVX1 U200 ( .A(in_17bit[2]), .Y(n184) );
  INVX1 U201 ( .A(in_17bit[4]), .Y(n186) );
  INVX1 U202 ( .A(in_17bit[0]), .Y(n182) );
  NAND2X1 U203 ( .A(n237), .B(n236), .Y(N447) );
  AOI22X1 U204 ( .A0(N108), .A1(n281), .B0(N205), .B1(n37), .Y(n236) );
  AOI22X1 U205 ( .A0(N347), .A1(n36), .B0(n198), .B1(in_17bit_b[0]), .Y(n237)
         );
  NAND2X1 U206 ( .A(n240), .B(n239), .Y(N448) );
  AOI22X1 U207 ( .A0(N109), .A1(n281), .B0(N206), .B1(n37), .Y(n239) );
  AOI22X1 U208 ( .A0(N348), .A1(n36), .B0(n198), .B1(in_17bit_b[1]), .Y(n240)
         );
  NAND2X1 U209 ( .A(n243), .B(n242), .Y(N449) );
  AOI22X1 U210 ( .A0(N110), .A1(n281), .B0(N207), .B1(n37), .Y(n242) );
  AOI22X1 U211 ( .A0(N349), .A1(n36), .B0(n198), .B1(in_17bit_b[2]), .Y(n243)
         );
  NAND2X1 U212 ( .A(n246), .B(n245), .Y(N450) );
  AOI22X1 U213 ( .A0(N111), .A1(n281), .B0(N208), .B1(n37), .Y(n245) );
  AOI22X1 U214 ( .A0(N350), .A1(n36), .B0(n198), .B1(in_17bit_b[3]), .Y(n246)
         );
  NAND2X1 U215 ( .A(n249), .B(n248), .Y(N451) );
  AOI22X1 U216 ( .A0(N112), .A1(n281), .B0(N209), .B1(n37), .Y(n248) );
  AOI22X1 U217 ( .A0(N351), .A1(n36), .B0(n198), .B1(in_17bit_b[4]), .Y(n249)
         );
  NAND2X1 U218 ( .A(n252), .B(n251), .Y(N452) );
  AOI22X1 U219 ( .A0(N113), .A1(n281), .B0(N210), .B1(n37), .Y(n251) );
  AOI22X1 U220 ( .A0(N352), .A1(n36), .B0(n198), .B1(in_17bit_b[5]), .Y(n252)
         );
  NAND2X1 U221 ( .A(n255), .B(n254), .Y(N453) );
  AOI22X1 U222 ( .A0(N114), .A1(n281), .B0(N211), .B1(n37), .Y(n254) );
  AOI22X1 U223 ( .A0(N353), .A1(n36), .B0(n198), .B1(in_17bit_b[6]), .Y(n255)
         );
  NAND2X1 U224 ( .A(n258), .B(n257), .Y(N454) );
  AOI22X1 U225 ( .A0(N115), .A1(n281), .B0(N212), .B1(n37), .Y(n257) );
  AOI22X1 U226 ( .A0(N354), .A1(n36), .B0(n198), .B1(in_17bit_b[7]), .Y(n258)
         );
  NAND2X1 U227 ( .A(n261), .B(n260), .Y(N455) );
  AOI22X1 U228 ( .A0(N116), .A1(n281), .B0(N213), .B1(n37), .Y(n260) );
  AOI22X1 U229 ( .A0(N355), .A1(n36), .B0(n198), .B1(in_17bit_b[8]), .Y(n261)
         );
  NAND2X1 U230 ( .A(n264), .B(n263), .Y(N456) );
  AOI22X1 U231 ( .A0(N117), .A1(n281), .B0(N214), .B1(n37), .Y(n263) );
  AOI22X1 U232 ( .A0(N356), .A1(n36), .B0(n198), .B1(in_17bit_b[9]), .Y(n264)
         );
  NAND2X1 U233 ( .A(n267), .B(n266), .Y(N457) );
  AOI22X1 U234 ( .A0(N118), .A1(n281), .B0(N215), .B1(n37), .Y(n266) );
  AOI22X1 U235 ( .A0(N357), .A1(n36), .B0(n198), .B1(in_17bit_b[10]), .Y(n267)
         );
  NAND2X1 U236 ( .A(n270), .B(n269), .Y(N458) );
  AOI22X1 U237 ( .A0(N119), .A1(n281), .B0(N216), .B1(n37), .Y(n269) );
  AOI22X1 U238 ( .A0(N358), .A1(n36), .B0(n198), .B1(in_17bit_b[11]), .Y(n270)
         );
  NAND2X1 U239 ( .A(n273), .B(n272), .Y(N459) );
  AOI22X1 U240 ( .A0(N120), .A1(n281), .B0(N217), .B1(n37), .Y(n272) );
  AOI22X1 U241 ( .A0(N359), .A1(n36), .B0(n198), .B1(in_17bit_b[12]), .Y(n273)
         );
  NAND2X1 U242 ( .A(n276), .B(n275), .Y(N460) );
  AOI22X1 U243 ( .A0(N121), .A1(n281), .B0(N218), .B1(n37), .Y(n275) );
  AOI22X1 U244 ( .A0(N360), .A1(n36), .B0(n198), .B1(in_17bit_b[13]), .Y(n276)
         );
  NAND2X1 U245 ( .A(n279), .B(n278), .Y(N461) );
  AOI22X1 U246 ( .A0(N122), .A1(n281), .B0(N219), .B1(n37), .Y(n278) );
  AOI22X1 U247 ( .A0(N361), .A1(n36), .B0(n198), .B1(in_17bit_b[14]), .Y(n279)
         );
  NAND2X1 U248 ( .A(n283), .B(n282), .Y(N462) );
  AOI22X1 U249 ( .A0(N123), .A1(n281), .B0(N220), .B1(n37), .Y(n282) );
  AOI22X1 U250 ( .A0(N362), .A1(n36), .B0(n198), .B1(in_17bit_b[15]), .Y(n283)
         );
  OAI21XL U251 ( .A0(in_8bit[7]), .A1(n76), .B0(n75), .Y(n82) );
  NAND2BX1 U252 ( .AN(neg_mul[12]), .B(in_8bit[7]), .Y(n75) );
  OAI21XL U253 ( .A0(in_8bit[7]), .A1(n94), .B0(n93), .Y(n100) );
  NAND2BX1 U254 ( .AN(neg_mul[14]), .B(in_8bit[7]), .Y(n93) );
  XNOR2X1 U255 ( .A(n11), .B(sub_add_75_b0_carry[13]), .Y(n28) );
  OAI21XL U256 ( .A0(in_8bit[7]), .A1(n57), .B0(n56), .Y(n62) );
  NAND2BX1 U257 ( .AN(neg_mul[9]), .B(in_8bit[7]), .Y(n56) );
  OAI21XL U258 ( .A0(in_8bit[7]), .A1(n48), .B0(n47), .Y(n54) );
  NAND2BX1 U259 ( .AN(neg_mul[8]), .B(in_8bit[7]), .Y(n47) );
  OAI21XL U260 ( .A0(in_8bit[7]), .A1(n65), .B0(n64), .Y(n70) );
  NAND2BX1 U261 ( .AN(neg_mul[10]), .B(in_8bit[7]), .Y(n64) );
  OAI21XL U262 ( .A0(in_8bit[7]), .A1(n171), .B0(n170), .Y(n176) );
  NAND2BX1 U263 ( .AN(neg_mul[15]), .B(in_8bit[7]), .Y(n170) );
  OAI21XL U264 ( .A0(in_8bit[7]), .A1(n85), .B0(n84), .Y(n91) );
  NAND2BX1 U265 ( .AN(neg_mul[13]), .B(in_8bit[7]), .Y(n84) );
  MX2X1 U266 ( .A(neg_mul[22]), .B(N480), .S0(n181), .Y(out[15]) );
  NAND4BBX1 U267 ( .AN(n36), .BN(n37), .C(n234), .D(n287), .Y(N446) );
  AOI2BB1X1 U268 ( .A0N(n229), .A1N(n228), .B0(n281), .Y(n234) );
  OR4X2 U269 ( .A(in_8bit[4]), .B(in_8bit[5]), .C(n39), .D(in_8bit[7]), .Y(
        n229) );
  OR4XL U270 ( .A(n38), .B(in_8bit[0]), .C(in_8bit[2]), .D(in_8bit[3]), .Y(
        n228) );
  NOR3X1 U271 ( .A(in_8bit[4]), .B(in_8bit[5]), .C(n200), .Y(n232) );
  NAND4X1 U272 ( .A(n39), .B(in_8bit[4]), .C(n38), .D(n200), .Y(n230) );
  NOR2BX1 U273 ( .AN(n98), .B(neg_mul[15]), .Y(n29) );
  NAND4X1 U274 ( .A(n38), .B(in_8bit[7]), .C(n221), .D(n40), .Y(n222) );
  NOR2X1 U275 ( .A(n39), .B(in_8bit[4]), .Y(n221) );
  NAND2X1 U276 ( .A(n55), .B(n14), .Y(n63) );
  NAND2X1 U277 ( .A(out[0]), .B(neg_mul[8]), .Y(n48) );
  NAND2X1 U278 ( .A(neg_mul[10]), .B(n63), .Y(n65) );
  NAND2X1 U279 ( .A(neg_mul[12]), .B(n74), .Y(n76) );
  NAND2X1 U280 ( .A(neg_mul[14]), .B(n92), .Y(n94) );
  AOI21X1 U281 ( .A0(n59), .A1(in_8bit[7]), .B0(n58), .Y(n60) );
  INVX1 U282 ( .A(n57), .Y(n59) );
  NOR2X1 U283 ( .A(in_8bit[7]), .B(neg_mul[9]), .Y(n58) );
  NAND2BX1 U284 ( .AN(n55), .B(neg_mul[9]), .Y(n57) );
  AOI21X1 U285 ( .A0(n173), .A1(in_8bit[7]), .B0(n172), .Y(n174) );
  INVX1 U286 ( .A(n171), .Y(n173) );
  NOR2X1 U287 ( .A(in_8bit[7]), .B(neg_mul[15]), .Y(n172) );
  AOI21X1 U288 ( .A0(n87), .A1(in_8bit[7]), .B0(n86), .Y(n88) );
  INVX1 U289 ( .A(n85), .Y(n87) );
  NOR2X1 U290 ( .A(in_8bit[7]), .B(neg_mul[13]), .Y(n86) );
  NAND2X1 U291 ( .A(n227), .B(n226), .Y(n281) );
  NAND4X1 U292 ( .A(n232), .B(n233), .C(n39), .D(n38), .Y(n226) );
  NAND4X1 U293 ( .A(n231), .B(in_8bit[5]), .C(in_8bit[4]), .D(n200), .Y(n227)
         );
  NAND2X1 U294 ( .A(neg_mul[15]), .B(n101), .Y(n171) );
  NAND2X1 U295 ( .A(neg_mul[13]), .B(n83), .Y(n85) );
  OR2X2 U296 ( .A(n63), .B(neg_mul[10]), .Y(n68) );
  OR2X2 U297 ( .A(n74), .B(neg_mul[12]), .Y(n83) );
  NAND2X1 U298 ( .A(n80), .B(n12), .Y(n92) );
  NAND2X1 U299 ( .A(n89), .B(n13), .Y(n101) );
  NOR2X1 U300 ( .A(n50), .B(n49), .Y(n52) );
  NOR2X1 U301 ( .A(in_8bit[7]), .B(neg_mul[8]), .Y(n49) );
  NOR2X1 U302 ( .A(n200), .B(n48), .Y(n50) );
  NOR2X1 U303 ( .A(in_8bit[7]), .B(neg_mul[10]), .Y(n66) );
  NOR2X1 U304 ( .A(n200), .B(n65), .Y(n67) );
  NOR2X1 U305 ( .A(n78), .B(n77), .Y(n79) );
  NOR2X1 U306 ( .A(in_8bit[7]), .B(neg_mul[12]), .Y(n77) );
  NOR2X1 U307 ( .A(n200), .B(n76), .Y(n78) );
  NOR2X1 U308 ( .A(n96), .B(n95), .Y(n97) );
  NOR2X1 U309 ( .A(in_8bit[7]), .B(neg_mul[14]), .Y(n95) );
  NOR2X1 U310 ( .A(n200), .B(n94), .Y(n96) );
  OR2X2 U311 ( .A(out[0]), .B(neg_mul[8]), .Y(n51) );
  NAND2X1 U312 ( .A(sub_add_75_b0_carry[15]), .B(n9), .Y(n30) );
  INVX1 U313 ( .A(in_8bit[7]), .Y(n200) );
  AOI21X4 U314 ( .A0(n42), .A1(n54), .B0(n53), .Y(out[1]) );
  OAI21X4 U315 ( .A0(n44), .A1(n60), .B0(n63), .Y(n61) );
  AOI21X4 U316 ( .A0(n42), .A1(n62), .B0(n61), .Y(out[2]) );
  AOI21X4 U317 ( .A0(n43), .A1(n70), .B0(n69), .Y(out[3]) );
  XNOR2X4 U318 ( .A(n44), .B(in_8bit[7]), .Y(n71) );
  MXI2X4 U319 ( .A(n11), .B(n28), .S0(n181), .Y(out[13]) );
  AND2X1 U320 ( .A(add_1_root_r112_carry_20_), .B(in_17bit_b[16]), .Y(
        add_1_root_r112_SUM_21_) );
  XOR2X1 U321 ( .A(in_17bit_b[16]), .B(add_1_root_r112_carry_20_), .Y(
        add_1_root_r112_SUM_20_) );
  AND2X1 U322 ( .A(add_1_root_r112_carry_19_), .B(in_17bit_b[15]), .Y(
        add_1_root_r112_carry_20_) );
  XOR2X1 U323 ( .A(in_17bit_b[15]), .B(add_1_root_r112_carry_19_), .Y(
        add_1_root_r112_SUM_19_) );
  AND2X1 U324 ( .A(add_1_root_r112_carry_18_), .B(in_17bit_b[14]), .Y(
        add_1_root_r112_carry_19_) );
  XOR2X1 U325 ( .A(in_17bit_b[14]), .B(add_1_root_r112_carry_18_), .Y(
        add_1_root_r112_SUM_18_) );
  AND2X1 U326 ( .A(add_1_root_r112_carry_17_), .B(in_17bit_b[13]), .Y(
        add_1_root_r112_carry_18_) );
  XOR2X1 U327 ( .A(in_17bit_b[13]), .B(add_1_root_r112_carry_17_), .Y(
        add_1_root_r112_SUM_17_) );
  AND2X1 U328 ( .A(add_2_root_r119_carry_21_), .B(in_17bit_b[16]), .Y(
        add_2_root_r119_SUM_22_) );
  XOR2X1 U329 ( .A(in_17bit_b[16]), .B(add_2_root_r119_carry_21_), .Y(
        add_2_root_r119_SUM_21_) );
  AND2X1 U330 ( .A(add_1_root_r119_carry[22]), .B(in_17bit_b[16]), .Y(
        add_1_root_r119_SUM_23_) );
  XOR2X1 U331 ( .A(in_17bit_b[16]), .B(add_1_root_r119_carry[22]), .Y(
        add_1_root_r119_SUM_22_) );
  AND2X1 U332 ( .A(add_1_root_r119_carry[21]), .B(in_17bit_b[15]), .Y(
        add_1_root_r119_carry[22]) );
  XOR2X1 U333 ( .A(in_17bit_b[15]), .B(add_1_root_r119_carry[21]), .Y(
        add_1_root_r119_SUM_21_) );
  AND2X1 U334 ( .A(add_1_root_r119_carry[20]), .B(in_17bit_b[14]), .Y(
        add_1_root_r119_carry[21]) );
  XOR2X1 U335 ( .A(in_17bit_b[14]), .B(add_1_root_r119_carry[20]), .Y(
        add_1_root_r119_SUM_20_) );
  AND2X1 U336 ( .A(add_1_root_r119_A_6_), .B(in_17bit_b[0]), .Y(
        add_1_root_r119_carry[7]) );
  XOR2X1 U337 ( .A(in_17bit_b[0]), .B(add_1_root_r119_A_6_), .Y(
        add_1_root_r119_SUM_6_) );
  AND2X1 U338 ( .A(add_3_root_r119_carry_18_), .B(in_17bit_b[16]), .Y(
        add_1_root_r119_A_19_) );
  XOR2X1 U339 ( .A(in_17bit_b[16]), .B(add_3_root_r119_carry_18_), .Y(
        add_1_root_r119_A_18_) );
  AND2X1 U340 ( .A(in_17bit_b[1]), .B(in_17bit_b[0]), .Y(
        add_3_root_r119_carry_3_) );
  XOR2X1 U341 ( .A(in_17bit_b[0]), .B(in_17bit_b[1]), .Y(add_1_root_r119_A_2_)
         );
  AND2X1 U342 ( .A(add_2_root_r115_carry_19_), .B(in_17bit_b[16]), .Y(
        add_2_root_r115_SUM_20_) );
  XOR2X1 U343 ( .A(in_17bit_b[16]), .B(add_2_root_r115_carry_19_), .Y(
        add_2_root_r115_SUM_19_) );
  AND2X1 U344 ( .A(add_2_root_r115_carry_18_), .B(in_17bit_b[15]), .Y(
        add_2_root_r115_carry_19_) );
  XOR2X1 U345 ( .A(in_17bit_b[15]), .B(add_2_root_r115_carry_18_), .Y(
        add_2_root_r115_SUM_18_) );
  AND2X1 U346 ( .A(add_1_root_r115_carry_22_), .B(in_17bit_b[16]), .Y(
        add_1_root_r115_SUM_23_) );
  XOR2X1 U347 ( .A(in_17bit_b[16]), .B(add_1_root_r115_carry_22_), .Y(
        add_1_root_r115_SUM_22_) );
  AND2X1 U348 ( .A(add_1_root_r115_carry_21_), .B(in_17bit_b[15]), .Y(
        add_1_root_r115_carry_22_) );
  XOR2X1 U349 ( .A(in_17bit_b[15]), .B(add_1_root_r115_carry_21_), .Y(
        add_1_root_r115_SUM_21_) );
  AND2X1 U350 ( .A(in_17bit_b[2]), .B(in_17bit_b[0]), .Y(
        add_1_root_r115_carry_7_) );
  XOR2X1 U351 ( .A(in_17bit_b[0]), .B(in_17bit_b[2]), .Y(
        add_1_root_r115_SUM_6_) );
  XOR2X1 U352 ( .A(n45), .B(sub_add_54_b0_carry[16]), .Y(N29) );
  AND2X1 U353 ( .A(sub_add_54_b0_carry[15]), .B(n197), .Y(
        sub_add_54_b0_carry[16]) );
  XOR2X1 U354 ( .A(n197), .B(sub_add_54_b0_carry[15]), .Y(N28) );
  AND2X1 U355 ( .A(sub_add_54_b0_carry[14]), .B(n196), .Y(
        sub_add_54_b0_carry[15]) );
  XOR2X1 U356 ( .A(n196), .B(sub_add_54_b0_carry[14]), .Y(N27) );
  AND2X1 U357 ( .A(sub_add_54_b0_carry[13]), .B(n195), .Y(
        sub_add_54_b0_carry[14]) );
  XOR2X1 U358 ( .A(n195), .B(sub_add_54_b0_carry[13]), .Y(N26) );
  AND2X1 U359 ( .A(sub_add_54_b0_carry[12]), .B(n194), .Y(
        sub_add_54_b0_carry[13]) );
  XOR2X1 U360 ( .A(n194), .B(sub_add_54_b0_carry[12]), .Y(N25) );
  AND2X1 U361 ( .A(sub_add_54_b0_carry[11]), .B(n193), .Y(
        sub_add_54_b0_carry[12]) );
  XOR2X1 U362 ( .A(n193), .B(sub_add_54_b0_carry[11]), .Y(N24) );
  AND2X1 U363 ( .A(sub_add_54_b0_carry[10]), .B(n192), .Y(
        sub_add_54_b0_carry[11]) );
  XOR2X1 U364 ( .A(n192), .B(sub_add_54_b0_carry[10]), .Y(N23) );
  AND2X1 U365 ( .A(sub_add_54_b0_carry[9]), .B(n191), .Y(
        sub_add_54_b0_carry[10]) );
  XOR2X1 U366 ( .A(n191), .B(sub_add_54_b0_carry[9]), .Y(N22) );
  AND2X1 U367 ( .A(sub_add_54_b0_carry[8]), .B(n190), .Y(
        sub_add_54_b0_carry[9]) );
  XOR2X1 U368 ( .A(n190), .B(sub_add_54_b0_carry[8]), .Y(N21) );
  AND2X1 U369 ( .A(sub_add_54_b0_carry[7]), .B(n189), .Y(
        sub_add_54_b0_carry[8]) );
  XOR2X1 U370 ( .A(n189), .B(sub_add_54_b0_carry[7]), .Y(N20) );
  AND2X1 U371 ( .A(sub_add_54_b0_carry[6]), .B(n188), .Y(
        sub_add_54_b0_carry[7]) );
  XOR2X1 U372 ( .A(n188), .B(sub_add_54_b0_carry[6]), .Y(N19) );
  AND2X1 U373 ( .A(sub_add_54_b0_carry[5]), .B(n187), .Y(
        sub_add_54_b0_carry[6]) );
  XOR2X1 U374 ( .A(n187), .B(sub_add_54_b0_carry[5]), .Y(N18) );
  AND2X1 U375 ( .A(sub_add_54_b0_carry[4]), .B(n186), .Y(
        sub_add_54_b0_carry[5]) );
  XOR2X1 U376 ( .A(n186), .B(sub_add_54_b0_carry[4]), .Y(N17) );
  AND2X1 U377 ( .A(sub_add_54_b0_carry[3]), .B(n185), .Y(
        sub_add_54_b0_carry[4]) );
  XOR2X1 U378 ( .A(n185), .B(sub_add_54_b0_carry[3]), .Y(N16) );
  AND2X1 U379 ( .A(sub_add_54_b0_carry[2]), .B(n184), .Y(
        sub_add_54_b0_carry[3]) );
  XOR2X1 U380 ( .A(n184), .B(sub_add_54_b0_carry[2]), .Y(N15) );
  AND2X1 U381 ( .A(n182), .B(n183), .Y(sub_add_54_b0_carry[2]) );
  XOR2X1 U382 ( .A(n183), .B(n182), .Y(N14) );
  XOR2X1 U383 ( .A(n9), .B(sub_add_75_b0_carry[15]), .Y(N480) );
  AND2X1 U384 ( .A(sub_add_75_b0_carry[14]), .B(n10), .Y(
        sub_add_75_b0_carry[15]) );
  XOR2X1 U385 ( .A(n10), .B(sub_add_75_b0_carry[14]), .Y(N479) );
  AND2X1 U386 ( .A(sub_add_75_b0_carry[13]), .B(n11), .Y(
        sub_add_75_b0_carry[14]) );
  AND2X1 U387 ( .A(n27), .B(n8), .Y(sub_add_75_b0_carry[13]) );
  AND2X1 U388 ( .A(in_17bit_b[0]), .B(in_17bit_b[4]), .Y(
        add_1_root_r112_carry_5_) );
endmodule


module multi16_8_DW01_add_0 ( A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, 
        A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, 
        A_4_, B_23_, B_22_, B_21_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, 
        B_14_, B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, 
        SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, 
        SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, 
        SUM_7_ );
  input A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_,
         A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, B_23_, B_22_,
         B_21_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_,
         B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_;
  output SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_,
         SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_,
         SUM_8_, SUM_7_;
  wire   n1, n2, n3, n4;
  wire   [23:7] carry;

  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry[7]), .CO(carry[8]), .S(SUM_7_)
         );
  ADDFX2 U1_21 ( .A(A_21_), .B(B_21_), .CI(carry[21]), .CO(carry[22]), .S(
        SUM_21_) );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry[20]), .CO(carry[21]), .S(
        SUM_20_) );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry[19]), .CO(carry[20]), .S(
        SUM_19_) );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry[18]), .CO(carry[19]), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry[17]), .CO(carry[18]), .S(
        SUM_17_) );
  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry[16]), .CO(carry[17]), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry[15]), .CO(carry[16]), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry[14]), .CO(carry[15]), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry[13]), .CO(carry[14]), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry[12]), .CO(carry[13]), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry[11]), .CO(carry[12]), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry[10]), .CO(carry[11]), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry[9]), .CO(carry[10]), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry[8]), .CO(carry[9]), .S(SUM_8_)
         );
  ADDFX2 U1_22 ( .A(A_22_), .B(B_22_), .CI(carry[22]), .CO(carry[23]), .S(
        SUM_22_) );
  AND2X2 U1 ( .A(A_4_), .B(B_4_), .Y(n1) );
  XOR2X1 U2 ( .A(B_23_), .B(carry[23]), .Y(SUM_23_) );
  OAI2BB1X1 U3 ( .A0N(n2), .A1N(A_6_), .B0(n3), .Y(carry[7]) );
  OAI21XL U4 ( .A0(A_6_), .A1(n2), .B0(B_6_), .Y(n3) );
  OAI2BB1X1 U5 ( .A0N(n1), .A1N(A_5_), .B0(n4), .Y(n2) );
  OAI21XL U6 ( .A0(A_5_), .A1(n1), .B0(B_5_), .Y(n4) );
endmodule


module multi16_8_DW01_add_4 ( A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, 
        A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, 
        B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, 
        B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, SUM_22_, SUM_21_, SUM_20_, 
        SUM_19_, SUM_18_, SUM_17_, SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, 
        SUM_11_, SUM_10_, SUM_9_, SUM_8_, SUM_7_ );
  input A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_,
         A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, B_20_, B_19_,
         B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, B_10_, B_9_,
         B_8_, B_7_, B_6_, B_5_;
  output SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_,
         SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_,
         SUM_7_;
  wire   carry_21_, carry_20_, carry_19_, carry_18_, carry_17_, carry_16_,
         carry_15_, carry_14_, carry_13_, carry_12_, carry_11_, carry_10_,
         carry_9_, carry_8_, carry_7_, n1;

  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry_16_), .CO(carry_17_), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry_15_), .CO(carry_16_), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry_14_), .CO(carry_15_), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry_13_), .CO(carry_14_), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry_12_), .CO(carry_13_), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry_11_), .CO(carry_12_), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry_10_), .CO(carry_11_), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry_9_), .CO(carry_10_), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry_8_), .CO(carry_9_), .S(SUM_8_)
         );
  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry_7_), .CO(carry_8_), .S(SUM_7_)
         );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry_20_), .CO(carry_21_), .S(
        SUM_20_) );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry_19_), .CO(carry_20_), .S(
        SUM_19_) );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry_18_), .CO(carry_19_), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry_17_), .CO(carry_18_), .S(
        SUM_17_) );
  ADDFX2 U1_21 ( .A(A_21_), .B(B_21_), .CI(carry_21_), .CO(SUM_22_), .S(
        SUM_21_) );
  OAI2BB1X1 U1 ( .A0N(A_6_), .A1N(B_6_), .B0(n1), .Y(carry_7_) );
  OAI211X1 U2 ( .A0(B_6_), .A1(A_6_), .B0(A_5_), .C0(B_5_), .Y(n1) );
endmodule


module multi16_8_DW01_add_6 ( A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, 
        A_16_, A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, 
        A_6_, A_5_, A_4_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, 
        B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, 
        SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, 
        SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, 
        SUM_7_ );
  input A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_,
         A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, B_20_,
         B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, B_10_,
         B_9_, B_8_, B_7_, B_6_, B_5_, B_4_;
  output SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_,
         SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_,
         SUM_8_, SUM_7_;
  wire   n1, n2, n3, n4, n5, n6;
  wire   [21:7] carry;

  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry[7]), .CO(carry[8]), .S(SUM_7_)
         );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry[18]), .CO(carry[19]), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry[17]), .CO(carry[18]), .S(
        SUM_17_) );
  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry[16]), .CO(carry[17]), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry[15]), .CO(carry[16]), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry[14]), .CO(carry[15]), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry[13]), .CO(carry[14]), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry[12]), .CO(carry[13]), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry[11]), .CO(carry[12]), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry[10]), .CO(carry[11]), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry[9]), .CO(carry[10]), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry[8]), .CO(carry[9]), .S(SUM_8_)
         );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry[19]), .CO(carry[20]), .S(
        SUM_19_) );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry[20]), .CO(carry[21]), .S(
        SUM_20_) );
  AND2X2 U1 ( .A(A_22_), .B(n2), .Y(n1) );
  AND2X2 U2 ( .A(A_21_), .B(carry[21]), .Y(n2) );
  XOR2X1 U3 ( .A(A_23_), .B(n1), .Y(SUM_23_) );
  AND2X2 U4 ( .A(A_4_), .B(B_4_), .Y(n3) );
  XOR2X1 U5 ( .A(A_21_), .B(carry[21]), .Y(SUM_21_) );
  XOR2X1 U6 ( .A(A_22_), .B(n2), .Y(SUM_22_) );
  OAI2BB1X1 U7 ( .A0N(n4), .A1N(A_6_), .B0(n5), .Y(carry[7]) );
  OAI21XL U8 ( .A0(A_6_), .A1(n4), .B0(B_6_), .Y(n5) );
  OAI2BB1X1 U9 ( .A0N(n3), .A1N(A_5_), .B0(n6), .Y(n4) );
  OAI21XL U10 ( .A0(A_5_), .A1(n3), .B0(B_5_), .Y(n6) );
endmodule


module multi16_8 ( in_17bit, in_8bit, out );
  input [16:0] in_17bit;
  input [7:0] in_8bit;
  output [16:0] out;
  wire   n291, n292, n293, n294, n295, n296, N14, N15, N16, N17, N18, N19, N20,
         N21, N22, N23, N24, N25, N26, N27, N28, N29, N108, N109, N110, N111,
         N112, N113, N114, N115, N116, N117, N118, N119, N120, N121, N122,
         N123, N205, N206, N207, N208, N209, N210, N211, N212, N213, N214,
         N215, N216, N217, N218, N219, N220, N221, N347, N348, N349, N350,
         N351, N352, N353, N354, N355, N356, N357, N358, N359, N360, N361,
         N362, N363, N446, N447, N448, N449, N450, N451, N452, N453, N454,
         N455, N456, N457, N458, N459, N460, N461, N462, N463, N480, N481,
         add_2_root_r119_carry_10_, add_2_root_r119_carry_11_,
         add_2_root_r119_carry_12_, add_2_root_r119_carry_13_,
         add_2_root_r119_carry_14_, add_2_root_r119_carry_15_,
         add_2_root_r119_carry_16_, add_2_root_r119_carry_17_,
         add_2_root_r119_carry_18_, add_2_root_r119_carry_19_,
         add_2_root_r119_carry_20_, add_2_root_r119_carry_21_,
         add_2_root_r119_carry_7_, add_2_root_r119_carry_8_,
         add_2_root_r119_carry_9_, add_2_root_r119_SUM_6_,
         add_2_root_r119_SUM_7_, add_2_root_r119_SUM_8_,
         add_2_root_r119_SUM_9_, add_2_root_r119_SUM_10_,
         add_2_root_r119_SUM_11_, add_2_root_r119_SUM_12_,
         add_2_root_r119_SUM_13_, add_2_root_r119_SUM_14_,
         add_2_root_r119_SUM_15_, add_2_root_r119_SUM_16_,
         add_2_root_r119_SUM_17_, add_2_root_r119_SUM_18_,
         add_2_root_r119_SUM_19_, add_2_root_r119_SUM_20_,
         add_2_root_r119_SUM_21_, add_2_root_r119_SUM_22_,
         add_1_root_r119_SUM_6_, add_1_root_r119_SUM_7_,
         add_1_root_r119_SUM_8_, add_1_root_r119_SUM_9_,
         add_1_root_r119_SUM_10_, add_1_root_r119_SUM_11_,
         add_1_root_r119_SUM_12_, add_1_root_r119_SUM_13_,
         add_1_root_r119_SUM_14_, add_1_root_r119_SUM_15_,
         add_1_root_r119_SUM_16_, add_1_root_r119_SUM_17_,
         add_1_root_r119_SUM_18_, add_1_root_r119_SUM_19_,
         add_1_root_r119_SUM_20_, add_1_root_r119_SUM_21_,
         add_1_root_r119_SUM_22_, add_1_root_r119_SUM_23_,
         add_1_root_r119_A_2_, add_1_root_r119_A_3_, add_1_root_r119_A_4_,
         add_1_root_r119_A_5_, add_1_root_r119_A_6_, add_1_root_r119_A_7_,
         add_1_root_r119_A_8_, add_1_root_r119_A_9_, add_1_root_r119_A_10_,
         add_1_root_r119_A_11_, add_1_root_r119_A_12_, add_1_root_r119_A_13_,
         add_1_root_r119_A_14_, add_1_root_r119_A_15_, add_1_root_r119_A_16_,
         add_1_root_r119_A_17_, add_1_root_r119_A_18_, add_1_root_r119_A_19_,
         add_3_root_r119_carry_10_, add_3_root_r119_carry_11_,
         add_3_root_r119_carry_12_, add_3_root_r119_carry_13_,
         add_3_root_r119_carry_14_, add_3_root_r119_carry_15_,
         add_3_root_r119_carry_16_, add_3_root_r119_carry_17_,
         add_3_root_r119_carry_18_, add_3_root_r119_carry_3_,
         add_3_root_r119_carry_4_, add_3_root_r119_carry_5_,
         add_3_root_r119_carry_6_, add_3_root_r119_carry_7_,
         add_3_root_r119_carry_8_, add_3_root_r119_carry_9_,
         add_1_root_r112_carry_10_, add_1_root_r112_carry_11_,
         add_1_root_r112_carry_12_, add_1_root_r112_carry_13_,
         add_1_root_r112_carry_14_, add_1_root_r112_carry_15_,
         add_1_root_r112_carry_16_, add_1_root_r112_carry_17_,
         add_1_root_r112_carry_18_, add_1_root_r112_carry_19_,
         add_1_root_r112_carry_20_, add_1_root_r112_carry_5_,
         add_1_root_r112_carry_6_, add_1_root_r112_carry_7_,
         add_1_root_r112_carry_8_, add_1_root_r112_carry_9_,
         add_1_root_r112_SUM_1_, add_1_root_r112_SUM_2_,
         add_1_root_r112_SUM_3_, add_1_root_r112_SUM_4_,
         add_1_root_r112_SUM_5_, add_1_root_r112_SUM_6_,
         add_1_root_r112_SUM_7_, add_1_root_r112_SUM_8_,
         add_1_root_r112_SUM_9_, add_1_root_r112_SUM_10_,
         add_1_root_r112_SUM_11_, add_1_root_r112_SUM_12_,
         add_1_root_r112_SUM_13_, add_1_root_r112_SUM_14_,
         add_1_root_r112_SUM_15_, add_1_root_r112_SUM_16_,
         add_1_root_r112_SUM_17_, add_1_root_r112_SUM_18_,
         add_1_root_r112_SUM_19_, add_1_root_r112_SUM_20_,
         add_1_root_r112_SUM_21_, add_2_root_r115_carry_10_,
         add_2_root_r115_carry_11_, add_2_root_r115_carry_12_,
         add_2_root_r115_carry_13_, add_2_root_r115_carry_14_,
         add_2_root_r115_carry_15_, add_2_root_r115_carry_16_,
         add_2_root_r115_carry_17_, add_2_root_r115_carry_18_,
         add_2_root_r115_carry_19_, add_2_root_r115_carry_4_,
         add_2_root_r115_carry_5_, add_2_root_r115_carry_6_,
         add_2_root_r115_carry_7_, add_2_root_r115_carry_8_,
         add_2_root_r115_carry_9_, add_2_root_r115_SUM_3_,
         add_2_root_r115_SUM_4_, add_2_root_r115_SUM_5_,
         add_2_root_r115_SUM_6_, add_2_root_r115_SUM_7_,
         add_2_root_r115_SUM_8_, add_2_root_r115_SUM_9_,
         add_2_root_r115_SUM_10_, add_2_root_r115_SUM_11_,
         add_2_root_r115_SUM_12_, add_2_root_r115_SUM_13_,
         add_2_root_r115_SUM_14_, add_2_root_r115_SUM_15_,
         add_2_root_r115_SUM_16_, add_2_root_r115_SUM_17_,
         add_2_root_r115_SUM_18_, add_2_root_r115_SUM_19_,
         add_2_root_r115_SUM_20_, add_1_root_r115_carry_10_,
         add_1_root_r115_carry_11_, add_1_root_r115_carry_12_,
         add_1_root_r115_carry_13_, add_1_root_r115_carry_14_,
         add_1_root_r115_carry_15_, add_1_root_r115_carry_16_,
         add_1_root_r115_carry_17_, add_1_root_r115_carry_18_,
         add_1_root_r115_carry_19_, add_1_root_r115_carry_20_,
         add_1_root_r115_carry_21_, add_1_root_r115_carry_22_,
         add_1_root_r115_carry_8_, add_1_root_r115_carry_9_,
         add_1_root_r115_SUM_7_, add_1_root_r115_SUM_8_,
         add_1_root_r115_SUM_9_, add_1_root_r115_SUM_10_,
         add_1_root_r115_SUM_11_, add_1_root_r115_SUM_12_,
         add_1_root_r115_SUM_13_, add_1_root_r115_SUM_14_,
         add_1_root_r115_SUM_15_, add_1_root_r115_SUM_16_,
         add_1_root_r115_SUM_17_, add_1_root_r115_SUM_18_,
         add_1_root_r115_SUM_19_, add_1_root_r115_SUM_20_,
         add_1_root_r115_SUM_21_, add_1_root_r115_SUM_22_,
         add_1_root_r115_SUM_23_, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n24, n25, n27, n28, n29, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n158, n160, n161, n162, n163, n164, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290;
  wire   [16:0] in_17bit_b;
  wire   [23:8] neg_mul;
  wire   [16:13] sub_add_75_b0_carry;
  wire   [16:2] sub_add_54_b0_carry;
  wire   [22:7] add_1_root_r119_carry;

  multi16_8_DW01_add_0 add_0_root_r119 ( .A_22_(add_2_root_r119_SUM_22_), 
        .A_21_(add_2_root_r119_SUM_21_), .A_20_(add_2_root_r119_SUM_20_), 
        .A_19_(add_2_root_r119_SUM_19_), .A_18_(add_2_root_r119_SUM_18_), 
        .A_17_(add_2_root_r119_SUM_17_), .A_16_(add_2_root_r119_SUM_16_), 
        .A_15_(add_2_root_r119_SUM_15_), .A_14_(add_2_root_r119_SUM_14_), 
        .A_13_(add_2_root_r119_SUM_13_), .A_12_(add_2_root_r119_SUM_12_), 
        .A_11_(add_2_root_r119_SUM_11_), .A_10_(add_2_root_r119_SUM_10_), 
        .A_9_(add_2_root_r119_SUM_9_), .A_8_(add_2_root_r119_SUM_8_), .A_7_(
        add_2_root_r119_SUM_7_), .A_6_(add_2_root_r119_SUM_6_), .A_5_(
        add_1_root_r119_A_2_), .A_4_(in_17bit_b[0]), .B_23_(
        add_1_root_r119_SUM_23_), .B_22_(add_1_root_r119_SUM_22_), .B_21_(
        add_1_root_r119_SUM_21_), .B_20_(add_1_root_r119_SUM_20_), .B_19_(
        add_1_root_r119_SUM_19_), .B_18_(add_1_root_r119_SUM_18_), .B_17_(
        add_1_root_r119_SUM_17_), .B_16_(add_1_root_r119_SUM_16_), .B_15_(
        add_1_root_r119_SUM_15_), .B_14_(add_1_root_r119_SUM_14_), .B_13_(
        add_1_root_r119_SUM_13_), .B_12_(add_1_root_r119_SUM_12_), .B_11_(
        add_1_root_r119_SUM_11_), .B_10_(add_1_root_r119_SUM_10_), .B_9_(
        add_1_root_r119_SUM_9_), .B_8_(add_1_root_r119_SUM_8_), .B_7_(
        add_1_root_r119_SUM_7_), .B_6_(add_1_root_r119_SUM_6_), .B_5_(
        add_1_root_r119_A_5_), .B_4_(add_1_root_r119_A_4_), .SUM_23_(N363), 
        .SUM_22_(N362), .SUM_21_(N361), .SUM_20_(N360), .SUM_19_(N359), 
        .SUM_18_(N358), .SUM_17_(N357), .SUM_16_(N356), .SUM_15_(N355), 
        .SUM_14_(N354), .SUM_13_(N353), .SUM_12_(N352), .SUM_11_(N351), 
        .SUM_10_(N350), .SUM_9_(N349), .SUM_8_(N348), .SUM_7_(N347) );
  multi16_8_DW01_add_4 add_0_root_r112 ( .A_21_(in_17bit_b[16]), .A_20_(
        in_17bit_b[15]), .A_19_(in_17bit_b[14]), .A_18_(in_17bit_b[13]), 
        .A_17_(in_17bit_b[12]), .A_16_(in_17bit_b[11]), .A_15_(in_17bit_b[10]), 
        .A_14_(in_17bit_b[9]), .A_13_(in_17bit_b[8]), .A_12_(in_17bit_b[7]), 
        .A_11_(in_17bit_b[6]), .A_10_(in_17bit_b[5]), .A_9_(in_17bit_b[4]), 
        .A_8_(in_17bit_b[3]), .A_7_(in_17bit_b[2]), .A_6_(in_17bit_b[1]), 
        .A_5_(in_17bit_b[0]), .B_21_(add_1_root_r112_SUM_21_), .B_20_(
        add_1_root_r112_SUM_20_), .B_19_(add_1_root_r112_SUM_19_), .B_18_(
        add_1_root_r112_SUM_18_), .B_17_(add_1_root_r112_SUM_17_), .B_16_(
        add_1_root_r112_SUM_16_), .B_15_(add_1_root_r112_SUM_15_), .B_14_(
        add_1_root_r112_SUM_14_), .B_13_(add_1_root_r112_SUM_13_), .B_12_(
        add_1_root_r112_SUM_12_), .B_11_(add_1_root_r112_SUM_11_), .B_10_(
        add_1_root_r112_SUM_10_), .B_9_(add_1_root_r112_SUM_9_), .B_8_(
        add_1_root_r112_SUM_8_), .B_7_(add_1_root_r112_SUM_7_), .B_6_(
        add_1_root_r112_SUM_6_), .B_5_(add_1_root_r112_SUM_5_), .SUM_22_(N123), 
        .SUM_21_(N122), .SUM_20_(N121), .SUM_19_(N120), .SUM_18_(N119), 
        .SUM_17_(N118), .SUM_16_(N117), .SUM_15_(N116), .SUM_14_(N115), 
        .SUM_13_(N114), .SUM_12_(N113), .SUM_11_(N112), .SUM_10_(N111), 
        .SUM_9_(N110), .SUM_8_(N109), .SUM_7_(N108) );
  multi16_8_DW01_add_6 add_0_root_r115 ( .A_23_(add_1_root_r115_SUM_23_), 
        .A_22_(add_1_root_r115_SUM_22_), .A_21_(add_1_root_r115_SUM_21_), 
        .A_20_(add_1_root_r115_SUM_20_), .A_19_(add_1_root_r115_SUM_19_), 
        .A_18_(add_1_root_r115_SUM_18_), .A_17_(add_1_root_r115_SUM_17_), 
        .A_16_(add_1_root_r115_SUM_16_), .A_15_(add_1_root_r115_SUM_15_), 
        .A_14_(add_1_root_r115_SUM_14_), .A_13_(add_1_root_r115_SUM_13_), 
        .A_12_(add_1_root_r115_SUM_12_), .A_11_(add_1_root_r115_SUM_11_), 
        .A_10_(add_1_root_r115_SUM_10_), .A_9_(add_1_root_r115_SUM_9_), .A_8_(
        add_1_root_r115_SUM_8_), .A_7_(add_1_root_r115_SUM_7_), .A_6_(
        add_2_root_r115_SUM_3_), .A_5_(in_17bit_b[1]), .A_4_(in_17bit_b[0]), 
        .B_20_(add_2_root_r115_SUM_20_), .B_19_(add_2_root_r115_SUM_19_), 
        .B_18_(add_2_root_r115_SUM_18_), .B_17_(add_2_root_r115_SUM_17_), 
        .B_16_(add_2_root_r115_SUM_16_), .B_15_(add_2_root_r115_SUM_15_), 
        .B_14_(add_2_root_r115_SUM_14_), .B_13_(add_2_root_r115_SUM_13_), 
        .B_12_(add_2_root_r115_SUM_12_), .B_11_(add_2_root_r115_SUM_11_), 
        .B_10_(add_2_root_r115_SUM_10_), .B_9_(add_2_root_r115_SUM_9_), .B_8_(
        add_2_root_r115_SUM_8_), .B_7_(add_2_root_r115_SUM_7_), .B_6_(
        add_2_root_r115_SUM_6_), .B_5_(add_2_root_r115_SUM_5_), .B_4_(
        add_2_root_r115_SUM_4_), .SUM_23_(N221), .SUM_22_(N220), .SUM_21_(N219), .SUM_20_(N218), .SUM_19_(N217), .SUM_18_(N216), .SUM_17_(N215), .SUM_16_(
        N214), .SUM_15_(N213), .SUM_14_(N212), .SUM_13_(N211), .SUM_12_(N210), 
        .SUM_11_(N209), .SUM_10_(N208), .SUM_9_(N207), .SUM_8_(N206), .SUM_7_(
        N205) );
  TLATX1 neg_mul_reg_19_ ( .G(N446), .D(N459), .QN(n5) );
  TLATX1 neg_mul_reg_18_ ( .G(N446), .D(N458), .QN(n1) );
  TLATX1 neg_mul_reg_17_ ( .G(N446), .D(N457), .QN(n4) );
  TLATX1 neg_mul_reg_16_ ( .G(N446), .D(N456), .QN(n3) );
  TLATX1 neg_mul_reg_15_ ( .G(N446), .D(N455), .QN(n2) );
  TLATX1 neg_mul_reg_23_ ( .G(N446), .D(N463), .Q(neg_mul[23]), .QN(n16) );
  TLATX1 neg_mul_reg_22_ ( .G(N446), .D(N462), .Q(neg_mul[22]), .QN(n8) );
  TLATX1 neg_mul_reg_21_ ( .G(N446), .D(N461), .QN(n35) );
  TLATX1 neg_mul_reg_20_ ( .G(N446), .D(N460), .QN(n12) );
  TLATX1 neg_mul_reg_9_ ( .G(N446), .D(N449), .Q(neg_mul[9]), .QN(n15) );
  TLATX1 neg_mul_reg_14_ ( .G(N446), .D(N454), .Q(neg_mul[14]), .QN(n11) );
  TLATX1 neg_mul_reg_13_ ( .G(N446), .D(N453), .Q(neg_mul[13]), .QN(n10) );
  TLATX1 neg_mul_reg_12_ ( .G(N446), .D(N452), .Q(neg_mul[12]), .QN(n9) );
  TLATX1 neg_mul_reg_11_ ( .G(N446), .D(N451), .Q(neg_mul[11]), .QN(n7) );
  TLATX1 neg_mul_reg_10_ ( .G(N446), .D(N450), .Q(neg_mul[10]), .QN(n14) );
  TLATX1 neg_mul_reg_8_ ( .G(N446), .D(N448), .Q(neg_mul[8]), .QN(n13) );
  TLATX1 neg_mul_reg_7_ ( .G(N446), .D(N447), .Q(out[0]) );
  NAND2X1 U2 ( .A(n45), .B(n9), .Y(n86) );
  NOR2X2 U3 ( .A(n38), .B(n172), .Y(n174) );
  INVX1 U4 ( .A(n57), .Y(n55) );
  CLKINVX3 U5 ( .A(n24), .Y(n57) );
  CLKINVX3 U6 ( .A(n290), .Y(in_17bit_b[16]) );
  AOI2BB2X2 U7 ( .B0(n80), .B1(n44), .A0N(n45), .A1N(neg_mul[11]), .Y(n81) );
  CLKINVX8 U8 ( .A(n47), .Y(n44) );
  OAI21X2 U9 ( .A0(n27), .A1(n64), .B0(n63), .Y(n69) );
  INVX12 U10 ( .A(n47), .Y(n27) );
  XNOR2X4 U11 ( .A(n176), .B(n5), .Y(out[12]) );
  NOR2X2 U12 ( .A(n177), .B(n40), .Y(n176) );
  INVX8 U13 ( .A(in_8bit[7]), .Y(n47) );
  AOI2BB2X1 U14 ( .B0(n88), .B1(n31), .A0N(n44), .A1N(neg_mul[12]), .Y(n89) );
  OAI21XL U15 ( .A0(n31), .A1(n79), .B0(n78), .Y(n84) );
  NOR2X2 U16 ( .A(n28), .B(n81), .Y(n83) );
  AOI2BB2X2 U17 ( .B0(n65), .B1(n27), .A0N(n45), .A1N(neg_mul[9]), .Y(n66) );
  OAI2BB1X1 U18 ( .A0N(n47), .A1N(n6), .B0(n59), .Y(n62) );
  MXI2X1 U19 ( .A(n35), .B(n17), .S0(n178), .Y(out[14]) );
  INVX1 U20 ( .A(n18), .Y(n76) );
  XNOR2X2 U21 ( .A(n28), .B(n27), .Y(n177) );
  INVX4 U22 ( .A(n177), .Y(n178) );
  NAND4BXL U23 ( .AN(n44), .B(n53), .C(in_8bit[1]), .D(in_8bit[4]), .Y(n189)
         );
  AND2X2 U24 ( .A(out[0]), .B(neg_mul[8]), .Y(n6) );
  XNOR2X1 U25 ( .A(n35), .B(sub_add_75_b0_carry[14]), .Y(n17) );
  NAND2X2 U26 ( .A(n45), .B(n7), .Y(n78) );
  CLKINVX8 U27 ( .A(n19), .Y(out[2]) );
  OR2X2 U28 ( .A(neg_mul[9]), .B(n46), .Y(n63) );
  MX2X1 U29 ( .A(n71), .B(neg_mul[10]), .S0(in_8bit[7]), .Y(n18) );
  INVX4 U30 ( .A(n295), .Y(n19) );
  AOI211X2 U31 ( .A0(n56), .A1(n69), .B0(n68), .C0(n67), .Y(n295) );
  NOR2BX2 U32 ( .AN(n58), .B(n97), .Y(n99) );
  INVX8 U33 ( .A(n25), .Y(out[1]) );
  BUFX8 U34 ( .A(n293), .Y(out[5]) );
  AOI211X2 U35 ( .A0(n56), .A1(n92), .B0(n91), .C0(n90), .Y(n293) );
  NAND2X2 U36 ( .A(n45), .B(n13), .Y(n59) );
  BUFX8 U37 ( .A(n292), .Y(out[6]) );
  AOI211X2 U38 ( .A0(n24), .A1(n100), .B0(n99), .C0(n98), .Y(n292) );
  BUFX8 U39 ( .A(n291), .Y(out[7]) );
  AOI211X2 U40 ( .A0(n24), .A1(n164), .B0(n163), .C0(n36), .Y(n291) );
  NOR4BXL U41 ( .AN(n233), .B(n209), .C(in_8bit[1]), .D(in_8bit[2]), .Y(n234)
         );
  NOR2BX4 U42 ( .AN(n58), .B(n73), .Y(n75) );
  NOR2BX4 U43 ( .AN(n58), .B(n66), .Y(n68) );
  INVX4 U44 ( .A(n296), .Y(n25) );
  OAI21X1 U45 ( .A0(n44), .A1(n160), .B0(n158), .Y(n164) );
  NOR2BX2 U46 ( .AN(n58), .B(n162), .Y(n163) );
  CLKINVX8 U47 ( .A(n46), .Y(n45) );
  INVX8 U48 ( .A(n29), .Y(n24) );
  CLKINVX8 U49 ( .A(n28), .Y(n29) );
  AOI211X2 U50 ( .A0(n28), .A1(n62), .B0(n61), .C0(n42), .Y(n296) );
  BUFX20 U51 ( .A(in_17bit[16]), .Y(n28) );
  NOR2X4 U52 ( .A(n28), .B(n60), .Y(n61) );
  NAND3XL U53 ( .A(n44), .B(n52), .C(n50), .Y(n188) );
  NOR2BX2 U54 ( .AN(n58), .B(n89), .Y(n91) );
  OAI21X1 U55 ( .A0(n44), .A1(n95), .B0(n94), .Y(n100) );
  BUFX8 U56 ( .A(n294), .Y(out[3]) );
  AOI211X2 U57 ( .A0(n56), .A1(n76), .B0(n75), .C0(n74), .Y(n294) );
  INVX8 U58 ( .A(in_8bit[7]), .Y(n46) );
  AOI2BB2X1 U59 ( .B0(n96), .B1(n45), .A0N(n45), .A1N(neg_mul[13]), .Y(n97) );
  XNOR2X4 U60 ( .A(n28), .B(n31), .Y(n170) );
  XNOR2X2 U61 ( .A(n28), .B(n31), .Y(n175) );
  INVX8 U62 ( .A(n58), .Y(n56) );
  AOI2BB2X2 U63 ( .B0(n161), .B1(n31), .A0N(n31), .A1N(neg_mul[14]), .Y(n162)
         );
  XNOR2X4 U64 ( .A(n28), .B(n27), .Y(n172) );
  CLKINVX8 U65 ( .A(n46), .Y(n31) );
  INVX1 U66 ( .A(n240), .Y(in_17bit_b[1]) );
  INVX1 U67 ( .A(n279), .Y(in_17bit_b[14]) );
  INVX1 U68 ( .A(n276), .Y(in_17bit_b[13]) );
  INVX1 U69 ( .A(n243), .Y(in_17bit_b[2]) );
  INVX1 U70 ( .A(n252), .Y(in_17bit_b[5]) );
  INVX1 U71 ( .A(n255), .Y(in_17bit_b[6]) );
  INVX1 U72 ( .A(n258), .Y(in_17bit_b[7]) );
  INVX1 U73 ( .A(n261), .Y(in_17bit_b[8]) );
  INVX1 U74 ( .A(n264), .Y(in_17bit_b[9]) );
  INVX1 U75 ( .A(n267), .Y(in_17bit_b[10]) );
  INVX1 U76 ( .A(n270), .Y(in_17bit_b[11]) );
  INVX1 U77 ( .A(n273), .Y(in_17bit_b[12]) );
  INVX1 U78 ( .A(n249), .Y(in_17bit_b[4]) );
  INVX1 U79 ( .A(n246), .Y(in_17bit_b[3]) );
  XNOR2X4 U80 ( .A(n32), .B(n1), .Y(out[11]) );
  NOR2X4 U81 ( .A(n39), .B(n175), .Y(n32) );
  AOI21X1 U82 ( .A0(n33), .A1(n34), .B0(n283), .Y(n236) );
  NOR4XL U83 ( .A(in_8bit[4]), .B(n49), .C(n53), .D(n27), .Y(n33) );
  NOR4XL U84 ( .A(in_8bit[1]), .B(in_8bit[0]), .C(in_8bit[2]), .D(in_8bit[3]), 
        .Y(n34) );
  NAND3X1 U85 ( .A(in_8bit[2]), .B(n51), .C(n49), .Y(n231) );
  NAND3BX1 U86 ( .AN(n49), .B(n48), .C(in_8bit[3]), .Y(n232) );
  INVX1 U87 ( .A(n50), .Y(n49) );
  INVX1 U88 ( .A(n54), .Y(n53) );
  INVX1 U89 ( .A(n208), .Y(n289) );
  OAI21XL U90 ( .A0(n289), .A1(n290), .B0(n288), .Y(N463) );
  AOI22X1 U91 ( .A0(N221), .A1(n287), .B0(N363), .B1(n286), .Y(n288) );
  ADDFX2 U92 ( .A(in_17bit_b[16]), .B(in_17bit_b[12]), .CI(
        add_1_root_r112_carry_16_), .CO(add_1_root_r112_carry_17_), .S(
        add_1_root_r112_SUM_16_) );
  ADDFX2 U93 ( .A(add_1_root_r119_A_19_), .B(in_17bit_b[13]), .CI(
        add_1_root_r119_carry[19]), .CO(add_1_root_r119_carry[20]), .S(
        add_1_root_r119_SUM_19_) );
  ADDFX2 U94 ( .A(in_17bit_b[16]), .B(in_17bit_b[15]), .CI(
        add_3_root_r119_carry_17_), .CO(add_3_root_r119_carry_18_), .S(
        add_1_root_r119_A_17_) );
  ADDFX2 U95 ( .A(in_17bit_b[16]), .B(in_17bit_b[14]), .CI(
        add_2_root_r115_carry_17_), .CO(add_2_root_r115_carry_18_), .S(
        add_2_root_r115_SUM_17_) );
  ADDFX2 U96 ( .A(in_17bit_b[16]), .B(in_17bit_b[14]), .CI(
        add_1_root_r115_carry_20_), .CO(add_1_root_r115_carry_21_), .S(
        add_1_root_r115_SUM_20_) );
  ADDFX2 U97 ( .A(in_17bit_b[16]), .B(in_17bit_b[15]), .CI(
        add_2_root_r119_carry_20_), .CO(add_2_root_r119_carry_21_), .S(
        add_2_root_r119_SUM_20_) );
  ADDFX2 U98 ( .A(in_17bit_b[3]), .B(in_17bit_b[1]), .CI(
        add_2_root_r115_carry_4_), .CO(add_2_root_r115_carry_5_), .S(
        add_2_root_r115_SUM_4_) );
  ADDFX2 U99 ( .A(in_17bit_b[4]), .B(in_17bit_b[2]), .CI(
        add_2_root_r115_carry_5_), .CO(add_2_root_r115_carry_6_), .S(
        add_2_root_r115_SUM_5_) );
  ADDFX2 U100 ( .A(in_17bit_b[5]), .B(in_17bit_b[1]), .CI(
        add_1_root_r112_carry_5_), .CO(add_1_root_r112_carry_6_), .S(
        add_1_root_r112_SUM_5_) );
  ADDFX2 U101 ( .A(in_17bit_b[6]), .B(in_17bit_b[5]), .CI(
        add_3_root_r119_carry_7_), .CO(add_3_root_r119_carry_8_), .S(
        add_1_root_r119_A_7_) );
  ADDFX2 U102 ( .A(in_17bit_b[6]), .B(in_17bit_b[2]), .CI(
        add_1_root_r112_carry_6_), .CO(add_1_root_r112_carry_7_), .S(
        add_1_root_r112_SUM_6_) );
  ADDFX2 U103 ( .A(in_17bit_b[3]), .B(in_17bit_b[1]), .CI(
        add_2_root_r115_carry_4_), .CO(add_1_root_r115_carry_8_), .S(
        add_1_root_r115_SUM_7_) );
  ADDFX2 U104 ( .A(in_17bit_b[7]), .B(in_17bit_b[6]), .CI(
        add_3_root_r119_carry_8_), .CO(add_3_root_r119_carry_9_), .S(
        add_1_root_r119_A_8_) );
  ADDFX2 U105 ( .A(add_1_root_r119_A_7_), .B(in_17bit_b[1]), .CI(
        add_1_root_r119_carry[7]), .CO(add_1_root_r119_carry[8]), .S(
        add_1_root_r119_SUM_7_) );
  ADDFX2 U106 ( .A(in_17bit_b[2]), .B(in_17bit_b[1]), .CI(
        add_3_root_r119_carry_3_), .CO(add_2_root_r119_carry_7_), .S(
        add_2_root_r119_SUM_6_) );
  ADDFX2 U107 ( .A(in_17bit_b[4]), .B(in_17bit_b[2]), .CI(
        add_1_root_r115_carry_8_), .CO(add_1_root_r115_carry_9_), .S(
        add_1_root_r115_SUM_8_) );
  ADDFX2 U108 ( .A(in_17bit_b[8]), .B(in_17bit_b[7]), .CI(
        add_3_root_r119_carry_9_), .CO(add_3_root_r119_carry_10_), .S(
        add_1_root_r119_A_9_) );
  ADDFX2 U109 ( .A(add_1_root_r119_A_8_), .B(in_17bit_b[2]), .CI(
        add_1_root_r119_carry[8]), .CO(add_1_root_r119_carry[9]), .S(
        add_1_root_r119_SUM_8_) );
  ADDFX2 U110 ( .A(in_17bit_b[3]), .B(in_17bit_b[2]), .CI(
        add_2_root_r119_carry_7_), .CO(add_2_root_r119_carry_8_), .S(
        add_2_root_r119_SUM_7_) );
  ADDFX2 U111 ( .A(in_17bit_b[6]), .B(in_17bit_b[4]), .CI(
        add_2_root_r115_carry_7_), .CO(add_2_root_r115_carry_8_), .S(
        add_2_root_r115_SUM_7_) );
  ADDFX2 U112 ( .A(in_17bit_b[9]), .B(in_17bit_b[8]), .CI(
        add_3_root_r119_carry_10_), .CO(add_3_root_r119_carry_11_), .S(
        add_1_root_r119_A_10_) );
  ADDFX2 U113 ( .A(in_17bit_b[7]), .B(in_17bit_b[5]), .CI(
        add_2_root_r115_carry_8_), .CO(add_2_root_r115_carry_9_), .S(
        add_2_root_r115_SUM_8_) );
  ADDFX2 U114 ( .A(in_17bit_b[9]), .B(in_17bit_b[5]), .CI(
        add_1_root_r112_carry_9_), .CO(add_1_root_r112_carry_10_), .S(
        add_1_root_r112_SUM_9_) );
  ADDFX2 U115 ( .A(in_17bit_b[6]), .B(in_17bit_b[4]), .CI(
        add_1_root_r115_carry_10_), .CO(add_1_root_r115_carry_11_), .S(
        add_1_root_r115_SUM_10_) );
  ADDFX2 U116 ( .A(in_17bit_b[10]), .B(in_17bit_b[9]), .CI(
        add_3_root_r119_carry_11_), .CO(add_3_root_r119_carry_12_), .S(
        add_1_root_r119_A_11_) );
  ADDFX2 U117 ( .A(in_17bit_b[8]), .B(in_17bit_b[4]), .CI(
        add_1_root_r112_carry_8_), .CO(add_1_root_r112_carry_9_), .S(
        add_1_root_r112_SUM_8_) );
  ADDFX2 U118 ( .A(add_1_root_r119_A_10_), .B(in_17bit_b[4]), .CI(
        add_1_root_r119_carry[10]), .CO(add_1_root_r119_carry[11]), .S(
        add_1_root_r119_SUM_10_) );
  ADDFX2 U119 ( .A(in_17bit_b[5]), .B(in_17bit_b[4]), .CI(
        add_2_root_r119_carry_9_), .CO(add_2_root_r119_carry_10_), .S(
        add_2_root_r119_SUM_9_) );
  ADDFX2 U120 ( .A(in_17bit_b[8]), .B(in_17bit_b[6]), .CI(
        add_2_root_r115_carry_9_), .CO(add_2_root_r115_carry_10_), .S(
        add_2_root_r115_SUM_9_) );
  ADDFX2 U121 ( .A(in_17bit_b[10]), .B(in_17bit_b[6]), .CI(
        add_1_root_r112_carry_10_), .CO(add_1_root_r112_carry_11_), .S(
        add_1_root_r112_SUM_10_) );
  ADDFX2 U122 ( .A(in_17bit_b[7]), .B(in_17bit_b[5]), .CI(
        add_1_root_r115_carry_11_), .CO(add_1_root_r115_carry_12_), .S(
        add_1_root_r115_SUM_11_) );
  ADDFX2 U123 ( .A(in_17bit_b[11]), .B(in_17bit_b[10]), .CI(
        add_3_root_r119_carry_12_), .CO(add_3_root_r119_carry_13_), .S(
        add_1_root_r119_A_12_) );
  ADDFX2 U124 ( .A(add_1_root_r119_A_11_), .B(in_17bit_b[5]), .CI(
        add_1_root_r119_carry[11]), .CO(add_1_root_r119_carry[12]), .S(
        add_1_root_r119_SUM_11_) );
  ADDFX2 U125 ( .A(in_17bit_b[6]), .B(in_17bit_b[5]), .CI(
        add_2_root_r119_carry_10_), .CO(add_2_root_r119_carry_11_), .S(
        add_2_root_r119_SUM_10_) );
  ADDFX2 U126 ( .A(in_17bit_b[9]), .B(in_17bit_b[7]), .CI(
        add_2_root_r115_carry_10_), .CO(add_2_root_r115_carry_11_), .S(
        add_2_root_r115_SUM_10_) );
  ADDFX2 U127 ( .A(in_17bit_b[11]), .B(in_17bit_b[7]), .CI(
        add_1_root_r112_carry_11_), .CO(add_1_root_r112_carry_12_), .S(
        add_1_root_r112_SUM_11_) );
  ADDFX2 U128 ( .A(in_17bit_b[8]), .B(in_17bit_b[6]), .CI(
        add_1_root_r115_carry_12_), .CO(add_1_root_r115_carry_13_), .S(
        add_1_root_r115_SUM_12_) );
  ADDFX2 U129 ( .A(in_17bit_b[12]), .B(in_17bit_b[11]), .CI(
        add_3_root_r119_carry_13_), .CO(add_3_root_r119_carry_14_), .S(
        add_1_root_r119_A_13_) );
  ADDFX2 U130 ( .A(add_1_root_r119_A_12_), .B(in_17bit_b[6]), .CI(
        add_1_root_r119_carry[12]), .CO(add_1_root_r119_carry[13]), .S(
        add_1_root_r119_SUM_12_) );
  ADDFX2 U131 ( .A(in_17bit_b[7]), .B(in_17bit_b[6]), .CI(
        add_2_root_r119_carry_11_), .CO(add_2_root_r119_carry_12_), .S(
        add_2_root_r119_SUM_11_) );
  ADDFX2 U132 ( .A(in_17bit_b[10]), .B(in_17bit_b[8]), .CI(
        add_2_root_r115_carry_11_), .CO(add_2_root_r115_carry_12_), .S(
        add_2_root_r115_SUM_11_) );
  ADDFX2 U133 ( .A(in_17bit_b[12]), .B(in_17bit_b[8]), .CI(
        add_1_root_r112_carry_12_), .CO(add_1_root_r112_carry_13_), .S(
        add_1_root_r112_SUM_12_) );
  ADDFX2 U134 ( .A(in_17bit_b[9]), .B(in_17bit_b[7]), .CI(
        add_1_root_r115_carry_13_), .CO(add_1_root_r115_carry_14_), .S(
        add_1_root_r115_SUM_13_) );
  ADDFX2 U135 ( .A(in_17bit_b[13]), .B(in_17bit_b[12]), .CI(
        add_3_root_r119_carry_14_), .CO(add_3_root_r119_carry_15_), .S(
        add_1_root_r119_A_14_) );
  ADDFX2 U136 ( .A(add_1_root_r119_A_13_), .B(in_17bit_b[7]), .CI(
        add_1_root_r119_carry[13]), .CO(add_1_root_r119_carry[14]), .S(
        add_1_root_r119_SUM_13_) );
  ADDFX2 U137 ( .A(in_17bit_b[8]), .B(in_17bit_b[7]), .CI(
        add_2_root_r119_carry_12_), .CO(add_2_root_r119_carry_13_), .S(
        add_2_root_r119_SUM_12_) );
  ADDFX2 U138 ( .A(in_17bit_b[11]), .B(in_17bit_b[9]), .CI(
        add_2_root_r115_carry_12_), .CO(add_2_root_r115_carry_13_), .S(
        add_2_root_r115_SUM_12_) );
  ADDFX2 U139 ( .A(in_17bit_b[13]), .B(in_17bit_b[9]), .CI(
        add_1_root_r112_carry_13_), .CO(add_1_root_r112_carry_14_), .S(
        add_1_root_r112_SUM_13_) );
  ADDFX2 U140 ( .A(in_17bit_b[10]), .B(in_17bit_b[8]), .CI(
        add_1_root_r115_carry_14_), .CO(add_1_root_r115_carry_15_), .S(
        add_1_root_r115_SUM_14_) );
  ADDFX2 U141 ( .A(in_17bit_b[14]), .B(in_17bit_b[13]), .CI(
        add_3_root_r119_carry_15_), .CO(add_3_root_r119_carry_16_), .S(
        add_1_root_r119_A_15_) );
  ADDFX2 U142 ( .A(add_1_root_r119_A_14_), .B(in_17bit_b[8]), .CI(
        add_1_root_r119_carry[14]), .CO(add_1_root_r119_carry[15]), .S(
        add_1_root_r119_SUM_14_) );
  ADDFX2 U143 ( .A(in_17bit_b[9]), .B(in_17bit_b[8]), .CI(
        add_2_root_r119_carry_13_), .CO(add_2_root_r119_carry_14_), .S(
        add_2_root_r119_SUM_13_) );
  ADDFX2 U144 ( .A(in_17bit_b[12]), .B(in_17bit_b[10]), .CI(
        add_2_root_r115_carry_13_), .CO(add_2_root_r115_carry_14_), .S(
        add_2_root_r115_SUM_13_) );
  ADDFX2 U145 ( .A(in_17bit_b[14]), .B(in_17bit_b[10]), .CI(
        add_1_root_r112_carry_14_), .CO(add_1_root_r112_carry_15_), .S(
        add_1_root_r112_SUM_14_) );
  ADDFX2 U146 ( .A(in_17bit_b[11]), .B(in_17bit_b[9]), .CI(
        add_1_root_r115_carry_15_), .CO(add_1_root_r115_carry_16_), .S(
        add_1_root_r115_SUM_15_) );
  ADDFX2 U147 ( .A(add_1_root_r119_A_15_), .B(in_17bit_b[9]), .CI(
        add_1_root_r119_carry[15]), .CO(add_1_root_r119_carry[16]), .S(
        add_1_root_r119_SUM_15_) );
  ADDFX2 U148 ( .A(in_17bit_b[3]), .B(in_17bit_b[2]), .CI(
        add_3_root_r119_carry_4_), .CO(add_3_root_r119_carry_5_), .S(
        add_1_root_r119_A_4_) );
  ADDFX2 U149 ( .A(in_17bit_b[2]), .B(in_17bit_b[1]), .CI(
        add_3_root_r119_carry_3_), .CO(add_3_root_r119_carry_4_), .S(
        add_1_root_r119_A_3_) );
  ADDFX2 U150 ( .A(in_17bit_b[10]), .B(in_17bit_b[9]), .CI(
        add_2_root_r119_carry_14_), .CO(add_2_root_r119_carry_15_), .S(
        add_2_root_r119_SUM_14_) );
  ADDFX2 U151 ( .A(in_17bit_b[13]), .B(in_17bit_b[11]), .CI(
        add_2_root_r115_carry_14_), .CO(add_2_root_r115_carry_15_), .S(
        add_2_root_r115_SUM_14_) );
  ADDFX2 U152 ( .A(in_17bit_b[15]), .B(in_17bit_b[11]), .CI(
        add_1_root_r112_carry_15_), .CO(add_1_root_r112_carry_16_), .S(
        add_1_root_r112_SUM_15_) );
  ADDFX2 U153 ( .A(in_17bit_b[12]), .B(in_17bit_b[10]), .CI(
        add_1_root_r115_carry_16_), .CO(add_1_root_r115_carry_17_), .S(
        add_1_root_r115_SUM_16_) );
  ADDFX2 U154 ( .A(add_1_root_r119_A_16_), .B(in_17bit_b[10]), .CI(
        add_1_root_r119_carry[16]), .CO(add_1_root_r119_carry[17]), .S(
        add_1_root_r119_SUM_16_) );
  ADDFX2 U155 ( .A(in_17bit_b[11]), .B(in_17bit_b[10]), .CI(
        add_2_root_r119_carry_15_), .CO(add_2_root_r119_carry_16_), .S(
        add_2_root_r119_SUM_15_) );
  ADDFX2 U156 ( .A(in_17bit_b[14]), .B(in_17bit_b[12]), .CI(
        add_2_root_r115_carry_15_), .CO(add_2_root_r115_carry_16_), .S(
        add_2_root_r115_SUM_15_) );
  ADDFX2 U157 ( .A(in_17bit_b[13]), .B(in_17bit_b[11]), .CI(
        add_1_root_r115_carry_17_), .CO(add_1_root_r115_carry_18_), .S(
        add_1_root_r115_SUM_17_) );
  ADDFX2 U158 ( .A(add_1_root_r119_A_17_), .B(in_17bit_b[11]), .CI(
        add_1_root_r119_carry[17]), .CO(add_1_root_r119_carry[18]), .S(
        add_1_root_r119_SUM_17_) );
  ADDFX2 U159 ( .A(in_17bit_b[12]), .B(in_17bit_b[11]), .CI(
        add_2_root_r119_carry_16_), .CO(add_2_root_r119_carry_17_), .S(
        add_2_root_r119_SUM_16_) );
  ADDFX2 U160 ( .A(in_17bit_b[15]), .B(in_17bit_b[13]), .CI(
        add_2_root_r115_carry_16_), .CO(add_2_root_r115_carry_17_), .S(
        add_2_root_r115_SUM_16_) );
  ADDFX2 U161 ( .A(add_1_root_r119_A_18_), .B(in_17bit_b[12]), .CI(
        add_1_root_r119_carry[18]), .CO(add_1_root_r119_carry[19]), .S(
        add_1_root_r119_SUM_18_) );
  ADDFX2 U162 ( .A(in_17bit_b[13]), .B(in_17bit_b[12]), .CI(
        add_2_root_r119_carry_17_), .CO(add_2_root_r119_carry_18_), .S(
        add_2_root_r119_SUM_17_) );
  ADDFX2 U163 ( .A(in_17bit_b[15]), .B(in_17bit_b[13]), .CI(
        add_1_root_r115_carry_19_), .CO(add_1_root_r115_carry_20_), .S(
        add_1_root_r115_SUM_19_) );
  ADDFX2 U164 ( .A(in_17bit_b[5]), .B(in_17bit_b[3]), .CI(
        add_2_root_r115_carry_6_), .CO(add_2_root_r115_carry_7_), .S(
        add_2_root_r115_SUM_6_) );
  ADDFX2 U165 ( .A(in_17bit_b[7]), .B(in_17bit_b[3]), .CI(
        add_1_root_r112_carry_7_), .CO(add_1_root_r112_carry_8_), .S(
        add_1_root_r112_SUM_7_) );
  ADDFX2 U166 ( .A(in_17bit_b[5]), .B(in_17bit_b[3]), .CI(
        add_1_root_r115_carry_9_), .CO(add_1_root_r115_carry_10_), .S(
        add_1_root_r115_SUM_9_) );
  ADDFX2 U167 ( .A(add_1_root_r119_A_9_), .B(in_17bit_b[3]), .CI(
        add_1_root_r119_carry[9]), .CO(add_1_root_r119_carry[10]), .S(
        add_1_root_r119_SUM_9_) );
  ADDFX2 U168 ( .A(in_17bit_b[4]), .B(in_17bit_b[3]), .CI(
        add_2_root_r119_carry_8_), .CO(add_2_root_r119_carry_9_), .S(
        add_2_root_r119_SUM_8_) );
  ADDFX2 U169 ( .A(in_17bit_b[15]), .B(in_17bit_b[14]), .CI(
        add_3_root_r119_carry_16_), .CO(add_3_root_r119_carry_17_), .S(
        add_1_root_r119_A_16_) );
  ADDFX2 U170 ( .A(in_17bit_b[14]), .B(in_17bit_b[12]), .CI(
        add_1_root_r115_carry_18_), .CO(add_1_root_r115_carry_19_), .S(
        add_1_root_r115_SUM_18_) );
  ADDFX2 U171 ( .A(in_17bit_b[5]), .B(in_17bit_b[4]), .CI(
        add_3_root_r119_carry_6_), .CO(add_3_root_r119_carry_7_), .S(
        add_1_root_r119_A_6_) );
  ADDFX2 U172 ( .A(in_17bit_b[14]), .B(in_17bit_b[13]), .CI(
        add_2_root_r119_carry_18_), .CO(add_2_root_r119_carry_19_), .S(
        add_2_root_r119_SUM_18_) );
  ADDFX2 U173 ( .A(in_17bit_b[4]), .B(in_17bit_b[3]), .CI(
        add_3_root_r119_carry_5_), .CO(add_3_root_r119_carry_6_), .S(
        add_1_root_r119_A_5_) );
  ADDFX2 U174 ( .A(in_17bit_b[15]), .B(in_17bit_b[14]), .CI(
        add_2_root_r119_carry_19_), .CO(add_2_root_r119_carry_20_), .S(
        add_2_root_r119_SUM_19_) );
  INVX1 U175 ( .A(in_8bit[2]), .Y(n48) );
  INVX1 U176 ( .A(in_8bit[4]), .Y(n52) );
  INVX1 U177 ( .A(in_8bit[3]), .Y(n51) );
  INVX1 U178 ( .A(in_8bit[6]), .Y(n54) );
  INVX1 U179 ( .A(in_8bit[5]), .Y(n50) );
  NOR3X1 U180 ( .A(n48), .B(n51), .C(n209), .Y(n235) );
  CLKINVX3 U181 ( .A(n237), .Y(in_17bit_b[0]) );
  NAND2XL U182 ( .A(N29), .B(n24), .Y(n290) );
  INVX1 U183 ( .A(n85), .Y(n82) );
  CLKINVX3 U184 ( .A(n282), .Y(in_17bit_b[15]) );
  OR2X2 U185 ( .A(n184), .B(n183), .Y(n286) );
  NOR2X1 U186 ( .A(n185), .B(n231), .Y(n183) );
  NOR2X1 U187 ( .A(n232), .B(n230), .Y(n184) );
  OR2X2 U188 ( .A(n187), .B(n186), .Y(n287) );
  NOR2X1 U189 ( .A(n185), .B(n232), .Y(n186) );
  NOR2X1 U190 ( .A(n231), .B(n230), .Y(n187) );
  OAI2BB1X1 U191 ( .A0N(n234), .A1N(n191), .B0(n190), .Y(n208) );
  INVX1 U192 ( .A(n188), .Y(n191) );
  NAND3BX1 U193 ( .AN(n189), .B(n235), .C(n49), .Y(n190) );
  NAND3X1 U194 ( .A(n234), .B(n49), .C(n179), .Y(n180) );
  NOR2XL U195 ( .A(n27), .B(n52), .Y(n179) );
  INVX1 U196 ( .A(n77), .Y(n74) );
  INVX1 U197 ( .A(n93), .Y(n90) );
  INVX1 U198 ( .A(n101), .Y(n98) );
  NAND2X1 U199 ( .A(n239), .B(n238), .Y(N447) );
  AOI22X1 U200 ( .A0(N108), .A1(n283), .B0(N205), .B1(n287), .Y(n238) );
  AOI22X1 U201 ( .A0(N347), .A1(n286), .B0(n208), .B1(in_17bit_b[0]), .Y(n239)
         );
  NAND2X1 U202 ( .A(n242), .B(n241), .Y(N448) );
  AOI22X1 U203 ( .A0(N109), .A1(n283), .B0(N206), .B1(n287), .Y(n241) );
  AOI22X1 U204 ( .A0(N348), .A1(n286), .B0(n208), .B1(in_17bit_b[1]), .Y(n242)
         );
  NAND2X1 U205 ( .A(n245), .B(n244), .Y(N449) );
  AOI22X1 U206 ( .A0(N110), .A1(n283), .B0(N207), .B1(n287), .Y(n244) );
  AOI22X1 U207 ( .A0(N349), .A1(n286), .B0(n208), .B1(in_17bit_b[2]), .Y(n245)
         );
  NAND2X1 U208 ( .A(n248), .B(n247), .Y(N450) );
  AOI22X1 U209 ( .A0(N111), .A1(n283), .B0(N208), .B1(n287), .Y(n247) );
  AOI22X1 U210 ( .A0(N350), .A1(n286), .B0(n208), .B1(in_17bit_b[3]), .Y(n248)
         );
  NAND2X1 U211 ( .A(n251), .B(n250), .Y(N451) );
  AOI22X1 U212 ( .A0(N112), .A1(n283), .B0(N209), .B1(n287), .Y(n250) );
  AOI22X1 U213 ( .A0(N351), .A1(n286), .B0(n208), .B1(in_17bit_b[4]), .Y(n251)
         );
  NAND2X1 U214 ( .A(n254), .B(n253), .Y(N452) );
  AOI22X1 U215 ( .A0(N113), .A1(n283), .B0(N210), .B1(n287), .Y(n253) );
  AOI22X1 U216 ( .A0(N352), .A1(n286), .B0(n208), .B1(in_17bit_b[5]), .Y(n254)
         );
  NAND2X1 U217 ( .A(n257), .B(n256), .Y(N453) );
  AOI22X1 U218 ( .A0(N114), .A1(n283), .B0(N211), .B1(n287), .Y(n256) );
  AOI22X1 U219 ( .A0(N353), .A1(n286), .B0(n208), .B1(in_17bit_b[6]), .Y(n257)
         );
  NAND2X1 U220 ( .A(n260), .B(n259), .Y(N454) );
  AOI22X1 U221 ( .A0(N115), .A1(n283), .B0(N212), .B1(n287), .Y(n259) );
  AOI22X1 U222 ( .A0(N354), .A1(n286), .B0(n208), .B1(in_17bit_b[7]), .Y(n260)
         );
  NAND2X1 U223 ( .A(n263), .B(n262), .Y(N455) );
  AOI22X1 U224 ( .A0(N116), .A1(n283), .B0(N213), .B1(n287), .Y(n262) );
  AOI22X1 U225 ( .A0(N355), .A1(n286), .B0(n208), .B1(in_17bit_b[8]), .Y(n263)
         );
  NAND2X1 U226 ( .A(n266), .B(n265), .Y(N456) );
  AOI22X1 U227 ( .A0(N117), .A1(n283), .B0(N214), .B1(n287), .Y(n265) );
  AOI22X1 U228 ( .A0(N356), .A1(n286), .B0(n208), .B1(in_17bit_b[9]), .Y(n266)
         );
  NAND2X1 U229 ( .A(n269), .B(n268), .Y(N457) );
  AOI22X1 U230 ( .A0(N118), .A1(n283), .B0(N215), .B1(n287), .Y(n268) );
  AOI22X1 U231 ( .A0(N357), .A1(n286), .B0(n208), .B1(in_17bit_b[10]), .Y(n269) );
  NAND2X1 U232 ( .A(n272), .B(n271), .Y(N458) );
  AOI22X1 U233 ( .A0(N119), .A1(n283), .B0(N216), .B1(n287), .Y(n271) );
  AOI22X1 U234 ( .A0(N358), .A1(n286), .B0(n208), .B1(in_17bit_b[11]), .Y(n272) );
  NAND2X1 U235 ( .A(n275), .B(n274), .Y(N459) );
  AOI22X1 U236 ( .A0(N120), .A1(n283), .B0(N217), .B1(n287), .Y(n274) );
  AOI22X1 U237 ( .A0(N359), .A1(n286), .B0(n208), .B1(in_17bit_b[12]), .Y(n275) );
  NAND2X1 U238 ( .A(n278), .B(n277), .Y(N460) );
  AOI22X1 U239 ( .A0(N121), .A1(n283), .B0(N218), .B1(n287), .Y(n277) );
  AOI22X1 U240 ( .A0(N360), .A1(n286), .B0(n208), .B1(in_17bit_b[13]), .Y(n278) );
  NAND2X1 U241 ( .A(n281), .B(n280), .Y(N461) );
  AOI22X1 U242 ( .A0(N122), .A1(n283), .B0(N219), .B1(n287), .Y(n280) );
  AOI22X1 U243 ( .A0(N361), .A1(n286), .B0(n208), .B1(in_17bit_b[14]), .Y(n281) );
  NAND2X1 U244 ( .A(n285), .B(n284), .Y(N462) );
  AOI22X1 U245 ( .A0(N123), .A1(n283), .B0(N220), .B1(n287), .Y(n284) );
  AOI22X1 U246 ( .A0(N362), .A1(n286), .B0(n208), .B1(in_17bit_b[15]), .Y(n285) );
  OAI21X1 U247 ( .A0(n44), .A1(n87), .B0(n86), .Y(n92) );
  NAND2XL U248 ( .A(n45), .B(n10), .Y(n94) );
  NAND2XL U249 ( .A(n45), .B(n11), .Y(n158) );
  INVX1 U250 ( .A(n70), .Y(n67) );
  NAND4BBX1 U251 ( .AN(n286), .BN(n287), .C(n236), .D(n289), .Y(N446) );
  NAND4XL U252 ( .A(in_8bit[1]), .B(n44), .C(n229), .D(n209), .Y(n230) );
  NOR2X1 U253 ( .A(n53), .B(in_8bit[4]), .Y(n229) );
  NOR2X1 U254 ( .A(n53), .B(in_8bit[3]), .Y(n233) );
  AOI22XL U255 ( .A0(in_17bit[0]), .A1(n55), .B0(in_17bit[0]), .B1(n57), .Y(
        n237) );
  AOI22X1 U256 ( .A0(N27), .A1(n55), .B0(in_17bit[14]), .B1(n57), .Y(n279) );
  AOI22X1 U257 ( .A0(N28), .A1(n55), .B0(in_17bit[15]), .B1(n57), .Y(n282) );
  AOI22X1 U258 ( .A0(N16), .A1(n55), .B0(in_17bit[3]), .B1(n57), .Y(n246) );
  AOI22X1 U259 ( .A0(N17), .A1(n55), .B0(in_17bit[4]), .B1(n57), .Y(n249) );
  AOI22X1 U260 ( .A0(N18), .A1(n55), .B0(in_17bit[5]), .B1(n57), .Y(n252) );
  AOI22X1 U261 ( .A0(N19), .A1(n55), .B0(in_17bit[6]), .B1(n57), .Y(n255) );
  AOI22X1 U262 ( .A0(N20), .A1(n55), .B0(in_17bit[7]), .B1(n57), .Y(n258) );
  AOI22X1 U263 ( .A0(N21), .A1(n55), .B0(in_17bit[8]), .B1(n57), .Y(n261) );
  AOI22X1 U264 ( .A0(N22), .A1(n55), .B0(in_17bit[9]), .B1(n57), .Y(n264) );
  AOI22X1 U265 ( .A0(N23), .A1(n55), .B0(in_17bit[10]), .B1(n57), .Y(n267) );
  AOI22X1 U266 ( .A0(N24), .A1(n55), .B0(in_17bit[11]), .B1(n57), .Y(n270) );
  AOI22X1 U267 ( .A0(N25), .A1(n55), .B0(in_17bit[12]), .B1(n57), .Y(n273) );
  AOI22X1 U268 ( .A0(N26), .A1(n55), .B0(in_17bit[13]), .B1(n57), .Y(n276) );
  AOI22XL U269 ( .A0(N14), .A1(n24), .B0(in_17bit[1]), .B1(n57), .Y(n240) );
  AOI22XL U270 ( .A0(N15), .A1(n55), .B0(in_17bit[2]), .B1(n57), .Y(n243) );
  INVXL U271 ( .A(in_8bit[0]), .Y(n209) );
  AND2X2 U272 ( .A(n98), .B(n11), .Y(n36) );
  NAND2X1 U273 ( .A(n42), .B(n15), .Y(n70) );
  AND2X2 U274 ( .A(n36), .B(n2), .Y(n37) );
  AND2X2 U275 ( .A(n37), .B(n3), .Y(n38) );
  AND2X2 U276 ( .A(n38), .B(n4), .Y(n39) );
  OR2XL U277 ( .A(n189), .B(in_8bit[0]), .Y(n185) );
  OAI2BB1X1 U278 ( .A0N(n182), .A1N(n181), .B0(n180), .Y(n283) );
  NOR2BX1 U279 ( .AN(n235), .B(n54), .Y(n182) );
  NOR2BX1 U280 ( .AN(in_8bit[1]), .B(n188), .Y(n181) );
  NAND2BX1 U281 ( .AN(n70), .B(n14), .Y(n77) );
  NAND2X1 U282 ( .A(n74), .B(n7), .Y(n85) );
  NAND2X1 U283 ( .A(n82), .B(n9), .Y(n93) );
  NAND2X1 U284 ( .A(n90), .B(n10), .Y(n101) );
  AND2X2 U285 ( .A(n39), .B(n1), .Y(n40) );
  INVX1 U286 ( .A(in_17bit[3]), .Y(n195) );
  INVX1 U287 ( .A(in_17bit[4]), .Y(n196) );
  INVX1 U288 ( .A(in_17bit[5]), .Y(n197) );
  INVX1 U289 ( .A(in_17bit[6]), .Y(n198) );
  INVX1 U290 ( .A(in_17bit[7]), .Y(n199) );
  INVX1 U291 ( .A(in_17bit[8]), .Y(n200) );
  INVX1 U292 ( .A(in_17bit[9]), .Y(n201) );
  INVX1 U293 ( .A(in_17bit[10]), .Y(n202) );
  INVX1 U294 ( .A(in_17bit[11]), .Y(n203) );
  INVX1 U295 ( .A(in_17bit[12]), .Y(n204) );
  INVX1 U296 ( .A(in_17bit[13]), .Y(n205) );
  INVX1 U297 ( .A(in_17bit[14]), .Y(n206) );
  INVX1 U298 ( .A(in_17bit[15]), .Y(n207) );
  INVX1 U299 ( .A(in_17bit[1]), .Y(n193) );
  INVX1 U300 ( .A(in_17bit[2]), .Y(n194) );
  INVX1 U301 ( .A(in_17bit[0]), .Y(n192) );
  XNOR2X1 U302 ( .A(n12), .B(sub_add_75_b0_carry[13]), .Y(n41) );
  INVX1 U303 ( .A(n79), .Y(n80) );
  INVX1 U304 ( .A(n87), .Y(n88) );
  INVX1 U305 ( .A(n71), .Y(n72) );
  INVX1 U306 ( .A(n160), .Y(n161) );
  INVX1 U307 ( .A(n95), .Y(n96) );
  INVX1 U308 ( .A(n64), .Y(n65) );
  MX2X1 U309 ( .A(neg_mul[22]), .B(N480), .S0(n178), .Y(out[15]) );
  MX2X1 U310 ( .A(neg_mul[23]), .B(N481), .S0(n178), .Y(out[16]) );
  NOR2X1 U311 ( .A(out[0]), .B(neg_mul[8]), .Y(n42) );
  NAND2BX1 U312 ( .AN(n42), .B(neg_mul[9]), .Y(n64) );
  NAND2X1 U313 ( .A(neg_mul[10]), .B(n70), .Y(n71) );
  NAND2X1 U314 ( .A(neg_mul[11]), .B(n77), .Y(n79) );
  NAND2X1 U315 ( .A(neg_mul[13]), .B(n93), .Y(n95) );
  NAND2X1 U316 ( .A(neg_mul[14]), .B(n101), .Y(n160) );
  NAND2X1 U317 ( .A(neg_mul[12]), .B(n85), .Y(n87) );
  INVX8 U318 ( .A(in_17bit[16]), .Y(n58) );
  AOI2BB2X4 U319 ( .B0(n6), .B1(n27), .A0N(n44), .A1N(neg_mul[8]), .Y(n60) );
  AOI2BB2X4 U320 ( .B0(n72), .B1(n31), .A0N(n31), .A1N(neg_mul[10]), .Y(n73)
         );
  AOI211X2 U321 ( .A0(n56), .A1(n84), .B0(n83), .C0(n82), .Y(out[4]) );
  NOR2X4 U322 ( .A(n36), .B(n170), .Y(n171) );
  XNOR2X4 U323 ( .A(n171), .B(n2), .Y(out[8]) );
  NOR2X4 U324 ( .A(n37), .B(n172), .Y(n173) );
  XNOR2X4 U325 ( .A(n173), .B(n3), .Y(out[9]) );
  XNOR2X4 U326 ( .A(n174), .B(n4), .Y(out[10]) );
  MXI2X4 U327 ( .A(n12), .B(n41), .S0(n178), .Y(out[13]) );
  AND2X1 U328 ( .A(add_1_root_r112_carry_20_), .B(in_17bit_b[16]), .Y(
        add_1_root_r112_SUM_21_) );
  XOR2X1 U329 ( .A(in_17bit_b[16]), .B(add_1_root_r112_carry_20_), .Y(
        add_1_root_r112_SUM_20_) );
  AND2X1 U330 ( .A(add_1_root_r112_carry_19_), .B(in_17bit_b[15]), .Y(
        add_1_root_r112_carry_20_) );
  XOR2X1 U331 ( .A(in_17bit_b[15]), .B(add_1_root_r112_carry_19_), .Y(
        add_1_root_r112_SUM_19_) );
  AND2X1 U332 ( .A(add_1_root_r112_carry_18_), .B(in_17bit_b[14]), .Y(
        add_1_root_r112_carry_19_) );
  XOR2X1 U333 ( .A(in_17bit_b[14]), .B(add_1_root_r112_carry_18_), .Y(
        add_1_root_r112_SUM_18_) );
  AND2X1 U334 ( .A(add_1_root_r112_carry_17_), .B(in_17bit_b[13]), .Y(
        add_1_root_r112_carry_18_) );
  XOR2X1 U335 ( .A(in_17bit_b[13]), .B(add_1_root_r112_carry_17_), .Y(
        add_1_root_r112_SUM_17_) );
  AND2X1 U336 ( .A(add_2_root_r119_carry_21_), .B(in_17bit_b[16]), .Y(
        add_2_root_r119_SUM_22_) );
  XOR2X1 U337 ( .A(in_17bit_b[16]), .B(add_2_root_r119_carry_21_), .Y(
        add_2_root_r119_SUM_21_) );
  AND2X1 U338 ( .A(add_1_root_r119_carry[22]), .B(in_17bit_b[16]), .Y(
        add_1_root_r119_SUM_23_) );
  XOR2X1 U339 ( .A(in_17bit_b[16]), .B(add_1_root_r119_carry[22]), .Y(
        add_1_root_r119_SUM_22_) );
  AND2X1 U340 ( .A(add_1_root_r119_carry[21]), .B(in_17bit_b[15]), .Y(
        add_1_root_r119_carry[22]) );
  XOR2X1 U341 ( .A(in_17bit_b[15]), .B(add_1_root_r119_carry[21]), .Y(
        add_1_root_r119_SUM_21_) );
  AND2X1 U342 ( .A(add_1_root_r119_carry[20]), .B(in_17bit_b[14]), .Y(
        add_1_root_r119_carry[21]) );
  XOR2X1 U343 ( .A(in_17bit_b[14]), .B(add_1_root_r119_carry[20]), .Y(
        add_1_root_r119_SUM_20_) );
  AND2X1 U344 ( .A(add_1_root_r119_A_6_), .B(in_17bit_b[0]), .Y(
        add_1_root_r119_carry[7]) );
  XOR2X1 U345 ( .A(in_17bit_b[0]), .B(add_1_root_r119_A_6_), .Y(
        add_1_root_r119_SUM_6_) );
  AND2X1 U346 ( .A(add_3_root_r119_carry_18_), .B(in_17bit_b[16]), .Y(
        add_1_root_r119_A_19_) );
  XOR2X1 U347 ( .A(in_17bit_b[16]), .B(add_3_root_r119_carry_18_), .Y(
        add_1_root_r119_A_18_) );
  AND2X1 U348 ( .A(in_17bit_b[1]), .B(in_17bit_b[0]), .Y(
        add_3_root_r119_carry_3_) );
  XOR2X1 U349 ( .A(in_17bit_b[0]), .B(in_17bit_b[1]), .Y(add_1_root_r119_A_2_)
         );
  AND2X1 U350 ( .A(add_2_root_r115_carry_19_), .B(in_17bit_b[16]), .Y(
        add_2_root_r115_SUM_20_) );
  XOR2X1 U351 ( .A(in_17bit_b[16]), .B(add_2_root_r115_carry_19_), .Y(
        add_2_root_r115_SUM_19_) );
  AND2X1 U352 ( .A(add_2_root_r115_carry_18_), .B(in_17bit_b[15]), .Y(
        add_2_root_r115_carry_19_) );
  XOR2X1 U353 ( .A(in_17bit_b[15]), .B(add_2_root_r115_carry_18_), .Y(
        add_2_root_r115_SUM_18_) );
  AND2X1 U354 ( .A(in_17bit_b[2]), .B(in_17bit_b[0]), .Y(
        add_2_root_r115_carry_4_) );
  XOR2X1 U355 ( .A(in_17bit_b[0]), .B(in_17bit_b[2]), .Y(
        add_2_root_r115_SUM_3_) );
  AND2X1 U356 ( .A(add_1_root_r115_carry_22_), .B(in_17bit_b[16]), .Y(
        add_1_root_r115_SUM_23_) );
  XOR2X1 U357 ( .A(in_17bit_b[16]), .B(add_1_root_r115_carry_22_), .Y(
        add_1_root_r115_SUM_22_) );
  AND2X1 U358 ( .A(add_1_root_r115_carry_21_), .B(in_17bit_b[15]), .Y(
        add_1_root_r115_carry_22_) );
  XOR2X1 U359 ( .A(in_17bit_b[15]), .B(add_1_root_r115_carry_21_), .Y(
        add_1_root_r115_SUM_21_) );
  XOR2X1 U360 ( .A(n57), .B(sub_add_54_b0_carry[16]), .Y(N29) );
  AND2X1 U361 ( .A(sub_add_54_b0_carry[15]), .B(n207), .Y(
        sub_add_54_b0_carry[16]) );
  XOR2X1 U362 ( .A(n207), .B(sub_add_54_b0_carry[15]), .Y(N28) );
  AND2X1 U363 ( .A(sub_add_54_b0_carry[14]), .B(n206), .Y(
        sub_add_54_b0_carry[15]) );
  XOR2X1 U364 ( .A(n206), .B(sub_add_54_b0_carry[14]), .Y(N27) );
  AND2X1 U365 ( .A(sub_add_54_b0_carry[13]), .B(n205), .Y(
        sub_add_54_b0_carry[14]) );
  XOR2X1 U366 ( .A(n205), .B(sub_add_54_b0_carry[13]), .Y(N26) );
  AND2X1 U367 ( .A(sub_add_54_b0_carry[12]), .B(n204), .Y(
        sub_add_54_b0_carry[13]) );
  XOR2X1 U368 ( .A(n204), .B(sub_add_54_b0_carry[12]), .Y(N25) );
  AND2X1 U369 ( .A(sub_add_54_b0_carry[11]), .B(n203), .Y(
        sub_add_54_b0_carry[12]) );
  XOR2X1 U370 ( .A(n203), .B(sub_add_54_b0_carry[11]), .Y(N24) );
  AND2X1 U371 ( .A(sub_add_54_b0_carry[10]), .B(n202), .Y(
        sub_add_54_b0_carry[11]) );
  XOR2X1 U372 ( .A(n202), .B(sub_add_54_b0_carry[10]), .Y(N23) );
  AND2X1 U373 ( .A(sub_add_54_b0_carry[9]), .B(n201), .Y(
        sub_add_54_b0_carry[10]) );
  XOR2X1 U374 ( .A(n201), .B(sub_add_54_b0_carry[9]), .Y(N22) );
  AND2X1 U375 ( .A(sub_add_54_b0_carry[8]), .B(n200), .Y(
        sub_add_54_b0_carry[9]) );
  XOR2X1 U376 ( .A(n200), .B(sub_add_54_b0_carry[8]), .Y(N21) );
  AND2X1 U377 ( .A(sub_add_54_b0_carry[7]), .B(n199), .Y(
        sub_add_54_b0_carry[8]) );
  XOR2X1 U378 ( .A(n199), .B(sub_add_54_b0_carry[7]), .Y(N20) );
  AND2X1 U379 ( .A(sub_add_54_b0_carry[6]), .B(n198), .Y(
        sub_add_54_b0_carry[7]) );
  XOR2X1 U380 ( .A(n198), .B(sub_add_54_b0_carry[6]), .Y(N19) );
  AND2X1 U381 ( .A(sub_add_54_b0_carry[5]), .B(n197), .Y(
        sub_add_54_b0_carry[6]) );
  XOR2X1 U382 ( .A(n197), .B(sub_add_54_b0_carry[5]), .Y(N18) );
  AND2X1 U383 ( .A(sub_add_54_b0_carry[4]), .B(n196), .Y(
        sub_add_54_b0_carry[5]) );
  XOR2X1 U384 ( .A(n196), .B(sub_add_54_b0_carry[4]), .Y(N17) );
  AND2X1 U385 ( .A(sub_add_54_b0_carry[3]), .B(n195), .Y(
        sub_add_54_b0_carry[4]) );
  XOR2X1 U386 ( .A(n195), .B(sub_add_54_b0_carry[3]), .Y(N16) );
  AND2X1 U387 ( .A(sub_add_54_b0_carry[2]), .B(n194), .Y(
        sub_add_54_b0_carry[3]) );
  XOR2X1 U388 ( .A(n194), .B(sub_add_54_b0_carry[2]), .Y(N15) );
  AND2X1 U389 ( .A(n192), .B(n193), .Y(sub_add_54_b0_carry[2]) );
  XOR2X1 U390 ( .A(n193), .B(n192), .Y(N14) );
  XOR2X1 U391 ( .A(n16), .B(sub_add_75_b0_carry[16]), .Y(N481) );
  AND2X1 U392 ( .A(sub_add_75_b0_carry[15]), .B(n8), .Y(
        sub_add_75_b0_carry[16]) );
  XOR2X1 U393 ( .A(n8), .B(sub_add_75_b0_carry[15]), .Y(N480) );
  AND2X1 U394 ( .A(sub_add_75_b0_carry[14]), .B(n35), .Y(
        sub_add_75_b0_carry[15]) );
  AND2X1 U395 ( .A(sub_add_75_b0_carry[13]), .B(n12), .Y(
        sub_add_75_b0_carry[14]) );
  AND2X1 U396 ( .A(n40), .B(n5), .Y(sub_add_75_b0_carry[13]) );
  AND2X1 U397 ( .A(in_17bit_b[0]), .B(in_17bit_b[4]), .Y(
        add_1_root_r112_carry_5_) );
endmodule


module multi16_7_DW01_add_0 ( A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, 
        A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, 
        A_4_, B_23_, B_22_, B_21_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, 
        B_14_, B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, 
        SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, 
        SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, 
        SUM_7_ );
  input A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_,
         A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, B_23_, B_22_,
         B_21_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_,
         B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_;
  output SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_,
         SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_,
         SUM_8_, SUM_7_;
  wire   n1, n2, n3, n4;
  wire   [23:7] carry;

  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry[7]), .CO(carry[8]), .S(SUM_7_)
         );
  ADDFX2 U1_21 ( .A(A_21_), .B(B_21_), .CI(carry[21]), .CO(carry[22]), .S(
        SUM_21_) );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry[20]), .CO(carry[21]), .S(
        SUM_20_) );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry[19]), .CO(carry[20]), .S(
        SUM_19_) );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry[18]), .CO(carry[19]), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry[17]), .CO(carry[18]), .S(
        SUM_17_) );
  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry[16]), .CO(carry[17]), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry[15]), .CO(carry[16]), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry[14]), .CO(carry[15]), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry[13]), .CO(carry[14]), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry[12]), .CO(carry[13]), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry[11]), .CO(carry[12]), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry[10]), .CO(carry[11]), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry[9]), .CO(carry[10]), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry[8]), .CO(carry[9]), .S(SUM_8_)
         );
  ADDFX2 U1_22 ( .A(A_22_), .B(B_22_), .CI(carry[22]), .CO(carry[23]), .S(
        SUM_22_) );
  AND2X2 U1 ( .A(A_4_), .B(B_4_), .Y(n1) );
  XOR2X1 U2 ( .A(B_23_), .B(carry[23]), .Y(SUM_23_) );
  OAI2BB1X1 U3 ( .A0N(n2), .A1N(A_6_), .B0(n3), .Y(carry[7]) );
  OAI21XL U4 ( .A0(A_6_), .A1(n2), .B0(B_6_), .Y(n3) );
  OAI2BB1X1 U5 ( .A0N(n1), .A1N(A_5_), .B0(n4), .Y(n2) );
  OAI21XL U6 ( .A0(A_5_), .A1(n1), .B0(B_5_), .Y(n4) );
endmodule


module multi16_7_DW01_add_4 ( A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, 
        A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, 
        B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, 
        B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, SUM_22_, SUM_21_, SUM_20_, 
        SUM_19_, SUM_18_, SUM_17_, SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, 
        SUM_11_, SUM_10_, SUM_9_, SUM_8_, SUM_7_ );
  input A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_,
         A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, B_20_, B_19_,
         B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, B_10_, B_9_,
         B_8_, B_7_, B_6_, B_5_;
  output SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_,
         SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_,
         SUM_7_;
  wire   carry_21_, carry_20_, carry_19_, carry_18_, carry_17_, carry_16_,
         carry_15_, carry_14_, carry_13_, carry_12_, carry_11_, carry_10_,
         carry_9_, carry_8_, carry_7_, n1;

  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry_16_), .CO(carry_17_), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry_15_), .CO(carry_16_), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry_14_), .CO(carry_15_), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry_13_), .CO(carry_14_), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry_12_), .CO(carry_13_), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry_11_), .CO(carry_12_), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry_10_), .CO(carry_11_), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry_9_), .CO(carry_10_), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry_8_), .CO(carry_9_), .S(SUM_8_)
         );
  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry_7_), .CO(carry_8_), .S(SUM_7_)
         );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry_20_), .CO(carry_21_), .S(
        SUM_20_) );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry_19_), .CO(carry_20_), .S(
        SUM_19_) );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry_18_), .CO(carry_19_), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry_17_), .CO(carry_18_), .S(
        SUM_17_) );
  ADDFX2 U1_21 ( .A(A_21_), .B(B_21_), .CI(carry_21_), .CO(SUM_22_), .S(
        SUM_21_) );
  OAI2BB1X1 U1 ( .A0N(A_6_), .A1N(B_6_), .B0(n1), .Y(carry_7_) );
  OAI211X1 U2 ( .A0(B_6_), .A1(A_6_), .B0(A_5_), .C0(B_5_), .Y(n1) );
endmodule


module multi16_7_DW01_add_6 ( A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, 
        A_16_, A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, 
        A_6_, A_5_, A_4_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, 
        B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, 
        SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, 
        SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, 
        SUM_7_ );
  input A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_,
         A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, B_20_,
         B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, B_10_,
         B_9_, B_8_, B_7_, B_6_, B_5_, B_4_;
  output SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_,
         SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_,
         SUM_8_, SUM_7_;
  wire   n1, n2, n3, n4, n5, n6;
  wire   [21:7] carry;

  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry[7]), .CO(carry[8]), .S(SUM_7_)
         );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry[18]), .CO(carry[19]), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry[17]), .CO(carry[18]), .S(
        SUM_17_) );
  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry[16]), .CO(carry[17]), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry[15]), .CO(carry[16]), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry[14]), .CO(carry[15]), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry[13]), .CO(carry[14]), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry[12]), .CO(carry[13]), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry[11]), .CO(carry[12]), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry[10]), .CO(carry[11]), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry[9]), .CO(carry[10]), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry[8]), .CO(carry[9]), .S(SUM_8_)
         );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry[19]), .CO(carry[20]), .S(
        SUM_19_) );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry[20]), .CO(carry[21]), .S(
        SUM_20_) );
  AND2X2 U1 ( .A(A_22_), .B(n2), .Y(n1) );
  AND2X2 U2 ( .A(A_21_), .B(carry[21]), .Y(n2) );
  AND2X2 U3 ( .A(A_4_), .B(B_4_), .Y(n3) );
  XOR2X1 U4 ( .A(A_23_), .B(n1), .Y(SUM_23_) );
  XOR2X1 U5 ( .A(A_21_), .B(carry[21]), .Y(SUM_21_) );
  XOR2X1 U6 ( .A(A_22_), .B(n2), .Y(SUM_22_) );
  OAI2BB1X1 U7 ( .A0N(n4), .A1N(A_6_), .B0(n5), .Y(carry[7]) );
  OAI21XL U8 ( .A0(A_6_), .A1(n4), .B0(B_6_), .Y(n5) );
  OAI2BB1X1 U9 ( .A0N(n3), .A1N(A_5_), .B0(n6), .Y(n4) );
  OAI21XL U10 ( .A0(A_5_), .A1(n3), .B0(B_5_), .Y(n6) );
endmodule


module multi16_7 ( in_17bit, in_8bit, out );
  input [16:0] in_17bit;
  input [7:0] in_8bit;
  output [16:0] out;
  wire   n258, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26,
         N27, N28, N29, N108, N109, N110, N111, N112, N113, N114, N115, N116,
         N117, N118, N119, N120, N121, N122, N123, N205, N206, N207, N208,
         N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, N219,
         N220, N221, N347, N348, N349, N350, N351, N352, N353, N354, N355,
         N356, N357, N358, N359, N360, N361, N362, N363, N446, N447, N448,
         N449, N450, N451, N452, N453, N454, N455, N456, N457, N458, N459,
         N460, N461, N462, N463, N480, add_2_root_r119_carry_10_,
         add_2_root_r119_carry_11_, add_2_root_r119_carry_12_,
         add_2_root_r119_carry_13_, add_2_root_r119_carry_14_,
         add_2_root_r119_carry_15_, add_2_root_r119_carry_16_,
         add_2_root_r119_carry_17_, add_2_root_r119_carry_18_,
         add_2_root_r119_carry_19_, add_2_root_r119_carry_20_,
         add_2_root_r119_carry_21_, add_2_root_r119_carry_6_,
         add_2_root_r119_carry_7_, add_2_root_r119_carry_8_,
         add_2_root_r119_carry_9_, add_2_root_r119_SUM_5_,
         add_2_root_r119_SUM_6_, add_2_root_r119_SUM_7_,
         add_2_root_r119_SUM_8_, add_2_root_r119_SUM_9_,
         add_2_root_r119_SUM_10_, add_2_root_r119_SUM_11_,
         add_2_root_r119_SUM_12_, add_2_root_r119_SUM_13_,
         add_2_root_r119_SUM_14_, add_2_root_r119_SUM_15_,
         add_2_root_r119_SUM_16_, add_2_root_r119_SUM_17_,
         add_2_root_r119_SUM_18_, add_2_root_r119_SUM_19_,
         add_2_root_r119_SUM_20_, add_2_root_r119_SUM_21_,
         add_2_root_r119_SUM_22_, add_1_root_r119_SUM_6_,
         add_1_root_r119_SUM_7_, add_1_root_r119_SUM_8_,
         add_1_root_r119_SUM_9_, add_1_root_r119_SUM_10_,
         add_1_root_r119_SUM_11_, add_1_root_r119_SUM_12_,
         add_1_root_r119_SUM_13_, add_1_root_r119_SUM_14_,
         add_1_root_r119_SUM_15_, add_1_root_r119_SUM_16_,
         add_1_root_r119_SUM_17_, add_1_root_r119_SUM_18_,
         add_1_root_r119_SUM_19_, add_1_root_r119_SUM_20_,
         add_1_root_r119_SUM_21_, add_1_root_r119_SUM_22_,
         add_1_root_r119_SUM_23_, add_1_root_r119_A_3_, add_1_root_r119_A_4_,
         add_1_root_r119_A_5_, add_1_root_r119_A_6_, add_1_root_r119_A_7_,
         add_1_root_r119_A_8_, add_1_root_r119_A_9_, add_1_root_r119_A_10_,
         add_1_root_r119_A_11_, add_1_root_r119_A_12_, add_1_root_r119_A_13_,
         add_1_root_r119_A_14_, add_1_root_r119_A_15_, add_1_root_r119_A_16_,
         add_1_root_r119_A_17_, add_1_root_r119_A_18_, add_1_root_r119_A_19_,
         add_3_root_r119_carry_10_, add_3_root_r119_carry_11_,
         add_3_root_r119_carry_12_, add_3_root_r119_carry_13_,
         add_3_root_r119_carry_14_, add_3_root_r119_carry_15_,
         add_3_root_r119_carry_16_, add_3_root_r119_carry_17_,
         add_3_root_r119_carry_18_, add_3_root_r119_carry_4_,
         add_3_root_r119_carry_5_, add_3_root_r119_carry_6_,
         add_3_root_r119_carry_7_, add_3_root_r119_carry_8_,
         add_3_root_r119_carry_9_, add_1_root_r112_carry_10_,
         add_1_root_r112_carry_11_, add_1_root_r112_carry_12_,
         add_1_root_r112_carry_13_, add_1_root_r112_carry_14_,
         add_1_root_r112_carry_15_, add_1_root_r112_carry_16_,
         add_1_root_r112_carry_17_, add_1_root_r112_carry_18_,
         add_1_root_r112_carry_19_, add_1_root_r112_carry_20_,
         add_1_root_r112_carry_5_, add_1_root_r112_carry_6_,
         add_1_root_r112_carry_7_, add_1_root_r112_carry_8_,
         add_1_root_r112_carry_9_, add_1_root_r112_SUM_1_,
         add_1_root_r112_SUM_2_, add_1_root_r112_SUM_3_,
         add_1_root_r112_SUM_4_, add_1_root_r112_SUM_5_,
         add_1_root_r112_SUM_6_, add_1_root_r112_SUM_7_,
         add_1_root_r112_SUM_8_, add_1_root_r112_SUM_9_,
         add_1_root_r112_SUM_10_, add_1_root_r112_SUM_11_,
         add_1_root_r112_SUM_12_, add_1_root_r112_SUM_13_,
         add_1_root_r112_SUM_14_, add_1_root_r112_SUM_15_,
         add_1_root_r112_SUM_16_, add_1_root_r112_SUM_17_,
         add_1_root_r112_SUM_18_, add_1_root_r112_SUM_19_,
         add_1_root_r112_SUM_20_, add_1_root_r112_SUM_21_,
         add_2_root_r115_carry_10_, add_2_root_r115_carry_11_,
         add_2_root_r115_carry_12_, add_2_root_r115_carry_13_,
         add_2_root_r115_carry_14_, add_2_root_r115_carry_15_,
         add_2_root_r115_carry_16_, add_2_root_r115_carry_17_,
         add_2_root_r115_carry_18_, add_2_root_r115_carry_19_,
         add_2_root_r115_carry_4_, add_2_root_r115_carry_5_,
         add_2_root_r115_carry_6_, add_2_root_r115_carry_7_,
         add_2_root_r115_carry_8_, add_2_root_r115_carry_9_,
         add_2_root_r115_SUM_4_, add_2_root_r115_SUM_5_,
         add_2_root_r115_SUM_6_, add_2_root_r115_SUM_7_,
         add_2_root_r115_SUM_8_, add_2_root_r115_SUM_9_,
         add_2_root_r115_SUM_10_, add_2_root_r115_SUM_11_,
         add_2_root_r115_SUM_12_, add_2_root_r115_SUM_13_,
         add_2_root_r115_SUM_14_, add_2_root_r115_SUM_15_,
         add_2_root_r115_SUM_16_, add_2_root_r115_SUM_17_,
         add_2_root_r115_SUM_18_, add_2_root_r115_SUM_19_,
         add_2_root_r115_SUM_20_, add_1_root_r115_carry_10_,
         add_1_root_r115_carry_11_, add_1_root_r115_carry_12_,
         add_1_root_r115_carry_13_, add_1_root_r115_carry_14_,
         add_1_root_r115_carry_15_, add_1_root_r115_carry_16_,
         add_1_root_r115_carry_17_, add_1_root_r115_carry_18_,
         add_1_root_r115_carry_19_, add_1_root_r115_carry_20_,
         add_1_root_r115_carry_21_, add_1_root_r115_carry_22_,
         add_1_root_r115_carry_8_, add_1_root_r115_carry_9_,
         add_1_root_r115_SUM_6_, add_1_root_r115_SUM_7_,
         add_1_root_r115_SUM_8_, add_1_root_r115_SUM_9_,
         add_1_root_r115_SUM_10_, add_1_root_r115_SUM_11_,
         add_1_root_r115_SUM_12_, add_1_root_r115_SUM_13_,
         add_1_root_r115_SUM_14_, add_1_root_r115_SUM_15_,
         add_1_root_r115_SUM_16_, add_1_root_r115_SUM_17_,
         add_1_root_r115_SUM_18_, add_1_root_r115_SUM_19_,
         add_1_root_r115_SUM_20_, add_1_root_r115_SUM_21_,
         add_1_root_r115_SUM_22_, add_1_root_r115_SUM_23_, n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n24, n26, n27, n28, n29, n30, n31, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n158, n160, n161, n162, n163, n164,
         n167, n168, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257;
  wire   [16:0] in_17bit_b;
  wire   [23:8] neg_mul;
  wire   [15:13] sub_add_75_b0_carry;
  wire   [15:2] sub_add_54_b0_carry;
  wire   [22:7] add_1_root_r119_carry;

  multi16_7_DW01_add_0 add_0_root_r119 ( .A_22_(add_2_root_r119_SUM_22_), 
        .A_21_(add_2_root_r119_SUM_21_), .A_20_(add_2_root_r119_SUM_20_), 
        .A_19_(add_2_root_r119_SUM_19_), .A_18_(add_2_root_r119_SUM_18_), 
        .A_17_(add_2_root_r119_SUM_17_), .A_16_(add_2_root_r119_SUM_16_), 
        .A_15_(add_2_root_r119_SUM_15_), .A_14_(add_2_root_r119_SUM_14_), 
        .A_13_(add_2_root_r119_SUM_13_), .A_12_(add_2_root_r119_SUM_12_), 
        .A_11_(add_2_root_r119_SUM_11_), .A_10_(add_2_root_r119_SUM_10_), 
        .A_9_(add_2_root_r119_SUM_9_), .A_8_(add_2_root_r119_SUM_8_), .A_7_(
        add_2_root_r119_SUM_7_), .A_6_(add_2_root_r119_SUM_6_), .A_5_(
        add_2_root_r119_SUM_5_), .A_4_(in_17bit_b[0]), .B_23_(
        add_1_root_r119_SUM_23_), .B_22_(add_1_root_r119_SUM_22_), .B_21_(
        add_1_root_r119_SUM_21_), .B_20_(add_1_root_r119_SUM_20_), .B_19_(
        add_1_root_r119_SUM_19_), .B_18_(add_1_root_r119_SUM_18_), .B_17_(
        add_1_root_r119_SUM_17_), .B_16_(add_1_root_r119_SUM_16_), .B_15_(
        add_1_root_r119_SUM_15_), .B_14_(add_1_root_r119_SUM_14_), .B_13_(
        add_1_root_r119_SUM_13_), .B_12_(add_1_root_r119_SUM_12_), .B_11_(
        add_1_root_r119_SUM_11_), .B_10_(add_1_root_r119_SUM_10_), .B_9_(
        add_1_root_r119_SUM_9_), .B_8_(add_1_root_r119_SUM_8_), .B_7_(
        add_1_root_r119_SUM_7_), .B_6_(add_1_root_r119_SUM_6_), .B_5_(
        add_1_root_r119_A_5_), .B_4_(add_1_root_r119_A_4_), .SUM_23_(N363), 
        .SUM_22_(N362), .SUM_21_(N361), .SUM_20_(N360), .SUM_19_(N359), 
        .SUM_18_(N358), .SUM_17_(N357), .SUM_16_(N356), .SUM_15_(N355), 
        .SUM_14_(N354), .SUM_13_(N353), .SUM_12_(N352), .SUM_11_(N351), 
        .SUM_10_(N350), .SUM_9_(N349), .SUM_8_(N348), .SUM_7_(N347) );
  multi16_7_DW01_add_4 add_0_root_r112 ( .A_21_(in_17bit_b[16]), .A_20_(
        in_17bit_b[15]), .A_19_(in_17bit_b[14]), .A_18_(in_17bit_b[13]), 
        .A_17_(in_17bit_b[12]), .A_16_(in_17bit_b[11]), .A_15_(in_17bit_b[10]), 
        .A_14_(in_17bit_b[9]), .A_13_(in_17bit_b[8]), .A_12_(in_17bit_b[7]), 
        .A_11_(in_17bit_b[6]), .A_10_(in_17bit_b[5]), .A_9_(in_17bit_b[4]), 
        .A_8_(in_17bit_b[3]), .A_7_(in_17bit_b[2]), .A_6_(n176), .A_5_(
        in_17bit_b[0]), .B_21_(add_1_root_r112_SUM_21_), .B_20_(
        add_1_root_r112_SUM_20_), .B_19_(add_1_root_r112_SUM_19_), .B_18_(
        add_1_root_r112_SUM_18_), .B_17_(add_1_root_r112_SUM_17_), .B_16_(
        add_1_root_r112_SUM_16_), .B_15_(add_1_root_r112_SUM_15_), .B_14_(
        add_1_root_r112_SUM_14_), .B_13_(add_1_root_r112_SUM_13_), .B_12_(
        add_1_root_r112_SUM_12_), .B_11_(add_1_root_r112_SUM_11_), .B_10_(
        add_1_root_r112_SUM_10_), .B_9_(add_1_root_r112_SUM_9_), .B_8_(
        add_1_root_r112_SUM_8_), .B_7_(add_1_root_r112_SUM_7_), .B_6_(
        add_1_root_r112_SUM_6_), .B_5_(add_1_root_r112_SUM_5_), .SUM_22_(N123), 
        .SUM_21_(N122), .SUM_20_(N121), .SUM_19_(N120), .SUM_18_(N119), 
        .SUM_17_(N118), .SUM_16_(N117), .SUM_15_(N116), .SUM_14_(N115), 
        .SUM_13_(N114), .SUM_12_(N113), .SUM_11_(N112), .SUM_10_(N111), 
        .SUM_9_(N110), .SUM_8_(N109), .SUM_7_(N108) );
  multi16_7_DW01_add_6 add_0_root_r115 ( .A_23_(add_1_root_r115_SUM_23_), 
        .A_22_(add_1_root_r115_SUM_22_), .A_21_(add_1_root_r115_SUM_21_), 
        .A_20_(add_1_root_r115_SUM_20_), .A_19_(add_1_root_r115_SUM_19_), 
        .A_18_(add_1_root_r115_SUM_18_), .A_17_(add_1_root_r115_SUM_17_), 
        .A_16_(add_1_root_r115_SUM_16_), .A_15_(add_1_root_r115_SUM_15_), 
        .A_14_(add_1_root_r115_SUM_14_), .A_13_(add_1_root_r115_SUM_13_), 
        .A_12_(add_1_root_r115_SUM_12_), .A_11_(add_1_root_r115_SUM_11_), 
        .A_10_(add_1_root_r115_SUM_10_), .A_9_(add_1_root_r115_SUM_9_), .A_8_(
        add_1_root_r115_SUM_8_), .A_7_(add_1_root_r115_SUM_7_), .A_6_(
        add_1_root_r115_SUM_6_), .A_5_(n176), .A_4_(in_17bit_b[0]), .B_20_(
        add_2_root_r115_SUM_20_), .B_19_(add_2_root_r115_SUM_19_), .B_18_(
        add_2_root_r115_SUM_18_), .B_17_(add_2_root_r115_SUM_17_), .B_16_(
        add_2_root_r115_SUM_16_), .B_15_(add_2_root_r115_SUM_15_), .B_14_(
        add_2_root_r115_SUM_14_), .B_13_(add_2_root_r115_SUM_13_), .B_12_(
        add_2_root_r115_SUM_12_), .B_11_(add_2_root_r115_SUM_11_), .B_10_(
        add_2_root_r115_SUM_10_), .B_9_(add_2_root_r115_SUM_9_), .B_8_(
        add_2_root_r115_SUM_8_), .B_7_(add_2_root_r115_SUM_7_), .B_6_(
        add_2_root_r115_SUM_6_), .B_5_(add_2_root_r115_SUM_5_), .B_4_(
        add_2_root_r115_SUM_4_), .SUM_23_(N221), .SUM_22_(N220), .SUM_21_(N219), .SUM_20_(N218), .SUM_19_(N217), .SUM_18_(N216), .SUM_17_(N215), .SUM_16_(
        N214), .SUM_15_(N213), .SUM_14_(N212), .SUM_13_(N211), .SUM_12_(N210), 
        .SUM_11_(N209), .SUM_10_(N208), .SUM_9_(N207), .SUM_8_(N206), .SUM_7_(
        N205) );
  TLATX1 neg_mul_reg_19_ ( .G(N446), .D(N459), .Q(n3), .QN(n12) );
  TLATX1 neg_mul_reg_18_ ( .G(N446), .D(N458), .QN(n9) );
  TLATX1 neg_mul_reg_17_ ( .G(N446), .D(N457), .QN(n6) );
  TLATX1 neg_mul_reg_16_ ( .G(N446), .D(N456), .QN(n8) );
  TLATX1 neg_mul_reg_15_ ( .G(N446), .D(N455), .QN(n7) );
  TLATX1 neg_mul_reg_14_ ( .G(N446), .D(N454), .Q(n2), .QN(n11) );
  TLATX1 neg_mul_reg_13_ ( .G(N446), .D(N453), .Q(neg_mul[13]), .QN(n17) );
  TLATX1 neg_mul_reg_12_ ( .G(N446), .D(N452), .Q(neg_mul[12]), .QN(n16) );
  TLATX1 neg_mul_reg_11_ ( .G(N446), .D(N451), .Q(neg_mul[11]), .QN(n18) );
  TLATX1 neg_mul_reg_10_ ( .G(N446), .D(N450), .Q(neg_mul[10]), .QN(n15) );
  TLATX1 neg_mul_reg_23_ ( .G(N446), .D(N463), .Q(neg_mul[23]), .QN(n4) );
  TLATX1 neg_mul_reg_22_ ( .G(N446), .D(N462), .Q(neg_mul[22]), .QN(n10) );
  TLATX1 neg_mul_reg_21_ ( .G(N446), .D(N461), .QN(n36) );
  TLATX1 neg_mul_reg_20_ ( .G(N446), .D(N460), .QN(n13) );
  TLATX1 neg_mul_reg_9_ ( .G(N446), .D(N449), .Q(neg_mul[9]) );
  TLATX1 neg_mul_reg_8_ ( .G(N446), .D(N448), .Q(neg_mul[8]), .QN(n14) );
  TLATX1 neg_mul_reg_7_ ( .G(N446), .D(N447), .Q(out[0]) );
  CLKINVX3 U2 ( .A(n257), .Y(in_17bit_b[16]) );
  INVX12 U3 ( .A(n90), .Y(n91) );
  AOI2BB2X2 U4 ( .B0(n65), .B1(n14), .A0N(n65), .A1N(n77), .Y(n78) );
  BUFX16 U5 ( .A(n258), .Y(out[6]) );
  INVX2 U6 ( .A(n65), .Y(n29) );
  OR2X2 U7 ( .A(n90), .B(n56), .Y(n41) );
  MXI2X1 U8 ( .A(n36), .B(n20), .S0(n91), .Y(out[14]) );
  MX2X1 U9 ( .A(neg_mul[22]), .B(N480), .S0(n91), .Y(out[15]) );
  XNOR2X2 U10 ( .A(n70), .B(n29), .Y(n83) );
  INVX1 U11 ( .A(n60), .Y(n30) );
  OR2X2 U12 ( .A(n71), .B(n76), .Y(n5) );
  XNOR2X2 U13 ( .A(n71), .B(n65), .Y(n90) );
  XNOR2X4 U14 ( .A(n84), .B(neg_mul[12]), .Y(n1) );
  AOI22X1 U15 ( .A0(N27), .A1(n21), .B0(in_17bit[14]), .B1(n73), .Y(n246) );
  XNOR2X1 U16 ( .A(neg_mul[23]), .B(n61), .Y(n19) );
  INVX1 U17 ( .A(n59), .Y(n28) );
  XNOR2X1 U18 ( .A(n36), .B(sub_add_75_b0_carry[14]), .Y(n20) );
  INVX8 U19 ( .A(n69), .Y(n71) );
  CLKINVX1 U20 ( .A(in_17bit[16]), .Y(n70) );
  INVX1 U21 ( .A(n73), .Y(n21) );
  NAND3X4 U22 ( .A(n24), .B(n28), .C(n5), .Y(n22) );
  INVX8 U23 ( .A(n22), .Y(out[1]) );
  CLKINVX4 U24 ( .A(n68), .Y(n74) );
  NAND2BX4 U25 ( .AN(n82), .B(neg_mul[11]), .Y(n27) );
  NOR2X2 U26 ( .A(n52), .B(n88), .Y(n33) );
  XNOR2X4 U27 ( .A(n71), .B(n65), .Y(n80) );
  INVX8 U28 ( .A(in_17bit[16]), .Y(n69) );
  XNOR2X4 U29 ( .A(n68), .B(n65), .Y(n86) );
  NAND2X2 U30 ( .A(n82), .B(n18), .Y(n26) );
  CLKINVX8 U31 ( .A(n69), .Y(n68) );
  OR2X4 U32 ( .A(n74), .B(n78), .Y(n24) );
  INVX8 U33 ( .A(n1), .Y(out[5]) );
  NOR2X4 U34 ( .A(n80), .B(n59), .Y(n79) );
  NAND2X4 U35 ( .A(n26), .B(n27), .Y(out[4]) );
  BUFX16 U36 ( .A(in_8bit[7]), .Y(n65) );
  XOR2X4 U37 ( .A(n81), .B(neg_mul[10]), .Y(out[3]) );
  XNOR2X4 U38 ( .A(n69), .B(n65), .Y(n31) );
  NOR2BX4 U39 ( .AN(n30), .B(n86), .Y(n81) );
  INVX8 U40 ( .A(n31), .Y(n88) );
  NOR2X4 U41 ( .A(n43), .B(n83), .Y(n84) );
  XOR2X4 U42 ( .A(n85), .B(neg_mul[13]), .Y(n258) );
  NOR2X2 U43 ( .A(n88), .B(n54), .Y(n34) );
  XNOR2X4 U44 ( .A(n33), .B(n7), .Y(out[8]) );
  XNOR2X4 U45 ( .A(n34), .B(n6), .Y(out[10]) );
  NOR2X4 U46 ( .A(n86), .B(n45), .Y(n35) );
  AOI2BB2X2 U47 ( .B0(n75), .B1(n65), .A0N(n65), .A1N(neg_mul[8]), .Y(n76) );
  NOR2X4 U48 ( .A(n88), .B(n42), .Y(n82) );
  AOI22XL U49 ( .A0(N355), .A1(n253), .B0(n177), .B1(in_17bit_b[8]), .Y(n230)
         );
  AOI22XL U50 ( .A0(N356), .A1(n253), .B0(n177), .B1(in_17bit_b[9]), .Y(n233)
         );
  AOI22XL U51 ( .A0(N357), .A1(n253), .B0(n177), .B1(in_17bit_b[10]), .Y(n236)
         );
  AOI22XL U52 ( .A0(N358), .A1(n253), .B0(n177), .B1(in_17bit_b[11]), .Y(n239)
         );
  AOI22XL U53 ( .A0(N120), .A1(n250), .B0(N217), .B1(n254), .Y(n241) );
  AOI22XL U54 ( .A0(N359), .A1(n253), .B0(n177), .B1(in_17bit_b[12]), .Y(n242)
         );
  AOI22XL U55 ( .A0(N121), .A1(n250), .B0(N218), .B1(n254), .Y(n244) );
  AOI22XL U56 ( .A0(N360), .A1(n253), .B0(n177), .B1(in_17bit_b[13]), .Y(n245)
         );
  AOI22XL U57 ( .A0(N122), .A1(n250), .B0(N219), .B1(n254), .Y(n247) );
  AOI22XL U58 ( .A0(N361), .A1(n253), .B0(n177), .B1(in_17bit_b[14]), .Y(n248)
         );
  AOI22XL U59 ( .A0(N123), .A1(n250), .B0(N220), .B1(n254), .Y(n251) );
  AOI22XL U60 ( .A0(N362), .A1(n253), .B0(n177), .B1(in_17bit_b[15]), .Y(n252)
         );
  INVXL U61 ( .A(n68), .Y(n73) );
  INVX1 U62 ( .A(n246), .Y(in_17bit_b[14]) );
  INVX1 U63 ( .A(n243), .Y(in_17bit_b[13]) );
  INVX1 U64 ( .A(n210), .Y(in_17bit_b[2]) );
  INVX1 U65 ( .A(n219), .Y(in_17bit_b[5]) );
  INVX1 U66 ( .A(n222), .Y(in_17bit_b[6]) );
  INVX1 U67 ( .A(n225), .Y(in_17bit_b[7]) );
  INVX1 U68 ( .A(n228), .Y(in_17bit_b[8]) );
  INVX1 U69 ( .A(n231), .Y(in_17bit_b[9]) );
  INVX1 U70 ( .A(n234), .Y(in_17bit_b[10]) );
  INVX1 U71 ( .A(n237), .Y(in_17bit_b[11]) );
  INVX1 U72 ( .A(n240), .Y(in_17bit_b[12]) );
  INVX1 U73 ( .A(n216), .Y(in_17bit_b[4]) );
  INVX1 U74 ( .A(n213), .Y(in_17bit_b[3]) );
  XOR2X4 U75 ( .A(n35), .B(n2), .Y(out[7]) );
  AOI21X1 U76 ( .A0(n37), .A1(n38), .B0(n250), .Y(n203) );
  NOR4XL U77 ( .A(in_8bit[4]), .B(in_8bit[5]), .C(in_8bit[6]), .D(n65), .Y(n37) );
  NOR4X1 U78 ( .A(in_8bit[1]), .B(in_8bit[0]), .C(in_8bit[2]), .D(in_8bit[3]), 
        .Y(n38) );
  AND4X1 U79 ( .A(in_8bit[1]), .B(n65), .C(n198), .D(n64), .Y(n39) );
  ADDFX2 U80 ( .A(in_17bit_b[16]), .B(in_17bit_b[12]), .CI(
        add_1_root_r112_carry_16_), .CO(add_1_root_r112_carry_17_), .S(
        add_1_root_r112_SUM_16_) );
  ADDFX2 U81 ( .A(add_1_root_r119_A_19_), .B(in_17bit_b[13]), .CI(
        add_1_root_r119_carry[19]), .CO(add_1_root_r119_carry[20]), .S(
        add_1_root_r119_SUM_19_) );
  ADDFX2 U82 ( .A(in_17bit_b[16]), .B(in_17bit_b[15]), .CI(
        add_3_root_r119_carry_17_), .CO(add_3_root_r119_carry_18_), .S(
        add_1_root_r119_A_17_) );
  ADDFX2 U83 ( .A(in_17bit_b[16]), .B(in_17bit_b[14]), .CI(
        add_2_root_r115_carry_17_), .CO(add_2_root_r115_carry_18_), .S(
        add_2_root_r115_SUM_17_) );
  ADDFX2 U84 ( .A(in_17bit_b[16]), .B(in_17bit_b[14]), .CI(
        add_1_root_r115_carry_20_), .CO(add_1_root_r115_carry_21_), .S(
        add_1_root_r115_SUM_20_) );
  ADDFX2 U85 ( .A(in_17bit_b[16]), .B(in_17bit_b[15]), .CI(
        add_2_root_r119_carry_20_), .CO(add_2_root_r119_carry_21_), .S(
        add_2_root_r119_SUM_20_) );
  ADDFX2 U86 ( .A(in_17bit_b[3]), .B(n176), .CI(add_2_root_r115_carry_4_), 
        .CO(add_2_root_r115_carry_5_), .S(add_2_root_r115_SUM_4_) );
  ADDFX2 U87 ( .A(in_17bit_b[4]), .B(in_17bit_b[2]), .CI(
        add_2_root_r115_carry_5_), .CO(add_2_root_r115_carry_6_), .S(
        add_2_root_r115_SUM_5_) );
  ADDFX2 U88 ( .A(in_17bit_b[5]), .B(n176), .CI(add_1_root_r112_carry_5_), 
        .CO(add_1_root_r112_carry_6_), .S(add_1_root_r112_SUM_5_) );
  ADDFX2 U89 ( .A(in_17bit_b[6]), .B(in_17bit_b[5]), .CI(
        add_3_root_r119_carry_7_), .CO(add_3_root_r119_carry_8_), .S(
        add_1_root_r119_A_7_) );
  ADDFX2 U90 ( .A(in_17bit_b[6]), .B(in_17bit_b[2]), .CI(
        add_1_root_r112_carry_6_), .CO(add_1_root_r112_carry_7_), .S(
        add_1_root_r112_SUM_6_) );
  ADDFX2 U91 ( .A(in_17bit_b[3]), .B(n176), .CI(add_2_root_r115_carry_4_), 
        .CO(add_1_root_r115_carry_8_), .S(add_1_root_r115_SUM_7_) );
  ADDFX2 U92 ( .A(in_17bit_b[7]), .B(in_17bit_b[6]), .CI(
        add_3_root_r119_carry_8_), .CO(add_3_root_r119_carry_9_), .S(
        add_1_root_r119_A_8_) );
  ADDFX2 U93 ( .A(add_1_root_r119_A_7_), .B(n176), .CI(
        add_1_root_r119_carry[7]), .CO(add_1_root_r119_carry[8]), .S(
        add_1_root_r119_SUM_7_) );
  ADDFX2 U94 ( .A(in_17bit_b[2]), .B(n176), .CI(add_2_root_r119_carry_6_), 
        .CO(add_2_root_r119_carry_7_), .S(add_2_root_r119_SUM_6_) );
  ADDFX2 U95 ( .A(in_17bit_b[4]), .B(in_17bit_b[2]), .CI(
        add_1_root_r115_carry_8_), .CO(add_1_root_r115_carry_9_), .S(
        add_1_root_r115_SUM_8_) );
  ADDFX2 U96 ( .A(in_17bit_b[8]), .B(in_17bit_b[7]), .CI(
        add_3_root_r119_carry_9_), .CO(add_3_root_r119_carry_10_), .S(
        add_1_root_r119_A_9_) );
  ADDFX2 U97 ( .A(add_1_root_r119_A_8_), .B(in_17bit_b[2]), .CI(
        add_1_root_r119_carry[8]), .CO(add_1_root_r119_carry[9]), .S(
        add_1_root_r119_SUM_8_) );
  ADDFX2 U98 ( .A(in_17bit_b[6]), .B(in_17bit_b[4]), .CI(
        add_2_root_r115_carry_7_), .CO(add_2_root_r115_carry_8_), .S(
        add_2_root_r115_SUM_7_) );
  ADDFX2 U99 ( .A(in_17bit_b[8]), .B(in_17bit_b[4]), .CI(
        add_1_root_r112_carry_8_), .CO(add_1_root_r112_carry_9_), .S(
        add_1_root_r112_SUM_8_) );
  ADDFX2 U100 ( .A(in_17bit_b[9]), .B(in_17bit_b[8]), .CI(
        add_3_root_r119_carry_10_), .CO(add_3_root_r119_carry_11_), .S(
        add_1_root_r119_A_10_) );
  ADDFX2 U101 ( .A(in_17bit_b[7]), .B(in_17bit_b[5]), .CI(
        add_2_root_r115_carry_8_), .CO(add_2_root_r115_carry_9_), .S(
        add_2_root_r115_SUM_8_) );
  ADDFX2 U102 ( .A(in_17bit_b[10]), .B(in_17bit_b[9]), .CI(
        add_3_root_r119_carry_11_), .CO(add_3_root_r119_carry_12_), .S(
        add_1_root_r119_A_11_) );
  ADDFX2 U103 ( .A(in_17bit_b[3]), .B(in_17bit_b[2]), .CI(
        add_2_root_r119_carry_7_), .CO(add_2_root_r119_carry_8_), .S(
        add_2_root_r119_SUM_7_) );
  ADDFX2 U104 ( .A(in_17bit_b[9]), .B(in_17bit_b[5]), .CI(
        add_1_root_r112_carry_9_), .CO(add_1_root_r112_carry_10_), .S(
        add_1_root_r112_SUM_9_) );
  ADDFX2 U105 ( .A(add_1_root_r119_A_10_), .B(in_17bit_b[4]), .CI(
        add_1_root_r119_carry[10]), .CO(add_1_root_r119_carry[11]), .S(
        add_1_root_r119_SUM_10_) );
  ADDFX2 U106 ( .A(in_17bit_b[5]), .B(in_17bit_b[4]), .CI(
        add_2_root_r119_carry_9_), .CO(add_2_root_r119_carry_10_), .S(
        add_2_root_r119_SUM_9_) );
  ADDFX2 U107 ( .A(in_17bit_b[8]), .B(in_17bit_b[6]), .CI(
        add_2_root_r115_carry_9_), .CO(add_2_root_r115_carry_10_), .S(
        add_2_root_r115_SUM_9_) );
  ADDFX2 U108 ( .A(in_17bit_b[10]), .B(in_17bit_b[6]), .CI(
        add_1_root_r112_carry_10_), .CO(add_1_root_r112_carry_11_), .S(
        add_1_root_r112_SUM_10_) );
  ADDFX2 U109 ( .A(in_17bit_b[7]), .B(in_17bit_b[5]), .CI(
        add_1_root_r115_carry_11_), .CO(add_1_root_r115_carry_12_), .S(
        add_1_root_r115_SUM_11_) );
  ADDFX2 U110 ( .A(in_17bit_b[11]), .B(in_17bit_b[10]), .CI(
        add_3_root_r119_carry_12_), .CO(add_3_root_r119_carry_13_), .S(
        add_1_root_r119_A_12_) );
  ADDFX2 U111 ( .A(add_1_root_r119_A_11_), .B(in_17bit_b[5]), .CI(
        add_1_root_r119_carry[11]), .CO(add_1_root_r119_carry[12]), .S(
        add_1_root_r119_SUM_11_) );
  ADDFX2 U112 ( .A(in_17bit_b[6]), .B(in_17bit_b[5]), .CI(
        add_2_root_r119_carry_10_), .CO(add_2_root_r119_carry_11_), .S(
        add_2_root_r119_SUM_10_) );
  ADDFX2 U113 ( .A(in_17bit_b[9]), .B(in_17bit_b[7]), .CI(
        add_2_root_r115_carry_10_), .CO(add_2_root_r115_carry_11_), .S(
        add_2_root_r115_SUM_10_) );
  ADDFX2 U114 ( .A(in_17bit_b[11]), .B(in_17bit_b[7]), .CI(
        add_1_root_r112_carry_11_), .CO(add_1_root_r112_carry_12_), .S(
        add_1_root_r112_SUM_11_) );
  ADDFX2 U115 ( .A(in_17bit_b[8]), .B(in_17bit_b[6]), .CI(
        add_1_root_r115_carry_12_), .CO(add_1_root_r115_carry_13_), .S(
        add_1_root_r115_SUM_12_) );
  ADDFX2 U116 ( .A(in_17bit_b[12]), .B(in_17bit_b[11]), .CI(
        add_3_root_r119_carry_13_), .CO(add_3_root_r119_carry_14_), .S(
        add_1_root_r119_A_13_) );
  ADDFX2 U117 ( .A(add_1_root_r119_A_12_), .B(in_17bit_b[6]), .CI(
        add_1_root_r119_carry[12]), .CO(add_1_root_r119_carry[13]), .S(
        add_1_root_r119_SUM_12_) );
  ADDFX2 U118 ( .A(in_17bit_b[10]), .B(in_17bit_b[8]), .CI(
        add_2_root_r115_carry_11_), .CO(add_2_root_r115_carry_12_), .S(
        add_2_root_r115_SUM_11_) );
  ADDFX2 U119 ( .A(in_17bit_b[12]), .B(in_17bit_b[8]), .CI(
        add_1_root_r112_carry_12_), .CO(add_1_root_r112_carry_13_), .S(
        add_1_root_r112_SUM_12_) );
  ADDFX2 U120 ( .A(in_17bit_b[9]), .B(in_17bit_b[7]), .CI(
        add_1_root_r115_carry_13_), .CO(add_1_root_r115_carry_14_), .S(
        add_1_root_r115_SUM_13_) );
  ADDFX2 U121 ( .A(in_17bit_b[13]), .B(in_17bit_b[12]), .CI(
        add_3_root_r119_carry_14_), .CO(add_3_root_r119_carry_15_), .S(
        add_1_root_r119_A_14_) );
  ADDFX2 U122 ( .A(add_1_root_r119_A_13_), .B(in_17bit_b[7]), .CI(
        add_1_root_r119_carry[13]), .CO(add_1_root_r119_carry[14]), .S(
        add_1_root_r119_SUM_13_) );
  ADDFX2 U123 ( .A(in_17bit_b[8]), .B(in_17bit_b[7]), .CI(
        add_2_root_r119_carry_12_), .CO(add_2_root_r119_carry_13_), .S(
        add_2_root_r119_SUM_12_) );
  ADDFX2 U124 ( .A(in_17bit_b[13]), .B(in_17bit_b[9]), .CI(
        add_1_root_r112_carry_13_), .CO(add_1_root_r112_carry_14_), .S(
        add_1_root_r112_SUM_13_) );
  ADDFX2 U125 ( .A(in_17bit_b[10]), .B(in_17bit_b[8]), .CI(
        add_1_root_r115_carry_14_), .CO(add_1_root_r115_carry_15_), .S(
        add_1_root_r115_SUM_14_) );
  ADDFX2 U126 ( .A(in_17bit_b[14]), .B(in_17bit_b[13]), .CI(
        add_3_root_r119_carry_15_), .CO(add_3_root_r119_carry_16_), .S(
        add_1_root_r119_A_15_) );
  ADDFX2 U127 ( .A(add_1_root_r119_A_14_), .B(in_17bit_b[8]), .CI(
        add_1_root_r119_carry[14]), .CO(add_1_root_r119_carry[15]), .S(
        add_1_root_r119_SUM_14_) );
  ADDFX2 U128 ( .A(in_17bit_b[3]), .B(in_17bit_b[2]), .CI(
        add_3_root_r119_carry_4_), .CO(add_3_root_r119_carry_5_), .S(
        add_1_root_r119_A_4_) );
  ADDFX2 U129 ( .A(in_17bit_b[2]), .B(n176), .CI(add_2_root_r119_carry_6_), 
        .CO(add_3_root_r119_carry_4_), .S(add_1_root_r119_A_3_) );
  ADDFX2 U130 ( .A(in_17bit_b[9]), .B(in_17bit_b[8]), .CI(
        add_2_root_r119_carry_13_), .CO(add_2_root_r119_carry_14_), .S(
        add_2_root_r119_SUM_13_) );
  ADDFX2 U131 ( .A(in_17bit_b[12]), .B(in_17bit_b[10]), .CI(
        add_2_root_r115_carry_13_), .CO(add_2_root_r115_carry_14_), .S(
        add_2_root_r115_SUM_13_) );
  ADDFX2 U132 ( .A(in_17bit_b[14]), .B(in_17bit_b[10]), .CI(
        add_1_root_r112_carry_14_), .CO(add_1_root_r112_carry_15_), .S(
        add_1_root_r112_SUM_14_) );
  ADDFX2 U133 ( .A(in_17bit_b[11]), .B(in_17bit_b[9]), .CI(
        add_1_root_r115_carry_15_), .CO(add_1_root_r115_carry_16_), .S(
        add_1_root_r115_SUM_15_) );
  ADDFX2 U134 ( .A(add_1_root_r119_A_15_), .B(in_17bit_b[9]), .CI(
        add_1_root_r119_carry[15]), .CO(add_1_root_r119_carry[16]), .S(
        add_1_root_r119_SUM_15_) );
  ADDFX2 U135 ( .A(in_17bit_b[10]), .B(in_17bit_b[9]), .CI(
        add_2_root_r119_carry_14_), .CO(add_2_root_r119_carry_15_), .S(
        add_2_root_r119_SUM_14_) );
  ADDFX2 U136 ( .A(in_17bit_b[13]), .B(in_17bit_b[11]), .CI(
        add_2_root_r115_carry_14_), .CO(add_2_root_r115_carry_15_), .S(
        add_2_root_r115_SUM_14_) );
  ADDFX2 U137 ( .A(in_17bit_b[15]), .B(in_17bit_b[11]), .CI(
        add_1_root_r112_carry_15_), .CO(add_1_root_r112_carry_16_), .S(
        add_1_root_r112_SUM_15_) );
  ADDFX2 U138 ( .A(in_17bit_b[12]), .B(in_17bit_b[10]), .CI(
        add_1_root_r115_carry_16_), .CO(add_1_root_r115_carry_17_), .S(
        add_1_root_r115_SUM_16_) );
  ADDFX2 U139 ( .A(add_1_root_r119_A_16_), .B(in_17bit_b[10]), .CI(
        add_1_root_r119_carry[16]), .CO(add_1_root_r119_carry[17]), .S(
        add_1_root_r119_SUM_16_) );
  ADDFX2 U140 ( .A(in_17bit_b[11]), .B(in_17bit_b[10]), .CI(
        add_2_root_r119_carry_15_), .CO(add_2_root_r119_carry_16_), .S(
        add_2_root_r119_SUM_15_) );
  ADDFX2 U141 ( .A(in_17bit_b[14]), .B(in_17bit_b[12]), .CI(
        add_2_root_r115_carry_15_), .CO(add_2_root_r115_carry_16_), .S(
        add_2_root_r115_SUM_15_) );
  ADDFX2 U142 ( .A(in_17bit_b[13]), .B(in_17bit_b[11]), .CI(
        add_1_root_r115_carry_17_), .CO(add_1_root_r115_carry_18_), .S(
        add_1_root_r115_SUM_17_) );
  ADDFX2 U143 ( .A(add_1_root_r119_A_17_), .B(in_17bit_b[11]), .CI(
        add_1_root_r119_carry[17]), .CO(add_1_root_r119_carry[18]), .S(
        add_1_root_r119_SUM_17_) );
  ADDFX2 U144 ( .A(in_17bit_b[5]), .B(in_17bit_b[4]), .CI(
        add_3_root_r119_carry_6_), .CO(add_3_root_r119_carry_7_), .S(
        add_1_root_r119_A_6_) );
  ADDFX2 U145 ( .A(in_17bit_b[15]), .B(in_17bit_b[13]), .CI(
        add_2_root_r115_carry_16_), .CO(add_2_root_r115_carry_17_), .S(
        add_2_root_r115_SUM_16_) );
  ADDFX2 U146 ( .A(in_17bit_b[14]), .B(in_17bit_b[12]), .CI(
        add_1_root_r115_carry_18_), .CO(add_1_root_r115_carry_19_), .S(
        add_1_root_r115_SUM_18_) );
  ADDFX2 U147 ( .A(add_1_root_r119_A_18_), .B(in_17bit_b[12]), .CI(
        add_1_root_r119_carry[18]), .CO(add_1_root_r119_carry[19]), .S(
        add_1_root_r119_SUM_18_) );
  ADDFX2 U148 ( .A(in_17bit_b[15]), .B(in_17bit_b[13]), .CI(
        add_1_root_r115_carry_19_), .CO(add_1_root_r115_carry_20_), .S(
        add_1_root_r115_SUM_19_) );
  ADDFX2 U149 ( .A(in_17bit_b[5]), .B(in_17bit_b[3]), .CI(
        add_2_root_r115_carry_6_), .CO(add_2_root_r115_carry_7_), .S(
        add_2_root_r115_SUM_6_) );
  ADDFX2 U150 ( .A(in_17bit_b[7]), .B(in_17bit_b[3]), .CI(
        add_1_root_r112_carry_7_), .CO(add_1_root_r112_carry_8_), .S(
        add_1_root_r112_SUM_7_) );
  ADDFX2 U151 ( .A(in_17bit_b[14]), .B(in_17bit_b[13]), .CI(
        add_2_root_r119_carry_18_), .CO(add_2_root_r119_carry_19_), .S(
        add_2_root_r119_SUM_18_) );
  ADDFX2 U152 ( .A(in_17bit_b[5]), .B(in_17bit_b[3]), .CI(
        add_1_root_r115_carry_9_), .CO(add_1_root_r115_carry_10_), .S(
        add_1_root_r115_SUM_9_) );
  ADDFX2 U153 ( .A(add_1_root_r119_A_9_), .B(in_17bit_b[3]), .CI(
        add_1_root_r119_carry[9]), .CO(add_1_root_r119_carry[10]), .S(
        add_1_root_r119_SUM_9_) );
  ADDFX2 U154 ( .A(in_17bit_b[4]), .B(in_17bit_b[3]), .CI(
        add_2_root_r119_carry_8_), .CO(add_2_root_r119_carry_9_), .S(
        add_2_root_r119_SUM_8_) );
  ADDFX2 U155 ( .A(in_17bit_b[6]), .B(in_17bit_b[4]), .CI(
        add_1_root_r115_carry_10_), .CO(add_1_root_r115_carry_11_), .S(
        add_1_root_r115_SUM_10_) );
  ADDFX2 U156 ( .A(in_17bit_b[7]), .B(in_17bit_b[6]), .CI(
        add_2_root_r119_carry_11_), .CO(add_2_root_r119_carry_12_), .S(
        add_2_root_r119_SUM_11_) );
  ADDFX2 U157 ( .A(in_17bit_b[11]), .B(in_17bit_b[9]), .CI(
        add_2_root_r115_carry_12_), .CO(add_2_root_r115_carry_13_), .S(
        add_2_root_r115_SUM_12_) );
  ADDFX2 U158 ( .A(in_17bit_b[15]), .B(in_17bit_b[14]), .CI(
        add_3_root_r119_carry_16_), .CO(add_3_root_r119_carry_17_), .S(
        add_1_root_r119_A_16_) );
  ADDFX2 U159 ( .A(in_17bit_b[4]), .B(in_17bit_b[3]), .CI(
        add_3_root_r119_carry_5_), .CO(add_3_root_r119_carry_6_), .S(
        add_1_root_r119_A_5_) );
  ADDFX2 U160 ( .A(in_17bit_b[12]), .B(in_17bit_b[11]), .CI(
        add_2_root_r119_carry_16_), .CO(add_2_root_r119_carry_17_), .S(
        add_2_root_r119_SUM_16_) );
  ADDFX2 U161 ( .A(in_17bit_b[13]), .B(in_17bit_b[12]), .CI(
        add_2_root_r119_carry_17_), .CO(add_2_root_r119_carry_18_), .S(
        add_2_root_r119_SUM_17_) );
  ADDFX2 U162 ( .A(in_17bit_b[15]), .B(in_17bit_b[14]), .CI(
        add_2_root_r119_carry_19_), .CO(add_2_root_r119_carry_20_), .S(
        add_2_root_r119_SUM_19_) );
  INVX1 U163 ( .A(n21), .Y(n72) );
  XNOR2X1 U164 ( .A(n74), .B(n40), .Y(N29) );
  NAND2X1 U165 ( .A(sub_add_54_b0_carry[15]), .B(n175), .Y(n40) );
  CLKINVX3 U166 ( .A(n204), .Y(in_17bit_b[0]) );
  OAI21XL U167 ( .A0(n256), .A1(n257), .B0(n255), .Y(N463) );
  AOI22XL U168 ( .A0(N221), .A1(n254), .B0(N363), .B1(n253), .Y(n255) );
  INVX1 U169 ( .A(n177), .Y(n256) );
  CLKINVX3 U170 ( .A(n249), .Y(in_17bit_b[15]) );
  NAND2X1 U171 ( .A(n55), .B(in_8bit[1]), .Y(n92) );
  INVX1 U172 ( .A(in_8bit[0]), .Y(n64) );
  INVX1 U173 ( .A(in_8bit[2]), .Y(n66) );
  INVX1 U174 ( .A(in_8bit[5]), .Y(n67) );
  XNOR2X4 U175 ( .A(n41), .B(n3), .Y(out[12]) );
  MXI2XL U176 ( .A(n4), .B(n19), .S0(n91), .Y(out[16]) );
  AOI22XL U177 ( .A0(N28), .A1(n21), .B0(in_17bit[15]), .B1(n73), .Y(n249) );
  AOI22XL U178 ( .A0(N16), .A1(n21), .B0(in_17bit[3]), .B1(n72), .Y(n213) );
  AOI22XL U179 ( .A0(N17), .A1(n21), .B0(in_17bit[4]), .B1(n73), .Y(n216) );
  AOI22XL U180 ( .A0(N18), .A1(n21), .B0(in_17bit[5]), .B1(n73), .Y(n219) );
  AOI22XL U181 ( .A0(N19), .A1(n21), .B0(in_17bit[6]), .B1(n72), .Y(n222) );
  AOI22XL U182 ( .A0(N20), .A1(n21), .B0(in_17bit[7]), .B1(n73), .Y(n225) );
  AOI22XL U183 ( .A0(N21), .A1(n21), .B0(in_17bit[8]), .B1(n73), .Y(n228) );
  AOI22XL U184 ( .A0(N22), .A1(n21), .B0(in_17bit[9]), .B1(n72), .Y(n231) );
  AOI22XL U185 ( .A0(N23), .A1(n21), .B0(in_17bit[10]), .B1(n72), .Y(n234) );
  AOI22XL U186 ( .A0(N24), .A1(n21), .B0(in_17bit[11]), .B1(n72), .Y(n237) );
  AOI22XL U187 ( .A0(N25), .A1(n21), .B0(in_17bit[12]), .B1(n72), .Y(n240) );
  AOI22XL U188 ( .A0(N26), .A1(n21), .B0(in_17bit[13]), .B1(n73), .Y(n243) );
  NOR3X1 U189 ( .A(n66), .B(n178), .C(n64), .Y(n202) );
  AND2X2 U190 ( .A(n60), .B(n15), .Y(n42) );
  AND2X2 U191 ( .A(n42), .B(n18), .Y(n43) );
  AND2X2 U192 ( .A(n43), .B(n16), .Y(n44) );
  AND2X2 U193 ( .A(n44), .B(n17), .Y(n45) );
  NOR2X1 U194 ( .A(in_8bit[0]), .B(n98), .Y(n46) );
  AOI21X1 U195 ( .A0(n97), .A1(n39), .B0(n48), .Y(n47) );
  INVX1 U196 ( .A(n47), .Y(n253) );
  AND2X2 U197 ( .A(n46), .B(n57), .Y(n48) );
  AND2X2 U198 ( .A(n54), .B(n6), .Y(n49) );
  AOI21X1 U199 ( .A0(n57), .A1(n39), .B0(n51), .Y(n50) );
  INVX1 U200 ( .A(n50), .Y(n254) );
  AND2X2 U201 ( .A(n46), .B(n97), .Y(n51) );
  AND2X2 U202 ( .A(n45), .B(n11), .Y(n52) );
  AND2X2 U203 ( .A(n52), .B(n7), .Y(n53) );
  AND2X2 U204 ( .A(n53), .B(n8), .Y(n54) );
  OAI2BB1X1 U205 ( .A0N(n201), .A1N(n55), .B0(n99), .Y(n177) );
  NAND3BX1 U206 ( .AN(n98), .B(n202), .C(in_8bit[5]), .Y(n99) );
  AND3X1 U207 ( .A(n65), .B(n93), .C(n67), .Y(n55) );
  NOR2XL U208 ( .A(n65), .B(n93), .Y(n94) );
  AND2X2 U209 ( .A(n49), .B(n9), .Y(n56) );
  INVX1 U210 ( .A(in_17bit[3]), .Y(n160) );
  INVX1 U211 ( .A(in_17bit[4]), .Y(n161) );
  INVX1 U212 ( .A(in_17bit[5]), .Y(n162) );
  INVX1 U213 ( .A(in_17bit[6]), .Y(n163) );
  INVX1 U214 ( .A(in_17bit[7]), .Y(n164) );
  INVX1 U215 ( .A(in_17bit[8]), .Y(n167) );
  INVX1 U216 ( .A(in_17bit[9]), .Y(n168) );
  INVX1 U217 ( .A(in_17bit[10]), .Y(n170) );
  INVX1 U218 ( .A(in_17bit[11]), .Y(n171) );
  INVX1 U219 ( .A(in_17bit[12]), .Y(n172) );
  INVX1 U220 ( .A(in_17bit[13]), .Y(n173) );
  INVX1 U221 ( .A(in_17bit[14]), .Y(n174) );
  INVX1 U222 ( .A(in_17bit[15]), .Y(n175) );
  INVX1 U223 ( .A(in_17bit[1]), .Y(n101) );
  INVX1 U224 ( .A(in_17bit[2]), .Y(n158) );
  INVX1 U225 ( .A(in_17bit[0]), .Y(n100) );
  AND3X2 U226 ( .A(in_8bit[2]), .B(n178), .C(in_8bit[5]), .Y(n57) );
  INVX1 U227 ( .A(n77), .Y(n75) );
  NAND2X1 U228 ( .A(n206), .B(n205), .Y(N447) );
  AOI22X1 U229 ( .A0(N108), .A1(n250), .B0(N205), .B1(n254), .Y(n205) );
  AOI22X1 U230 ( .A0(N347), .A1(n253), .B0(n177), .B1(in_17bit_b[0]), .Y(n206)
         );
  NAND2X1 U231 ( .A(n209), .B(n208), .Y(N448) );
  AOI22X1 U232 ( .A0(N109), .A1(n250), .B0(N206), .B1(n254), .Y(n208) );
  AOI22X1 U233 ( .A0(N348), .A1(n253), .B0(n177), .B1(n176), .Y(n209) );
  INVX1 U234 ( .A(n207), .Y(n176) );
  NAND2X1 U235 ( .A(n212), .B(n211), .Y(N449) );
  AOI22X1 U236 ( .A0(N110), .A1(n250), .B0(N207), .B1(n254), .Y(n211) );
  AOI22X1 U237 ( .A0(N349), .A1(n253), .B0(n177), .B1(in_17bit_b[2]), .Y(n212)
         );
  NAND2X1 U238 ( .A(n215), .B(n214), .Y(N450) );
  AOI22X1 U239 ( .A0(N111), .A1(n250), .B0(N208), .B1(n254), .Y(n214) );
  AOI22X1 U240 ( .A0(N350), .A1(n253), .B0(n177), .B1(in_17bit_b[3]), .Y(n215)
         );
  NAND2X1 U241 ( .A(n218), .B(n217), .Y(N451) );
  AOI22X1 U242 ( .A0(N112), .A1(n250), .B0(N209), .B1(n254), .Y(n217) );
  AOI22X1 U243 ( .A0(N351), .A1(n253), .B0(n177), .B1(in_17bit_b[4]), .Y(n218)
         );
  NAND2X1 U244 ( .A(n221), .B(n220), .Y(N452) );
  AOI22X1 U245 ( .A0(N113), .A1(n250), .B0(N210), .B1(n254), .Y(n220) );
  AOI22X1 U246 ( .A0(N352), .A1(n253), .B0(n177), .B1(in_17bit_b[5]), .Y(n221)
         );
  NAND2X1 U247 ( .A(n224), .B(n223), .Y(N453) );
  AOI22X1 U248 ( .A0(N114), .A1(n250), .B0(N211), .B1(n254), .Y(n223) );
  AOI22X1 U249 ( .A0(N353), .A1(n253), .B0(n177), .B1(in_17bit_b[6]), .Y(n224)
         );
  NAND2X1 U250 ( .A(n227), .B(n226), .Y(N454) );
  AOI22X1 U251 ( .A0(N115), .A1(n250), .B0(N212), .B1(n254), .Y(n226) );
  AOI22X1 U252 ( .A0(N354), .A1(n253), .B0(n177), .B1(in_17bit_b[7]), .Y(n227)
         );
  NAND2X1 U253 ( .A(n230), .B(n229), .Y(N455) );
  AOI22X1 U254 ( .A0(N116), .A1(n250), .B0(N213), .B1(n254), .Y(n229) );
  NAND2X1 U255 ( .A(n233), .B(n232), .Y(N456) );
  AOI22X1 U256 ( .A0(N117), .A1(n250), .B0(N214), .B1(n254), .Y(n232) );
  NAND2X1 U257 ( .A(n236), .B(n235), .Y(N457) );
  AOI22X1 U258 ( .A0(N118), .A1(n250), .B0(N215), .B1(n254), .Y(n235) );
  NAND2X1 U259 ( .A(n239), .B(n238), .Y(N458) );
  AOI22X1 U260 ( .A0(N119), .A1(n250), .B0(N216), .B1(n254), .Y(n238) );
  NAND2X1 U261 ( .A(n242), .B(n241), .Y(N459) );
  NAND2X1 U262 ( .A(n245), .B(n244), .Y(N460) );
  NAND2X1 U263 ( .A(n248), .B(n247), .Y(N461) );
  NAND2X1 U264 ( .A(n252), .B(n251), .Y(N462) );
  XNOR2X1 U265 ( .A(n13), .B(sub_add_75_b0_carry[13]), .Y(n58) );
  NAND4BBX1 U266 ( .AN(n253), .BN(n254), .C(n203), .D(n256), .Y(N446) );
  NOR4BX1 U267 ( .AN(n200), .B(n64), .C(in_8bit[1]), .D(in_8bit[2]), .Y(n201)
         );
  NOR2X1 U268 ( .A(in_8bit[6]), .B(in_8bit[3]), .Y(n200) );
  NOR2X1 U269 ( .A(out[0]), .B(neg_mul[8]), .Y(n59) );
  NOR2BX1 U270 ( .AN(n59), .B(neg_mul[9]), .Y(n60) );
  NAND4BXL U271 ( .AN(n65), .B(in_8bit[6]), .C(in_8bit[1]), .D(in_8bit[4]), 
        .Y(n98) );
  NAND2X1 U272 ( .A(n96), .B(n95), .Y(n250) );
  NAND3BX1 U273 ( .AN(n92), .B(n202), .C(in_8bit[6]), .Y(n96) );
  NAND3X1 U274 ( .A(n201), .B(in_8bit[5]), .C(n94), .Y(n95) );
  NAND2X1 U275 ( .A(out[0]), .B(neg_mul[8]), .Y(n77) );
  INVX1 U276 ( .A(n199), .Y(n97) );
  NAND3BX1 U277 ( .AN(in_8bit[5]), .B(n66), .C(in_8bit[3]), .Y(n199) );
  NOR2X1 U278 ( .A(in_8bit[6]), .B(in_8bit[4]), .Y(n198) );
  NAND2X1 U279 ( .A(sub_add_75_b0_carry[15]), .B(n10), .Y(n61) );
  INVX1 U280 ( .A(in_8bit[4]), .Y(n93) );
  INVX1 U281 ( .A(in_8bit[3]), .Y(n178) );
  NOR2X2 U282 ( .A(n90), .B(n49), .Y(n89) );
  XOR2X4 U283 ( .A(n79), .B(neg_mul[9]), .Y(out[2]) );
  NAND2XL U284 ( .A(N29), .B(n71), .Y(n257) );
  AOI22XL U285 ( .A0(N15), .A1(n71), .B0(in_17bit[2]), .B1(n73), .Y(n210) );
  AOI22XL U286 ( .A0(N14), .A1(n71), .B0(in_17bit[1]), .B1(n73), .Y(n207) );
  AOI22XL U287 ( .A0(in_17bit[0]), .A1(n71), .B0(in_17bit[0]), .B1(n73), .Y(
        n204) );
  NOR2X2 U288 ( .A(n53), .B(n88), .Y(n87) );
  NOR2X4 U289 ( .A(n44), .B(n88), .Y(n85) );
  XNOR2X4 U290 ( .A(n87), .B(n8), .Y(out[9]) );
  XNOR2X4 U291 ( .A(n89), .B(n9), .Y(out[11]) );
  MXI2X4 U292 ( .A(n13), .B(n58), .S0(n91), .Y(out[13]) );
  AND2X1 U293 ( .A(add_1_root_r112_carry_20_), .B(in_17bit_b[16]), .Y(
        add_1_root_r112_SUM_21_) );
  XOR2X1 U294 ( .A(in_17bit_b[16]), .B(add_1_root_r112_carry_20_), .Y(
        add_1_root_r112_SUM_20_) );
  AND2X1 U295 ( .A(add_1_root_r112_carry_19_), .B(in_17bit_b[15]), .Y(
        add_1_root_r112_carry_20_) );
  XOR2X1 U296 ( .A(in_17bit_b[15]), .B(add_1_root_r112_carry_19_), .Y(
        add_1_root_r112_SUM_19_) );
  AND2X1 U297 ( .A(add_1_root_r112_carry_18_), .B(in_17bit_b[14]), .Y(
        add_1_root_r112_carry_19_) );
  XOR2X1 U298 ( .A(in_17bit_b[14]), .B(add_1_root_r112_carry_18_), .Y(
        add_1_root_r112_SUM_18_) );
  AND2X1 U299 ( .A(add_1_root_r112_carry_17_), .B(in_17bit_b[13]), .Y(
        add_1_root_r112_carry_18_) );
  XOR2X1 U300 ( .A(in_17bit_b[13]), .B(add_1_root_r112_carry_17_), .Y(
        add_1_root_r112_SUM_17_) );
  AND2X1 U301 ( .A(add_2_root_r119_carry_21_), .B(in_17bit_b[16]), .Y(
        add_2_root_r119_SUM_22_) );
  XOR2X1 U302 ( .A(in_17bit_b[16]), .B(add_2_root_r119_carry_21_), .Y(
        add_2_root_r119_SUM_21_) );
  AND2X1 U303 ( .A(n176), .B(in_17bit_b[0]), .Y(add_2_root_r119_carry_6_) );
  XOR2X1 U304 ( .A(in_17bit_b[0]), .B(n176), .Y(add_2_root_r119_SUM_5_) );
  AND2X1 U305 ( .A(add_1_root_r119_carry[22]), .B(in_17bit_b[16]), .Y(
        add_1_root_r119_SUM_23_) );
  XOR2X1 U306 ( .A(in_17bit_b[16]), .B(add_1_root_r119_carry[22]), .Y(
        add_1_root_r119_SUM_22_) );
  AND2X1 U307 ( .A(add_1_root_r119_carry[21]), .B(in_17bit_b[15]), .Y(
        add_1_root_r119_carry[22]) );
  XOR2X1 U308 ( .A(in_17bit_b[15]), .B(add_1_root_r119_carry[21]), .Y(
        add_1_root_r119_SUM_21_) );
  AND2X1 U309 ( .A(add_1_root_r119_carry[20]), .B(in_17bit_b[14]), .Y(
        add_1_root_r119_carry[21]) );
  XOR2X1 U310 ( .A(in_17bit_b[14]), .B(add_1_root_r119_carry[20]), .Y(
        add_1_root_r119_SUM_20_) );
  AND2X1 U311 ( .A(add_1_root_r119_A_6_), .B(in_17bit_b[0]), .Y(
        add_1_root_r119_carry[7]) );
  XOR2X1 U312 ( .A(in_17bit_b[0]), .B(add_1_root_r119_A_6_), .Y(
        add_1_root_r119_SUM_6_) );
  AND2X1 U313 ( .A(add_3_root_r119_carry_18_), .B(in_17bit_b[16]), .Y(
        add_1_root_r119_A_19_) );
  XOR2X1 U314 ( .A(in_17bit_b[16]), .B(add_3_root_r119_carry_18_), .Y(
        add_1_root_r119_A_18_) );
  AND2X1 U315 ( .A(add_2_root_r115_carry_19_), .B(in_17bit_b[16]), .Y(
        add_2_root_r115_SUM_20_) );
  XOR2X1 U316 ( .A(in_17bit_b[16]), .B(add_2_root_r115_carry_19_), .Y(
        add_2_root_r115_SUM_19_) );
  AND2X1 U317 ( .A(add_2_root_r115_carry_18_), .B(in_17bit_b[15]), .Y(
        add_2_root_r115_carry_19_) );
  XOR2X1 U318 ( .A(in_17bit_b[15]), .B(add_2_root_r115_carry_18_), .Y(
        add_2_root_r115_SUM_18_) );
  AND2X1 U319 ( .A(in_17bit_b[2]), .B(in_17bit_b[0]), .Y(
        add_2_root_r115_carry_4_) );
  AND2X1 U320 ( .A(add_1_root_r115_carry_22_), .B(in_17bit_b[16]), .Y(
        add_1_root_r115_SUM_23_) );
  XOR2X1 U321 ( .A(in_17bit_b[16]), .B(add_1_root_r115_carry_22_), .Y(
        add_1_root_r115_SUM_22_) );
  AND2X1 U322 ( .A(add_1_root_r115_carry_21_), .B(in_17bit_b[15]), .Y(
        add_1_root_r115_carry_22_) );
  XOR2X1 U323 ( .A(in_17bit_b[15]), .B(add_1_root_r115_carry_21_), .Y(
        add_1_root_r115_SUM_21_) );
  XOR2X1 U324 ( .A(in_17bit_b[0]), .B(in_17bit_b[2]), .Y(
        add_1_root_r115_SUM_6_) );
  XOR2X1 U325 ( .A(n175), .B(sub_add_54_b0_carry[15]), .Y(N28) );
  AND2X1 U326 ( .A(sub_add_54_b0_carry[14]), .B(n174), .Y(
        sub_add_54_b0_carry[15]) );
  XOR2X1 U327 ( .A(n174), .B(sub_add_54_b0_carry[14]), .Y(N27) );
  AND2X1 U328 ( .A(sub_add_54_b0_carry[13]), .B(n173), .Y(
        sub_add_54_b0_carry[14]) );
  XOR2X1 U329 ( .A(n173), .B(sub_add_54_b0_carry[13]), .Y(N26) );
  AND2X1 U330 ( .A(sub_add_54_b0_carry[12]), .B(n172), .Y(
        sub_add_54_b0_carry[13]) );
  XOR2X1 U331 ( .A(n172), .B(sub_add_54_b0_carry[12]), .Y(N25) );
  AND2X1 U332 ( .A(sub_add_54_b0_carry[11]), .B(n171), .Y(
        sub_add_54_b0_carry[12]) );
  XOR2X1 U333 ( .A(n171), .B(sub_add_54_b0_carry[11]), .Y(N24) );
  AND2X1 U334 ( .A(sub_add_54_b0_carry[10]), .B(n170), .Y(
        sub_add_54_b0_carry[11]) );
  XOR2X1 U335 ( .A(n170), .B(sub_add_54_b0_carry[10]), .Y(N23) );
  AND2X1 U336 ( .A(sub_add_54_b0_carry[9]), .B(n168), .Y(
        sub_add_54_b0_carry[10]) );
  XOR2X1 U337 ( .A(n168), .B(sub_add_54_b0_carry[9]), .Y(N22) );
  AND2X1 U338 ( .A(sub_add_54_b0_carry[8]), .B(n167), .Y(
        sub_add_54_b0_carry[9]) );
  XOR2X1 U339 ( .A(n167), .B(sub_add_54_b0_carry[8]), .Y(N21) );
  AND2X1 U340 ( .A(sub_add_54_b0_carry[7]), .B(n164), .Y(
        sub_add_54_b0_carry[8]) );
  XOR2X1 U341 ( .A(n164), .B(sub_add_54_b0_carry[7]), .Y(N20) );
  AND2X1 U342 ( .A(sub_add_54_b0_carry[6]), .B(n163), .Y(
        sub_add_54_b0_carry[7]) );
  XOR2X1 U343 ( .A(n163), .B(sub_add_54_b0_carry[6]), .Y(N19) );
  AND2X1 U344 ( .A(sub_add_54_b0_carry[5]), .B(n162), .Y(
        sub_add_54_b0_carry[6]) );
  XOR2X1 U345 ( .A(n162), .B(sub_add_54_b0_carry[5]), .Y(N18) );
  AND2X1 U346 ( .A(sub_add_54_b0_carry[4]), .B(n161), .Y(
        sub_add_54_b0_carry[5]) );
  XOR2X1 U347 ( .A(n161), .B(sub_add_54_b0_carry[4]), .Y(N17) );
  AND2X1 U348 ( .A(sub_add_54_b0_carry[3]), .B(n160), .Y(
        sub_add_54_b0_carry[4]) );
  XOR2X1 U349 ( .A(n160), .B(sub_add_54_b0_carry[3]), .Y(N16) );
  AND2X1 U350 ( .A(sub_add_54_b0_carry[2]), .B(n158), .Y(
        sub_add_54_b0_carry[3]) );
  XOR2X1 U351 ( .A(n158), .B(sub_add_54_b0_carry[2]), .Y(N15) );
  AND2X1 U352 ( .A(n100), .B(n101), .Y(sub_add_54_b0_carry[2]) );
  XOR2X1 U353 ( .A(n101), .B(n100), .Y(N14) );
  XOR2X1 U354 ( .A(n10), .B(sub_add_75_b0_carry[15]), .Y(N480) );
  AND2X1 U355 ( .A(sub_add_75_b0_carry[14]), .B(n36), .Y(
        sub_add_75_b0_carry[15]) );
  AND2X1 U356 ( .A(sub_add_75_b0_carry[13]), .B(n13), .Y(
        sub_add_75_b0_carry[14]) );
  AND2X1 U357 ( .A(n56), .B(n12), .Y(sub_add_75_b0_carry[13]) );
  AND2X1 U358 ( .A(in_17bit_b[0]), .B(in_17bit_b[4]), .Y(
        add_1_root_r112_carry_5_) );
endmodule


module multi16_6_DW01_add_0 ( A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, 
        A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, 
        A_4_, B_23_, B_22_, B_21_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, 
        B_14_, B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, 
        SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, 
        SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, 
        SUM_7_ );
  input A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_,
         A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, B_23_, B_22_,
         B_21_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_,
         B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_;
  output SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_,
         SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_,
         SUM_8_, SUM_7_;
  wire   n1, n2, n3, n4;
  wire   [23:7] carry;

  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry[7]), .CO(carry[8]), .S(SUM_7_)
         );
  ADDFX2 U1_21 ( .A(A_21_), .B(B_21_), .CI(carry[21]), .CO(carry[22]), .S(
        SUM_21_) );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry[20]), .CO(carry[21]), .S(
        SUM_20_) );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry[19]), .CO(carry[20]), .S(
        SUM_19_) );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry[18]), .CO(carry[19]), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry[17]), .CO(carry[18]), .S(
        SUM_17_) );
  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry[16]), .CO(carry[17]), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry[15]), .CO(carry[16]), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry[14]), .CO(carry[15]), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry[13]), .CO(carry[14]), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry[12]), .CO(carry[13]), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry[11]), .CO(carry[12]), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry[10]), .CO(carry[11]), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry[9]), .CO(carry[10]), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry[8]), .CO(carry[9]), .S(SUM_8_)
         );
  ADDFX2 U1_22 ( .A(A_22_), .B(B_22_), .CI(carry[22]), .CO(carry[23]), .S(
        SUM_22_) );
  AND2X2 U1 ( .A(A_4_), .B(B_4_), .Y(n1) );
  XOR2X1 U2 ( .A(B_23_), .B(carry[23]), .Y(SUM_23_) );
  OAI2BB1X1 U3 ( .A0N(n2), .A1N(A_6_), .B0(n3), .Y(carry[7]) );
  OAI21XL U4 ( .A0(A_6_), .A1(n2), .B0(B_6_), .Y(n3) );
  OAI2BB1X1 U5 ( .A0N(n1), .A1N(A_5_), .B0(n4), .Y(n2) );
  OAI21XL U6 ( .A0(A_5_), .A1(n1), .B0(B_5_), .Y(n4) );
endmodule


module multi16_6_DW01_add_4 ( A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, 
        A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, 
        B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, 
        B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, SUM_22_, SUM_21_, SUM_20_, 
        SUM_19_, SUM_18_, SUM_17_, SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, 
        SUM_11_, SUM_10_, SUM_9_, SUM_8_, SUM_7_ );
  input A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_,
         A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, B_20_, B_19_,
         B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, B_10_, B_9_,
         B_8_, B_7_, B_6_, B_5_;
  output SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_,
         SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_,
         SUM_7_;
  wire   carry_21_, carry_20_, carry_19_, carry_18_, carry_17_, carry_16_,
         carry_15_, carry_14_, carry_13_, carry_12_, carry_11_, carry_10_,
         carry_9_, carry_8_, carry_7_, n1;

  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry_16_), .CO(carry_17_), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry_15_), .CO(carry_16_), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry_14_), .CO(carry_15_), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry_13_), .CO(carry_14_), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry_12_), .CO(carry_13_), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry_11_), .CO(carry_12_), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry_10_), .CO(carry_11_), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry_9_), .CO(carry_10_), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry_8_), .CO(carry_9_), .S(SUM_8_)
         );
  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry_7_), .CO(carry_8_), .S(SUM_7_)
         );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry_20_), .CO(carry_21_), .S(
        SUM_20_) );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry_19_), .CO(carry_20_), .S(
        SUM_19_) );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry_18_), .CO(carry_19_), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry_17_), .CO(carry_18_), .S(
        SUM_17_) );
  ADDFX2 U1_21 ( .A(A_21_), .B(B_21_), .CI(carry_21_), .CO(SUM_22_), .S(
        SUM_21_) );
  OAI2BB1X1 U1 ( .A0N(A_6_), .A1N(B_6_), .B0(n1), .Y(carry_7_) );
  OAI211X1 U2 ( .A0(B_6_), .A1(A_6_), .B0(A_5_), .C0(B_5_), .Y(n1) );
endmodule


module multi16_6_DW01_add_6 ( A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, 
        A_16_, A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, 
        A_6_, A_5_, A_4_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, 
        B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, 
        SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, 
        SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, 
        SUM_7_ );
  input A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_,
         A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, B_20_,
         B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, B_10_,
         B_9_, B_8_, B_7_, B_6_, B_5_, B_4_;
  output SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_,
         SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_,
         SUM_8_, SUM_7_;
  wire   n1, n2, n3, n4, n5, n6;
  wire   [21:7] carry;

  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry[7]), .CO(carry[8]), .S(SUM_7_)
         );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry[18]), .CO(carry[19]), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry[17]), .CO(carry[18]), .S(
        SUM_17_) );
  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry[16]), .CO(carry[17]), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry[15]), .CO(carry[16]), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry[14]), .CO(carry[15]), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry[13]), .CO(carry[14]), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry[12]), .CO(carry[13]), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry[11]), .CO(carry[12]), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry[10]), .CO(carry[11]), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry[9]), .CO(carry[10]), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry[8]), .CO(carry[9]), .S(SUM_8_)
         );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry[19]), .CO(carry[20]), .S(
        SUM_19_) );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry[20]), .CO(carry[21]), .S(
        SUM_20_) );
  AND2X2 U1 ( .A(A_22_), .B(n2), .Y(n1) );
  AND2X2 U2 ( .A(A_21_), .B(carry[21]), .Y(n2) );
  AND2X2 U3 ( .A(A_4_), .B(B_4_), .Y(n3) );
  XOR2X1 U4 ( .A(A_23_), .B(n1), .Y(SUM_23_) );
  XOR2X1 U5 ( .A(A_21_), .B(carry[21]), .Y(SUM_21_) );
  XOR2X1 U6 ( .A(A_22_), .B(n2), .Y(SUM_22_) );
  OAI2BB1X1 U7 ( .A0N(n4), .A1N(A_6_), .B0(n5), .Y(carry[7]) );
  OAI21XL U8 ( .A0(A_6_), .A1(n4), .B0(B_6_), .Y(n5) );
  OAI2BB1X1 U9 ( .A0N(n3), .A1N(A_5_), .B0(n6), .Y(n4) );
  OAI21XL U10 ( .A0(A_5_), .A1(n3), .B0(B_5_), .Y(n6) );
endmodule


module multi16_6 ( in_17bit, in_8bit, out );
  input [16:0] in_17bit;
  input [7:0] in_8bit;
  output [16:0] out;
  wire   n286, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26,
         N27, N28, N29, N108, N109, N110, N111, N112, N113, N114, N115, N116,
         N117, N118, N119, N120, N121, N122, N123, N205, N206, N207, N208,
         N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, N219,
         N220, N221, N347, N348, N349, N350, N351, N352, N353, N354, N355,
         N356, N357, N358, N359, N360, N361, N362, N363, N446, N447, N448,
         N449, N450, N451, N452, N453, N454, N455, N456, N457, N458, N459,
         N460, N461, N462, N463, N479, N480, N481, add_2_root_r119_carry_10_,
         add_2_root_r119_carry_11_, add_2_root_r119_carry_12_,
         add_2_root_r119_carry_13_, add_2_root_r119_carry_14_,
         add_2_root_r119_carry_15_, add_2_root_r119_carry_16_,
         add_2_root_r119_carry_17_, add_2_root_r119_carry_18_,
         add_2_root_r119_carry_19_, add_2_root_r119_carry_20_,
         add_2_root_r119_carry_21_, add_2_root_r119_carry_7_,
         add_2_root_r119_carry_8_, add_2_root_r119_carry_9_,
         add_2_root_r119_SUM_5_, add_2_root_r119_SUM_6_,
         add_2_root_r119_SUM_7_, add_2_root_r119_SUM_8_,
         add_2_root_r119_SUM_9_, add_2_root_r119_SUM_10_,
         add_2_root_r119_SUM_11_, add_2_root_r119_SUM_12_,
         add_2_root_r119_SUM_13_, add_2_root_r119_SUM_14_,
         add_2_root_r119_SUM_15_, add_2_root_r119_SUM_16_,
         add_2_root_r119_SUM_17_, add_2_root_r119_SUM_18_,
         add_2_root_r119_SUM_19_, add_2_root_r119_SUM_20_,
         add_2_root_r119_SUM_21_, add_2_root_r119_SUM_22_,
         add_1_root_r119_SUM_6_, add_1_root_r119_SUM_7_,
         add_1_root_r119_SUM_8_, add_1_root_r119_SUM_9_,
         add_1_root_r119_SUM_10_, add_1_root_r119_SUM_11_,
         add_1_root_r119_SUM_12_, add_1_root_r119_SUM_13_,
         add_1_root_r119_SUM_14_, add_1_root_r119_SUM_15_,
         add_1_root_r119_SUM_16_, add_1_root_r119_SUM_17_,
         add_1_root_r119_SUM_18_, add_1_root_r119_SUM_19_,
         add_1_root_r119_SUM_20_, add_1_root_r119_SUM_21_,
         add_1_root_r119_SUM_22_, add_1_root_r119_SUM_23_,
         add_1_root_r119_A_3_, add_1_root_r119_A_4_, add_1_root_r119_A_5_,
         add_1_root_r119_A_6_, add_1_root_r119_A_7_, add_1_root_r119_A_8_,
         add_1_root_r119_A_9_, add_1_root_r119_A_10_, add_1_root_r119_A_11_,
         add_1_root_r119_A_12_, add_1_root_r119_A_13_, add_1_root_r119_A_14_,
         add_1_root_r119_A_15_, add_1_root_r119_A_16_, add_1_root_r119_A_17_,
         add_1_root_r119_A_18_, add_1_root_r119_A_19_,
         add_3_root_r119_carry_10_, add_3_root_r119_carry_11_,
         add_3_root_r119_carry_12_, add_3_root_r119_carry_13_,
         add_3_root_r119_carry_14_, add_3_root_r119_carry_15_,
         add_3_root_r119_carry_16_, add_3_root_r119_carry_17_,
         add_3_root_r119_carry_18_, add_3_root_r119_carry_3_,
         add_3_root_r119_carry_4_, add_3_root_r119_carry_5_,
         add_3_root_r119_carry_6_, add_3_root_r119_carry_7_,
         add_3_root_r119_carry_8_, add_3_root_r119_carry_9_,
         add_1_root_r112_carry_10_, add_1_root_r112_carry_11_,
         add_1_root_r112_carry_12_, add_1_root_r112_carry_13_,
         add_1_root_r112_carry_14_, add_1_root_r112_carry_15_,
         add_1_root_r112_carry_16_, add_1_root_r112_carry_17_,
         add_1_root_r112_carry_18_, add_1_root_r112_carry_19_,
         add_1_root_r112_carry_20_, add_1_root_r112_carry_5_,
         add_1_root_r112_carry_6_, add_1_root_r112_carry_7_,
         add_1_root_r112_carry_8_, add_1_root_r112_carry_9_,
         add_1_root_r112_SUM_1_, add_1_root_r112_SUM_2_,
         add_1_root_r112_SUM_3_, add_1_root_r112_SUM_4_,
         add_1_root_r112_SUM_5_, add_1_root_r112_SUM_6_,
         add_1_root_r112_SUM_7_, add_1_root_r112_SUM_8_,
         add_1_root_r112_SUM_9_, add_1_root_r112_SUM_10_,
         add_1_root_r112_SUM_11_, add_1_root_r112_SUM_12_,
         add_1_root_r112_SUM_13_, add_1_root_r112_SUM_14_,
         add_1_root_r112_SUM_15_, add_1_root_r112_SUM_16_,
         add_1_root_r112_SUM_17_, add_1_root_r112_SUM_18_,
         add_1_root_r112_SUM_19_, add_1_root_r112_SUM_20_,
         add_1_root_r112_SUM_21_, add_2_root_r115_carry_10_,
         add_2_root_r115_carry_11_, add_2_root_r115_carry_12_,
         add_2_root_r115_carry_13_, add_2_root_r115_carry_14_,
         add_2_root_r115_carry_15_, add_2_root_r115_carry_16_,
         add_2_root_r115_carry_17_, add_2_root_r115_carry_18_,
         add_2_root_r115_carry_19_, add_2_root_r115_carry_4_,
         add_2_root_r115_carry_5_, add_2_root_r115_carry_6_,
         add_2_root_r115_carry_7_, add_2_root_r115_carry_8_,
         add_2_root_r115_carry_9_, add_2_root_r115_SUM_3_,
         add_2_root_r115_SUM_4_, add_2_root_r115_SUM_5_,
         add_2_root_r115_SUM_6_, add_2_root_r115_SUM_7_,
         add_2_root_r115_SUM_8_, add_2_root_r115_SUM_9_,
         add_2_root_r115_SUM_10_, add_2_root_r115_SUM_11_,
         add_2_root_r115_SUM_12_, add_2_root_r115_SUM_13_,
         add_2_root_r115_SUM_14_, add_2_root_r115_SUM_15_,
         add_2_root_r115_SUM_16_, add_2_root_r115_SUM_17_,
         add_2_root_r115_SUM_18_, add_2_root_r115_SUM_19_,
         add_2_root_r115_SUM_20_, add_1_root_r115_carry_10_,
         add_1_root_r115_carry_11_, add_1_root_r115_carry_12_,
         add_1_root_r115_carry_13_, add_1_root_r115_carry_14_,
         add_1_root_r115_carry_15_, add_1_root_r115_carry_16_,
         add_1_root_r115_carry_17_, add_1_root_r115_carry_18_,
         add_1_root_r115_carry_19_, add_1_root_r115_carry_20_,
         add_1_root_r115_carry_21_, add_1_root_r115_carry_22_,
         add_1_root_r115_carry_8_, add_1_root_r115_carry_9_,
         add_1_root_r115_SUM_7_, add_1_root_r115_SUM_8_,
         add_1_root_r115_SUM_9_, add_1_root_r115_SUM_10_,
         add_1_root_r115_SUM_11_, add_1_root_r115_SUM_12_,
         add_1_root_r115_SUM_13_, add_1_root_r115_SUM_14_,
         add_1_root_r115_SUM_15_, add_1_root_r115_SUM_16_,
         add_1_root_r115_SUM_17_, add_1_root_r115_SUM_18_,
         add_1_root_r115_SUM_19_, add_1_root_r115_SUM_20_,
         add_1_root_r115_SUM_21_, add_1_root_r115_SUM_22_,
         add_1_root_r115_SUM_23_, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n158, n160, n163, n164, n167, n168, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285;
  wire   [16:0] in_17bit_b;
  wire   [23:8] neg_mul;
  wire   [16:13] sub_add_75_b0_carry;
  wire   [16:2] sub_add_54_b0_carry;
  wire   [22:7] add_1_root_r119_carry;

  multi16_6_DW01_add_0 add_0_root_r119 ( .A_22_(add_2_root_r119_SUM_22_), 
        .A_21_(add_2_root_r119_SUM_21_), .A_20_(add_2_root_r119_SUM_20_), 
        .A_19_(add_2_root_r119_SUM_19_), .A_18_(add_2_root_r119_SUM_18_), 
        .A_17_(add_2_root_r119_SUM_17_), .A_16_(add_2_root_r119_SUM_16_), 
        .A_15_(add_2_root_r119_SUM_15_), .A_14_(add_2_root_r119_SUM_14_), 
        .A_13_(add_2_root_r119_SUM_13_), .A_12_(add_2_root_r119_SUM_12_), 
        .A_11_(add_2_root_r119_SUM_11_), .A_10_(add_2_root_r119_SUM_10_), 
        .A_9_(add_2_root_r119_SUM_9_), .A_8_(add_2_root_r119_SUM_8_), .A_7_(
        add_2_root_r119_SUM_7_), .A_6_(add_2_root_r119_SUM_6_), .A_5_(
        add_2_root_r119_SUM_5_), .A_4_(in_17bit_b[0]), .B_23_(
        add_1_root_r119_SUM_23_), .B_22_(add_1_root_r119_SUM_22_), .B_21_(
        add_1_root_r119_SUM_21_), .B_20_(add_1_root_r119_SUM_20_), .B_19_(
        add_1_root_r119_SUM_19_), .B_18_(add_1_root_r119_SUM_18_), .B_17_(
        add_1_root_r119_SUM_17_), .B_16_(add_1_root_r119_SUM_16_), .B_15_(
        add_1_root_r119_SUM_15_), .B_14_(add_1_root_r119_SUM_14_), .B_13_(
        add_1_root_r119_SUM_13_), .B_12_(add_1_root_r119_SUM_12_), .B_11_(
        add_1_root_r119_SUM_11_), .B_10_(add_1_root_r119_SUM_10_), .B_9_(
        add_1_root_r119_SUM_9_), .B_8_(add_1_root_r119_SUM_8_), .B_7_(
        add_1_root_r119_SUM_7_), .B_6_(add_1_root_r119_SUM_6_), .B_5_(
        add_1_root_r119_A_5_), .B_4_(add_1_root_r119_A_4_), .SUM_23_(N363), 
        .SUM_22_(N362), .SUM_21_(N361), .SUM_20_(N360), .SUM_19_(N359), 
        .SUM_18_(N358), .SUM_17_(N357), .SUM_16_(N356), .SUM_15_(N355), 
        .SUM_14_(N354), .SUM_13_(N353), .SUM_12_(N352), .SUM_11_(N351), 
        .SUM_10_(N350), .SUM_9_(N349), .SUM_8_(N348), .SUM_7_(N347) );
  multi16_6_DW01_add_4 add_0_root_r112 ( .A_21_(in_17bit_b[16]), .A_20_(
        in_17bit_b[15]), .A_19_(in_17bit_b[14]), .A_18_(in_17bit_b[13]), 
        .A_17_(in_17bit_b[12]), .A_16_(in_17bit_b[11]), .A_15_(in_17bit_b[10]), 
        .A_14_(in_17bit_b[9]), .A_13_(in_17bit_b[8]), .A_12_(in_17bit_b[7]), 
        .A_11_(in_17bit_b[6]), .A_10_(in_17bit_b[5]), .A_9_(in_17bit_b[4]), 
        .A_8_(in_17bit_b[3]), .A_7_(in_17bit_b[2]), .A_6_(n202), .A_5_(
        in_17bit_b[0]), .B_21_(add_1_root_r112_SUM_21_), .B_20_(
        add_1_root_r112_SUM_20_), .B_19_(add_1_root_r112_SUM_19_), .B_18_(
        add_1_root_r112_SUM_18_), .B_17_(add_1_root_r112_SUM_17_), .B_16_(
        add_1_root_r112_SUM_16_), .B_15_(add_1_root_r112_SUM_15_), .B_14_(
        add_1_root_r112_SUM_14_), .B_13_(add_1_root_r112_SUM_13_), .B_12_(
        add_1_root_r112_SUM_12_), .B_11_(add_1_root_r112_SUM_11_), .B_10_(
        add_1_root_r112_SUM_10_), .B_9_(add_1_root_r112_SUM_9_), .B_8_(
        add_1_root_r112_SUM_8_), .B_7_(add_1_root_r112_SUM_7_), .B_6_(
        add_1_root_r112_SUM_6_), .B_5_(add_1_root_r112_SUM_5_), .SUM_22_(N123), 
        .SUM_21_(N122), .SUM_20_(N121), .SUM_19_(N120), .SUM_18_(N119), 
        .SUM_17_(N118), .SUM_16_(N117), .SUM_15_(N116), .SUM_14_(N115), 
        .SUM_13_(N114), .SUM_12_(N113), .SUM_11_(N112), .SUM_10_(N111), 
        .SUM_9_(N110), .SUM_8_(N109), .SUM_7_(N108) );
  multi16_6_DW01_add_6 add_0_root_r115 ( .A_23_(add_1_root_r115_SUM_23_), 
        .A_22_(add_1_root_r115_SUM_22_), .A_21_(add_1_root_r115_SUM_21_), 
        .A_20_(add_1_root_r115_SUM_20_), .A_19_(add_1_root_r115_SUM_19_), 
        .A_18_(add_1_root_r115_SUM_18_), .A_17_(add_1_root_r115_SUM_17_), 
        .A_16_(add_1_root_r115_SUM_16_), .A_15_(add_1_root_r115_SUM_15_), 
        .A_14_(add_1_root_r115_SUM_14_), .A_13_(add_1_root_r115_SUM_13_), 
        .A_12_(add_1_root_r115_SUM_12_), .A_11_(add_1_root_r115_SUM_11_), 
        .A_10_(add_1_root_r115_SUM_10_), .A_9_(add_1_root_r115_SUM_9_), .A_8_(
        add_1_root_r115_SUM_8_), .A_7_(add_1_root_r115_SUM_7_), .A_6_(
        add_2_root_r115_SUM_3_), .A_5_(n202), .A_4_(in_17bit_b[0]), .B_20_(
        add_2_root_r115_SUM_20_), .B_19_(add_2_root_r115_SUM_19_), .B_18_(
        add_2_root_r115_SUM_18_), .B_17_(add_2_root_r115_SUM_17_), .B_16_(
        add_2_root_r115_SUM_16_), .B_15_(add_2_root_r115_SUM_15_), .B_14_(
        add_2_root_r115_SUM_14_), .B_13_(add_2_root_r115_SUM_13_), .B_12_(
        add_2_root_r115_SUM_12_), .B_11_(add_2_root_r115_SUM_11_), .B_10_(
        add_2_root_r115_SUM_10_), .B_9_(add_2_root_r115_SUM_9_), .B_8_(
        add_2_root_r115_SUM_8_), .B_7_(add_2_root_r115_SUM_7_), .B_6_(
        add_2_root_r115_SUM_6_), .B_5_(add_2_root_r115_SUM_5_), .B_4_(
        add_2_root_r115_SUM_4_), .SUM_23_(N221), .SUM_22_(N220), .SUM_21_(N219), .SUM_20_(N218), .SUM_19_(N217), .SUM_18_(N216), .SUM_17_(N215), .SUM_16_(
        N214), .SUM_15_(N213), .SUM_14_(N212), .SUM_13_(N211), .SUM_12_(N210), 
        .SUM_11_(N209), .SUM_10_(N208), .SUM_9_(N207), .SUM_8_(N206), .SUM_7_(
        N205) );
  TLATX1 neg_mul_reg_19_ ( .G(N446), .D(N459), .QN(n4) );
  TLATX1 neg_mul_reg_18_ ( .G(N446), .D(N458), .QN(n3) );
  TLATX1 neg_mul_reg_16_ ( .G(N446), .D(N456), .Q(neg_mul[16]), .QN(n1) );
  TLATX1 neg_mul_reg_15_ ( .G(N446), .D(N455), .Q(neg_mul[15]), .QN(n2) );
  TLATX1 neg_mul_reg_23_ ( .G(N446), .D(N463), .Q(neg_mul[23]), .QN(n17) );
  TLATX1 neg_mul_reg_22_ ( .G(N446), .D(N462), .Q(neg_mul[22]), .QN(n12) );
  TLATX1 neg_mul_reg_21_ ( .G(N446), .D(N461), .Q(neg_mul[21]), .QN(n11) );
  TLATX1 neg_mul_reg_20_ ( .G(N446), .D(N460), .QN(n16) );
  TLATX1 neg_mul_reg_11_ ( .G(N446), .D(N451), .Q(neg_mul[11]), .QN(n7) );
  TLATX1 neg_mul_reg_14_ ( .G(N446), .D(N454), .Q(neg_mul[14]), .QN(n8) );
  TLATX1 neg_mul_reg_13_ ( .G(N446), .D(N453), .Q(neg_mul[13]), .QN(n10) );
  TLATX1 neg_mul_reg_9_ ( .G(N446), .D(N449), .Q(neg_mul[9]), .QN(n6) );
  TLATX1 neg_mul_reg_17_ ( .G(N446), .D(N457), .Q(neg_mul[17]), .QN(n15) );
  TLATX1 neg_mul_reg_12_ ( .G(N446), .D(N452), .Q(neg_mul[12]), .QN(n13) );
  TLATX1 neg_mul_reg_10_ ( .G(N446), .D(N450), .Q(neg_mul[10]), .QN(n5) );
  TLATX1 neg_mul_reg_8_ ( .G(N446), .D(N448), .Q(neg_mul[8]), .QN(n14) );
  TLATX1 neg_mul_reg_7_ ( .G(N446), .D(N447), .Q(out[0]) );
  OAI21X1 U2 ( .A0(n42), .A1(n60), .B0(n59), .Y(n65) );
  NOR2XL U3 ( .A(n100), .B(n51), .Y(n101) );
  MX2X2 U4 ( .A(neg_mul[21]), .B(N479), .S0(n177), .Y(out[14]) );
  NOR2X2 U5 ( .A(n51), .B(n56), .Y(n57) );
  INVX1 U6 ( .A(n20), .Y(n21) );
  CLKINVX3 U7 ( .A(n285), .Y(in_17bit_b[16]) );
  NOR2X2 U8 ( .A(n50), .B(n70), .Y(n72) );
  AOI2BB2X4 U9 ( .B0(n55), .B1(n42), .A0N(n44), .A1N(neg_mul[8]), .Y(n56) );
  AOI2BB2X4 U10 ( .B0(n61), .B1(n42), .A0N(n44), .A1N(neg_mul[9]), .Y(n62) );
  AOI2BB2X4 U11 ( .B0(n69), .B1(n43), .A0N(n44), .A1N(neg_mul[10]), .Y(n70) );
  AOI2BB2X4 U12 ( .B0(n39), .B1(n43), .A0N(n44), .A1N(neg_mul[11]), .Y(n76) );
  INVX12 U13 ( .A(n45), .Y(n44) );
  OAI21X1 U14 ( .A0(n42), .A1(n82), .B0(n81), .Y(n87) );
  INVX1 U15 ( .A(n168), .Y(n52) );
  NAND2X1 U16 ( .A(n43), .B(n7), .Y(n75) );
  OAI21XL U17 ( .A0(n42), .A1(n98), .B0(n97), .Y(n158) );
  OAI21X1 U18 ( .A0(n42), .A1(n90), .B0(n89), .Y(n95) );
  NOR2X1 U19 ( .A(n23), .B(n173), .Y(n174) );
  INVX1 U20 ( .A(n26), .Y(n22) );
  OAI21X1 U21 ( .A0(n42), .A1(n68), .B0(n67), .Y(n73) );
  INVX1 U22 ( .A(n66), .Y(n63) );
  INVX16 U23 ( .A(n45), .Y(n42) );
  CLKINVX3 U24 ( .A(n176), .Y(n177) );
  CLKBUFX3 U25 ( .A(n19), .Y(n20) );
  NOR2X2 U26 ( .A(n51), .B(n62), .Y(n64) );
  AND4X1 U27 ( .A(in_8bit[1]), .B(n43), .C(n224), .D(n41), .Y(n9) );
  NAND2X2 U28 ( .A(n43), .B(n8), .Y(n97) );
  AOI2BB2X2 U29 ( .B0(n83), .B1(n43), .A0N(n44), .A1N(neg_mul[12]), .Y(n84) );
  OAI21X2 U30 ( .A0(n43), .A1(n54), .B0(n53), .Y(n58) );
  NOR2X2 U31 ( .A(n92), .B(n50), .Y(n94) );
  NAND2X1 U32 ( .A(n43), .B(n10), .Y(n89) );
  OR4XL U33 ( .A(in_8bit[4]), .B(in_8bit[5]), .C(in_8bit[6]), .D(n43), .Y(n228) );
  AOI2BB2X2 U34 ( .B0(n91), .B1(n43), .A0N(n43), .A1N(neg_mul[13]), .Y(n92) );
  CLKBUFX8 U35 ( .A(n50), .Y(n19) );
  INVX8 U36 ( .A(n49), .Y(n50) );
  NAND2X2 U37 ( .A(n43), .B(n5), .Y(n67) );
  BUFX8 U38 ( .A(n286), .Y(out[5]) );
  INVX4 U39 ( .A(in_8bit[7]), .Y(n45) );
  INVXL U40 ( .A(in_8bit[7]), .Y(n46) );
  OAI2BB1X1 U41 ( .A0N(n46), .A1N(n39), .B0(n75), .Y(n79) );
  NAND2X4 U42 ( .A(n43), .B(n14), .Y(n53) );
  XOR2X4 U43 ( .A(n167), .B(neg_mul[16]), .Y(out[9]) );
  XOR2X4 U44 ( .A(n163), .B(neg_mul[15]), .Y(out[8]) );
  NOR2BX4 U45 ( .AN(n22), .B(n160), .Y(n24) );
  XNOR2X4 U46 ( .A(n23), .B(n42), .Y(n160) );
  AOI211X2 U47 ( .A0(n23), .A1(n87), .B0(n86), .C0(n85), .Y(n286) );
  XNOR2X4 U48 ( .A(n19), .B(n42), .Y(n176) );
  AOI22XL U49 ( .A0(N16), .A1(n19), .B0(in_17bit[3]), .B1(n21), .Y(n241) );
  AOI22XL U50 ( .A0(N27), .A1(n19), .B0(in_17bit[14]), .B1(n21), .Y(n274) );
  AOI22XL U51 ( .A0(N22), .A1(n19), .B0(in_17bit[9]), .B1(n21), .Y(n259) );
  AOI22XL U52 ( .A0(N28), .A1(n19), .B0(in_17bit[15]), .B1(n21), .Y(n277) );
  AOI22XL U53 ( .A0(N18), .A1(n19), .B0(in_17bit[5]), .B1(n21), .Y(n247) );
  AOI22XL U54 ( .A0(N24), .A1(n19), .B0(in_17bit[11]), .B1(n21), .Y(n265) );
  AOI22XL U55 ( .A0(N20), .A1(n19), .B0(in_17bit[7]), .B1(n21), .Y(n253) );
  INVX20 U56 ( .A(n45), .Y(n43) );
  NOR2X4 U57 ( .A(n23), .B(n84), .Y(n86) );
  NOR2X2 U58 ( .A(n51), .B(n76), .Y(n78) );
  NOR2X4 U59 ( .A(n27), .B(n160), .Y(n163) );
  NAND2X2 U60 ( .A(n43), .B(n6), .Y(n59) );
  INVX8 U61 ( .A(n49), .Y(n51) );
  AOI22XL U62 ( .A0(N23), .A1(n20), .B0(in_17bit[10]), .B1(n21), .Y(n262) );
  AOI22XL U63 ( .A0(N17), .A1(n20), .B0(in_17bit[4]), .B1(n21), .Y(n244) );
  AOI22XL U64 ( .A0(N25), .A1(n20), .B0(in_17bit[12]), .B1(n21), .Y(n268) );
  AOI22XL U65 ( .A0(N21), .A1(n20), .B0(in_17bit[8]), .B1(n21), .Y(n256) );
  AOI22XL U66 ( .A0(N19), .A1(n20), .B0(in_17bit[6]), .B1(n21), .Y(n250) );
  AOI22XL U67 ( .A0(N26), .A1(n20), .B0(in_17bit[13]), .B1(n21), .Y(n271) );
  AOI211X4 U68 ( .A0(n23), .A1(n175), .B0(n174), .C0(n26), .Y(out[10]) );
  AOI211X4 U69 ( .A0(n50), .A1(n158), .B0(n101), .C0(n27), .Y(out[7]) );
  NOR2X4 U70 ( .A(n28), .B(n164), .Y(n167) );
  XNOR2X4 U71 ( .A(n23), .B(n42), .Y(n164) );
  AOI2BB2X2 U72 ( .B0(n99), .B1(n43), .A0N(n44), .A1N(neg_mul[14]), .Y(n100)
         );
  AOI2BB2X1 U73 ( .B0(n172), .B1(n42), .A0N(n44), .A1N(neg_mul[17]), .Y(n173)
         );
  NAND4BX1 U74 ( .AN(n44), .B(in_8bit[6]), .C(in_8bit[1]), .D(in_8bit[4]), .Y(
        n184) );
  AOI211X4 U75 ( .A0(n50), .A1(n58), .B0(n57), .C0(n38), .Y(out[1]) );
  BUFX20 U76 ( .A(n50), .Y(n23) );
  AOI211X4 U77 ( .A0(n79), .A1(n51), .B0(n78), .C0(n77), .Y(out[4]) );
  AOI211X4 U78 ( .A0(n73), .A1(n50), .B0(n72), .C0(n71), .Y(out[3]) );
  AOI211X4 U79 ( .A0(n95), .A1(n50), .B0(n94), .C0(n93), .Y(out[6]) );
  OR2X4 U80 ( .A(n176), .B(n35), .Y(n25) );
  AOI22XL U81 ( .A0(N355), .A1(n281), .B0(n203), .B1(in_17bit_b[8]), .Y(n258)
         );
  AOI22XL U82 ( .A0(N356), .A1(n281), .B0(n203), .B1(in_17bit_b[9]), .Y(n261)
         );
  AOI22XL U83 ( .A0(N357), .A1(n281), .B0(n203), .B1(in_17bit_b[10]), .Y(n264)
         );
  AOI22XL U84 ( .A0(N358), .A1(n281), .B0(n203), .B1(in_17bit_b[11]), .Y(n267)
         );
  AOI22XL U85 ( .A0(N120), .A1(n278), .B0(N217), .B1(n282), .Y(n269) );
  AOI22XL U86 ( .A0(N359), .A1(n281), .B0(n203), .B1(in_17bit_b[12]), .Y(n270)
         );
  AOI22XL U87 ( .A0(N121), .A1(n278), .B0(N218), .B1(n282), .Y(n272) );
  AOI22XL U88 ( .A0(N360), .A1(n281), .B0(n203), .B1(in_17bit_b[13]), .Y(n273)
         );
  AOI22XL U89 ( .A0(N122), .A1(n278), .B0(N219), .B1(n282), .Y(n275) );
  AOI22XL U90 ( .A0(N361), .A1(n281), .B0(n203), .B1(in_17bit_b[14]), .Y(n276)
         );
  AOI22XL U91 ( .A0(N123), .A1(n278), .B0(N220), .B1(n282), .Y(n279) );
  AOI22XL U92 ( .A0(N362), .A1(n281), .B0(n203), .B1(in_17bit_b[15]), .Y(n280)
         );
  INVX8 U93 ( .A(in_17bit[16]), .Y(n49) );
  INVX1 U94 ( .A(n274), .Y(in_17bit_b[14]) );
  INVX1 U95 ( .A(n271), .Y(in_17bit_b[13]) );
  INVX1 U96 ( .A(n238), .Y(in_17bit_b[2]) );
  INVX1 U97 ( .A(n247), .Y(in_17bit_b[5]) );
  INVX1 U98 ( .A(n250), .Y(in_17bit_b[6]) );
  INVX1 U99 ( .A(n256), .Y(in_17bit_b[8]) );
  INVX1 U100 ( .A(n259), .Y(in_17bit_b[9]) );
  INVX1 U101 ( .A(n262), .Y(in_17bit_b[10]) );
  INVX1 U102 ( .A(n265), .Y(in_17bit_b[11]) );
  INVX1 U103 ( .A(n268), .Y(in_17bit_b[12]) );
  INVX1 U104 ( .A(n253), .Y(in_17bit_b[7]) );
  INVX1 U105 ( .A(n244), .Y(in_17bit_b[4]) );
  INVX1 U106 ( .A(n241), .Y(in_17bit_b[3]) );
  XNOR2X4 U107 ( .A(n24), .B(n3), .Y(out[11]) );
  OAI21XL U108 ( .A0(n42), .A1(n171), .B0(n170), .Y(n175) );
  ADDFX2 U109 ( .A(in_17bit_b[16]), .B(in_17bit_b[12]), .CI(
        add_1_root_r112_carry_16_), .CO(add_1_root_r112_carry_17_), .S(
        add_1_root_r112_SUM_16_) );
  ADDFX2 U110 ( .A(add_1_root_r119_A_19_), .B(in_17bit_b[13]), .CI(
        add_1_root_r119_carry[19]), .CO(add_1_root_r119_carry[20]), .S(
        add_1_root_r119_SUM_19_) );
  ADDFX2 U111 ( .A(in_17bit_b[16]), .B(in_17bit_b[15]), .CI(
        add_3_root_r119_carry_17_), .CO(add_3_root_r119_carry_18_), .S(
        add_1_root_r119_A_17_) );
  ADDFX2 U112 ( .A(in_17bit_b[16]), .B(in_17bit_b[14]), .CI(
        add_2_root_r115_carry_17_), .CO(add_2_root_r115_carry_18_), .S(
        add_2_root_r115_SUM_17_) );
  ADDFX2 U113 ( .A(in_17bit_b[16]), .B(in_17bit_b[14]), .CI(
        add_1_root_r115_carry_20_), .CO(add_1_root_r115_carry_21_), .S(
        add_1_root_r115_SUM_20_) );
  ADDFX2 U114 ( .A(in_17bit_b[16]), .B(in_17bit_b[15]), .CI(
        add_2_root_r119_carry_20_), .CO(add_2_root_r119_carry_21_), .S(
        add_2_root_r119_SUM_20_) );
  ADDFX2 U115 ( .A(in_17bit_b[3]), .B(n202), .CI(add_2_root_r115_carry_4_), 
        .CO(add_2_root_r115_carry_5_), .S(add_2_root_r115_SUM_4_) );
  ADDFX2 U116 ( .A(in_17bit_b[4]), .B(in_17bit_b[2]), .CI(
        add_2_root_r115_carry_5_), .CO(add_2_root_r115_carry_6_), .S(
        add_2_root_r115_SUM_5_) );
  ADDFX2 U117 ( .A(in_17bit_b[5]), .B(n202), .CI(add_1_root_r112_carry_5_), 
        .CO(add_1_root_r112_carry_6_), .S(add_1_root_r112_SUM_5_) );
  ADDFX2 U118 ( .A(in_17bit_b[6]), .B(in_17bit_b[5]), .CI(
        add_3_root_r119_carry_7_), .CO(add_3_root_r119_carry_8_), .S(
        add_1_root_r119_A_7_) );
  ADDFX2 U119 ( .A(in_17bit_b[6]), .B(in_17bit_b[2]), .CI(
        add_1_root_r112_carry_6_), .CO(add_1_root_r112_carry_7_), .S(
        add_1_root_r112_SUM_6_) );
  ADDFX2 U120 ( .A(in_17bit_b[3]), .B(n202), .CI(add_2_root_r115_carry_4_), 
        .CO(add_1_root_r115_carry_8_), .S(add_1_root_r115_SUM_7_) );
  ADDFX2 U121 ( .A(in_17bit_b[7]), .B(in_17bit_b[6]), .CI(
        add_3_root_r119_carry_8_), .CO(add_3_root_r119_carry_9_), .S(
        add_1_root_r119_A_8_) );
  ADDFX2 U122 ( .A(add_1_root_r119_A_7_), .B(n202), .CI(
        add_1_root_r119_carry[7]), .CO(add_1_root_r119_carry[8]), .S(
        add_1_root_r119_SUM_7_) );
  ADDFX2 U123 ( .A(in_17bit_b[2]), .B(n202), .CI(add_3_root_r119_carry_3_), 
        .CO(add_2_root_r119_carry_7_), .S(add_2_root_r119_SUM_6_) );
  ADDFX2 U124 ( .A(in_17bit_b[4]), .B(in_17bit_b[2]), .CI(
        add_1_root_r115_carry_8_), .CO(add_1_root_r115_carry_9_), .S(
        add_1_root_r115_SUM_8_) );
  ADDFX2 U125 ( .A(in_17bit_b[8]), .B(in_17bit_b[7]), .CI(
        add_3_root_r119_carry_9_), .CO(add_3_root_r119_carry_10_), .S(
        add_1_root_r119_A_9_) );
  ADDFX2 U126 ( .A(add_1_root_r119_A_8_), .B(in_17bit_b[2]), .CI(
        add_1_root_r119_carry[8]), .CO(add_1_root_r119_carry[9]), .S(
        add_1_root_r119_SUM_8_) );
  ADDFX2 U127 ( .A(in_17bit_b[3]), .B(in_17bit_b[2]), .CI(
        add_2_root_r119_carry_7_), .CO(add_2_root_r119_carry_8_), .S(
        add_2_root_r119_SUM_7_) );
  ADDFX2 U128 ( .A(in_17bit_b[6]), .B(in_17bit_b[4]), .CI(
        add_2_root_r115_carry_7_), .CO(add_2_root_r115_carry_8_), .S(
        add_2_root_r115_SUM_7_) );
  ADDFX2 U129 ( .A(in_17bit_b[9]), .B(in_17bit_b[8]), .CI(
        add_3_root_r119_carry_10_), .CO(add_3_root_r119_carry_11_), .S(
        add_1_root_r119_A_10_) );
  ADDFX2 U130 ( .A(in_17bit_b[8]), .B(in_17bit_b[4]), .CI(
        add_1_root_r112_carry_8_), .CO(add_1_root_r112_carry_9_), .S(
        add_1_root_r112_SUM_8_) );
  ADDFX2 U131 ( .A(in_17bit_b[7]), .B(in_17bit_b[5]), .CI(
        add_2_root_r115_carry_8_), .CO(add_2_root_r115_carry_9_), .S(
        add_2_root_r115_SUM_8_) );
  ADDFX2 U132 ( .A(in_17bit_b[9]), .B(in_17bit_b[5]), .CI(
        add_1_root_r112_carry_9_), .CO(add_1_root_r112_carry_10_), .S(
        add_1_root_r112_SUM_9_) );
  ADDFX2 U133 ( .A(in_17bit_b[10]), .B(in_17bit_b[9]), .CI(
        add_3_root_r119_carry_11_), .CO(add_3_root_r119_carry_12_), .S(
        add_1_root_r119_A_11_) );
  ADDFX2 U134 ( .A(add_1_root_r119_A_10_), .B(in_17bit_b[4]), .CI(
        add_1_root_r119_carry[10]), .CO(add_1_root_r119_carry[11]), .S(
        add_1_root_r119_SUM_10_) );
  ADDFX2 U135 ( .A(in_17bit_b[5]), .B(in_17bit_b[4]), .CI(
        add_2_root_r119_carry_9_), .CO(add_2_root_r119_carry_10_), .S(
        add_2_root_r119_SUM_9_) );
  ADDFX2 U136 ( .A(in_17bit_b[8]), .B(in_17bit_b[6]), .CI(
        add_2_root_r115_carry_9_), .CO(add_2_root_r115_carry_10_), .S(
        add_2_root_r115_SUM_9_) );
  ADDFX2 U137 ( .A(in_17bit_b[10]), .B(in_17bit_b[6]), .CI(
        add_1_root_r112_carry_10_), .CO(add_1_root_r112_carry_11_), .S(
        add_1_root_r112_SUM_10_) );
  ADDFX2 U138 ( .A(in_17bit_b[7]), .B(in_17bit_b[5]), .CI(
        add_1_root_r115_carry_11_), .CO(add_1_root_r115_carry_12_), .S(
        add_1_root_r115_SUM_11_) );
  ADDFX2 U139 ( .A(in_17bit_b[11]), .B(in_17bit_b[10]), .CI(
        add_3_root_r119_carry_12_), .CO(add_3_root_r119_carry_13_), .S(
        add_1_root_r119_A_12_) );
  ADDFX2 U140 ( .A(add_1_root_r119_A_11_), .B(in_17bit_b[5]), .CI(
        add_1_root_r119_carry[11]), .CO(add_1_root_r119_carry[12]), .S(
        add_1_root_r119_SUM_11_) );
  ADDFX2 U141 ( .A(in_17bit_b[6]), .B(in_17bit_b[5]), .CI(
        add_2_root_r119_carry_10_), .CO(add_2_root_r119_carry_11_), .S(
        add_2_root_r119_SUM_10_) );
  ADDFX2 U142 ( .A(in_17bit_b[9]), .B(in_17bit_b[7]), .CI(
        add_2_root_r115_carry_10_), .CO(add_2_root_r115_carry_11_), .S(
        add_2_root_r115_SUM_10_) );
  ADDFX2 U143 ( .A(in_17bit_b[11]), .B(in_17bit_b[7]), .CI(
        add_1_root_r112_carry_11_), .CO(add_1_root_r112_carry_12_), .S(
        add_1_root_r112_SUM_11_) );
  ADDFX2 U144 ( .A(in_17bit_b[8]), .B(in_17bit_b[6]), .CI(
        add_1_root_r115_carry_12_), .CO(add_1_root_r115_carry_13_), .S(
        add_1_root_r115_SUM_12_) );
  ADDFX2 U145 ( .A(in_17bit_b[12]), .B(in_17bit_b[11]), .CI(
        add_3_root_r119_carry_13_), .CO(add_3_root_r119_carry_14_), .S(
        add_1_root_r119_A_13_) );
  ADDFX2 U146 ( .A(add_1_root_r119_A_12_), .B(in_17bit_b[6]), .CI(
        add_1_root_r119_carry[12]), .CO(add_1_root_r119_carry[13]), .S(
        add_1_root_r119_SUM_12_) );
  ADDFX2 U147 ( .A(in_17bit_b[7]), .B(in_17bit_b[6]), .CI(
        add_2_root_r119_carry_11_), .CO(add_2_root_r119_carry_12_), .S(
        add_2_root_r119_SUM_11_) );
  ADDFX2 U148 ( .A(in_17bit_b[10]), .B(in_17bit_b[8]), .CI(
        add_2_root_r115_carry_11_), .CO(add_2_root_r115_carry_12_), .S(
        add_2_root_r115_SUM_11_) );
  ADDFX2 U149 ( .A(in_17bit_b[12]), .B(in_17bit_b[8]), .CI(
        add_1_root_r112_carry_12_), .CO(add_1_root_r112_carry_13_), .S(
        add_1_root_r112_SUM_12_) );
  ADDFX2 U150 ( .A(in_17bit_b[9]), .B(in_17bit_b[7]), .CI(
        add_1_root_r115_carry_13_), .CO(add_1_root_r115_carry_14_), .S(
        add_1_root_r115_SUM_13_) );
  ADDFX2 U151 ( .A(in_17bit_b[13]), .B(in_17bit_b[12]), .CI(
        add_3_root_r119_carry_14_), .CO(add_3_root_r119_carry_15_), .S(
        add_1_root_r119_A_14_) );
  ADDFX2 U152 ( .A(add_1_root_r119_A_13_), .B(in_17bit_b[7]), .CI(
        add_1_root_r119_carry[13]), .CO(add_1_root_r119_carry[14]), .S(
        add_1_root_r119_SUM_13_) );
  ADDFX2 U153 ( .A(in_17bit_b[8]), .B(in_17bit_b[7]), .CI(
        add_2_root_r119_carry_12_), .CO(add_2_root_r119_carry_13_), .S(
        add_2_root_r119_SUM_12_) );
  ADDFX2 U154 ( .A(in_17bit_b[11]), .B(in_17bit_b[9]), .CI(
        add_2_root_r115_carry_12_), .CO(add_2_root_r115_carry_13_), .S(
        add_2_root_r115_SUM_12_) );
  ADDFX2 U155 ( .A(in_17bit_b[13]), .B(in_17bit_b[9]), .CI(
        add_1_root_r112_carry_13_), .CO(add_1_root_r112_carry_14_), .S(
        add_1_root_r112_SUM_13_) );
  ADDFX2 U156 ( .A(in_17bit_b[10]), .B(in_17bit_b[8]), .CI(
        add_1_root_r115_carry_14_), .CO(add_1_root_r115_carry_15_), .S(
        add_1_root_r115_SUM_14_) );
  ADDFX2 U157 ( .A(in_17bit_b[14]), .B(in_17bit_b[13]), .CI(
        add_3_root_r119_carry_15_), .CO(add_3_root_r119_carry_16_), .S(
        add_1_root_r119_A_15_) );
  ADDFX2 U158 ( .A(add_1_root_r119_A_14_), .B(in_17bit_b[8]), .CI(
        add_1_root_r119_carry[14]), .CO(add_1_root_r119_carry[15]), .S(
        add_1_root_r119_SUM_14_) );
  ADDFX2 U159 ( .A(in_17bit_b[3]), .B(in_17bit_b[2]), .CI(
        add_3_root_r119_carry_4_), .CO(add_3_root_r119_carry_5_), .S(
        add_1_root_r119_A_4_) );
  ADDFX2 U160 ( .A(in_17bit_b[2]), .B(n202), .CI(add_3_root_r119_carry_3_), 
        .CO(add_3_root_r119_carry_4_), .S(add_1_root_r119_A_3_) );
  ADDFX2 U161 ( .A(in_17bit_b[9]), .B(in_17bit_b[8]), .CI(
        add_2_root_r119_carry_13_), .CO(add_2_root_r119_carry_14_), .S(
        add_2_root_r119_SUM_13_) );
  ADDFX2 U162 ( .A(in_17bit_b[12]), .B(in_17bit_b[10]), .CI(
        add_2_root_r115_carry_13_), .CO(add_2_root_r115_carry_14_), .S(
        add_2_root_r115_SUM_13_) );
  ADDFX2 U163 ( .A(in_17bit_b[14]), .B(in_17bit_b[10]), .CI(
        add_1_root_r112_carry_14_), .CO(add_1_root_r112_carry_15_), .S(
        add_1_root_r112_SUM_14_) );
  ADDFX2 U164 ( .A(in_17bit_b[11]), .B(in_17bit_b[9]), .CI(
        add_1_root_r115_carry_15_), .CO(add_1_root_r115_carry_16_), .S(
        add_1_root_r115_SUM_15_) );
  ADDFX2 U165 ( .A(add_1_root_r119_A_15_), .B(in_17bit_b[9]), .CI(
        add_1_root_r119_carry[15]), .CO(add_1_root_r119_carry[16]), .S(
        add_1_root_r119_SUM_15_) );
  ADDFX2 U166 ( .A(in_17bit_b[10]), .B(in_17bit_b[9]), .CI(
        add_2_root_r119_carry_14_), .CO(add_2_root_r119_carry_15_), .S(
        add_2_root_r119_SUM_14_) );
  ADDFX2 U167 ( .A(in_17bit_b[13]), .B(in_17bit_b[11]), .CI(
        add_2_root_r115_carry_14_), .CO(add_2_root_r115_carry_15_), .S(
        add_2_root_r115_SUM_14_) );
  ADDFX2 U168 ( .A(in_17bit_b[15]), .B(in_17bit_b[11]), .CI(
        add_1_root_r112_carry_15_), .CO(add_1_root_r112_carry_16_), .S(
        add_1_root_r112_SUM_15_) );
  ADDFX2 U169 ( .A(in_17bit_b[12]), .B(in_17bit_b[10]), .CI(
        add_1_root_r115_carry_16_), .CO(add_1_root_r115_carry_17_), .S(
        add_1_root_r115_SUM_16_) );
  ADDFX2 U170 ( .A(add_1_root_r119_A_16_), .B(in_17bit_b[10]), .CI(
        add_1_root_r119_carry[16]), .CO(add_1_root_r119_carry[17]), .S(
        add_1_root_r119_SUM_16_) );
  ADDFX2 U171 ( .A(in_17bit_b[11]), .B(in_17bit_b[10]), .CI(
        add_2_root_r119_carry_15_), .CO(add_2_root_r119_carry_16_), .S(
        add_2_root_r119_SUM_15_) );
  ADDFX2 U172 ( .A(in_17bit_b[14]), .B(in_17bit_b[12]), .CI(
        add_2_root_r115_carry_15_), .CO(add_2_root_r115_carry_16_), .S(
        add_2_root_r115_SUM_15_) );
  ADDFX2 U173 ( .A(in_17bit_b[13]), .B(in_17bit_b[11]), .CI(
        add_1_root_r115_carry_17_), .CO(add_1_root_r115_carry_18_), .S(
        add_1_root_r115_SUM_17_) );
  ADDFX2 U174 ( .A(add_1_root_r119_A_17_), .B(in_17bit_b[11]), .CI(
        add_1_root_r119_carry[17]), .CO(add_1_root_r119_carry[18]), .S(
        add_1_root_r119_SUM_17_) );
  ADDFX2 U175 ( .A(in_17bit_b[12]), .B(in_17bit_b[11]), .CI(
        add_2_root_r119_carry_16_), .CO(add_2_root_r119_carry_17_), .S(
        add_2_root_r119_SUM_16_) );
  ADDFX2 U176 ( .A(in_17bit_b[15]), .B(in_17bit_b[13]), .CI(
        add_2_root_r115_carry_16_), .CO(add_2_root_r115_carry_17_), .S(
        add_2_root_r115_SUM_16_) );
  ADDFX2 U177 ( .A(in_17bit_b[14]), .B(in_17bit_b[12]), .CI(
        add_1_root_r115_carry_18_), .CO(add_1_root_r115_carry_19_), .S(
        add_1_root_r115_SUM_18_) );
  ADDFX2 U178 ( .A(add_1_root_r119_A_18_), .B(in_17bit_b[12]), .CI(
        add_1_root_r119_carry[18]), .CO(add_1_root_r119_carry[19]), .S(
        add_1_root_r119_SUM_18_) );
  ADDFX2 U179 ( .A(in_17bit_b[13]), .B(in_17bit_b[12]), .CI(
        add_2_root_r119_carry_17_), .CO(add_2_root_r119_carry_18_), .S(
        add_2_root_r119_SUM_17_) );
  ADDFX2 U180 ( .A(in_17bit_b[15]), .B(in_17bit_b[13]), .CI(
        add_1_root_r115_carry_19_), .CO(add_1_root_r115_carry_20_), .S(
        add_1_root_r115_SUM_19_) );
  ADDFX2 U181 ( .A(in_17bit_b[14]), .B(in_17bit_b[13]), .CI(
        add_2_root_r119_carry_18_), .CO(add_2_root_r119_carry_19_), .S(
        add_2_root_r119_SUM_18_) );
  ADDFX2 U182 ( .A(in_17bit_b[5]), .B(in_17bit_b[3]), .CI(
        add_2_root_r115_carry_6_), .CO(add_2_root_r115_carry_7_), .S(
        add_2_root_r115_SUM_6_) );
  ADDFX2 U183 ( .A(in_17bit_b[7]), .B(in_17bit_b[3]), .CI(
        add_1_root_r112_carry_7_), .CO(add_1_root_r112_carry_8_), .S(
        add_1_root_r112_SUM_7_) );
  ADDFX2 U184 ( .A(in_17bit_b[5]), .B(in_17bit_b[3]), .CI(
        add_1_root_r115_carry_9_), .CO(add_1_root_r115_carry_10_), .S(
        add_1_root_r115_SUM_9_) );
  ADDFX2 U185 ( .A(add_1_root_r119_A_9_), .B(in_17bit_b[3]), .CI(
        add_1_root_r119_carry[9]), .CO(add_1_root_r119_carry[10]), .S(
        add_1_root_r119_SUM_9_) );
  ADDFX2 U186 ( .A(in_17bit_b[4]), .B(in_17bit_b[3]), .CI(
        add_2_root_r119_carry_8_), .CO(add_2_root_r119_carry_9_), .S(
        add_2_root_r119_SUM_8_) );
  ADDFX2 U187 ( .A(in_17bit_b[6]), .B(in_17bit_b[4]), .CI(
        add_1_root_r115_carry_10_), .CO(add_1_root_r115_carry_11_), .S(
        add_1_root_r115_SUM_10_) );
  ADDFX2 U188 ( .A(in_17bit_b[15]), .B(in_17bit_b[14]), .CI(
        add_3_root_r119_carry_16_), .CO(add_3_root_r119_carry_17_), .S(
        add_1_root_r119_A_16_) );
  ADDFX2 U189 ( .A(in_17bit_b[5]), .B(in_17bit_b[4]), .CI(
        add_3_root_r119_carry_6_), .CO(add_3_root_r119_carry_7_), .S(
        add_1_root_r119_A_6_) );
  ADDFX2 U190 ( .A(in_17bit_b[4]), .B(in_17bit_b[3]), .CI(
        add_3_root_r119_carry_5_), .CO(add_3_root_r119_carry_6_), .S(
        add_1_root_r119_A_5_) );
  ADDFX2 U191 ( .A(in_17bit_b[15]), .B(in_17bit_b[14]), .CI(
        add_2_root_r119_carry_19_), .CO(add_2_root_r119_carry_20_), .S(
        add_2_root_r119_SUM_19_) );
  CLKINVX3 U192 ( .A(n232), .Y(in_17bit_b[0]) );
  INVX1 U193 ( .A(n203), .Y(n284) );
  NAND2XL U194 ( .A(N29), .B(n19), .Y(n285) );
  OAI21XL U195 ( .A0(n284), .A1(n285), .B0(n283), .Y(N463) );
  AOI22XL U196 ( .A0(N221), .A1(n282), .B0(N363), .B1(n281), .Y(n283) );
  INVX1 U197 ( .A(n80), .Y(n77) );
  CLKINVX3 U198 ( .A(n277), .Y(in_17bit_b[15]) );
  INVX1 U199 ( .A(n96), .Y(n93) );
  INVX1 U200 ( .A(n88), .Y(n85) );
  INVX1 U201 ( .A(n74), .Y(n71) );
  NAND2X1 U202 ( .A(n30), .B(in_8bit[1]), .Y(n178) );
  INVX1 U203 ( .A(in_8bit[2]), .Y(n47) );
  INVX1 U204 ( .A(in_8bit[0]), .Y(n41) );
  INVX1 U205 ( .A(in_8bit[5]), .Y(n48) );
  XOR2X2 U206 ( .A(n25), .B(n4), .Y(out[12]) );
  NAND2XL U207 ( .A(n43), .B(n13), .Y(n81) );
  NOR3X1 U208 ( .A(n47), .B(n204), .C(n41), .Y(n230) );
  AND2X2 U209 ( .A(n52), .B(n15), .Y(n26) );
  AND2X2 U210 ( .A(n93), .B(n8), .Y(n27) );
  NAND2X1 U211 ( .A(n38), .B(n6), .Y(n66) );
  AND2X2 U212 ( .A(n27), .B(n2), .Y(n28) );
  NOR2X1 U213 ( .A(in_8bit[0]), .B(n184), .Y(n29) );
  AND3X1 U214 ( .A(n43), .B(n179), .C(n48), .Y(n30) );
  AOI21X1 U215 ( .A0(n183), .A1(n9), .B0(n32), .Y(n31) );
  INVX1 U216 ( .A(n31), .Y(n281) );
  AND2X2 U217 ( .A(n29), .B(n36), .Y(n32) );
  AOI21X1 U218 ( .A0(n36), .A1(n9), .B0(n34), .Y(n33) );
  INVX1 U219 ( .A(n33), .Y(n282) );
  AND2X2 U220 ( .A(n29), .B(n183), .Y(n34) );
  NAND2X1 U221 ( .A(n28), .B(n1), .Y(n168) );
  NAND2X1 U222 ( .A(n85), .B(n10), .Y(n96) );
  NAND2X1 U223 ( .A(n71), .B(n7), .Y(n80) );
  OAI2BB1X1 U224 ( .A0N(n229), .A1N(n30), .B0(n185), .Y(n203) );
  NAND3BX1 U225 ( .AN(n184), .B(n230), .C(in_8bit[5]), .Y(n185) );
  NAND2X1 U226 ( .A(n77), .B(n13), .Y(n88) );
  AND2X2 U227 ( .A(n26), .B(n3), .Y(n35) );
  INVX1 U228 ( .A(in_17bit[3]), .Y(n189) );
  INVX1 U229 ( .A(in_17bit[4]), .Y(n190) );
  INVX1 U230 ( .A(in_17bit[5]), .Y(n191) );
  INVX1 U231 ( .A(in_17bit[6]), .Y(n192) );
  INVX1 U232 ( .A(in_17bit[7]), .Y(n193) );
  INVX1 U233 ( .A(in_17bit[8]), .Y(n194) );
  INVX1 U234 ( .A(in_17bit[9]), .Y(n195) );
  INVX1 U235 ( .A(in_17bit[10]), .Y(n196) );
  INVX1 U236 ( .A(in_17bit[11]), .Y(n197) );
  INVX1 U237 ( .A(in_17bit[12]), .Y(n198) );
  INVX1 U238 ( .A(in_17bit[13]), .Y(n199) );
  INVX1 U239 ( .A(in_17bit[14]), .Y(n200) );
  INVX1 U240 ( .A(in_17bit[15]), .Y(n201) );
  NAND2BX1 U241 ( .AN(n66), .B(n5), .Y(n74) );
  INVX1 U242 ( .A(in_17bit[1]), .Y(n187) );
  INVX1 U243 ( .A(in_17bit[2]), .Y(n188) );
  INVX1 U244 ( .A(in_17bit[0]), .Y(n186) );
  AND3X2 U245 ( .A(in_8bit[2]), .B(n204), .C(in_8bit[5]), .Y(n36) );
  INVX1 U246 ( .A(n171), .Y(n172) );
  NAND2X1 U247 ( .A(n234), .B(n233), .Y(N447) );
  AOI22X1 U248 ( .A0(N108), .A1(n278), .B0(N205), .B1(n282), .Y(n233) );
  AOI22X1 U249 ( .A0(N347), .A1(n281), .B0(n203), .B1(in_17bit_b[0]), .Y(n234)
         );
  NAND2X1 U250 ( .A(n237), .B(n236), .Y(N448) );
  AOI22X1 U251 ( .A0(N109), .A1(n278), .B0(N206), .B1(n282), .Y(n236) );
  AOI22X1 U252 ( .A0(N348), .A1(n281), .B0(n203), .B1(n202), .Y(n237) );
  INVX1 U253 ( .A(n235), .Y(n202) );
  NAND2X1 U254 ( .A(n240), .B(n239), .Y(N449) );
  AOI22X1 U255 ( .A0(N110), .A1(n278), .B0(N207), .B1(n282), .Y(n239) );
  AOI22X1 U256 ( .A0(N349), .A1(n281), .B0(n203), .B1(in_17bit_b[2]), .Y(n240)
         );
  NAND2X1 U257 ( .A(n243), .B(n242), .Y(N450) );
  AOI22X1 U258 ( .A0(N111), .A1(n278), .B0(N208), .B1(n282), .Y(n242) );
  AOI22X1 U259 ( .A0(N350), .A1(n281), .B0(n203), .B1(in_17bit_b[3]), .Y(n243)
         );
  NAND2X1 U260 ( .A(n246), .B(n245), .Y(N451) );
  AOI22X1 U261 ( .A0(N112), .A1(n278), .B0(N209), .B1(n282), .Y(n245) );
  AOI22X1 U262 ( .A0(N351), .A1(n281), .B0(n203), .B1(in_17bit_b[4]), .Y(n246)
         );
  NAND2X1 U263 ( .A(n249), .B(n248), .Y(N452) );
  AOI22X1 U264 ( .A0(N113), .A1(n278), .B0(N210), .B1(n282), .Y(n248) );
  AOI22X1 U265 ( .A0(N352), .A1(n281), .B0(n203), .B1(in_17bit_b[5]), .Y(n249)
         );
  NAND2X1 U266 ( .A(n252), .B(n251), .Y(N453) );
  AOI22X1 U267 ( .A0(N114), .A1(n278), .B0(N211), .B1(n282), .Y(n251) );
  AOI22X1 U268 ( .A0(N353), .A1(n281), .B0(n203), .B1(in_17bit_b[6]), .Y(n252)
         );
  NAND2X1 U269 ( .A(n255), .B(n254), .Y(N454) );
  AOI22X1 U270 ( .A0(N115), .A1(n278), .B0(N212), .B1(n282), .Y(n254) );
  AOI22X1 U271 ( .A0(N354), .A1(n281), .B0(n203), .B1(in_17bit_b[7]), .Y(n255)
         );
  NAND2X1 U272 ( .A(n258), .B(n257), .Y(N455) );
  AOI22X1 U273 ( .A0(N116), .A1(n278), .B0(N213), .B1(n282), .Y(n257) );
  NAND2X1 U274 ( .A(n261), .B(n260), .Y(N456) );
  AOI22X1 U275 ( .A0(N117), .A1(n278), .B0(N214), .B1(n282), .Y(n260) );
  NAND2X1 U276 ( .A(n264), .B(n263), .Y(N457) );
  AOI22X1 U277 ( .A0(N118), .A1(n278), .B0(N215), .B1(n282), .Y(n263) );
  NAND2X1 U278 ( .A(n267), .B(n266), .Y(N458) );
  AOI22X1 U279 ( .A0(N119), .A1(n278), .B0(N216), .B1(n282), .Y(n266) );
  NAND2X1 U280 ( .A(n270), .B(n269), .Y(N459) );
  NAND2X1 U281 ( .A(n273), .B(n272), .Y(N460) );
  NAND2X1 U282 ( .A(n276), .B(n275), .Y(N461) );
  NAND2X1 U283 ( .A(n280), .B(n279), .Y(N462) );
  INVX1 U284 ( .A(n98), .Y(n99) );
  XNOR2X1 U285 ( .A(n16), .B(sub_add_75_b0_carry[13]), .Y(n37) );
  INVX1 U286 ( .A(n90), .Y(n91) );
  INVX1 U287 ( .A(n68), .Y(n69) );
  INVX1 U288 ( .A(n54), .Y(n55) );
  INVX1 U289 ( .A(n60), .Y(n61) );
  INVX1 U290 ( .A(n82), .Y(n83) );
  MX2X1 U291 ( .A(neg_mul[22]), .B(N480), .S0(n177), .Y(out[15]) );
  MX2X1 U292 ( .A(neg_mul[23]), .B(N481), .S0(n177), .Y(out[16]) );
  NAND4BBX1 U293 ( .AN(n281), .BN(n282), .C(n231), .D(n284), .Y(N446) );
  AOI2BB1X1 U294 ( .A0N(n228), .A1N(n227), .B0(n278), .Y(n231) );
  OR4X2 U295 ( .A(in_8bit[1]), .B(in_8bit[0]), .C(in_8bit[2]), .D(in_8bit[3]), 
        .Y(n227) );
  NOR4BX1 U296 ( .AN(n226), .B(n41), .C(in_8bit[1]), .D(in_8bit[2]), .Y(n229)
         );
  NOR2X1 U297 ( .A(in_8bit[6]), .B(in_8bit[3]), .Y(n226) );
  NOR2X1 U298 ( .A(out[0]), .B(neg_mul[8]), .Y(n38) );
  AND2X2 U299 ( .A(neg_mul[11]), .B(n74), .Y(n39) );
  NAND2BX1 U300 ( .AN(n38), .B(neg_mul[9]), .Y(n60) );
  NAND2X1 U301 ( .A(out[0]), .B(neg_mul[8]), .Y(n54) );
  NAND2X1 U302 ( .A(neg_mul[10]), .B(n66), .Y(n68) );
  NAND2X1 U303 ( .A(n182), .B(n181), .Y(n278) );
  NAND3BX1 U304 ( .AN(n178), .B(n230), .C(in_8bit[6]), .Y(n182) );
  NAND3X1 U305 ( .A(n229), .B(in_8bit[5]), .C(n180), .Y(n181) );
  NAND2X1 U306 ( .A(neg_mul[13]), .B(n88), .Y(n90) );
  NAND2X1 U307 ( .A(neg_mul[14]), .B(n96), .Y(n98) );
  NAND2X1 U308 ( .A(neg_mul[12]), .B(n80), .Y(n82) );
  NOR2X1 U309 ( .A(in_8bit[6]), .B(in_8bit[4]), .Y(n224) );
  NAND2X1 U310 ( .A(neg_mul[17]), .B(n168), .Y(n171) );
  INVX1 U311 ( .A(n225), .Y(n183) );
  NAND3BX1 U312 ( .AN(in_8bit[5]), .B(n47), .C(in_8bit[3]), .Y(n225) );
  INVX1 U313 ( .A(in_8bit[3]), .Y(n204) );
  INVX1 U314 ( .A(in_8bit[4]), .Y(n179) );
  NOR2XL U315 ( .A(n43), .B(n179), .Y(n180) );
  NAND2XL U316 ( .A(n43), .B(n15), .Y(n170) );
  AOI22XL U317 ( .A0(N15), .A1(n20), .B0(in_17bit[2]), .B1(n21), .Y(n238) );
  AOI22XL U318 ( .A0(N14), .A1(n19), .B0(in_17bit[1]), .B1(n21), .Y(n235) );
  AOI22XL U319 ( .A0(in_17bit[0]), .A1(n20), .B0(in_17bit[0]), .B1(n21), .Y(
        n232) );
  AOI211X4 U320 ( .A0(n65), .A1(n51), .B0(n64), .C0(n63), .Y(out[2]) );
  MXI2X4 U321 ( .A(n16), .B(n37), .S0(n177), .Y(out[13]) );
  AND2X1 U322 ( .A(add_1_root_r112_carry_20_), .B(in_17bit_b[16]), .Y(
        add_1_root_r112_SUM_21_) );
  XOR2X1 U323 ( .A(in_17bit_b[16]), .B(add_1_root_r112_carry_20_), .Y(
        add_1_root_r112_SUM_20_) );
  AND2X1 U324 ( .A(add_1_root_r112_carry_19_), .B(in_17bit_b[15]), .Y(
        add_1_root_r112_carry_20_) );
  XOR2X1 U325 ( .A(in_17bit_b[15]), .B(add_1_root_r112_carry_19_), .Y(
        add_1_root_r112_SUM_19_) );
  AND2X1 U326 ( .A(add_1_root_r112_carry_18_), .B(in_17bit_b[14]), .Y(
        add_1_root_r112_carry_19_) );
  XOR2X1 U327 ( .A(in_17bit_b[14]), .B(add_1_root_r112_carry_18_), .Y(
        add_1_root_r112_SUM_18_) );
  AND2X1 U328 ( .A(add_1_root_r112_carry_17_), .B(in_17bit_b[13]), .Y(
        add_1_root_r112_carry_18_) );
  XOR2X1 U329 ( .A(in_17bit_b[13]), .B(add_1_root_r112_carry_17_), .Y(
        add_1_root_r112_SUM_17_) );
  AND2X1 U330 ( .A(add_2_root_r119_carry_21_), .B(in_17bit_b[16]), .Y(
        add_2_root_r119_SUM_22_) );
  XOR2X1 U331 ( .A(in_17bit_b[16]), .B(add_2_root_r119_carry_21_), .Y(
        add_2_root_r119_SUM_21_) );
  XOR2X1 U332 ( .A(in_17bit_b[0]), .B(n202), .Y(add_2_root_r119_SUM_5_) );
  AND2X1 U333 ( .A(add_1_root_r119_carry[22]), .B(in_17bit_b[16]), .Y(
        add_1_root_r119_SUM_23_) );
  XOR2X1 U334 ( .A(in_17bit_b[16]), .B(add_1_root_r119_carry[22]), .Y(
        add_1_root_r119_SUM_22_) );
  AND2X1 U335 ( .A(add_1_root_r119_carry[21]), .B(in_17bit_b[15]), .Y(
        add_1_root_r119_carry[22]) );
  XOR2X1 U336 ( .A(in_17bit_b[15]), .B(add_1_root_r119_carry[21]), .Y(
        add_1_root_r119_SUM_21_) );
  AND2X1 U337 ( .A(add_1_root_r119_carry[20]), .B(in_17bit_b[14]), .Y(
        add_1_root_r119_carry[21]) );
  XOR2X1 U338 ( .A(in_17bit_b[14]), .B(add_1_root_r119_carry[20]), .Y(
        add_1_root_r119_SUM_20_) );
  AND2X1 U339 ( .A(add_1_root_r119_A_6_), .B(in_17bit_b[0]), .Y(
        add_1_root_r119_carry[7]) );
  XOR2X1 U340 ( .A(in_17bit_b[0]), .B(add_1_root_r119_A_6_), .Y(
        add_1_root_r119_SUM_6_) );
  AND2X1 U341 ( .A(add_3_root_r119_carry_18_), .B(in_17bit_b[16]), .Y(
        add_1_root_r119_A_19_) );
  XOR2X1 U342 ( .A(in_17bit_b[16]), .B(add_3_root_r119_carry_18_), .Y(
        add_1_root_r119_A_18_) );
  AND2X1 U343 ( .A(n202), .B(in_17bit_b[0]), .Y(add_3_root_r119_carry_3_) );
  AND2X1 U344 ( .A(add_2_root_r115_carry_19_), .B(in_17bit_b[16]), .Y(
        add_2_root_r115_SUM_20_) );
  XOR2X1 U345 ( .A(in_17bit_b[16]), .B(add_2_root_r115_carry_19_), .Y(
        add_2_root_r115_SUM_19_) );
  AND2X1 U346 ( .A(add_2_root_r115_carry_18_), .B(in_17bit_b[15]), .Y(
        add_2_root_r115_carry_19_) );
  XOR2X1 U347 ( .A(in_17bit_b[15]), .B(add_2_root_r115_carry_18_), .Y(
        add_2_root_r115_SUM_18_) );
  AND2X1 U348 ( .A(in_17bit_b[2]), .B(in_17bit_b[0]), .Y(
        add_2_root_r115_carry_4_) );
  XOR2X1 U349 ( .A(in_17bit_b[0]), .B(in_17bit_b[2]), .Y(
        add_2_root_r115_SUM_3_) );
  AND2X1 U350 ( .A(add_1_root_r115_carry_22_), .B(in_17bit_b[16]), .Y(
        add_1_root_r115_SUM_23_) );
  XOR2X1 U351 ( .A(in_17bit_b[16]), .B(add_1_root_r115_carry_22_), .Y(
        add_1_root_r115_SUM_22_) );
  AND2X1 U352 ( .A(add_1_root_r115_carry_21_), .B(in_17bit_b[15]), .Y(
        add_1_root_r115_carry_22_) );
  XOR2X1 U353 ( .A(in_17bit_b[15]), .B(add_1_root_r115_carry_21_), .Y(
        add_1_root_r115_SUM_21_) );
  XOR2X1 U354 ( .A(n21), .B(sub_add_54_b0_carry[16]), .Y(N29) );
  AND2X1 U355 ( .A(sub_add_54_b0_carry[15]), .B(n201), .Y(
        sub_add_54_b0_carry[16]) );
  XOR2X1 U356 ( .A(n201), .B(sub_add_54_b0_carry[15]), .Y(N28) );
  AND2X1 U357 ( .A(sub_add_54_b0_carry[14]), .B(n200), .Y(
        sub_add_54_b0_carry[15]) );
  XOR2X1 U358 ( .A(n200), .B(sub_add_54_b0_carry[14]), .Y(N27) );
  AND2X1 U359 ( .A(sub_add_54_b0_carry[13]), .B(n199), .Y(
        sub_add_54_b0_carry[14]) );
  XOR2X1 U360 ( .A(n199), .B(sub_add_54_b0_carry[13]), .Y(N26) );
  AND2X1 U361 ( .A(sub_add_54_b0_carry[12]), .B(n198), .Y(
        sub_add_54_b0_carry[13]) );
  XOR2X1 U362 ( .A(n198), .B(sub_add_54_b0_carry[12]), .Y(N25) );
  AND2X1 U363 ( .A(sub_add_54_b0_carry[11]), .B(n197), .Y(
        sub_add_54_b0_carry[12]) );
  XOR2X1 U364 ( .A(n197), .B(sub_add_54_b0_carry[11]), .Y(N24) );
  AND2X1 U365 ( .A(sub_add_54_b0_carry[10]), .B(n196), .Y(
        sub_add_54_b0_carry[11]) );
  XOR2X1 U366 ( .A(n196), .B(sub_add_54_b0_carry[10]), .Y(N23) );
  AND2X1 U367 ( .A(sub_add_54_b0_carry[9]), .B(n195), .Y(
        sub_add_54_b0_carry[10]) );
  XOR2X1 U368 ( .A(n195), .B(sub_add_54_b0_carry[9]), .Y(N22) );
  AND2X1 U369 ( .A(sub_add_54_b0_carry[8]), .B(n194), .Y(
        sub_add_54_b0_carry[9]) );
  XOR2X1 U370 ( .A(n194), .B(sub_add_54_b0_carry[8]), .Y(N21) );
  AND2X1 U371 ( .A(sub_add_54_b0_carry[7]), .B(n193), .Y(
        sub_add_54_b0_carry[8]) );
  XOR2X1 U372 ( .A(n193), .B(sub_add_54_b0_carry[7]), .Y(N20) );
  AND2X1 U373 ( .A(sub_add_54_b0_carry[6]), .B(n192), .Y(
        sub_add_54_b0_carry[7]) );
  XOR2X1 U374 ( .A(n192), .B(sub_add_54_b0_carry[6]), .Y(N19) );
  AND2X1 U375 ( .A(sub_add_54_b0_carry[5]), .B(n191), .Y(
        sub_add_54_b0_carry[6]) );
  XOR2X1 U376 ( .A(n191), .B(sub_add_54_b0_carry[5]), .Y(N18) );
  AND2X1 U377 ( .A(sub_add_54_b0_carry[4]), .B(n190), .Y(
        sub_add_54_b0_carry[5]) );
  XOR2X1 U378 ( .A(n190), .B(sub_add_54_b0_carry[4]), .Y(N17) );
  AND2X1 U379 ( .A(sub_add_54_b0_carry[3]), .B(n189), .Y(
        sub_add_54_b0_carry[4]) );
  XOR2X1 U380 ( .A(n189), .B(sub_add_54_b0_carry[3]), .Y(N16) );
  AND2X1 U381 ( .A(sub_add_54_b0_carry[2]), .B(n188), .Y(
        sub_add_54_b0_carry[3]) );
  XOR2X1 U382 ( .A(n188), .B(sub_add_54_b0_carry[2]), .Y(N15) );
  AND2X1 U383 ( .A(n186), .B(n187), .Y(sub_add_54_b0_carry[2]) );
  XOR2X1 U384 ( .A(n187), .B(n186), .Y(N14) );
  XOR2X1 U385 ( .A(n17), .B(sub_add_75_b0_carry[16]), .Y(N481) );
  AND2X1 U386 ( .A(sub_add_75_b0_carry[15]), .B(n12), .Y(
        sub_add_75_b0_carry[16]) );
  XOR2X1 U387 ( .A(n12), .B(sub_add_75_b0_carry[15]), .Y(N480) );
  AND2X1 U388 ( .A(sub_add_75_b0_carry[14]), .B(n11), .Y(
        sub_add_75_b0_carry[15]) );
  XOR2X1 U389 ( .A(n11), .B(sub_add_75_b0_carry[14]), .Y(N479) );
  AND2X1 U390 ( .A(sub_add_75_b0_carry[13]), .B(n16), .Y(
        sub_add_75_b0_carry[14]) );
  AND2X1 U391 ( .A(n35), .B(n4), .Y(sub_add_75_b0_carry[13]) );
  AND2X1 U392 ( .A(in_17bit_b[0]), .B(in_17bit_b[4]), .Y(
        add_1_root_r112_carry_5_) );
endmodule


module multi16_5_DW01_add_0 ( A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, 
        A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, 
        A_4_, B_23_, B_22_, B_21_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, 
        B_14_, B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, 
        SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, 
        SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, 
        SUM_7_ );
  input A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_,
         A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, B_23_, B_22_,
         B_21_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_,
         B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_;
  output SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_,
         SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_,
         SUM_8_, SUM_7_;
  wire   n1, n2, n3, n4;
  wire   [23:7] carry;

  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry[7]), .CO(carry[8]), .S(SUM_7_)
         );
  ADDFX2 U1_21 ( .A(A_21_), .B(B_21_), .CI(carry[21]), .CO(carry[22]), .S(
        SUM_21_) );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry[20]), .CO(carry[21]), .S(
        SUM_20_) );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry[19]), .CO(carry[20]), .S(
        SUM_19_) );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry[18]), .CO(carry[19]), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry[17]), .CO(carry[18]), .S(
        SUM_17_) );
  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry[16]), .CO(carry[17]), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry[15]), .CO(carry[16]), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry[14]), .CO(carry[15]), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry[13]), .CO(carry[14]), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry[12]), .CO(carry[13]), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry[11]), .CO(carry[12]), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry[10]), .CO(carry[11]), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry[9]), .CO(carry[10]), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry[8]), .CO(carry[9]), .S(SUM_8_)
         );
  ADDFX2 U1_22 ( .A(A_22_), .B(B_22_), .CI(carry[22]), .CO(carry[23]), .S(
        SUM_22_) );
  AND2X2 U1 ( .A(A_4_), .B(B_4_), .Y(n1) );
  XOR2X1 U2 ( .A(B_23_), .B(carry[23]), .Y(SUM_23_) );
  OAI2BB1X1 U3 ( .A0N(n2), .A1N(A_6_), .B0(n3), .Y(carry[7]) );
  OAI21XL U4 ( .A0(A_6_), .A1(n2), .B0(B_6_), .Y(n3) );
  OAI2BB1X1 U5 ( .A0N(n1), .A1N(A_5_), .B0(n4), .Y(n2) );
  OAI21XL U6 ( .A0(A_5_), .A1(n1), .B0(B_5_), .Y(n4) );
endmodule


module multi16_5_DW01_add_4 ( A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, 
        A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, 
        B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, 
        B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, SUM_22_, SUM_21_, SUM_20_, 
        SUM_19_, SUM_18_, SUM_17_, SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, 
        SUM_11_, SUM_10_, SUM_9_, SUM_8_, SUM_7_ );
  input A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_,
         A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, B_20_, B_19_,
         B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, B_10_, B_9_,
         B_8_, B_7_, B_6_, B_5_;
  output SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_,
         SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_,
         SUM_7_;
  wire   carry_21_, carry_20_, carry_19_, carry_18_, carry_17_, carry_16_,
         carry_15_, carry_14_, carry_13_, carry_12_, carry_11_, carry_10_,
         carry_9_, carry_8_, carry_7_, n1;

  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry_16_), .CO(carry_17_), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry_15_), .CO(carry_16_), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry_14_), .CO(carry_15_), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry_13_), .CO(carry_14_), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry_12_), .CO(carry_13_), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry_11_), .CO(carry_12_), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry_10_), .CO(carry_11_), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry_9_), .CO(carry_10_), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry_8_), .CO(carry_9_), .S(SUM_8_)
         );
  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry_7_), .CO(carry_8_), .S(SUM_7_)
         );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry_20_), .CO(carry_21_), .S(
        SUM_20_) );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry_19_), .CO(carry_20_), .S(
        SUM_19_) );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry_18_), .CO(carry_19_), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry_17_), .CO(carry_18_), .S(
        SUM_17_) );
  ADDFX2 U1_21 ( .A(A_21_), .B(B_21_), .CI(carry_21_), .CO(SUM_22_), .S(
        SUM_21_) );
  OAI2BB1X1 U1 ( .A0N(A_6_), .A1N(B_6_), .B0(n1), .Y(carry_7_) );
  OAI211X1 U2 ( .A0(B_6_), .A1(A_6_), .B0(A_5_), .C0(B_5_), .Y(n1) );
endmodule


module multi16_5_DW01_add_6 ( A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, 
        A_16_, A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, 
        A_6_, A_5_, A_4_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, 
        B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, 
        SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, 
        SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, 
        SUM_7_ );
  input A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_,
         A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, B_20_,
         B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, B_10_,
         B_9_, B_8_, B_7_, B_6_, B_5_, B_4_;
  output SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_,
         SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_,
         SUM_8_, SUM_7_;
  wire   n1, n2, n3, n4, n5, n6;
  wire   [21:7] carry;

  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry[7]), .CO(carry[8]), .S(SUM_7_)
         );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry[18]), .CO(carry[19]), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry[17]), .CO(carry[18]), .S(
        SUM_17_) );
  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry[16]), .CO(carry[17]), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry[15]), .CO(carry[16]), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry[14]), .CO(carry[15]), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry[13]), .CO(carry[14]), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry[12]), .CO(carry[13]), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry[11]), .CO(carry[12]), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry[10]), .CO(carry[11]), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry[9]), .CO(carry[10]), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry[8]), .CO(carry[9]), .S(SUM_8_)
         );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry[19]), .CO(carry[20]), .S(
        SUM_19_) );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry[20]), .CO(carry[21]), .S(
        SUM_20_) );
  AND2X2 U1 ( .A(A_22_), .B(n2), .Y(n1) );
  AND2X2 U2 ( .A(A_21_), .B(carry[21]), .Y(n2) );
  XOR2X1 U3 ( .A(A_23_), .B(n1), .Y(SUM_23_) );
  AND2X2 U4 ( .A(A_4_), .B(B_4_), .Y(n3) );
  XOR2X1 U5 ( .A(A_21_), .B(carry[21]), .Y(SUM_21_) );
  XOR2X1 U6 ( .A(A_22_), .B(n2), .Y(SUM_22_) );
  OAI2BB1X1 U7 ( .A0N(n4), .A1N(A_6_), .B0(n5), .Y(carry[7]) );
  OAI21XL U8 ( .A0(A_6_), .A1(n4), .B0(B_6_), .Y(n5) );
  OAI2BB1X1 U9 ( .A0N(n3), .A1N(A_5_), .B0(n6), .Y(n4) );
  OAI21XL U10 ( .A0(A_5_), .A1(n3), .B0(B_5_), .Y(n6) );
endmodule


module multi16_5 ( in_17bit, in_8bit, out );
  input [16:0] in_17bit;
  input [7:0] in_8bit;
  output [16:0] out;
  wire   N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27,
         N28, N29, N108, N109, N110, N111, N112, N113, N114, N115, N116, N117,
         N118, N119, N120, N121, N122, N123, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220,
         N221, N347, N348, N349, N350, N351, N352, N353, N354, N355, N356,
         N357, N358, N359, N360, N361, N362, N363, N446, N447, N448, N449,
         N450, N451, N452, N453, N454, N455, N456, N457, N458, N459, N460,
         N461, N462, N463, N478, N479, N480, add_2_root_r119_carry_10_,
         add_2_root_r119_carry_11_, add_2_root_r119_carry_12_,
         add_2_root_r119_carry_13_, add_2_root_r119_carry_14_,
         add_2_root_r119_carry_15_, add_2_root_r119_carry_16_,
         add_2_root_r119_carry_17_, add_2_root_r119_carry_18_,
         add_2_root_r119_carry_19_, add_2_root_r119_carry_20_,
         add_2_root_r119_carry_21_, add_2_root_r119_carry_6_,
         add_2_root_r119_carry_7_, add_2_root_r119_carry_8_,
         add_2_root_r119_carry_9_, add_2_root_r119_SUM_6_,
         add_2_root_r119_SUM_7_, add_2_root_r119_SUM_8_,
         add_2_root_r119_SUM_9_, add_2_root_r119_SUM_10_,
         add_2_root_r119_SUM_11_, add_2_root_r119_SUM_12_,
         add_2_root_r119_SUM_13_, add_2_root_r119_SUM_14_,
         add_2_root_r119_SUM_15_, add_2_root_r119_SUM_16_,
         add_2_root_r119_SUM_17_, add_2_root_r119_SUM_18_,
         add_2_root_r119_SUM_19_, add_2_root_r119_SUM_20_,
         add_2_root_r119_SUM_21_, add_2_root_r119_SUM_22_,
         add_1_root_r119_SUM_6_, add_1_root_r119_SUM_7_,
         add_1_root_r119_SUM_8_, add_1_root_r119_SUM_9_,
         add_1_root_r119_SUM_10_, add_1_root_r119_SUM_11_,
         add_1_root_r119_SUM_12_, add_1_root_r119_SUM_13_,
         add_1_root_r119_SUM_14_, add_1_root_r119_SUM_15_,
         add_1_root_r119_SUM_16_, add_1_root_r119_SUM_17_,
         add_1_root_r119_SUM_18_, add_1_root_r119_SUM_19_,
         add_1_root_r119_SUM_20_, add_1_root_r119_SUM_21_,
         add_1_root_r119_SUM_22_, add_1_root_r119_SUM_23_,
         add_1_root_r119_A_2_, add_1_root_r119_A_3_, add_1_root_r119_A_4_,
         add_1_root_r119_A_5_, add_1_root_r119_A_6_, add_1_root_r119_A_7_,
         add_1_root_r119_A_8_, add_1_root_r119_A_9_, add_1_root_r119_A_10_,
         add_1_root_r119_A_11_, add_1_root_r119_A_12_, add_1_root_r119_A_13_,
         add_1_root_r119_A_14_, add_1_root_r119_A_15_, add_1_root_r119_A_16_,
         add_1_root_r119_A_17_, add_1_root_r119_A_18_, add_1_root_r119_A_19_,
         add_3_root_r119_carry_10_, add_3_root_r119_carry_11_,
         add_3_root_r119_carry_12_, add_3_root_r119_carry_13_,
         add_3_root_r119_carry_14_, add_3_root_r119_carry_15_,
         add_3_root_r119_carry_16_, add_3_root_r119_carry_17_,
         add_3_root_r119_carry_18_, add_3_root_r119_carry_4_,
         add_3_root_r119_carry_5_, add_3_root_r119_carry_6_,
         add_3_root_r119_carry_7_, add_3_root_r119_carry_8_,
         add_3_root_r119_carry_9_, add_1_root_r112_carry_10_,
         add_1_root_r112_carry_11_, add_1_root_r112_carry_12_,
         add_1_root_r112_carry_13_, add_1_root_r112_carry_14_,
         add_1_root_r112_carry_15_, add_1_root_r112_carry_16_,
         add_1_root_r112_carry_17_, add_1_root_r112_carry_18_,
         add_1_root_r112_carry_19_, add_1_root_r112_carry_20_,
         add_1_root_r112_carry_5_, add_1_root_r112_carry_6_,
         add_1_root_r112_carry_7_, add_1_root_r112_carry_8_,
         add_1_root_r112_carry_9_, add_1_root_r112_SUM_1_,
         add_1_root_r112_SUM_2_, add_1_root_r112_SUM_3_,
         add_1_root_r112_SUM_4_, add_1_root_r112_SUM_5_,
         add_1_root_r112_SUM_6_, add_1_root_r112_SUM_7_,
         add_1_root_r112_SUM_8_, add_1_root_r112_SUM_9_,
         add_1_root_r112_SUM_10_, add_1_root_r112_SUM_11_,
         add_1_root_r112_SUM_12_, add_1_root_r112_SUM_13_,
         add_1_root_r112_SUM_14_, add_1_root_r112_SUM_15_,
         add_1_root_r112_SUM_16_, add_1_root_r112_SUM_17_,
         add_1_root_r112_SUM_18_, add_1_root_r112_SUM_19_,
         add_1_root_r112_SUM_20_, add_1_root_r112_SUM_21_,
         add_2_root_r115_carry_10_, add_2_root_r115_carry_11_,
         add_2_root_r115_carry_12_, add_2_root_r115_carry_13_,
         add_2_root_r115_carry_14_, add_2_root_r115_carry_15_,
         add_2_root_r115_carry_16_, add_2_root_r115_carry_17_,
         add_2_root_r115_carry_18_, add_2_root_r115_carry_19_,
         add_2_root_r115_carry_4_, add_2_root_r115_carry_5_,
         add_2_root_r115_carry_6_, add_2_root_r115_carry_7_,
         add_2_root_r115_carry_8_, add_2_root_r115_carry_9_,
         add_2_root_r115_SUM_4_, add_2_root_r115_SUM_5_,
         add_2_root_r115_SUM_6_, add_2_root_r115_SUM_7_,
         add_2_root_r115_SUM_8_, add_2_root_r115_SUM_9_,
         add_2_root_r115_SUM_10_, add_2_root_r115_SUM_11_,
         add_2_root_r115_SUM_12_, add_2_root_r115_SUM_13_,
         add_2_root_r115_SUM_14_, add_2_root_r115_SUM_15_,
         add_2_root_r115_SUM_16_, add_2_root_r115_SUM_17_,
         add_2_root_r115_SUM_18_, add_2_root_r115_SUM_19_,
         add_2_root_r115_SUM_20_, add_1_root_r115_carry_10_,
         add_1_root_r115_carry_11_, add_1_root_r115_carry_12_,
         add_1_root_r115_carry_13_, add_1_root_r115_carry_14_,
         add_1_root_r115_carry_15_, add_1_root_r115_carry_16_,
         add_1_root_r115_carry_17_, add_1_root_r115_carry_18_,
         add_1_root_r115_carry_19_, add_1_root_r115_carry_20_,
         add_1_root_r115_carry_21_, add_1_root_r115_carry_22_,
         add_1_root_r115_carry_8_, add_1_root_r115_carry_9_,
         add_1_root_r115_SUM_6_, add_1_root_r115_SUM_7_,
         add_1_root_r115_SUM_8_, add_1_root_r115_SUM_9_,
         add_1_root_r115_SUM_10_, add_1_root_r115_SUM_11_,
         add_1_root_r115_SUM_12_, add_1_root_r115_SUM_13_,
         add_1_root_r115_SUM_14_, add_1_root_r115_SUM_15_,
         add_1_root_r115_SUM_16_, add_1_root_r115_SUM_17_,
         add_1_root_r115_SUM_18_, add_1_root_r115_SUM_19_,
         add_1_root_r115_SUM_20_, add_1_root_r115_SUM_21_,
         add_1_root_r115_SUM_22_, add_1_root_r115_SUM_23_, n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n158, n160, n161, n162,
         n163, n164, n170, n171, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252;
  wire   [16:0] in_17bit_b;
  wire   [23:8] neg_mul;
  wire   [15:12] sub_add_75_b0_carry;
  wire   [16:2] sub_add_54_b0_carry;
  wire   [22:7] add_1_root_r119_carry;

  multi16_5_DW01_add_0 add_0_root_r119 ( .A_22_(add_2_root_r119_SUM_22_), 
        .A_21_(add_2_root_r119_SUM_21_), .A_20_(add_2_root_r119_SUM_20_), 
        .A_19_(add_2_root_r119_SUM_19_), .A_18_(add_2_root_r119_SUM_18_), 
        .A_17_(add_2_root_r119_SUM_17_), .A_16_(add_2_root_r119_SUM_16_), 
        .A_15_(add_2_root_r119_SUM_15_), .A_14_(add_2_root_r119_SUM_14_), 
        .A_13_(add_2_root_r119_SUM_13_), .A_12_(add_2_root_r119_SUM_12_), 
        .A_11_(add_2_root_r119_SUM_11_), .A_10_(add_2_root_r119_SUM_10_), 
        .A_9_(add_2_root_r119_SUM_9_), .A_8_(add_2_root_r119_SUM_8_), .A_7_(
        add_2_root_r119_SUM_7_), .A_6_(add_2_root_r119_SUM_6_), .A_5_(
        add_1_root_r119_A_2_), .A_4_(in_17bit_b[0]), .B_23_(
        add_1_root_r119_SUM_23_), .B_22_(add_1_root_r119_SUM_22_), .B_21_(
        add_1_root_r119_SUM_21_), .B_20_(add_1_root_r119_SUM_20_), .B_19_(
        add_1_root_r119_SUM_19_), .B_18_(add_1_root_r119_SUM_18_), .B_17_(
        add_1_root_r119_SUM_17_), .B_16_(add_1_root_r119_SUM_16_), .B_15_(
        add_1_root_r119_SUM_15_), .B_14_(add_1_root_r119_SUM_14_), .B_13_(
        add_1_root_r119_SUM_13_), .B_12_(add_1_root_r119_SUM_12_), .B_11_(
        add_1_root_r119_SUM_11_), .B_10_(add_1_root_r119_SUM_10_), .B_9_(
        add_1_root_r119_SUM_9_), .B_8_(add_1_root_r119_SUM_8_), .B_7_(
        add_1_root_r119_SUM_7_), .B_6_(add_1_root_r119_SUM_6_), .B_5_(
        add_1_root_r119_A_5_), .B_4_(add_1_root_r119_A_4_), .SUM_23_(N363), 
        .SUM_22_(N362), .SUM_21_(N361), .SUM_20_(N360), .SUM_19_(N359), 
        .SUM_18_(N358), .SUM_17_(N357), .SUM_16_(N356), .SUM_15_(N355), 
        .SUM_14_(N354), .SUM_13_(N353), .SUM_12_(N352), .SUM_11_(N351), 
        .SUM_10_(N350), .SUM_9_(N349), .SUM_8_(N348), .SUM_7_(N347) );
  multi16_5_DW01_add_4 add_0_root_r112 ( .A_21_(in_17bit_b[16]), .A_20_(
        in_17bit_b[15]), .A_19_(in_17bit_b[14]), .A_18_(in_17bit_b[13]), 
        .A_17_(in_17bit_b[12]), .A_16_(in_17bit_b[11]), .A_15_(in_17bit_b[10]), 
        .A_14_(in_17bit_b[9]), .A_13_(in_17bit_b[8]), .A_12_(in_17bit_b[7]), 
        .A_11_(in_17bit_b[6]), .A_10_(in_17bit_b[5]), .A_9_(in_17bit_b[4]), 
        .A_8_(in_17bit_b[3]), .A_7_(in_17bit_b[2]), .A_6_(in_17bit_b[1]), 
        .A_5_(in_17bit_b[0]), .B_21_(add_1_root_r112_SUM_21_), .B_20_(
        add_1_root_r112_SUM_20_), .B_19_(add_1_root_r112_SUM_19_), .B_18_(
        add_1_root_r112_SUM_18_), .B_17_(add_1_root_r112_SUM_17_), .B_16_(
        add_1_root_r112_SUM_16_), .B_15_(add_1_root_r112_SUM_15_), .B_14_(
        add_1_root_r112_SUM_14_), .B_13_(add_1_root_r112_SUM_13_), .B_12_(
        add_1_root_r112_SUM_12_), .B_11_(add_1_root_r112_SUM_11_), .B_10_(
        add_1_root_r112_SUM_10_), .B_9_(add_1_root_r112_SUM_9_), .B_8_(
        add_1_root_r112_SUM_8_), .B_7_(add_1_root_r112_SUM_7_), .B_6_(
        add_1_root_r112_SUM_6_), .B_5_(add_1_root_r112_SUM_5_), .SUM_22_(N123), 
        .SUM_21_(N122), .SUM_20_(N121), .SUM_19_(N120), .SUM_18_(N119), 
        .SUM_17_(N118), .SUM_16_(N117), .SUM_15_(N116), .SUM_14_(N115), 
        .SUM_13_(N114), .SUM_12_(N113), .SUM_11_(N112), .SUM_10_(N111), 
        .SUM_9_(N110), .SUM_8_(N109), .SUM_7_(N108) );
  multi16_5_DW01_add_6 add_0_root_r115 ( .A_23_(add_1_root_r115_SUM_23_), 
        .A_22_(add_1_root_r115_SUM_22_), .A_21_(add_1_root_r115_SUM_21_), 
        .A_20_(add_1_root_r115_SUM_20_), .A_19_(add_1_root_r115_SUM_19_), 
        .A_18_(add_1_root_r115_SUM_18_), .A_17_(add_1_root_r115_SUM_17_), 
        .A_16_(add_1_root_r115_SUM_16_), .A_15_(add_1_root_r115_SUM_15_), 
        .A_14_(add_1_root_r115_SUM_14_), .A_13_(add_1_root_r115_SUM_13_), 
        .A_12_(add_1_root_r115_SUM_12_), .A_11_(add_1_root_r115_SUM_11_), 
        .A_10_(add_1_root_r115_SUM_10_), .A_9_(add_1_root_r115_SUM_9_), .A_8_(
        add_1_root_r115_SUM_8_), .A_7_(add_1_root_r115_SUM_7_), .A_6_(
        add_1_root_r115_SUM_6_), .A_5_(in_17bit_b[1]), .A_4_(in_17bit_b[0]), 
        .B_20_(add_2_root_r115_SUM_20_), .B_19_(add_2_root_r115_SUM_19_), 
        .B_18_(add_2_root_r115_SUM_18_), .B_17_(add_2_root_r115_SUM_17_), 
        .B_16_(add_2_root_r115_SUM_16_), .B_15_(add_2_root_r115_SUM_15_), 
        .B_14_(add_2_root_r115_SUM_14_), .B_13_(add_2_root_r115_SUM_13_), 
        .B_12_(add_2_root_r115_SUM_12_), .B_11_(add_2_root_r115_SUM_11_), 
        .B_10_(add_2_root_r115_SUM_10_), .B_9_(add_2_root_r115_SUM_9_), .B_8_(
        add_2_root_r115_SUM_8_), .B_7_(add_2_root_r115_SUM_7_), .B_6_(
        add_2_root_r115_SUM_6_), .B_5_(add_2_root_r115_SUM_5_), .B_4_(
        add_2_root_r115_SUM_4_), .SUM_23_(N221), .SUM_22_(N220), .SUM_21_(N219), .SUM_20_(N218), .SUM_19_(N217), .SUM_18_(N216), .SUM_17_(N215), .SUM_16_(
        N214), .SUM_15_(N213), .SUM_14_(N212), .SUM_13_(N211), .SUM_12_(N210), 
        .SUM_11_(N209), .SUM_10_(N208), .SUM_9_(N207), .SUM_8_(N206), .SUM_7_(
        N205) );
  TLATX1 neg_mul_reg_18_ ( .G(N446), .D(N458), .QN(n18) );
  TLATX1 neg_mul_reg_17_ ( .G(N446), .D(N457), .QN(n17) );
  TLATX1 neg_mul_reg_16_ ( .G(N446), .D(N456), .QN(n16) );
  TLATX1 neg_mul_reg_15_ ( .G(N446), .D(N455), .QN(n12) );
  TLATX1 neg_mul_reg_14_ ( .G(N446), .D(N454), .QN(n15) );
  TLATX1 neg_mul_reg_13_ ( .G(N446), .D(N453), .Q(n3), .QN(n14) );
  TLATX1 neg_mul_reg_12_ ( .G(N446), .D(N452), .QN(n13) );
  TLATX1 neg_mul_reg_11_ ( .G(N446), .D(N451), .Q(neg_mul[11]), .QN(n9) );
  TLATX1 neg_mul_reg_9_ ( .G(N446), .D(N449), .Q(neg_mul[9]), .QN(n8) );
  TLATX1 neg_mul_reg_23_ ( .G(N446), .D(N463), .Q(neg_mul[23]), .QN(n10) );
  TLATX1 neg_mul_reg_22_ ( .G(N446), .D(N462), .Q(neg_mul[22]), .QN(n19) );
  TLATX1 neg_mul_reg_21_ ( .G(N446), .D(N461), .Q(neg_mul[21]), .QN(n21) );
  TLATX1 neg_mul_reg_20_ ( .G(N446), .D(N460), .Q(neg_mul[20]), .QN(n22) );
  TLATX1 neg_mul_reg_19_ ( .G(N446), .D(N459), .QN(n23) );
  TLATX1 neg_mul_reg_8_ ( .G(N446), .D(N448), .Q(neg_mul[8]) );
  TLATX1 neg_mul_reg_10_ ( .G(N446), .D(N450), .Q(neg_mul[10]), .QN(n7) );
  TLATX1 neg_mul_reg_7_ ( .G(N446), .D(N447), .Q(out[0]), .QN(n20) );
  INVXL U2 ( .A(n56), .Y(n1) );
  CLKINVX3 U3 ( .A(n45), .Y(n5) );
  XOR2X4 U4 ( .A(n74), .B(n2), .Y(out[7]) );
  CLKINVX20 U5 ( .A(n15), .Y(n2) );
  XOR2X4 U6 ( .A(n72), .B(n3), .Y(out[6]) );
  BUFX2 U7 ( .A(n77), .Y(n4) );
  INVX4 U8 ( .A(n4), .Y(n78) );
  XNOR2X4 U9 ( .A(in_8bit[7]), .B(n27), .Y(n77) );
  INVX4 U10 ( .A(in_8bit[7]), .Y(n45) );
  XNOR2X4 U11 ( .A(n5), .B(n27), .Y(n59) );
  CLKINVX3 U12 ( .A(n252), .Y(in_17bit_b[16]) );
  NOR2X4 U13 ( .A(n6), .B(n68), .Y(n70) );
  CLKINVX20 U14 ( .A(n57), .Y(n6) );
  XNOR2X4 U15 ( .A(n75), .B(n16), .Y(out[9]) );
  NOR2X2 U16 ( .A(n73), .B(n32), .Y(n71) );
  XNOR2X2 U17 ( .A(n28), .B(n12), .Y(out[8]) );
  OR3X4 U18 ( .A(n67), .B(n69), .C(n66), .Y(n11) );
  XNOR2X1 U19 ( .A(neg_mul[23]), .B(n41), .Y(n24) );
  BUFX20 U20 ( .A(in_17bit[16]), .Y(n25) );
  NOR2X1 U21 ( .A(n77), .B(n38), .Y(n29) );
  AOI2BB2X2 U22 ( .B0(n62), .B1(n43), .A0N(n43), .A1N(neg_mul[10]), .Y(n63) );
  INVXL U23 ( .A(n1), .Y(n53) );
  INVX8 U24 ( .A(n25), .Y(n56) );
  INVX8 U25 ( .A(n11), .Y(out[3]) );
  XNOR2X4 U26 ( .A(n56), .B(n45), .Y(n73) );
  BUFX20 U27 ( .A(n25), .Y(n27) );
  NOR2X2 U28 ( .A(n77), .B(n35), .Y(n28) );
  XOR2X4 U29 ( .A(n70), .B(neg_mul[11]), .Y(out[4]) );
  NOR2X4 U30 ( .A(n34), .B(n77), .Y(n74) );
  NOR2X4 U31 ( .A(n40), .B(n73), .Y(n60) );
  AOI2BB2X2 U32 ( .B0(n43), .B1(n7), .A0N(n43), .A1N(n64), .Y(n65) );
  CLKINVX4 U33 ( .A(n45), .Y(n43) );
  INVX8 U34 ( .A(n56), .Y(n54) );
  NOR2X1 U35 ( .A(n59), .B(n36), .Y(n75) );
  XNOR2X4 U36 ( .A(n29), .B(n18), .Y(out[11]) );
  XOR2X4 U37 ( .A(n60), .B(neg_mul[9]), .Y(out[2]) );
  XOR2X4 U38 ( .A(n45), .B(n27), .Y(n68) );
  NOR2X4 U39 ( .A(n33), .B(n68), .Y(n72) );
  NOR2BX4 U40 ( .AN(n54), .B(n65), .Y(n66) );
  NOR2X2 U41 ( .A(n77), .B(n37), .Y(n76) );
  MX2X1 U42 ( .A(neg_mul[21]), .B(N479), .S0(n78), .Y(out[14]) );
  INVXL U43 ( .A(n45), .Y(n44) );
  INVX1 U44 ( .A(n202), .Y(in_17bit_b[1]) );
  INVX1 U45 ( .A(n241), .Y(in_17bit_b[14]) );
  INVX1 U46 ( .A(n238), .Y(in_17bit_b[13]) );
  INVX1 U47 ( .A(n205), .Y(in_17bit_b[2]) );
  INVX1 U48 ( .A(n214), .Y(in_17bit_b[5]) );
  INVX1 U49 ( .A(n217), .Y(in_17bit_b[6]) );
  INVX1 U50 ( .A(n220), .Y(in_17bit_b[7]) );
  INVX1 U51 ( .A(n229), .Y(in_17bit_b[10]) );
  INVX1 U52 ( .A(n223), .Y(in_17bit_b[8]) );
  INVX1 U53 ( .A(n226), .Y(in_17bit_b[9]) );
  INVX1 U54 ( .A(n232), .Y(in_17bit_b[11]) );
  INVX1 U55 ( .A(n235), .Y(in_17bit_b[12]) );
  INVX1 U56 ( .A(n211), .Y(in_17bit_b[4]) );
  INVX1 U57 ( .A(n208), .Y(in_17bit_b[3]) );
  AOI21X1 U58 ( .A0(n30), .A1(n31), .B0(n245), .Y(n198) );
  NOR4XL U59 ( .A(in_8bit[4]), .B(n47), .C(in_8bit[6]), .D(n44), .Y(n30) );
  NOR4XL U60 ( .A(in_8bit[1]), .B(in_8bit[0]), .C(in_8bit[2]), .D(in_8bit[3]), 
        .Y(n31) );
  NOR2X2 U61 ( .A(n54), .B(n63), .Y(n67) );
  MX2X1 U62 ( .A(neg_mul[20]), .B(N478), .S0(n78), .Y(out[13]) );
  NAND3X1 U63 ( .A(in_8bit[2]), .B(n49), .C(n47), .Y(n193) );
  NAND3BX1 U64 ( .AN(n47), .B(n46), .C(in_8bit[3]), .Y(n194) );
  NAND3X1 U65 ( .A(n44), .B(n50), .C(n48), .Y(n88) );
  INVX1 U66 ( .A(n48), .Y(n47) );
  INVX1 U67 ( .A(n170), .Y(n251) );
  OAI21XL U68 ( .A0(n251), .A1(n252), .B0(n250), .Y(N463) );
  AOI22X1 U69 ( .A0(N221), .A1(n249), .B0(N363), .B1(n248), .Y(n250) );
  ADDFX2 U70 ( .A(in_17bit_b[16]), .B(in_17bit_b[12]), .CI(
        add_1_root_r112_carry_16_), .CO(add_1_root_r112_carry_17_), .S(
        add_1_root_r112_SUM_16_) );
  ADDFX2 U71 ( .A(add_1_root_r119_A_19_), .B(in_17bit_b[13]), .CI(
        add_1_root_r119_carry[19]), .CO(add_1_root_r119_carry[20]), .S(
        add_1_root_r119_SUM_19_) );
  ADDFX2 U72 ( .A(in_17bit_b[16]), .B(in_17bit_b[15]), .CI(
        add_3_root_r119_carry_17_), .CO(add_3_root_r119_carry_18_), .S(
        add_1_root_r119_A_17_) );
  ADDFX2 U73 ( .A(in_17bit_b[16]), .B(in_17bit_b[14]), .CI(
        add_2_root_r115_carry_17_), .CO(add_2_root_r115_carry_18_), .S(
        add_2_root_r115_SUM_17_) );
  ADDFX2 U74 ( .A(in_17bit_b[16]), .B(in_17bit_b[14]), .CI(
        add_1_root_r115_carry_20_), .CO(add_1_root_r115_carry_21_), .S(
        add_1_root_r115_SUM_20_) );
  ADDFX2 U75 ( .A(in_17bit_b[16]), .B(in_17bit_b[15]), .CI(
        add_2_root_r119_carry_20_), .CO(add_2_root_r119_carry_21_), .S(
        add_2_root_r119_SUM_20_) );
  ADDFX2 U76 ( .A(in_17bit_b[3]), .B(in_17bit_b[1]), .CI(
        add_2_root_r115_carry_4_), .CO(add_2_root_r115_carry_5_), .S(
        add_2_root_r115_SUM_4_) );
  ADDFX2 U77 ( .A(in_17bit_b[4]), .B(in_17bit_b[2]), .CI(
        add_2_root_r115_carry_5_), .CO(add_2_root_r115_carry_6_), .S(
        add_2_root_r115_SUM_5_) );
  ADDFX2 U78 ( .A(in_17bit_b[5]), .B(in_17bit_b[1]), .CI(
        add_1_root_r112_carry_5_), .CO(add_1_root_r112_carry_6_), .S(
        add_1_root_r112_SUM_5_) );
  ADDFX2 U79 ( .A(in_17bit_b[6]), .B(in_17bit_b[5]), .CI(
        add_3_root_r119_carry_7_), .CO(add_3_root_r119_carry_8_), .S(
        add_1_root_r119_A_7_) );
  ADDFX2 U80 ( .A(in_17bit_b[6]), .B(in_17bit_b[2]), .CI(
        add_1_root_r112_carry_6_), .CO(add_1_root_r112_carry_7_), .S(
        add_1_root_r112_SUM_6_) );
  ADDFX2 U81 ( .A(in_17bit_b[3]), .B(in_17bit_b[1]), .CI(
        add_2_root_r115_carry_4_), .CO(add_1_root_r115_carry_8_), .S(
        add_1_root_r115_SUM_7_) );
  ADDFX2 U82 ( .A(in_17bit_b[7]), .B(in_17bit_b[6]), .CI(
        add_3_root_r119_carry_8_), .CO(add_3_root_r119_carry_9_), .S(
        add_1_root_r119_A_8_) );
  ADDFX2 U83 ( .A(add_1_root_r119_A_7_), .B(in_17bit_b[1]), .CI(
        add_1_root_r119_carry[7]), .CO(add_1_root_r119_carry[8]), .S(
        add_1_root_r119_SUM_7_) );
  ADDFX2 U84 ( .A(in_17bit_b[2]), .B(in_17bit_b[1]), .CI(
        add_2_root_r119_carry_6_), .CO(add_2_root_r119_carry_7_), .S(
        add_2_root_r119_SUM_6_) );
  ADDFX2 U85 ( .A(in_17bit_b[4]), .B(in_17bit_b[2]), .CI(
        add_1_root_r115_carry_8_), .CO(add_1_root_r115_carry_9_), .S(
        add_1_root_r115_SUM_8_) );
  ADDFX2 U86 ( .A(in_17bit_b[8]), .B(in_17bit_b[7]), .CI(
        add_3_root_r119_carry_9_), .CO(add_3_root_r119_carry_10_), .S(
        add_1_root_r119_A_9_) );
  ADDFX2 U87 ( .A(add_1_root_r119_A_8_), .B(in_17bit_b[2]), .CI(
        add_1_root_r119_carry[8]), .CO(add_1_root_r119_carry[9]), .S(
        add_1_root_r119_SUM_8_) );
  ADDFX2 U88 ( .A(in_17bit_b[3]), .B(in_17bit_b[2]), .CI(
        add_2_root_r119_carry_7_), .CO(add_2_root_r119_carry_8_), .S(
        add_2_root_r119_SUM_7_) );
  ADDFX2 U89 ( .A(in_17bit_b[6]), .B(in_17bit_b[4]), .CI(
        add_2_root_r115_carry_7_), .CO(add_2_root_r115_carry_8_), .S(
        add_2_root_r115_SUM_7_) );
  ADDFX2 U90 ( .A(in_17bit_b[9]), .B(in_17bit_b[8]), .CI(
        add_3_root_r119_carry_10_), .CO(add_3_root_r119_carry_11_), .S(
        add_1_root_r119_A_10_) );
  ADDFX2 U91 ( .A(in_17bit_b[7]), .B(in_17bit_b[5]), .CI(
        add_2_root_r115_carry_8_), .CO(add_2_root_r115_carry_9_), .S(
        add_2_root_r115_SUM_8_) );
  ADDFX2 U92 ( .A(in_17bit_b[9]), .B(in_17bit_b[5]), .CI(
        add_1_root_r112_carry_9_), .CO(add_1_root_r112_carry_10_), .S(
        add_1_root_r112_SUM_9_) );
  ADDFX2 U93 ( .A(in_17bit_b[6]), .B(in_17bit_b[4]), .CI(
        add_1_root_r115_carry_10_), .CO(add_1_root_r115_carry_11_), .S(
        add_1_root_r115_SUM_10_) );
  ADDFX2 U94 ( .A(in_17bit_b[10]), .B(in_17bit_b[9]), .CI(
        add_3_root_r119_carry_11_), .CO(add_3_root_r119_carry_12_), .S(
        add_1_root_r119_A_11_) );
  ADDFX2 U95 ( .A(add_1_root_r119_A_10_), .B(in_17bit_b[4]), .CI(
        add_1_root_r119_carry[10]), .CO(add_1_root_r119_carry[11]), .S(
        add_1_root_r119_SUM_10_) );
  ADDFX2 U96 ( .A(in_17bit_b[8]), .B(in_17bit_b[6]), .CI(
        add_2_root_r115_carry_9_), .CO(add_2_root_r115_carry_10_), .S(
        add_2_root_r115_SUM_9_) );
  ADDFX2 U97 ( .A(in_17bit_b[7]), .B(in_17bit_b[5]), .CI(
        add_1_root_r115_carry_11_), .CO(add_1_root_r115_carry_12_), .S(
        add_1_root_r115_SUM_11_) );
  ADDFX2 U98 ( .A(in_17bit_b[11]), .B(in_17bit_b[10]), .CI(
        add_3_root_r119_carry_12_), .CO(add_3_root_r119_carry_13_), .S(
        add_1_root_r119_A_12_) );
  ADDFX2 U99 ( .A(add_1_root_r119_A_11_), .B(in_17bit_b[5]), .CI(
        add_1_root_r119_carry[11]), .CO(add_1_root_r119_carry[12]), .S(
        add_1_root_r119_SUM_11_) );
  ADDFX2 U100 ( .A(in_17bit_b[6]), .B(in_17bit_b[5]), .CI(
        add_2_root_r119_carry_10_), .CO(add_2_root_r119_carry_11_), .S(
        add_2_root_r119_SUM_10_) );
  ADDFX2 U101 ( .A(in_17bit_b[9]), .B(in_17bit_b[7]), .CI(
        add_2_root_r115_carry_10_), .CO(add_2_root_r115_carry_11_), .S(
        add_2_root_r115_SUM_10_) );
  ADDFX2 U102 ( .A(in_17bit_b[11]), .B(in_17bit_b[7]), .CI(
        add_1_root_r112_carry_11_), .CO(add_1_root_r112_carry_12_), .S(
        add_1_root_r112_SUM_11_) );
  ADDFX2 U103 ( .A(in_17bit_b[8]), .B(in_17bit_b[6]), .CI(
        add_1_root_r115_carry_12_), .CO(add_1_root_r115_carry_13_), .S(
        add_1_root_r115_SUM_12_) );
  ADDFX2 U104 ( .A(in_17bit_b[12]), .B(in_17bit_b[11]), .CI(
        add_3_root_r119_carry_13_), .CO(add_3_root_r119_carry_14_), .S(
        add_1_root_r119_A_13_) );
  ADDFX2 U105 ( .A(add_1_root_r119_A_12_), .B(in_17bit_b[6]), .CI(
        add_1_root_r119_carry[12]), .CO(add_1_root_r119_carry[13]), .S(
        add_1_root_r119_SUM_12_) );
  ADDFX2 U106 ( .A(in_17bit_b[7]), .B(in_17bit_b[6]), .CI(
        add_2_root_r119_carry_11_), .CO(add_2_root_r119_carry_12_), .S(
        add_2_root_r119_SUM_11_) );
  ADDFX2 U107 ( .A(in_17bit_b[10]), .B(in_17bit_b[8]), .CI(
        add_2_root_r115_carry_11_), .CO(add_2_root_r115_carry_12_), .S(
        add_2_root_r115_SUM_11_) );
  ADDFX2 U108 ( .A(in_17bit_b[12]), .B(in_17bit_b[8]), .CI(
        add_1_root_r112_carry_12_), .CO(add_1_root_r112_carry_13_), .S(
        add_1_root_r112_SUM_12_) );
  ADDFX2 U109 ( .A(in_17bit_b[9]), .B(in_17bit_b[7]), .CI(
        add_1_root_r115_carry_13_), .CO(add_1_root_r115_carry_14_), .S(
        add_1_root_r115_SUM_13_) );
  ADDFX2 U110 ( .A(in_17bit_b[13]), .B(in_17bit_b[12]), .CI(
        add_3_root_r119_carry_14_), .CO(add_3_root_r119_carry_15_), .S(
        add_1_root_r119_A_14_) );
  ADDFX2 U111 ( .A(add_1_root_r119_A_13_), .B(in_17bit_b[7]), .CI(
        add_1_root_r119_carry[13]), .CO(add_1_root_r119_carry[14]), .S(
        add_1_root_r119_SUM_13_) );
  ADDFX2 U112 ( .A(in_17bit_b[8]), .B(in_17bit_b[7]), .CI(
        add_2_root_r119_carry_12_), .CO(add_2_root_r119_carry_13_), .S(
        add_2_root_r119_SUM_12_) );
  ADDFX2 U113 ( .A(in_17bit_b[11]), .B(in_17bit_b[9]), .CI(
        add_2_root_r115_carry_12_), .CO(add_2_root_r115_carry_13_), .S(
        add_2_root_r115_SUM_12_) );
  ADDFX2 U114 ( .A(in_17bit_b[13]), .B(in_17bit_b[9]), .CI(
        add_1_root_r112_carry_13_), .CO(add_1_root_r112_carry_14_), .S(
        add_1_root_r112_SUM_13_) );
  ADDFX2 U115 ( .A(in_17bit_b[14]), .B(in_17bit_b[13]), .CI(
        add_3_root_r119_carry_15_), .CO(add_3_root_r119_carry_16_), .S(
        add_1_root_r119_A_15_) );
  ADDFX2 U116 ( .A(add_1_root_r119_A_14_), .B(in_17bit_b[8]), .CI(
        add_1_root_r119_carry[14]), .CO(add_1_root_r119_carry[15]), .S(
        add_1_root_r119_SUM_14_) );
  ADDFX2 U117 ( .A(in_17bit_b[9]), .B(in_17bit_b[8]), .CI(
        add_2_root_r119_carry_13_), .CO(add_2_root_r119_carry_14_), .S(
        add_2_root_r119_SUM_13_) );
  ADDFX2 U118 ( .A(in_17bit_b[12]), .B(in_17bit_b[10]), .CI(
        add_2_root_r115_carry_13_), .CO(add_2_root_r115_carry_14_), .S(
        add_2_root_r115_SUM_13_) );
  ADDFX2 U119 ( .A(in_17bit_b[14]), .B(in_17bit_b[10]), .CI(
        add_1_root_r112_carry_14_), .CO(add_1_root_r112_carry_15_), .S(
        add_1_root_r112_SUM_14_) );
  ADDFX2 U120 ( .A(in_17bit_b[11]), .B(in_17bit_b[9]), .CI(
        add_1_root_r115_carry_15_), .CO(add_1_root_r115_carry_16_), .S(
        add_1_root_r115_SUM_15_) );
  ADDFX2 U121 ( .A(add_1_root_r119_A_15_), .B(in_17bit_b[9]), .CI(
        add_1_root_r119_carry[15]), .CO(add_1_root_r119_carry[16]), .S(
        add_1_root_r119_SUM_15_) );
  ADDFX2 U122 ( .A(in_17bit_b[3]), .B(in_17bit_b[2]), .CI(
        add_3_root_r119_carry_4_), .CO(add_3_root_r119_carry_5_), .S(
        add_1_root_r119_A_4_) );
  ADDFX2 U123 ( .A(in_17bit_b[2]), .B(in_17bit_b[1]), .CI(
        add_2_root_r119_carry_6_), .CO(add_3_root_r119_carry_4_), .S(
        add_1_root_r119_A_3_) );
  ADDFX2 U124 ( .A(in_17bit_b[10]), .B(in_17bit_b[9]), .CI(
        add_2_root_r119_carry_14_), .CO(add_2_root_r119_carry_15_), .S(
        add_2_root_r119_SUM_14_) );
  ADDFX2 U125 ( .A(in_17bit_b[13]), .B(in_17bit_b[11]), .CI(
        add_2_root_r115_carry_14_), .CO(add_2_root_r115_carry_15_), .S(
        add_2_root_r115_SUM_14_) );
  ADDFX2 U126 ( .A(in_17bit_b[15]), .B(in_17bit_b[11]), .CI(
        add_1_root_r112_carry_15_), .CO(add_1_root_r112_carry_16_), .S(
        add_1_root_r112_SUM_15_) );
  ADDFX2 U127 ( .A(in_17bit_b[12]), .B(in_17bit_b[10]), .CI(
        add_1_root_r115_carry_16_), .CO(add_1_root_r115_carry_17_), .S(
        add_1_root_r115_SUM_16_) );
  ADDFX2 U128 ( .A(add_1_root_r119_A_16_), .B(in_17bit_b[10]), .CI(
        add_1_root_r119_carry[16]), .CO(add_1_root_r119_carry[17]), .S(
        add_1_root_r119_SUM_16_) );
  ADDFX2 U129 ( .A(in_17bit_b[11]), .B(in_17bit_b[10]), .CI(
        add_2_root_r119_carry_15_), .CO(add_2_root_r119_carry_16_), .S(
        add_2_root_r119_SUM_15_) );
  ADDFX2 U130 ( .A(in_17bit_b[14]), .B(in_17bit_b[12]), .CI(
        add_2_root_r115_carry_15_), .CO(add_2_root_r115_carry_16_), .S(
        add_2_root_r115_SUM_15_) );
  ADDFX2 U131 ( .A(add_1_root_r119_A_17_), .B(in_17bit_b[11]), .CI(
        add_1_root_r119_carry[17]), .CO(add_1_root_r119_carry[18]), .S(
        add_1_root_r119_SUM_17_) );
  ADDFX2 U132 ( .A(in_17bit_b[12]), .B(in_17bit_b[11]), .CI(
        add_2_root_r119_carry_16_), .CO(add_2_root_r119_carry_17_), .S(
        add_2_root_r119_SUM_16_) );
  ADDFX2 U133 ( .A(in_17bit_b[15]), .B(in_17bit_b[13]), .CI(
        add_2_root_r115_carry_16_), .CO(add_2_root_r115_carry_17_), .S(
        add_2_root_r115_SUM_16_) );
  ADDFX2 U134 ( .A(in_17bit_b[14]), .B(in_17bit_b[12]), .CI(
        add_1_root_r115_carry_18_), .CO(add_1_root_r115_carry_19_), .S(
        add_1_root_r115_SUM_18_) );
  ADDFX2 U135 ( .A(add_1_root_r119_A_18_), .B(in_17bit_b[12]), .CI(
        add_1_root_r119_carry[18]), .CO(add_1_root_r119_carry[19]), .S(
        add_1_root_r119_SUM_18_) );
  ADDFX2 U136 ( .A(in_17bit_b[13]), .B(in_17bit_b[12]), .CI(
        add_2_root_r119_carry_17_), .CO(add_2_root_r119_carry_18_), .S(
        add_2_root_r119_SUM_17_) );
  ADDFX2 U137 ( .A(in_17bit_b[13]), .B(in_17bit_b[11]), .CI(
        add_1_root_r115_carry_17_), .CO(add_1_root_r115_carry_18_), .S(
        add_1_root_r115_SUM_17_) );
  ADDFX2 U138 ( .A(in_17bit_b[7]), .B(in_17bit_b[3]), .CI(
        add_1_root_r112_carry_7_), .CO(add_1_root_r112_carry_8_), .S(
        add_1_root_r112_SUM_7_) );
  ADDFX2 U139 ( .A(in_17bit_b[8]), .B(in_17bit_b[4]), .CI(
        add_1_root_r112_carry_8_), .CO(add_1_root_r112_carry_9_), .S(
        add_1_root_r112_SUM_8_) );
  ADDFX2 U140 ( .A(in_17bit_b[5]), .B(in_17bit_b[3]), .CI(
        add_1_root_r115_carry_9_), .CO(add_1_root_r115_carry_10_), .S(
        add_1_root_r115_SUM_9_) );
  ADDFX2 U141 ( .A(add_1_root_r119_A_9_), .B(in_17bit_b[3]), .CI(
        add_1_root_r119_carry[9]), .CO(add_1_root_r119_carry[10]), .S(
        add_1_root_r119_SUM_9_) );
  ADDFX2 U142 ( .A(in_17bit_b[4]), .B(in_17bit_b[3]), .CI(
        add_2_root_r119_carry_8_), .CO(add_2_root_r119_carry_9_), .S(
        add_2_root_r119_SUM_8_) );
  ADDFX2 U143 ( .A(in_17bit_b[5]), .B(in_17bit_b[4]), .CI(
        add_2_root_r119_carry_9_), .CO(add_2_root_r119_carry_10_), .S(
        add_2_root_r119_SUM_9_) );
  ADDFX2 U144 ( .A(in_17bit_b[10]), .B(in_17bit_b[6]), .CI(
        add_1_root_r112_carry_10_), .CO(add_1_root_r112_carry_11_), .S(
        add_1_root_r112_SUM_10_) );
  ADDFX2 U145 ( .A(in_17bit_b[10]), .B(in_17bit_b[8]), .CI(
        add_1_root_r115_carry_14_), .CO(add_1_root_r115_carry_15_), .S(
        add_1_root_r115_SUM_14_) );
  ADDFX2 U146 ( .A(in_17bit_b[15]), .B(in_17bit_b[14]), .CI(
        add_3_root_r119_carry_16_), .CO(add_3_root_r119_carry_17_), .S(
        add_1_root_r119_A_16_) );
  ADDFX2 U147 ( .A(in_17bit_b[5]), .B(in_17bit_b[3]), .CI(
        add_2_root_r115_carry_6_), .CO(add_2_root_r115_carry_7_), .S(
        add_2_root_r115_SUM_6_) );
  ADDFX2 U148 ( .A(in_17bit_b[4]), .B(in_17bit_b[3]), .CI(
        add_3_root_r119_carry_5_), .CO(add_3_root_r119_carry_6_), .S(
        add_1_root_r119_A_5_) );
  ADDFX2 U149 ( .A(in_17bit_b[5]), .B(in_17bit_b[4]), .CI(
        add_3_root_r119_carry_6_), .CO(add_3_root_r119_carry_7_), .S(
        add_1_root_r119_A_6_) );
  ADDFX2 U150 ( .A(in_17bit_b[15]), .B(in_17bit_b[13]), .CI(
        add_1_root_r115_carry_19_), .CO(add_1_root_r115_carry_20_), .S(
        add_1_root_r115_SUM_19_) );
  ADDFX2 U151 ( .A(in_17bit_b[14]), .B(in_17bit_b[13]), .CI(
        add_2_root_r119_carry_18_), .CO(add_2_root_r119_carry_19_), .S(
        add_2_root_r119_SUM_18_) );
  ADDFX2 U152 ( .A(in_17bit_b[15]), .B(in_17bit_b[14]), .CI(
        add_2_root_r119_carry_19_), .CO(add_2_root_r119_carry_20_), .S(
        add_2_root_r119_SUM_19_) );
  INVXL U153 ( .A(n53), .Y(n52) );
  INVX1 U154 ( .A(in_8bit[2]), .Y(n46) );
  INVX1 U155 ( .A(n52), .Y(n55) );
  INVX1 U156 ( .A(in_8bit[4]), .Y(n50) );
  INVX1 U157 ( .A(in_8bit[3]), .Y(n49) );
  INVX1 U158 ( .A(in_8bit[6]), .Y(n51) );
  INVX1 U159 ( .A(in_8bit[5]), .Y(n48) );
  NOR3X1 U160 ( .A(n46), .B(n49), .C(n171), .Y(n197) );
  CLKINVX3 U161 ( .A(n199), .Y(in_17bit_b[0]) );
  NAND2XL U162 ( .A(N29), .B(n1), .Y(n252) );
  CLKINVX3 U163 ( .A(n244), .Y(in_17bit_b[15]) );
  OR2X2 U164 ( .A(n84), .B(n83), .Y(n248) );
  NOR2X1 U165 ( .A(n85), .B(n193), .Y(n83) );
  NOR2X1 U166 ( .A(n194), .B(n192), .Y(n84) );
  OR2X2 U167 ( .A(n87), .B(n86), .Y(n249) );
  NOR2X1 U168 ( .A(n85), .B(n194), .Y(n86) );
  NOR2X1 U169 ( .A(n193), .B(n192), .Y(n87) );
  OAI2BB1X1 U170 ( .A0N(n196), .A1N(n91), .B0(n90), .Y(n170) );
  INVX1 U171 ( .A(n88), .Y(n91) );
  NAND3BX1 U172 ( .AN(n89), .B(n197), .C(n47), .Y(n90) );
  NAND3X1 U173 ( .A(n196), .B(n47), .C(n79), .Y(n80) );
  NOR2X1 U174 ( .A(n44), .B(n50), .Y(n79) );
  NAND2X1 U175 ( .A(n201), .B(n200), .Y(N447) );
  AOI22X1 U176 ( .A0(N108), .A1(n245), .B0(N205), .B1(n249), .Y(n200) );
  AOI22X1 U177 ( .A0(N347), .A1(n248), .B0(n170), .B1(in_17bit_b[0]), .Y(n201)
         );
  NAND2X1 U178 ( .A(n204), .B(n203), .Y(N448) );
  AOI22X1 U179 ( .A0(N109), .A1(n245), .B0(N206), .B1(n249), .Y(n203) );
  AOI22X1 U180 ( .A0(N348), .A1(n248), .B0(n170), .B1(in_17bit_b[1]), .Y(n204)
         );
  NAND2X1 U181 ( .A(n207), .B(n206), .Y(N449) );
  AOI22X1 U182 ( .A0(N110), .A1(n245), .B0(N207), .B1(n249), .Y(n206) );
  AOI22X1 U183 ( .A0(N349), .A1(n248), .B0(n170), .B1(in_17bit_b[2]), .Y(n207)
         );
  NAND2X1 U184 ( .A(n210), .B(n209), .Y(N450) );
  AOI22X1 U185 ( .A0(N111), .A1(n245), .B0(N208), .B1(n249), .Y(n209) );
  AOI22X1 U186 ( .A0(N350), .A1(n248), .B0(n170), .B1(in_17bit_b[3]), .Y(n210)
         );
  NAND2X1 U187 ( .A(n213), .B(n212), .Y(N451) );
  AOI22X1 U188 ( .A0(N112), .A1(n245), .B0(N209), .B1(n249), .Y(n212) );
  AOI22X1 U189 ( .A0(N351), .A1(n248), .B0(n170), .B1(in_17bit_b[4]), .Y(n213)
         );
  NAND2X1 U190 ( .A(n216), .B(n215), .Y(N452) );
  AOI22X1 U191 ( .A0(N113), .A1(n245), .B0(N210), .B1(n249), .Y(n215) );
  AOI22X1 U192 ( .A0(N352), .A1(n248), .B0(n170), .B1(in_17bit_b[5]), .Y(n216)
         );
  NAND2X1 U193 ( .A(n219), .B(n218), .Y(N453) );
  AOI22X1 U194 ( .A0(N114), .A1(n245), .B0(N211), .B1(n249), .Y(n218) );
  AOI22X1 U195 ( .A0(N353), .A1(n248), .B0(n170), .B1(in_17bit_b[6]), .Y(n219)
         );
  NAND2X1 U196 ( .A(n222), .B(n221), .Y(N454) );
  AOI22X1 U197 ( .A0(N115), .A1(n245), .B0(N212), .B1(n249), .Y(n221) );
  AOI22X1 U198 ( .A0(N354), .A1(n248), .B0(n170), .B1(in_17bit_b[7]), .Y(n222)
         );
  NAND2X1 U199 ( .A(n225), .B(n224), .Y(N455) );
  AOI22X1 U200 ( .A0(N116), .A1(n245), .B0(N213), .B1(n249), .Y(n224) );
  AOI22X1 U201 ( .A0(N355), .A1(n248), .B0(n170), .B1(in_17bit_b[8]), .Y(n225)
         );
  NAND2X1 U202 ( .A(n228), .B(n227), .Y(N456) );
  AOI22X1 U203 ( .A0(N117), .A1(n245), .B0(N214), .B1(n249), .Y(n227) );
  AOI22X1 U204 ( .A0(N356), .A1(n248), .B0(n170), .B1(in_17bit_b[9]), .Y(n228)
         );
  NAND2X1 U205 ( .A(n231), .B(n230), .Y(N457) );
  AOI22X1 U206 ( .A0(N118), .A1(n245), .B0(N215), .B1(n249), .Y(n230) );
  AOI22X1 U207 ( .A0(N357), .A1(n248), .B0(n170), .B1(in_17bit_b[10]), .Y(n231) );
  NAND2X1 U208 ( .A(n234), .B(n233), .Y(N458) );
  AOI22X1 U209 ( .A0(N119), .A1(n245), .B0(N216), .B1(n249), .Y(n233) );
  AOI22X1 U210 ( .A0(N358), .A1(n248), .B0(n170), .B1(in_17bit_b[11]), .Y(n234) );
  NAND2X1 U211 ( .A(n237), .B(n236), .Y(N459) );
  AOI22X1 U212 ( .A0(N120), .A1(n245), .B0(N217), .B1(n249), .Y(n236) );
  AOI22X1 U213 ( .A0(N359), .A1(n248), .B0(n170), .B1(in_17bit_b[12]), .Y(n237) );
  NAND2X1 U214 ( .A(n240), .B(n239), .Y(N460) );
  AOI22X1 U215 ( .A0(N121), .A1(n245), .B0(N218), .B1(n249), .Y(n239) );
  AOI22X1 U216 ( .A0(N360), .A1(n248), .B0(n170), .B1(in_17bit_b[13]), .Y(n240) );
  NAND2X1 U217 ( .A(n243), .B(n242), .Y(N461) );
  AOI22X1 U218 ( .A0(N122), .A1(n245), .B0(N219), .B1(n249), .Y(n242) );
  AOI22X1 U219 ( .A0(N361), .A1(n248), .B0(n170), .B1(in_17bit_b[14]), .Y(n243) );
  NAND2X1 U220 ( .A(n247), .B(n246), .Y(N462) );
  AOI22X1 U221 ( .A0(N123), .A1(n245), .B0(N220), .B1(n249), .Y(n246) );
  AOI22X1 U222 ( .A0(N362), .A1(n248), .B0(n170), .B1(in_17bit_b[15]), .Y(n247) );
  MXI2XL U223 ( .A(n10), .B(n24), .S0(n78), .Y(out[16]) );
  NAND4BBX1 U224 ( .AN(n248), .BN(n249), .C(n198), .D(n251), .Y(N446) );
  NAND4XL U225 ( .A(in_8bit[1]), .B(n44), .C(n191), .D(n171), .Y(n192) );
  NOR2X1 U226 ( .A(in_8bit[6]), .B(in_8bit[4]), .Y(n191) );
  NOR4BX1 U227 ( .AN(n195), .B(n171), .C(in_8bit[1]), .D(in_8bit[2]), .Y(n196)
         );
  NOR2X1 U228 ( .A(in_8bit[6]), .B(in_8bit[3]), .Y(n195) );
  AOI22XL U229 ( .A0(in_17bit[0]), .A1(n54), .B0(in_17bit[0]), .B1(n53), .Y(
        n199) );
  NAND4BXL U230 ( .AN(n44), .B(in_8bit[6]), .C(in_8bit[1]), .D(in_8bit[4]), 
        .Y(n89) );
  INVX1 U231 ( .A(n57), .Y(n69) );
  NAND2BX1 U232 ( .AN(n61), .B(n7), .Y(n57) );
  AOI22XL U233 ( .A0(N27), .A1(n54), .B0(in_17bit[14]), .B1(n55), .Y(n241) );
  AOI22XL U234 ( .A0(N28), .A1(n54), .B0(in_17bit[15]), .B1(n55), .Y(n244) );
  AOI22XL U235 ( .A0(N21), .A1(n54), .B0(in_17bit[8]), .B1(n55), .Y(n223) );
  AOI22XL U236 ( .A0(N22), .A1(n54), .B0(in_17bit[9]), .B1(n53), .Y(n226) );
  AOI22XL U237 ( .A0(N24), .A1(n54), .B0(in_17bit[11]), .B1(n55), .Y(n232) );
  AOI22XL U238 ( .A0(N25), .A1(n54), .B0(in_17bit[12]), .B1(n53), .Y(n235) );
  AOI22XL U239 ( .A0(N26), .A1(n54), .B0(in_17bit[13]), .B1(n55), .Y(n238) );
  AOI22XL U240 ( .A0(N14), .A1(n54), .B0(in_17bit[1]), .B1(n55), .Y(n202) );
  AOI22XL U241 ( .A0(N15), .A1(n54), .B0(in_17bit[2]), .B1(n55), .Y(n205) );
  AOI22XL U242 ( .A0(N16), .A1(n54), .B0(in_17bit[3]), .B1(n53), .Y(n208) );
  AOI22XL U243 ( .A0(N17), .A1(n54), .B0(in_17bit[4]), .B1(n53), .Y(n211) );
  AOI22XL U244 ( .A0(N18), .A1(n54), .B0(in_17bit[5]), .B1(n55), .Y(n214) );
  AOI22XL U245 ( .A0(N19), .A1(n54), .B0(in_17bit[6]), .B1(n53), .Y(n217) );
  AOI22XL U246 ( .A0(N20), .A1(n54), .B0(in_17bit[7]), .B1(n53), .Y(n220) );
  AOI22XL U247 ( .A0(N23), .A1(n54), .B0(in_17bit[10]), .B1(n53), .Y(n229) );
  INVXL U248 ( .A(in_8bit[0]), .Y(n171) );
  AND2X2 U249 ( .A(n69), .B(n9), .Y(n32) );
  AND2X2 U250 ( .A(n32), .B(n13), .Y(n33) );
  AND2X2 U251 ( .A(n33), .B(n14), .Y(n34) );
  AND2X2 U252 ( .A(n34), .B(n15), .Y(n35) );
  AND2X2 U253 ( .A(n35), .B(n12), .Y(n36) );
  AND2X2 U254 ( .A(n36), .B(n16), .Y(n37) );
  OR2XL U255 ( .A(n89), .B(in_8bit[0]), .Y(n85) );
  OAI2BB1X1 U256 ( .A0N(n82), .A1N(n81), .B0(n80), .Y(n245) );
  NOR2BX1 U257 ( .AN(n197), .B(n51), .Y(n82) );
  NOR2BX1 U258 ( .AN(in_8bit[1]), .B(n88), .Y(n81) );
  NAND2X1 U259 ( .A(n40), .B(n8), .Y(n61) );
  AND2X2 U260 ( .A(n37), .B(n17), .Y(n38) );
  INVX1 U261 ( .A(in_17bit[3]), .Y(n95) );
  INVX1 U262 ( .A(in_17bit[4]), .Y(n96) );
  INVX1 U263 ( .A(in_17bit[5]), .Y(n97) );
  INVX1 U264 ( .A(in_17bit[6]), .Y(n98) );
  INVX1 U265 ( .A(in_17bit[7]), .Y(n99) );
  INVX1 U266 ( .A(in_17bit[8]), .Y(n100) );
  INVX1 U267 ( .A(in_17bit[9]), .Y(n101) );
  INVX1 U268 ( .A(in_17bit[10]), .Y(n158) );
  INVX1 U269 ( .A(in_17bit[11]), .Y(n160) );
  INVX1 U270 ( .A(in_17bit[12]), .Y(n161) );
  INVX1 U271 ( .A(in_17bit[13]), .Y(n162) );
  INVX1 U272 ( .A(in_17bit[14]), .Y(n163) );
  INVX1 U273 ( .A(in_17bit[15]), .Y(n164) );
  INVX1 U274 ( .A(in_17bit[1]), .Y(n93) );
  INVX1 U275 ( .A(in_17bit[2]), .Y(n94) );
  INVX1 U276 ( .A(in_17bit[0]), .Y(n92) );
  INVX1 U277 ( .A(n64), .Y(n62) );
  XNOR2X1 U278 ( .A(n23), .B(sub_add_75_b0_carry[12]), .Y(n39) );
  MX2X1 U279 ( .A(neg_mul[22]), .B(N480), .S0(n78), .Y(out[15]) );
  NOR2X1 U280 ( .A(out[0]), .B(neg_mul[8]), .Y(n40) );
  NAND2X1 U281 ( .A(neg_mul[10]), .B(n61), .Y(n64) );
  NAND2X1 U282 ( .A(sub_add_75_b0_carry[15]), .B(n19), .Y(n41) );
  NOR2X4 U283 ( .A(n59), .B(n20), .Y(n58) );
  XOR2X4 U284 ( .A(n58), .B(neg_mul[8]), .Y(out[1]) );
  XNOR2X4 U285 ( .A(n71), .B(n13), .Y(out[5]) );
  XNOR2X4 U286 ( .A(n76), .B(n17), .Y(out[10]) );
  MXI2X4 U287 ( .A(n23), .B(n39), .S0(n78), .Y(out[12]) );
  AND2X1 U288 ( .A(add_1_root_r112_carry_20_), .B(in_17bit_b[16]), .Y(
        add_1_root_r112_SUM_21_) );
  XOR2X1 U289 ( .A(in_17bit_b[16]), .B(add_1_root_r112_carry_20_), .Y(
        add_1_root_r112_SUM_20_) );
  AND2X1 U290 ( .A(add_1_root_r112_carry_19_), .B(in_17bit_b[15]), .Y(
        add_1_root_r112_carry_20_) );
  XOR2X1 U291 ( .A(in_17bit_b[15]), .B(add_1_root_r112_carry_19_), .Y(
        add_1_root_r112_SUM_19_) );
  AND2X1 U292 ( .A(add_1_root_r112_carry_18_), .B(in_17bit_b[14]), .Y(
        add_1_root_r112_carry_19_) );
  XOR2X1 U293 ( .A(in_17bit_b[14]), .B(add_1_root_r112_carry_18_), .Y(
        add_1_root_r112_SUM_18_) );
  AND2X1 U294 ( .A(add_1_root_r112_carry_17_), .B(in_17bit_b[13]), .Y(
        add_1_root_r112_carry_18_) );
  XOR2X1 U295 ( .A(in_17bit_b[13]), .B(add_1_root_r112_carry_17_), .Y(
        add_1_root_r112_SUM_17_) );
  AND2X1 U296 ( .A(add_2_root_r119_carry_21_), .B(in_17bit_b[16]), .Y(
        add_2_root_r119_SUM_22_) );
  XOR2X1 U297 ( .A(in_17bit_b[16]), .B(add_2_root_r119_carry_21_), .Y(
        add_2_root_r119_SUM_21_) );
  AND2X1 U298 ( .A(in_17bit_b[1]), .B(in_17bit_b[0]), .Y(
        add_2_root_r119_carry_6_) );
  AND2X1 U299 ( .A(add_1_root_r119_carry[22]), .B(in_17bit_b[16]), .Y(
        add_1_root_r119_SUM_23_) );
  XOR2X1 U300 ( .A(in_17bit_b[16]), .B(add_1_root_r119_carry[22]), .Y(
        add_1_root_r119_SUM_22_) );
  AND2X1 U301 ( .A(add_1_root_r119_carry[21]), .B(in_17bit_b[15]), .Y(
        add_1_root_r119_carry[22]) );
  XOR2X1 U302 ( .A(in_17bit_b[15]), .B(add_1_root_r119_carry[21]), .Y(
        add_1_root_r119_SUM_21_) );
  AND2X1 U303 ( .A(add_1_root_r119_carry[20]), .B(in_17bit_b[14]), .Y(
        add_1_root_r119_carry[21]) );
  XOR2X1 U304 ( .A(in_17bit_b[14]), .B(add_1_root_r119_carry[20]), .Y(
        add_1_root_r119_SUM_20_) );
  AND2X1 U305 ( .A(add_1_root_r119_A_6_), .B(in_17bit_b[0]), .Y(
        add_1_root_r119_carry[7]) );
  XOR2X1 U306 ( .A(in_17bit_b[0]), .B(add_1_root_r119_A_6_), .Y(
        add_1_root_r119_SUM_6_) );
  AND2X1 U307 ( .A(add_3_root_r119_carry_18_), .B(in_17bit_b[16]), .Y(
        add_1_root_r119_A_19_) );
  XOR2X1 U308 ( .A(in_17bit_b[16]), .B(add_3_root_r119_carry_18_), .Y(
        add_1_root_r119_A_18_) );
  XOR2X1 U309 ( .A(in_17bit_b[0]), .B(in_17bit_b[1]), .Y(add_1_root_r119_A_2_)
         );
  AND2X1 U310 ( .A(add_2_root_r115_carry_19_), .B(in_17bit_b[16]), .Y(
        add_2_root_r115_SUM_20_) );
  XOR2X1 U311 ( .A(in_17bit_b[16]), .B(add_2_root_r115_carry_19_), .Y(
        add_2_root_r115_SUM_19_) );
  AND2X1 U312 ( .A(add_2_root_r115_carry_18_), .B(in_17bit_b[15]), .Y(
        add_2_root_r115_carry_19_) );
  XOR2X1 U313 ( .A(in_17bit_b[15]), .B(add_2_root_r115_carry_18_), .Y(
        add_2_root_r115_SUM_18_) );
  AND2X1 U314 ( .A(in_17bit_b[2]), .B(in_17bit_b[0]), .Y(
        add_2_root_r115_carry_4_) );
  AND2X1 U315 ( .A(add_1_root_r115_carry_22_), .B(in_17bit_b[16]), .Y(
        add_1_root_r115_SUM_23_) );
  XOR2X1 U316 ( .A(in_17bit_b[16]), .B(add_1_root_r115_carry_22_), .Y(
        add_1_root_r115_SUM_22_) );
  AND2X1 U317 ( .A(add_1_root_r115_carry_21_), .B(in_17bit_b[15]), .Y(
        add_1_root_r115_carry_22_) );
  XOR2X1 U318 ( .A(in_17bit_b[15]), .B(add_1_root_r115_carry_21_), .Y(
        add_1_root_r115_SUM_21_) );
  XOR2X1 U319 ( .A(in_17bit_b[0]), .B(in_17bit_b[2]), .Y(
        add_1_root_r115_SUM_6_) );
  XOR2X1 U320 ( .A(n56), .B(sub_add_54_b0_carry[16]), .Y(N29) );
  AND2X1 U321 ( .A(sub_add_54_b0_carry[15]), .B(n164), .Y(
        sub_add_54_b0_carry[16]) );
  XOR2X1 U322 ( .A(n164), .B(sub_add_54_b0_carry[15]), .Y(N28) );
  AND2X1 U323 ( .A(sub_add_54_b0_carry[14]), .B(n163), .Y(
        sub_add_54_b0_carry[15]) );
  XOR2X1 U324 ( .A(n163), .B(sub_add_54_b0_carry[14]), .Y(N27) );
  AND2X1 U325 ( .A(sub_add_54_b0_carry[13]), .B(n162), .Y(
        sub_add_54_b0_carry[14]) );
  XOR2X1 U326 ( .A(n162), .B(sub_add_54_b0_carry[13]), .Y(N26) );
  AND2X1 U327 ( .A(sub_add_54_b0_carry[12]), .B(n161), .Y(
        sub_add_54_b0_carry[13]) );
  XOR2X1 U328 ( .A(n161), .B(sub_add_54_b0_carry[12]), .Y(N25) );
  AND2X1 U329 ( .A(sub_add_54_b0_carry[11]), .B(n160), .Y(
        sub_add_54_b0_carry[12]) );
  XOR2X1 U330 ( .A(n160), .B(sub_add_54_b0_carry[11]), .Y(N24) );
  AND2X1 U331 ( .A(sub_add_54_b0_carry[10]), .B(n158), .Y(
        sub_add_54_b0_carry[11]) );
  XOR2X1 U332 ( .A(n158), .B(sub_add_54_b0_carry[10]), .Y(N23) );
  AND2X1 U333 ( .A(sub_add_54_b0_carry[9]), .B(n101), .Y(
        sub_add_54_b0_carry[10]) );
  XOR2X1 U334 ( .A(n101), .B(sub_add_54_b0_carry[9]), .Y(N22) );
  AND2X1 U335 ( .A(sub_add_54_b0_carry[8]), .B(n100), .Y(
        sub_add_54_b0_carry[9]) );
  XOR2X1 U336 ( .A(n100), .B(sub_add_54_b0_carry[8]), .Y(N21) );
  AND2X1 U337 ( .A(sub_add_54_b0_carry[7]), .B(n99), .Y(sub_add_54_b0_carry[8]) );
  XOR2X1 U338 ( .A(n99), .B(sub_add_54_b0_carry[7]), .Y(N20) );
  AND2X1 U339 ( .A(sub_add_54_b0_carry[6]), .B(n98), .Y(sub_add_54_b0_carry[7]) );
  XOR2X1 U340 ( .A(n98), .B(sub_add_54_b0_carry[6]), .Y(N19) );
  AND2X1 U341 ( .A(sub_add_54_b0_carry[5]), .B(n97), .Y(sub_add_54_b0_carry[6]) );
  XOR2X1 U342 ( .A(n97), .B(sub_add_54_b0_carry[5]), .Y(N18) );
  AND2X1 U343 ( .A(sub_add_54_b0_carry[4]), .B(n96), .Y(sub_add_54_b0_carry[5]) );
  XOR2X1 U344 ( .A(n96), .B(sub_add_54_b0_carry[4]), .Y(N17) );
  AND2X1 U345 ( .A(sub_add_54_b0_carry[3]), .B(n95), .Y(sub_add_54_b0_carry[4]) );
  XOR2X1 U346 ( .A(n95), .B(sub_add_54_b0_carry[3]), .Y(N16) );
  AND2X1 U347 ( .A(sub_add_54_b0_carry[2]), .B(n94), .Y(sub_add_54_b0_carry[3]) );
  XOR2X1 U348 ( .A(n94), .B(sub_add_54_b0_carry[2]), .Y(N15) );
  AND2X1 U349 ( .A(n92), .B(n93), .Y(sub_add_54_b0_carry[2]) );
  XOR2X1 U350 ( .A(n93), .B(n92), .Y(N14) );
  XOR2X1 U351 ( .A(n19), .B(sub_add_75_b0_carry[15]), .Y(N480) );
  AND2X1 U352 ( .A(sub_add_75_b0_carry[14]), .B(n21), .Y(
        sub_add_75_b0_carry[15]) );
  XOR2X1 U353 ( .A(n21), .B(sub_add_75_b0_carry[14]), .Y(N479) );
  AND2X1 U354 ( .A(sub_add_75_b0_carry[13]), .B(n22), .Y(
        sub_add_75_b0_carry[14]) );
  XOR2X1 U355 ( .A(n22), .B(sub_add_75_b0_carry[13]), .Y(N478) );
  AND2X1 U356 ( .A(sub_add_75_b0_carry[12]), .B(n23), .Y(
        sub_add_75_b0_carry[13]) );
  AND2X1 U357 ( .A(n38), .B(n18), .Y(sub_add_75_b0_carry[12]) );
  AND2X1 U358 ( .A(in_17bit_b[0]), .B(in_17bit_b[4]), .Y(
        add_1_root_r112_carry_5_) );
endmodule


module multi16_4_DW01_add_0 ( A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, 
        A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, 
        A_4_, B_23_, B_22_, B_21_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, 
        B_14_, B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, 
        SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, 
        SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, 
        SUM_7_ );
  input A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_,
         A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, B_23_, B_22_,
         B_21_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_,
         B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_;
  output SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_,
         SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_,
         SUM_8_, SUM_7_;
  wire   n1, n2, n3, n4;
  wire   [23:7] carry;

  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry[7]), .CO(carry[8]), .S(SUM_7_)
         );
  ADDFX2 U1_21 ( .A(A_21_), .B(B_21_), .CI(carry[21]), .CO(carry[22]), .S(
        SUM_21_) );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry[20]), .CO(carry[21]), .S(
        SUM_20_) );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry[19]), .CO(carry[20]), .S(
        SUM_19_) );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry[18]), .CO(carry[19]), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry[17]), .CO(carry[18]), .S(
        SUM_17_) );
  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry[16]), .CO(carry[17]), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry[15]), .CO(carry[16]), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry[14]), .CO(carry[15]), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry[13]), .CO(carry[14]), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry[12]), .CO(carry[13]), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry[11]), .CO(carry[12]), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry[10]), .CO(carry[11]), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry[9]), .CO(carry[10]), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry[8]), .CO(carry[9]), .S(SUM_8_)
         );
  ADDFX2 U1_22 ( .A(A_22_), .B(B_22_), .CI(carry[22]), .CO(carry[23]), .S(
        SUM_22_) );
  AND2X2 U1 ( .A(A_4_), .B(B_4_), .Y(n1) );
  XOR2X1 U2 ( .A(B_23_), .B(carry[23]), .Y(SUM_23_) );
  OAI2BB1X1 U3 ( .A0N(n2), .A1N(A_6_), .B0(n3), .Y(carry[7]) );
  OAI21XL U4 ( .A0(A_6_), .A1(n2), .B0(B_6_), .Y(n3) );
  OAI2BB1X1 U5 ( .A0N(n1), .A1N(A_5_), .B0(n4), .Y(n2) );
  OAI21XL U6 ( .A0(A_5_), .A1(n1), .B0(B_5_), .Y(n4) );
endmodule


module multi16_4_DW01_add_4 ( A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, 
        A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, 
        B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, 
        B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, SUM_22_, SUM_21_, SUM_20_, 
        SUM_19_, SUM_18_, SUM_17_, SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, 
        SUM_11_, SUM_10_, SUM_9_, SUM_8_, SUM_7_ );
  input A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_,
         A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, B_20_, B_19_,
         B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, B_10_, B_9_,
         B_8_, B_7_, B_6_, B_5_;
  output SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_,
         SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_,
         SUM_7_;
  wire   carry_21_, carry_20_, carry_19_, carry_18_, carry_17_, carry_16_,
         carry_15_, carry_14_, carry_13_, carry_12_, carry_11_, carry_10_,
         carry_9_, carry_8_, carry_7_, n1;

  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry_16_), .CO(carry_17_), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry_15_), .CO(carry_16_), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry_14_), .CO(carry_15_), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry_13_), .CO(carry_14_), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry_12_), .CO(carry_13_), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry_11_), .CO(carry_12_), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry_10_), .CO(carry_11_), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry_9_), .CO(carry_10_), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry_8_), .CO(carry_9_), .S(SUM_8_)
         );
  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry_7_), .CO(carry_8_), .S(SUM_7_)
         );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry_20_), .CO(carry_21_), .S(
        SUM_20_) );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry_19_), .CO(carry_20_), .S(
        SUM_19_) );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry_18_), .CO(carry_19_), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry_17_), .CO(carry_18_), .S(
        SUM_17_) );
  ADDFX2 U1_21 ( .A(A_21_), .B(B_21_), .CI(carry_21_), .CO(SUM_22_), .S(
        SUM_21_) );
  OAI2BB1X1 U1 ( .A0N(A_6_), .A1N(B_6_), .B0(n1), .Y(carry_7_) );
  OAI211X1 U2 ( .A0(B_6_), .A1(A_6_), .B0(A_5_), .C0(B_5_), .Y(n1) );
endmodule


module multi16_4_DW01_add_6 ( A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, 
        A_16_, A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, 
        A_6_, A_5_, A_4_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, 
        B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, 
        SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, 
        SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, 
        SUM_7_ );
  input A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_,
         A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, B_20_,
         B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, B_10_,
         B_9_, B_8_, B_7_, B_6_, B_5_, B_4_;
  output SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_,
         SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_,
         SUM_8_, SUM_7_;
  wire   n1, n2, n3, n4, n5, n6;
  wire   [21:7] carry;

  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry[7]), .CO(carry[8]), .S(SUM_7_)
         );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry[18]), .CO(carry[19]), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry[17]), .CO(carry[18]), .S(
        SUM_17_) );
  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry[16]), .CO(carry[17]), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry[15]), .CO(carry[16]), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry[14]), .CO(carry[15]), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry[13]), .CO(carry[14]), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry[12]), .CO(carry[13]), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry[11]), .CO(carry[12]), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry[10]), .CO(carry[11]), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry[9]), .CO(carry[10]), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry[8]), .CO(carry[9]), .S(SUM_8_)
         );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry[19]), .CO(carry[20]), .S(
        SUM_19_) );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry[20]), .CO(carry[21]), .S(
        SUM_20_) );
  AND2X2 U1 ( .A(A_22_), .B(n2), .Y(n1) );
  AND2X2 U2 ( .A(A_21_), .B(carry[21]), .Y(n2) );
  XOR2X1 U3 ( .A(A_23_), .B(n1), .Y(SUM_23_) );
  XOR2X1 U4 ( .A(A_21_), .B(carry[21]), .Y(SUM_21_) );
  XOR2X1 U5 ( .A(A_22_), .B(n2), .Y(SUM_22_) );
  AND2X2 U6 ( .A(A_4_), .B(B_4_), .Y(n3) );
  OAI2BB1X1 U7 ( .A0N(n4), .A1N(A_6_), .B0(n5), .Y(carry[7]) );
  OAI21XL U8 ( .A0(A_6_), .A1(n4), .B0(B_6_), .Y(n5) );
  OAI2BB1X1 U9 ( .A0N(n3), .A1N(A_5_), .B0(n6), .Y(n4) );
  OAI21XL U10 ( .A0(A_5_), .A1(n3), .B0(B_5_), .Y(n6) );
endmodule


module multi16_4 ( in_17bit, in_8bit, out );
  input [16:0] in_17bit;
  input [7:0] in_8bit;
  output [16:0] out;
  wire   n295, n296, n297, n298, n299, N14, N15, N16, N17, N18, N19, N20, N21,
         N22, N23, N24, N25, N26, N27, N28, N29, N108, N109, N110, N111, N112,
         N113, N114, N115, N116, N117, N118, N119, N120, N121, N122, N123,
         N205, N206, N207, N208, N209, N210, N211, N212, N213, N214, N215,
         N216, N217, N218, N219, N220, N221, N347, N348, N349, N350, N351,
         N352, N353, N354, N355, N356, N357, N358, N359, N360, N361, N362,
         N363, N446, N447, N448, N449, N450, N451, N452, N453, N454, N455,
         N456, N457, N458, N459, N460, N461, N462, N463, N479, N480, N481,
         add_2_root_r119_carry_10_, add_2_root_r119_carry_11_,
         add_2_root_r119_carry_12_, add_2_root_r119_carry_13_,
         add_2_root_r119_carry_14_, add_2_root_r119_carry_15_,
         add_2_root_r119_carry_16_, add_2_root_r119_carry_17_,
         add_2_root_r119_carry_18_, add_2_root_r119_carry_19_,
         add_2_root_r119_carry_20_, add_2_root_r119_carry_21_,
         add_2_root_r119_carry_7_, add_2_root_r119_carry_8_,
         add_2_root_r119_carry_9_, add_2_root_r119_SUM_6_,
         add_2_root_r119_SUM_7_, add_2_root_r119_SUM_8_,
         add_2_root_r119_SUM_9_, add_2_root_r119_SUM_10_,
         add_2_root_r119_SUM_11_, add_2_root_r119_SUM_12_,
         add_2_root_r119_SUM_13_, add_2_root_r119_SUM_14_,
         add_2_root_r119_SUM_15_, add_2_root_r119_SUM_16_,
         add_2_root_r119_SUM_17_, add_2_root_r119_SUM_18_,
         add_2_root_r119_SUM_19_, add_2_root_r119_SUM_20_,
         add_2_root_r119_SUM_21_, add_2_root_r119_SUM_22_,
         add_1_root_r119_SUM_6_, add_1_root_r119_SUM_7_,
         add_1_root_r119_SUM_8_, add_1_root_r119_SUM_9_,
         add_1_root_r119_SUM_10_, add_1_root_r119_SUM_11_,
         add_1_root_r119_SUM_12_, add_1_root_r119_SUM_13_,
         add_1_root_r119_SUM_14_, add_1_root_r119_SUM_15_,
         add_1_root_r119_SUM_16_, add_1_root_r119_SUM_17_,
         add_1_root_r119_SUM_18_, add_1_root_r119_SUM_19_,
         add_1_root_r119_SUM_20_, add_1_root_r119_SUM_21_,
         add_1_root_r119_SUM_22_, add_1_root_r119_SUM_23_,
         add_1_root_r119_A_2_, add_1_root_r119_A_3_, add_1_root_r119_A_4_,
         add_1_root_r119_A_5_, add_1_root_r119_A_6_, add_1_root_r119_A_7_,
         add_1_root_r119_A_8_, add_1_root_r119_A_9_, add_1_root_r119_A_10_,
         add_1_root_r119_A_11_, add_1_root_r119_A_12_, add_1_root_r119_A_13_,
         add_1_root_r119_A_14_, add_1_root_r119_A_15_, add_1_root_r119_A_16_,
         add_1_root_r119_A_17_, add_1_root_r119_A_18_, add_1_root_r119_A_19_,
         add_3_root_r119_carry_10_, add_3_root_r119_carry_11_,
         add_3_root_r119_carry_12_, add_3_root_r119_carry_13_,
         add_3_root_r119_carry_14_, add_3_root_r119_carry_15_,
         add_3_root_r119_carry_16_, add_3_root_r119_carry_17_,
         add_3_root_r119_carry_18_, add_3_root_r119_carry_3_,
         add_3_root_r119_carry_4_, add_3_root_r119_carry_5_,
         add_3_root_r119_carry_6_, add_3_root_r119_carry_7_,
         add_3_root_r119_carry_8_, add_3_root_r119_carry_9_,
         add_1_root_r112_carry_10_, add_1_root_r112_carry_11_,
         add_1_root_r112_carry_12_, add_1_root_r112_carry_13_,
         add_1_root_r112_carry_14_, add_1_root_r112_carry_15_,
         add_1_root_r112_carry_16_, add_1_root_r112_carry_17_,
         add_1_root_r112_carry_18_, add_1_root_r112_carry_19_,
         add_1_root_r112_carry_20_, add_1_root_r112_carry_5_,
         add_1_root_r112_carry_6_, add_1_root_r112_carry_7_,
         add_1_root_r112_carry_8_, add_1_root_r112_carry_9_,
         add_1_root_r112_SUM_1_, add_1_root_r112_SUM_2_,
         add_1_root_r112_SUM_3_, add_1_root_r112_SUM_4_,
         add_1_root_r112_SUM_5_, add_1_root_r112_SUM_6_,
         add_1_root_r112_SUM_7_, add_1_root_r112_SUM_8_,
         add_1_root_r112_SUM_9_, add_1_root_r112_SUM_10_,
         add_1_root_r112_SUM_11_, add_1_root_r112_SUM_12_,
         add_1_root_r112_SUM_13_, add_1_root_r112_SUM_14_,
         add_1_root_r112_SUM_15_, add_1_root_r112_SUM_16_,
         add_1_root_r112_SUM_17_, add_1_root_r112_SUM_18_,
         add_1_root_r112_SUM_19_, add_1_root_r112_SUM_20_,
         add_1_root_r112_SUM_21_, add_2_root_r115_carry_10_,
         add_2_root_r115_carry_11_, add_2_root_r115_carry_12_,
         add_2_root_r115_carry_13_, add_2_root_r115_carry_14_,
         add_2_root_r115_carry_15_, add_2_root_r115_carry_16_,
         add_2_root_r115_carry_17_, add_2_root_r115_carry_18_,
         add_2_root_r115_carry_19_, add_2_root_r115_carry_5_,
         add_2_root_r115_carry_6_, add_2_root_r115_carry_7_,
         add_2_root_r115_carry_8_, add_2_root_r115_carry_9_,
         add_2_root_r115_SUM_4_, add_2_root_r115_SUM_5_,
         add_2_root_r115_SUM_6_, add_2_root_r115_SUM_7_,
         add_2_root_r115_SUM_8_, add_2_root_r115_SUM_9_,
         add_2_root_r115_SUM_10_, add_2_root_r115_SUM_11_,
         add_2_root_r115_SUM_12_, add_2_root_r115_SUM_13_,
         add_2_root_r115_SUM_14_, add_2_root_r115_SUM_15_,
         add_2_root_r115_SUM_16_, add_2_root_r115_SUM_17_,
         add_2_root_r115_SUM_18_, add_2_root_r115_SUM_19_,
         add_2_root_r115_SUM_20_, add_1_root_r115_carry_10_,
         add_1_root_r115_carry_11_, add_1_root_r115_carry_12_,
         add_1_root_r115_carry_13_, add_1_root_r115_carry_14_,
         add_1_root_r115_carry_15_, add_1_root_r115_carry_16_,
         add_1_root_r115_carry_17_, add_1_root_r115_carry_18_,
         add_1_root_r115_carry_19_, add_1_root_r115_carry_20_,
         add_1_root_r115_carry_21_, add_1_root_r115_carry_22_,
         add_1_root_r115_carry_7_, add_1_root_r115_carry_8_,
         add_1_root_r115_carry_9_, add_1_root_r115_SUM_6_,
         add_1_root_r115_SUM_7_, add_1_root_r115_SUM_8_,
         add_1_root_r115_SUM_9_, add_1_root_r115_SUM_10_,
         add_1_root_r115_SUM_11_, add_1_root_r115_SUM_12_,
         add_1_root_r115_SUM_13_, add_1_root_r115_SUM_14_,
         add_1_root_r115_SUM_15_, add_1_root_r115_SUM_16_,
         add_1_root_r115_SUM_17_, add_1_root_r115_SUM_18_,
         add_1_root_r115_SUM_19_, add_1_root_r115_SUM_20_,
         add_1_root_r115_SUM_21_, add_1_root_r115_SUM_22_,
         add_1_root_r115_SUM_23_, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n22, n23, n26, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n158, n160, n161, n162, n163, n164, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294;
  wire   [16:0] in_17bit_b;
  wire   [23:8] neg_mul;
  wire   [16:13] sub_add_75_b0_carry;
  wire   [15:2] sub_add_54_b0_carry;
  wire   [22:7] add_1_root_r119_carry;

  multi16_4_DW01_add_0 add_0_root_r119 ( .A_22_(add_2_root_r119_SUM_22_), 
        .A_21_(add_2_root_r119_SUM_21_), .A_20_(add_2_root_r119_SUM_20_), 
        .A_19_(add_2_root_r119_SUM_19_), .A_18_(add_2_root_r119_SUM_18_), 
        .A_17_(add_2_root_r119_SUM_17_), .A_16_(add_2_root_r119_SUM_16_), 
        .A_15_(add_2_root_r119_SUM_15_), .A_14_(add_2_root_r119_SUM_14_), 
        .A_13_(add_2_root_r119_SUM_13_), .A_12_(add_2_root_r119_SUM_12_), 
        .A_11_(add_2_root_r119_SUM_11_), .A_10_(add_2_root_r119_SUM_10_), 
        .A_9_(add_2_root_r119_SUM_9_), .A_8_(add_2_root_r119_SUM_8_), .A_7_(
        add_2_root_r119_SUM_7_), .A_6_(add_2_root_r119_SUM_6_), .A_5_(
        add_1_root_r119_A_2_), .A_4_(in_17bit_b[0]), .B_23_(
        add_1_root_r119_SUM_23_), .B_22_(add_1_root_r119_SUM_22_), .B_21_(
        add_1_root_r119_SUM_21_), .B_20_(add_1_root_r119_SUM_20_), .B_19_(
        add_1_root_r119_SUM_19_), .B_18_(add_1_root_r119_SUM_18_), .B_17_(
        add_1_root_r119_SUM_17_), .B_16_(add_1_root_r119_SUM_16_), .B_15_(
        add_1_root_r119_SUM_15_), .B_14_(add_1_root_r119_SUM_14_), .B_13_(
        add_1_root_r119_SUM_13_), .B_12_(add_1_root_r119_SUM_12_), .B_11_(
        add_1_root_r119_SUM_11_), .B_10_(add_1_root_r119_SUM_10_), .B_9_(
        add_1_root_r119_SUM_9_), .B_8_(add_1_root_r119_SUM_8_), .B_7_(
        add_1_root_r119_SUM_7_), .B_6_(add_1_root_r119_SUM_6_), .B_5_(
        add_1_root_r119_A_5_), .B_4_(add_1_root_r119_A_4_), .SUM_23_(N363), 
        .SUM_22_(N362), .SUM_21_(N361), .SUM_20_(N360), .SUM_19_(N359), 
        .SUM_18_(N358), .SUM_17_(N357), .SUM_16_(N356), .SUM_15_(N355), 
        .SUM_14_(N354), .SUM_13_(N353), .SUM_12_(N352), .SUM_11_(N351), 
        .SUM_10_(N350), .SUM_9_(N349), .SUM_8_(N348), .SUM_7_(N347) );
  multi16_4_DW01_add_4 add_0_root_r112 ( .A_21_(in_17bit_b[16]), .A_20_(
        in_17bit_b[15]), .A_19_(in_17bit_b[14]), .A_18_(in_17bit_b[13]), 
        .A_17_(in_17bit_b[12]), .A_16_(in_17bit_b[11]), .A_15_(in_17bit_b[10]), 
        .A_14_(in_17bit_b[9]), .A_13_(in_17bit_b[8]), .A_12_(in_17bit_b[7]), 
        .A_11_(in_17bit_b[6]), .A_10_(in_17bit_b[5]), .A_9_(in_17bit_b[4]), 
        .A_8_(in_17bit_b[3]), .A_7_(in_17bit_b[2]), .A_6_(in_17bit_b[1]), 
        .A_5_(in_17bit_b[0]), .B_21_(add_1_root_r112_SUM_21_), .B_20_(
        add_1_root_r112_SUM_20_), .B_19_(add_1_root_r112_SUM_19_), .B_18_(
        add_1_root_r112_SUM_18_), .B_17_(add_1_root_r112_SUM_17_), .B_16_(
        add_1_root_r112_SUM_16_), .B_15_(add_1_root_r112_SUM_15_), .B_14_(
        add_1_root_r112_SUM_14_), .B_13_(add_1_root_r112_SUM_13_), .B_12_(
        add_1_root_r112_SUM_12_), .B_11_(add_1_root_r112_SUM_11_), .B_10_(
        add_1_root_r112_SUM_10_), .B_9_(add_1_root_r112_SUM_9_), .B_8_(
        add_1_root_r112_SUM_8_), .B_7_(add_1_root_r112_SUM_7_), .B_6_(
        add_1_root_r112_SUM_6_), .B_5_(add_1_root_r112_SUM_5_), .SUM_22_(N123), 
        .SUM_21_(N122), .SUM_20_(N121), .SUM_19_(N120), .SUM_18_(N119), 
        .SUM_17_(N118), .SUM_16_(N117), .SUM_15_(N116), .SUM_14_(N115), 
        .SUM_13_(N114), .SUM_12_(N113), .SUM_11_(N112), .SUM_10_(N111), 
        .SUM_9_(N110), .SUM_8_(N109), .SUM_7_(N108) );
  multi16_4_DW01_add_6 add_0_root_r115 ( .A_23_(add_1_root_r115_SUM_23_), 
        .A_22_(add_1_root_r115_SUM_22_), .A_21_(add_1_root_r115_SUM_21_), 
        .A_20_(add_1_root_r115_SUM_20_), .A_19_(add_1_root_r115_SUM_19_), 
        .A_18_(add_1_root_r115_SUM_18_), .A_17_(add_1_root_r115_SUM_17_), 
        .A_16_(add_1_root_r115_SUM_16_), .A_15_(add_1_root_r115_SUM_15_), 
        .A_14_(add_1_root_r115_SUM_14_), .A_13_(add_1_root_r115_SUM_13_), 
        .A_12_(add_1_root_r115_SUM_12_), .A_11_(add_1_root_r115_SUM_11_), 
        .A_10_(add_1_root_r115_SUM_10_), .A_9_(add_1_root_r115_SUM_9_), .A_8_(
        add_1_root_r115_SUM_8_), .A_7_(add_1_root_r115_SUM_7_), .A_6_(
        add_1_root_r115_SUM_6_), .A_5_(in_17bit_b[1]), .A_4_(in_17bit_b[0]), 
        .B_20_(add_2_root_r115_SUM_20_), .B_19_(add_2_root_r115_SUM_19_), 
        .B_18_(add_2_root_r115_SUM_18_), .B_17_(add_2_root_r115_SUM_17_), 
        .B_16_(add_2_root_r115_SUM_16_), .B_15_(add_2_root_r115_SUM_15_), 
        .B_14_(add_2_root_r115_SUM_14_), .B_13_(add_2_root_r115_SUM_13_), 
        .B_12_(add_2_root_r115_SUM_12_), .B_11_(add_2_root_r115_SUM_11_), 
        .B_10_(add_2_root_r115_SUM_10_), .B_9_(add_2_root_r115_SUM_9_), .B_8_(
        add_2_root_r115_SUM_8_), .B_7_(add_2_root_r115_SUM_7_), .B_6_(
        add_2_root_r115_SUM_6_), .B_5_(add_2_root_r115_SUM_5_), .B_4_(
        add_2_root_r115_SUM_4_), .SUM_23_(N221), .SUM_22_(N220), .SUM_21_(N219), .SUM_20_(N218), .SUM_19_(N217), .SUM_18_(N216), .SUM_17_(N215), .SUM_16_(
        N214), .SUM_15_(N213), .SUM_14_(N212), .SUM_13_(N211), .SUM_12_(N210), 
        .SUM_11_(N209), .SUM_10_(N208), .SUM_9_(N207), .SUM_8_(N206), .SUM_7_(
        N205) );
  TLATX1 neg_mul_reg_19_ ( .G(N446), .D(N459), .QN(n5) );
  TLATX1 neg_mul_reg_18_ ( .G(N446), .D(N458), .QN(n4) );
  TLATX1 neg_mul_reg_17_ ( .G(N446), .D(N457), .QN(n3) );
  TLATX1 neg_mul_reg_16_ ( .G(N446), .D(N456), .Q(neg_mul[16]), .QN(n18) );
  TLATX1 neg_mul_reg_23_ ( .G(N446), .D(N463), .Q(neg_mul[23]), .QN(n17) );
  TLATX1 neg_mul_reg_22_ ( .G(N446), .D(N462), .Q(neg_mul[22]), .QN(n10) );
  TLATX1 neg_mul_reg_21_ ( .G(N446), .D(N461), .Q(neg_mul[21]), .QN(n9) );
  TLATX1 neg_mul_reg_20_ ( .G(N446), .D(N460), .QN(n16) );
  TLATX1 neg_mul_reg_9_ ( .G(N446), .D(N449), .Q(neg_mul[9]), .QN(n11) );
  TLATX1 neg_mul_reg_15_ ( .G(N446), .D(N455), .Q(neg_mul[15]), .QN(n15) );
  TLATX1 neg_mul_reg_14_ ( .G(N446), .D(N454), .Q(neg_mul[14]), .QN(n14) );
  TLATX1 neg_mul_reg_13_ ( .G(N446), .D(N453), .Q(neg_mul[13]), .QN(n13) );
  TLATX1 neg_mul_reg_12_ ( .G(N446), .D(N452), .Q(neg_mul[12]), .QN(n7) );
  TLATX1 neg_mul_reg_11_ ( .G(N446), .D(N451), .Q(neg_mul[11]), .QN(n12) );
  TLATX1 neg_mul_reg_10_ ( .G(N446), .D(N450), .Q(neg_mul[10]), .QN(n6) );
  TLATX1 neg_mul_reg_8_ ( .G(N446), .D(N448), .Q(neg_mul[8]), .QN(n19) );
  TLATX1 neg_mul_reg_7_ ( .G(N446), .D(N447), .Q(out[0]) );
  NAND2X1 U2 ( .A(n2), .B(n11), .Y(n59) );
  CLKBUFX8 U3 ( .A(n298), .Y(out[2]) );
  BUFX8 U4 ( .A(in_17bit[16]), .Y(n20) );
  CLKINVX3 U5 ( .A(n54), .Y(n51) );
  CLKINVX3 U6 ( .A(n294), .Y(in_17bit_b[16]) );
  NOR2X1 U7 ( .A(n172), .B(n20), .Y(n173) );
  BUFX8 U8 ( .A(n43), .Y(n1) );
  BUFX16 U9 ( .A(n43), .Y(n2) );
  OAI21X1 U10 ( .A0(n42), .A1(n84), .B0(n83), .Y(n89) );
  NAND2XL U11 ( .A(n2), .B(n7), .Y(n83) );
  INVX20 U12 ( .A(n46), .Y(n42) );
  NOR2X2 U13 ( .A(n53), .B(n70), .Y(n72) );
  AOI2BB2X1 U14 ( .B0(n69), .B1(n42), .A0N(n44), .A1N(neg_mul[10]), .Y(n70) );
  NAND2XL U15 ( .A(n1), .B(n6), .Y(n67) );
  AOI2BB2X1 U16 ( .B0(n61), .B1(n42), .A0N(n44), .A1N(neg_mul[9]), .Y(n62) );
  OAI21XL U17 ( .A0(n42), .A1(n68), .B0(n67), .Y(n73) );
  CLKINVX2 U18 ( .A(in_8bit[7]), .Y(n46) );
  MXI2X1 U19 ( .A(n16), .B(n35), .S0(n181), .Y(out[13]) );
  XNOR2X2 U20 ( .A(n179), .B(n5), .Y(out[12]) );
  MX2X2 U21 ( .A(neg_mul[21]), .B(N479), .S0(n181), .Y(out[14]) );
  INVX8 U22 ( .A(n45), .Y(n43) );
  AND2X2 U23 ( .A(out[0]), .B(neg_mul[8]), .Y(n8) );
  CLKINVX3 U24 ( .A(n53), .Y(n22) );
  NOR2X1 U25 ( .A(n94), .B(n52), .Y(n96) );
  CLKINVX8 U26 ( .A(n49), .Y(n53) );
  OAI2BB1X2 U27 ( .A0N(n46), .A1N(n8), .B0(n55), .Y(n58) );
  AOI2BB2X1 U28 ( .B0(n93), .B1(n2), .A0N(n2), .A1N(neg_mul[13]), .Y(n94) );
  BUFX16 U29 ( .A(n296), .Y(out[4]) );
  XNOR2X2 U30 ( .A(n52), .B(n42), .Y(n177) );
  INVX12 U31 ( .A(n180), .Y(n181) );
  NOR2X2 U32 ( .A(n20), .B(n158), .Y(n161) );
  AOI211X2 U33 ( .A0(n20), .A1(n89), .B0(n88), .C0(n87), .Y(out[5]) );
  BUFX8 U34 ( .A(n295), .Y(out[7]) );
  AOI211X2 U35 ( .A0(n23), .A1(n162), .B0(n161), .C0(n160), .Y(n295) );
  AOI211X2 U36 ( .A0(n65), .A1(n20), .B0(n64), .C0(n63), .Y(n298) );
  INVX4 U37 ( .A(n22), .Y(n23) );
  NOR2X2 U38 ( .A(n53), .B(n86), .Y(n88) );
  XOR2X4 U39 ( .A(n175), .B(neg_mul[16]), .Y(out[9]) );
  NOR2X4 U40 ( .A(n52), .B(n56), .Y(n57) );
  INVX8 U41 ( .A(in_17bit[16]), .Y(n49) );
  NOR2X2 U42 ( .A(n53), .B(n78), .Y(n80) );
  INVXL U43 ( .A(n23), .Y(n54) );
  XNOR2X4 U44 ( .A(n53), .B(n42), .Y(n180) );
  INVX8 U45 ( .A(n49), .Y(n52) );
  NOR2X2 U46 ( .A(n20), .B(n62), .Y(n64) );
  CLKINVX8 U47 ( .A(n26), .Y(out[3]) );
  AOI2BB2X2 U48 ( .B0(n8), .B1(n42), .A0N(n44), .A1N(neg_mul[8]), .Y(n56) );
  CLKINVX8 U49 ( .A(n45), .Y(n44) );
  INVX4 U50 ( .A(in_8bit[7]), .Y(n45) );
  INVX4 U51 ( .A(n297), .Y(n26) );
  AOI211X2 U52 ( .A0(n20), .A1(n73), .B0(n72), .C0(n71), .Y(n297) );
  NOR2X4 U53 ( .A(n32), .B(n177), .Y(n176) );
  AOI2BB2XL U54 ( .B0(n85), .B1(n1), .A0N(n44), .A1N(neg_mul[12]), .Y(n86) );
  AOI2BB2XL U55 ( .B0(n171), .B1(n2), .A0N(n44), .A1N(neg_mul[15]), .Y(n172)
         );
  OAI21XL U56 ( .A0(n42), .A1(n60), .B0(n59), .Y(n65) );
  NOR2X2 U57 ( .A(n180), .B(n34), .Y(n179) );
  NOR4XL U58 ( .A(in_8bit[1]), .B(in_8bit[0]), .C(in_8bit[2]), .D(in_8bit[3]), 
        .Y(n29) );
  INVX1 U59 ( .A(n244), .Y(in_17bit_b[1]) );
  INVX1 U60 ( .A(n283), .Y(in_17bit_b[14]) );
  INVX1 U61 ( .A(n280), .Y(in_17bit_b[13]) );
  INVX1 U62 ( .A(n247), .Y(in_17bit_b[2]) );
  INVX1 U63 ( .A(n256), .Y(in_17bit_b[5]) );
  INVX1 U64 ( .A(n259), .Y(in_17bit_b[6]) );
  INVX1 U65 ( .A(n262), .Y(in_17bit_b[7]) );
  INVX1 U66 ( .A(n265), .Y(in_17bit_b[8]) );
  INVX1 U67 ( .A(n268), .Y(in_17bit_b[9]) );
  INVX1 U68 ( .A(n271), .Y(in_17bit_b[10]) );
  INVX1 U69 ( .A(n274), .Y(in_17bit_b[11]) );
  INVX1 U70 ( .A(n277), .Y(in_17bit_b[12]) );
  INVX1 U71 ( .A(n253), .Y(in_17bit_b[4]) );
  INVX1 U72 ( .A(n250), .Y(in_17bit_b[3]) );
  NAND2XL U73 ( .A(n2), .B(n12), .Y(n75) );
  NOR2X2 U74 ( .A(n33), .B(n177), .Y(n178) );
  NAND2XL U75 ( .A(n2), .B(n15), .Y(n164) );
  AOI21X1 U76 ( .A0(n28), .A1(n29), .B0(n287), .Y(n240) );
  NOR4XL U77 ( .A(in_8bit[4]), .B(n39), .C(in_8bit[6]), .D(n2), .Y(n28) );
  NAND2XL U78 ( .A(n1), .B(n19), .Y(n55) );
  OAI21XL U79 ( .A0(n293), .A1(n294), .B0(n292), .Y(N463) );
  AOI22X1 U80 ( .A0(N221), .A1(n291), .B0(N363), .B1(n290), .Y(n292) );
  INVX1 U81 ( .A(n212), .Y(n293) );
  NAND3XL U82 ( .A(n2), .B(n48), .C(n40), .Y(n192) );
  ADDFX2 U83 ( .A(in_17bit_b[16]), .B(in_17bit_b[12]), .CI(
        add_1_root_r112_carry_16_), .CO(add_1_root_r112_carry_17_), .S(
        add_1_root_r112_SUM_16_) );
  ADDFX2 U84 ( .A(add_1_root_r119_A_19_), .B(in_17bit_b[13]), .CI(
        add_1_root_r119_carry[19]), .CO(add_1_root_r119_carry[20]), .S(
        add_1_root_r119_SUM_19_) );
  ADDFX2 U85 ( .A(in_17bit_b[16]), .B(in_17bit_b[15]), .CI(
        add_3_root_r119_carry_17_), .CO(add_3_root_r119_carry_18_), .S(
        add_1_root_r119_A_17_) );
  ADDFX2 U86 ( .A(in_17bit_b[16]), .B(in_17bit_b[14]), .CI(
        add_2_root_r115_carry_17_), .CO(add_2_root_r115_carry_18_), .S(
        add_2_root_r115_SUM_17_) );
  ADDFX2 U87 ( .A(in_17bit_b[16]), .B(in_17bit_b[14]), .CI(
        add_1_root_r115_carry_20_), .CO(add_1_root_r115_carry_21_), .S(
        add_1_root_r115_SUM_20_) );
  ADDFX2 U88 ( .A(in_17bit_b[16]), .B(in_17bit_b[15]), .CI(
        add_2_root_r119_carry_20_), .CO(add_2_root_r119_carry_21_), .S(
        add_2_root_r119_SUM_20_) );
  ADDFX2 U89 ( .A(in_17bit_b[3]), .B(in_17bit_b[1]), .CI(
        add_1_root_r115_carry_7_), .CO(add_2_root_r115_carry_5_), .S(
        add_2_root_r115_SUM_4_) );
  ADDFX2 U90 ( .A(in_17bit_b[4]), .B(in_17bit_b[2]), .CI(
        add_2_root_r115_carry_5_), .CO(add_2_root_r115_carry_6_), .S(
        add_2_root_r115_SUM_5_) );
  ADDFX2 U91 ( .A(in_17bit_b[5]), .B(in_17bit_b[1]), .CI(
        add_1_root_r112_carry_5_), .CO(add_1_root_r112_carry_6_), .S(
        add_1_root_r112_SUM_5_) );
  ADDFX2 U92 ( .A(in_17bit_b[6]), .B(in_17bit_b[5]), .CI(
        add_3_root_r119_carry_7_), .CO(add_3_root_r119_carry_8_), .S(
        add_1_root_r119_A_7_) );
  ADDFX2 U93 ( .A(in_17bit_b[6]), .B(in_17bit_b[2]), .CI(
        add_1_root_r112_carry_6_), .CO(add_1_root_r112_carry_7_), .S(
        add_1_root_r112_SUM_6_) );
  ADDFX2 U94 ( .A(in_17bit_b[3]), .B(in_17bit_b[1]), .CI(
        add_1_root_r115_carry_7_), .CO(add_1_root_r115_carry_8_), .S(
        add_1_root_r115_SUM_7_) );
  ADDFX2 U95 ( .A(in_17bit_b[7]), .B(in_17bit_b[6]), .CI(
        add_3_root_r119_carry_8_), .CO(add_3_root_r119_carry_9_), .S(
        add_1_root_r119_A_8_) );
  ADDFX2 U96 ( .A(add_1_root_r119_A_7_), .B(in_17bit_b[1]), .CI(
        add_1_root_r119_carry[7]), .CO(add_1_root_r119_carry[8]), .S(
        add_1_root_r119_SUM_7_) );
  ADDFX2 U97 ( .A(in_17bit_b[2]), .B(in_17bit_b[1]), .CI(
        add_3_root_r119_carry_3_), .CO(add_2_root_r119_carry_7_), .S(
        add_2_root_r119_SUM_6_) );
  ADDFX2 U98 ( .A(in_17bit_b[4]), .B(in_17bit_b[2]), .CI(
        add_1_root_r115_carry_8_), .CO(add_1_root_r115_carry_9_), .S(
        add_1_root_r115_SUM_8_) );
  ADDFX2 U99 ( .A(in_17bit_b[8]), .B(in_17bit_b[7]), .CI(
        add_3_root_r119_carry_9_), .CO(add_3_root_r119_carry_10_), .S(
        add_1_root_r119_A_9_) );
  ADDFX2 U100 ( .A(add_1_root_r119_A_8_), .B(in_17bit_b[2]), .CI(
        add_1_root_r119_carry[8]), .CO(add_1_root_r119_carry[9]), .S(
        add_1_root_r119_SUM_8_) );
  ADDFX2 U101 ( .A(in_17bit_b[3]), .B(in_17bit_b[2]), .CI(
        add_2_root_r119_carry_7_), .CO(add_2_root_r119_carry_8_), .S(
        add_2_root_r119_SUM_7_) );
  ADDFX2 U102 ( .A(in_17bit_b[6]), .B(in_17bit_b[4]), .CI(
        add_2_root_r115_carry_7_), .CO(add_2_root_r115_carry_8_), .S(
        add_2_root_r115_SUM_7_) );
  ADDFX2 U103 ( .A(in_17bit_b[9]), .B(in_17bit_b[8]), .CI(
        add_3_root_r119_carry_10_), .CO(add_3_root_r119_carry_11_), .S(
        add_1_root_r119_A_10_) );
  ADDFX2 U104 ( .A(in_17bit_b[7]), .B(in_17bit_b[5]), .CI(
        add_2_root_r115_carry_8_), .CO(add_2_root_r115_carry_9_), .S(
        add_2_root_r115_SUM_8_) );
  ADDFX2 U105 ( .A(in_17bit_b[9]), .B(in_17bit_b[5]), .CI(
        add_1_root_r112_carry_9_), .CO(add_1_root_r112_carry_10_), .S(
        add_1_root_r112_SUM_9_) );
  ADDFX2 U106 ( .A(in_17bit_b[6]), .B(in_17bit_b[4]), .CI(
        add_1_root_r115_carry_10_), .CO(add_1_root_r115_carry_11_), .S(
        add_1_root_r115_SUM_10_) );
  ADDFX2 U107 ( .A(in_17bit_b[10]), .B(in_17bit_b[9]), .CI(
        add_3_root_r119_carry_11_), .CO(add_3_root_r119_carry_12_), .S(
        add_1_root_r119_A_11_) );
  ADDFX2 U108 ( .A(add_1_root_r119_A_10_), .B(in_17bit_b[4]), .CI(
        add_1_root_r119_carry[10]), .CO(add_1_root_r119_carry[11]), .S(
        add_1_root_r119_SUM_10_) );
  ADDFX2 U109 ( .A(in_17bit_b[5]), .B(in_17bit_b[4]), .CI(
        add_2_root_r119_carry_9_), .CO(add_2_root_r119_carry_10_), .S(
        add_2_root_r119_SUM_9_) );
  ADDFX2 U110 ( .A(in_17bit_b[8]), .B(in_17bit_b[6]), .CI(
        add_2_root_r115_carry_9_), .CO(add_2_root_r115_carry_10_), .S(
        add_2_root_r115_SUM_9_) );
  ADDFX2 U111 ( .A(in_17bit_b[10]), .B(in_17bit_b[6]), .CI(
        add_1_root_r112_carry_10_), .CO(add_1_root_r112_carry_11_), .S(
        add_1_root_r112_SUM_10_) );
  ADDFX2 U112 ( .A(in_17bit_b[7]), .B(in_17bit_b[5]), .CI(
        add_1_root_r115_carry_11_), .CO(add_1_root_r115_carry_12_), .S(
        add_1_root_r115_SUM_11_) );
  ADDFX2 U113 ( .A(in_17bit_b[11]), .B(in_17bit_b[10]), .CI(
        add_3_root_r119_carry_12_), .CO(add_3_root_r119_carry_13_), .S(
        add_1_root_r119_A_12_) );
  ADDFX2 U114 ( .A(add_1_root_r119_A_11_), .B(in_17bit_b[5]), .CI(
        add_1_root_r119_carry[11]), .CO(add_1_root_r119_carry[12]), .S(
        add_1_root_r119_SUM_11_) );
  ADDFX2 U115 ( .A(in_17bit_b[6]), .B(in_17bit_b[5]), .CI(
        add_2_root_r119_carry_10_), .CO(add_2_root_r119_carry_11_), .S(
        add_2_root_r119_SUM_10_) );
  ADDFX2 U116 ( .A(in_17bit_b[9]), .B(in_17bit_b[7]), .CI(
        add_2_root_r115_carry_10_), .CO(add_2_root_r115_carry_11_), .S(
        add_2_root_r115_SUM_10_) );
  ADDFX2 U117 ( .A(in_17bit_b[11]), .B(in_17bit_b[7]), .CI(
        add_1_root_r112_carry_11_), .CO(add_1_root_r112_carry_12_), .S(
        add_1_root_r112_SUM_11_) );
  ADDFX2 U118 ( .A(in_17bit_b[8]), .B(in_17bit_b[6]), .CI(
        add_1_root_r115_carry_12_), .CO(add_1_root_r115_carry_13_), .S(
        add_1_root_r115_SUM_12_) );
  ADDFX2 U119 ( .A(in_17bit_b[12]), .B(in_17bit_b[11]), .CI(
        add_3_root_r119_carry_13_), .CO(add_3_root_r119_carry_14_), .S(
        add_1_root_r119_A_13_) );
  ADDFX2 U120 ( .A(add_1_root_r119_A_12_), .B(in_17bit_b[6]), .CI(
        add_1_root_r119_carry[12]), .CO(add_1_root_r119_carry[13]), .S(
        add_1_root_r119_SUM_12_) );
  ADDFX2 U121 ( .A(in_17bit_b[7]), .B(in_17bit_b[6]), .CI(
        add_2_root_r119_carry_11_), .CO(add_2_root_r119_carry_12_), .S(
        add_2_root_r119_SUM_11_) );
  ADDFX2 U122 ( .A(in_17bit_b[10]), .B(in_17bit_b[8]), .CI(
        add_2_root_r115_carry_11_), .CO(add_2_root_r115_carry_12_), .S(
        add_2_root_r115_SUM_11_) );
  ADDFX2 U123 ( .A(in_17bit_b[12]), .B(in_17bit_b[8]), .CI(
        add_1_root_r112_carry_12_), .CO(add_1_root_r112_carry_13_), .S(
        add_1_root_r112_SUM_12_) );
  ADDFX2 U124 ( .A(in_17bit_b[9]), .B(in_17bit_b[7]), .CI(
        add_1_root_r115_carry_13_), .CO(add_1_root_r115_carry_14_), .S(
        add_1_root_r115_SUM_13_) );
  ADDFX2 U125 ( .A(in_17bit_b[13]), .B(in_17bit_b[12]), .CI(
        add_3_root_r119_carry_14_), .CO(add_3_root_r119_carry_15_), .S(
        add_1_root_r119_A_14_) );
  ADDFX2 U126 ( .A(add_1_root_r119_A_13_), .B(in_17bit_b[7]), .CI(
        add_1_root_r119_carry[13]), .CO(add_1_root_r119_carry[14]), .S(
        add_1_root_r119_SUM_13_) );
  ADDFX2 U127 ( .A(in_17bit_b[8]), .B(in_17bit_b[7]), .CI(
        add_2_root_r119_carry_12_), .CO(add_2_root_r119_carry_13_), .S(
        add_2_root_r119_SUM_12_) );
  ADDFX2 U128 ( .A(in_17bit_b[11]), .B(in_17bit_b[9]), .CI(
        add_2_root_r115_carry_12_), .CO(add_2_root_r115_carry_13_), .S(
        add_2_root_r115_SUM_12_) );
  ADDFX2 U129 ( .A(in_17bit_b[13]), .B(in_17bit_b[9]), .CI(
        add_1_root_r112_carry_13_), .CO(add_1_root_r112_carry_14_), .S(
        add_1_root_r112_SUM_13_) );
  ADDFX2 U130 ( .A(in_17bit_b[10]), .B(in_17bit_b[8]), .CI(
        add_1_root_r115_carry_14_), .CO(add_1_root_r115_carry_15_), .S(
        add_1_root_r115_SUM_14_) );
  ADDFX2 U131 ( .A(in_17bit_b[14]), .B(in_17bit_b[13]), .CI(
        add_3_root_r119_carry_15_), .CO(add_3_root_r119_carry_16_), .S(
        add_1_root_r119_A_15_) );
  ADDFX2 U132 ( .A(add_1_root_r119_A_14_), .B(in_17bit_b[8]), .CI(
        add_1_root_r119_carry[14]), .CO(add_1_root_r119_carry[15]), .S(
        add_1_root_r119_SUM_14_) );
  ADDFX2 U133 ( .A(in_17bit_b[9]), .B(in_17bit_b[8]), .CI(
        add_2_root_r119_carry_13_), .CO(add_2_root_r119_carry_14_), .S(
        add_2_root_r119_SUM_13_) );
  ADDFX2 U134 ( .A(in_17bit_b[12]), .B(in_17bit_b[10]), .CI(
        add_2_root_r115_carry_13_), .CO(add_2_root_r115_carry_14_), .S(
        add_2_root_r115_SUM_13_) );
  ADDFX2 U135 ( .A(in_17bit_b[14]), .B(in_17bit_b[10]), .CI(
        add_1_root_r112_carry_14_), .CO(add_1_root_r112_carry_15_), .S(
        add_1_root_r112_SUM_14_) );
  ADDFX2 U136 ( .A(in_17bit_b[11]), .B(in_17bit_b[9]), .CI(
        add_1_root_r115_carry_15_), .CO(add_1_root_r115_carry_16_), .S(
        add_1_root_r115_SUM_15_) );
  ADDFX2 U137 ( .A(add_1_root_r119_A_15_), .B(in_17bit_b[9]), .CI(
        add_1_root_r119_carry[15]), .CO(add_1_root_r119_carry[16]), .S(
        add_1_root_r119_SUM_15_) );
  ADDFX2 U138 ( .A(in_17bit_b[3]), .B(in_17bit_b[2]), .CI(
        add_3_root_r119_carry_4_), .CO(add_3_root_r119_carry_5_), .S(
        add_1_root_r119_A_4_) );
  ADDFX2 U139 ( .A(in_17bit_b[2]), .B(in_17bit_b[1]), .CI(
        add_3_root_r119_carry_3_), .CO(add_3_root_r119_carry_4_), .S(
        add_1_root_r119_A_3_) );
  ADDFX2 U140 ( .A(in_17bit_b[10]), .B(in_17bit_b[9]), .CI(
        add_2_root_r119_carry_14_), .CO(add_2_root_r119_carry_15_), .S(
        add_2_root_r119_SUM_14_) );
  ADDFX2 U141 ( .A(in_17bit_b[13]), .B(in_17bit_b[11]), .CI(
        add_2_root_r115_carry_14_), .CO(add_2_root_r115_carry_15_), .S(
        add_2_root_r115_SUM_14_) );
  ADDFX2 U142 ( .A(in_17bit_b[15]), .B(in_17bit_b[11]), .CI(
        add_1_root_r112_carry_15_), .CO(add_1_root_r112_carry_16_), .S(
        add_1_root_r112_SUM_15_) );
  ADDFX2 U143 ( .A(in_17bit_b[12]), .B(in_17bit_b[10]), .CI(
        add_1_root_r115_carry_16_), .CO(add_1_root_r115_carry_17_), .S(
        add_1_root_r115_SUM_16_) );
  ADDFX2 U144 ( .A(add_1_root_r119_A_16_), .B(in_17bit_b[10]), .CI(
        add_1_root_r119_carry[16]), .CO(add_1_root_r119_carry[17]), .S(
        add_1_root_r119_SUM_16_) );
  ADDFX2 U145 ( .A(in_17bit_b[11]), .B(in_17bit_b[10]), .CI(
        add_2_root_r119_carry_15_), .CO(add_2_root_r119_carry_16_), .S(
        add_2_root_r119_SUM_15_) );
  ADDFX2 U146 ( .A(in_17bit_b[14]), .B(in_17bit_b[12]), .CI(
        add_2_root_r115_carry_15_), .CO(add_2_root_r115_carry_16_), .S(
        add_2_root_r115_SUM_15_) );
  ADDFX2 U147 ( .A(in_17bit_b[13]), .B(in_17bit_b[11]), .CI(
        add_1_root_r115_carry_17_), .CO(add_1_root_r115_carry_18_), .S(
        add_1_root_r115_SUM_17_) );
  ADDFX2 U148 ( .A(add_1_root_r119_A_17_), .B(in_17bit_b[11]), .CI(
        add_1_root_r119_carry[17]), .CO(add_1_root_r119_carry[18]), .S(
        add_1_root_r119_SUM_17_) );
  ADDFX2 U149 ( .A(in_17bit_b[12]), .B(in_17bit_b[11]), .CI(
        add_2_root_r119_carry_16_), .CO(add_2_root_r119_carry_17_), .S(
        add_2_root_r119_SUM_16_) );
  ADDFX2 U150 ( .A(in_17bit_b[14]), .B(in_17bit_b[12]), .CI(
        add_1_root_r115_carry_18_), .CO(add_1_root_r115_carry_19_), .S(
        add_1_root_r115_SUM_18_) );
  ADDFX2 U151 ( .A(add_1_root_r119_A_18_), .B(in_17bit_b[12]), .CI(
        add_1_root_r119_carry[18]), .CO(add_1_root_r119_carry[19]), .S(
        add_1_root_r119_SUM_18_) );
  ADDFX2 U152 ( .A(in_17bit_b[15]), .B(in_17bit_b[13]), .CI(
        add_2_root_r115_carry_16_), .CO(add_2_root_r115_carry_17_), .S(
        add_2_root_r115_SUM_16_) );
  ADDFX2 U153 ( .A(in_17bit_b[13]), .B(in_17bit_b[12]), .CI(
        add_2_root_r119_carry_17_), .CO(add_2_root_r119_carry_18_), .S(
        add_2_root_r119_SUM_17_) );
  ADDFX2 U154 ( .A(in_17bit_b[5]), .B(in_17bit_b[3]), .CI(
        add_2_root_r115_carry_6_), .CO(add_2_root_r115_carry_7_), .S(
        add_2_root_r115_SUM_6_) );
  ADDFX2 U155 ( .A(in_17bit_b[7]), .B(in_17bit_b[3]), .CI(
        add_1_root_r112_carry_7_), .CO(add_1_root_r112_carry_8_), .S(
        add_1_root_r112_SUM_7_) );
  ADDFX2 U156 ( .A(in_17bit_b[8]), .B(in_17bit_b[4]), .CI(
        add_1_root_r112_carry_8_), .CO(add_1_root_r112_carry_9_), .S(
        add_1_root_r112_SUM_8_) );
  ADDFX2 U157 ( .A(in_17bit_b[5]), .B(in_17bit_b[3]), .CI(
        add_1_root_r115_carry_9_), .CO(add_1_root_r115_carry_10_), .S(
        add_1_root_r115_SUM_9_) );
  ADDFX2 U158 ( .A(in_17bit_b[4]), .B(in_17bit_b[3]), .CI(
        add_2_root_r119_carry_8_), .CO(add_2_root_r119_carry_9_), .S(
        add_2_root_r119_SUM_8_) );
  ADDFX2 U159 ( .A(in_17bit_b[15]), .B(in_17bit_b[14]), .CI(
        add_3_root_r119_carry_16_), .CO(add_3_root_r119_carry_17_), .S(
        add_1_root_r119_A_16_) );
  ADDFX2 U160 ( .A(in_17bit_b[4]), .B(in_17bit_b[3]), .CI(
        add_3_root_r119_carry_5_), .CO(add_3_root_r119_carry_6_), .S(
        add_1_root_r119_A_5_) );
  ADDFX2 U161 ( .A(in_17bit_b[5]), .B(in_17bit_b[4]), .CI(
        add_3_root_r119_carry_6_), .CO(add_3_root_r119_carry_7_), .S(
        add_1_root_r119_A_6_) );
  ADDFX2 U162 ( .A(in_17bit_b[15]), .B(in_17bit_b[13]), .CI(
        add_1_root_r115_carry_19_), .CO(add_1_root_r115_carry_20_), .S(
        add_1_root_r115_SUM_19_) );
  ADDFX2 U163 ( .A(in_17bit_b[14]), .B(in_17bit_b[13]), .CI(
        add_2_root_r119_carry_18_), .CO(add_2_root_r119_carry_19_), .S(
        add_2_root_r119_SUM_18_) );
  ADDFX2 U164 ( .A(add_1_root_r119_A_9_), .B(in_17bit_b[3]), .CI(
        add_1_root_r119_carry[9]), .CO(add_1_root_r119_carry[10]), .S(
        add_1_root_r119_SUM_9_) );
  ADDFX2 U165 ( .A(in_17bit_b[15]), .B(in_17bit_b[14]), .CI(
        add_2_root_r119_carry_19_), .CO(add_2_root_r119_carry_20_), .S(
        add_2_root_r119_SUM_19_) );
  NAND2X1 U166 ( .A(n285), .B(n284), .Y(N461) );
  AOI22X1 U167 ( .A0(N122), .A1(n287), .B0(N219), .B1(n291), .Y(n284) );
  AOI22X1 U168 ( .A0(N361), .A1(n290), .B0(n212), .B1(in_17bit_b[14]), .Y(n285) );
  NAND2X1 U169 ( .A(n289), .B(n288), .Y(N462) );
  AOI22X1 U170 ( .A0(N123), .A1(n287), .B0(N220), .B1(n291), .Y(n288) );
  AOI22X1 U171 ( .A0(N362), .A1(n290), .B0(n212), .B1(in_17bit_b[15]), .Y(n289) );
  INVX1 U172 ( .A(n40), .Y(n39) );
  INVX1 U173 ( .A(in_8bit[0]), .Y(n47) );
  INVX1 U174 ( .A(in_8bit[3]), .Y(n41) );
  INVX1 U175 ( .A(in_8bit[4]), .Y(n48) );
  XNOR2X1 U176 ( .A(n54), .B(n30), .Y(N29) );
  NAND2X1 U177 ( .A(sub_add_54_b0_carry[15]), .B(n211), .Y(n30) );
  NOR3X1 U178 ( .A(n213), .B(n41), .C(n47), .Y(n239) );
  CLKINVX3 U179 ( .A(n241), .Y(in_17bit_b[0]) );
  NAND3BX1 U180 ( .AN(n39), .B(n213), .C(in_8bit[3]), .Y(n236) );
  NAND3X1 U181 ( .A(n238), .B(n39), .C(n183), .Y(n184) );
  NOR2XL U182 ( .A(n2), .B(n48), .Y(n183) );
  NAND2BX1 U183 ( .AN(n193), .B(n47), .Y(n189) );
  CLKINVX3 U184 ( .A(n286), .Y(in_17bit_b[15]) );
  OR2X2 U185 ( .A(n188), .B(n187), .Y(n290) );
  NOR2X1 U186 ( .A(n236), .B(n234), .Y(n187) );
  NOR2X1 U187 ( .A(n189), .B(n235), .Y(n188) );
  OR2X2 U188 ( .A(n191), .B(n190), .Y(n291) );
  NOR2X1 U189 ( .A(n189), .B(n236), .Y(n190) );
  NOR2X1 U190 ( .A(n234), .B(n235), .Y(n191) );
  OAI2BB1X1 U191 ( .A0N(n186), .A1N(n185), .B0(n184), .Y(n287) );
  NOR2BX1 U192 ( .AN(in_8bit[1]), .B(n192), .Y(n185) );
  NOR2BX1 U193 ( .AN(n239), .B(n182), .Y(n186) );
  OAI2BB1X1 U194 ( .A0N(n238), .A1N(n195), .B0(n194), .Y(n212) );
  INVX1 U195 ( .A(n192), .Y(n195) );
  NAND3BX1 U196 ( .AN(n193), .B(n239), .C(n39), .Y(n194) );
  INVX1 U197 ( .A(n74), .Y(n71) );
  INVX1 U198 ( .A(n82), .Y(n79) );
  INVX1 U199 ( .A(n90), .Y(n87) );
  INVX1 U200 ( .A(n98), .Y(n95) );
  INVX1 U201 ( .A(n163), .Y(n160) );
  NAND2X1 U202 ( .A(n243), .B(n242), .Y(N447) );
  AOI22X1 U203 ( .A0(N108), .A1(n287), .B0(N205), .B1(n291), .Y(n242) );
  AOI22X1 U204 ( .A0(N347), .A1(n290), .B0(n212), .B1(in_17bit_b[0]), .Y(n243)
         );
  NAND2X1 U205 ( .A(n246), .B(n245), .Y(N448) );
  AOI22X1 U206 ( .A0(N109), .A1(n287), .B0(N206), .B1(n291), .Y(n245) );
  AOI22X1 U207 ( .A0(N348), .A1(n290), .B0(n212), .B1(in_17bit_b[1]), .Y(n246)
         );
  NAND2X1 U208 ( .A(n249), .B(n248), .Y(N449) );
  AOI22X1 U209 ( .A0(N110), .A1(n287), .B0(N207), .B1(n291), .Y(n248) );
  AOI22X1 U210 ( .A0(N349), .A1(n290), .B0(n212), .B1(in_17bit_b[2]), .Y(n249)
         );
  NAND2X1 U211 ( .A(n252), .B(n251), .Y(N450) );
  AOI22X1 U212 ( .A0(N111), .A1(n287), .B0(N208), .B1(n291), .Y(n251) );
  AOI22X1 U213 ( .A0(N350), .A1(n290), .B0(n212), .B1(in_17bit_b[3]), .Y(n252)
         );
  NAND2X1 U214 ( .A(n255), .B(n254), .Y(N451) );
  AOI22X1 U215 ( .A0(N112), .A1(n287), .B0(N209), .B1(n291), .Y(n254) );
  AOI22X1 U216 ( .A0(N351), .A1(n290), .B0(n212), .B1(in_17bit_b[4]), .Y(n255)
         );
  NAND2X1 U217 ( .A(n258), .B(n257), .Y(N452) );
  AOI22X1 U218 ( .A0(N113), .A1(n287), .B0(N210), .B1(n291), .Y(n257) );
  AOI22X1 U219 ( .A0(N352), .A1(n290), .B0(n212), .B1(in_17bit_b[5]), .Y(n258)
         );
  NAND2X1 U220 ( .A(n261), .B(n260), .Y(N453) );
  AOI22X1 U221 ( .A0(N114), .A1(n287), .B0(N211), .B1(n291), .Y(n260) );
  AOI22X1 U222 ( .A0(N353), .A1(n290), .B0(n212), .B1(in_17bit_b[6]), .Y(n261)
         );
  NAND2X1 U223 ( .A(n264), .B(n263), .Y(N454) );
  AOI22X1 U224 ( .A0(N115), .A1(n287), .B0(N212), .B1(n291), .Y(n263) );
  AOI22X1 U225 ( .A0(N354), .A1(n290), .B0(n212), .B1(in_17bit_b[7]), .Y(n264)
         );
  NAND2X1 U226 ( .A(n267), .B(n266), .Y(N455) );
  AOI22X1 U227 ( .A0(N116), .A1(n287), .B0(N213), .B1(n291), .Y(n266) );
  AOI22X1 U228 ( .A0(N355), .A1(n290), .B0(n212), .B1(in_17bit_b[8]), .Y(n267)
         );
  NAND2X1 U229 ( .A(n270), .B(n269), .Y(N456) );
  AOI22X1 U230 ( .A0(N117), .A1(n287), .B0(N214), .B1(n291), .Y(n269) );
  AOI22X1 U231 ( .A0(N356), .A1(n290), .B0(n212), .B1(in_17bit_b[9]), .Y(n270)
         );
  NAND2X1 U232 ( .A(n273), .B(n272), .Y(N457) );
  AOI22X1 U233 ( .A0(N118), .A1(n287), .B0(N215), .B1(n291), .Y(n272) );
  AOI22X1 U234 ( .A0(N357), .A1(n290), .B0(n212), .B1(in_17bit_b[10]), .Y(n273) );
  NAND2X1 U235 ( .A(n276), .B(n275), .Y(N458) );
  AOI22X1 U236 ( .A0(N119), .A1(n287), .B0(N216), .B1(n291), .Y(n275) );
  AOI22X1 U237 ( .A0(N358), .A1(n290), .B0(n212), .B1(in_17bit_b[11]), .Y(n276) );
  NAND2X1 U238 ( .A(n279), .B(n278), .Y(N459) );
  AOI22X1 U239 ( .A0(N120), .A1(n287), .B0(N217), .B1(n291), .Y(n278) );
  AOI22X1 U240 ( .A0(N359), .A1(n290), .B0(n212), .B1(in_17bit_b[12]), .Y(n279) );
  NAND2X1 U241 ( .A(n282), .B(n281), .Y(N460) );
  AOI22X1 U242 ( .A0(N121), .A1(n287), .B0(N218), .B1(n291), .Y(n281) );
  AOI22X1 U243 ( .A0(N360), .A1(n290), .B0(n212), .B1(in_17bit_b[13]), .Y(n282) );
  INVX1 U244 ( .A(in_8bit[5]), .Y(n40) );
  INVX1 U245 ( .A(n66), .Y(n63) );
  OAI21XL U246 ( .A0(n42), .A1(n76), .B0(n75), .Y(n81) );
  OAI21XL U247 ( .A0(n42), .A1(n100), .B0(n99), .Y(n162) );
  NAND2XL U248 ( .A(n2), .B(n14), .Y(n99) );
  OAI21XL U249 ( .A0(n42), .A1(n92), .B0(n91), .Y(n97) );
  NAND2XL U250 ( .A(n2), .B(n13), .Y(n91) );
  OAI21XL U251 ( .A0(n42), .A1(n170), .B0(n164), .Y(n174) );
  NOR4BXL U252 ( .AN(n237), .B(n47), .C(in_8bit[1]), .D(in_8bit[2]), .Y(n238)
         );
  NOR2XL U253 ( .A(in_8bit[6]), .B(in_8bit[3]), .Y(n237) );
  NAND3XL U254 ( .A(in_8bit[2]), .B(n41), .C(n39), .Y(n235) );
  INVXL U255 ( .A(in_8bit[2]), .Y(n213) );
  NAND4BBX1 U256 ( .AN(n290), .BN(n291), .C(n240), .D(n293), .Y(N446) );
  NAND4XL U257 ( .A(in_8bit[1]), .B(n2), .C(n233), .D(n47), .Y(n234) );
  NOR2XL U258 ( .A(in_8bit[6]), .B(in_8bit[4]), .Y(n233) );
  AOI22XL U259 ( .A0(in_17bit[0]), .A1(n51), .B0(in_17bit[0]), .B1(n54), .Y(
        n241) );
  AOI22X1 U260 ( .A0(N27), .A1(n51), .B0(in_17bit[14]), .B1(n50), .Y(n283) );
  AOI22X1 U261 ( .A0(N26), .A1(n51), .B0(in_17bit[13]), .B1(n54), .Y(n280) );
  AOI22X1 U262 ( .A0(N28), .A1(n51), .B0(in_17bit[15]), .B1(n54), .Y(n286) );
  AOI22XL U263 ( .A0(N14), .A1(n51), .B0(in_17bit[1]), .B1(n54), .Y(n244) );
  AOI22XL U264 ( .A0(N15), .A1(n51), .B0(in_17bit[2]), .B1(n54), .Y(n247) );
  AOI22X1 U265 ( .A0(N16), .A1(n51), .B0(in_17bit[3]), .B1(n50), .Y(n250) );
  AOI22X1 U266 ( .A0(N17), .A1(n51), .B0(in_17bit[4]), .B1(n50), .Y(n253) );
  AOI22X1 U267 ( .A0(N18), .A1(n51), .B0(in_17bit[5]), .B1(n54), .Y(n256) );
  AOI22X1 U268 ( .A0(N19), .A1(n51), .B0(in_17bit[6]), .B1(n50), .Y(n259) );
  AOI22X1 U269 ( .A0(N20), .A1(n51), .B0(in_17bit[7]), .B1(n50), .Y(n262) );
  AOI22X1 U270 ( .A0(N21), .A1(n51), .B0(in_17bit[8]), .B1(n50), .Y(n265) );
  AOI22X1 U271 ( .A0(N22), .A1(n51), .B0(in_17bit[9]), .B1(n54), .Y(n268) );
  AOI22X1 U272 ( .A0(N23), .A1(n51), .B0(in_17bit[10]), .B1(n50), .Y(n271) );
  AOI22X1 U273 ( .A0(N24), .A1(n51), .B0(in_17bit[11]), .B1(n54), .Y(n274) );
  AOI22X1 U274 ( .A0(N25), .A1(n51), .B0(in_17bit[12]), .B1(n50), .Y(n277) );
  AND2X2 U275 ( .A(n160), .B(n15), .Y(n31) );
  NAND4BXL U276 ( .AN(n44), .B(in_8bit[4]), .C(in_8bit[1]), .D(in_8bit[6]), 
        .Y(n193) );
  NAND2X1 U277 ( .A(n36), .B(n11), .Y(n66) );
  AND2X2 U278 ( .A(n31), .B(n18), .Y(n32) );
  AND2X2 U279 ( .A(n32), .B(n3), .Y(n33) );
  NAND2BX1 U280 ( .AN(n66), .B(n6), .Y(n74) );
  NAND2X1 U281 ( .A(n71), .B(n12), .Y(n82) );
  NAND2X1 U282 ( .A(n79), .B(n7), .Y(n90) );
  NAND2X1 U283 ( .A(n87), .B(n13), .Y(n98) );
  NAND2X1 U284 ( .A(n95), .B(n14), .Y(n163) );
  INVXL U285 ( .A(in_8bit[6]), .Y(n182) );
  AND2X2 U286 ( .A(n33), .B(n4), .Y(n34) );
  INVX1 U287 ( .A(in_17bit[0]), .Y(n196) );
  INVX1 U288 ( .A(in_17bit[1]), .Y(n197) );
  INVX1 U289 ( .A(in_17bit[2]), .Y(n198) );
  INVX1 U290 ( .A(in_17bit[3]), .Y(n199) );
  INVX1 U291 ( .A(in_17bit[4]), .Y(n200) );
  INVX1 U292 ( .A(in_17bit[5]), .Y(n201) );
  INVX1 U293 ( .A(in_17bit[6]), .Y(n202) );
  INVX1 U294 ( .A(in_17bit[7]), .Y(n203) );
  INVX1 U295 ( .A(in_17bit[8]), .Y(n204) );
  INVX1 U296 ( .A(in_17bit[9]), .Y(n205) );
  INVX1 U297 ( .A(in_17bit[10]), .Y(n206) );
  INVX1 U298 ( .A(in_17bit[11]), .Y(n207) );
  INVX1 U299 ( .A(in_17bit[12]), .Y(n208) );
  INVX1 U300 ( .A(in_17bit[13]), .Y(n209) );
  INVX1 U301 ( .A(in_17bit[14]), .Y(n210) );
  INVX1 U302 ( .A(in_17bit[15]), .Y(n211) );
  INVXL U303 ( .A(n51), .Y(n50) );
  XNOR2X1 U304 ( .A(n16), .B(sub_add_75_b0_carry[13]), .Y(n35) );
  AOI2BB2X1 U305 ( .B0(n101), .B1(n2), .A0N(n44), .A1N(neg_mul[14]), .Y(n158)
         );
  INVX1 U306 ( .A(n100), .Y(n101) );
  INVX1 U307 ( .A(n92), .Y(n93) );
  INVX1 U308 ( .A(n84), .Y(n85) );
  INVX1 U309 ( .A(n170), .Y(n171) );
  INVX1 U310 ( .A(n68), .Y(n69) );
  INVX1 U311 ( .A(n60), .Y(n61) );
  AOI2BB2X1 U312 ( .B0(n77), .B1(n2), .A0N(n44), .A1N(neg_mul[11]), .Y(n78) );
  INVX1 U313 ( .A(n76), .Y(n77) );
  MX2X1 U314 ( .A(neg_mul[22]), .B(N480), .S0(n181), .Y(out[15]) );
  MX2X1 U315 ( .A(neg_mul[23]), .B(N481), .S0(n181), .Y(out[16]) );
  NOR2X1 U316 ( .A(out[0]), .B(neg_mul[8]), .Y(n36) );
  NAND2BX1 U317 ( .AN(n36), .B(neg_mul[9]), .Y(n60) );
  NAND2X1 U318 ( .A(neg_mul[10]), .B(n66), .Y(n68) );
  NAND2X1 U319 ( .A(neg_mul[11]), .B(n74), .Y(n76) );
  NAND2X1 U320 ( .A(neg_mul[12]), .B(n82), .Y(n84) );
  NAND2X1 U321 ( .A(neg_mul[13]), .B(n90), .Y(n92) );
  NAND2X1 U322 ( .A(neg_mul[15]), .B(n163), .Y(n170) );
  NAND2X1 U323 ( .A(neg_mul[14]), .B(n98), .Y(n100) );
  BUFX8 U324 ( .A(n299), .Y(out[1]) );
  AOI211X2 U325 ( .A0(n52), .A1(n58), .B0(n57), .C0(n36), .Y(n299) );
  NAND2XL U326 ( .A(N29), .B(n51), .Y(n294) );
  AOI211X4 U327 ( .A0(n23), .A1(n174), .B0(n173), .C0(n31), .Y(out[8]) );
  AOI211X4 U328 ( .A0(n20), .A1(n97), .B0(n96), .C0(n95), .Y(out[6]) );
  AOI211X4 U329 ( .A0(n20), .A1(n81), .B0(n80), .C0(n79), .Y(n296) );
  NOR2X4 U330 ( .A(n31), .B(n180), .Y(n175) );
  XNOR2X4 U331 ( .A(n176), .B(n3), .Y(out[10]) );
  XNOR2X4 U332 ( .A(n178), .B(n4), .Y(out[11]) );
  AND2X1 U333 ( .A(add_1_root_r112_carry_20_), .B(in_17bit_b[16]), .Y(
        add_1_root_r112_SUM_21_) );
  XOR2X1 U334 ( .A(in_17bit_b[16]), .B(add_1_root_r112_carry_20_), .Y(
        add_1_root_r112_SUM_20_) );
  AND2X1 U335 ( .A(add_1_root_r112_carry_19_), .B(in_17bit_b[15]), .Y(
        add_1_root_r112_carry_20_) );
  XOR2X1 U336 ( .A(in_17bit_b[15]), .B(add_1_root_r112_carry_19_), .Y(
        add_1_root_r112_SUM_19_) );
  AND2X1 U337 ( .A(add_1_root_r112_carry_18_), .B(in_17bit_b[14]), .Y(
        add_1_root_r112_carry_19_) );
  XOR2X1 U338 ( .A(in_17bit_b[14]), .B(add_1_root_r112_carry_18_), .Y(
        add_1_root_r112_SUM_18_) );
  AND2X1 U339 ( .A(add_1_root_r112_carry_17_), .B(in_17bit_b[13]), .Y(
        add_1_root_r112_carry_18_) );
  XOR2X1 U340 ( .A(in_17bit_b[13]), .B(add_1_root_r112_carry_17_), .Y(
        add_1_root_r112_SUM_17_) );
  AND2X1 U341 ( .A(add_2_root_r119_carry_21_), .B(in_17bit_b[16]), .Y(
        add_2_root_r119_SUM_22_) );
  XOR2X1 U342 ( .A(in_17bit_b[16]), .B(add_2_root_r119_carry_21_), .Y(
        add_2_root_r119_SUM_21_) );
  AND2X1 U343 ( .A(add_1_root_r119_carry[22]), .B(in_17bit_b[16]), .Y(
        add_1_root_r119_SUM_23_) );
  XOR2X1 U344 ( .A(in_17bit_b[16]), .B(add_1_root_r119_carry[22]), .Y(
        add_1_root_r119_SUM_22_) );
  AND2X1 U345 ( .A(add_1_root_r119_carry[21]), .B(in_17bit_b[15]), .Y(
        add_1_root_r119_carry[22]) );
  XOR2X1 U346 ( .A(in_17bit_b[15]), .B(add_1_root_r119_carry[21]), .Y(
        add_1_root_r119_SUM_21_) );
  AND2X1 U347 ( .A(add_1_root_r119_carry[20]), .B(in_17bit_b[14]), .Y(
        add_1_root_r119_carry[21]) );
  XOR2X1 U348 ( .A(in_17bit_b[14]), .B(add_1_root_r119_carry[20]), .Y(
        add_1_root_r119_SUM_20_) );
  AND2X1 U349 ( .A(add_1_root_r119_A_6_), .B(in_17bit_b[0]), .Y(
        add_1_root_r119_carry[7]) );
  XOR2X1 U350 ( .A(in_17bit_b[0]), .B(add_1_root_r119_A_6_), .Y(
        add_1_root_r119_SUM_6_) );
  AND2X1 U351 ( .A(add_3_root_r119_carry_18_), .B(in_17bit_b[16]), .Y(
        add_1_root_r119_A_19_) );
  XOR2X1 U352 ( .A(in_17bit_b[16]), .B(add_3_root_r119_carry_18_), .Y(
        add_1_root_r119_A_18_) );
  AND2X1 U353 ( .A(in_17bit_b[1]), .B(in_17bit_b[0]), .Y(
        add_3_root_r119_carry_3_) );
  XOR2X1 U354 ( .A(in_17bit_b[0]), .B(in_17bit_b[1]), .Y(add_1_root_r119_A_2_)
         );
  AND2X1 U355 ( .A(add_2_root_r115_carry_19_), .B(in_17bit_b[16]), .Y(
        add_2_root_r115_SUM_20_) );
  XOR2X1 U356 ( .A(in_17bit_b[16]), .B(add_2_root_r115_carry_19_), .Y(
        add_2_root_r115_SUM_19_) );
  AND2X1 U357 ( .A(add_2_root_r115_carry_18_), .B(in_17bit_b[15]), .Y(
        add_2_root_r115_carry_19_) );
  XOR2X1 U358 ( .A(in_17bit_b[15]), .B(add_2_root_r115_carry_18_), .Y(
        add_2_root_r115_SUM_18_) );
  AND2X1 U359 ( .A(add_1_root_r115_carry_22_), .B(in_17bit_b[16]), .Y(
        add_1_root_r115_SUM_23_) );
  XOR2X1 U360 ( .A(in_17bit_b[16]), .B(add_1_root_r115_carry_22_), .Y(
        add_1_root_r115_SUM_22_) );
  AND2X1 U361 ( .A(add_1_root_r115_carry_21_), .B(in_17bit_b[15]), .Y(
        add_1_root_r115_carry_22_) );
  XOR2X1 U362 ( .A(in_17bit_b[15]), .B(add_1_root_r115_carry_21_), .Y(
        add_1_root_r115_SUM_21_) );
  AND2X1 U363 ( .A(in_17bit_b[2]), .B(in_17bit_b[0]), .Y(
        add_1_root_r115_carry_7_) );
  XOR2X1 U364 ( .A(in_17bit_b[0]), .B(in_17bit_b[2]), .Y(
        add_1_root_r115_SUM_6_) );
  XOR2X1 U365 ( .A(n211), .B(sub_add_54_b0_carry[15]), .Y(N28) );
  AND2X1 U366 ( .A(sub_add_54_b0_carry[14]), .B(n210), .Y(
        sub_add_54_b0_carry[15]) );
  XOR2X1 U367 ( .A(n210), .B(sub_add_54_b0_carry[14]), .Y(N27) );
  AND2X1 U368 ( .A(sub_add_54_b0_carry[13]), .B(n209), .Y(
        sub_add_54_b0_carry[14]) );
  XOR2X1 U369 ( .A(n209), .B(sub_add_54_b0_carry[13]), .Y(N26) );
  AND2X1 U370 ( .A(sub_add_54_b0_carry[12]), .B(n208), .Y(
        sub_add_54_b0_carry[13]) );
  XOR2X1 U371 ( .A(n208), .B(sub_add_54_b0_carry[12]), .Y(N25) );
  AND2X1 U372 ( .A(sub_add_54_b0_carry[11]), .B(n207), .Y(
        sub_add_54_b0_carry[12]) );
  XOR2X1 U373 ( .A(n207), .B(sub_add_54_b0_carry[11]), .Y(N24) );
  AND2X1 U374 ( .A(sub_add_54_b0_carry[10]), .B(n206), .Y(
        sub_add_54_b0_carry[11]) );
  XOR2X1 U375 ( .A(n206), .B(sub_add_54_b0_carry[10]), .Y(N23) );
  AND2X1 U376 ( .A(sub_add_54_b0_carry[9]), .B(n205), .Y(
        sub_add_54_b0_carry[10]) );
  XOR2X1 U377 ( .A(n205), .B(sub_add_54_b0_carry[9]), .Y(N22) );
  AND2X1 U378 ( .A(sub_add_54_b0_carry[8]), .B(n204), .Y(
        sub_add_54_b0_carry[9]) );
  XOR2X1 U379 ( .A(n204), .B(sub_add_54_b0_carry[8]), .Y(N21) );
  AND2X1 U380 ( .A(sub_add_54_b0_carry[7]), .B(n203), .Y(
        sub_add_54_b0_carry[8]) );
  XOR2X1 U381 ( .A(n203), .B(sub_add_54_b0_carry[7]), .Y(N20) );
  AND2X1 U382 ( .A(sub_add_54_b0_carry[6]), .B(n202), .Y(
        sub_add_54_b0_carry[7]) );
  XOR2X1 U383 ( .A(n202), .B(sub_add_54_b0_carry[6]), .Y(N19) );
  AND2X1 U384 ( .A(sub_add_54_b0_carry[5]), .B(n201), .Y(
        sub_add_54_b0_carry[6]) );
  XOR2X1 U385 ( .A(n201), .B(sub_add_54_b0_carry[5]), .Y(N18) );
  AND2X1 U386 ( .A(sub_add_54_b0_carry[4]), .B(n200), .Y(
        sub_add_54_b0_carry[5]) );
  XOR2X1 U387 ( .A(n200), .B(sub_add_54_b0_carry[4]), .Y(N17) );
  AND2X1 U388 ( .A(sub_add_54_b0_carry[3]), .B(n199), .Y(
        sub_add_54_b0_carry[4]) );
  XOR2X1 U389 ( .A(n199), .B(sub_add_54_b0_carry[3]), .Y(N16) );
  AND2X1 U390 ( .A(sub_add_54_b0_carry[2]), .B(n198), .Y(
        sub_add_54_b0_carry[3]) );
  XOR2X1 U391 ( .A(n198), .B(sub_add_54_b0_carry[2]), .Y(N15) );
  AND2X1 U392 ( .A(n196), .B(n197), .Y(sub_add_54_b0_carry[2]) );
  XOR2X1 U393 ( .A(n197), .B(n196), .Y(N14) );
  XOR2X1 U394 ( .A(n17), .B(sub_add_75_b0_carry[16]), .Y(N481) );
  AND2X1 U395 ( .A(sub_add_75_b0_carry[15]), .B(n10), .Y(
        sub_add_75_b0_carry[16]) );
  XOR2X1 U396 ( .A(n10), .B(sub_add_75_b0_carry[15]), .Y(N480) );
  AND2X1 U397 ( .A(sub_add_75_b0_carry[14]), .B(n9), .Y(
        sub_add_75_b0_carry[15]) );
  XOR2X1 U398 ( .A(n9), .B(sub_add_75_b0_carry[14]), .Y(N479) );
  AND2X1 U399 ( .A(sub_add_75_b0_carry[13]), .B(n16), .Y(
        sub_add_75_b0_carry[14]) );
  AND2X1 U400 ( .A(n34), .B(n5), .Y(sub_add_75_b0_carry[13]) );
  AND2X1 U401 ( .A(in_17bit_b[0]), .B(in_17bit_b[4]), .Y(
        add_1_root_r112_carry_5_) );
endmodule


module multi16_3_DW01_add_0 ( A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, 
        A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, 
        A_4_, B_23_, B_22_, B_21_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, 
        B_14_, B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, 
        SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, 
        SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, 
        SUM_7_ );
  input A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_,
         A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, B_23_, B_22_,
         B_21_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_,
         B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_;
  output SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_,
         SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_,
         SUM_8_, SUM_7_;
  wire   n1, n2, n3, n4;
  wire   [23:7] carry;

  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry[7]), .CO(carry[8]), .S(SUM_7_)
         );
  ADDFX2 U1_21 ( .A(A_21_), .B(B_21_), .CI(carry[21]), .CO(carry[22]), .S(
        SUM_21_) );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry[20]), .CO(carry[21]), .S(
        SUM_20_) );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry[19]), .CO(carry[20]), .S(
        SUM_19_) );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry[18]), .CO(carry[19]), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry[17]), .CO(carry[18]), .S(
        SUM_17_) );
  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry[16]), .CO(carry[17]), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry[15]), .CO(carry[16]), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry[14]), .CO(carry[15]), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry[13]), .CO(carry[14]), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry[12]), .CO(carry[13]), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry[11]), .CO(carry[12]), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry[10]), .CO(carry[11]), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry[9]), .CO(carry[10]), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry[8]), .CO(carry[9]), .S(SUM_8_)
         );
  ADDFX2 U1_22 ( .A(A_22_), .B(B_22_), .CI(carry[22]), .CO(carry[23]), .S(
        SUM_22_) );
  AND2X2 U1 ( .A(A_4_), .B(B_4_), .Y(n1) );
  XOR2X1 U2 ( .A(B_23_), .B(carry[23]), .Y(SUM_23_) );
  OAI2BB1X1 U3 ( .A0N(n2), .A1N(A_6_), .B0(n3), .Y(carry[7]) );
  OAI21XL U4 ( .A0(A_6_), .A1(n2), .B0(B_6_), .Y(n3) );
  OAI2BB1X1 U5 ( .A0N(n1), .A1N(A_5_), .B0(n4), .Y(n2) );
  OAI21XL U6 ( .A0(A_5_), .A1(n1), .B0(B_5_), .Y(n4) );
endmodule


module multi16_3_DW01_add_4 ( A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, 
        A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, 
        B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, 
        B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, SUM_22_, SUM_21_, SUM_20_, 
        SUM_19_, SUM_18_, SUM_17_, SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, 
        SUM_11_, SUM_10_, SUM_9_, SUM_8_, SUM_7_ );
  input A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_,
         A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, B_20_, B_19_,
         B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, B_10_, B_9_,
         B_8_, B_7_, B_6_, B_5_;
  output SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_,
         SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_,
         SUM_7_;
  wire   carry_21_, carry_20_, carry_19_, carry_18_, carry_17_, carry_16_,
         carry_15_, carry_14_, carry_13_, carry_12_, carry_11_, carry_10_,
         carry_9_, carry_8_, carry_7_, n1;

  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry_16_), .CO(carry_17_), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry_15_), .CO(carry_16_), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry_14_), .CO(carry_15_), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry_13_), .CO(carry_14_), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry_12_), .CO(carry_13_), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry_11_), .CO(carry_12_), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry_10_), .CO(carry_11_), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry_9_), .CO(carry_10_), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry_8_), .CO(carry_9_), .S(SUM_8_)
         );
  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry_7_), .CO(carry_8_), .S(SUM_7_)
         );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry_20_), .CO(carry_21_), .S(
        SUM_20_) );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry_19_), .CO(carry_20_), .S(
        SUM_19_) );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry_18_), .CO(carry_19_), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry_17_), .CO(carry_18_), .S(
        SUM_17_) );
  ADDFX2 U1_21 ( .A(A_21_), .B(B_21_), .CI(carry_21_), .CO(SUM_22_), .S(
        SUM_21_) );
  OAI2BB1X1 U1 ( .A0N(A_6_), .A1N(B_6_), .B0(n1), .Y(carry_7_) );
  OAI211X1 U2 ( .A0(B_6_), .A1(A_6_), .B0(A_5_), .C0(B_5_), .Y(n1) );
endmodule


module multi16_3_DW01_add_6 ( A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, 
        A_16_, A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, 
        A_6_, A_5_, A_4_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, 
        B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, 
        SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, 
        SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, 
        SUM_7_ );
  input A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_,
         A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, B_20_,
         B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, B_10_,
         B_9_, B_8_, B_7_, B_6_, B_5_, B_4_;
  output SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_,
         SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_,
         SUM_8_, SUM_7_;
  wire   n1, n2, n3, n4, n5, n6;
  wire   [21:7] carry;

  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry[7]), .CO(carry[8]), .S(SUM_7_)
         );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry[18]), .CO(carry[19]), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry[17]), .CO(carry[18]), .S(
        SUM_17_) );
  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry[16]), .CO(carry[17]), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry[15]), .CO(carry[16]), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry[14]), .CO(carry[15]), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry[13]), .CO(carry[14]), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry[12]), .CO(carry[13]), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry[11]), .CO(carry[12]), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry[10]), .CO(carry[11]), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry[9]), .CO(carry[10]), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry[8]), .CO(carry[9]), .S(SUM_8_)
         );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry[19]), .CO(carry[20]), .S(
        SUM_19_) );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry[20]), .CO(carry[21]), .S(
        SUM_20_) );
  AND2X2 U1 ( .A(A_22_), .B(n2), .Y(n1) );
  AND2X2 U2 ( .A(A_21_), .B(carry[21]), .Y(n2) );
  AND2X2 U3 ( .A(A_4_), .B(B_4_), .Y(n3) );
  XOR2X1 U4 ( .A(A_23_), .B(n1), .Y(SUM_23_) );
  XOR2X1 U5 ( .A(A_21_), .B(carry[21]), .Y(SUM_21_) );
  XOR2X1 U6 ( .A(A_22_), .B(n2), .Y(SUM_22_) );
  OAI2BB1X1 U7 ( .A0N(n4), .A1N(A_6_), .B0(n5), .Y(carry[7]) );
  OAI21XL U8 ( .A0(A_6_), .A1(n4), .B0(B_6_), .Y(n5) );
  OAI2BB1X1 U9 ( .A0N(n3), .A1N(A_5_), .B0(n6), .Y(n4) );
  OAI21XL U10 ( .A0(A_5_), .A1(n3), .B0(B_5_), .Y(n6) );
endmodule


module multi16_3 ( in_17bit, in_8bit, out );
  input [16:0] in_17bit;
  input [7:0] in_8bit;
  output [16:0] out;
  wire   n256, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26,
         N27, N28, N29, N108, N109, N110, N111, N112, N113, N114, N115, N116,
         N117, N118, N119, N120, N121, N122, N123, N205, N206, N207, N208,
         N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, N219,
         N220, N221, N347, N348, N349, N350, N351, N352, N353, N354, N355,
         N356, N357, N358, N359, N360, N361, N362, N363, N446, N447, N448,
         N449, N450, N451, N452, N453, N454, N455, N456, N457, N458, N459,
         N460, N461, N462, N463, N480, add_2_root_r119_carry_10_,
         add_2_root_r119_carry_11_, add_2_root_r119_carry_12_,
         add_2_root_r119_carry_13_, add_2_root_r119_carry_14_,
         add_2_root_r119_carry_15_, add_2_root_r119_carry_16_,
         add_2_root_r119_carry_17_, add_2_root_r119_carry_18_,
         add_2_root_r119_carry_19_, add_2_root_r119_carry_20_,
         add_2_root_r119_carry_21_, add_2_root_r119_carry_7_,
         add_2_root_r119_carry_8_, add_2_root_r119_carry_9_,
         add_2_root_r119_SUM_6_, add_2_root_r119_SUM_7_,
         add_2_root_r119_SUM_8_, add_2_root_r119_SUM_9_,
         add_2_root_r119_SUM_10_, add_2_root_r119_SUM_11_,
         add_2_root_r119_SUM_12_, add_2_root_r119_SUM_13_,
         add_2_root_r119_SUM_14_, add_2_root_r119_SUM_15_,
         add_2_root_r119_SUM_16_, add_2_root_r119_SUM_17_,
         add_2_root_r119_SUM_18_, add_2_root_r119_SUM_19_,
         add_2_root_r119_SUM_20_, add_2_root_r119_SUM_21_,
         add_2_root_r119_SUM_22_, add_1_root_r119_SUM_6_,
         add_1_root_r119_SUM_7_, add_1_root_r119_SUM_8_,
         add_1_root_r119_SUM_9_, add_1_root_r119_SUM_10_,
         add_1_root_r119_SUM_11_, add_1_root_r119_SUM_12_,
         add_1_root_r119_SUM_13_, add_1_root_r119_SUM_14_,
         add_1_root_r119_SUM_15_, add_1_root_r119_SUM_16_,
         add_1_root_r119_SUM_17_, add_1_root_r119_SUM_18_,
         add_1_root_r119_SUM_19_, add_1_root_r119_SUM_20_,
         add_1_root_r119_SUM_21_, add_1_root_r119_SUM_22_,
         add_1_root_r119_SUM_23_, add_1_root_r119_A_2_, add_1_root_r119_A_3_,
         add_1_root_r119_A_4_, add_1_root_r119_A_5_, add_1_root_r119_A_6_,
         add_1_root_r119_A_7_, add_1_root_r119_A_8_, add_1_root_r119_A_9_,
         add_1_root_r119_A_10_, add_1_root_r119_A_11_, add_1_root_r119_A_12_,
         add_1_root_r119_A_13_, add_1_root_r119_A_14_, add_1_root_r119_A_15_,
         add_1_root_r119_A_16_, add_1_root_r119_A_17_, add_1_root_r119_A_18_,
         add_1_root_r119_A_19_, add_3_root_r119_carry_10_,
         add_3_root_r119_carry_11_, add_3_root_r119_carry_12_,
         add_3_root_r119_carry_13_, add_3_root_r119_carry_14_,
         add_3_root_r119_carry_15_, add_3_root_r119_carry_16_,
         add_3_root_r119_carry_17_, add_3_root_r119_carry_18_,
         add_3_root_r119_carry_3_, add_3_root_r119_carry_4_,
         add_3_root_r119_carry_5_, add_3_root_r119_carry_6_,
         add_3_root_r119_carry_7_, add_3_root_r119_carry_8_,
         add_3_root_r119_carry_9_, add_1_root_r112_carry_10_,
         add_1_root_r112_carry_11_, add_1_root_r112_carry_12_,
         add_1_root_r112_carry_13_, add_1_root_r112_carry_14_,
         add_1_root_r112_carry_15_, add_1_root_r112_carry_16_,
         add_1_root_r112_carry_17_, add_1_root_r112_carry_18_,
         add_1_root_r112_carry_19_, add_1_root_r112_carry_20_,
         add_1_root_r112_carry_5_, add_1_root_r112_carry_6_,
         add_1_root_r112_carry_7_, add_1_root_r112_carry_8_,
         add_1_root_r112_carry_9_, add_1_root_r112_SUM_1_,
         add_1_root_r112_SUM_2_, add_1_root_r112_SUM_3_,
         add_1_root_r112_SUM_4_, add_1_root_r112_SUM_5_,
         add_1_root_r112_SUM_6_, add_1_root_r112_SUM_7_,
         add_1_root_r112_SUM_8_, add_1_root_r112_SUM_9_,
         add_1_root_r112_SUM_10_, add_1_root_r112_SUM_11_,
         add_1_root_r112_SUM_12_, add_1_root_r112_SUM_13_,
         add_1_root_r112_SUM_14_, add_1_root_r112_SUM_15_,
         add_1_root_r112_SUM_16_, add_1_root_r112_SUM_17_,
         add_1_root_r112_SUM_18_, add_1_root_r112_SUM_19_,
         add_1_root_r112_SUM_20_, add_1_root_r112_SUM_21_,
         add_2_root_r115_carry_10_, add_2_root_r115_carry_11_,
         add_2_root_r115_carry_12_, add_2_root_r115_carry_13_,
         add_2_root_r115_carry_14_, add_2_root_r115_carry_15_,
         add_2_root_r115_carry_16_, add_2_root_r115_carry_17_,
         add_2_root_r115_carry_18_, add_2_root_r115_carry_19_,
         add_2_root_r115_carry_5_, add_2_root_r115_carry_6_,
         add_2_root_r115_carry_7_, add_2_root_r115_carry_8_,
         add_2_root_r115_carry_9_, add_2_root_r115_SUM_4_,
         add_2_root_r115_SUM_5_, add_2_root_r115_SUM_6_,
         add_2_root_r115_SUM_7_, add_2_root_r115_SUM_8_,
         add_2_root_r115_SUM_9_, add_2_root_r115_SUM_10_,
         add_2_root_r115_SUM_11_, add_2_root_r115_SUM_12_,
         add_2_root_r115_SUM_13_, add_2_root_r115_SUM_14_,
         add_2_root_r115_SUM_15_, add_2_root_r115_SUM_16_,
         add_2_root_r115_SUM_17_, add_2_root_r115_SUM_18_,
         add_2_root_r115_SUM_19_, add_2_root_r115_SUM_20_,
         add_1_root_r115_carry_10_, add_1_root_r115_carry_11_,
         add_1_root_r115_carry_12_, add_1_root_r115_carry_13_,
         add_1_root_r115_carry_14_, add_1_root_r115_carry_15_,
         add_1_root_r115_carry_16_, add_1_root_r115_carry_17_,
         add_1_root_r115_carry_18_, add_1_root_r115_carry_19_,
         add_1_root_r115_carry_20_, add_1_root_r115_carry_21_,
         add_1_root_r115_carry_22_, add_1_root_r115_carry_7_,
         add_1_root_r115_carry_8_, add_1_root_r115_carry_9_,
         add_1_root_r115_SUM_6_, add_1_root_r115_SUM_7_,
         add_1_root_r115_SUM_8_, add_1_root_r115_SUM_9_,
         add_1_root_r115_SUM_10_, add_1_root_r115_SUM_11_,
         add_1_root_r115_SUM_12_, add_1_root_r115_SUM_13_,
         add_1_root_r115_SUM_14_, add_1_root_r115_SUM_15_,
         add_1_root_r115_SUM_16_, add_1_root_r115_SUM_17_,
         add_1_root_r115_SUM_18_, add_1_root_r115_SUM_19_,
         add_1_root_r115_SUM_20_, add_1_root_r115_SUM_21_,
         add_1_root_r115_SUM_22_, add_1_root_r115_SUM_23_, n2, n3, n4, n5, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n158, n160, n161, n162,
         n163, n164, n168, n170, n171, n172, n173, n174, n175, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255;
  wire   [16:0] in_17bit_b;
  wire   [23:8] neg_mul;
  wire   [15:13] sub_add_75_b0_carry;
  wire   [16:2] sub_add_54_b0_carry;
  wire   [22:7] add_1_root_r119_carry;

  multi16_3_DW01_add_0 add_0_root_r119 ( .A_22_(add_2_root_r119_SUM_22_), 
        .A_21_(add_2_root_r119_SUM_21_), .A_20_(add_2_root_r119_SUM_20_), 
        .A_19_(add_2_root_r119_SUM_19_), .A_18_(add_2_root_r119_SUM_18_), 
        .A_17_(add_2_root_r119_SUM_17_), .A_16_(add_2_root_r119_SUM_16_), 
        .A_15_(add_2_root_r119_SUM_15_), .A_14_(add_2_root_r119_SUM_14_), 
        .A_13_(add_2_root_r119_SUM_13_), .A_12_(add_2_root_r119_SUM_12_), 
        .A_11_(add_2_root_r119_SUM_11_), .A_10_(add_2_root_r119_SUM_10_), 
        .A_9_(add_2_root_r119_SUM_9_), .A_8_(add_2_root_r119_SUM_8_), .A_7_(
        add_2_root_r119_SUM_7_), .A_6_(add_2_root_r119_SUM_6_), .A_5_(
        add_1_root_r119_A_2_), .A_4_(in_17bit_b[0]), .B_23_(
        add_1_root_r119_SUM_23_), .B_22_(add_1_root_r119_SUM_22_), .B_21_(
        add_1_root_r119_SUM_21_), .B_20_(add_1_root_r119_SUM_20_), .B_19_(
        add_1_root_r119_SUM_19_), .B_18_(add_1_root_r119_SUM_18_), .B_17_(
        add_1_root_r119_SUM_17_), .B_16_(add_1_root_r119_SUM_16_), .B_15_(
        add_1_root_r119_SUM_15_), .B_14_(add_1_root_r119_SUM_14_), .B_13_(
        add_1_root_r119_SUM_13_), .B_12_(add_1_root_r119_SUM_12_), .B_11_(
        add_1_root_r119_SUM_11_), .B_10_(add_1_root_r119_SUM_10_), .B_9_(
        add_1_root_r119_SUM_9_), .B_8_(add_1_root_r119_SUM_8_), .B_7_(
        add_1_root_r119_SUM_7_), .B_6_(add_1_root_r119_SUM_6_), .B_5_(
        add_1_root_r119_A_5_), .B_4_(add_1_root_r119_A_4_), .SUM_23_(N363), 
        .SUM_22_(N362), .SUM_21_(N361), .SUM_20_(N360), .SUM_19_(N359), 
        .SUM_18_(N358), .SUM_17_(N357), .SUM_16_(N356), .SUM_15_(N355), 
        .SUM_14_(N354), .SUM_13_(N353), .SUM_12_(N352), .SUM_11_(N351), 
        .SUM_10_(N350), .SUM_9_(N349), .SUM_8_(N348), .SUM_7_(N347) );
  multi16_3_DW01_add_4 add_0_root_r112 ( .A_21_(in_17bit_b[16]), .A_20_(
        in_17bit_b[15]), .A_19_(in_17bit_b[14]), .A_18_(in_17bit_b[13]), 
        .A_17_(in_17bit_b[12]), .A_16_(in_17bit_b[11]), .A_15_(in_17bit_b[10]), 
        .A_14_(in_17bit_b[9]), .A_13_(in_17bit_b[8]), .A_12_(in_17bit_b[7]), 
        .A_11_(in_17bit_b[6]), .A_10_(in_17bit_b[5]), .A_9_(in_17bit_b[4]), 
        .A_8_(in_17bit_b[3]), .A_7_(in_17bit_b[2]), .A_6_(in_17bit_b[1]), 
        .A_5_(in_17bit_b[0]), .B_21_(add_1_root_r112_SUM_21_), .B_20_(
        add_1_root_r112_SUM_20_), .B_19_(add_1_root_r112_SUM_19_), .B_18_(
        add_1_root_r112_SUM_18_), .B_17_(add_1_root_r112_SUM_17_), .B_16_(
        add_1_root_r112_SUM_16_), .B_15_(add_1_root_r112_SUM_15_), .B_14_(
        add_1_root_r112_SUM_14_), .B_13_(add_1_root_r112_SUM_13_), .B_12_(
        add_1_root_r112_SUM_12_), .B_11_(add_1_root_r112_SUM_11_), .B_10_(
        add_1_root_r112_SUM_10_), .B_9_(add_1_root_r112_SUM_9_), .B_8_(
        add_1_root_r112_SUM_8_), .B_7_(add_1_root_r112_SUM_7_), .B_6_(
        add_1_root_r112_SUM_6_), .B_5_(add_1_root_r112_SUM_5_), .SUM_22_(N123), 
        .SUM_21_(N122), .SUM_20_(N121), .SUM_19_(N120), .SUM_18_(N119), 
        .SUM_17_(N118), .SUM_16_(N117), .SUM_15_(N116), .SUM_14_(N115), 
        .SUM_13_(N114), .SUM_12_(N113), .SUM_11_(N112), .SUM_10_(N111), 
        .SUM_9_(N110), .SUM_8_(N109), .SUM_7_(N108) );
  multi16_3_DW01_add_6 add_0_root_r115 ( .A_23_(add_1_root_r115_SUM_23_), 
        .A_22_(add_1_root_r115_SUM_22_), .A_21_(add_1_root_r115_SUM_21_), 
        .A_20_(add_1_root_r115_SUM_20_), .A_19_(add_1_root_r115_SUM_19_), 
        .A_18_(add_1_root_r115_SUM_18_), .A_17_(add_1_root_r115_SUM_17_), 
        .A_16_(add_1_root_r115_SUM_16_), .A_15_(add_1_root_r115_SUM_15_), 
        .A_14_(add_1_root_r115_SUM_14_), .A_13_(add_1_root_r115_SUM_13_), 
        .A_12_(add_1_root_r115_SUM_12_), .A_11_(add_1_root_r115_SUM_11_), 
        .A_10_(add_1_root_r115_SUM_10_), .A_9_(add_1_root_r115_SUM_9_), .A_8_(
        add_1_root_r115_SUM_8_), .A_7_(add_1_root_r115_SUM_7_), .A_6_(
        add_1_root_r115_SUM_6_), .A_5_(in_17bit_b[1]), .A_4_(in_17bit_b[0]), 
        .B_20_(add_2_root_r115_SUM_20_), .B_19_(add_2_root_r115_SUM_19_), 
        .B_18_(add_2_root_r115_SUM_18_), .B_17_(add_2_root_r115_SUM_17_), 
        .B_16_(add_2_root_r115_SUM_16_), .B_15_(add_2_root_r115_SUM_15_), 
        .B_14_(add_2_root_r115_SUM_14_), .B_13_(add_2_root_r115_SUM_13_), 
        .B_12_(add_2_root_r115_SUM_12_), .B_11_(add_2_root_r115_SUM_11_), 
        .B_10_(add_2_root_r115_SUM_10_), .B_9_(add_2_root_r115_SUM_9_), .B_8_(
        add_2_root_r115_SUM_8_), .B_7_(add_2_root_r115_SUM_7_), .B_6_(
        add_2_root_r115_SUM_6_), .B_5_(add_2_root_r115_SUM_5_), .B_4_(
        add_2_root_r115_SUM_4_), .SUM_23_(N221), .SUM_22_(N220), .SUM_21_(N219), .SUM_20_(N218), .SUM_19_(N217), .SUM_18_(N216), .SUM_17_(N215), .SUM_16_(
        N214), .SUM_15_(N213), .SUM_14_(N212), .SUM_13_(N211), .SUM_12_(N210), 
        .SUM_11_(N209), .SUM_10_(N208), .SUM_9_(N207), .SUM_8_(N206), .SUM_7_(
        N205) );
  TLATX1 neg_mul_reg_19_ ( .G(N446), .D(N459), .QN(n10) );
  TLATX1 neg_mul_reg_18_ ( .G(N446), .D(N458), .QN(n5) );
  TLATX1 neg_mul_reg_17_ ( .G(N446), .D(N457), .Q(neg_mul[17]), .QN(n16) );
  TLATX1 neg_mul_reg_16_ ( .G(N446), .D(N456), .QN(n8) );
  TLATX1 neg_mul_reg_15_ ( .G(N446), .D(N455), .QN(n7) );
  TLATX1 neg_mul_reg_14_ ( .G(N446), .D(N454), .QN(n6) );
  TLATX1 neg_mul_reg_12_ ( .G(N446), .D(N452), .Q(neg_mul[12]), .QN(n3) );
  TLATX1 neg_mul_reg_11_ ( .G(N446), .D(N451), .Q(neg_mul[11]), .QN(n15) );
  TLATX1 neg_mul_reg_10_ ( .G(N446), .D(N450), .QN(n18) );
  TLATX1 neg_mul_reg_9_ ( .G(N446), .D(N449), .Q(n2), .QN(n12) );
  TLATX1 neg_mul_reg_8_ ( .G(N446), .D(N448), .Q(neg_mul[8]) );
  TLATX1 neg_mul_reg_23_ ( .G(N446), .D(N463), .Q(neg_mul[23]), .QN(n4) );
  TLATX1 neg_mul_reg_22_ ( .G(N446), .D(N462), .Q(neg_mul[22]), .QN(n11) );
  TLATX1 neg_mul_reg_21_ ( .G(N446), .D(N461), .QN(n28) );
  TLATX1 neg_mul_reg_20_ ( .G(N446), .D(N460), .QN(n13) );
  TLATX1 neg_mul_reg_13_ ( .G(N446), .D(N453), .Q(neg_mul[13]), .QN(n9) );
  TLATX1 neg_mul_reg_7_ ( .G(N446), .D(N447), .Q(out[0]), .QN(n20) );
  CLKINVX1 U2 ( .A(n63), .Y(n61) );
  INVX1 U3 ( .A(n61), .Y(n62) );
  CLKINVX8 U4 ( .A(n58), .Y(n63) );
  CLKINVX3 U5 ( .A(n255), .Y(in_17bit_b[16]) );
  XOR2X2 U6 ( .A(n25), .B(in_17bit[16]), .Y(n65) );
  BUFX3 U7 ( .A(n256), .Y(out[13]) );
  MXI2XL U8 ( .A(n13), .B(n44), .S0(n87), .Y(n256) );
  CLKINVX3 U9 ( .A(n56), .Y(n55) );
  INVX1 U10 ( .A(in_8bit[7]), .Y(n56) );
  AOI2BB2X2 U11 ( .B0(n25), .B1(n9), .A0N(n55), .A1N(n76), .Y(n78) );
  INVX1 U12 ( .A(n45), .Y(n24) );
  MXI2X1 U13 ( .A(n28), .B(n14), .S0(n87), .Y(out[14]) );
  CLKINVX2 U14 ( .A(n21), .Y(n87) );
  INVX1 U15 ( .A(n96), .Y(n92) );
  AOI22X1 U16 ( .A0(N27), .A1(n61), .B0(in_17bit[14]), .B1(n62), .Y(n244) );
  XNOR2X1 U17 ( .A(n28), .B(sub_add_75_b0_carry[14]), .Y(n14) );
  XNOR2X1 U18 ( .A(neg_mul[23]), .B(n46), .Y(n17) );
  XNOR2X4 U19 ( .A(n25), .B(n63), .Y(n68) );
  XNOR2X4 U20 ( .A(n25), .B(n58), .Y(n67) );
  OAI21X2 U21 ( .A0(n78), .A1(n63), .B0(n77), .Y(n79) );
  XNOR2X2 U22 ( .A(n25), .B(n59), .Y(n70) );
  NOR2X4 U23 ( .A(n73), .B(n71), .Y(n72) );
  XOR2X4 U24 ( .A(n26), .B(n18), .Y(out[3]) );
  XOR2X4 U25 ( .A(n66), .B(neg_mul[8]), .Y(n19) );
  INVX8 U26 ( .A(n19), .Y(out[1]) );
  NAND2BX4 U27 ( .AN(n20), .B(n65), .Y(n66) );
  INVX8 U28 ( .A(n60), .Y(n59) );
  XNOR2X2 U29 ( .A(n25), .B(n59), .Y(n21) );
  NAND2X4 U30 ( .A(n69), .B(n68), .Y(n26) );
  XOR2X4 U31 ( .A(n74), .B(neg_mul[12]), .Y(out[5]) );
  CLKINVX3 U32 ( .A(n60), .Y(n23) );
  NOR2BX4 U33 ( .AN(n24), .B(n67), .Y(n27) );
  XOR2X4 U34 ( .A(n85), .B(neg_mul[17]), .Y(out[10]) );
  OR2X4 U35 ( .A(n21), .B(n40), .Y(n34) );
  INVXL U36 ( .A(in_8bit[0]), .Y(n53) );
  INVXL U37 ( .A(in_8bit[4]), .Y(n52) );
  XOR2X4 U38 ( .A(n72), .B(neg_mul[11]), .Y(out[4]) );
  BUFX20 U39 ( .A(in_8bit[7]), .Y(n25) );
  NOR2X4 U40 ( .A(n81), .B(n70), .Y(n82) );
  INVX8 U41 ( .A(n60), .Y(n58) );
  NOR2X4 U42 ( .A(n86), .B(n39), .Y(n85) );
  NOR2X4 U43 ( .A(n36), .B(n86), .Y(n84) );
  INVX8 U44 ( .A(n33), .Y(out[11]) );
  INVX8 U45 ( .A(in_17bit[16]), .Y(n60) );
  XNOR2X4 U46 ( .A(n25), .B(n23), .Y(n86) );
  NOR2X2 U47 ( .A(n21), .B(n38), .Y(n83) );
  OR2X2 U48 ( .A(n86), .B(n43), .Y(n35) );
  AOI2BB2X2 U49 ( .B0(n75), .B1(n25), .A0N(n55), .A1N(neg_mul[13]), .Y(n80) );
  CLKBUFXL U50 ( .A(in_8bit[1]), .Y(n54) );
  INVX1 U51 ( .A(n205), .Y(in_17bit_b[1]) );
  INVX1 U52 ( .A(n244), .Y(in_17bit_b[14]) );
  INVX1 U53 ( .A(n241), .Y(in_17bit_b[13]) );
  INVX1 U54 ( .A(n208), .Y(in_17bit_b[2]) );
  INVX1 U55 ( .A(n229), .Y(in_17bit_b[9]) );
  INVX1 U56 ( .A(n235), .Y(in_17bit_b[11]) );
  INVX1 U57 ( .A(n238), .Y(in_17bit_b[12]) );
  INVX1 U58 ( .A(n217), .Y(in_17bit_b[5]) );
  INVX1 U59 ( .A(n220), .Y(in_17bit_b[6]) );
  INVX1 U60 ( .A(n223), .Y(in_17bit_b[7]) );
  INVX1 U61 ( .A(n226), .Y(in_17bit_b[8]) );
  INVX1 U62 ( .A(n232), .Y(in_17bit_b[10]) );
  INVX1 U63 ( .A(n214), .Y(in_17bit_b[4]) );
  INVX1 U64 ( .A(n211), .Y(in_17bit_b[3]) );
  XOR2X4 U65 ( .A(n27), .B(n2), .Y(out[2]) );
  XOR2X2 U66 ( .A(n35), .B(n10), .Y(out[12]) );
  AOI21X1 U67 ( .A0(n29), .A1(n30), .B0(n248), .Y(n201) );
  NOR4XL U68 ( .A(in_8bit[4]), .B(in_8bit[5]), .C(in_8bit[6]), .D(n25), .Y(n29) );
  NOR4XL U69 ( .A(n54), .B(in_8bit[0]), .C(in_8bit[2]), .D(in_8bit[3]), .Y(n30) );
  AND4X1 U70 ( .A(n54), .B(n25), .C(n195), .D(n53), .Y(n31) );
  NAND2X1 U71 ( .A(n32), .B(n54), .Y(n88) );
  NOR3X1 U72 ( .A(n50), .B(n51), .C(n53), .Y(n200) );
  NAND3X1 U73 ( .A(in_8bit[2]), .B(n51), .C(in_8bit[5]), .Y(n196) );
  ADDFX2 U74 ( .A(in_17bit_b[16]), .B(in_17bit_b[12]), .CI(
        add_1_root_r112_carry_16_), .CO(add_1_root_r112_carry_17_), .S(
        add_1_root_r112_SUM_16_) );
  ADDFX2 U75 ( .A(add_1_root_r119_A_19_), .B(in_17bit_b[13]), .CI(
        add_1_root_r119_carry[19]), .CO(add_1_root_r119_carry[20]), .S(
        add_1_root_r119_SUM_19_) );
  ADDFX2 U76 ( .A(in_17bit_b[16]), .B(in_17bit_b[15]), .CI(
        add_3_root_r119_carry_17_), .CO(add_3_root_r119_carry_18_), .S(
        add_1_root_r119_A_17_) );
  ADDFX2 U77 ( .A(in_17bit_b[16]), .B(in_17bit_b[14]), .CI(
        add_2_root_r115_carry_17_), .CO(add_2_root_r115_carry_18_), .S(
        add_2_root_r115_SUM_17_) );
  ADDFX2 U78 ( .A(in_17bit_b[16]), .B(in_17bit_b[14]), .CI(
        add_1_root_r115_carry_20_), .CO(add_1_root_r115_carry_21_), .S(
        add_1_root_r115_SUM_20_) );
  ADDFX2 U79 ( .A(in_17bit_b[16]), .B(in_17bit_b[15]), .CI(
        add_2_root_r119_carry_20_), .CO(add_2_root_r119_carry_21_), .S(
        add_2_root_r119_SUM_20_) );
  AND3X1 U80 ( .A(n25), .B(n52), .C(n57), .Y(n32) );
  NOR2XL U81 ( .A(n25), .B(n52), .Y(n89) );
  ADDFX2 U82 ( .A(in_17bit_b[3]), .B(in_17bit_b[1]), .CI(
        add_1_root_r115_carry_7_), .CO(add_2_root_r115_carry_5_), .S(
        add_2_root_r115_SUM_4_) );
  ADDFX2 U83 ( .A(in_17bit_b[4]), .B(in_17bit_b[2]), .CI(
        add_2_root_r115_carry_5_), .CO(add_2_root_r115_carry_6_), .S(
        add_2_root_r115_SUM_5_) );
  ADDFX2 U84 ( .A(in_17bit_b[5]), .B(in_17bit_b[1]), .CI(
        add_1_root_r112_carry_5_), .CO(add_1_root_r112_carry_6_), .S(
        add_1_root_r112_SUM_5_) );
  ADDFX2 U85 ( .A(in_17bit_b[6]), .B(in_17bit_b[5]), .CI(
        add_3_root_r119_carry_7_), .CO(add_3_root_r119_carry_8_), .S(
        add_1_root_r119_A_7_) );
  ADDFX2 U86 ( .A(in_17bit_b[6]), .B(in_17bit_b[2]), .CI(
        add_1_root_r112_carry_6_), .CO(add_1_root_r112_carry_7_), .S(
        add_1_root_r112_SUM_6_) );
  ADDFX2 U87 ( .A(in_17bit_b[3]), .B(in_17bit_b[1]), .CI(
        add_1_root_r115_carry_7_), .CO(add_1_root_r115_carry_8_), .S(
        add_1_root_r115_SUM_7_) );
  ADDFX2 U88 ( .A(in_17bit_b[7]), .B(in_17bit_b[6]), .CI(
        add_3_root_r119_carry_8_), .CO(add_3_root_r119_carry_9_), .S(
        add_1_root_r119_A_8_) );
  ADDFX2 U89 ( .A(add_1_root_r119_A_7_), .B(in_17bit_b[1]), .CI(
        add_1_root_r119_carry[7]), .CO(add_1_root_r119_carry[8]), .S(
        add_1_root_r119_SUM_7_) );
  ADDFX2 U90 ( .A(in_17bit_b[2]), .B(in_17bit_b[1]), .CI(
        add_3_root_r119_carry_3_), .CO(add_2_root_r119_carry_7_), .S(
        add_2_root_r119_SUM_6_) );
  ADDFX2 U91 ( .A(in_17bit_b[4]), .B(in_17bit_b[2]), .CI(
        add_1_root_r115_carry_8_), .CO(add_1_root_r115_carry_9_), .S(
        add_1_root_r115_SUM_8_) );
  ADDFX2 U92 ( .A(in_17bit_b[8]), .B(in_17bit_b[7]), .CI(
        add_3_root_r119_carry_9_), .CO(add_3_root_r119_carry_10_), .S(
        add_1_root_r119_A_9_) );
  ADDFX2 U93 ( .A(add_1_root_r119_A_8_), .B(in_17bit_b[2]), .CI(
        add_1_root_r119_carry[8]), .CO(add_1_root_r119_carry[9]), .S(
        add_1_root_r119_SUM_8_) );
  ADDFX2 U94 ( .A(in_17bit_b[3]), .B(in_17bit_b[2]), .CI(
        add_2_root_r119_carry_7_), .CO(add_2_root_r119_carry_8_), .S(
        add_2_root_r119_SUM_7_) );
  ADDFX2 U95 ( .A(in_17bit_b[6]), .B(in_17bit_b[4]), .CI(
        add_2_root_r115_carry_7_), .CO(add_2_root_r115_carry_8_), .S(
        add_2_root_r115_SUM_7_) );
  ADDFX2 U96 ( .A(in_17bit_b[8]), .B(in_17bit_b[4]), .CI(
        add_1_root_r112_carry_8_), .CO(add_1_root_r112_carry_9_), .S(
        add_1_root_r112_SUM_8_) );
  ADDFX2 U97 ( .A(in_17bit_b[9]), .B(in_17bit_b[8]), .CI(
        add_3_root_r119_carry_10_), .CO(add_3_root_r119_carry_11_), .S(
        add_1_root_r119_A_10_) );
  ADDFX2 U98 ( .A(in_17bit_b[7]), .B(in_17bit_b[5]), .CI(
        add_2_root_r115_carry_8_), .CO(add_2_root_r115_carry_9_), .S(
        add_2_root_r115_SUM_8_) );
  ADDFX2 U99 ( .A(in_17bit_b[9]), .B(in_17bit_b[5]), .CI(
        add_1_root_r112_carry_9_), .CO(add_1_root_r112_carry_10_), .S(
        add_1_root_r112_SUM_9_) );
  ADDFX2 U100 ( .A(in_17bit_b[6]), .B(in_17bit_b[4]), .CI(
        add_1_root_r115_carry_10_), .CO(add_1_root_r115_carry_11_), .S(
        add_1_root_r115_SUM_10_) );
  ADDFX2 U101 ( .A(in_17bit_b[10]), .B(in_17bit_b[9]), .CI(
        add_3_root_r119_carry_11_), .CO(add_3_root_r119_carry_12_), .S(
        add_1_root_r119_A_11_) );
  ADDFX2 U102 ( .A(in_17bit_b[5]), .B(in_17bit_b[4]), .CI(
        add_2_root_r119_carry_9_), .CO(add_2_root_r119_carry_10_), .S(
        add_2_root_r119_SUM_9_) );
  ADDFX2 U103 ( .A(in_17bit_b[10]), .B(in_17bit_b[6]), .CI(
        add_1_root_r112_carry_10_), .CO(add_1_root_r112_carry_11_), .S(
        add_1_root_r112_SUM_10_) );
  ADDFX2 U104 ( .A(in_17bit_b[7]), .B(in_17bit_b[5]), .CI(
        add_1_root_r115_carry_11_), .CO(add_1_root_r115_carry_12_), .S(
        add_1_root_r115_SUM_11_) );
  ADDFX2 U105 ( .A(in_17bit_b[11]), .B(in_17bit_b[10]), .CI(
        add_3_root_r119_carry_12_), .CO(add_3_root_r119_carry_13_), .S(
        add_1_root_r119_A_12_) );
  ADDFX2 U106 ( .A(add_1_root_r119_A_11_), .B(in_17bit_b[5]), .CI(
        add_1_root_r119_carry[11]), .CO(add_1_root_r119_carry[12]), .S(
        add_1_root_r119_SUM_11_) );
  ADDFX2 U107 ( .A(in_17bit_b[6]), .B(in_17bit_b[5]), .CI(
        add_2_root_r119_carry_10_), .CO(add_2_root_r119_carry_11_), .S(
        add_2_root_r119_SUM_10_) );
  ADDFX2 U108 ( .A(in_17bit_b[9]), .B(in_17bit_b[7]), .CI(
        add_2_root_r115_carry_10_), .CO(add_2_root_r115_carry_11_), .S(
        add_2_root_r115_SUM_10_) );
  ADDFX2 U109 ( .A(in_17bit_b[11]), .B(in_17bit_b[7]), .CI(
        add_1_root_r112_carry_11_), .CO(add_1_root_r112_carry_12_), .S(
        add_1_root_r112_SUM_11_) );
  ADDFX2 U110 ( .A(in_17bit_b[8]), .B(in_17bit_b[6]), .CI(
        add_1_root_r115_carry_12_), .CO(add_1_root_r115_carry_13_), .S(
        add_1_root_r115_SUM_12_) );
  ADDFX2 U111 ( .A(in_17bit_b[12]), .B(in_17bit_b[11]), .CI(
        add_3_root_r119_carry_13_), .CO(add_3_root_r119_carry_14_), .S(
        add_1_root_r119_A_13_) );
  ADDFX2 U112 ( .A(add_1_root_r119_A_12_), .B(in_17bit_b[6]), .CI(
        add_1_root_r119_carry[12]), .CO(add_1_root_r119_carry[13]), .S(
        add_1_root_r119_SUM_12_) );
  ADDFX2 U113 ( .A(in_17bit_b[7]), .B(in_17bit_b[6]), .CI(
        add_2_root_r119_carry_11_), .CO(add_2_root_r119_carry_12_), .S(
        add_2_root_r119_SUM_11_) );
  ADDFX2 U114 ( .A(in_17bit_b[10]), .B(in_17bit_b[8]), .CI(
        add_2_root_r115_carry_11_), .CO(add_2_root_r115_carry_12_), .S(
        add_2_root_r115_SUM_11_) );
  ADDFX2 U115 ( .A(in_17bit_b[12]), .B(in_17bit_b[8]), .CI(
        add_1_root_r112_carry_12_), .CO(add_1_root_r112_carry_13_), .S(
        add_1_root_r112_SUM_12_) );
  ADDFX2 U116 ( .A(in_17bit_b[9]), .B(in_17bit_b[7]), .CI(
        add_1_root_r115_carry_13_), .CO(add_1_root_r115_carry_14_), .S(
        add_1_root_r115_SUM_13_) );
  ADDFX2 U117 ( .A(in_17bit_b[13]), .B(in_17bit_b[12]), .CI(
        add_3_root_r119_carry_14_), .CO(add_3_root_r119_carry_15_), .S(
        add_1_root_r119_A_14_) );
  ADDFX2 U118 ( .A(add_1_root_r119_A_13_), .B(in_17bit_b[7]), .CI(
        add_1_root_r119_carry[13]), .CO(add_1_root_r119_carry[14]), .S(
        add_1_root_r119_SUM_13_) );
  ADDFX2 U119 ( .A(in_17bit_b[8]), .B(in_17bit_b[7]), .CI(
        add_2_root_r119_carry_12_), .CO(add_2_root_r119_carry_13_), .S(
        add_2_root_r119_SUM_12_) );
  ADDFX2 U120 ( .A(in_17bit_b[13]), .B(in_17bit_b[9]), .CI(
        add_1_root_r112_carry_13_), .CO(add_1_root_r112_carry_14_), .S(
        add_1_root_r112_SUM_13_) );
  ADDFX2 U121 ( .A(in_17bit_b[10]), .B(in_17bit_b[8]), .CI(
        add_1_root_r115_carry_14_), .CO(add_1_root_r115_carry_15_), .S(
        add_1_root_r115_SUM_14_) );
  ADDFX2 U122 ( .A(in_17bit_b[14]), .B(in_17bit_b[13]), .CI(
        add_3_root_r119_carry_15_), .CO(add_3_root_r119_carry_16_), .S(
        add_1_root_r119_A_15_) );
  ADDFX2 U123 ( .A(add_1_root_r119_A_14_), .B(in_17bit_b[8]), .CI(
        add_1_root_r119_carry[14]), .CO(add_1_root_r119_carry[15]), .S(
        add_1_root_r119_SUM_14_) );
  ADDFX2 U124 ( .A(in_17bit_b[9]), .B(in_17bit_b[8]), .CI(
        add_2_root_r119_carry_13_), .CO(add_2_root_r119_carry_14_), .S(
        add_2_root_r119_SUM_13_) );
  ADDFX2 U125 ( .A(in_17bit_b[12]), .B(in_17bit_b[10]), .CI(
        add_2_root_r115_carry_13_), .CO(add_2_root_r115_carry_14_), .S(
        add_2_root_r115_SUM_13_) );
  ADDFX2 U126 ( .A(in_17bit_b[14]), .B(in_17bit_b[10]), .CI(
        add_1_root_r112_carry_14_), .CO(add_1_root_r112_carry_15_), .S(
        add_1_root_r112_SUM_14_) );
  ADDFX2 U127 ( .A(in_17bit_b[11]), .B(in_17bit_b[9]), .CI(
        add_1_root_r115_carry_15_), .CO(add_1_root_r115_carry_16_), .S(
        add_1_root_r115_SUM_15_) );
  ADDFX2 U128 ( .A(add_1_root_r119_A_15_), .B(in_17bit_b[9]), .CI(
        add_1_root_r119_carry[15]), .CO(add_1_root_r119_carry[16]), .S(
        add_1_root_r119_SUM_15_) );
  ADDFX2 U129 ( .A(in_17bit_b[3]), .B(in_17bit_b[2]), .CI(
        add_3_root_r119_carry_4_), .CO(add_3_root_r119_carry_5_), .S(
        add_1_root_r119_A_4_) );
  ADDFX2 U130 ( .A(in_17bit_b[2]), .B(in_17bit_b[1]), .CI(
        add_3_root_r119_carry_3_), .CO(add_3_root_r119_carry_4_), .S(
        add_1_root_r119_A_3_) );
  ADDFX2 U131 ( .A(in_17bit_b[10]), .B(in_17bit_b[9]), .CI(
        add_2_root_r119_carry_14_), .CO(add_2_root_r119_carry_15_), .S(
        add_2_root_r119_SUM_14_) );
  ADDFX2 U132 ( .A(in_17bit_b[13]), .B(in_17bit_b[11]), .CI(
        add_2_root_r115_carry_14_), .CO(add_2_root_r115_carry_15_), .S(
        add_2_root_r115_SUM_14_) );
  ADDFX2 U133 ( .A(in_17bit_b[15]), .B(in_17bit_b[11]), .CI(
        add_1_root_r112_carry_15_), .CO(add_1_root_r112_carry_16_), .S(
        add_1_root_r112_SUM_15_) );
  ADDFX2 U134 ( .A(in_17bit_b[12]), .B(in_17bit_b[10]), .CI(
        add_1_root_r115_carry_16_), .CO(add_1_root_r115_carry_17_), .S(
        add_1_root_r115_SUM_16_) );
  ADDFX2 U135 ( .A(add_1_root_r119_A_16_), .B(in_17bit_b[10]), .CI(
        add_1_root_r119_carry[16]), .CO(add_1_root_r119_carry[17]), .S(
        add_1_root_r119_SUM_16_) );
  ADDFX2 U136 ( .A(in_17bit_b[11]), .B(in_17bit_b[10]), .CI(
        add_2_root_r119_carry_15_), .CO(add_2_root_r119_carry_16_), .S(
        add_2_root_r119_SUM_15_) );
  ADDFX2 U137 ( .A(in_17bit_b[14]), .B(in_17bit_b[12]), .CI(
        add_2_root_r115_carry_15_), .CO(add_2_root_r115_carry_16_), .S(
        add_2_root_r115_SUM_15_) );
  ADDFX2 U138 ( .A(in_17bit_b[13]), .B(in_17bit_b[11]), .CI(
        add_1_root_r115_carry_17_), .CO(add_1_root_r115_carry_18_), .S(
        add_1_root_r115_SUM_17_) );
  ADDFX2 U139 ( .A(add_1_root_r119_A_17_), .B(in_17bit_b[11]), .CI(
        add_1_root_r119_carry[17]), .CO(add_1_root_r119_carry[18]), .S(
        add_1_root_r119_SUM_17_) );
  ADDFX2 U140 ( .A(in_17bit_b[12]), .B(in_17bit_b[11]), .CI(
        add_2_root_r119_carry_16_), .CO(add_2_root_r119_carry_17_), .S(
        add_2_root_r119_SUM_16_) );
  ADDFX2 U141 ( .A(in_17bit_b[14]), .B(in_17bit_b[12]), .CI(
        add_1_root_r115_carry_18_), .CO(add_1_root_r115_carry_19_), .S(
        add_1_root_r115_SUM_18_) );
  ADDFX2 U142 ( .A(add_1_root_r119_A_18_), .B(in_17bit_b[12]), .CI(
        add_1_root_r119_carry[18]), .CO(add_1_root_r119_carry[19]), .S(
        add_1_root_r119_SUM_18_) );
  ADDFX2 U143 ( .A(in_17bit_b[13]), .B(in_17bit_b[12]), .CI(
        add_2_root_r119_carry_17_), .CO(add_2_root_r119_carry_18_), .S(
        add_2_root_r119_SUM_17_) );
  ADDFX2 U144 ( .A(in_17bit_b[15]), .B(in_17bit_b[13]), .CI(
        add_1_root_r115_carry_19_), .CO(add_1_root_r115_carry_20_), .S(
        add_1_root_r115_SUM_19_) );
  ADDFX2 U145 ( .A(in_17bit_b[5]), .B(in_17bit_b[3]), .CI(
        add_2_root_r115_carry_6_), .CO(add_2_root_r115_carry_7_), .S(
        add_2_root_r115_SUM_6_) );
  ADDFX2 U146 ( .A(in_17bit_b[7]), .B(in_17bit_b[3]), .CI(
        add_1_root_r112_carry_7_), .CO(add_1_root_r112_carry_8_), .S(
        add_1_root_r112_SUM_7_) );
  ADDFX2 U147 ( .A(in_17bit_b[5]), .B(in_17bit_b[3]), .CI(
        add_1_root_r115_carry_9_), .CO(add_1_root_r115_carry_10_), .S(
        add_1_root_r115_SUM_9_) );
  ADDFX2 U148 ( .A(add_1_root_r119_A_9_), .B(in_17bit_b[3]), .CI(
        add_1_root_r119_carry[9]), .CO(add_1_root_r119_carry[10]), .S(
        add_1_root_r119_SUM_9_) );
  ADDFX2 U149 ( .A(in_17bit_b[11]), .B(in_17bit_b[9]), .CI(
        add_2_root_r115_carry_12_), .CO(add_2_root_r115_carry_13_), .S(
        add_2_root_r115_SUM_12_) );
  ADDFX2 U150 ( .A(add_1_root_r119_A_10_), .B(in_17bit_b[4]), .CI(
        add_1_root_r119_carry[10]), .CO(add_1_root_r119_carry[11]), .S(
        add_1_root_r119_SUM_10_) );
  ADDFX2 U151 ( .A(in_17bit_b[8]), .B(in_17bit_b[6]), .CI(
        add_2_root_r115_carry_9_), .CO(add_2_root_r115_carry_10_), .S(
        add_2_root_r115_SUM_9_) );
  ADDFX2 U152 ( .A(in_17bit_b[4]), .B(in_17bit_b[3]), .CI(
        add_2_root_r119_carry_8_), .CO(add_2_root_r119_carry_9_), .S(
        add_2_root_r119_SUM_8_) );
  ADDFX2 U153 ( .A(in_17bit_b[15]), .B(in_17bit_b[14]), .CI(
        add_3_root_r119_carry_16_), .CO(add_3_root_r119_carry_17_), .S(
        add_1_root_r119_A_16_) );
  ADDFX2 U154 ( .A(in_17bit_b[15]), .B(in_17bit_b[13]), .CI(
        add_2_root_r115_carry_16_), .CO(add_2_root_r115_carry_17_), .S(
        add_2_root_r115_SUM_16_) );
  ADDFX2 U155 ( .A(in_17bit_b[4]), .B(in_17bit_b[3]), .CI(
        add_3_root_r119_carry_5_), .CO(add_3_root_r119_carry_6_), .S(
        add_1_root_r119_A_5_) );
  ADDFX2 U156 ( .A(in_17bit_b[5]), .B(in_17bit_b[4]), .CI(
        add_3_root_r119_carry_6_), .CO(add_3_root_r119_carry_7_), .S(
        add_1_root_r119_A_6_) );
  ADDFX2 U157 ( .A(in_17bit_b[14]), .B(in_17bit_b[13]), .CI(
        add_2_root_r119_carry_18_), .CO(add_2_root_r119_carry_19_), .S(
        add_2_root_r119_SUM_18_) );
  ADDFX2 U158 ( .A(in_17bit_b[15]), .B(in_17bit_b[14]), .CI(
        add_2_root_r119_carry_19_), .CO(add_2_root_r119_carry_20_), .S(
        add_2_root_r119_SUM_19_) );
  INVX1 U159 ( .A(n197), .Y(n95) );
  NAND3BX1 U160 ( .AN(in_8bit[5]), .B(n50), .C(in_8bit[3]), .Y(n197) );
  INVX1 U161 ( .A(in_8bit[3]), .Y(n51) );
  CLKINVX3 U162 ( .A(n202), .Y(in_17bit_b[0]) );
  INVX1 U163 ( .A(n175), .Y(n254) );
  NAND2XL U164 ( .A(N29), .B(n61), .Y(n255) );
  INVX1 U165 ( .A(n77), .Y(n81) );
  OAI21XL U166 ( .A0(n254), .A1(n255), .B0(n253), .Y(N463) );
  AOI22X1 U167 ( .A0(N221), .A1(n49), .B0(N363), .B1(n48), .Y(n253) );
  CLKINVX3 U168 ( .A(n247), .Y(in_17bit_b[15]) );
  INVX1 U169 ( .A(in_8bit[2]), .Y(n50) );
  INVX1 U170 ( .A(in_8bit[5]), .Y(n57) );
  XNOR2X4 U171 ( .A(n34), .B(n5), .Y(n33) );
  MXI2XL U172 ( .A(n4), .B(n17), .S0(n87), .Y(out[16]) );
  AOI22XL U173 ( .A0(in_17bit[0]), .A1(n61), .B0(in_17bit[0]), .B1(n62), .Y(
        n202) );
  AOI22XL U174 ( .A0(N28), .A1(n61), .B0(in_17bit[15]), .B1(n62), .Y(n247) );
  AOI22XL U175 ( .A0(N22), .A1(n61), .B0(in_17bit[9]), .B1(n62), .Y(n229) );
  AOI22XL U176 ( .A0(N24), .A1(n61), .B0(in_17bit[11]), .B1(n62), .Y(n235) );
  AOI22XL U177 ( .A0(N25), .A1(n61), .B0(in_17bit[12]), .B1(n62), .Y(n238) );
  AOI22XL U178 ( .A0(N26), .A1(n61), .B0(in_17bit[13]), .B1(n62), .Y(n241) );
  AOI22XL U179 ( .A0(N14), .A1(n61), .B0(in_17bit[1]), .B1(n62), .Y(n205) );
  AOI22XL U180 ( .A0(N15), .A1(n61), .B0(in_17bit[2]), .B1(n62), .Y(n208) );
  AOI22XL U181 ( .A0(N16), .A1(n61), .B0(in_17bit[3]), .B1(n62), .Y(n211) );
  AOI22XL U182 ( .A0(N17), .A1(n61), .B0(in_17bit[4]), .B1(n62), .Y(n214) );
  AOI22XL U183 ( .A0(N18), .A1(n61), .B0(in_17bit[5]), .B1(n62), .Y(n217) );
  AOI22XL U184 ( .A0(N19), .A1(n61), .B0(in_17bit[6]), .B1(n62), .Y(n220) );
  AOI22XL U185 ( .A0(N20), .A1(n61), .B0(in_17bit[7]), .B1(n62), .Y(n223) );
  AOI22XL U186 ( .A0(N21), .A1(n61), .B0(in_17bit[8]), .B1(n62), .Y(n226) );
  AOI22XL U187 ( .A0(N23), .A1(n61), .B0(in_17bit[10]), .B1(n62), .Y(n232) );
  INVX1 U188 ( .A(n64), .Y(n71) );
  NAND2BX1 U189 ( .AN(n69), .B(n18), .Y(n64) );
  AND2X2 U190 ( .A(n38), .B(n7), .Y(n36) );
  AND2X2 U191 ( .A(n71), .B(n15), .Y(n37) );
  AND2X2 U192 ( .A(n81), .B(n6), .Y(n38) );
  AND2X2 U193 ( .A(n36), .B(n8), .Y(n39) );
  AND2X2 U194 ( .A(n39), .B(n16), .Y(n40) );
  BUFX3 U195 ( .A(n251), .Y(n48) );
  OAI2BB1X1 U196 ( .A0N(n95), .A1N(n31), .B0(n93), .Y(n251) );
  NAND2BX1 U197 ( .AN(n196), .B(n42), .Y(n93) );
  BUFX3 U198 ( .A(n252), .Y(n49) );
  OAI2BB1X1 U199 ( .A0N(n42), .A1N(n95), .B0(n94), .Y(n252) );
  NAND2BX1 U200 ( .AN(n196), .B(n31), .Y(n94) );
  AND2X2 U201 ( .A(n37), .B(n3), .Y(n41) );
  NAND2X1 U202 ( .A(n41), .B(n9), .Y(n77) );
  OAI2BB1X1 U203 ( .A0N(n199), .A1N(n32), .B0(n97), .Y(n175) );
  NAND3BX1 U204 ( .AN(n96), .B(n200), .C(in_8bit[5]), .Y(n97) );
  NAND2X1 U205 ( .A(n45), .B(n12), .Y(n69) );
  AND2X2 U206 ( .A(n92), .B(n53), .Y(n42) );
  AND2X2 U207 ( .A(n40), .B(n5), .Y(n43) );
  INVX1 U208 ( .A(in_17bit[0]), .Y(n98) );
  INVX1 U209 ( .A(in_17bit[1]), .Y(n99) );
  INVX1 U210 ( .A(in_17bit[2]), .Y(n100) );
  INVX1 U211 ( .A(in_17bit[3]), .Y(n101) );
  INVX1 U212 ( .A(in_17bit[4]), .Y(n158) );
  INVX1 U213 ( .A(in_17bit[5]), .Y(n160) );
  INVX1 U214 ( .A(in_17bit[6]), .Y(n161) );
  INVX1 U215 ( .A(in_17bit[7]), .Y(n162) );
  INVX1 U216 ( .A(in_17bit[8]), .Y(n163) );
  INVX1 U217 ( .A(in_17bit[9]), .Y(n164) );
  INVX1 U218 ( .A(in_17bit[10]), .Y(n168) );
  INVX1 U219 ( .A(in_17bit[11]), .Y(n170) );
  INVX1 U220 ( .A(in_17bit[12]), .Y(n171) );
  INVX1 U221 ( .A(in_17bit[13]), .Y(n172) );
  INVX1 U222 ( .A(in_17bit[14]), .Y(n173) );
  INVX1 U223 ( .A(in_17bit[15]), .Y(n174) );
  NAND2X1 U224 ( .A(n204), .B(n203), .Y(N447) );
  AOI22X1 U225 ( .A0(N108), .A1(n248), .B0(N205), .B1(n49), .Y(n203) );
  AOI22X1 U226 ( .A0(N347), .A1(n48), .B0(n175), .B1(in_17bit_b[0]), .Y(n204)
         );
  NAND2X1 U227 ( .A(n207), .B(n206), .Y(N448) );
  AOI22X1 U228 ( .A0(N109), .A1(n248), .B0(N206), .B1(n49), .Y(n206) );
  AOI22X1 U229 ( .A0(N348), .A1(n48), .B0(n175), .B1(in_17bit_b[1]), .Y(n207)
         );
  NAND2X1 U230 ( .A(n210), .B(n209), .Y(N449) );
  AOI22X1 U231 ( .A0(N110), .A1(n248), .B0(N207), .B1(n49), .Y(n209) );
  AOI22X1 U232 ( .A0(N349), .A1(n48), .B0(n175), .B1(in_17bit_b[2]), .Y(n210)
         );
  NAND2X1 U233 ( .A(n213), .B(n212), .Y(N450) );
  AOI22X1 U234 ( .A0(N111), .A1(n248), .B0(N208), .B1(n49), .Y(n212) );
  AOI22X1 U235 ( .A0(N350), .A1(n48), .B0(n175), .B1(in_17bit_b[3]), .Y(n213)
         );
  NAND2X1 U236 ( .A(n216), .B(n215), .Y(N451) );
  AOI22X1 U237 ( .A0(N112), .A1(n248), .B0(N209), .B1(n49), .Y(n215) );
  AOI22X1 U238 ( .A0(N351), .A1(n48), .B0(n175), .B1(in_17bit_b[4]), .Y(n216)
         );
  NAND2X1 U239 ( .A(n219), .B(n218), .Y(N452) );
  AOI22X1 U240 ( .A0(N113), .A1(n248), .B0(N210), .B1(n49), .Y(n218) );
  AOI22X1 U241 ( .A0(N352), .A1(n48), .B0(n175), .B1(in_17bit_b[5]), .Y(n219)
         );
  NAND2X1 U242 ( .A(n222), .B(n221), .Y(N453) );
  AOI22X1 U243 ( .A0(N114), .A1(n248), .B0(N211), .B1(n49), .Y(n221) );
  AOI22X1 U244 ( .A0(N353), .A1(n48), .B0(n175), .B1(in_17bit_b[6]), .Y(n222)
         );
  NAND2X1 U245 ( .A(n225), .B(n224), .Y(N454) );
  AOI22X1 U246 ( .A0(N115), .A1(n248), .B0(N212), .B1(n49), .Y(n224) );
  AOI22X1 U247 ( .A0(N354), .A1(n48), .B0(n175), .B1(in_17bit_b[7]), .Y(n225)
         );
  NAND2X1 U248 ( .A(n228), .B(n227), .Y(N455) );
  AOI22X1 U249 ( .A0(N116), .A1(n248), .B0(N213), .B1(n49), .Y(n227) );
  AOI22X1 U250 ( .A0(N355), .A1(n48), .B0(n175), .B1(in_17bit_b[8]), .Y(n228)
         );
  NAND2X1 U251 ( .A(n231), .B(n230), .Y(N456) );
  AOI22X1 U252 ( .A0(N117), .A1(n248), .B0(N214), .B1(n49), .Y(n230) );
  AOI22X1 U253 ( .A0(N356), .A1(n48), .B0(n175), .B1(in_17bit_b[9]), .Y(n231)
         );
  NAND2X1 U254 ( .A(n234), .B(n233), .Y(N457) );
  AOI22X1 U255 ( .A0(N118), .A1(n248), .B0(N215), .B1(n49), .Y(n233) );
  AOI22X1 U256 ( .A0(N357), .A1(n48), .B0(n175), .B1(in_17bit_b[10]), .Y(n234)
         );
  NAND2X1 U257 ( .A(n237), .B(n236), .Y(N458) );
  AOI22X1 U258 ( .A0(N119), .A1(n248), .B0(N216), .B1(n49), .Y(n236) );
  AOI22X1 U259 ( .A0(N358), .A1(n48), .B0(n175), .B1(in_17bit_b[11]), .Y(n237)
         );
  NAND2X1 U260 ( .A(n240), .B(n239), .Y(N459) );
  AOI22X1 U261 ( .A0(N120), .A1(n248), .B0(N217), .B1(n49), .Y(n239) );
  AOI22X1 U262 ( .A0(N359), .A1(n48), .B0(n175), .B1(in_17bit_b[12]), .Y(n240)
         );
  NAND2X1 U263 ( .A(n243), .B(n242), .Y(N460) );
  AOI22X1 U264 ( .A0(N121), .A1(n248), .B0(N218), .B1(n49), .Y(n242) );
  AOI22X1 U265 ( .A0(N360), .A1(n48), .B0(n175), .B1(in_17bit_b[13]), .Y(n243)
         );
  NAND2X1 U266 ( .A(n246), .B(n245), .Y(N461) );
  AOI22X1 U267 ( .A0(N122), .A1(n248), .B0(N219), .B1(n49), .Y(n245) );
  AOI22X1 U268 ( .A0(N361), .A1(n48), .B0(n175), .B1(in_17bit_b[14]), .Y(n246)
         );
  NAND2X1 U269 ( .A(n250), .B(n249), .Y(N462) );
  AOI22X1 U270 ( .A0(N123), .A1(n248), .B0(N220), .B1(n49), .Y(n249) );
  AOI22X1 U271 ( .A0(N362), .A1(n48), .B0(n175), .B1(in_17bit_b[15]), .Y(n250)
         );
  XNOR2X1 U272 ( .A(n13), .B(sub_add_75_b0_carry[13]), .Y(n44) );
  INVX1 U273 ( .A(n76), .Y(n75) );
  MX2X1 U274 ( .A(neg_mul[22]), .B(N480), .S0(n87), .Y(out[15]) );
  NAND4BBX1 U275 ( .AN(n48), .BN(n49), .C(n201), .D(n254), .Y(N446) );
  NOR4BX1 U276 ( .AN(n198), .B(n53), .C(n54), .D(in_8bit[2]), .Y(n199) );
  NOR2X1 U277 ( .A(in_8bit[6]), .B(in_8bit[3]), .Y(n198) );
  NAND4BXL U278 ( .AN(n55), .B(in_8bit[6]), .C(n54), .D(in_8bit[4]), .Y(n96)
         );
  NOR2X1 U279 ( .A(out[0]), .B(neg_mul[8]), .Y(n45) );
  NOR2X1 U280 ( .A(in_8bit[6]), .B(in_8bit[4]), .Y(n195) );
  NAND2X1 U281 ( .A(n91), .B(n90), .Y(n248) );
  NAND3BX1 U282 ( .AN(n88), .B(n200), .C(in_8bit[6]), .Y(n91) );
  NAND3X1 U283 ( .A(n199), .B(in_8bit[5]), .C(n89), .Y(n90) );
  NAND2BX1 U284 ( .AN(n41), .B(neg_mul[13]), .Y(n76) );
  NAND2X1 U285 ( .A(sub_add_75_b0_carry[15]), .B(n11), .Y(n46) );
  XNOR2X4 U286 ( .A(n25), .B(n59), .Y(n73) );
  NOR2X4 U287 ( .A(n73), .B(n37), .Y(n74) );
  AOI2BB1X4 U288 ( .A0N(n23), .A1N(n80), .B0(n79), .Y(out[6]) );
  XNOR2X4 U289 ( .A(n82), .B(n6), .Y(out[7]) );
  XNOR2X4 U290 ( .A(n83), .B(n7), .Y(out[8]) );
  XNOR2X4 U291 ( .A(n84), .B(n8), .Y(out[9]) );
  AND2X1 U292 ( .A(add_1_root_r112_carry_20_), .B(in_17bit_b[16]), .Y(
        add_1_root_r112_SUM_21_) );
  XOR2X1 U293 ( .A(in_17bit_b[16]), .B(add_1_root_r112_carry_20_), .Y(
        add_1_root_r112_SUM_20_) );
  AND2X1 U294 ( .A(add_1_root_r112_carry_19_), .B(in_17bit_b[15]), .Y(
        add_1_root_r112_carry_20_) );
  XOR2X1 U295 ( .A(in_17bit_b[15]), .B(add_1_root_r112_carry_19_), .Y(
        add_1_root_r112_SUM_19_) );
  AND2X1 U296 ( .A(add_1_root_r112_carry_18_), .B(in_17bit_b[14]), .Y(
        add_1_root_r112_carry_19_) );
  XOR2X1 U297 ( .A(in_17bit_b[14]), .B(add_1_root_r112_carry_18_), .Y(
        add_1_root_r112_SUM_18_) );
  AND2X1 U298 ( .A(add_1_root_r112_carry_17_), .B(in_17bit_b[13]), .Y(
        add_1_root_r112_carry_18_) );
  XOR2X1 U299 ( .A(in_17bit_b[13]), .B(add_1_root_r112_carry_17_), .Y(
        add_1_root_r112_SUM_17_) );
  AND2X1 U300 ( .A(add_2_root_r119_carry_21_), .B(in_17bit_b[16]), .Y(
        add_2_root_r119_SUM_22_) );
  XOR2X1 U301 ( .A(in_17bit_b[16]), .B(add_2_root_r119_carry_21_), .Y(
        add_2_root_r119_SUM_21_) );
  AND2X1 U302 ( .A(add_1_root_r119_carry[22]), .B(in_17bit_b[16]), .Y(
        add_1_root_r119_SUM_23_) );
  XOR2X1 U303 ( .A(in_17bit_b[16]), .B(add_1_root_r119_carry[22]), .Y(
        add_1_root_r119_SUM_22_) );
  AND2X1 U304 ( .A(add_1_root_r119_carry[21]), .B(in_17bit_b[15]), .Y(
        add_1_root_r119_carry[22]) );
  XOR2X1 U305 ( .A(in_17bit_b[15]), .B(add_1_root_r119_carry[21]), .Y(
        add_1_root_r119_SUM_21_) );
  AND2X1 U306 ( .A(add_1_root_r119_carry[20]), .B(in_17bit_b[14]), .Y(
        add_1_root_r119_carry[21]) );
  XOR2X1 U307 ( .A(in_17bit_b[14]), .B(add_1_root_r119_carry[20]), .Y(
        add_1_root_r119_SUM_20_) );
  AND2X1 U308 ( .A(add_1_root_r119_A_6_), .B(in_17bit_b[0]), .Y(
        add_1_root_r119_carry[7]) );
  XOR2X1 U309 ( .A(in_17bit_b[0]), .B(add_1_root_r119_A_6_), .Y(
        add_1_root_r119_SUM_6_) );
  AND2X1 U310 ( .A(add_3_root_r119_carry_18_), .B(in_17bit_b[16]), .Y(
        add_1_root_r119_A_19_) );
  XOR2X1 U311 ( .A(in_17bit_b[16]), .B(add_3_root_r119_carry_18_), .Y(
        add_1_root_r119_A_18_) );
  AND2X1 U312 ( .A(in_17bit_b[1]), .B(in_17bit_b[0]), .Y(
        add_3_root_r119_carry_3_) );
  XOR2X1 U313 ( .A(in_17bit_b[0]), .B(in_17bit_b[1]), .Y(add_1_root_r119_A_2_)
         );
  AND2X1 U314 ( .A(add_2_root_r115_carry_19_), .B(in_17bit_b[16]), .Y(
        add_2_root_r115_SUM_20_) );
  XOR2X1 U315 ( .A(in_17bit_b[16]), .B(add_2_root_r115_carry_19_), .Y(
        add_2_root_r115_SUM_19_) );
  AND2X1 U316 ( .A(add_2_root_r115_carry_18_), .B(in_17bit_b[15]), .Y(
        add_2_root_r115_carry_19_) );
  XOR2X1 U317 ( .A(in_17bit_b[15]), .B(add_2_root_r115_carry_18_), .Y(
        add_2_root_r115_SUM_18_) );
  AND2X1 U318 ( .A(add_1_root_r115_carry_22_), .B(in_17bit_b[16]), .Y(
        add_1_root_r115_SUM_23_) );
  XOR2X1 U319 ( .A(in_17bit_b[16]), .B(add_1_root_r115_carry_22_), .Y(
        add_1_root_r115_SUM_22_) );
  AND2X1 U320 ( .A(add_1_root_r115_carry_21_), .B(in_17bit_b[15]), .Y(
        add_1_root_r115_carry_22_) );
  XOR2X1 U321 ( .A(in_17bit_b[15]), .B(add_1_root_r115_carry_21_), .Y(
        add_1_root_r115_SUM_21_) );
  AND2X1 U322 ( .A(in_17bit_b[2]), .B(in_17bit_b[0]), .Y(
        add_1_root_r115_carry_7_) );
  XOR2X1 U323 ( .A(in_17bit_b[0]), .B(in_17bit_b[2]), .Y(
        add_1_root_r115_SUM_6_) );
  XOR2X1 U324 ( .A(n63), .B(sub_add_54_b0_carry[16]), .Y(N29) );
  AND2X1 U325 ( .A(sub_add_54_b0_carry[15]), .B(n174), .Y(
        sub_add_54_b0_carry[16]) );
  XOR2X1 U326 ( .A(n174), .B(sub_add_54_b0_carry[15]), .Y(N28) );
  AND2X1 U327 ( .A(sub_add_54_b0_carry[14]), .B(n173), .Y(
        sub_add_54_b0_carry[15]) );
  XOR2X1 U328 ( .A(n173), .B(sub_add_54_b0_carry[14]), .Y(N27) );
  AND2X1 U329 ( .A(sub_add_54_b0_carry[13]), .B(n172), .Y(
        sub_add_54_b0_carry[14]) );
  XOR2X1 U330 ( .A(n172), .B(sub_add_54_b0_carry[13]), .Y(N26) );
  AND2X1 U331 ( .A(sub_add_54_b0_carry[12]), .B(n171), .Y(
        sub_add_54_b0_carry[13]) );
  XOR2X1 U332 ( .A(n171), .B(sub_add_54_b0_carry[12]), .Y(N25) );
  AND2X1 U333 ( .A(sub_add_54_b0_carry[11]), .B(n170), .Y(
        sub_add_54_b0_carry[12]) );
  XOR2X1 U334 ( .A(n170), .B(sub_add_54_b0_carry[11]), .Y(N24) );
  AND2X1 U335 ( .A(sub_add_54_b0_carry[10]), .B(n168), .Y(
        sub_add_54_b0_carry[11]) );
  XOR2X1 U336 ( .A(n168), .B(sub_add_54_b0_carry[10]), .Y(N23) );
  AND2X1 U337 ( .A(sub_add_54_b0_carry[9]), .B(n164), .Y(
        sub_add_54_b0_carry[10]) );
  XOR2X1 U338 ( .A(n164), .B(sub_add_54_b0_carry[9]), .Y(N22) );
  AND2X1 U339 ( .A(sub_add_54_b0_carry[8]), .B(n163), .Y(
        sub_add_54_b0_carry[9]) );
  XOR2X1 U340 ( .A(n163), .B(sub_add_54_b0_carry[8]), .Y(N21) );
  AND2X1 U341 ( .A(sub_add_54_b0_carry[7]), .B(n162), .Y(
        sub_add_54_b0_carry[8]) );
  XOR2X1 U342 ( .A(n162), .B(sub_add_54_b0_carry[7]), .Y(N20) );
  AND2X1 U343 ( .A(sub_add_54_b0_carry[6]), .B(n161), .Y(
        sub_add_54_b0_carry[7]) );
  XOR2X1 U344 ( .A(n161), .B(sub_add_54_b0_carry[6]), .Y(N19) );
  AND2X1 U345 ( .A(sub_add_54_b0_carry[5]), .B(n160), .Y(
        sub_add_54_b0_carry[6]) );
  XOR2X1 U346 ( .A(n160), .B(sub_add_54_b0_carry[5]), .Y(N18) );
  AND2X1 U347 ( .A(sub_add_54_b0_carry[4]), .B(n158), .Y(
        sub_add_54_b0_carry[5]) );
  XOR2X1 U348 ( .A(n158), .B(sub_add_54_b0_carry[4]), .Y(N17) );
  AND2X1 U349 ( .A(sub_add_54_b0_carry[3]), .B(n101), .Y(
        sub_add_54_b0_carry[4]) );
  XOR2X1 U350 ( .A(n101), .B(sub_add_54_b0_carry[3]), .Y(N16) );
  AND2X1 U351 ( .A(sub_add_54_b0_carry[2]), .B(n100), .Y(
        sub_add_54_b0_carry[3]) );
  XOR2X1 U352 ( .A(n100), .B(sub_add_54_b0_carry[2]), .Y(N15) );
  AND2X1 U353 ( .A(n98), .B(n99), .Y(sub_add_54_b0_carry[2]) );
  XOR2X1 U354 ( .A(n99), .B(n98), .Y(N14) );
  XOR2X1 U355 ( .A(n11), .B(sub_add_75_b0_carry[15]), .Y(N480) );
  AND2X1 U356 ( .A(sub_add_75_b0_carry[14]), .B(n28), .Y(
        sub_add_75_b0_carry[15]) );
  AND2X1 U357 ( .A(sub_add_75_b0_carry[13]), .B(n13), .Y(
        sub_add_75_b0_carry[14]) );
  AND2X1 U358 ( .A(n43), .B(n10), .Y(sub_add_75_b0_carry[13]) );
  AND2X1 U359 ( .A(in_17bit_b[0]), .B(in_17bit_b[4]), .Y(
        add_1_root_r112_carry_5_) );
endmodule


module multi16_2_DW01_add_0 ( A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, 
        A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, 
        A_4_, B_23_, B_22_, B_21_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, 
        B_14_, B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, 
        SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, 
        SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, 
        SUM_7_ );
  input A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_,
         A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, B_23_, B_22_,
         B_21_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_,
         B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_;
  output SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_,
         SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_,
         SUM_8_, SUM_7_;
  wire   n1, n2, n3, n4;
  wire   [23:7] carry;

  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry[7]), .CO(carry[8]), .S(SUM_7_)
         );
  ADDFX2 U1_21 ( .A(A_21_), .B(B_21_), .CI(carry[21]), .CO(carry[22]), .S(
        SUM_21_) );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry[20]), .CO(carry[21]), .S(
        SUM_20_) );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry[19]), .CO(carry[20]), .S(
        SUM_19_) );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry[18]), .CO(carry[19]), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry[17]), .CO(carry[18]), .S(
        SUM_17_) );
  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry[16]), .CO(carry[17]), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry[15]), .CO(carry[16]), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry[14]), .CO(carry[15]), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry[13]), .CO(carry[14]), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry[12]), .CO(carry[13]), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry[11]), .CO(carry[12]), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry[10]), .CO(carry[11]), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry[9]), .CO(carry[10]), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry[8]), .CO(carry[9]), .S(SUM_8_)
         );
  ADDFX2 U1_22 ( .A(A_22_), .B(B_22_), .CI(carry[22]), .CO(carry[23]), .S(
        SUM_22_) );
  AND2X2 U1 ( .A(A_4_), .B(B_4_), .Y(n1) );
  XOR2X1 U2 ( .A(B_23_), .B(carry[23]), .Y(SUM_23_) );
  OAI2BB1X1 U3 ( .A0N(n2), .A1N(A_6_), .B0(n3), .Y(carry[7]) );
  OAI21XL U4 ( .A0(A_6_), .A1(n2), .B0(B_6_), .Y(n3) );
  OAI2BB1X1 U5 ( .A0N(n1), .A1N(A_5_), .B0(n4), .Y(n2) );
  OAI21XL U6 ( .A0(A_5_), .A1(n1), .B0(B_5_), .Y(n4) );
endmodule


module multi16_2_DW01_add_4 ( A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, 
        A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, 
        B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, 
        B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, SUM_22_, SUM_21_, SUM_20_, 
        SUM_19_, SUM_18_, SUM_17_, SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, 
        SUM_11_, SUM_10_, SUM_9_, SUM_8_, SUM_7_ );
  input A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_,
         A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, B_20_, B_19_,
         B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, B_10_, B_9_,
         B_8_, B_7_, B_6_, B_5_;
  output SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_,
         SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_,
         SUM_7_;
  wire   carry_21_, carry_20_, carry_19_, carry_18_, carry_17_, carry_16_,
         carry_15_, carry_14_, carry_13_, carry_12_, carry_11_, carry_10_,
         carry_9_, carry_8_, carry_7_, n1;

  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry_16_), .CO(carry_17_), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry_15_), .CO(carry_16_), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry_14_), .CO(carry_15_), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry_13_), .CO(carry_14_), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry_12_), .CO(carry_13_), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry_11_), .CO(carry_12_), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry_10_), .CO(carry_11_), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry_9_), .CO(carry_10_), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry_8_), .CO(carry_9_), .S(SUM_8_)
         );
  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry_7_), .CO(carry_8_), .S(SUM_7_)
         );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry_20_), .CO(carry_21_), .S(
        SUM_20_) );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry_19_), .CO(carry_20_), .S(
        SUM_19_) );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry_18_), .CO(carry_19_), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry_17_), .CO(carry_18_), .S(
        SUM_17_) );
  ADDFX2 U1_21 ( .A(A_21_), .B(B_21_), .CI(carry_21_), .CO(SUM_22_), .S(
        SUM_21_) );
  OAI2BB1X1 U1 ( .A0N(A_6_), .A1N(B_6_), .B0(n1), .Y(carry_7_) );
  OAI211X1 U2 ( .A0(B_6_), .A1(A_6_), .B0(A_5_), .C0(B_5_), .Y(n1) );
endmodule


module multi16_2_DW01_add_6 ( A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, 
        A_16_, A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, 
        A_6_, A_5_, A_4_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, 
        B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, 
        SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, 
        SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, 
        SUM_7_ );
  input A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_,
         A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, B_20_,
         B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, B_10_,
         B_9_, B_8_, B_7_, B_6_, B_5_, B_4_;
  output SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_,
         SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_,
         SUM_8_, SUM_7_;
  wire   n1, n2, n3, n4, n5, n6;
  wire   [21:7] carry;

  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry[7]), .CO(carry[8]), .S(SUM_7_)
         );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry[18]), .CO(carry[19]), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry[17]), .CO(carry[18]), .S(
        SUM_17_) );
  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry[16]), .CO(carry[17]), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry[15]), .CO(carry[16]), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry[14]), .CO(carry[15]), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry[13]), .CO(carry[14]), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry[12]), .CO(carry[13]), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry[11]), .CO(carry[12]), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry[10]), .CO(carry[11]), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry[9]), .CO(carry[10]), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry[8]), .CO(carry[9]), .S(SUM_8_)
         );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry[19]), .CO(carry[20]), .S(
        SUM_19_) );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry[20]), .CO(carry[21]), .S(
        SUM_20_) );
  AND2X2 U1 ( .A(A_22_), .B(n2), .Y(n1) );
  AND2X2 U2 ( .A(A_21_), .B(carry[21]), .Y(n2) );
  AND2X2 U3 ( .A(A_4_), .B(B_4_), .Y(n3) );
  XOR2X1 U4 ( .A(A_23_), .B(n1), .Y(SUM_23_) );
  XOR2X1 U5 ( .A(A_21_), .B(carry[21]), .Y(SUM_21_) );
  XOR2X1 U6 ( .A(A_22_), .B(n2), .Y(SUM_22_) );
  OAI2BB1X1 U7 ( .A0N(n4), .A1N(A_6_), .B0(n5), .Y(carry[7]) );
  OAI21XL U8 ( .A0(A_6_), .A1(n4), .B0(B_6_), .Y(n5) );
  OAI2BB1X1 U9 ( .A0N(n3), .A1N(A_5_), .B0(n6), .Y(n4) );
  OAI21XL U10 ( .A0(A_5_), .A1(n3), .B0(B_5_), .Y(n6) );
endmodule


module multi16_2 ( in_17bit, in_8bit, out );
  input [16:0] in_17bit;
  input [7:0] in_8bit;
  output [16:0] out;
  wire   n269, n270, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24,
         N25, N26, N27, N28, N29, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, N205, N206,
         N207, N208, N209, N210, N211, N212, N213, N214, N215, N216, N217,
         N218, N219, N220, N221, N347, N348, N349, N350, N351, N352, N353,
         N354, N355, N356, N357, N358, N359, N360, N361, N362, N363, N446,
         N447, N448, N449, N450, N451, N452, N453, N454, N455, N456, N457,
         N458, N459, N460, N461, N462, N463, N480, N481,
         add_2_root_r119_carry_10_, add_2_root_r119_carry_11_,
         add_2_root_r119_carry_12_, add_2_root_r119_carry_13_,
         add_2_root_r119_carry_14_, add_2_root_r119_carry_15_,
         add_2_root_r119_carry_16_, add_2_root_r119_carry_17_,
         add_2_root_r119_carry_18_, add_2_root_r119_carry_19_,
         add_2_root_r119_carry_20_, add_2_root_r119_carry_21_,
         add_2_root_r119_carry_7_, add_2_root_r119_carry_8_,
         add_2_root_r119_carry_9_, add_2_root_r119_SUM_6_,
         add_2_root_r119_SUM_7_, add_2_root_r119_SUM_8_,
         add_2_root_r119_SUM_9_, add_2_root_r119_SUM_10_,
         add_2_root_r119_SUM_11_, add_2_root_r119_SUM_12_,
         add_2_root_r119_SUM_13_, add_2_root_r119_SUM_14_,
         add_2_root_r119_SUM_15_, add_2_root_r119_SUM_16_,
         add_2_root_r119_SUM_17_, add_2_root_r119_SUM_18_,
         add_2_root_r119_SUM_19_, add_2_root_r119_SUM_20_,
         add_2_root_r119_SUM_21_, add_2_root_r119_SUM_22_,
         add_1_root_r119_SUM_6_, add_1_root_r119_SUM_7_,
         add_1_root_r119_SUM_8_, add_1_root_r119_SUM_9_,
         add_1_root_r119_SUM_10_, add_1_root_r119_SUM_11_,
         add_1_root_r119_SUM_12_, add_1_root_r119_SUM_13_,
         add_1_root_r119_SUM_14_, add_1_root_r119_SUM_15_,
         add_1_root_r119_SUM_16_, add_1_root_r119_SUM_17_,
         add_1_root_r119_SUM_18_, add_1_root_r119_SUM_19_,
         add_1_root_r119_SUM_20_, add_1_root_r119_SUM_21_,
         add_1_root_r119_SUM_22_, add_1_root_r119_SUM_23_,
         add_1_root_r119_A_2_, add_1_root_r119_A_3_, add_1_root_r119_A_4_,
         add_1_root_r119_A_5_, add_1_root_r119_A_6_, add_1_root_r119_A_7_,
         add_1_root_r119_A_8_, add_1_root_r119_A_9_, add_1_root_r119_A_10_,
         add_1_root_r119_A_11_, add_1_root_r119_A_12_, add_1_root_r119_A_13_,
         add_1_root_r119_A_14_, add_1_root_r119_A_15_, add_1_root_r119_A_16_,
         add_1_root_r119_A_17_, add_1_root_r119_A_18_, add_1_root_r119_A_19_,
         add_3_root_r119_carry_10_, add_3_root_r119_carry_11_,
         add_3_root_r119_carry_12_, add_3_root_r119_carry_13_,
         add_3_root_r119_carry_14_, add_3_root_r119_carry_15_,
         add_3_root_r119_carry_16_, add_3_root_r119_carry_17_,
         add_3_root_r119_carry_18_, add_3_root_r119_carry_3_,
         add_3_root_r119_carry_4_, add_3_root_r119_carry_5_,
         add_3_root_r119_carry_6_, add_3_root_r119_carry_7_,
         add_3_root_r119_carry_8_, add_3_root_r119_carry_9_,
         add_1_root_r112_carry_10_, add_1_root_r112_carry_11_,
         add_1_root_r112_carry_12_, add_1_root_r112_carry_13_,
         add_1_root_r112_carry_14_, add_1_root_r112_carry_15_,
         add_1_root_r112_carry_16_, add_1_root_r112_carry_17_,
         add_1_root_r112_carry_18_, add_1_root_r112_carry_19_,
         add_1_root_r112_carry_20_, add_1_root_r112_carry_5_,
         add_1_root_r112_carry_6_, add_1_root_r112_carry_7_,
         add_1_root_r112_carry_8_, add_1_root_r112_carry_9_,
         add_1_root_r112_SUM_1_, add_1_root_r112_SUM_2_,
         add_1_root_r112_SUM_3_, add_1_root_r112_SUM_4_,
         add_1_root_r112_SUM_5_, add_1_root_r112_SUM_6_,
         add_1_root_r112_SUM_7_, add_1_root_r112_SUM_8_,
         add_1_root_r112_SUM_9_, add_1_root_r112_SUM_10_,
         add_1_root_r112_SUM_11_, add_1_root_r112_SUM_12_,
         add_1_root_r112_SUM_13_, add_1_root_r112_SUM_14_,
         add_1_root_r112_SUM_15_, add_1_root_r112_SUM_16_,
         add_1_root_r112_SUM_17_, add_1_root_r112_SUM_18_,
         add_1_root_r112_SUM_19_, add_1_root_r112_SUM_20_,
         add_1_root_r112_SUM_21_, add_2_root_r115_carry_10_,
         add_2_root_r115_carry_11_, add_2_root_r115_carry_12_,
         add_2_root_r115_carry_13_, add_2_root_r115_carry_14_,
         add_2_root_r115_carry_15_, add_2_root_r115_carry_16_,
         add_2_root_r115_carry_17_, add_2_root_r115_carry_18_,
         add_2_root_r115_carry_19_, add_2_root_r115_carry_5_,
         add_2_root_r115_carry_6_, add_2_root_r115_carry_7_,
         add_2_root_r115_carry_8_, add_2_root_r115_carry_9_,
         add_2_root_r115_SUM_4_, add_2_root_r115_SUM_5_,
         add_2_root_r115_SUM_6_, add_2_root_r115_SUM_7_,
         add_2_root_r115_SUM_8_, add_2_root_r115_SUM_9_,
         add_2_root_r115_SUM_10_, add_2_root_r115_SUM_11_,
         add_2_root_r115_SUM_12_, add_2_root_r115_SUM_13_,
         add_2_root_r115_SUM_14_, add_2_root_r115_SUM_15_,
         add_2_root_r115_SUM_16_, add_2_root_r115_SUM_17_,
         add_2_root_r115_SUM_18_, add_2_root_r115_SUM_19_,
         add_2_root_r115_SUM_20_, add_1_root_r115_carry_10_,
         add_1_root_r115_carry_11_, add_1_root_r115_carry_12_,
         add_1_root_r115_carry_13_, add_1_root_r115_carry_14_,
         add_1_root_r115_carry_15_, add_1_root_r115_carry_16_,
         add_1_root_r115_carry_17_, add_1_root_r115_carry_18_,
         add_1_root_r115_carry_19_, add_1_root_r115_carry_20_,
         add_1_root_r115_carry_21_, add_1_root_r115_carry_22_,
         add_1_root_r115_carry_7_, add_1_root_r115_carry_8_,
         add_1_root_r115_carry_9_, add_1_root_r115_SUM_6_,
         add_1_root_r115_SUM_7_, add_1_root_r115_SUM_8_,
         add_1_root_r115_SUM_9_, add_1_root_r115_SUM_10_,
         add_1_root_r115_SUM_11_, add_1_root_r115_SUM_12_,
         add_1_root_r115_SUM_13_, add_1_root_r115_SUM_14_,
         add_1_root_r115_SUM_15_, add_1_root_r115_SUM_16_,
         add_1_root_r115_SUM_17_, add_1_root_r115_SUM_18_,
         add_1_root_r115_SUM_19_, add_1_root_r115_SUM_20_,
         add_1_root_r115_SUM_21_, add_1_root_r115_SUM_22_,
         add_1_root_r115_SUM_23_, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n20, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n158, n160, n161, n162, n163, n164, n168, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268;
  wire   [16:0] in_17bit_b;
  wire   [23:8] neg_mul;
  wire   [16:13] sub_add_75_b0_carry;
  wire   [16:2] sub_add_54_b0_carry;
  wire   [22:7] add_1_root_r119_carry;

  multi16_2_DW01_add_0 add_0_root_r119 ( .A_22_(add_2_root_r119_SUM_22_), 
        .A_21_(add_2_root_r119_SUM_21_), .A_20_(add_2_root_r119_SUM_20_), 
        .A_19_(add_2_root_r119_SUM_19_), .A_18_(add_2_root_r119_SUM_18_), 
        .A_17_(add_2_root_r119_SUM_17_), .A_16_(add_2_root_r119_SUM_16_), 
        .A_15_(add_2_root_r119_SUM_15_), .A_14_(add_2_root_r119_SUM_14_), 
        .A_13_(add_2_root_r119_SUM_13_), .A_12_(add_2_root_r119_SUM_12_), 
        .A_11_(add_2_root_r119_SUM_11_), .A_10_(add_2_root_r119_SUM_10_), 
        .A_9_(add_2_root_r119_SUM_9_), .A_8_(add_2_root_r119_SUM_8_), .A_7_(
        add_2_root_r119_SUM_7_), .A_6_(add_2_root_r119_SUM_6_), .A_5_(
        add_1_root_r119_A_2_), .A_4_(in_17bit_b[0]), .B_23_(
        add_1_root_r119_SUM_23_), .B_22_(add_1_root_r119_SUM_22_), .B_21_(
        add_1_root_r119_SUM_21_), .B_20_(add_1_root_r119_SUM_20_), .B_19_(
        add_1_root_r119_SUM_19_), .B_18_(add_1_root_r119_SUM_18_), .B_17_(
        add_1_root_r119_SUM_17_), .B_16_(add_1_root_r119_SUM_16_), .B_15_(
        add_1_root_r119_SUM_15_), .B_14_(add_1_root_r119_SUM_14_), .B_13_(
        add_1_root_r119_SUM_13_), .B_12_(add_1_root_r119_SUM_12_), .B_11_(
        add_1_root_r119_SUM_11_), .B_10_(add_1_root_r119_SUM_10_), .B_9_(
        add_1_root_r119_SUM_9_), .B_8_(add_1_root_r119_SUM_8_), .B_7_(
        add_1_root_r119_SUM_7_), .B_6_(add_1_root_r119_SUM_6_), .B_5_(
        add_1_root_r119_A_5_), .B_4_(add_1_root_r119_A_4_), .SUM_23_(N363), 
        .SUM_22_(N362), .SUM_21_(N361), .SUM_20_(N360), .SUM_19_(N359), 
        .SUM_18_(N358), .SUM_17_(N357), .SUM_16_(N356), .SUM_15_(N355), 
        .SUM_14_(N354), .SUM_13_(N353), .SUM_12_(N352), .SUM_11_(N351), 
        .SUM_10_(N350), .SUM_9_(N349), .SUM_8_(N348), .SUM_7_(N347) );
  multi16_2_DW01_add_4 add_0_root_r112 ( .A_21_(in_17bit_b[16]), .A_20_(
        in_17bit_b[15]), .A_19_(in_17bit_b[14]), .A_18_(in_17bit_b[13]), 
        .A_17_(in_17bit_b[12]), .A_16_(in_17bit_b[11]), .A_15_(in_17bit_b[10]), 
        .A_14_(in_17bit_b[9]), .A_13_(in_17bit_b[8]), .A_12_(in_17bit_b[7]), 
        .A_11_(in_17bit_b[6]), .A_10_(in_17bit_b[5]), .A_9_(in_17bit_b[4]), 
        .A_8_(in_17bit_b[3]), .A_7_(in_17bit_b[2]), .A_6_(n187), .A_5_(
        in_17bit_b[0]), .B_21_(add_1_root_r112_SUM_21_), .B_20_(
        add_1_root_r112_SUM_20_), .B_19_(add_1_root_r112_SUM_19_), .B_18_(
        add_1_root_r112_SUM_18_), .B_17_(add_1_root_r112_SUM_17_), .B_16_(
        add_1_root_r112_SUM_16_), .B_15_(add_1_root_r112_SUM_15_), .B_14_(
        add_1_root_r112_SUM_14_), .B_13_(add_1_root_r112_SUM_13_), .B_12_(
        add_1_root_r112_SUM_12_), .B_11_(add_1_root_r112_SUM_11_), .B_10_(
        add_1_root_r112_SUM_10_), .B_9_(add_1_root_r112_SUM_9_), .B_8_(
        add_1_root_r112_SUM_8_), .B_7_(add_1_root_r112_SUM_7_), .B_6_(
        add_1_root_r112_SUM_6_), .B_5_(add_1_root_r112_SUM_5_), .SUM_22_(N123), 
        .SUM_21_(N122), .SUM_20_(N121), .SUM_19_(N120), .SUM_18_(N119), 
        .SUM_17_(N118), .SUM_16_(N117), .SUM_15_(N116), .SUM_14_(N115), 
        .SUM_13_(N114), .SUM_12_(N113), .SUM_11_(N112), .SUM_10_(N111), 
        .SUM_9_(N110), .SUM_8_(N109), .SUM_7_(N108) );
  multi16_2_DW01_add_6 add_0_root_r115 ( .A_23_(add_1_root_r115_SUM_23_), 
        .A_22_(add_1_root_r115_SUM_22_), .A_21_(add_1_root_r115_SUM_21_), 
        .A_20_(add_1_root_r115_SUM_20_), .A_19_(add_1_root_r115_SUM_19_), 
        .A_18_(add_1_root_r115_SUM_18_), .A_17_(add_1_root_r115_SUM_17_), 
        .A_16_(add_1_root_r115_SUM_16_), .A_15_(add_1_root_r115_SUM_15_), 
        .A_14_(add_1_root_r115_SUM_14_), .A_13_(add_1_root_r115_SUM_13_), 
        .A_12_(add_1_root_r115_SUM_12_), .A_11_(add_1_root_r115_SUM_11_), 
        .A_10_(add_1_root_r115_SUM_10_), .A_9_(add_1_root_r115_SUM_9_), .A_8_(
        add_1_root_r115_SUM_8_), .A_7_(add_1_root_r115_SUM_7_), .A_6_(
        add_1_root_r115_SUM_6_), .A_5_(n187), .A_4_(in_17bit_b[0]), .B_20_(
        add_2_root_r115_SUM_20_), .B_19_(add_2_root_r115_SUM_19_), .B_18_(
        add_2_root_r115_SUM_18_), .B_17_(add_2_root_r115_SUM_17_), .B_16_(
        add_2_root_r115_SUM_16_), .B_15_(add_2_root_r115_SUM_15_), .B_14_(
        add_2_root_r115_SUM_14_), .B_13_(add_2_root_r115_SUM_13_), .B_12_(
        add_2_root_r115_SUM_12_), .B_11_(add_2_root_r115_SUM_11_), .B_10_(
        add_2_root_r115_SUM_10_), .B_9_(add_2_root_r115_SUM_9_), .B_8_(
        add_2_root_r115_SUM_8_), .B_7_(add_2_root_r115_SUM_7_), .B_6_(
        add_2_root_r115_SUM_6_), .B_5_(add_2_root_r115_SUM_5_), .B_4_(
        add_2_root_r115_SUM_4_), .SUM_23_(N221), .SUM_22_(N220), .SUM_21_(N219), .SUM_20_(N218), .SUM_19_(N217), .SUM_18_(N216), .SUM_17_(N215), .SUM_16_(
        N214), .SUM_15_(N213), .SUM_14_(N212), .SUM_13_(N211), .SUM_12_(N210), 
        .SUM_11_(N209), .SUM_10_(N208), .SUM_9_(N207), .SUM_8_(N206), .SUM_7_(
        N205) );
  TLATX1 neg_mul_reg_19_ ( .G(N446), .D(N459), .Q(n1), .QN(n14) );
  TLATX1 neg_mul_reg_18_ ( .G(N446), .D(N458), .QN(n5) );
  TLATX1 neg_mul_reg_17_ ( .G(N446), .D(N457), .QN(n8) );
  TLATX1 neg_mul_reg_16_ ( .G(N446), .D(N456), .QN(n7) );
  TLATX1 neg_mul_reg_15_ ( .G(N446), .D(N455), .QN(n3) );
  TLATX1 neg_mul_reg_13_ ( .G(N446), .D(N453), .Q(neg_mul[13]), .QN(n2) );
  TLATX1 neg_mul_reg_12_ ( .G(N446), .D(N452), .QN(n4) );
  TLATX1 neg_mul_reg_11_ ( .G(N446), .D(N451), .QN(n6) );
  TLATX1 neg_mul_reg_23_ ( .G(N446), .D(N463), .Q(neg_mul[23]), .QN(n16) );
  TLATX1 neg_mul_reg_22_ ( .G(N446), .D(N462), .Q(neg_mul[22]), .QN(n13) );
  TLATX1 neg_mul_reg_21_ ( .G(N446), .D(N461), .QN(n27) );
  TLATX1 neg_mul_reg_20_ ( .G(N446), .D(N460), .QN(n15) );
  TLATX1 neg_mul_reg_14_ ( .G(N446), .D(N454), .Q(neg_mul[14]), .QN(n12) );
  TLATX1 neg_mul_reg_10_ ( .G(N446), .D(N450), .Q(neg_mul[10]), .QN(n9) );
  TLATX1 neg_mul_reg_9_ ( .G(N446), .D(N449), .Q(neg_mul[9]), .QN(n10) );
  TLATX1 neg_mul_reg_8_ ( .G(N446), .D(N448), .Q(neg_mul[8]), .QN(n11) );
  TLATX1 neg_mul_reg_7_ ( .G(N446), .D(N447), .Q(out[0]) );
  NOR2X4 U2 ( .A(n59), .B(n69), .Y(n70) );
  CLKINVX3 U3 ( .A(n61), .Y(n23) );
  CLKINVX1 U4 ( .A(n57), .Y(n61) );
  CLKINVX3 U5 ( .A(n268), .Y(in_17bit_b[16]) );
  MXI2X4 U6 ( .A(n15), .B(n41), .S0(n99), .Y(out[13]) );
  INVX1 U7 ( .A(n88), .Y(n65) );
  MXI2X1 U8 ( .A(n27), .B(n17), .S0(n99), .Y(out[14]) );
  INVX1 U9 ( .A(n168), .Y(n161) );
  XNOR2X1 U10 ( .A(n27), .B(sub_add_75_b0_carry[14]), .Y(n17) );
  BUFX8 U11 ( .A(in_17bit[16]), .Y(n24) );
  AOI2BB2X1 U12 ( .B0(n52), .B1(n12), .A0N(n20), .A1N(n91), .Y(n92) );
  AOI2BB2X1 U13 ( .B0(n89), .B1(n52), .A0N(n20), .A1N(neg_mul[14]), .Y(n90) );
  NAND4BX1 U14 ( .AN(n20), .B(in_8bit[6]), .C(n51), .D(in_8bit[4]), .Y(n168)
         );
  AOI2BB2X4 U15 ( .B0(n66), .B1(n53), .A0N(n53), .A1N(neg_mul[8]), .Y(n67) );
  OAI2BB1X2 U16 ( .A0N(n44), .A1N(n54), .B0(n72), .Y(n75) );
  NOR2BX2 U17 ( .AN(n58), .B(n92), .Y(n93) );
  XNOR2X4 U18 ( .A(n57), .B(n52), .Y(n95) );
  NOR2BX4 U19 ( .AN(n64), .B(n85), .Y(n84) );
  XNOR2X4 U20 ( .A(n18), .B(n5), .Y(out[11]) );
  NOR2X4 U21 ( .A(n98), .B(n38), .Y(n18) );
  CLKINVX8 U22 ( .A(n59), .Y(n60) );
  AOI2BB2X4 U23 ( .B0(n78), .B1(n52), .A0N(n52), .A1N(neg_mul[10]), .Y(n79) );
  XNOR2X2 U24 ( .A(n24), .B(n20), .Y(n86) );
  OAI2BB2X2 U25 ( .B0(neg_mul[9]), .B1(n20), .A0N(n53), .A1N(n44), .Y(n76) );
  BUFX12 U26 ( .A(n269), .Y(out[3]) );
  INVX4 U27 ( .A(n98), .Y(n99) );
  NOR2X4 U28 ( .A(n24), .B(n67), .Y(n71) );
  BUFX8 U29 ( .A(n270), .Y(out[2]) );
  AOI221X2 U30 ( .A0(n63), .A1(n76), .B0(n58), .B1(n75), .C0(n74), .Y(n270) );
  INVX8 U31 ( .A(n54), .Y(n20) );
  NOR2X4 U32 ( .A(n79), .B(n58), .Y(n22) );
  NOR3X4 U33 ( .A(n82), .B(n22), .C(n83), .Y(n269) );
  NOR2BX4 U34 ( .AN(n24), .B(n81), .Y(n82) );
  XOR2X4 U35 ( .A(n87), .B(neg_mul[13]), .Y(out[6]) );
  AOI2BB2X2 U36 ( .B0(n52), .B1(n9), .A0N(n53), .A1N(n80), .Y(n81) );
  NOR2X2 U37 ( .A(n57), .B(n90), .Y(n94) );
  INVX8 U38 ( .A(n54), .Y(n52) );
  NAND2X2 U39 ( .A(n53), .B(n10), .Y(n72) );
  INVX8 U40 ( .A(in_8bit[7]), .Y(n54) );
  INVXL U41 ( .A(in_8bit[0]), .Y(n50) );
  INVXL U42 ( .A(in_8bit[4]), .Y(n49) );
  INVX8 U43 ( .A(n59), .Y(n58) );
  INVX8 U44 ( .A(n54), .Y(n53) );
  INVXL U45 ( .A(n23), .Y(n62) );
  INVX8 U46 ( .A(in_17bit[16]), .Y(n59) );
  INVX8 U47 ( .A(n60), .Y(n63) );
  INVX8 U48 ( .A(n63), .Y(n57) );
  OR2X4 U49 ( .A(n98), .B(n40), .Y(n32) );
  XNOR2X4 U50 ( .A(n57), .B(n52), .Y(n98) );
  CLKBUFXL U51 ( .A(in_8bit[1]), .Y(n51) );
  INVX1 U52 ( .A(n257), .Y(in_17bit_b[14]) );
  INVX1 U53 ( .A(n254), .Y(in_17bit_b[13]) );
  INVX1 U54 ( .A(n221), .Y(in_17bit_b[2]) );
  INVX1 U55 ( .A(n230), .Y(in_17bit_b[5]) );
  INVX1 U56 ( .A(n233), .Y(in_17bit_b[6]) );
  INVX1 U57 ( .A(n236), .Y(in_17bit_b[7]) );
  INVX1 U58 ( .A(n239), .Y(in_17bit_b[8]) );
  INVX1 U59 ( .A(n242), .Y(in_17bit_b[9]) );
  INVX1 U60 ( .A(n245), .Y(in_17bit_b[10]) );
  INVX1 U61 ( .A(n248), .Y(in_17bit_b[11]) );
  INVX1 U62 ( .A(n251), .Y(in_17bit_b[12]) );
  INVX1 U63 ( .A(n227), .Y(in_17bit_b[4]) );
  INVX1 U64 ( .A(n224), .Y(in_17bit_b[3]) );
  XNOR2X4 U65 ( .A(n25), .B(n4), .Y(out[5]) );
  NOR2X4 U66 ( .A(n34), .B(n85), .Y(n25) );
  XNOR2X4 U67 ( .A(n26), .B(n3), .Y(out[8]) );
  NOR2X4 U68 ( .A(n33), .B(n95), .Y(n26) );
  AOI21X1 U69 ( .A0(n28), .A1(n29), .B0(n261), .Y(n214) );
  NOR4XL U70 ( .A(in_8bit[4]), .B(n55), .C(in_8bit[6]), .D(n20), .Y(n28) );
  NOR4XL U71 ( .A(n51), .B(in_8bit[0]), .C(in_8bit[2]), .D(in_8bit[3]), .Y(n29) );
  AND4X1 U72 ( .A(n51), .B(n20), .C(n208), .D(n50), .Y(n30) );
  NAND2X1 U73 ( .A(n31), .B(n51), .Y(n100) );
  NOR3X1 U74 ( .A(n47), .B(n48), .C(n50), .Y(n213) );
  NAND3X1 U75 ( .A(in_8bit[2]), .B(n48), .C(n55), .Y(n209) );
  ADDFX2 U76 ( .A(in_17bit_b[16]), .B(in_17bit_b[12]), .CI(
        add_1_root_r112_carry_16_), .CO(add_1_root_r112_carry_17_), .S(
        add_1_root_r112_SUM_16_) );
  ADDFX2 U77 ( .A(add_1_root_r119_A_19_), .B(in_17bit_b[13]), .CI(
        add_1_root_r119_carry[19]), .CO(add_1_root_r119_carry[20]), .S(
        add_1_root_r119_SUM_19_) );
  ADDFX2 U78 ( .A(in_17bit_b[16]), .B(in_17bit_b[15]), .CI(
        add_3_root_r119_carry_17_), .CO(add_3_root_r119_carry_18_), .S(
        add_1_root_r119_A_17_) );
  ADDFX2 U79 ( .A(in_17bit_b[16]), .B(in_17bit_b[14]), .CI(
        add_2_root_r115_carry_17_), .CO(add_2_root_r115_carry_18_), .S(
        add_2_root_r115_SUM_17_) );
  ADDFX2 U80 ( .A(in_17bit_b[16]), .B(in_17bit_b[14]), .CI(
        add_1_root_r115_carry_20_), .CO(add_1_root_r115_carry_21_), .S(
        add_1_root_r115_SUM_20_) );
  ADDFX2 U81 ( .A(in_17bit_b[16]), .B(in_17bit_b[15]), .CI(
        add_2_root_r119_carry_20_), .CO(add_2_root_r119_carry_21_), .S(
        add_2_root_r119_SUM_20_) );
  AND3X1 U82 ( .A(n20), .B(n49), .C(n56), .Y(n31) );
  NOR2XL U83 ( .A(n20), .B(n49), .Y(n101) );
  ADDFX2 U84 ( .A(in_17bit_b[3]), .B(n187), .CI(add_1_root_r115_carry_7_), 
        .CO(add_2_root_r115_carry_5_), .S(add_2_root_r115_SUM_4_) );
  ADDFX2 U85 ( .A(in_17bit_b[4]), .B(in_17bit_b[2]), .CI(
        add_2_root_r115_carry_5_), .CO(add_2_root_r115_carry_6_), .S(
        add_2_root_r115_SUM_5_) );
  ADDFX2 U86 ( .A(in_17bit_b[5]), .B(n187), .CI(add_1_root_r112_carry_5_), 
        .CO(add_1_root_r112_carry_6_), .S(add_1_root_r112_SUM_5_) );
  ADDFX2 U87 ( .A(in_17bit_b[6]), .B(in_17bit_b[5]), .CI(
        add_3_root_r119_carry_7_), .CO(add_3_root_r119_carry_8_), .S(
        add_1_root_r119_A_7_) );
  ADDFX2 U88 ( .A(in_17bit_b[6]), .B(in_17bit_b[2]), .CI(
        add_1_root_r112_carry_6_), .CO(add_1_root_r112_carry_7_), .S(
        add_1_root_r112_SUM_6_) );
  ADDFX2 U89 ( .A(in_17bit_b[3]), .B(n187), .CI(add_1_root_r115_carry_7_), 
        .CO(add_1_root_r115_carry_8_), .S(add_1_root_r115_SUM_7_) );
  ADDFX2 U90 ( .A(in_17bit_b[7]), .B(in_17bit_b[6]), .CI(
        add_3_root_r119_carry_8_), .CO(add_3_root_r119_carry_9_), .S(
        add_1_root_r119_A_8_) );
  ADDFX2 U91 ( .A(add_1_root_r119_A_7_), .B(n187), .CI(
        add_1_root_r119_carry[7]), .CO(add_1_root_r119_carry[8]), .S(
        add_1_root_r119_SUM_7_) );
  ADDFX2 U92 ( .A(in_17bit_b[2]), .B(n187), .CI(add_3_root_r119_carry_3_), 
        .CO(add_2_root_r119_carry_7_), .S(add_2_root_r119_SUM_6_) );
  ADDFX2 U93 ( .A(in_17bit_b[4]), .B(in_17bit_b[2]), .CI(
        add_1_root_r115_carry_8_), .CO(add_1_root_r115_carry_9_), .S(
        add_1_root_r115_SUM_8_) );
  ADDFX2 U94 ( .A(in_17bit_b[8]), .B(in_17bit_b[7]), .CI(
        add_3_root_r119_carry_9_), .CO(add_3_root_r119_carry_10_), .S(
        add_1_root_r119_A_9_) );
  ADDFX2 U95 ( .A(add_1_root_r119_A_8_), .B(in_17bit_b[2]), .CI(
        add_1_root_r119_carry[8]), .CO(add_1_root_r119_carry[9]), .S(
        add_1_root_r119_SUM_8_) );
  ADDFX2 U96 ( .A(in_17bit_b[3]), .B(in_17bit_b[2]), .CI(
        add_2_root_r119_carry_7_), .CO(add_2_root_r119_carry_8_), .S(
        add_2_root_r119_SUM_7_) );
  ADDFX2 U97 ( .A(in_17bit_b[6]), .B(in_17bit_b[4]), .CI(
        add_2_root_r115_carry_7_), .CO(add_2_root_r115_carry_8_), .S(
        add_2_root_r115_SUM_7_) );
  ADDFX2 U98 ( .A(in_17bit_b[8]), .B(in_17bit_b[4]), .CI(
        add_1_root_r112_carry_8_), .CO(add_1_root_r112_carry_9_), .S(
        add_1_root_r112_SUM_8_) );
  ADDFX2 U99 ( .A(in_17bit_b[9]), .B(in_17bit_b[8]), .CI(
        add_3_root_r119_carry_10_), .CO(add_3_root_r119_carry_11_), .S(
        add_1_root_r119_A_10_) );
  ADDFX2 U100 ( .A(in_17bit_b[7]), .B(in_17bit_b[5]), .CI(
        add_2_root_r115_carry_8_), .CO(add_2_root_r115_carry_9_), .S(
        add_2_root_r115_SUM_8_) );
  ADDFX2 U101 ( .A(in_17bit_b[9]), .B(in_17bit_b[5]), .CI(
        add_1_root_r112_carry_9_), .CO(add_1_root_r112_carry_10_), .S(
        add_1_root_r112_SUM_9_) );
  ADDFX2 U102 ( .A(in_17bit_b[10]), .B(in_17bit_b[9]), .CI(
        add_3_root_r119_carry_11_), .CO(add_3_root_r119_carry_12_), .S(
        add_1_root_r119_A_11_) );
  ADDFX2 U103 ( .A(add_1_root_r119_A_10_), .B(in_17bit_b[4]), .CI(
        add_1_root_r119_carry[10]), .CO(add_1_root_r119_carry[11]), .S(
        add_1_root_r119_SUM_10_) );
  ADDFX2 U104 ( .A(in_17bit_b[8]), .B(in_17bit_b[6]), .CI(
        add_2_root_r115_carry_9_), .CO(add_2_root_r115_carry_10_), .S(
        add_2_root_r115_SUM_9_) );
  ADDFX2 U105 ( .A(in_17bit_b[10]), .B(in_17bit_b[6]), .CI(
        add_1_root_r112_carry_10_), .CO(add_1_root_r112_carry_11_), .S(
        add_1_root_r112_SUM_10_) );
  ADDFX2 U106 ( .A(in_17bit_b[7]), .B(in_17bit_b[5]), .CI(
        add_1_root_r115_carry_11_), .CO(add_1_root_r115_carry_12_), .S(
        add_1_root_r115_SUM_11_) );
  ADDFX2 U107 ( .A(in_17bit_b[11]), .B(in_17bit_b[10]), .CI(
        add_3_root_r119_carry_12_), .CO(add_3_root_r119_carry_13_), .S(
        add_1_root_r119_A_12_) );
  ADDFX2 U108 ( .A(add_1_root_r119_A_11_), .B(in_17bit_b[5]), .CI(
        add_1_root_r119_carry[11]), .CO(add_1_root_r119_carry[12]), .S(
        add_1_root_r119_SUM_11_) );
  ADDFX2 U109 ( .A(in_17bit_b[6]), .B(in_17bit_b[5]), .CI(
        add_2_root_r119_carry_10_), .CO(add_2_root_r119_carry_11_), .S(
        add_2_root_r119_SUM_10_) );
  ADDFX2 U110 ( .A(in_17bit_b[9]), .B(in_17bit_b[7]), .CI(
        add_2_root_r115_carry_10_), .CO(add_2_root_r115_carry_11_), .S(
        add_2_root_r115_SUM_10_) );
  ADDFX2 U111 ( .A(in_17bit_b[8]), .B(in_17bit_b[6]), .CI(
        add_1_root_r115_carry_12_), .CO(add_1_root_r115_carry_13_), .S(
        add_1_root_r115_SUM_12_) );
  ADDFX2 U112 ( .A(in_17bit_b[12]), .B(in_17bit_b[11]), .CI(
        add_3_root_r119_carry_13_), .CO(add_3_root_r119_carry_14_), .S(
        add_1_root_r119_A_13_) );
  ADDFX2 U113 ( .A(in_17bit_b[7]), .B(in_17bit_b[6]), .CI(
        add_2_root_r119_carry_11_), .CO(add_2_root_r119_carry_12_), .S(
        add_2_root_r119_SUM_11_) );
  ADDFX2 U114 ( .A(in_17bit_b[10]), .B(in_17bit_b[8]), .CI(
        add_2_root_r115_carry_11_), .CO(add_2_root_r115_carry_12_), .S(
        add_2_root_r115_SUM_11_) );
  ADDFX2 U115 ( .A(in_17bit_b[12]), .B(in_17bit_b[8]), .CI(
        add_1_root_r112_carry_12_), .CO(add_1_root_r112_carry_13_), .S(
        add_1_root_r112_SUM_12_) );
  ADDFX2 U116 ( .A(in_17bit_b[9]), .B(in_17bit_b[7]), .CI(
        add_1_root_r115_carry_13_), .CO(add_1_root_r115_carry_14_), .S(
        add_1_root_r115_SUM_13_) );
  ADDFX2 U117 ( .A(in_17bit_b[13]), .B(in_17bit_b[12]), .CI(
        add_3_root_r119_carry_14_), .CO(add_3_root_r119_carry_15_), .S(
        add_1_root_r119_A_14_) );
  ADDFX2 U118 ( .A(add_1_root_r119_A_13_), .B(in_17bit_b[7]), .CI(
        add_1_root_r119_carry[13]), .CO(add_1_root_r119_carry[14]), .S(
        add_1_root_r119_SUM_13_) );
  ADDFX2 U119 ( .A(in_17bit_b[8]), .B(in_17bit_b[7]), .CI(
        add_2_root_r119_carry_12_), .CO(add_2_root_r119_carry_13_), .S(
        add_2_root_r119_SUM_12_) );
  ADDFX2 U120 ( .A(in_17bit_b[11]), .B(in_17bit_b[9]), .CI(
        add_2_root_r115_carry_12_), .CO(add_2_root_r115_carry_13_), .S(
        add_2_root_r115_SUM_12_) );
  ADDFX2 U121 ( .A(in_17bit_b[13]), .B(in_17bit_b[9]), .CI(
        add_1_root_r112_carry_13_), .CO(add_1_root_r112_carry_14_), .S(
        add_1_root_r112_SUM_13_) );
  ADDFX2 U122 ( .A(in_17bit_b[10]), .B(in_17bit_b[8]), .CI(
        add_1_root_r115_carry_14_), .CO(add_1_root_r115_carry_15_), .S(
        add_1_root_r115_SUM_14_) );
  ADDFX2 U123 ( .A(in_17bit_b[14]), .B(in_17bit_b[13]), .CI(
        add_3_root_r119_carry_15_), .CO(add_3_root_r119_carry_16_), .S(
        add_1_root_r119_A_15_) );
  ADDFX2 U124 ( .A(add_1_root_r119_A_14_), .B(in_17bit_b[8]), .CI(
        add_1_root_r119_carry[14]), .CO(add_1_root_r119_carry[15]), .S(
        add_1_root_r119_SUM_14_) );
  ADDFX2 U125 ( .A(in_17bit_b[9]), .B(in_17bit_b[8]), .CI(
        add_2_root_r119_carry_13_), .CO(add_2_root_r119_carry_14_), .S(
        add_2_root_r119_SUM_13_) );
  ADDFX2 U126 ( .A(in_17bit_b[12]), .B(in_17bit_b[10]), .CI(
        add_2_root_r115_carry_13_), .CO(add_2_root_r115_carry_14_), .S(
        add_2_root_r115_SUM_13_) );
  ADDFX2 U127 ( .A(in_17bit_b[14]), .B(in_17bit_b[10]), .CI(
        add_1_root_r112_carry_14_), .CO(add_1_root_r112_carry_15_), .S(
        add_1_root_r112_SUM_14_) );
  ADDFX2 U128 ( .A(in_17bit_b[11]), .B(in_17bit_b[9]), .CI(
        add_1_root_r115_carry_15_), .CO(add_1_root_r115_carry_16_), .S(
        add_1_root_r115_SUM_15_) );
  ADDFX2 U129 ( .A(add_1_root_r119_A_15_), .B(in_17bit_b[9]), .CI(
        add_1_root_r119_carry[15]), .CO(add_1_root_r119_carry[16]), .S(
        add_1_root_r119_SUM_15_) );
  ADDFX2 U130 ( .A(in_17bit_b[3]), .B(in_17bit_b[2]), .CI(
        add_3_root_r119_carry_4_), .CO(add_3_root_r119_carry_5_), .S(
        add_1_root_r119_A_4_) );
  ADDFX2 U131 ( .A(in_17bit_b[2]), .B(n187), .CI(add_3_root_r119_carry_3_), 
        .CO(add_3_root_r119_carry_4_), .S(add_1_root_r119_A_3_) );
  ADDFX2 U132 ( .A(in_17bit_b[10]), .B(in_17bit_b[9]), .CI(
        add_2_root_r119_carry_14_), .CO(add_2_root_r119_carry_15_), .S(
        add_2_root_r119_SUM_14_) );
  ADDFX2 U133 ( .A(in_17bit_b[15]), .B(in_17bit_b[11]), .CI(
        add_1_root_r112_carry_15_), .CO(add_1_root_r112_carry_16_), .S(
        add_1_root_r112_SUM_15_) );
  ADDFX2 U134 ( .A(add_1_root_r119_A_16_), .B(in_17bit_b[10]), .CI(
        add_1_root_r119_carry[16]), .CO(add_1_root_r119_carry[17]), .S(
        add_1_root_r119_SUM_16_) );
  ADDFX2 U135 ( .A(in_17bit_b[11]), .B(in_17bit_b[10]), .CI(
        add_2_root_r119_carry_15_), .CO(add_2_root_r119_carry_16_), .S(
        add_2_root_r119_SUM_15_) );
  ADDFX2 U136 ( .A(in_17bit_b[14]), .B(in_17bit_b[12]), .CI(
        add_2_root_r115_carry_15_), .CO(add_2_root_r115_carry_16_), .S(
        add_2_root_r115_SUM_15_) );
  ADDFX2 U137 ( .A(in_17bit_b[13]), .B(in_17bit_b[11]), .CI(
        add_1_root_r115_carry_17_), .CO(add_1_root_r115_carry_18_), .S(
        add_1_root_r115_SUM_17_) );
  ADDFX2 U138 ( .A(add_1_root_r119_A_17_), .B(in_17bit_b[11]), .CI(
        add_1_root_r119_carry[17]), .CO(add_1_root_r119_carry[18]), .S(
        add_1_root_r119_SUM_17_) );
  ADDFX2 U139 ( .A(in_17bit_b[12]), .B(in_17bit_b[11]), .CI(
        add_2_root_r119_carry_16_), .CO(add_2_root_r119_carry_17_), .S(
        add_2_root_r119_SUM_16_) );
  ADDFX2 U140 ( .A(in_17bit_b[15]), .B(in_17bit_b[13]), .CI(
        add_2_root_r115_carry_16_), .CO(add_2_root_r115_carry_17_), .S(
        add_2_root_r115_SUM_16_) );
  ADDFX2 U141 ( .A(in_17bit_b[14]), .B(in_17bit_b[12]), .CI(
        add_1_root_r115_carry_18_), .CO(add_1_root_r115_carry_19_), .S(
        add_1_root_r115_SUM_18_) );
  ADDFX2 U142 ( .A(add_1_root_r119_A_18_), .B(in_17bit_b[12]), .CI(
        add_1_root_r119_carry[18]), .CO(add_1_root_r119_carry[19]), .S(
        add_1_root_r119_SUM_18_) );
  ADDFX2 U143 ( .A(in_17bit_b[5]), .B(in_17bit_b[4]), .CI(
        add_3_root_r119_carry_6_), .CO(add_3_root_r119_carry_7_), .S(
        add_1_root_r119_A_6_) );
  ADDFX2 U144 ( .A(in_17bit_b[15]), .B(in_17bit_b[13]), .CI(
        add_1_root_r115_carry_19_), .CO(add_1_root_r115_carry_20_), .S(
        add_1_root_r115_SUM_19_) );
  ADDFX2 U145 ( .A(in_17bit_b[14]), .B(in_17bit_b[13]), .CI(
        add_2_root_r119_carry_18_), .CO(add_2_root_r119_carry_19_), .S(
        add_2_root_r119_SUM_18_) );
  ADDFX2 U146 ( .A(in_17bit_b[5]), .B(in_17bit_b[3]), .CI(
        add_2_root_r115_carry_6_), .CO(add_2_root_r115_carry_7_), .S(
        add_2_root_r115_SUM_6_) );
  ADDFX2 U147 ( .A(in_17bit_b[7]), .B(in_17bit_b[3]), .CI(
        add_1_root_r112_carry_7_), .CO(add_1_root_r112_carry_8_), .S(
        add_1_root_r112_SUM_7_) );
  ADDFX2 U148 ( .A(in_17bit_b[5]), .B(in_17bit_b[3]), .CI(
        add_1_root_r115_carry_9_), .CO(add_1_root_r115_carry_10_), .S(
        add_1_root_r115_SUM_9_) );
  ADDFX2 U149 ( .A(add_1_root_r119_A_9_), .B(in_17bit_b[3]), .CI(
        add_1_root_r119_carry[9]), .CO(add_1_root_r119_carry[10]), .S(
        add_1_root_r119_SUM_9_) );
  ADDFX2 U150 ( .A(in_17bit_b[4]), .B(in_17bit_b[3]), .CI(
        add_2_root_r119_carry_8_), .CO(add_2_root_r119_carry_9_), .S(
        add_2_root_r119_SUM_8_) );
  ADDFX2 U151 ( .A(in_17bit_b[6]), .B(in_17bit_b[4]), .CI(
        add_1_root_r115_carry_10_), .CO(add_1_root_r115_carry_11_), .S(
        add_1_root_r115_SUM_10_) );
  ADDFX2 U152 ( .A(in_17bit_b[5]), .B(in_17bit_b[4]), .CI(
        add_2_root_r119_carry_9_), .CO(add_2_root_r119_carry_10_), .S(
        add_2_root_r119_SUM_9_) );
  ADDFX2 U153 ( .A(in_17bit_b[11]), .B(in_17bit_b[7]), .CI(
        add_1_root_r112_carry_11_), .CO(add_1_root_r112_carry_12_), .S(
        add_1_root_r112_SUM_11_) );
  ADDFX2 U154 ( .A(add_1_root_r119_A_12_), .B(in_17bit_b[6]), .CI(
        add_1_root_r119_carry[12]), .CO(add_1_root_r119_carry[13]), .S(
        add_1_root_r119_SUM_12_) );
  ADDFX2 U155 ( .A(in_17bit_b[13]), .B(in_17bit_b[11]), .CI(
        add_2_root_r115_carry_14_), .CO(add_2_root_r115_carry_15_), .S(
        add_2_root_r115_SUM_14_) );
  ADDFX2 U156 ( .A(in_17bit_b[12]), .B(in_17bit_b[10]), .CI(
        add_1_root_r115_carry_16_), .CO(add_1_root_r115_carry_17_), .S(
        add_1_root_r115_SUM_16_) );
  ADDFX2 U157 ( .A(in_17bit_b[15]), .B(in_17bit_b[14]), .CI(
        add_3_root_r119_carry_16_), .CO(add_3_root_r119_carry_17_), .S(
        add_1_root_r119_A_16_) );
  ADDFX2 U158 ( .A(in_17bit_b[4]), .B(in_17bit_b[3]), .CI(
        add_3_root_r119_carry_5_), .CO(add_3_root_r119_carry_6_), .S(
        add_1_root_r119_A_5_) );
  ADDFX2 U159 ( .A(in_17bit_b[13]), .B(in_17bit_b[12]), .CI(
        add_2_root_r119_carry_17_), .CO(add_2_root_r119_carry_18_), .S(
        add_2_root_r119_SUM_17_) );
  ADDFX2 U160 ( .A(in_17bit_b[15]), .B(in_17bit_b[14]), .CI(
        add_2_root_r119_carry_19_), .CO(add_2_root_r119_carry_20_), .S(
        add_2_root_r119_SUM_19_) );
  INVX1 U161 ( .A(n210), .Y(n164) );
  NAND3BX1 U162 ( .AN(n55), .B(n47), .C(in_8bit[3]), .Y(n210) );
  INVX1 U163 ( .A(n56), .Y(n55) );
  INVX1 U164 ( .A(in_8bit[3]), .Y(n48) );
  CLKINVX3 U165 ( .A(n215), .Y(in_17bit_b[0]) );
  INVX1 U166 ( .A(n188), .Y(n267) );
  NAND2XL U167 ( .A(N29), .B(n23), .Y(n268) );
  OAI21XL U168 ( .A0(n267), .A1(n268), .B0(n266), .Y(N463) );
  AOI22X1 U169 ( .A0(N221), .A1(n46), .B0(N363), .B1(n45), .Y(n266) );
  CLKINVX3 U170 ( .A(n260), .Y(in_17bit_b[15]) );
  INVX1 U171 ( .A(in_8bit[2]), .Y(n47) );
  INVX1 U172 ( .A(in_8bit[5]), .Y(n56) );
  XNOR2X4 U173 ( .A(n32), .B(n1), .Y(out[12]) );
  AOI22X1 U174 ( .A0(in_17bit[0]), .A1(n23), .B0(in_17bit[0]), .B1(n62), .Y(
        n215) );
  AOI22X1 U175 ( .A0(N27), .A1(n23), .B0(in_17bit[14]), .B1(n61), .Y(n257) );
  AOI22X1 U176 ( .A0(N28), .A1(n23), .B0(in_17bit[15]), .B1(n61), .Y(n260) );
  AOI22X1 U177 ( .A0(N14), .A1(n23), .B0(in_17bit[1]), .B1(n62), .Y(n218) );
  AOI22X1 U178 ( .A0(N15), .A1(n23), .B0(in_17bit[2]), .B1(n61), .Y(n221) );
  AOI22X1 U179 ( .A0(N16), .A1(n23), .B0(in_17bit[3]), .B1(n61), .Y(n224) );
  AOI22X1 U180 ( .A0(N17), .A1(n23), .B0(in_17bit[4]), .B1(n61), .Y(n227) );
  AOI22X1 U181 ( .A0(N18), .A1(n23), .B0(in_17bit[5]), .B1(n61), .Y(n230) );
  AOI22X1 U182 ( .A0(N19), .A1(n23), .B0(in_17bit[6]), .B1(n61), .Y(n233) );
  AOI22X1 U183 ( .A0(N20), .A1(n23), .B0(in_17bit[7]), .B1(n61), .Y(n236) );
  AOI22X1 U184 ( .A0(N21), .A1(n23), .B0(in_17bit[8]), .B1(n61), .Y(n239) );
  AOI22X1 U185 ( .A0(N22), .A1(n23), .B0(in_17bit[9]), .B1(n61), .Y(n242) );
  AOI22X1 U186 ( .A0(N23), .A1(n23), .B0(in_17bit[10]), .B1(n61), .Y(n245) );
  AOI22X1 U187 ( .A0(N24), .A1(n23), .B0(in_17bit[11]), .B1(n61), .Y(n248) );
  AOI22X1 U188 ( .A0(N25), .A1(n23), .B0(in_17bit[12]), .B1(n61), .Y(n251) );
  AOI22X1 U189 ( .A0(N26), .A1(n23), .B0(in_17bit[13]), .B1(n61), .Y(n254) );
  INVX1 U190 ( .A(n64), .Y(n83) );
  NAND2BX1 U191 ( .AN(n77), .B(n9), .Y(n64) );
  AND2X2 U192 ( .A(n65), .B(n12), .Y(n33) );
  NAND2X1 U193 ( .A(n42), .B(n10), .Y(n77) );
  AND2X2 U194 ( .A(n83), .B(n6), .Y(n34) );
  AND2X2 U195 ( .A(n33), .B(n3), .Y(n35) );
  AND2X2 U196 ( .A(n34), .B(n4), .Y(n36) );
  AND2X2 U197 ( .A(n35), .B(n7), .Y(n37) );
  AND2X2 U198 ( .A(n37), .B(n8), .Y(n38) );
  BUFX3 U199 ( .A(n264), .Y(n45) );
  OAI2BB1X1 U200 ( .A0N(n164), .A1N(n30), .B0(n162), .Y(n264) );
  NAND2BX1 U201 ( .AN(n209), .B(n39), .Y(n162) );
  BUFX3 U202 ( .A(n265), .Y(n46) );
  OAI2BB1X1 U203 ( .A0N(n39), .A1N(n164), .B0(n163), .Y(n265) );
  NAND2BX1 U204 ( .AN(n209), .B(n30), .Y(n163) );
  NAND2X1 U205 ( .A(n36), .B(n2), .Y(n88) );
  OAI2BB1X1 U206 ( .A0N(n212), .A1N(n31), .B0(n170), .Y(n188) );
  NAND3BX1 U207 ( .AN(n168), .B(n213), .C(n55), .Y(n170) );
  AND2X2 U208 ( .A(n161), .B(n50), .Y(n39) );
  AND2X2 U209 ( .A(n38), .B(n5), .Y(n40) );
  INVX1 U210 ( .A(in_17bit[0]), .Y(n171) );
  INVX1 U211 ( .A(in_17bit[1]), .Y(n172) );
  INVX1 U212 ( .A(in_17bit[2]), .Y(n173) );
  INVX1 U213 ( .A(in_17bit[3]), .Y(n174) );
  INVX1 U214 ( .A(in_17bit[4]), .Y(n175) );
  INVX1 U215 ( .A(in_17bit[5]), .Y(n176) );
  INVX1 U216 ( .A(in_17bit[6]), .Y(n177) );
  INVX1 U217 ( .A(in_17bit[7]), .Y(n178) );
  INVX1 U218 ( .A(in_17bit[8]), .Y(n179) );
  INVX1 U219 ( .A(in_17bit[9]), .Y(n180) );
  INVX1 U220 ( .A(in_17bit[10]), .Y(n181) );
  INVX1 U221 ( .A(in_17bit[11]), .Y(n182) );
  INVX1 U222 ( .A(in_17bit[12]), .Y(n183) );
  INVX1 U223 ( .A(in_17bit[13]), .Y(n184) );
  INVX1 U224 ( .A(in_17bit[14]), .Y(n185) );
  INVX1 U225 ( .A(in_17bit[15]), .Y(n186) );
  INVX1 U226 ( .A(n80), .Y(n78) );
  INVX1 U227 ( .A(n68), .Y(n66) );
  NAND2X1 U228 ( .A(n217), .B(n216), .Y(N447) );
  AOI22X1 U229 ( .A0(N108), .A1(n261), .B0(N205), .B1(n46), .Y(n216) );
  AOI22X1 U230 ( .A0(N347), .A1(n45), .B0(n188), .B1(in_17bit_b[0]), .Y(n217)
         );
  NAND2X1 U231 ( .A(n220), .B(n219), .Y(N448) );
  AOI22X1 U232 ( .A0(N109), .A1(n261), .B0(N206), .B1(n46), .Y(n219) );
  AOI22X1 U233 ( .A0(N348), .A1(n45), .B0(n188), .B1(n187), .Y(n220) );
  INVX1 U234 ( .A(n218), .Y(n187) );
  NAND2X1 U235 ( .A(n223), .B(n222), .Y(N449) );
  AOI22X1 U236 ( .A0(N110), .A1(n261), .B0(N207), .B1(n46), .Y(n222) );
  AOI22X1 U237 ( .A0(N349), .A1(n45), .B0(n188), .B1(in_17bit_b[2]), .Y(n223)
         );
  NAND2X1 U238 ( .A(n226), .B(n225), .Y(N450) );
  AOI22X1 U239 ( .A0(N111), .A1(n261), .B0(N208), .B1(n46), .Y(n225) );
  AOI22X1 U240 ( .A0(N350), .A1(n45), .B0(n188), .B1(in_17bit_b[3]), .Y(n226)
         );
  NAND2X1 U241 ( .A(n229), .B(n228), .Y(N451) );
  AOI22X1 U242 ( .A0(N112), .A1(n261), .B0(N209), .B1(n46), .Y(n228) );
  AOI22X1 U243 ( .A0(N351), .A1(n45), .B0(n188), .B1(in_17bit_b[4]), .Y(n229)
         );
  NAND2X1 U244 ( .A(n232), .B(n231), .Y(N452) );
  AOI22X1 U245 ( .A0(N113), .A1(n261), .B0(N210), .B1(n46), .Y(n231) );
  AOI22X1 U246 ( .A0(N352), .A1(n45), .B0(n188), .B1(in_17bit_b[5]), .Y(n232)
         );
  NAND2X1 U247 ( .A(n235), .B(n234), .Y(N453) );
  AOI22X1 U248 ( .A0(N114), .A1(n261), .B0(N211), .B1(n46), .Y(n234) );
  AOI22X1 U249 ( .A0(N353), .A1(n45), .B0(n188), .B1(in_17bit_b[6]), .Y(n235)
         );
  NAND2X1 U250 ( .A(n238), .B(n237), .Y(N454) );
  AOI22X1 U251 ( .A0(N115), .A1(n261), .B0(N212), .B1(n46), .Y(n237) );
  AOI22X1 U252 ( .A0(N354), .A1(n45), .B0(n188), .B1(in_17bit_b[7]), .Y(n238)
         );
  NAND2X1 U253 ( .A(n241), .B(n240), .Y(N455) );
  AOI22X1 U254 ( .A0(N116), .A1(n261), .B0(N213), .B1(n46), .Y(n240) );
  AOI22X1 U255 ( .A0(N355), .A1(n45), .B0(n188), .B1(in_17bit_b[8]), .Y(n241)
         );
  NAND2X1 U256 ( .A(n244), .B(n243), .Y(N456) );
  AOI22X1 U257 ( .A0(N117), .A1(n261), .B0(N214), .B1(n46), .Y(n243) );
  AOI22X1 U258 ( .A0(N356), .A1(n45), .B0(n188), .B1(in_17bit_b[9]), .Y(n244)
         );
  NAND2X1 U259 ( .A(n247), .B(n246), .Y(N457) );
  AOI22X1 U260 ( .A0(N118), .A1(n261), .B0(N215), .B1(n46), .Y(n246) );
  AOI22X1 U261 ( .A0(N357), .A1(n45), .B0(n188), .B1(in_17bit_b[10]), .Y(n247)
         );
  NAND2X1 U262 ( .A(n250), .B(n249), .Y(N458) );
  AOI22X1 U263 ( .A0(N119), .A1(n261), .B0(N216), .B1(n46), .Y(n249) );
  AOI22X1 U264 ( .A0(N358), .A1(n45), .B0(n188), .B1(in_17bit_b[11]), .Y(n250)
         );
  NAND2X1 U265 ( .A(n253), .B(n252), .Y(N459) );
  AOI22X1 U266 ( .A0(N120), .A1(n261), .B0(N217), .B1(n46), .Y(n252) );
  AOI22X1 U267 ( .A0(N359), .A1(n45), .B0(n188), .B1(in_17bit_b[12]), .Y(n253)
         );
  NAND2X1 U268 ( .A(n256), .B(n255), .Y(N460) );
  AOI22X1 U269 ( .A0(N121), .A1(n261), .B0(N218), .B1(n46), .Y(n255) );
  AOI22X1 U270 ( .A0(N360), .A1(n45), .B0(n188), .B1(in_17bit_b[13]), .Y(n256)
         );
  NAND2X1 U271 ( .A(n259), .B(n258), .Y(N461) );
  AOI22X1 U272 ( .A0(N122), .A1(n261), .B0(N219), .B1(n46), .Y(n258) );
  AOI22X1 U273 ( .A0(N361), .A1(n45), .B0(n188), .B1(in_17bit_b[14]), .Y(n259)
         );
  NAND2X1 U274 ( .A(n263), .B(n262), .Y(N462) );
  AOI22X1 U275 ( .A0(N123), .A1(n261), .B0(N220), .B1(n46), .Y(n262) );
  AOI22X1 U276 ( .A0(N362), .A1(n45), .B0(n188), .B1(in_17bit_b[15]), .Y(n263)
         );
  INVX1 U277 ( .A(n73), .Y(n44) );
  XNOR2X1 U278 ( .A(n15), .B(sub_add_75_b0_carry[13]), .Y(n41) );
  INVX1 U279 ( .A(n77), .Y(n74) );
  INVX1 U280 ( .A(n91), .Y(n89) );
  MX2X1 U281 ( .A(neg_mul[22]), .B(N480), .S0(n99), .Y(out[15]) );
  MX2X1 U282 ( .A(neg_mul[23]), .B(N481), .S0(n99), .Y(out[16]) );
  NAND4BBX1 U283 ( .AN(n45), .BN(n46), .C(n214), .D(n267), .Y(N446) );
  NOR4BX1 U284 ( .AN(n211), .B(n50), .C(n51), .D(in_8bit[2]), .Y(n212) );
  NOR2X1 U285 ( .A(in_8bit[6]), .B(in_8bit[3]), .Y(n211) );
  NOR2X1 U286 ( .A(out[0]), .B(neg_mul[8]), .Y(n42) );
  NAND2BX1 U287 ( .AN(n42), .B(neg_mul[9]), .Y(n73) );
  NOR2X1 U288 ( .A(in_8bit[6]), .B(in_8bit[4]), .Y(n208) );
  NAND2X1 U289 ( .A(n160), .B(n158), .Y(n261) );
  NAND3BX1 U290 ( .AN(n100), .B(n213), .C(in_8bit[6]), .Y(n160) );
  NAND3X1 U291 ( .A(n212), .B(n55), .C(n101), .Y(n158) );
  NAND2X1 U292 ( .A(neg_mul[10]), .B(n77), .Y(n80) );
  NAND2X1 U293 ( .A(out[0]), .B(neg_mul[8]), .Y(n68) );
  NAND2X1 U294 ( .A(neg_mul[14]), .B(n88), .Y(n91) );
  AOI2BB2X4 U295 ( .B0(n20), .B1(n11), .A0N(n53), .A1N(n68), .Y(n69) );
  NOR3X4 U296 ( .A(n71), .B(n70), .C(n42), .Y(out[1]) );
  XNOR2X4 U297 ( .A(n84), .B(n6), .Y(out[4]) );
  XNOR2X4 U298 ( .A(n58), .B(n52), .Y(n85) );
  NOR2X4 U299 ( .A(n36), .B(n86), .Y(n87) );
  NOR3X4 U300 ( .A(n93), .B(n33), .C(n94), .Y(out[7]) );
  NOR2X4 U301 ( .A(n35), .B(n95), .Y(n96) );
  XNOR2X4 U302 ( .A(n96), .B(n7), .Y(out[9]) );
  NOR2X4 U303 ( .A(n37), .B(n95), .Y(n97) );
  XNOR2X4 U304 ( .A(n97), .B(n8), .Y(out[10]) );
  AND2X1 U305 ( .A(add_1_root_r112_carry_20_), .B(in_17bit_b[16]), .Y(
        add_1_root_r112_SUM_21_) );
  XOR2X1 U306 ( .A(in_17bit_b[16]), .B(add_1_root_r112_carry_20_), .Y(
        add_1_root_r112_SUM_20_) );
  AND2X1 U307 ( .A(add_1_root_r112_carry_19_), .B(in_17bit_b[15]), .Y(
        add_1_root_r112_carry_20_) );
  XOR2X1 U308 ( .A(in_17bit_b[15]), .B(add_1_root_r112_carry_19_), .Y(
        add_1_root_r112_SUM_19_) );
  AND2X1 U309 ( .A(add_1_root_r112_carry_18_), .B(in_17bit_b[14]), .Y(
        add_1_root_r112_carry_19_) );
  XOR2X1 U310 ( .A(in_17bit_b[14]), .B(add_1_root_r112_carry_18_), .Y(
        add_1_root_r112_SUM_18_) );
  AND2X1 U311 ( .A(add_1_root_r112_carry_17_), .B(in_17bit_b[13]), .Y(
        add_1_root_r112_carry_18_) );
  XOR2X1 U312 ( .A(in_17bit_b[13]), .B(add_1_root_r112_carry_17_), .Y(
        add_1_root_r112_SUM_17_) );
  AND2X1 U313 ( .A(add_2_root_r119_carry_21_), .B(in_17bit_b[16]), .Y(
        add_2_root_r119_SUM_22_) );
  XOR2X1 U314 ( .A(in_17bit_b[16]), .B(add_2_root_r119_carry_21_), .Y(
        add_2_root_r119_SUM_21_) );
  AND2X1 U315 ( .A(add_1_root_r119_carry[22]), .B(in_17bit_b[16]), .Y(
        add_1_root_r119_SUM_23_) );
  XOR2X1 U316 ( .A(in_17bit_b[16]), .B(add_1_root_r119_carry[22]), .Y(
        add_1_root_r119_SUM_22_) );
  AND2X1 U317 ( .A(add_1_root_r119_carry[21]), .B(in_17bit_b[15]), .Y(
        add_1_root_r119_carry[22]) );
  XOR2X1 U318 ( .A(in_17bit_b[15]), .B(add_1_root_r119_carry[21]), .Y(
        add_1_root_r119_SUM_21_) );
  AND2X1 U319 ( .A(add_1_root_r119_carry[20]), .B(in_17bit_b[14]), .Y(
        add_1_root_r119_carry[21]) );
  XOR2X1 U320 ( .A(in_17bit_b[14]), .B(add_1_root_r119_carry[20]), .Y(
        add_1_root_r119_SUM_20_) );
  AND2X1 U321 ( .A(add_1_root_r119_A_6_), .B(in_17bit_b[0]), .Y(
        add_1_root_r119_carry[7]) );
  XOR2X1 U322 ( .A(in_17bit_b[0]), .B(add_1_root_r119_A_6_), .Y(
        add_1_root_r119_SUM_6_) );
  AND2X1 U323 ( .A(add_3_root_r119_carry_18_), .B(in_17bit_b[16]), .Y(
        add_1_root_r119_A_19_) );
  XOR2X1 U324 ( .A(in_17bit_b[16]), .B(add_3_root_r119_carry_18_), .Y(
        add_1_root_r119_A_18_) );
  AND2X1 U325 ( .A(n187), .B(in_17bit_b[0]), .Y(add_3_root_r119_carry_3_) );
  XOR2X1 U326 ( .A(in_17bit_b[0]), .B(n187), .Y(add_1_root_r119_A_2_) );
  AND2X1 U327 ( .A(add_2_root_r115_carry_19_), .B(in_17bit_b[16]), .Y(
        add_2_root_r115_SUM_20_) );
  XOR2X1 U328 ( .A(in_17bit_b[16]), .B(add_2_root_r115_carry_19_), .Y(
        add_2_root_r115_SUM_19_) );
  AND2X1 U329 ( .A(add_2_root_r115_carry_18_), .B(in_17bit_b[15]), .Y(
        add_2_root_r115_carry_19_) );
  XOR2X1 U330 ( .A(in_17bit_b[15]), .B(add_2_root_r115_carry_18_), .Y(
        add_2_root_r115_SUM_18_) );
  AND2X1 U331 ( .A(add_1_root_r115_carry_22_), .B(in_17bit_b[16]), .Y(
        add_1_root_r115_SUM_23_) );
  XOR2X1 U332 ( .A(in_17bit_b[16]), .B(add_1_root_r115_carry_22_), .Y(
        add_1_root_r115_SUM_22_) );
  AND2X1 U333 ( .A(add_1_root_r115_carry_21_), .B(in_17bit_b[15]), .Y(
        add_1_root_r115_carry_22_) );
  XOR2X1 U334 ( .A(in_17bit_b[15]), .B(add_1_root_r115_carry_21_), .Y(
        add_1_root_r115_SUM_21_) );
  AND2X1 U335 ( .A(in_17bit_b[2]), .B(in_17bit_b[0]), .Y(
        add_1_root_r115_carry_7_) );
  XOR2X1 U336 ( .A(in_17bit_b[0]), .B(in_17bit_b[2]), .Y(
        add_1_root_r115_SUM_6_) );
  XOR2X1 U337 ( .A(n62), .B(sub_add_54_b0_carry[16]), .Y(N29) );
  AND2X1 U338 ( .A(sub_add_54_b0_carry[15]), .B(n186), .Y(
        sub_add_54_b0_carry[16]) );
  XOR2X1 U339 ( .A(n186), .B(sub_add_54_b0_carry[15]), .Y(N28) );
  AND2X1 U340 ( .A(sub_add_54_b0_carry[14]), .B(n185), .Y(
        sub_add_54_b0_carry[15]) );
  XOR2X1 U341 ( .A(n185), .B(sub_add_54_b0_carry[14]), .Y(N27) );
  AND2X1 U342 ( .A(sub_add_54_b0_carry[13]), .B(n184), .Y(
        sub_add_54_b0_carry[14]) );
  XOR2X1 U343 ( .A(n184), .B(sub_add_54_b0_carry[13]), .Y(N26) );
  AND2X1 U344 ( .A(sub_add_54_b0_carry[12]), .B(n183), .Y(
        sub_add_54_b0_carry[13]) );
  XOR2X1 U345 ( .A(n183), .B(sub_add_54_b0_carry[12]), .Y(N25) );
  AND2X1 U346 ( .A(sub_add_54_b0_carry[11]), .B(n182), .Y(
        sub_add_54_b0_carry[12]) );
  XOR2X1 U347 ( .A(n182), .B(sub_add_54_b0_carry[11]), .Y(N24) );
  AND2X1 U348 ( .A(sub_add_54_b0_carry[10]), .B(n181), .Y(
        sub_add_54_b0_carry[11]) );
  XOR2X1 U349 ( .A(n181), .B(sub_add_54_b0_carry[10]), .Y(N23) );
  AND2X1 U350 ( .A(sub_add_54_b0_carry[9]), .B(n180), .Y(
        sub_add_54_b0_carry[10]) );
  XOR2X1 U351 ( .A(n180), .B(sub_add_54_b0_carry[9]), .Y(N22) );
  AND2X1 U352 ( .A(sub_add_54_b0_carry[8]), .B(n179), .Y(
        sub_add_54_b0_carry[9]) );
  XOR2X1 U353 ( .A(n179), .B(sub_add_54_b0_carry[8]), .Y(N21) );
  AND2X1 U354 ( .A(sub_add_54_b0_carry[7]), .B(n178), .Y(
        sub_add_54_b0_carry[8]) );
  XOR2X1 U355 ( .A(n178), .B(sub_add_54_b0_carry[7]), .Y(N20) );
  AND2X1 U356 ( .A(sub_add_54_b0_carry[6]), .B(n177), .Y(
        sub_add_54_b0_carry[7]) );
  XOR2X1 U357 ( .A(n177), .B(sub_add_54_b0_carry[6]), .Y(N19) );
  AND2X1 U358 ( .A(sub_add_54_b0_carry[5]), .B(n176), .Y(
        sub_add_54_b0_carry[6]) );
  XOR2X1 U359 ( .A(n176), .B(sub_add_54_b0_carry[5]), .Y(N18) );
  AND2X1 U360 ( .A(sub_add_54_b0_carry[4]), .B(n175), .Y(
        sub_add_54_b0_carry[5]) );
  XOR2X1 U361 ( .A(n175), .B(sub_add_54_b0_carry[4]), .Y(N17) );
  AND2X1 U362 ( .A(sub_add_54_b0_carry[3]), .B(n174), .Y(
        sub_add_54_b0_carry[4]) );
  XOR2X1 U363 ( .A(n174), .B(sub_add_54_b0_carry[3]), .Y(N16) );
  AND2X1 U364 ( .A(sub_add_54_b0_carry[2]), .B(n173), .Y(
        sub_add_54_b0_carry[3]) );
  XOR2X1 U365 ( .A(n173), .B(sub_add_54_b0_carry[2]), .Y(N15) );
  AND2X1 U366 ( .A(n171), .B(n172), .Y(sub_add_54_b0_carry[2]) );
  XOR2X1 U367 ( .A(n172), .B(n171), .Y(N14) );
  XOR2X1 U368 ( .A(n16), .B(sub_add_75_b0_carry[16]), .Y(N481) );
  AND2X1 U369 ( .A(sub_add_75_b0_carry[15]), .B(n13), .Y(
        sub_add_75_b0_carry[16]) );
  XOR2X1 U370 ( .A(n13), .B(sub_add_75_b0_carry[15]), .Y(N480) );
  AND2X1 U371 ( .A(sub_add_75_b0_carry[14]), .B(n27), .Y(
        sub_add_75_b0_carry[15]) );
  AND2X1 U372 ( .A(sub_add_75_b0_carry[13]), .B(n15), .Y(
        sub_add_75_b0_carry[14]) );
  AND2X1 U373 ( .A(n40), .B(n14), .Y(sub_add_75_b0_carry[13]) );
  AND2X1 U374 ( .A(in_17bit_b[0]), .B(in_17bit_b[4]), .Y(
        add_1_root_r112_carry_5_) );
endmodule


module multi16_1_DW01_add_0 ( A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, 
        A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, 
        A_4_, B_23_, B_22_, B_21_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, 
        B_14_, B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, 
        SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, 
        SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, 
        SUM_7_ );
  input A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_,
         A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, B_23_, B_22_,
         B_21_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_,
         B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_;
  output SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_,
         SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_,
         SUM_8_, SUM_7_;
  wire   n1, n2, n3, n4;
  wire   [23:7] carry;

  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry[7]), .CO(carry[8]), .S(SUM_7_)
         );
  ADDFX2 U1_21 ( .A(A_21_), .B(B_21_), .CI(carry[21]), .CO(carry[22]), .S(
        SUM_21_) );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry[20]), .CO(carry[21]), .S(
        SUM_20_) );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry[19]), .CO(carry[20]), .S(
        SUM_19_) );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry[18]), .CO(carry[19]), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry[17]), .CO(carry[18]), .S(
        SUM_17_) );
  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry[16]), .CO(carry[17]), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry[15]), .CO(carry[16]), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry[14]), .CO(carry[15]), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry[13]), .CO(carry[14]), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry[12]), .CO(carry[13]), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry[11]), .CO(carry[12]), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry[10]), .CO(carry[11]), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry[9]), .CO(carry[10]), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry[8]), .CO(carry[9]), .S(SUM_8_)
         );
  ADDFX2 U1_22 ( .A(A_22_), .B(B_22_), .CI(carry[22]), .CO(carry[23]), .S(
        SUM_22_) );
  AND2X2 U1 ( .A(A_4_), .B(B_4_), .Y(n1) );
  XOR2X1 U2 ( .A(B_23_), .B(carry[23]), .Y(SUM_23_) );
  OAI2BB1X1 U3 ( .A0N(n2), .A1N(A_6_), .B0(n3), .Y(carry[7]) );
  OAI21XL U4 ( .A0(A_6_), .A1(n2), .B0(B_6_), .Y(n3) );
  OAI2BB1X1 U5 ( .A0N(n1), .A1N(A_5_), .B0(n4), .Y(n2) );
  OAI21XL U6 ( .A0(A_5_), .A1(n1), .B0(B_5_), .Y(n4) );
endmodule


module multi16_1_DW01_add_4 ( A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, 
        A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, 
        B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, 
        B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, SUM_22_, SUM_21_, SUM_20_, 
        SUM_19_, SUM_18_, SUM_17_, SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, 
        SUM_11_, SUM_10_, SUM_9_, SUM_8_, SUM_7_ );
  input A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_,
         A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, B_20_, B_19_,
         B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, B_10_, B_9_,
         B_8_, B_7_, B_6_, B_5_;
  output SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_,
         SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_,
         SUM_7_;
  wire   carry_21_, carry_20_, carry_19_, carry_18_, carry_17_, carry_16_,
         carry_15_, carry_14_, carry_13_, carry_12_, carry_11_, carry_10_,
         carry_9_, carry_8_, carry_7_, n1;

  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry_16_), .CO(carry_17_), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry_15_), .CO(carry_16_), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry_14_), .CO(carry_15_), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry_13_), .CO(carry_14_), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry_12_), .CO(carry_13_), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry_11_), .CO(carry_12_), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry_10_), .CO(carry_11_), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry_9_), .CO(carry_10_), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry_8_), .CO(carry_9_), .S(SUM_8_)
         );
  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry_7_), .CO(carry_8_), .S(SUM_7_)
         );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry_20_), .CO(carry_21_), .S(
        SUM_20_) );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry_19_), .CO(carry_20_), .S(
        SUM_19_) );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry_18_), .CO(carry_19_), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry_17_), .CO(carry_18_), .S(
        SUM_17_) );
  ADDFX2 U1_21 ( .A(A_21_), .B(B_21_), .CI(carry_21_), .CO(SUM_22_), .S(
        SUM_21_) );
  OAI2BB1X1 U1 ( .A0N(A_6_), .A1N(B_6_), .B0(n1), .Y(carry_7_) );
  OAI211X1 U2 ( .A0(B_6_), .A1(A_6_), .B0(A_5_), .C0(B_5_), .Y(n1) );
endmodule


module multi16_1_DW01_add_6 ( A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, 
        A_16_, A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, 
        A_6_, A_5_, A_4_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, 
        B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, 
        SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, 
        SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, 
        SUM_7_ );
  input A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_,
         A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, B_20_,
         B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, B_10_,
         B_9_, B_8_, B_7_, B_6_, B_5_, B_4_;
  output SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_,
         SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_,
         SUM_8_, SUM_7_;
  wire   n1, n2, n3, n4, n5, n6;
  wire   [21:7] carry;

  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry[7]), .CO(carry[8]), .S(SUM_7_)
         );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry[18]), .CO(carry[19]), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry[17]), .CO(carry[18]), .S(
        SUM_17_) );
  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry[16]), .CO(carry[17]), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry[15]), .CO(carry[16]), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry[14]), .CO(carry[15]), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry[13]), .CO(carry[14]), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry[12]), .CO(carry[13]), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry[11]), .CO(carry[12]), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry[10]), .CO(carry[11]), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry[9]), .CO(carry[10]), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry[8]), .CO(carry[9]), .S(SUM_8_)
         );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry[19]), .CO(carry[20]), .S(
        SUM_19_) );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry[20]), .CO(carry[21]), .S(
        SUM_20_) );
  AND2X2 U1 ( .A(A_22_), .B(n2), .Y(n1) );
  AND2X2 U2 ( .A(A_21_), .B(carry[21]), .Y(n2) );
  XOR2X1 U3 ( .A(A_23_), .B(n1), .Y(SUM_23_) );
  XOR2X1 U4 ( .A(A_21_), .B(carry[21]), .Y(SUM_21_) );
  XOR2X1 U5 ( .A(A_22_), .B(n2), .Y(SUM_22_) );
  AND2X2 U6 ( .A(A_4_), .B(B_4_), .Y(n3) );
  OAI2BB1X1 U7 ( .A0N(n4), .A1N(A_6_), .B0(n5), .Y(carry[7]) );
  OAI21XL U8 ( .A0(A_6_), .A1(n4), .B0(B_6_), .Y(n5) );
  OAI2BB1X1 U9 ( .A0N(n3), .A1N(A_5_), .B0(n6), .Y(n4) );
  OAI21XL U10 ( .A0(A_5_), .A1(n3), .B0(B_5_), .Y(n6) );
endmodule


module multi16_1 ( in_17bit, in_8bit, out );
  input [16:0] in_17bit;
  input [7:0] in_8bit;
  output [16:0] out;
  wire   N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27,
         N28, N29, N108, N109, N110, N111, N112, N113, N114, N115, N116, N117,
         N118, N119, N120, N121, N122, N123, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220,
         N221, N347, N348, N349, N350, N351, N352, N353, N354, N355, N356,
         N357, N358, N359, N360, N361, N362, N363, N446, N447, N448, N449,
         N450, N451, N452, N453, N454, N455, N456, N457, N458, N459, N460,
         N461, N462, N463, N479, N480, add_2_root_r119_carry_10_,
         add_2_root_r119_carry_11_, add_2_root_r119_carry_12_,
         add_2_root_r119_carry_13_, add_2_root_r119_carry_14_,
         add_2_root_r119_carry_15_, add_2_root_r119_carry_16_,
         add_2_root_r119_carry_17_, add_2_root_r119_carry_18_,
         add_2_root_r119_carry_19_, add_2_root_r119_carry_20_,
         add_2_root_r119_carry_21_, add_2_root_r119_carry_7_,
         add_2_root_r119_carry_8_, add_2_root_r119_carry_9_,
         add_2_root_r119_SUM_6_, add_2_root_r119_SUM_7_,
         add_2_root_r119_SUM_8_, add_2_root_r119_SUM_9_,
         add_2_root_r119_SUM_10_, add_2_root_r119_SUM_11_,
         add_2_root_r119_SUM_12_, add_2_root_r119_SUM_13_,
         add_2_root_r119_SUM_14_, add_2_root_r119_SUM_15_,
         add_2_root_r119_SUM_16_, add_2_root_r119_SUM_17_,
         add_2_root_r119_SUM_18_, add_2_root_r119_SUM_19_,
         add_2_root_r119_SUM_20_, add_2_root_r119_SUM_21_,
         add_2_root_r119_SUM_22_, add_1_root_r119_SUM_6_,
         add_1_root_r119_SUM_7_, add_1_root_r119_SUM_8_,
         add_1_root_r119_SUM_9_, add_1_root_r119_SUM_10_,
         add_1_root_r119_SUM_11_, add_1_root_r119_SUM_12_,
         add_1_root_r119_SUM_13_, add_1_root_r119_SUM_14_,
         add_1_root_r119_SUM_15_, add_1_root_r119_SUM_16_,
         add_1_root_r119_SUM_17_, add_1_root_r119_SUM_18_,
         add_1_root_r119_SUM_19_, add_1_root_r119_SUM_20_,
         add_1_root_r119_SUM_21_, add_1_root_r119_SUM_22_,
         add_1_root_r119_SUM_23_, add_1_root_r119_A_2_, add_1_root_r119_A_3_,
         add_1_root_r119_A_4_, add_1_root_r119_A_5_, add_1_root_r119_A_6_,
         add_1_root_r119_A_7_, add_1_root_r119_A_8_, add_1_root_r119_A_9_,
         add_1_root_r119_A_10_, add_1_root_r119_A_11_, add_1_root_r119_A_12_,
         add_1_root_r119_A_13_, add_1_root_r119_A_14_, add_1_root_r119_A_15_,
         add_1_root_r119_A_16_, add_1_root_r119_A_17_, add_1_root_r119_A_18_,
         add_1_root_r119_A_19_, add_3_root_r119_carry_10_,
         add_3_root_r119_carry_11_, add_3_root_r119_carry_12_,
         add_3_root_r119_carry_13_, add_3_root_r119_carry_14_,
         add_3_root_r119_carry_15_, add_3_root_r119_carry_16_,
         add_3_root_r119_carry_17_, add_3_root_r119_carry_18_,
         add_3_root_r119_carry_3_, add_3_root_r119_carry_4_,
         add_3_root_r119_carry_5_, add_3_root_r119_carry_6_,
         add_3_root_r119_carry_7_, add_3_root_r119_carry_8_,
         add_3_root_r119_carry_9_, add_1_root_r112_carry_10_,
         add_1_root_r112_carry_11_, add_1_root_r112_carry_12_,
         add_1_root_r112_carry_13_, add_1_root_r112_carry_14_,
         add_1_root_r112_carry_15_, add_1_root_r112_carry_16_,
         add_1_root_r112_carry_17_, add_1_root_r112_carry_18_,
         add_1_root_r112_carry_19_, add_1_root_r112_carry_20_,
         add_1_root_r112_carry_5_, add_1_root_r112_carry_6_,
         add_1_root_r112_carry_7_, add_1_root_r112_carry_8_,
         add_1_root_r112_carry_9_, add_1_root_r112_SUM_1_,
         add_1_root_r112_SUM_2_, add_1_root_r112_SUM_3_,
         add_1_root_r112_SUM_4_, add_1_root_r112_SUM_5_,
         add_1_root_r112_SUM_6_, add_1_root_r112_SUM_7_,
         add_1_root_r112_SUM_8_, add_1_root_r112_SUM_9_,
         add_1_root_r112_SUM_10_, add_1_root_r112_SUM_11_,
         add_1_root_r112_SUM_12_, add_1_root_r112_SUM_13_,
         add_1_root_r112_SUM_14_, add_1_root_r112_SUM_15_,
         add_1_root_r112_SUM_16_, add_1_root_r112_SUM_17_,
         add_1_root_r112_SUM_18_, add_1_root_r112_SUM_19_,
         add_1_root_r112_SUM_20_, add_1_root_r112_SUM_21_,
         add_2_root_r115_carry_10_, add_2_root_r115_carry_11_,
         add_2_root_r115_carry_12_, add_2_root_r115_carry_13_,
         add_2_root_r115_carry_14_, add_2_root_r115_carry_15_,
         add_2_root_r115_carry_16_, add_2_root_r115_carry_17_,
         add_2_root_r115_carry_18_, add_2_root_r115_carry_19_,
         add_2_root_r115_carry_5_, add_2_root_r115_carry_6_,
         add_2_root_r115_carry_7_, add_2_root_r115_carry_8_,
         add_2_root_r115_carry_9_, add_2_root_r115_SUM_4_,
         add_2_root_r115_SUM_5_, add_2_root_r115_SUM_6_,
         add_2_root_r115_SUM_7_, add_2_root_r115_SUM_8_,
         add_2_root_r115_SUM_9_, add_2_root_r115_SUM_10_,
         add_2_root_r115_SUM_11_, add_2_root_r115_SUM_12_,
         add_2_root_r115_SUM_13_, add_2_root_r115_SUM_14_,
         add_2_root_r115_SUM_15_, add_2_root_r115_SUM_16_,
         add_2_root_r115_SUM_17_, add_2_root_r115_SUM_18_,
         add_2_root_r115_SUM_19_, add_2_root_r115_SUM_20_,
         add_1_root_r115_carry_10_, add_1_root_r115_carry_11_,
         add_1_root_r115_carry_12_, add_1_root_r115_carry_13_,
         add_1_root_r115_carry_14_, add_1_root_r115_carry_15_,
         add_1_root_r115_carry_16_, add_1_root_r115_carry_17_,
         add_1_root_r115_carry_18_, add_1_root_r115_carry_19_,
         add_1_root_r115_carry_20_, add_1_root_r115_carry_21_,
         add_1_root_r115_carry_22_, add_1_root_r115_carry_7_,
         add_1_root_r115_carry_8_, add_1_root_r115_carry_9_,
         add_1_root_r115_SUM_6_, add_1_root_r115_SUM_7_,
         add_1_root_r115_SUM_8_, add_1_root_r115_SUM_9_,
         add_1_root_r115_SUM_10_, add_1_root_r115_SUM_11_,
         add_1_root_r115_SUM_12_, add_1_root_r115_SUM_13_,
         add_1_root_r115_SUM_14_, add_1_root_r115_SUM_15_,
         add_1_root_r115_SUM_16_, add_1_root_r115_SUM_17_,
         add_1_root_r115_SUM_18_, add_1_root_r115_SUM_19_,
         add_1_root_r115_SUM_20_, add_1_root_r115_SUM_21_,
         add_1_root_r115_SUM_22_, add_1_root_r115_SUM_23_, n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n158, n160, n161,
         n162, n163, n164, n167, n168, n170, n171, n172, n173, n174, n175,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254;
  wire   [16:0] in_17bit_b;
  wire   [23:8] neg_mul;
  wire   [15:13] sub_add_75_b0_carry;
  wire   [16:2] sub_add_54_b0_carry;
  wire   [22:7] add_1_root_r119_carry;

  multi16_1_DW01_add_0 add_0_root_r119 ( .A_22_(add_2_root_r119_SUM_22_), 
        .A_21_(add_2_root_r119_SUM_21_), .A_20_(add_2_root_r119_SUM_20_), 
        .A_19_(add_2_root_r119_SUM_19_), .A_18_(add_2_root_r119_SUM_18_), 
        .A_17_(add_2_root_r119_SUM_17_), .A_16_(add_2_root_r119_SUM_16_), 
        .A_15_(add_2_root_r119_SUM_15_), .A_14_(add_2_root_r119_SUM_14_), 
        .A_13_(add_2_root_r119_SUM_13_), .A_12_(add_2_root_r119_SUM_12_), 
        .A_11_(add_2_root_r119_SUM_11_), .A_10_(add_2_root_r119_SUM_10_), 
        .A_9_(add_2_root_r119_SUM_9_), .A_8_(add_2_root_r119_SUM_8_), .A_7_(
        add_2_root_r119_SUM_7_), .A_6_(add_2_root_r119_SUM_6_), .A_5_(
        add_1_root_r119_A_2_), .A_4_(in_17bit_b[0]), .B_23_(
        add_1_root_r119_SUM_23_), .B_22_(add_1_root_r119_SUM_22_), .B_21_(
        add_1_root_r119_SUM_21_), .B_20_(add_1_root_r119_SUM_20_), .B_19_(
        add_1_root_r119_SUM_19_), .B_18_(add_1_root_r119_SUM_18_), .B_17_(
        add_1_root_r119_SUM_17_), .B_16_(add_1_root_r119_SUM_16_), .B_15_(
        add_1_root_r119_SUM_15_), .B_14_(add_1_root_r119_SUM_14_), .B_13_(
        add_1_root_r119_SUM_13_), .B_12_(add_1_root_r119_SUM_12_), .B_11_(
        add_1_root_r119_SUM_11_), .B_10_(add_1_root_r119_SUM_10_), .B_9_(
        add_1_root_r119_SUM_9_), .B_8_(add_1_root_r119_SUM_8_), .B_7_(
        add_1_root_r119_SUM_7_), .B_6_(add_1_root_r119_SUM_6_), .B_5_(
        add_1_root_r119_A_5_), .B_4_(add_1_root_r119_A_4_), .SUM_23_(N363), 
        .SUM_22_(N362), .SUM_21_(N361), .SUM_20_(N360), .SUM_19_(N359), 
        .SUM_18_(N358), .SUM_17_(N357), .SUM_16_(N356), .SUM_15_(N355), 
        .SUM_14_(N354), .SUM_13_(N353), .SUM_12_(N352), .SUM_11_(N351), 
        .SUM_10_(N350), .SUM_9_(N349), .SUM_8_(N348), .SUM_7_(N347) );
  multi16_1_DW01_add_4 add_0_root_r112 ( .A_21_(in_17bit_b[16]), .A_20_(
        in_17bit_b[15]), .A_19_(in_17bit_b[14]), .A_18_(in_17bit_b[13]), 
        .A_17_(in_17bit_b[12]), .A_16_(in_17bit_b[11]), .A_15_(in_17bit_b[10]), 
        .A_14_(in_17bit_b[9]), .A_13_(in_17bit_b[8]), .A_12_(in_17bit_b[7]), 
        .A_11_(in_17bit_b[6]), .A_10_(in_17bit_b[5]), .A_9_(in_17bit_b[4]), 
        .A_8_(in_17bit_b[3]), .A_7_(in_17bit_b[2]), .A_6_(in_17bit_b[1]), 
        .A_5_(in_17bit_b[0]), .B_21_(add_1_root_r112_SUM_21_), .B_20_(
        add_1_root_r112_SUM_20_), .B_19_(add_1_root_r112_SUM_19_), .B_18_(
        add_1_root_r112_SUM_18_), .B_17_(add_1_root_r112_SUM_17_), .B_16_(
        add_1_root_r112_SUM_16_), .B_15_(add_1_root_r112_SUM_15_), .B_14_(
        add_1_root_r112_SUM_14_), .B_13_(add_1_root_r112_SUM_13_), .B_12_(
        add_1_root_r112_SUM_12_), .B_11_(add_1_root_r112_SUM_11_), .B_10_(
        add_1_root_r112_SUM_10_), .B_9_(add_1_root_r112_SUM_9_), .B_8_(
        add_1_root_r112_SUM_8_), .B_7_(add_1_root_r112_SUM_7_), .B_6_(
        add_1_root_r112_SUM_6_), .B_5_(add_1_root_r112_SUM_5_), .SUM_22_(N123), 
        .SUM_21_(N122), .SUM_20_(N121), .SUM_19_(N120), .SUM_18_(N119), 
        .SUM_17_(N118), .SUM_16_(N117), .SUM_15_(N116), .SUM_14_(N115), 
        .SUM_13_(N114), .SUM_12_(N113), .SUM_11_(N112), .SUM_10_(N111), 
        .SUM_9_(N110), .SUM_8_(N109), .SUM_7_(N108) );
  multi16_1_DW01_add_6 add_0_root_r115 ( .A_23_(add_1_root_r115_SUM_23_), 
        .A_22_(add_1_root_r115_SUM_22_), .A_21_(add_1_root_r115_SUM_21_), 
        .A_20_(add_1_root_r115_SUM_20_), .A_19_(add_1_root_r115_SUM_19_), 
        .A_18_(add_1_root_r115_SUM_18_), .A_17_(add_1_root_r115_SUM_17_), 
        .A_16_(add_1_root_r115_SUM_16_), .A_15_(add_1_root_r115_SUM_15_), 
        .A_14_(add_1_root_r115_SUM_14_), .A_13_(add_1_root_r115_SUM_13_), 
        .A_12_(add_1_root_r115_SUM_12_), .A_11_(add_1_root_r115_SUM_11_), 
        .A_10_(add_1_root_r115_SUM_10_), .A_9_(add_1_root_r115_SUM_9_), .A_8_(
        add_1_root_r115_SUM_8_), .A_7_(add_1_root_r115_SUM_7_), .A_6_(
        add_1_root_r115_SUM_6_), .A_5_(in_17bit_b[1]), .A_4_(in_17bit_b[0]), 
        .B_20_(add_2_root_r115_SUM_20_), .B_19_(add_2_root_r115_SUM_19_), 
        .B_18_(add_2_root_r115_SUM_18_), .B_17_(add_2_root_r115_SUM_17_), 
        .B_16_(add_2_root_r115_SUM_16_), .B_15_(add_2_root_r115_SUM_15_), 
        .B_14_(add_2_root_r115_SUM_14_), .B_13_(add_2_root_r115_SUM_13_), 
        .B_12_(add_2_root_r115_SUM_12_), .B_11_(add_2_root_r115_SUM_11_), 
        .B_10_(add_2_root_r115_SUM_10_), .B_9_(add_2_root_r115_SUM_9_), .B_8_(
        add_2_root_r115_SUM_8_), .B_7_(add_2_root_r115_SUM_7_), .B_6_(
        add_2_root_r115_SUM_6_), .B_5_(add_2_root_r115_SUM_5_), .B_4_(
        add_2_root_r115_SUM_4_), .SUM_23_(N221), .SUM_22_(N220), .SUM_21_(N219), .SUM_20_(N218), .SUM_19_(N217), .SUM_18_(N216), .SUM_17_(N215), .SUM_16_(
        N214), .SUM_15_(N213), .SUM_14_(N212), .SUM_13_(N211), .SUM_12_(N210), 
        .SUM_11_(N209), .SUM_10_(N208), .SUM_9_(N207), .SUM_8_(N206), .SUM_7_(
        N205) );
  TLATX1 neg_mul_reg_19_ ( .G(N446), .D(N459), .QN(n10) );
  TLATX1 neg_mul_reg_18_ ( .G(N446), .D(N458), .QN(n9) );
  TLATX1 neg_mul_reg_17_ ( .G(N446), .D(N457), .QN(n3) );
  TLATX1 neg_mul_reg_16_ ( .G(N446), .D(N456), .QN(n2) );
  TLATX1 neg_mul_reg_15_ ( .G(N446), .D(N455), .QN(n4) );
  TLATX1 neg_mul_reg_14_ ( .G(N446), .D(N454), .QN(n8) );
  TLATX1 neg_mul_reg_13_ ( .G(N446), .D(N453), .QN(n7) );
  TLATX1 neg_mul_reg_12_ ( .G(N446), .D(N452), .QN(n6) );
  TLATX1 neg_mul_reg_11_ ( .G(N446), .D(N451), .QN(n5) );
  TLATX1 neg_mul_reg_23_ ( .G(N446), .D(N463), .Q(neg_mul[23]), .QN(n1) );
  TLATX1 neg_mul_reg_22_ ( .G(N446), .D(N462), .Q(neg_mul[22]), .QN(n13) );
  TLATX1 neg_mul_reg_21_ ( .G(N446), .D(N461), .Q(neg_mul[21]), .QN(n14) );
  TLATX1 neg_mul_reg_20_ ( .G(N446), .D(N460), .QN(n16) );
  TLATX1 neg_mul_reg_9_ ( .G(N446), .D(N449), .Q(neg_mul[9]), .QN(n11) );
  TLATX1 neg_mul_reg_10_ ( .G(N446), .D(N450), .Q(neg_mul[10]), .QN(n12) );
  TLATX1 neg_mul_reg_8_ ( .G(N446), .D(N448), .Q(neg_mul[8]), .QN(n15) );
  TLATX1 neg_mul_reg_7_ ( .G(N446), .D(N447), .Q(out[0]) );
  CLKINVX3 U2 ( .A(n254), .Y(in_17bit_b[16]) );
  OAI21X1 U3 ( .A0(n46), .A1(n57), .B0(n56), .Y(n61) );
  NOR2X4 U4 ( .A(n28), .B(n78), .Y(n79) );
  INVX4 U5 ( .A(n81), .Y(n85) );
  MXI2X2 U6 ( .A(n16), .B(n37), .S0(n85), .Y(out[13]) );
  AOI2BB2X2 U7 ( .B0(n58), .B1(n46), .A0N(n47), .A1N(neg_mul[8]), .Y(n59) );
  AOI2BB2X2 U8 ( .B0(n72), .B1(n46), .A0N(n47), .A1N(neg_mul[10]), .Y(n73) );
  NAND2X2 U9 ( .A(n46), .B(n15), .Y(n56) );
  NAND2X2 U10 ( .A(n46), .B(n11), .Y(n62) );
  INVX1 U11 ( .A(n95), .Y(n91) );
  CLKINVX4 U12 ( .A(n48), .Y(n47) );
  NOR2XL U13 ( .A(n73), .B(in_17bit[16]), .Y(n74) );
  XNOR2X1 U14 ( .A(neg_mul[23]), .B(n39), .Y(n17) );
  XNOR2X4 U15 ( .A(n19), .B(n46), .Y(n81) );
  OAI21X1 U16 ( .A0(n46), .A1(n63), .B0(n62), .Y(n68) );
  NOR2X4 U17 ( .A(n29), .B(n83), .Y(n80) );
  NOR2X4 U18 ( .A(n53), .B(n59), .Y(n60) );
  INVX8 U19 ( .A(n51), .Y(n53) );
  INVXL U20 ( .A(n19), .Y(n18) );
  INVX8 U21 ( .A(in_8bit[7]), .Y(n48) );
  INVX8 U22 ( .A(in_17bit[16]), .Y(n51) );
  NOR2BX2 U23 ( .AN(n51), .B(n65), .Y(n67) );
  INVX8 U24 ( .A(n51), .Y(n19) );
  OR2X2 U25 ( .A(n33), .B(n83), .Y(n26) );
  XOR2X4 U26 ( .A(n27), .B(n2), .Y(out[9]) );
  XNOR2X2 U27 ( .A(n19), .B(n46), .Y(n78) );
  AOI2BB2X2 U28 ( .B0(n64), .B1(n46), .A0N(n47), .A1N(neg_mul[9]), .Y(n65) );
  AOI211X4 U29 ( .A0(n19), .A1(n75), .B0(n74), .C0(n76), .Y(out[3]) );
  XNOR2X4 U30 ( .A(n20), .B(n4), .Y(out[8]) );
  OAI21X1 U31 ( .A0(n46), .A1(n71), .B0(n70), .Y(n75) );
  NAND2X2 U32 ( .A(n46), .B(n12), .Y(n70) );
  XOR2X4 U33 ( .A(n26), .B(n3), .Y(out[10]) );
  OR2X2 U34 ( .A(n32), .B(n83), .Y(n27) );
  NOR2X4 U35 ( .A(n30), .B(n81), .Y(n82) );
  AOI211X4 U36 ( .A0(n53), .A1(n61), .B0(n60), .C0(n38), .Y(out[1]) );
  NOR2X2 U37 ( .A(n76), .B(n83), .Y(n77) );
  NOR2X2 U38 ( .A(n34), .B(n83), .Y(n84) );
  NOR2X2 U39 ( .A(n31), .B(n83), .Y(n20) );
  XNOR2X4 U40 ( .A(n53), .B(n46), .Y(n83) );
  CLKINVX20 U41 ( .A(n48), .Y(n46) );
  AND3X1 U42 ( .A(in_8bit[2]), .B(n45), .C(n43), .Y(n35) );
  NOR4XL U43 ( .A(in_8bit[1]), .B(in_8bit[0]), .C(in_8bit[2]), .D(in_8bit[3]), 
        .Y(n23) );
  MX2X1 U44 ( .A(neg_mul[21]), .B(N479), .S0(n85), .Y(out[14]) );
  INVX1 U45 ( .A(n204), .Y(in_17bit_b[1]) );
  INVX1 U46 ( .A(n243), .Y(in_17bit_b[14]) );
  INVX1 U47 ( .A(n240), .Y(in_17bit_b[13]) );
  INVX1 U48 ( .A(n207), .Y(in_17bit_b[2]) );
  INVX1 U49 ( .A(n216), .Y(in_17bit_b[5]) );
  INVX1 U50 ( .A(n219), .Y(in_17bit_b[6]) );
  INVX1 U51 ( .A(n222), .Y(in_17bit_b[7]) );
  INVX1 U52 ( .A(n225), .Y(in_17bit_b[8]) );
  INVX1 U53 ( .A(n228), .Y(in_17bit_b[9]) );
  INVX1 U54 ( .A(n231), .Y(in_17bit_b[10]) );
  INVX1 U55 ( .A(n234), .Y(in_17bit_b[11]) );
  INVX1 U56 ( .A(n237), .Y(in_17bit_b[12]) );
  INVX1 U57 ( .A(n213), .Y(in_17bit_b[4]) );
  INVX1 U58 ( .A(n210), .Y(in_17bit_b[3]) );
  XNOR2X4 U59 ( .A(n21), .B(n10), .Y(out[12]) );
  NOR2X2 U60 ( .A(n78), .B(n36), .Y(n21) );
  AOI21X1 U61 ( .A0(n22), .A1(n23), .B0(n247), .Y(n200) );
  NOR4XL U62 ( .A(in_8bit[4]), .B(n43), .C(in_8bit[6]), .D(n47), .Y(n22) );
  AND4X1 U63 ( .A(in_8bit[1]), .B(n47), .C(n195), .D(n49), .Y(n24) );
  INVX1 U64 ( .A(n18), .Y(n52) );
  INVX1 U65 ( .A(n52), .Y(n54) );
  INVX1 U66 ( .A(n174), .Y(n253) );
  NAND3XL U67 ( .A(n46), .B(n50), .C(n44), .Y(n94) );
  OAI21XL U68 ( .A0(n253), .A1(n254), .B0(n252), .Y(N463) );
  AOI22X1 U69 ( .A0(N221), .A1(n42), .B0(N363), .B1(n41), .Y(n252) );
  ADDFX2 U70 ( .A(in_17bit_b[16]), .B(in_17bit_b[12]), .CI(
        add_1_root_r112_carry_16_), .CO(add_1_root_r112_carry_17_), .S(
        add_1_root_r112_SUM_16_) );
  ADDFX2 U71 ( .A(add_1_root_r119_A_19_), .B(in_17bit_b[13]), .CI(
        add_1_root_r119_carry[19]), .CO(add_1_root_r119_carry[20]), .S(
        add_1_root_r119_SUM_19_) );
  ADDFX2 U72 ( .A(in_17bit_b[16]), .B(in_17bit_b[15]), .CI(
        add_3_root_r119_carry_17_), .CO(add_3_root_r119_carry_18_), .S(
        add_1_root_r119_A_17_) );
  ADDFX2 U73 ( .A(in_17bit_b[16]), .B(in_17bit_b[14]), .CI(
        add_2_root_r115_carry_17_), .CO(add_2_root_r115_carry_18_), .S(
        add_2_root_r115_SUM_17_) );
  ADDFX2 U74 ( .A(in_17bit_b[16]), .B(in_17bit_b[14]), .CI(
        add_1_root_r115_carry_20_), .CO(add_1_root_r115_carry_21_), .S(
        add_1_root_r115_SUM_20_) );
  ADDFX2 U75 ( .A(in_17bit_b[16]), .B(in_17bit_b[15]), .CI(
        add_2_root_r119_carry_20_), .CO(add_2_root_r119_carry_21_), .S(
        add_2_root_r119_SUM_20_) );
  ADDFX2 U76 ( .A(in_17bit_b[3]), .B(in_17bit_b[1]), .CI(
        add_1_root_r115_carry_7_), .CO(add_2_root_r115_carry_5_), .S(
        add_2_root_r115_SUM_4_) );
  ADDFX2 U77 ( .A(in_17bit_b[4]), .B(in_17bit_b[2]), .CI(
        add_2_root_r115_carry_5_), .CO(add_2_root_r115_carry_6_), .S(
        add_2_root_r115_SUM_5_) );
  ADDFX2 U78 ( .A(in_17bit_b[5]), .B(in_17bit_b[1]), .CI(
        add_1_root_r112_carry_5_), .CO(add_1_root_r112_carry_6_), .S(
        add_1_root_r112_SUM_5_) );
  ADDFX2 U79 ( .A(in_17bit_b[6]), .B(in_17bit_b[5]), .CI(
        add_3_root_r119_carry_7_), .CO(add_3_root_r119_carry_8_), .S(
        add_1_root_r119_A_7_) );
  ADDFX2 U80 ( .A(in_17bit_b[6]), .B(in_17bit_b[2]), .CI(
        add_1_root_r112_carry_6_), .CO(add_1_root_r112_carry_7_), .S(
        add_1_root_r112_SUM_6_) );
  ADDFX2 U81 ( .A(in_17bit_b[3]), .B(in_17bit_b[1]), .CI(
        add_1_root_r115_carry_7_), .CO(add_1_root_r115_carry_8_), .S(
        add_1_root_r115_SUM_7_) );
  ADDFX2 U82 ( .A(in_17bit_b[7]), .B(in_17bit_b[6]), .CI(
        add_3_root_r119_carry_8_), .CO(add_3_root_r119_carry_9_), .S(
        add_1_root_r119_A_8_) );
  ADDFX2 U83 ( .A(add_1_root_r119_A_7_), .B(in_17bit_b[1]), .CI(
        add_1_root_r119_carry[7]), .CO(add_1_root_r119_carry[8]), .S(
        add_1_root_r119_SUM_7_) );
  ADDFX2 U84 ( .A(in_17bit_b[2]), .B(in_17bit_b[1]), .CI(
        add_3_root_r119_carry_3_), .CO(add_2_root_r119_carry_7_), .S(
        add_2_root_r119_SUM_6_) );
  ADDFX2 U85 ( .A(in_17bit_b[4]), .B(in_17bit_b[2]), .CI(
        add_1_root_r115_carry_8_), .CO(add_1_root_r115_carry_9_), .S(
        add_1_root_r115_SUM_8_) );
  ADDFX2 U86 ( .A(in_17bit_b[8]), .B(in_17bit_b[7]), .CI(
        add_3_root_r119_carry_9_), .CO(add_3_root_r119_carry_10_), .S(
        add_1_root_r119_A_9_) );
  ADDFX2 U87 ( .A(add_1_root_r119_A_8_), .B(in_17bit_b[2]), .CI(
        add_1_root_r119_carry[8]), .CO(add_1_root_r119_carry[9]), .S(
        add_1_root_r119_SUM_8_) );
  ADDFX2 U88 ( .A(in_17bit_b[3]), .B(in_17bit_b[2]), .CI(
        add_2_root_r119_carry_7_), .CO(add_2_root_r119_carry_8_), .S(
        add_2_root_r119_SUM_7_) );
  ADDFX2 U89 ( .A(in_17bit_b[6]), .B(in_17bit_b[4]), .CI(
        add_2_root_r115_carry_7_), .CO(add_2_root_r115_carry_8_), .S(
        add_2_root_r115_SUM_7_) );
  ADDFX2 U90 ( .A(in_17bit_b[8]), .B(in_17bit_b[4]), .CI(
        add_1_root_r112_carry_8_), .CO(add_1_root_r112_carry_9_), .S(
        add_1_root_r112_SUM_8_) );
  ADDFX2 U91 ( .A(in_17bit_b[9]), .B(in_17bit_b[8]), .CI(
        add_3_root_r119_carry_10_), .CO(add_3_root_r119_carry_11_), .S(
        add_1_root_r119_A_10_) );
  ADDFX2 U92 ( .A(in_17bit_b[7]), .B(in_17bit_b[5]), .CI(
        add_2_root_r115_carry_8_), .CO(add_2_root_r115_carry_9_), .S(
        add_2_root_r115_SUM_8_) );
  ADDFX2 U93 ( .A(in_17bit_b[9]), .B(in_17bit_b[5]), .CI(
        add_1_root_r112_carry_9_), .CO(add_1_root_r112_carry_10_), .S(
        add_1_root_r112_SUM_9_) );
  ADDFX2 U94 ( .A(in_17bit_b[6]), .B(in_17bit_b[4]), .CI(
        add_1_root_r115_carry_10_), .CO(add_1_root_r115_carry_11_), .S(
        add_1_root_r115_SUM_10_) );
  ADDFX2 U95 ( .A(in_17bit_b[10]), .B(in_17bit_b[9]), .CI(
        add_3_root_r119_carry_11_), .CO(add_3_root_r119_carry_12_), .S(
        add_1_root_r119_A_11_) );
  ADDFX2 U96 ( .A(add_1_root_r119_A_10_), .B(in_17bit_b[4]), .CI(
        add_1_root_r119_carry[10]), .CO(add_1_root_r119_carry[11]), .S(
        add_1_root_r119_SUM_10_) );
  ADDFX2 U97 ( .A(in_17bit_b[5]), .B(in_17bit_b[4]), .CI(
        add_2_root_r119_carry_9_), .CO(add_2_root_r119_carry_10_), .S(
        add_2_root_r119_SUM_9_) );
  ADDFX2 U98 ( .A(in_17bit_b[8]), .B(in_17bit_b[6]), .CI(
        add_2_root_r115_carry_9_), .CO(add_2_root_r115_carry_10_), .S(
        add_2_root_r115_SUM_9_) );
  ADDFX2 U99 ( .A(in_17bit_b[10]), .B(in_17bit_b[6]), .CI(
        add_1_root_r112_carry_10_), .CO(add_1_root_r112_carry_11_), .S(
        add_1_root_r112_SUM_10_) );
  ADDFX2 U100 ( .A(in_17bit_b[7]), .B(in_17bit_b[5]), .CI(
        add_1_root_r115_carry_11_), .CO(add_1_root_r115_carry_12_), .S(
        add_1_root_r115_SUM_11_) );
  ADDFX2 U101 ( .A(in_17bit_b[11]), .B(in_17bit_b[10]), .CI(
        add_3_root_r119_carry_12_), .CO(add_3_root_r119_carry_13_), .S(
        add_1_root_r119_A_12_) );
  ADDFX2 U102 ( .A(add_1_root_r119_A_11_), .B(in_17bit_b[5]), .CI(
        add_1_root_r119_carry[11]), .CO(add_1_root_r119_carry[12]), .S(
        add_1_root_r119_SUM_11_) );
  ADDFX2 U103 ( .A(in_17bit_b[6]), .B(in_17bit_b[5]), .CI(
        add_2_root_r119_carry_10_), .CO(add_2_root_r119_carry_11_), .S(
        add_2_root_r119_SUM_10_) );
  ADDFX2 U104 ( .A(in_17bit_b[9]), .B(in_17bit_b[7]), .CI(
        add_2_root_r115_carry_10_), .CO(add_2_root_r115_carry_11_), .S(
        add_2_root_r115_SUM_10_) );
  ADDFX2 U105 ( .A(in_17bit_b[11]), .B(in_17bit_b[7]), .CI(
        add_1_root_r112_carry_11_), .CO(add_1_root_r112_carry_12_), .S(
        add_1_root_r112_SUM_11_) );
  ADDFX2 U106 ( .A(in_17bit_b[8]), .B(in_17bit_b[6]), .CI(
        add_1_root_r115_carry_12_), .CO(add_1_root_r115_carry_13_), .S(
        add_1_root_r115_SUM_12_) );
  ADDFX2 U107 ( .A(in_17bit_b[12]), .B(in_17bit_b[11]), .CI(
        add_3_root_r119_carry_13_), .CO(add_3_root_r119_carry_14_), .S(
        add_1_root_r119_A_13_) );
  ADDFX2 U108 ( .A(add_1_root_r119_A_12_), .B(in_17bit_b[6]), .CI(
        add_1_root_r119_carry[12]), .CO(add_1_root_r119_carry[13]), .S(
        add_1_root_r119_SUM_12_) );
  ADDFX2 U109 ( .A(in_17bit_b[7]), .B(in_17bit_b[6]), .CI(
        add_2_root_r119_carry_11_), .CO(add_2_root_r119_carry_12_), .S(
        add_2_root_r119_SUM_11_) );
  ADDFX2 U110 ( .A(in_17bit_b[10]), .B(in_17bit_b[8]), .CI(
        add_2_root_r115_carry_11_), .CO(add_2_root_r115_carry_12_), .S(
        add_2_root_r115_SUM_11_) );
  ADDFX2 U111 ( .A(in_17bit_b[12]), .B(in_17bit_b[8]), .CI(
        add_1_root_r112_carry_12_), .CO(add_1_root_r112_carry_13_), .S(
        add_1_root_r112_SUM_12_) );
  ADDFX2 U112 ( .A(in_17bit_b[9]), .B(in_17bit_b[7]), .CI(
        add_1_root_r115_carry_13_), .CO(add_1_root_r115_carry_14_), .S(
        add_1_root_r115_SUM_13_) );
  ADDFX2 U113 ( .A(in_17bit_b[13]), .B(in_17bit_b[12]), .CI(
        add_3_root_r119_carry_14_), .CO(add_3_root_r119_carry_15_), .S(
        add_1_root_r119_A_14_) );
  ADDFX2 U114 ( .A(add_1_root_r119_A_13_), .B(in_17bit_b[7]), .CI(
        add_1_root_r119_carry[13]), .CO(add_1_root_r119_carry[14]), .S(
        add_1_root_r119_SUM_13_) );
  ADDFX2 U115 ( .A(in_17bit_b[8]), .B(in_17bit_b[7]), .CI(
        add_2_root_r119_carry_12_), .CO(add_2_root_r119_carry_13_), .S(
        add_2_root_r119_SUM_12_) );
  ADDFX2 U116 ( .A(in_17bit_b[11]), .B(in_17bit_b[9]), .CI(
        add_2_root_r115_carry_12_), .CO(add_2_root_r115_carry_13_), .S(
        add_2_root_r115_SUM_12_) );
  ADDFX2 U117 ( .A(in_17bit_b[13]), .B(in_17bit_b[9]), .CI(
        add_1_root_r112_carry_13_), .CO(add_1_root_r112_carry_14_), .S(
        add_1_root_r112_SUM_13_) );
  ADDFX2 U118 ( .A(in_17bit_b[10]), .B(in_17bit_b[8]), .CI(
        add_1_root_r115_carry_14_), .CO(add_1_root_r115_carry_15_), .S(
        add_1_root_r115_SUM_14_) );
  ADDFX2 U119 ( .A(in_17bit_b[14]), .B(in_17bit_b[13]), .CI(
        add_3_root_r119_carry_15_), .CO(add_3_root_r119_carry_16_), .S(
        add_1_root_r119_A_15_) );
  ADDFX2 U120 ( .A(add_1_root_r119_A_14_), .B(in_17bit_b[8]), .CI(
        add_1_root_r119_carry[14]), .CO(add_1_root_r119_carry[15]), .S(
        add_1_root_r119_SUM_14_) );
  ADDFX2 U121 ( .A(in_17bit_b[9]), .B(in_17bit_b[8]), .CI(
        add_2_root_r119_carry_13_), .CO(add_2_root_r119_carry_14_), .S(
        add_2_root_r119_SUM_13_) );
  ADDFX2 U122 ( .A(in_17bit_b[12]), .B(in_17bit_b[10]), .CI(
        add_2_root_r115_carry_13_), .CO(add_2_root_r115_carry_14_), .S(
        add_2_root_r115_SUM_13_) );
  ADDFX2 U123 ( .A(in_17bit_b[14]), .B(in_17bit_b[10]), .CI(
        add_1_root_r112_carry_14_), .CO(add_1_root_r112_carry_15_), .S(
        add_1_root_r112_SUM_14_) );
  ADDFX2 U124 ( .A(in_17bit_b[11]), .B(in_17bit_b[9]), .CI(
        add_1_root_r115_carry_15_), .CO(add_1_root_r115_carry_16_), .S(
        add_1_root_r115_SUM_15_) );
  ADDFX2 U125 ( .A(add_1_root_r119_A_15_), .B(in_17bit_b[9]), .CI(
        add_1_root_r119_carry[15]), .CO(add_1_root_r119_carry[16]), .S(
        add_1_root_r119_SUM_15_) );
  ADDFX2 U126 ( .A(in_17bit_b[3]), .B(in_17bit_b[2]), .CI(
        add_3_root_r119_carry_4_), .CO(add_3_root_r119_carry_5_), .S(
        add_1_root_r119_A_4_) );
  ADDFX2 U127 ( .A(in_17bit_b[2]), .B(in_17bit_b[1]), .CI(
        add_3_root_r119_carry_3_), .CO(add_3_root_r119_carry_4_), .S(
        add_1_root_r119_A_3_) );
  ADDFX2 U128 ( .A(in_17bit_b[13]), .B(in_17bit_b[11]), .CI(
        add_2_root_r115_carry_14_), .CO(add_2_root_r115_carry_15_), .S(
        add_2_root_r115_SUM_14_) );
  ADDFX2 U129 ( .A(in_17bit_b[15]), .B(in_17bit_b[11]), .CI(
        add_1_root_r112_carry_15_), .CO(add_1_root_r112_carry_16_), .S(
        add_1_root_r112_SUM_15_) );
  ADDFX2 U130 ( .A(in_17bit_b[12]), .B(in_17bit_b[10]), .CI(
        add_1_root_r115_carry_16_), .CO(add_1_root_r115_carry_17_), .S(
        add_1_root_r115_SUM_16_) );
  ADDFX2 U131 ( .A(add_1_root_r119_A_16_), .B(in_17bit_b[10]), .CI(
        add_1_root_r119_carry[16]), .CO(add_1_root_r119_carry[17]), .S(
        add_1_root_r119_SUM_16_) );
  ADDFX2 U132 ( .A(in_17bit_b[11]), .B(in_17bit_b[10]), .CI(
        add_2_root_r119_carry_15_), .CO(add_2_root_r119_carry_16_), .S(
        add_2_root_r119_SUM_15_) );
  ADDFX2 U133 ( .A(in_17bit_b[14]), .B(in_17bit_b[12]), .CI(
        add_2_root_r115_carry_15_), .CO(add_2_root_r115_carry_16_), .S(
        add_2_root_r115_SUM_15_) );
  ADDFX2 U134 ( .A(in_17bit_b[13]), .B(in_17bit_b[11]), .CI(
        add_1_root_r115_carry_17_), .CO(add_1_root_r115_carry_18_), .S(
        add_1_root_r115_SUM_17_) );
  ADDFX2 U135 ( .A(add_1_root_r119_A_17_), .B(in_17bit_b[11]), .CI(
        add_1_root_r119_carry[17]), .CO(add_1_root_r119_carry[18]), .S(
        add_1_root_r119_SUM_17_) );
  ADDFX2 U136 ( .A(in_17bit_b[12]), .B(in_17bit_b[11]), .CI(
        add_2_root_r119_carry_16_), .CO(add_2_root_r119_carry_17_), .S(
        add_2_root_r119_SUM_16_) );
  ADDFX2 U137 ( .A(in_17bit_b[14]), .B(in_17bit_b[12]), .CI(
        add_1_root_r115_carry_18_), .CO(add_1_root_r115_carry_19_), .S(
        add_1_root_r115_SUM_18_) );
  ADDFX2 U138 ( .A(add_1_root_r119_A_18_), .B(in_17bit_b[12]), .CI(
        add_1_root_r119_carry[18]), .CO(add_1_root_r119_carry[19]), .S(
        add_1_root_r119_SUM_18_) );
  ADDFX2 U139 ( .A(in_17bit_b[13]), .B(in_17bit_b[12]), .CI(
        add_2_root_r119_carry_17_), .CO(add_2_root_r119_carry_18_), .S(
        add_2_root_r119_SUM_17_) );
  ADDFX2 U140 ( .A(in_17bit_b[15]), .B(in_17bit_b[13]), .CI(
        add_2_root_r115_carry_16_), .CO(add_2_root_r115_carry_17_), .S(
        add_2_root_r115_SUM_16_) );
  ADDFX2 U141 ( .A(in_17bit_b[15]), .B(in_17bit_b[13]), .CI(
        add_1_root_r115_carry_19_), .CO(add_1_root_r115_carry_20_), .S(
        add_1_root_r115_SUM_19_) );
  ADDFX2 U142 ( .A(in_17bit_b[14]), .B(in_17bit_b[13]), .CI(
        add_2_root_r119_carry_18_), .CO(add_2_root_r119_carry_19_), .S(
        add_2_root_r119_SUM_18_) );
  ADDFX2 U143 ( .A(in_17bit_b[5]), .B(in_17bit_b[3]), .CI(
        add_2_root_r115_carry_6_), .CO(add_2_root_r115_carry_7_), .S(
        add_2_root_r115_SUM_6_) );
  ADDFX2 U144 ( .A(in_17bit_b[7]), .B(in_17bit_b[3]), .CI(
        add_1_root_r112_carry_7_), .CO(add_1_root_r112_carry_8_), .S(
        add_1_root_r112_SUM_7_) );
  ADDFX2 U145 ( .A(in_17bit_b[5]), .B(in_17bit_b[3]), .CI(
        add_1_root_r115_carry_9_), .CO(add_1_root_r115_carry_10_), .S(
        add_1_root_r115_SUM_9_) );
  ADDFX2 U146 ( .A(add_1_root_r119_A_9_), .B(in_17bit_b[3]), .CI(
        add_1_root_r119_carry[9]), .CO(add_1_root_r119_carry[10]), .S(
        add_1_root_r119_SUM_9_) );
  ADDFX2 U147 ( .A(in_17bit_b[10]), .B(in_17bit_b[9]), .CI(
        add_2_root_r119_carry_14_), .CO(add_2_root_r119_carry_15_), .S(
        add_2_root_r119_SUM_14_) );
  ADDFX2 U148 ( .A(in_17bit_b[15]), .B(in_17bit_b[14]), .CI(
        add_3_root_r119_carry_16_), .CO(add_3_root_r119_carry_17_), .S(
        add_1_root_r119_A_16_) );
  ADDFX2 U149 ( .A(in_17bit_b[4]), .B(in_17bit_b[3]), .CI(
        add_3_root_r119_carry_5_), .CO(add_3_root_r119_carry_6_), .S(
        add_1_root_r119_A_5_) );
  ADDFX2 U150 ( .A(in_17bit_b[5]), .B(in_17bit_b[4]), .CI(
        add_3_root_r119_carry_6_), .CO(add_3_root_r119_carry_7_), .S(
        add_1_root_r119_A_6_) );
  ADDFX2 U151 ( .A(in_17bit_b[4]), .B(in_17bit_b[3]), .CI(
        add_2_root_r119_carry_8_), .CO(add_2_root_r119_carry_9_), .S(
        add_2_root_r119_SUM_8_) );
  ADDFX2 U152 ( .A(in_17bit_b[15]), .B(in_17bit_b[14]), .CI(
        add_2_root_r119_carry_19_), .CO(add_2_root_r119_carry_20_), .S(
        add_2_root_r119_SUM_19_) );
  NAND2X1 U153 ( .A(n245), .B(n244), .Y(N461) );
  AOI22X1 U154 ( .A0(N122), .A1(n247), .B0(N219), .B1(n42), .Y(n244) );
  AOI22X1 U155 ( .A0(N361), .A1(n41), .B0(n174), .B1(in_17bit_b[14]), .Y(n245)
         );
  NAND2X1 U156 ( .A(n249), .B(n248), .Y(N462) );
  AOI22X1 U157 ( .A0(N123), .A1(n247), .B0(N220), .B1(n42), .Y(n248) );
  AOI22X1 U158 ( .A0(N362), .A1(n41), .B0(n174), .B1(in_17bit_b[15]), .Y(n249)
         );
  INVX1 U159 ( .A(n44), .Y(n43) );
  INVX1 U160 ( .A(in_8bit[0]), .Y(n49) );
  INVX1 U161 ( .A(in_8bit[3]), .Y(n45) );
  INVX1 U162 ( .A(in_8bit[4]), .Y(n50) );
  NOR3X1 U163 ( .A(n175), .B(n45), .C(n49), .Y(n199) );
  CLKINVX3 U164 ( .A(n201), .Y(in_17bit_b[0]) );
  NAND3BX1 U165 ( .AN(n43), .B(n175), .C(in_8bit[3]), .Y(n196) );
  NAND3X1 U166 ( .A(n198), .B(n43), .C(n87), .Y(n88) );
  NOR2XL U167 ( .A(n46), .B(n50), .Y(n87) );
  NAND2XL U168 ( .A(N29), .B(n19), .Y(n254) );
  CLKINVX3 U169 ( .A(n246), .Y(in_17bit_b[15]) );
  BUFX3 U170 ( .A(n250), .Y(n41) );
  OAI2BB1X1 U171 ( .A0N(n25), .A1N(n35), .B0(n92), .Y(n250) );
  NAND2BX1 U172 ( .AN(n196), .B(n24), .Y(n92) );
  BUFX3 U173 ( .A(n251), .Y(n42) );
  OAI2BB1X1 U174 ( .A0N(n35), .A1N(n24), .B0(n93), .Y(n251) );
  NAND2BX1 U175 ( .AN(n196), .B(n25), .Y(n93) );
  OAI2BB1X1 U176 ( .A0N(n90), .A1N(n89), .B0(n88), .Y(n247) );
  NOR2BX1 U177 ( .AN(in_8bit[1]), .B(n94), .Y(n89) );
  NOR2BX1 U178 ( .AN(n199), .B(n86), .Y(n90) );
  OAI2BB1X1 U179 ( .A0N(n198), .A1N(n97), .B0(n96), .Y(n174) );
  INVX1 U180 ( .A(n94), .Y(n97) );
  NAND3BX1 U181 ( .AN(n95), .B(n199), .C(n43), .Y(n96) );
  AND2X2 U182 ( .A(n91), .B(n49), .Y(n25) );
  NAND2X1 U183 ( .A(n203), .B(n202), .Y(N447) );
  AOI22X1 U184 ( .A0(N108), .A1(n247), .B0(N205), .B1(n42), .Y(n202) );
  AOI22X1 U185 ( .A0(N347), .A1(n41), .B0(n174), .B1(in_17bit_b[0]), .Y(n203)
         );
  NAND2X1 U186 ( .A(n206), .B(n205), .Y(N448) );
  AOI22X1 U187 ( .A0(N109), .A1(n247), .B0(N206), .B1(n42), .Y(n205) );
  AOI22X1 U188 ( .A0(N348), .A1(n41), .B0(n174), .B1(in_17bit_b[1]), .Y(n206)
         );
  NAND2X1 U189 ( .A(n209), .B(n208), .Y(N449) );
  AOI22X1 U190 ( .A0(N110), .A1(n247), .B0(N207), .B1(n42), .Y(n208) );
  AOI22X1 U191 ( .A0(N349), .A1(n41), .B0(n174), .B1(in_17bit_b[2]), .Y(n209)
         );
  NAND2X1 U192 ( .A(n212), .B(n211), .Y(N450) );
  AOI22X1 U193 ( .A0(N111), .A1(n247), .B0(N208), .B1(n42), .Y(n211) );
  AOI22X1 U194 ( .A0(N350), .A1(n41), .B0(n174), .B1(in_17bit_b[3]), .Y(n212)
         );
  NAND2X1 U195 ( .A(n215), .B(n214), .Y(N451) );
  AOI22X1 U196 ( .A0(N112), .A1(n247), .B0(N209), .B1(n42), .Y(n214) );
  AOI22X1 U197 ( .A0(N351), .A1(n41), .B0(n174), .B1(in_17bit_b[4]), .Y(n215)
         );
  NAND2X1 U198 ( .A(n218), .B(n217), .Y(N452) );
  AOI22X1 U199 ( .A0(N113), .A1(n247), .B0(N210), .B1(n42), .Y(n217) );
  AOI22X1 U200 ( .A0(N352), .A1(n41), .B0(n174), .B1(in_17bit_b[5]), .Y(n218)
         );
  NAND2X1 U201 ( .A(n221), .B(n220), .Y(N453) );
  AOI22X1 U202 ( .A0(N114), .A1(n247), .B0(N211), .B1(n42), .Y(n220) );
  AOI22X1 U203 ( .A0(N353), .A1(n41), .B0(n174), .B1(in_17bit_b[6]), .Y(n221)
         );
  NAND2X1 U204 ( .A(n224), .B(n223), .Y(N454) );
  AOI22X1 U205 ( .A0(N115), .A1(n247), .B0(N212), .B1(n42), .Y(n223) );
  AOI22X1 U206 ( .A0(N354), .A1(n41), .B0(n174), .B1(in_17bit_b[7]), .Y(n224)
         );
  NAND2X1 U207 ( .A(n227), .B(n226), .Y(N455) );
  AOI22X1 U208 ( .A0(N116), .A1(n247), .B0(N213), .B1(n42), .Y(n226) );
  AOI22X1 U209 ( .A0(N355), .A1(n41), .B0(n174), .B1(in_17bit_b[8]), .Y(n227)
         );
  NAND2X1 U210 ( .A(n230), .B(n229), .Y(N456) );
  AOI22X1 U211 ( .A0(N117), .A1(n247), .B0(N214), .B1(n42), .Y(n229) );
  AOI22X1 U212 ( .A0(N356), .A1(n41), .B0(n174), .B1(in_17bit_b[9]), .Y(n230)
         );
  NAND2X1 U213 ( .A(n233), .B(n232), .Y(N457) );
  AOI22X1 U214 ( .A0(N118), .A1(n247), .B0(N215), .B1(n42), .Y(n232) );
  AOI22X1 U215 ( .A0(N357), .A1(n41), .B0(n174), .B1(in_17bit_b[10]), .Y(n233)
         );
  NAND2X1 U216 ( .A(n236), .B(n235), .Y(N458) );
  AOI22X1 U217 ( .A0(N119), .A1(n247), .B0(N216), .B1(n42), .Y(n235) );
  AOI22X1 U218 ( .A0(N358), .A1(n41), .B0(n174), .B1(in_17bit_b[11]), .Y(n236)
         );
  NAND2X1 U219 ( .A(n239), .B(n238), .Y(N459) );
  AOI22X1 U220 ( .A0(N120), .A1(n247), .B0(N217), .B1(n42), .Y(n238) );
  AOI22X1 U221 ( .A0(N359), .A1(n41), .B0(n174), .B1(in_17bit_b[12]), .Y(n239)
         );
  NAND2X1 U222 ( .A(n242), .B(n241), .Y(N460) );
  AOI22X1 U223 ( .A0(N121), .A1(n247), .B0(N218), .B1(n42), .Y(n241) );
  AOI22X1 U224 ( .A0(N360), .A1(n41), .B0(n174), .B1(in_17bit_b[13]), .Y(n242)
         );
  INVX1 U225 ( .A(in_8bit[5]), .Y(n44) );
  INVX1 U226 ( .A(n69), .Y(n66) );
  MXI2XL U227 ( .A(n1), .B(n17), .S0(n85), .Y(out[16]) );
  NOR4BXL U228 ( .AN(n197), .B(n49), .C(in_8bit[1]), .D(in_8bit[2]), .Y(n198)
         );
  NOR2XL U229 ( .A(in_8bit[6]), .B(in_8bit[3]), .Y(n197) );
  INVXL U230 ( .A(in_8bit[2]), .Y(n175) );
  NAND4BBX1 U231 ( .AN(n41), .BN(n42), .C(n200), .D(n253), .Y(N446) );
  AOI22XL U232 ( .A0(in_17bit[0]), .A1(n19), .B0(in_17bit[0]), .B1(n54), .Y(
        n201) );
  AOI22X1 U233 ( .A0(N22), .A1(n52), .B0(in_17bit[9]), .B1(n18), .Y(n228) );
  AOI22X1 U234 ( .A0(N23), .A1(n52), .B0(in_17bit[10]), .B1(n54), .Y(n231) );
  AOI22X1 U235 ( .A0(N27), .A1(n52), .B0(in_17bit[14]), .B1(n54), .Y(n243) );
  AOI22XL U236 ( .A0(N14), .A1(n19), .B0(in_17bit[1]), .B1(n54), .Y(n204) );
  AOI22XL U237 ( .A0(N15), .A1(n19), .B0(in_17bit[2]), .B1(n18), .Y(n207) );
  AOI22X1 U238 ( .A0(N28), .A1(n52), .B0(in_17bit[15]), .B1(n54), .Y(n246) );
  AOI22X1 U239 ( .A0(N16), .A1(n52), .B0(in_17bit[3]), .B1(n18), .Y(n210) );
  AOI22X1 U240 ( .A0(N17), .A1(n52), .B0(in_17bit[4]), .B1(n18), .Y(n213) );
  AOI22X1 U241 ( .A0(N18), .A1(n52), .B0(in_17bit[5]), .B1(n54), .Y(n216) );
  AOI22X1 U242 ( .A0(N19), .A1(n52), .B0(in_17bit[6]), .B1(n18), .Y(n219) );
  AOI22X1 U243 ( .A0(N20), .A1(n52), .B0(in_17bit[7]), .B1(n18), .Y(n222) );
  AOI22X1 U244 ( .A0(N21), .A1(n52), .B0(in_17bit[8]), .B1(n54), .Y(n225) );
  AOI22X1 U245 ( .A0(N24), .A1(n52), .B0(in_17bit[11]), .B1(n18), .Y(n234) );
  AOI22X1 U246 ( .A0(N25), .A1(n52), .B0(in_17bit[12]), .B1(n18), .Y(n237) );
  AOI22X1 U247 ( .A0(N26), .A1(n52), .B0(in_17bit[13]), .B1(n54), .Y(n240) );
  INVX1 U248 ( .A(n55), .Y(n76) );
  NAND2BX1 U249 ( .AN(n69), .B(n12), .Y(n55) );
  NAND4BXL U250 ( .AN(n47), .B(in_8bit[4]), .C(in_8bit[1]), .D(in_8bit[6]), 
        .Y(n95) );
  NAND2X1 U251 ( .A(n38), .B(n11), .Y(n69) );
  AND2X2 U252 ( .A(n76), .B(n5), .Y(n28) );
  AND2X2 U253 ( .A(n28), .B(n6), .Y(n29) );
  AND2X2 U254 ( .A(n29), .B(n7), .Y(n30) );
  AND2X2 U255 ( .A(n30), .B(n8), .Y(n31) );
  AND2X2 U256 ( .A(n31), .B(n4), .Y(n32) );
  AND2X2 U257 ( .A(n32), .B(n2), .Y(n33) );
  AND2X2 U258 ( .A(n33), .B(n3), .Y(n34) );
  NOR2XL U259 ( .A(in_8bit[6]), .B(in_8bit[4]), .Y(n195) );
  INVXL U260 ( .A(in_8bit[6]), .Y(n86) );
  AND2X2 U261 ( .A(n34), .B(n9), .Y(n36) );
  INVX1 U262 ( .A(in_17bit[0]), .Y(n98) );
  INVX1 U263 ( .A(in_17bit[1]), .Y(n99) );
  INVX1 U264 ( .A(in_17bit[2]), .Y(n100) );
  INVX1 U265 ( .A(in_17bit[3]), .Y(n101) );
  INVX1 U266 ( .A(in_17bit[4]), .Y(n158) );
  INVX1 U267 ( .A(in_17bit[5]), .Y(n160) );
  INVX1 U268 ( .A(in_17bit[6]), .Y(n161) );
  INVX1 U269 ( .A(in_17bit[7]), .Y(n162) );
  INVX1 U270 ( .A(in_17bit[8]), .Y(n163) );
  INVX1 U271 ( .A(in_17bit[9]), .Y(n164) );
  INVX1 U272 ( .A(in_17bit[10]), .Y(n167) );
  INVX1 U273 ( .A(in_17bit[11]), .Y(n168) );
  INVX1 U274 ( .A(in_17bit[12]), .Y(n170) );
  INVX1 U275 ( .A(in_17bit[13]), .Y(n171) );
  INVX1 U276 ( .A(in_17bit[14]), .Y(n172) );
  INVX1 U277 ( .A(in_17bit[15]), .Y(n173) );
  INVX1 U278 ( .A(n71), .Y(n72) );
  XNOR2X1 U279 ( .A(n16), .B(sub_add_75_b0_carry[13]), .Y(n37) );
  INVX1 U280 ( .A(n57), .Y(n58) );
  INVX1 U281 ( .A(n63), .Y(n64) );
  MX2X1 U282 ( .A(neg_mul[22]), .B(N480), .S0(n85), .Y(out[15]) );
  NOR2X1 U283 ( .A(out[0]), .B(neg_mul[8]), .Y(n38) );
  NAND2BX1 U284 ( .AN(n38), .B(neg_mul[9]), .Y(n63) );
  NAND2X1 U285 ( .A(out[0]), .B(neg_mul[8]), .Y(n57) );
  NAND2X1 U286 ( .A(neg_mul[10]), .B(n69), .Y(n71) );
  NAND2X1 U287 ( .A(sub_add_75_b0_carry[15]), .B(n13), .Y(n39) );
  AOI211X4 U288 ( .A0(n19), .A1(n68), .B0(n67), .C0(n66), .Y(out[2]) );
  XNOR2X4 U289 ( .A(n77), .B(n5), .Y(out[4]) );
  XNOR2X4 U290 ( .A(n79), .B(n6), .Y(out[5]) );
  XNOR2X4 U291 ( .A(n80), .B(n7), .Y(out[6]) );
  XNOR2X4 U292 ( .A(n82), .B(n8), .Y(out[7]) );
  XNOR2X4 U293 ( .A(n84), .B(n9), .Y(out[11]) );
  AND2X1 U294 ( .A(add_1_root_r112_carry_20_), .B(in_17bit_b[16]), .Y(
        add_1_root_r112_SUM_21_) );
  XOR2X1 U295 ( .A(in_17bit_b[16]), .B(add_1_root_r112_carry_20_), .Y(
        add_1_root_r112_SUM_20_) );
  AND2X1 U296 ( .A(add_1_root_r112_carry_19_), .B(in_17bit_b[15]), .Y(
        add_1_root_r112_carry_20_) );
  XOR2X1 U297 ( .A(in_17bit_b[15]), .B(add_1_root_r112_carry_19_), .Y(
        add_1_root_r112_SUM_19_) );
  AND2X1 U298 ( .A(add_1_root_r112_carry_18_), .B(in_17bit_b[14]), .Y(
        add_1_root_r112_carry_19_) );
  XOR2X1 U299 ( .A(in_17bit_b[14]), .B(add_1_root_r112_carry_18_), .Y(
        add_1_root_r112_SUM_18_) );
  AND2X1 U300 ( .A(add_1_root_r112_carry_17_), .B(in_17bit_b[13]), .Y(
        add_1_root_r112_carry_18_) );
  XOR2X1 U301 ( .A(in_17bit_b[13]), .B(add_1_root_r112_carry_17_), .Y(
        add_1_root_r112_SUM_17_) );
  AND2X1 U302 ( .A(add_2_root_r119_carry_21_), .B(in_17bit_b[16]), .Y(
        add_2_root_r119_SUM_22_) );
  XOR2X1 U303 ( .A(in_17bit_b[16]), .B(add_2_root_r119_carry_21_), .Y(
        add_2_root_r119_SUM_21_) );
  AND2X1 U304 ( .A(add_1_root_r119_carry[22]), .B(in_17bit_b[16]), .Y(
        add_1_root_r119_SUM_23_) );
  XOR2X1 U305 ( .A(in_17bit_b[16]), .B(add_1_root_r119_carry[22]), .Y(
        add_1_root_r119_SUM_22_) );
  AND2X1 U306 ( .A(add_1_root_r119_carry[21]), .B(in_17bit_b[15]), .Y(
        add_1_root_r119_carry[22]) );
  XOR2X1 U307 ( .A(in_17bit_b[15]), .B(add_1_root_r119_carry[21]), .Y(
        add_1_root_r119_SUM_21_) );
  AND2X1 U308 ( .A(add_1_root_r119_carry[20]), .B(in_17bit_b[14]), .Y(
        add_1_root_r119_carry[21]) );
  XOR2X1 U309 ( .A(in_17bit_b[14]), .B(add_1_root_r119_carry[20]), .Y(
        add_1_root_r119_SUM_20_) );
  AND2X1 U310 ( .A(add_1_root_r119_A_6_), .B(in_17bit_b[0]), .Y(
        add_1_root_r119_carry[7]) );
  XOR2X1 U311 ( .A(in_17bit_b[0]), .B(add_1_root_r119_A_6_), .Y(
        add_1_root_r119_SUM_6_) );
  AND2X1 U312 ( .A(add_3_root_r119_carry_18_), .B(in_17bit_b[16]), .Y(
        add_1_root_r119_A_19_) );
  XOR2X1 U313 ( .A(in_17bit_b[16]), .B(add_3_root_r119_carry_18_), .Y(
        add_1_root_r119_A_18_) );
  AND2X1 U314 ( .A(in_17bit_b[1]), .B(in_17bit_b[0]), .Y(
        add_3_root_r119_carry_3_) );
  XOR2X1 U315 ( .A(in_17bit_b[0]), .B(in_17bit_b[1]), .Y(add_1_root_r119_A_2_)
         );
  AND2X1 U316 ( .A(add_2_root_r115_carry_19_), .B(in_17bit_b[16]), .Y(
        add_2_root_r115_SUM_20_) );
  XOR2X1 U317 ( .A(in_17bit_b[16]), .B(add_2_root_r115_carry_19_), .Y(
        add_2_root_r115_SUM_19_) );
  AND2X1 U318 ( .A(add_2_root_r115_carry_18_), .B(in_17bit_b[15]), .Y(
        add_2_root_r115_carry_19_) );
  XOR2X1 U319 ( .A(in_17bit_b[15]), .B(add_2_root_r115_carry_18_), .Y(
        add_2_root_r115_SUM_18_) );
  AND2X1 U320 ( .A(add_1_root_r115_carry_22_), .B(in_17bit_b[16]), .Y(
        add_1_root_r115_SUM_23_) );
  XOR2X1 U321 ( .A(in_17bit_b[16]), .B(add_1_root_r115_carry_22_), .Y(
        add_1_root_r115_SUM_22_) );
  AND2X1 U322 ( .A(add_1_root_r115_carry_21_), .B(in_17bit_b[15]), .Y(
        add_1_root_r115_carry_22_) );
  XOR2X1 U323 ( .A(in_17bit_b[15]), .B(add_1_root_r115_carry_21_), .Y(
        add_1_root_r115_SUM_21_) );
  AND2X1 U324 ( .A(in_17bit_b[2]), .B(in_17bit_b[0]), .Y(
        add_1_root_r115_carry_7_) );
  XOR2X1 U325 ( .A(in_17bit_b[0]), .B(in_17bit_b[2]), .Y(
        add_1_root_r115_SUM_6_) );
  XOR2X1 U326 ( .A(n54), .B(sub_add_54_b0_carry[16]), .Y(N29) );
  AND2X1 U327 ( .A(sub_add_54_b0_carry[15]), .B(n173), .Y(
        sub_add_54_b0_carry[16]) );
  XOR2X1 U328 ( .A(n173), .B(sub_add_54_b0_carry[15]), .Y(N28) );
  AND2X1 U329 ( .A(sub_add_54_b0_carry[14]), .B(n172), .Y(
        sub_add_54_b0_carry[15]) );
  XOR2X1 U330 ( .A(n172), .B(sub_add_54_b0_carry[14]), .Y(N27) );
  AND2X1 U331 ( .A(sub_add_54_b0_carry[13]), .B(n171), .Y(
        sub_add_54_b0_carry[14]) );
  XOR2X1 U332 ( .A(n171), .B(sub_add_54_b0_carry[13]), .Y(N26) );
  AND2X1 U333 ( .A(sub_add_54_b0_carry[12]), .B(n170), .Y(
        sub_add_54_b0_carry[13]) );
  XOR2X1 U334 ( .A(n170), .B(sub_add_54_b0_carry[12]), .Y(N25) );
  AND2X1 U335 ( .A(sub_add_54_b0_carry[11]), .B(n168), .Y(
        sub_add_54_b0_carry[12]) );
  XOR2X1 U336 ( .A(n168), .B(sub_add_54_b0_carry[11]), .Y(N24) );
  AND2X1 U337 ( .A(sub_add_54_b0_carry[10]), .B(n167), .Y(
        sub_add_54_b0_carry[11]) );
  XOR2X1 U338 ( .A(n167), .B(sub_add_54_b0_carry[10]), .Y(N23) );
  AND2X1 U339 ( .A(sub_add_54_b0_carry[9]), .B(n164), .Y(
        sub_add_54_b0_carry[10]) );
  XOR2X1 U340 ( .A(n164), .B(sub_add_54_b0_carry[9]), .Y(N22) );
  AND2X1 U341 ( .A(sub_add_54_b0_carry[8]), .B(n163), .Y(
        sub_add_54_b0_carry[9]) );
  XOR2X1 U342 ( .A(n163), .B(sub_add_54_b0_carry[8]), .Y(N21) );
  AND2X1 U343 ( .A(sub_add_54_b0_carry[7]), .B(n162), .Y(
        sub_add_54_b0_carry[8]) );
  XOR2X1 U344 ( .A(n162), .B(sub_add_54_b0_carry[7]), .Y(N20) );
  AND2X1 U345 ( .A(sub_add_54_b0_carry[6]), .B(n161), .Y(
        sub_add_54_b0_carry[7]) );
  XOR2X1 U346 ( .A(n161), .B(sub_add_54_b0_carry[6]), .Y(N19) );
  AND2X1 U347 ( .A(sub_add_54_b0_carry[5]), .B(n160), .Y(
        sub_add_54_b0_carry[6]) );
  XOR2X1 U348 ( .A(n160), .B(sub_add_54_b0_carry[5]), .Y(N18) );
  AND2X1 U349 ( .A(sub_add_54_b0_carry[4]), .B(n158), .Y(
        sub_add_54_b0_carry[5]) );
  XOR2X1 U350 ( .A(n158), .B(sub_add_54_b0_carry[4]), .Y(N17) );
  AND2X1 U351 ( .A(sub_add_54_b0_carry[3]), .B(n101), .Y(
        sub_add_54_b0_carry[4]) );
  XOR2X1 U352 ( .A(n101), .B(sub_add_54_b0_carry[3]), .Y(N16) );
  AND2X1 U353 ( .A(sub_add_54_b0_carry[2]), .B(n100), .Y(
        sub_add_54_b0_carry[3]) );
  XOR2X1 U354 ( .A(n100), .B(sub_add_54_b0_carry[2]), .Y(N15) );
  AND2X1 U355 ( .A(n98), .B(n99), .Y(sub_add_54_b0_carry[2]) );
  XOR2X1 U356 ( .A(n99), .B(n98), .Y(N14) );
  XOR2X1 U357 ( .A(n13), .B(sub_add_75_b0_carry[15]), .Y(N480) );
  AND2X1 U358 ( .A(sub_add_75_b0_carry[14]), .B(n14), .Y(
        sub_add_75_b0_carry[15]) );
  XOR2X1 U359 ( .A(n14), .B(sub_add_75_b0_carry[14]), .Y(N479) );
  AND2X1 U360 ( .A(sub_add_75_b0_carry[13]), .B(n16), .Y(
        sub_add_75_b0_carry[14]) );
  AND2X1 U361 ( .A(n36), .B(n10), .Y(sub_add_75_b0_carry[13]) );
  AND2X1 U362 ( .A(in_17bit_b[0]), .B(in_17bit_b[4]), .Y(
        add_1_root_r112_carry_5_) );
endmodule


module butterfly_DW01_add_18 ( A, B, SUM );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  wire   n161, n162, n163, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n23, n24, n25, n26, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n44, n45, n46, n48, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160;

  INVX4 U2 ( .A(n69), .Y(n68) );
  INVX8 U3 ( .A(n92), .Y(n96) );
  NOR2X2 U4 ( .A(B[5]), .B(A[5]), .Y(n1) );
  INVX4 U5 ( .A(n105), .Y(n156) );
  BUFX2 U6 ( .A(n112), .Y(n20) );
  OAI2BB1X4 U7 ( .A0N(n42), .A1N(n58), .B0(n13), .Y(n2) );
  OAI2BB1X2 U8 ( .A0N(n42), .A1N(n58), .B0(n13), .Y(n149) );
  INVX4 U9 ( .A(n37), .Y(n114) );
  NAND2X2 U10 ( .A(B[1]), .B(A[1]), .Y(n94) );
  AND2X2 U11 ( .A(n116), .B(n113), .Y(n26) );
  BUFX8 U12 ( .A(B[11]), .Y(n23) );
  INVX1 U13 ( .A(n28), .Y(n33) );
  OAI2BB1X2 U14 ( .A0N(n111), .A1N(n130), .B0(n128), .Y(n127) );
  NAND2X1 U15 ( .A(B[0]), .B(A[0]), .Y(n97) );
  INVX1 U16 ( .A(n36), .Y(n144) );
  CLKINVX3 U17 ( .A(n9), .Y(SUM[4]) );
  INVX1 U18 ( .A(n66), .Y(n53) );
  INVX1 U19 ( .A(n11), .Y(n12) );
  AND2X2 U20 ( .A(n119), .B(n110), .Y(n3) );
  AND2X2 U21 ( .A(n124), .B(n12), .Y(n4) );
  XNOR2X4 U22 ( .A(n8), .B(n131), .Y(n5) );
  XNOR2X2 U23 ( .A(n73), .B(n74), .Y(n6) );
  XNOR2X2 U24 ( .A(n58), .B(n59), .Y(n7) );
  BUFX4 U25 ( .A(n63), .Y(n18) );
  OR2X4 U26 ( .A(A[6]), .B(B[6]), .Y(n24) );
  NAND2X4 U27 ( .A(n111), .B(n110), .Y(n122) );
  NAND2BX4 U28 ( .AN(n132), .B(n133), .Y(n8) );
  NAND3X4 U29 ( .A(n75), .B(n25), .C(n154), .Y(n153) );
  CLKINVX8 U30 ( .A(n40), .Y(n109) );
  INVX3 U31 ( .A(n135), .Y(n30) );
  XNOR2XL U32 ( .A(n81), .B(n105), .Y(n9) );
  NOR2X4 U33 ( .A(A[13]), .B(B[13]), .Y(n10) );
  INVXL U34 ( .A(n39), .Y(n11) );
  CLKBUFXL U35 ( .A(n1), .Y(n17) );
  INVXL U36 ( .A(n41), .Y(n42) );
  NAND2X1 U37 ( .A(n65), .B(n53), .Y(n54) );
  NAND2X4 U38 ( .A(n60), .B(n63), .Y(n142) );
  DLY1X1 U39 ( .A(n60), .Y(n13) );
  XOR2X4 U40 ( .A(n98), .B(n15), .Y(n14) );
  XNOR2X4 U41 ( .A(B[16]), .B(A[16]), .Y(n15) );
  NOR2BX4 U42 ( .AN(n88), .B(n160), .Y(n158) );
  OAI21X4 U43 ( .A0(n96), .A1(n97), .B0(n94), .Y(n160) );
  NAND2X4 U44 ( .A(n16), .B(n101), .Y(n100) );
  AND4X4 U45 ( .A(n111), .B(n110), .C(n109), .D(n20), .Y(n16) );
  NAND2XL U46 ( .A(n116), .B(n113), .Y(n139) );
  NAND2X4 U47 ( .A(n77), .B(n80), .Y(n154) );
  NOR2BXL U48 ( .AN(n77), .B(n1), .Y(n79) );
  NAND2X4 U49 ( .A(n39), .B(n28), .Y(n136) );
  INVX8 U50 ( .A(n121), .Y(n130) );
  INVXL U51 ( .A(n114), .Y(n19) );
  XOR2X2 U52 ( .A(n82), .B(n83), .Y(SUM[3]) );
  XOR2X1 U53 ( .A(n149), .B(n150), .Y(n162) );
  INVXL U54 ( .A(n61), .Y(n34) );
  CLKINVX4 U55 ( .A(n109), .Y(n21) );
  BUFX8 U56 ( .A(n162), .Y(SUM[10]) );
  INVX2 U57 ( .A(n107), .Y(n106) );
  NOR2BX1 U58 ( .AN(n72), .B(n71), .Y(n74) );
  XNOR2X2 U59 ( .A(n34), .B(n62), .Y(n163) );
  AOI2BB1X1 U60 ( .A0N(n108), .A1N(n156), .B0(n106), .Y(n102) );
  OAI21X4 U61 ( .A0(n102), .A1(n103), .B0(n104), .Y(n101) );
  OR2X2 U62 ( .A(B[5]), .B(A[5]), .Y(n25) );
  OAI21X4 U63 ( .A0(n70), .A1(n71), .B0(n72), .Y(n65) );
  NAND2X4 U64 ( .A(B[6]), .B(A[6]), .Y(n72) );
  NOR2X4 U65 ( .A(n10), .B(n124), .Y(n123) );
  NAND3X4 U66 ( .A(n134), .B(n61), .C(n26), .Y(n133) );
  XOR2X2 U67 ( .A(n78), .B(n79), .Y(SUM[5]) );
  INVX8 U68 ( .A(n5), .Y(SUM[13]) );
  OR2X4 U69 ( .A(A[11]), .B(B[11]), .Y(n28) );
  AOI21X4 U70 ( .A0(n23), .A1(A[11]), .B0(n36), .Y(n143) );
  INVX2 U71 ( .A(n67), .Y(n155) );
  OR2X4 U72 ( .A(A[9]), .B(B[9]), .Y(n113) );
  INVX4 U73 ( .A(n68), .Y(n29) );
  INVX8 U74 ( .A(n137), .Y(n135) );
  AND2X2 U75 ( .A(n111), .B(n128), .Y(n38) );
  NAND4BX2 U76 ( .AN(n64), .B(n113), .C(n114), .D(n115), .Y(n103) );
  INVX2 U77 ( .A(n113), .Y(n31) );
  NOR2XL U78 ( .A(B[14]), .B(A[14]), .Y(n32) );
  AND3X4 U79 ( .A(n112), .B(n114), .C(n115), .Y(n134) );
  NAND2BX4 U80 ( .AN(n132), .B(n133), .Y(n35) );
  AND2X4 U81 ( .A(A[10]), .B(B[10]), .Y(n36) );
  NAND2X2 U82 ( .A(B[15]), .B(A[15]), .Y(n119) );
  NAND2X1 U83 ( .A(B[14]), .B(A[14]), .Y(n128) );
  NAND2BX4 U84 ( .AN(n33), .B(n30), .Y(n104) );
  AND2X2 U85 ( .A(A[14]), .B(B[14]), .Y(n44) );
  NOR2BX1 U86 ( .AN(n60), .B(n31), .Y(n59) );
  NOR2BXL U87 ( .AN(n144), .B(n19), .Y(n150) );
  NAND2X4 U88 ( .A(B[13]), .B(A[13]), .Y(n121) );
  INVX4 U89 ( .A(n116), .Y(n64) );
  OAI21X4 U90 ( .A0(n135), .A1(n136), .B0(n124), .Y(n132) );
  NOR2X4 U91 ( .A(B[10]), .B(A[10]), .Y(n37) );
  XNOR2X4 U92 ( .A(n129), .B(n38), .Y(SUM[14]) );
  NAND2X4 U93 ( .A(n2), .B(n114), .Y(n148) );
  OR2X4 U94 ( .A(A[12]), .B(B[12]), .Y(n39) );
  OR2X4 U95 ( .A(n125), .B(n3), .Y(n45) );
  NOR2X4 U96 ( .A(n41), .B(n37), .Y(n141) );
  NOR2X4 U97 ( .A(A[13]), .B(B[13]), .Y(n40) );
  AND2X2 U98 ( .A(n121), .B(n109), .Y(n131) );
  NAND2X4 U99 ( .A(A[9]), .B(B[9]), .Y(n60) );
  BUFX20 U100 ( .A(n161), .Y(SUM[11]) );
  NAND2X4 U101 ( .A(B[7]), .B(A[7]), .Y(n67) );
  NOR2BX4 U102 ( .AN(n72), .B(n155), .Y(n152) );
  NOR2X4 U103 ( .A(B[9]), .B(A[9]), .Y(n41) );
  NAND2X4 U104 ( .A(A[5]), .B(B[5]), .Y(n77) );
  NOR2X4 U105 ( .A(n123), .B(n44), .Y(n120) );
  INVX4 U106 ( .A(n78), .Y(n76) );
  OAI21X4 U107 ( .A0(n57), .A1(n156), .B0(n80), .Y(n78) );
  NAND3XL U108 ( .A(n115), .B(n61), .C(n114), .Y(n140) );
  NAND2X4 U109 ( .A(n116), .B(n61), .Y(n151) );
  OR2X4 U110 ( .A(B[7]), .B(A[7]), .Y(n69) );
  NAND2X4 U111 ( .A(n148), .B(n144), .Y(n145) );
  NOR2X2 U112 ( .A(n32), .B(n21), .Y(n126) );
  NAND2X2 U113 ( .A(n125), .B(n3), .Y(n46) );
  XOR2X4 U114 ( .A(n138), .B(n4), .Y(SUM[12]) );
  AOI21X4 U115 ( .A0(n120), .A1(n121), .B0(n122), .Y(n117) );
  NOR2X4 U116 ( .A(A[4]), .B(B[4]), .Y(n57) );
  OR2X4 U117 ( .A(A[2]), .B(B[2]), .Y(n91) );
  NOR2BXL U118 ( .AN(n80), .B(n57), .Y(n81) );
  NAND4BBX4 U119 ( .AN(n1), .BN(n57), .C(n69), .D(n24), .Y(n108) );
  NAND2X4 U120 ( .A(n45), .B(n46), .Y(SUM[15]) );
  INVX8 U121 ( .A(n14), .Y(SUM[16]) );
  CLKINVX4 U122 ( .A(n163), .Y(n48) );
  INVX8 U123 ( .A(n48), .Y(SUM[8]) );
  INVX8 U124 ( .A(n6), .Y(SUM[6]) );
  INVX8 U125 ( .A(n7), .Y(SUM[9]) );
  NAND2X4 U126 ( .A(n151), .B(n18), .Y(n58) );
  NAND2X4 U127 ( .A(B[4]), .B(A[4]), .Y(n80) );
  NOR2BX1 U128 ( .AN(n67), .B(n68), .Y(n66) );
  NAND2X2 U129 ( .A(n52), .B(n66), .Y(n55) );
  NAND2X4 U130 ( .A(B[2]), .B(A[2]), .Y(n88) );
  NAND2X2 U131 ( .A(B[12]), .B(A[12]), .Y(n124) );
  NAND2X4 U132 ( .A(n54), .B(n55), .Y(SUM[7]) );
  INVX2 U133 ( .A(n65), .Y(n52) );
  INVX2 U134 ( .A(n73), .Y(n70) );
  NOR2BXL U135 ( .AN(n88), .B(n87), .Y(n90) );
  OAI21X2 U136 ( .A0(n139), .A1(n140), .B0(n104), .Y(n138) );
  NAND2X1 U137 ( .A(B[3]), .B(A[3]), .Y(n84) );
  OR2X4 U138 ( .A(A[8]), .B(B[8]), .Y(n116) );
  NOR2BX1 U139 ( .AN(n97), .B(n56), .Y(SUM[0]) );
  NOR2XL U140 ( .A(A[0]), .B(B[0]), .Y(n56) );
  XOR2X1 U141 ( .A(n89), .B(n90), .Y(SUM[2]) );
  INVX1 U142 ( .A(n91), .Y(n87) );
  NOR2BX1 U143 ( .AN(n18), .B(n64), .Y(n62) );
  INVX1 U144 ( .A(n119), .Y(n118) );
  OAI21XL U145 ( .A0(n86), .A1(n87), .B0(n88), .Y(n82) );
  NOR2BX1 U146 ( .AN(n84), .B(n85), .Y(n83) );
  INVX1 U147 ( .A(n89), .Y(n86) );
  XOR2X1 U148 ( .A(n93), .B(n95), .Y(SUM[1]) );
  NOR2BXL U149 ( .AN(n94), .B(n96), .Y(n95) );
  INVXL U150 ( .A(n75), .Y(n71) );
  OAI2BB1X1 U151 ( .A0N(n92), .A1N(n93), .B0(n94), .Y(n89) );
  INVXL U152 ( .A(n157), .Y(n85) );
  INVX1 U153 ( .A(n97), .Y(n93) );
  NAND2X4 U154 ( .A(n99), .B(n100), .Y(n98) );
  OAI2BB1X4 U155 ( .A0N(n152), .A1N(n153), .B0(n29), .Y(n107) );
  NAND2XL U156 ( .A(n28), .B(n147), .Y(n146) );
  NAND2XL U157 ( .A(A[11]), .B(n23), .Y(n147) );
  OAI21X4 U158 ( .A0(n76), .A1(n17), .B0(n77), .Y(n73) );
  NOR2X4 U159 ( .A(n117), .B(n118), .Y(n99) );
  AOI21X4 U160 ( .A0(n8), .A1(n126), .B0(n127), .Y(n125) );
  OR2X4 U161 ( .A(B[15]), .B(A[15]), .Y(n110) );
  AOI21X4 U162 ( .A0(n35), .A1(n109), .B0(n130), .Y(n129) );
  OR2X4 U163 ( .A(B[14]), .B(A[14]), .Y(n111) );
  OR2X4 U164 ( .A(A[12]), .B(B[12]), .Y(n112) );
  OAI2BB1X4 U165 ( .A0N(n141), .A1N(n142), .B0(n143), .Y(n137) );
  XNOR2X4 U166 ( .A(n145), .B(n146), .Y(n161) );
  OR2X4 U167 ( .A(A[11]), .B(B[11]), .Y(n115) );
  NAND2X4 U168 ( .A(A[8]), .B(B[8]), .Y(n63) );
  OAI21X4 U169 ( .A0(n108), .A1(n156), .B0(n107), .Y(n61) );
  OR2X4 U170 ( .A(B[6]), .B(A[6]), .Y(n75) );
  OAI21X4 U171 ( .A0(n158), .A1(n159), .B0(n84), .Y(n105) );
  NAND2X4 U172 ( .A(n91), .B(n157), .Y(n159) );
  OR2X4 U173 ( .A(A[3]), .B(B[3]), .Y(n157) );
  OR2X4 U174 ( .A(A[1]), .B(B[1]), .Y(n92) );
endmodule


module butterfly_DW01_add_49 ( A, B, SUM );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184;

  NAND4X2 U2 ( .A(n163), .B(n21), .C(n70), .D(n164), .Y(n182) );
  NAND2X1 U3 ( .A(A[5]), .B(B[5]), .Y(n6) );
  BUFX8 U4 ( .A(n35), .Y(n29) );
  OR2X4 U5 ( .A(B[6]), .B(A[6]), .Y(n1) );
  AND2X2 U6 ( .A(n121), .B(n149), .Y(n2) );
  OAI2BB1X2 U7 ( .A0N(n154), .A1N(n148), .B0(n149), .Y(n124) );
  OR2X2 U8 ( .A(n61), .B(n62), .Y(n51) );
  NAND2X4 U9 ( .A(n26), .B(n77), .Y(n86) );
  CLKINVX3 U10 ( .A(n139), .Y(n41) );
  AND2X2 U11 ( .A(n56), .B(n59), .Y(n47) );
  CLKINVX3 U12 ( .A(A[2]), .Y(n179) );
  NAND3X2 U13 ( .A(n5), .B(n170), .C(n172), .Y(n169) );
  CLKINVX3 U14 ( .A(A[11]), .Y(n7) );
  NOR2X2 U15 ( .A(n117), .B(n29), .Y(n140) );
  INVX4 U16 ( .A(n96), .Y(n100) );
  AND2X2 U17 ( .A(n73), .B(n82), .Y(n84) );
  INVX1 U18 ( .A(n31), .Y(n67) );
  AND2X2 U19 ( .A(B[4]), .B(A[4]), .Y(n184) );
  CLKINVX3 U20 ( .A(n149), .Y(n139) );
  OR2X1 U21 ( .A(A[2]), .B(B[2]), .Y(n95) );
  NAND2X2 U22 ( .A(B[7]), .B(A[7]), .Y(n163) );
  BUFX8 U23 ( .A(n86), .Y(n24) );
  INVX1 U24 ( .A(n81), .Y(n85) );
  INVX1 U25 ( .A(n73), .Y(n72) );
  INVX1 U26 ( .A(A[7]), .Y(n15) );
  INVX4 U27 ( .A(n86), .Y(n57) );
  NOR2BX2 U28 ( .AN(n32), .B(n140), .Y(n136) );
  NOR2X1 U29 ( .A(n122), .B(n123), .Y(n104) );
  INVX1 U30 ( .A(n107), .Y(n106) );
  OAI21XL U31 ( .A0(n108), .A1(n109), .B0(n110), .Y(n107) );
  NOR2X1 U32 ( .A(n113), .B(n114), .Y(n108) );
  NOR2BX2 U33 ( .AN(n98), .B(n100), .Y(n99) );
  AND2X1 U34 ( .A(n117), .B(n121), .Y(n3) );
  AND2X2 U35 ( .A(n110), .B(n112), .Y(n4) );
  AND2X4 U36 ( .A(n47), .B(n171), .Y(n5) );
  INVX1 U37 ( .A(n158), .Y(n156) );
  BUFX8 U38 ( .A(n116), .Y(n32) );
  NAND2BX4 U39 ( .AN(n6), .B(n42), .Y(n164) );
  AND2X4 U40 ( .A(n95), .B(n181), .Y(n52) );
  INVX1 U41 ( .A(n36), .Y(n153) );
  NAND4BX4 U42 ( .AN(n28), .B(n19), .C(n24), .D(n45), .Y(n177) );
  NOR2X2 U43 ( .A(A[13]), .B(B[13]), .Y(n35) );
  NAND2X4 U44 ( .A(n7), .B(n8), .Y(n9) );
  NAND2X4 U45 ( .A(n9), .B(n158), .Y(n160) );
  INVX4 U46 ( .A(B[11]), .Y(n8) );
  CLKINVX2 U47 ( .A(n42), .Y(n69) );
  BUFX8 U48 ( .A(n61), .Y(n28) );
  AND2X4 U49 ( .A(n165), .B(n60), .Y(n11) );
  INVX2 U50 ( .A(n151), .Y(n150) );
  AND2X2 U51 ( .A(n121), .B(n132), .Y(n10) );
  OR2X4 U52 ( .A(A[7]), .B(B[7]), .Y(n165) );
  NAND2X4 U53 ( .A(n60), .B(n165), .Y(n126) );
  INVX4 U54 ( .A(n34), .Y(n117) );
  AND2X4 U55 ( .A(B[12]), .B(A[12]), .Y(n34) );
  INVXL U56 ( .A(n11), .Y(n40) );
  AND2X2 U57 ( .A(n56), .B(n19), .Y(n55) );
  CLKINVX4 U58 ( .A(n161), .Y(n174) );
  NAND3X4 U59 ( .A(n39), .B(n10), .C(n41), .Y(n137) );
  NAND2X4 U60 ( .A(n147), .B(n23), .Y(n12) );
  NAND2X2 U61 ( .A(n148), .B(n13), .Y(n22) );
  INVX4 U62 ( .A(n12), .Y(n13) );
  INVX3 U63 ( .A(n121), .Y(n37) );
  AND4X2 U64 ( .A(n21), .B(n70), .C(n164), .D(n163), .Y(n18) );
  OAI21X4 U65 ( .A0(n57), .A1(n85), .B0(n79), .Y(n83) );
  XOR2X4 U66 ( .A(n175), .B(n14), .Y(SUM[10]) );
  AND2X1 U67 ( .A(n146), .B(n158), .Y(n14) );
  NAND3BX4 U68 ( .AN(n28), .B(n45), .C(n24), .Y(n172) );
  NAND2X2 U69 ( .A(B[1]), .B(A[1]), .Y(n98) );
  NAND2BX4 U70 ( .AN(n163), .B(n45), .Y(n171) );
  INVX8 U71 ( .A(n62), .Y(n45) );
  XOR2X2 U72 ( .A(n93), .B(n94), .Y(SUM[2]) );
  NOR2BX1 U73 ( .AN(n15), .B(B[7]), .Y(n16) );
  NAND4BX4 U74 ( .AN(n16), .B(n76), .C(n82), .D(n81), .Y(n61) );
  NAND4X2 U75 ( .A(n177), .B(n176), .C(n17), .D(n56), .Y(n175) );
  OR2X2 U76 ( .A(n174), .B(n59), .Y(n17) );
  NAND3X1 U77 ( .A(n164), .B(n70), .C(n162), .Y(n173) );
  AOI21X4 U78 ( .A0(n133), .A1(n20), .B0(n134), .Y(n129) );
  NAND3X4 U79 ( .A(n82), .B(n76), .C(n184), .Y(n162) );
  NAND3X2 U80 ( .A(n82), .B(n1), .C(n184), .Y(n21) );
  INVX4 U81 ( .A(n174), .Y(n19) );
  BUFX8 U82 ( .A(n111), .Y(n20) );
  NOR2X1 U83 ( .A(n29), .B(n117), .Y(n113) );
  NAND2X4 U84 ( .A(n158), .B(n44), .Y(n148) );
  NOR2X2 U85 ( .A(A[9]), .B(B[9]), .Y(n157) );
  NOR2BX2 U86 ( .AN(n161), .B(n58), .Y(n183) );
  BUFX8 U87 ( .A(n146), .Y(n23) );
  OAI2BB1X4 U88 ( .A0N(n50), .A1N(n71), .B0(n73), .Y(n74) );
  NAND2X4 U89 ( .A(B[0]), .B(A[0]), .Y(n101) );
  NAND3BX2 U90 ( .AN(n120), .B(n39), .C(n2), .Y(n130) );
  INVX4 U91 ( .A(n30), .Y(n70) );
  NAND4X4 U92 ( .A(n162), .B(n70), .C(n164), .D(n163), .Y(n60) );
  AND2X4 U93 ( .A(n126), .B(n151), .Y(n25) );
  OAI2BB1X4 U94 ( .A0N(B[9]), .A1N(A[9]), .B0(n59), .Y(n155) );
  CLKBUFX8 U95 ( .A(n80), .Y(n26) );
  NAND2XL U96 ( .A(B[3]), .B(A[3]), .Y(n80) );
  INVX4 U97 ( .A(n25), .Y(n27) );
  INVXL U98 ( .A(n28), .Y(n127) );
  AND2X2 U99 ( .A(B[6]), .B(A[6]), .Y(n30) );
  NAND3X4 U100 ( .A(n148), .B(n147), .C(n23), .Y(n39) );
  OAI2BB1X1 U101 ( .A0N(B[7]), .A1N(A[7]), .B0(n165), .Y(n31) );
  NAND2XL U102 ( .A(B[13]), .B(A[13]), .Y(n116) );
  NAND2X4 U103 ( .A(B[11]), .B(A[11]), .Y(n147) );
  NAND2BX4 U104 ( .AN(n160), .B(n53), .Y(n33) );
  OAI2BB1X2 U105 ( .A0N(n153), .A1N(n63), .B0(n124), .Y(n152) );
  NOR2BX1 U106 ( .AN(n146), .B(n159), .Y(n154) );
  NOR2XL U107 ( .A(n174), .B(n156), .Y(n168) );
  NAND2BX4 U108 ( .AN(n160), .B(n53), .Y(n36) );
  AND2X4 U109 ( .A(n161), .B(n65), .Y(n53) );
  XNOR2X4 U110 ( .A(n57), .B(n87), .Y(SUM[4]) );
  CLKINVX8 U111 ( .A(n37), .Y(n38) );
  NAND4BX4 U112 ( .AN(n33), .B(n63), .C(n38), .D(n132), .Y(n138) );
  AND2X4 U113 ( .A(n81), .B(n82), .Y(n50) );
  NAND2X2 U114 ( .A(B[10]), .B(A[10]), .Y(n146) );
  OR2X4 U115 ( .A(B[6]), .B(A[6]), .Y(n42) );
  OR2X2 U116 ( .A(A[3]), .B(B[3]), .Y(n181) );
  NAND2X2 U117 ( .A(B[5]), .B(A[5]), .Y(n73) );
  XOR2X4 U118 ( .A(n27), .B(n64), .Y(SUM[8]) );
  AOI21X1 U119 ( .A0(n125), .A1(n40), .B0(n33), .Y(n122) );
  NAND2X2 U120 ( .A(B[9]), .B(A[9]), .Y(n56) );
  NAND2BX4 U121 ( .AN(n61), .B(n24), .Y(n151) );
  NAND3X4 U122 ( .A(n131), .B(n129), .C(n130), .Y(n128) );
  INVX4 U123 ( .A(n155), .Y(n43) );
  NOR2X4 U124 ( .A(n157), .B(n43), .Y(n44) );
  OR2X4 U125 ( .A(A[1]), .B(B[1]), .Y(n96) );
  INVX8 U126 ( .A(n65), .Y(n62) );
  NAND2X4 U127 ( .A(B[8]), .B(A[8]), .Y(n59) );
  NAND2X2 U128 ( .A(n77), .B(n78), .Y(n71) );
  XOR2X1 U129 ( .A(B[16]), .B(A[16]), .Y(n103) );
  AND2X1 U130 ( .A(n26), .B(n181), .Y(n89) );
  OAI21X2 U131 ( .A0(n68), .A1(n69), .B0(n70), .Y(n66) );
  NAND2X2 U132 ( .A(n173), .B(n49), .Y(n170) );
  NAND2X2 U133 ( .A(B[14]), .B(A[14]), .Y(n115) );
  NAND2X4 U134 ( .A(B[4]), .B(A[4]), .Y(n79) );
  NAND2X2 U135 ( .A(B[15]), .B(A[15]), .Y(n110) );
  OR2X4 U136 ( .A(B[5]), .B(A[5]), .Y(n82) );
  AOI21X2 U137 ( .A0(B[11]), .A1(A[11]), .B0(n139), .Y(n167) );
  NOR2X4 U138 ( .A(n11), .B(n150), .Y(n143) );
  AND2X2 U139 ( .A(n79), .B(n26), .Y(n78) );
  NAND4BBX2 U140 ( .AN(n120), .BN(n33), .C(n63), .D(n38), .Y(n131) );
  OAI21X2 U141 ( .A0(n29), .A1(n117), .B0(n32), .Y(n133) );
  NOR2BX2 U142 ( .AN(n79), .B(n85), .Y(n87) );
  OR2X4 U143 ( .A(A[11]), .B(B[11]), .Y(n149) );
  NAND2X2 U144 ( .A(n65), .B(n165), .Y(n58) );
  OR2X4 U145 ( .A(A[4]), .B(B[4]), .Y(n81) );
  XOR2X4 U146 ( .A(n83), .B(n84), .Y(SUM[5]) );
  OR2X4 U147 ( .A(A[14]), .B(B[14]), .Y(n111) );
  NAND2X4 U148 ( .A(n132), .B(n111), .Y(n120) );
  OR2X4 U149 ( .A(B[10]), .B(A[10]), .Y(n158) );
  NAND2BX4 U150 ( .AN(n36), .B(n38), .Y(n144) );
  CLKINVX3 U151 ( .A(n147), .Y(n159) );
  OAI21X1 U152 ( .A0(n90), .A1(n91), .B0(n92), .Y(n88) );
  NAND2XL U153 ( .A(n115), .B(n32), .Y(n114) );
  AOI21X2 U154 ( .A0(n50), .A1(n71), .B0(n72), .Y(n68) );
  OAI21X4 U155 ( .A0(n104), .A1(n105), .B0(n106), .Y(n102) );
  NAND2X2 U156 ( .A(n118), .B(n119), .Y(n105) );
  OAI2BB1X1 U157 ( .A0N(n26), .A1N(n77), .B0(n127), .Y(n125) );
  AND2X2 U158 ( .A(n115), .B(n111), .Y(n46) );
  XOR2X2 U159 ( .A(n97), .B(n99), .Y(SUM[1]) );
  NOR2BX2 U160 ( .AN(n92), .B(n91), .Y(n94) );
  NAND2X2 U161 ( .A(n182), .B(n183), .Y(n176) );
  OAI2BB1X4 U162 ( .A0N(n96), .A1N(n97), .B0(n98), .Y(n93) );
  AND2X1 U163 ( .A(n112), .B(n38), .Y(n118) );
  NOR2BX1 U164 ( .AN(n101), .B(n48), .Y(SUM[0]) );
  NOR2XL U165 ( .A(A[0]), .B(B[0]), .Y(n48) );
  INVX1 U166 ( .A(n93), .Y(n90) );
  INVX1 U167 ( .A(n120), .Y(n119) );
  NOR2BX2 U168 ( .AN(n32), .B(n29), .Y(n142) );
  NOR2BX1 U169 ( .AN(n59), .B(n62), .Y(n64) );
  INVX1 U170 ( .A(n95), .Y(n91) );
  INVX1 U171 ( .A(n115), .Y(n134) );
  AND2X1 U172 ( .A(n65), .B(n165), .Y(n49) );
  INVXL U173 ( .A(B[2]), .Y(n180) );
  INVX1 U174 ( .A(n101), .Y(n97) );
  INVX1 U175 ( .A(n124), .Y(n123) );
  NAND2X4 U176 ( .A(n52), .B(n178), .Y(n77) );
  NAND2XL U177 ( .A(B[2]), .B(A[2]), .Y(n92) );
  NAND2XL U178 ( .A(n20), .B(n112), .Y(n109) );
  AOI21X4 U179 ( .A0(n22), .A1(n2), .B0(n34), .Y(n145) );
  XOR2X4 U180 ( .A(n54), .B(n55), .Y(SUM[9]) );
  OAI221X2 U181 ( .A0(n57), .A1(n51), .B0(n18), .B1(n58), .C0(n59), .Y(n54) );
  XOR2X4 U182 ( .A(n66), .B(n67), .Y(SUM[7]) );
  XOR2X4 U183 ( .A(n74), .B(n75), .Y(SUM[6]) );
  NOR2BX4 U184 ( .AN(n70), .B(n69), .Y(n75) );
  XOR2X4 U185 ( .A(n88), .B(n89), .Y(SUM[3]) );
  XOR2X4 U186 ( .A(n102), .B(n103), .Y(SUM[16]) );
  XOR2X4 U187 ( .A(n128), .B(n4), .Y(SUM[15]) );
  OR2X4 U188 ( .A(A[15]), .B(B[15]), .Y(n112) );
  XOR2X4 U189 ( .A(n135), .B(n46), .Y(SUM[14]) );
  NAND3X4 U190 ( .A(n138), .B(n137), .C(n136), .Y(n135) );
  XOR2X4 U191 ( .A(n141), .B(n142), .Y(SUM[13]) );
  OR2X4 U192 ( .A(A[13]), .B(B[13]), .Y(n132) );
  OAI21X4 U193 ( .A0(n143), .A1(n144), .B0(n145), .Y(n141) );
  XOR2X4 U194 ( .A(n152), .B(n3), .Y(SUM[12]) );
  OR2X4 U195 ( .A(A[12]), .B(B[12]), .Y(n121) );
  NAND2X4 U196 ( .A(n151), .B(n126), .Y(n63) );
  XOR2X4 U197 ( .A(n166), .B(n167), .Y(SUM[11]) );
  OAI2BB1X4 U198 ( .A0N(n168), .A1N(n169), .B0(n23), .Y(n166) );
  OAI221X2 U199 ( .A0(n100), .A1(n101), .B0(n179), .B1(n180), .C0(n98), .Y(
        n178) );
  OR2X4 U200 ( .A(A[8]), .B(B[8]), .Y(n65) );
  OR2X4 U201 ( .A(B[6]), .B(A[6]), .Y(n76) );
  OR2X4 U202 ( .A(B[9]), .B(A[9]), .Y(n161) );
endmodule


module butterfly_DW01_add_50 ( A, B, SUM );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  wire   n193, n194, n195, n196, n197, n198, n199, n2, n3, n4, n5, n6, n8, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n38, n39,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n62, n63, n64, n66, n67, n68, n69, n70, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192;

  AND2X4 U2 ( .A(n49), .B(n148), .Y(n120) );
  BUFX20 U3 ( .A(n66), .Y(SUM[15]) );
  NOR2BX4 U4 ( .AN(n164), .B(n166), .Y(n165) );
  CLKINVXL U5 ( .A(n178), .Y(n25) );
  NAND3X2 U6 ( .A(n136), .B(n52), .C(n46), .Y(n135) );
  CLKINVX3 U7 ( .A(n76), .Y(n187) );
  NAND2X4 U8 ( .A(n144), .B(n142), .Y(n174) );
  NAND2X1 U9 ( .A(B[12]), .B(A[12]), .Y(n164) );
  NAND3X2 U10 ( .A(A[12]), .B(B[12]), .C(n128), .Y(n162) );
  NOR2BX1 U11 ( .AN(n114), .B(n116), .Y(n115) );
  INVX4 U12 ( .A(n112), .Y(n116) );
  NAND2X1 U13 ( .A(n31), .B(n144), .Y(n182) );
  OR2X2 U14 ( .A(A[8]), .B(B[8]), .Y(n80) );
  BUFX12 U15 ( .A(A[8]), .Y(n6) );
  BUFX12 U16 ( .A(n198), .Y(SUM[5]) );
  XOR2X1 U17 ( .A(n94), .B(n95), .Y(n198) );
  INVX4 U18 ( .A(n30), .Y(n31) );
  INVX1 U19 ( .A(n36), .Y(n166) );
  INVX2 U20 ( .A(n142), .Y(n30) );
  INVX1 U21 ( .A(n47), .Y(n48) );
  OR2X2 U22 ( .A(A[1]), .B(B[1]), .Y(n112) );
  INVX1 U23 ( .A(n149), .Y(n159) );
  BUFX4 U24 ( .A(n28), .Y(n73) );
  CLKINVX3 U25 ( .A(n26), .Y(n27) );
  INVX2 U26 ( .A(n89), .Y(n86) );
  BUFX3 U27 ( .A(n199), .Y(SUM[0]) );
  BUFX16 U28 ( .A(n194), .Y(SUM[12]) );
  CLKINVX3 U29 ( .A(n20), .Y(SUM[2]) );
  XOR2X2 U30 ( .A(n102), .B(n103), .Y(SUM[3]) );
  CLKINVX3 U31 ( .A(n16), .Y(SUM[4]) );
  NOR2BX1 U32 ( .AN(n98), .B(n96), .Y(n100) );
  NOR2BX1 U33 ( .AN(n93), .B(n92), .Y(n95) );
  NAND2X2 U34 ( .A(n161), .B(n154), .Y(n153) );
  AND2X4 U35 ( .A(n101), .B(n190), .Y(n2) );
  NAND2X1 U36 ( .A(n163), .B(n29), .Y(n3) );
  AND2X1 U37 ( .A(n140), .B(n25), .Y(n4) );
  INVX1 U38 ( .A(n18), .Y(n56) );
  INVX4 U39 ( .A(n83), .Y(n169) );
  CLKBUFX2 U40 ( .A(A[11]), .Y(n34) );
  NAND3X4 U41 ( .A(n52), .B(n136), .C(n46), .Y(n170) );
  INVX2 U42 ( .A(n52), .Y(n53) );
  INVX2 U43 ( .A(B[10]), .Y(n47) );
  NAND3X4 U44 ( .A(n5), .B(n129), .C(n130), .Y(n122) );
  AND2X4 U45 ( .A(n8), .B(n140), .Y(n5) );
  NAND2X4 U46 ( .A(n39), .B(n160), .Y(n58) );
  CLKINVX2 U47 ( .A(n39), .Y(n22) );
  CLKBUFX4 U48 ( .A(A[13]), .Y(n13) );
  NAND2X2 U49 ( .A(n175), .B(n176), .Y(n8) );
  NAND4X4 U50 ( .A(n52), .B(n2), .C(n99), .D(n46), .Y(n15) );
  BUFX8 U51 ( .A(B[8]), .Y(n42) );
  NOR3X4 U52 ( .A(n143), .B(n30), .C(n73), .Y(n133) );
  NAND3BX4 U53 ( .AN(n187), .B(n177), .C(n185), .Y(n184) );
  NAND3X4 U54 ( .A(n150), .B(n163), .C(n149), .Y(n147) );
  NAND3X2 U55 ( .A(n128), .B(B[12]), .C(A[12]), .Y(n150) );
  NAND2BX1 U56 ( .AN(n47), .B(n41), .Y(n183) );
  BUFX2 U57 ( .A(B[7]), .Y(n54) );
  CLKBUFX2 U58 ( .A(A[7]), .Y(n72) );
  INVX4 U59 ( .A(n75), .Y(n12) );
  NAND3BX4 U60 ( .AN(n87), .B(n46), .C(n136), .Y(n35) );
  NAND3BX4 U61 ( .AN(n169), .B(n135), .C(n134), .Y(n79) );
  BUFX12 U62 ( .A(n196), .Y(SUM[10]) );
  INVX8 U63 ( .A(n99), .Y(n97) );
  NAND4X4 U64 ( .A(n2), .B(n52), .C(n99), .D(n46), .Y(n171) );
  CLKINVX4 U65 ( .A(A[6]), .Y(n32) );
  CLKINVX8 U66 ( .A(n15), .Y(n78) );
  NOR2BX1 U67 ( .AN(n83), .B(n84), .Y(n82) );
  OAI21X2 U68 ( .A0(n6), .A1(n42), .B0(n131), .Y(n143) );
  BUFX20 U69 ( .A(n193), .Y(SUM[14]) );
  XOR2X4 U70 ( .A(n119), .B(n11), .Y(n10) );
  XOR2X4 U71 ( .A(B[16]), .B(n118), .Y(n11) );
  XOR2X4 U72 ( .A(n23), .B(n165), .Y(n194) );
  XNOR2X4 U73 ( .A(n74), .B(n12), .Y(SUM[9]) );
  NAND2BX4 U74 ( .AN(n14), .B(n29), .Y(n155) );
  NOR2X4 U75 ( .A(A[12]), .B(B[12]), .Y(n14) );
  INVX2 U76 ( .A(n155), .Y(n160) );
  CLKINVX8 U77 ( .A(n32), .Y(n33) );
  AND3X4 U78 ( .A(n35), .B(n83), .C(n172), .Y(n38) );
  NAND2X4 U79 ( .A(n148), .B(n19), .Y(n151) );
  XOR2X1 U80 ( .A(n97), .B(n100), .Y(n16) );
  NAND4X4 U81 ( .A(n171), .B(n170), .C(n83), .D(n172), .Y(n168) );
  DLY1X1 U82 ( .A(B[6]), .Y(n17) );
  OR2X4 U83 ( .A(A[8]), .B(B[8]), .Y(n18) );
  OR2X4 U84 ( .A(B[15]), .B(A[15]), .Y(n19) );
  AND2X4 U85 ( .A(n33), .B(B[6]), .Y(n69) );
  BUFX2 U86 ( .A(A[10]), .Y(n41) );
  XNOR2X4 U87 ( .A(n62), .B(n3), .Y(SUM[13]) );
  NAND2X4 U88 ( .A(n42), .B(n6), .Y(n24) );
  XOR2X1 U89 ( .A(n107), .B(n111), .Y(n20) );
  INVX2 U90 ( .A(n110), .Y(n107) );
  AND2X4 U91 ( .A(n69), .B(n85), .Y(n21) );
  BUFX20 U92 ( .A(n85), .Y(n46) );
  NAND2XL U93 ( .A(B[6]), .B(n33), .Y(n88) );
  NAND2X2 U94 ( .A(n42), .B(n6), .Y(n177) );
  AOI21X4 U95 ( .A0(n158), .A1(n127), .B0(n159), .Y(n152) );
  CLKINVX3 U96 ( .A(n22), .Y(n23) );
  CLKINVX2 U97 ( .A(B[11]), .Y(n26) );
  NAND2X4 U98 ( .A(n27), .B(n34), .Y(n140) );
  AND2X2 U99 ( .A(n149), .B(n127), .Y(n51) );
  NOR2X2 U100 ( .A(B[9]), .B(A[9]), .Y(n28) );
  NAND2X4 U101 ( .A(n44), .B(n13), .Y(n163) );
  OR2X4 U102 ( .A(B[13]), .B(A[13]), .Y(n29) );
  OR2X4 U103 ( .A(A[12]), .B(B[12]), .Y(n36) );
  BUFX12 U104 ( .A(n197), .Y(SUM[7]) );
  NAND3BX4 U105 ( .AN(n156), .B(n141), .C(n157), .Y(n39) );
  NAND3X1 U106 ( .A(n33), .B(n17), .C(n46), .Y(n134) );
  INVX8 U107 ( .A(n63), .Y(SUM[8]) );
  XOR2X2 U108 ( .A(n64), .B(n77), .Y(n63) );
  INVX8 U109 ( .A(n10), .Y(SUM[16]) );
  AND2X1 U110 ( .A(n18), .B(n177), .Y(n64) );
  NOR2BX4 U111 ( .AN(n45), .B(n155), .Y(n154) );
  OAI2BB1X4 U112 ( .A0N(n35), .A1N(n189), .B0(n18), .Y(n188) );
  NAND2X2 U113 ( .A(B[15]), .B(A[15]), .Y(n148) );
  INVX8 U114 ( .A(n87), .Y(n52) );
  NOR2X4 U115 ( .A(n21), .B(n169), .Y(n189) );
  INVX2 U116 ( .A(B[13]), .Y(n43) );
  CLKINVX4 U117 ( .A(n43), .Y(n44) );
  NAND3BX1 U118 ( .AN(n87), .B(n2), .C(n46), .Y(n139) );
  INVX8 U119 ( .A(n190), .Y(n92) );
  AND2X4 U120 ( .A(n126), .B(n45), .Y(n146) );
  OR2X4 U121 ( .A(B[14]), .B(A[14]), .Y(n45) );
  NAND2XL U122 ( .A(A[10]), .B(B[10]), .Y(n179) );
  NAND2X4 U123 ( .A(n131), .B(n80), .Y(n173) );
  NAND2X4 U124 ( .A(A[14]), .B(B[14]), .Y(n149) );
  NAND3X4 U125 ( .A(n188), .B(n177), .C(n185), .Y(n74) );
  NAND2X4 U126 ( .A(n146), .B(n147), .Y(n49) );
  OAI21X4 U127 ( .A0(n79), .A1(n132), .B0(n133), .Y(n129) );
  NAND2X4 U128 ( .A(n163), .B(n162), .Y(n158) );
  BUFX20 U129 ( .A(n195), .Y(SUM[11]) );
  INVX4 U130 ( .A(A[16]), .Y(n118) );
  XOR2X4 U131 ( .A(n50), .B(n51), .Y(n193) );
  NAND2X4 U132 ( .A(n58), .B(n59), .Y(n50) );
  NAND2X4 U133 ( .A(B[4]), .B(A[4]), .Y(n98) );
  AOI21X2 U134 ( .A0(n138), .A1(n104), .B0(n139), .Y(n132) );
  NOR2BX2 U135 ( .AN(n76), .B(n73), .Y(n75) );
  NAND2X4 U136 ( .A(n78), .B(n18), .Y(n185) );
  NAND2X4 U137 ( .A(n153), .B(n152), .Y(n67) );
  NAND2X2 U138 ( .A(n19), .B(n36), .Y(n125) );
  NOR2X4 U139 ( .A(n125), .B(n124), .Y(n123) );
  NAND2X4 U140 ( .A(n121), .B(n120), .Y(n119) );
  NAND2X4 U141 ( .A(n123), .B(n122), .Y(n121) );
  XNOR2X4 U142 ( .A(n55), .B(n186), .Y(n196) );
  AND2X1 U143 ( .A(n31), .B(n183), .Y(n55) );
  NAND2X2 U144 ( .A(n127), .B(n29), .Y(n124) );
  AOI21X4 U145 ( .A0(n24), .A1(n76), .B0(n28), .Y(n176) );
  NOR2X4 U146 ( .A(n184), .B(n57), .Y(n181) );
  OAI21X4 U147 ( .A0(n178), .A1(n179), .B0(n140), .Y(n156) );
  INVX8 U148 ( .A(n145), .Y(n178) );
  NOR2BX4 U149 ( .AN(n142), .B(n178), .Y(n175) );
  NOR2X4 U150 ( .A(n173), .B(n174), .Y(n167) );
  OAI2BB1X4 U151 ( .A0N(n36), .A1N(n161), .B0(n164), .Y(n62) );
  INVX2 U152 ( .A(n158), .Y(n59) );
  XOR2X4 U153 ( .A(n81), .B(n82), .Y(n197) );
  INVX8 U154 ( .A(n137), .Y(n87) );
  NAND2X4 U155 ( .A(n46), .B(n69), .Y(n172) );
  INVX4 U156 ( .A(n94), .Y(n91) );
  XOR2X4 U157 ( .A(n89), .B(n90), .Y(SUM[6]) );
  NOR2BX2 U158 ( .AN(n88), .B(n53), .Y(n90) );
  OAI21X4 U159 ( .A0(n92), .A1(n98), .B0(n93), .Y(n136) );
  NAND2X2 U160 ( .A(B[5]), .B(A[5]), .Y(n93) );
  NOR2X4 U161 ( .A(n56), .B(n38), .Y(n57) );
  OAI21X4 U162 ( .A0(n181), .A1(n182), .B0(n183), .Y(n180) );
  NAND2X4 U163 ( .A(n72), .B(n54), .Y(n83) );
  OR2X4 U164 ( .A(A[3]), .B(B[3]), .Y(n106) );
  OR2X4 U165 ( .A(A[2]), .B(B[2]), .Y(n192) );
  NOR2XL U166 ( .A(A[0]), .B(B[0]), .Y(n68) );
  XNOR2X4 U167 ( .A(n67), .B(n151), .Y(n66) );
  OAI21X2 U168 ( .A0(n86), .A1(n53), .B0(n88), .Y(n81) );
  OAI21X4 U169 ( .A0(n96), .A1(n97), .B0(n98), .Y(n94) );
  OR2X4 U170 ( .A(B[11]), .B(A[11]), .Y(n145) );
  AND2X4 U171 ( .A(n192), .B(n106), .Y(n70) );
  NAND2X4 U172 ( .A(n70), .B(n191), .Y(n138) );
  INVXL U173 ( .A(n117), .Y(n113) );
  NOR2BX1 U174 ( .AN(n117), .B(n68), .Y(n199) );
  INVXL U175 ( .A(n46), .Y(n84) );
  NOR2X1 U176 ( .A(n78), .B(n79), .Y(n77) );
  OAI21XL U177 ( .A0(n107), .A1(n108), .B0(n109), .Y(n102) );
  NOR2BX1 U178 ( .AN(n104), .B(n105), .Y(n103) );
  NOR2BX1 U179 ( .AN(n109), .B(n108), .Y(n111) );
  INVX1 U180 ( .A(n192), .Y(n108) );
  XOR2X1 U181 ( .A(n113), .B(n115), .Y(SUM[1]) );
  OAI2BB1X1 U182 ( .A0N(n112), .A1N(n113), .B0(n114), .Y(n110) );
  INVX1 U183 ( .A(n106), .Y(n105) );
  NAND2X1 U184 ( .A(B[1]), .B(A[1]), .Y(n114) );
  NAND2X1 U185 ( .A(B[0]), .B(A[0]), .Y(n117) );
  NAND2X4 U186 ( .A(n104), .B(n138), .Y(n99) );
  NAND3XL U187 ( .A(n41), .B(n131), .C(n48), .Y(n130) );
  NAND2X2 U188 ( .A(A[9]), .B(B[9]), .Y(n76) );
  OAI21X4 U189 ( .A0(n91), .A1(n92), .B0(n93), .Y(n89) );
  CLKINVX3 U190 ( .A(n101), .Y(n96) );
  OR2X4 U191 ( .A(B[15]), .B(A[15]), .Y(n126) );
  OR2X4 U192 ( .A(A[14]), .B(B[14]), .Y(n127) );
  OR2X4 U193 ( .A(B[13]), .B(A[13]), .Y(n128) );
  NAND3BX4 U194 ( .AN(n156), .B(n141), .C(n157), .Y(n161) );
  NAND2X4 U195 ( .A(n167), .B(n168), .Y(n157) );
  NAND2X4 U196 ( .A(n176), .B(n175), .Y(n141) );
  XOR2X4 U197 ( .A(n180), .B(n4), .Y(n195) );
  OR2X4 U198 ( .A(B[11]), .B(A[11]), .Y(n131) );
  AOI21X4 U199 ( .A0(n74), .A1(n144), .B0(n187), .Y(n186) );
  OR2X4 U200 ( .A(A[7]), .B(B[7]), .Y(n85) );
  OAI211X2 U201 ( .A0(n116), .A1(n117), .B0(n114), .C0(n109), .Y(n191) );
  NAND2X4 U202 ( .A(B[2]), .B(A[2]), .Y(n109) );
  NAND2X4 U203 ( .A(B[3]), .B(A[3]), .Y(n104) );
  OR2X4 U204 ( .A(A[6]), .B(B[6]), .Y(n137) );
  OR2X4 U205 ( .A(A[5]), .B(B[5]), .Y(n190) );
  OR2X4 U206 ( .A(A[4]), .B(B[4]), .Y(n101) );
  OR2X4 U207 ( .A(B[9]), .B(A[9]), .Y(n144) );
  OR2X4 U208 ( .A(B[10]), .B(A[10]), .Y(n142) );
endmodule


module butterfly_DW01_add_52 ( A, B, SUM );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  wire   n173, n174, n175, n176, n1, n2, n3, n4, n5, n6, n7, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n34, n35, n36, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172;

  OR2XL U2 ( .A(A[15]), .B(B[15]), .Y(n1) );
  OR2XL U3 ( .A(B[7]), .B(A[7]), .Y(n56) );
  NOR2BX4 U4 ( .AN(n152), .B(n169), .Y(n167) );
  NOR2X2 U5 ( .A(A[9]), .B(B[9]), .Y(n158) );
  INVX4 U6 ( .A(n124), .Y(n123) );
  AOI21XL U7 ( .A0(n122), .A1(n78), .B0(n98), .Y(n117) );
  NOR2BX4 U8 ( .AN(n2), .B(n103), .Y(n156) );
  NAND2X4 U9 ( .A(n157), .B(n53), .Y(n2) );
  NOR2X4 U10 ( .A(n158), .B(n26), .Y(n155) );
  NOR2BX4 U11 ( .AN(n73), .B(n71), .Y(n75) );
  INVX4 U12 ( .A(n152), .Y(n71) );
  NAND3BX2 U13 ( .AN(n143), .B(n108), .C(n141), .Y(n105) );
  NAND3BX2 U14 ( .AN(B[13]), .B(n108), .C(n107), .Y(n106) );
  CLKINVX3 U15 ( .A(n29), .Y(n28) );
  OR2X2 U16 ( .A(A[4]), .B(B[4]), .Y(n152) );
  INVX4 U17 ( .A(n109), .Y(n143) );
  OR2X2 U18 ( .A(B[13]), .B(A[13]), .Y(n100) );
  BUFX3 U19 ( .A(B[4]), .Y(n34) );
  CLKBUFX8 U20 ( .A(n50), .Y(n10) );
  INVX2 U21 ( .A(n22), .Y(n61) );
  BUFX16 U22 ( .A(n174), .Y(SUM[14]) );
  OAI21XL U23 ( .A0(n81), .A1(n82), .B0(n83), .Y(n76) );
  INVX1 U24 ( .A(n5), .Y(n23) );
  NOR2BXL U25 ( .AN(n109), .B(n145), .Y(n144) );
  NOR2BX1 U26 ( .AN(n83), .B(n82), .Y(n85) );
  OAI2BB1X2 U27 ( .A0N(n10), .A1N(n47), .B0(n49), .Y(n6) );
  INVX8 U28 ( .A(n35), .Y(n36) );
  OAI2BB1X4 U29 ( .A0N(n139), .A1N(n138), .B0(n140), .Y(n136) );
  CLKBUFX2 U30 ( .A(n154), .Y(n17) );
  XNOR2X4 U31 ( .A(n6), .B(n162), .Y(n3) );
  NOR2BX1 U32 ( .AN(n126), .B(n29), .Y(n160) );
  CLKINVX3 U33 ( .A(n26), .Y(n4) );
  NOR2X4 U34 ( .A(B[11]), .B(A[11]), .Y(n26) );
  CLKBUFX8 U35 ( .A(n19), .Y(n16) );
  AND2X1 U36 ( .A(n36), .B(n163), .Y(n5) );
  INVX3 U37 ( .A(n114), .Y(n27) );
  NAND3X2 U38 ( .A(A[5]), .B(B[5]), .C(n150), .Y(n172) );
  INVX3 U39 ( .A(n103), .Y(n30) );
  NAND2X1 U40 ( .A(A[9]), .B(B[9]), .Y(n49) );
  NAND2XL U41 ( .A(n151), .B(n152), .Y(n15) );
  XOR2X4 U42 ( .A(n23), .B(n48), .Y(SUM[9]) );
  NAND2X2 U43 ( .A(n95), .B(n1), .Y(n128) );
  AND2X2 U44 ( .A(n125), .B(n25), .Y(n110) );
  INVX8 U45 ( .A(n7), .Y(SUM[12]) );
  NAND2BX4 U46 ( .AN(n55), .B(n57), .Y(n148) );
  NAND4BBX4 U47 ( .AN(n15), .BN(n67), .C(n9), .D(n74), .Y(n57) );
  NOR2BXL U48 ( .AN(n63), .B(n16), .Y(n65) );
  XOR2X2 U49 ( .A(n64), .B(n65), .Y(SUM[6]) );
  CLKINVX3 U50 ( .A(n175), .Y(n7) );
  XOR2X1 U51 ( .A(n138), .B(n144), .Y(n175) );
  AND2X1 U52 ( .A(n17), .B(n30), .Y(n162) );
  INVX8 U53 ( .A(n16), .Y(n9) );
  OAI21X4 U54 ( .A0(n62), .A1(n16), .B0(n63), .Y(n58) );
  INVXL U55 ( .A(n158), .Y(n11) );
  INVX2 U56 ( .A(n11), .Y(n12) );
  NAND2X4 U57 ( .A(n21), .B(n45), .Y(n134) );
  INVX8 U58 ( .A(n145), .Y(n21) );
  NAND2X4 U59 ( .A(n99), .B(n22), .Y(n13) );
  NAND2X2 U60 ( .A(n14), .B(n55), .Y(n163) );
  INVX4 U61 ( .A(n13), .Y(n14) );
  NOR2X2 U62 ( .A(B[15]), .B(A[15]), .Y(n115) );
  OR2X4 U63 ( .A(n159), .B(n39), .Y(n41) );
  NAND2X1 U64 ( .A(B[5]), .B(A[5]), .Y(n68) );
  CLKINVX4 U65 ( .A(n126), .Y(n24) );
  NAND2X2 U66 ( .A(n63), .B(n60), .Y(n170) );
  NAND2X4 U67 ( .A(A[9]), .B(B[9]), .Y(n157) );
  NAND2X4 U68 ( .A(A[12]), .B(B[12]), .Y(n109) );
  NAND2X4 U69 ( .A(n30), .B(n10), .Y(n120) );
  AND3X4 U70 ( .A(n121), .B(n4), .C(n50), .Y(n43) );
  INVX1 U71 ( .A(n132), .Y(n140) );
  OAI2BB1X1 U72 ( .A0N(n22), .A1N(n55), .B0(n57), .Y(n51) );
  AOI21X4 U73 ( .A0(n132), .A1(n27), .B0(n133), .Y(n131) );
  AND2X2 U74 ( .A(n100), .B(n141), .Y(n31) );
  NAND3X4 U75 ( .A(n113), .B(n18), .C(n100), .Y(n112) );
  AND2X4 U76 ( .A(n28), .B(n97), .Y(n18) );
  NOR2X2 U77 ( .A(A[6]), .B(B[6]), .Y(n19) );
  BUFX20 U78 ( .A(n173), .Y(SUM[15]) );
  INVX1 U79 ( .A(n134), .Y(n139) );
  CLKBUFX2 U80 ( .A(n55), .Y(n20) );
  INVXL U81 ( .A(n108), .Y(n133) );
  BUFX4 U82 ( .A(n26), .Y(n29) );
  INVX8 U83 ( .A(n97), .Y(n145) );
  BUFX8 U84 ( .A(n56), .Y(n22) );
  NAND2BX4 U85 ( .AN(n134), .B(n27), .Y(n130) );
  NAND2X4 U86 ( .A(A[13]), .B(B[13]), .Y(n141) );
  INVX8 U87 ( .A(n121), .Y(n103) );
  NOR2X4 U88 ( .A(n123), .B(n24), .Y(n25) );
  NAND2X2 U89 ( .A(B[11]), .B(A[11]), .Y(n126) );
  NOR2X2 U90 ( .A(B[14]), .B(A[14]), .Y(n114) );
  NOR2X4 U91 ( .A(n120), .B(n119), .Y(n118) );
  NOR2X4 U92 ( .A(n114), .B(n115), .Y(n113) );
  NAND2X2 U93 ( .A(A[7]), .B(B[7]), .Y(n60) );
  OAI21X4 U94 ( .A0(n117), .A1(n20), .B0(n118), .Y(n111) );
  NAND2X1 U95 ( .A(A[15]), .B(B[15]), .Y(n95) );
  NOR2BX2 U96 ( .AN(n60), .B(n61), .Y(n59) );
  NAND2X2 U97 ( .A(B[6]), .B(A[6]), .Y(n63) );
  NAND3BX2 U98 ( .AN(n73), .B(n150), .C(n149), .Y(n171) );
  INVX8 U99 ( .A(n149), .Y(n67) );
  BUFX16 U100 ( .A(n176), .Y(SUM[7]) );
  INVX4 U101 ( .A(n64), .Y(n62) );
  AND3X4 U102 ( .A(n125), .B(n124), .C(n126), .Y(n44) );
  NAND2X4 U103 ( .A(n164), .B(n53), .Y(n35) );
  AOI21X4 U104 ( .A0(n138), .A1(n21), .B0(n143), .Y(n142) );
  OAI2BB1X4 U105 ( .A0N(n30), .A1N(n161), .B0(n17), .Y(n159) );
  NAND2X2 U106 ( .A(n124), .B(n126), .Y(n153) );
  OR2X4 U107 ( .A(B[13]), .B(A[13]), .Y(n45) );
  INVX2 U108 ( .A(n99), .Y(n54) );
  NAND2XL U109 ( .A(n108), .B(n101), .Y(n137) );
  INVX8 U110 ( .A(n74), .Y(n72) );
  NAND3X4 U111 ( .A(n43), .B(n147), .C(n148), .Y(n135) );
  NAND2X2 U112 ( .A(n159), .B(n39), .Y(n40) );
  NOR2BX4 U113 ( .AN(n53), .B(n54), .Y(n52) );
  NAND2X4 U114 ( .A(n101), .B(n102), .Y(n104) );
  NAND3BX4 U115 ( .AN(n98), .B(n74), .C(n99), .Y(n164) );
  NAND2X4 U116 ( .A(n96), .B(n95), .Y(n94) );
  NAND2BX4 U117 ( .AN(n154), .B(n116), .Y(n124) );
  AND2X4 U118 ( .A(n44), .B(n135), .Y(n129) );
  NOR2X4 U119 ( .A(n19), .B(n67), .Y(n168) );
  XNOR2X4 U120 ( .A(n142), .B(n31), .Y(SUM[13]) );
  OAI21X4 U121 ( .A0(n71), .A1(n72), .B0(n73), .Y(n69) );
  XOR2X2 U122 ( .A(n69), .B(n70), .Y(SUM[5]) );
  INVX4 U123 ( .A(n69), .Y(n66) );
  NAND3BX4 U124 ( .AN(n104), .B(n105), .C(n106), .Y(n96) );
  NAND2X4 U125 ( .A(A[14]), .B(B[14]), .Y(n108) );
  INVX4 U126 ( .A(n151), .Y(n169) );
  XOR2X4 U127 ( .A(n58), .B(n59), .Y(n176) );
  NAND2X2 U128 ( .A(B[2]), .B(A[2]), .Y(n83) );
  AOI21X4 U129 ( .A0(n111), .A1(n110), .B0(n112), .Y(n93) );
  NAND2X1 U130 ( .A(n99), .B(n22), .Y(n119) );
  NAND2X4 U131 ( .A(n167), .B(n168), .Y(n98) );
  NOR2X4 U132 ( .A(n93), .B(n94), .Y(n92) );
  OR2X4 U133 ( .A(A[2]), .B(B[2]), .Y(n166) );
  OAI2BB1X4 U134 ( .A0N(n10), .A1N(n47), .B0(n49), .Y(n161) );
  NAND2X4 U135 ( .A(n34), .B(A[4]), .Y(n73) );
  XOR2X4 U136 ( .A(n51), .B(n52), .Y(SUM[8]) );
  NAND2X4 U137 ( .A(n36), .B(n163), .Y(n47) );
  NAND2X4 U138 ( .A(B[8]), .B(A[8]), .Y(n53) );
  INVX8 U139 ( .A(n3), .Y(SUM[10]) );
  NAND2X4 U140 ( .A(n40), .B(n41), .Y(SUM[11]) );
  INVX1 U141 ( .A(n160), .Y(n39) );
  OAI21X4 U142 ( .A0(n66), .A1(n67), .B0(n68), .Y(n64) );
  NAND2X2 U143 ( .A(B[10]), .B(A[10]), .Y(n154) );
  NOR2BX1 U144 ( .AN(n49), .B(n12), .Y(n48) );
  NOR2XL U145 ( .A(A[0]), .B(B[0]), .Y(n42) );
  NAND2X1 U146 ( .A(B[3]), .B(A[3]), .Y(n78) );
  INVXL U147 ( .A(n166), .Y(n82) );
  INVXL U148 ( .A(n91), .Y(n87) );
  NAND2X4 U149 ( .A(n78), .B(n122), .Y(n74) );
  NOR2BX1 U150 ( .AN(n91), .B(n42), .Y(SUM[0]) );
  XOR2X1 U151 ( .A(n84), .B(n85), .Y(SUM[2]) );
  XNOR2X4 U152 ( .A(n127), .B(n128), .Y(n173) );
  XNOR2X4 U153 ( .A(n136), .B(n137), .Y(n174) );
  NOR2BXL U154 ( .AN(n68), .B(n67), .Y(n70) );
  XOR2X1 U155 ( .A(n74), .B(n75), .Y(SUM[4]) );
  XOR2X1 U156 ( .A(n87), .B(n89), .Y(SUM[1]) );
  NOR2BXL U157 ( .AN(n88), .B(n90), .Y(n89) );
  OAI2BB1X1 U158 ( .A0N(n86), .A1N(n87), .B0(n88), .Y(n84) );
  OAI2BB1X4 U159 ( .A0N(n45), .A1N(n143), .B0(n141), .Y(n132) );
  NAND2X1 U160 ( .A(B[1]), .B(A[1]), .Y(n88) );
  NAND2X4 U161 ( .A(n46), .B(n165), .Y(n122) );
  AND2X4 U162 ( .A(n166), .B(n80), .Y(n46) );
  INVX1 U163 ( .A(A[13]), .Y(n107) );
  XOR2X1 U164 ( .A(n76), .B(n77), .Y(SUM[3]) );
  NOR2BX1 U165 ( .AN(n78), .B(n79), .Y(n77) );
  INVX1 U166 ( .A(n84), .Y(n81) );
  NAND2X1 U167 ( .A(B[0]), .B(A[0]), .Y(n91) );
  INVXL U168 ( .A(n80), .Y(n79) );
  XNOR3X4 U169 ( .A(B[16]), .B(A[16]), .C(n92), .Y(SUM[16]) );
  OR2X4 U170 ( .A(A[15]), .B(B[15]), .Y(n102) );
  OAI21X4 U171 ( .A0(n129), .A1(n130), .B0(n131), .Y(n127) );
  OR2X4 U172 ( .A(B[14]), .B(A[14]), .Y(n101) );
  OR2X4 U173 ( .A(B[12]), .B(A[12]), .Y(n97) );
  NAND2X4 U174 ( .A(n146), .B(n135), .Y(n138) );
  NOR2X4 U175 ( .A(n61), .B(n54), .Y(n147) );
  NOR2BX4 U176 ( .AN(n125), .B(n153), .Y(n146) );
  NAND2X4 U177 ( .A(n156), .B(n155), .Y(n125) );
  OR2X4 U178 ( .A(B[11]), .B(A[11]), .Y(n116) );
  OR2X4 U179 ( .A(B[10]), .B(A[10]), .Y(n121) );
  OAI211X2 U180 ( .A0(n90), .A1(n91), .B0(n88), .C0(n83), .Y(n165) );
  CLKINVX3 U181 ( .A(n86), .Y(n90) );
  OR2X4 U182 ( .A(A[3]), .B(B[3]), .Y(n80) );
  OR2X4 U183 ( .A(A[1]), .B(B[1]), .Y(n86) );
  OR2X4 U184 ( .A(B[7]), .B(A[7]), .Y(n151) );
  NAND3BX4 U185 ( .AN(n170), .B(n171), .C(n172), .Y(n55) );
  OR2X4 U186 ( .A(A[5]), .B(B[5]), .Y(n149) );
  OR2X4 U187 ( .A(A[6]), .B(B[6]), .Y(n150) );
  OR2X4 U188 ( .A(A[8]), .B(B[8]), .Y(n99) );
  OR2X4 U189 ( .A(A[9]), .B(B[9]), .Y(n50) );
endmodule


module butterfly_DW01_add_56 ( A, B, SUM );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  wire   n189, n190, n191, n192, n193, n194, n195, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188;

  INVX8 U2 ( .A(n170), .Y(n167) );
  NOR2X2 U3 ( .A(n167), .B(n162), .Y(n1) );
  NAND3X2 U4 ( .A(n20), .B(n157), .C(n159), .Y(n155) );
  INVX4 U5 ( .A(n5), .Y(n27) );
  NAND2X2 U6 ( .A(B[14]), .B(A[14]), .Y(n126) );
  BUFX8 U7 ( .A(n62), .Y(n11) );
  INVX3 U8 ( .A(n81), .Y(n77) );
  INVX1 U9 ( .A(n4), .Y(n89) );
  NAND3X4 U10 ( .A(n156), .B(n155), .C(n128), .Y(n153) );
  OAI21X4 U11 ( .A0(n62), .A1(n60), .B0(n59), .Y(n95) );
  OAI2BB1X4 U12 ( .A0N(n151), .A1N(n122), .B0(n126), .Y(n149) );
  NAND2X2 U13 ( .A(n69), .B(n175), .Y(n172) );
  NOR2X4 U14 ( .A(n62), .B(n60), .Y(n186) );
  OAI21X4 U15 ( .A0(n172), .A1(n67), .B0(n173), .Y(n30) );
  BUFX8 U16 ( .A(n166), .Y(n2) );
  OR2X4 U17 ( .A(B[9]), .B(A[9]), .Y(n175) );
  AOI2BB1X4 U18 ( .A0N(B[9]), .A1N(A[9]), .B0(n167), .Y(n163) );
  INVX20 U19 ( .A(n44), .Y(SUM[1]) );
  CLKINVX2 U20 ( .A(n73), .Y(n148) );
  INVX1 U21 ( .A(n12), .Y(n87) );
  INVX1 U22 ( .A(n55), .Y(n38) );
  BUFX4 U23 ( .A(n79), .Y(n18) );
  INVX4 U24 ( .A(n175), .Y(n66) );
  NAND2X1 U25 ( .A(B[10]), .B(A[10]), .Y(n166) );
  INVX1 U26 ( .A(n139), .Y(n138) );
  INVX1 U27 ( .A(n118), .Y(n117) );
  OAI21XL U28 ( .A0(n119), .A1(n120), .B0(n121), .Y(n118) );
  NAND2X1 U29 ( .A(n132), .B(n133), .Y(n116) );
  BUFX20 U30 ( .A(B[2]), .Y(n60) );
  NAND2X1 U31 ( .A(n146), .B(n145), .Y(n101) );
  AND2X4 U32 ( .A(n82), .B(n83), .Y(n3) );
  BUFX8 U33 ( .A(n107), .Y(n14) );
  NOR2X2 U34 ( .A(n62), .B(n60), .Y(n147) );
  NOR2X4 U35 ( .A(B[3]), .B(A[3]), .Y(n4) );
  NOR2X2 U36 ( .A(A[3]), .B(B[3]), .Y(n31) );
  OR2X4 U37 ( .A(n61), .B(n59), .Y(n185) );
  NAND2BX4 U38 ( .AN(n143), .B(n100), .Y(n75) );
  NOR2BXL U39 ( .AN(n73), .B(n54), .Y(n72) );
  OAI21X2 U40 ( .A0(n18), .A1(n7), .B0(n23), .Y(n78) );
  XOR2X4 U41 ( .A(n108), .B(n109), .Y(n50) );
  NAND3X4 U42 ( .A(n178), .B(n180), .C(n179), .Y(n5) );
  OAI2BB1X4 U43 ( .A0N(n170), .A1N(n171), .B0(n2), .Y(n32) );
  AOI21X4 U44 ( .A0(n146), .A1(n145), .B0(n102), .Y(n100) );
  NAND2X2 U45 ( .A(B[7]), .B(A[7]), .Y(n73) );
  NAND3X4 U46 ( .A(n181), .B(n182), .C(n14), .Y(n177) );
  CLKINVX4 U47 ( .A(n57), .Y(n6) );
  INVX8 U48 ( .A(n61), .Y(n57) );
  CLKBUFX2 U49 ( .A(n80), .Y(n23) );
  BUFX20 U50 ( .A(n193), .Y(SUM[9]) );
  INVX2 U51 ( .A(n83), .Y(n7) );
  OR2X4 U52 ( .A(A[6]), .B(B[6]), .Y(n83) );
  INVX8 U53 ( .A(n47), .Y(SUM[8]) );
  XOR2X4 U54 ( .A(n48), .B(n37), .Y(n47) );
  INVX8 U55 ( .A(n50), .Y(SUM[2]) );
  AND2X2 U56 ( .A(n23), .B(n83), .Y(n8) );
  NOR2X4 U57 ( .A(n59), .B(n61), .Y(n130) );
  NAND2X2 U58 ( .A(n1), .B(n169), .Y(n9) );
  DLY1X1 U59 ( .A(n143), .Y(n10) );
  NAND2X2 U60 ( .A(n65), .B(n68), .Y(n164) );
  OAI21XL U61 ( .A0(n142), .A1(n10), .B0(n144), .Y(n141) );
  OR2X2 U62 ( .A(n77), .B(n102), .Y(n90) );
  NAND2BXL U63 ( .AN(n12), .B(n82), .Y(n86) );
  NAND2X4 U64 ( .A(n103), .B(n104), .Y(n143) );
  AOI21X2 U65 ( .A0(n77), .A1(n3), .B0(n78), .Y(n76) );
  OR2X4 U66 ( .A(n60), .B(n62), .Y(n26) );
  NAND2XL U67 ( .A(n60), .B(n62), .Y(n92) );
  INVXL U68 ( .A(n69), .Y(n15) );
  AND2X4 U69 ( .A(n59), .B(n61), .Y(n29) );
  AND2X2 U70 ( .A(n3), .B(n87), .Y(n74) );
  AOI2BB1X4 U71 ( .A0N(n66), .A1N(n68), .B0(n174), .Y(n173) );
  NOR2X4 U72 ( .A(A[4]), .B(B[4]), .Y(n12) );
  INVX2 U73 ( .A(n82), .Y(n13) );
  OR2X4 U74 ( .A(B[5]), .B(A[5]), .Y(n82) );
  OAI21X4 U75 ( .A0(n15), .A1(n67), .B0(n68), .Y(n63) );
  NOR2X2 U76 ( .A(n129), .B(n4), .Y(n16) );
  NOR2BX1 U77 ( .AN(n81), .B(n12), .Y(n99) );
  NOR2BX1 U78 ( .AN(n18), .B(n13), .Y(n98) );
  NAND3X4 U79 ( .A(n80), .B(n79), .C(n81), .Y(n180) );
  INVX2 U80 ( .A(n99), .Y(n46) );
  NAND2BX4 U81 ( .AN(n143), .B(n100), .Y(n17) );
  OAI211X2 U82 ( .A0(n60), .A1(n62), .B0(n6), .C0(n59), .Y(n182) );
  BUFX20 U83 ( .A(n189), .Y(SUM[15]) );
  NAND2XL U84 ( .A(n68), .B(n69), .Y(n48) );
  CLKINVX4 U85 ( .A(n57), .Y(n58) );
  AND2X2 U86 ( .A(B[11]), .B(A[11]), .Y(n19) );
  INVXL U87 ( .A(n162), .Y(n20) );
  INVXL U88 ( .A(n19), .Y(n21) );
  INVXL U89 ( .A(n102), .Y(n22) );
  CLKINVX8 U90 ( .A(n91), .Y(n102) );
  DLY1X1 U91 ( .A(n140), .Y(n24) );
  NAND2X2 U92 ( .A(B[9]), .B(A[9]), .Y(n65) );
  AND2X2 U93 ( .A(n21), .B(n158), .Y(n33) );
  OR2X4 U94 ( .A(n62), .B(n60), .Y(n28) );
  NOR2X4 U95 ( .A(n130), .B(n96), .Y(n94) );
  INVX8 U96 ( .A(n158), .Y(n162) );
  OAI2BB1X4 U97 ( .A0N(n26), .A1N(n108), .B0(n14), .Y(n105) );
  NOR2BX2 U98 ( .AN(n91), .B(n4), .Y(n106) );
  NOR2X4 U99 ( .A(n27), .B(n148), .Y(n140) );
  OAI21X2 U100 ( .A0(n9), .A1(n67), .B0(n139), .Y(n160) );
  OAI21X4 U101 ( .A0(n58), .A1(n59), .B0(n110), .Y(n113) );
  NAND3BX4 U102 ( .AN(n31), .B(n28), .C(n29), .Y(n103) );
  NOR2BX4 U103 ( .AN(n69), .B(n66), .Y(n169) );
  NOR2X4 U104 ( .A(n129), .B(n4), .Y(n176) );
  NOR2BX4 U105 ( .AN(n2), .B(n19), .Y(n165) );
  OAI2BB1X4 U106 ( .A0N(n16), .A1N(n177), .B0(n140), .Y(n37) );
  NAND2X4 U107 ( .A(n61), .B(n59), .Y(n110) );
  OAI21X4 U108 ( .A0(n61), .A1(n59), .B0(n112), .Y(n111) );
  AOI2BB2X4 U109 ( .B0(n26), .B1(n94), .A0N(n95), .A1N(n57), .Y(n93) );
  OAI21X4 U110 ( .A0(n115), .A1(n116), .B0(n117), .Y(n114) );
  XNOR2X4 U111 ( .A(n32), .B(n33), .Y(n51) );
  BUFX20 U112 ( .A(A[1]), .Y(n61) );
  INVX8 U113 ( .A(n52), .Y(SUM[10]) );
  XNOR2X4 U114 ( .A(n30), .B(n53), .Y(n52) );
  BUFX20 U115 ( .A(n194), .Y(SUM[7]) );
  INVX20 U116 ( .A(n45), .Y(SUM[4]) );
  INVX4 U117 ( .A(n157), .Y(n136) );
  NOR2BX2 U118 ( .AN(n128), .B(n136), .Y(n161) );
  NAND2X4 U119 ( .A(B[12]), .B(A[12]), .Y(n128) );
  AOI21X4 U120 ( .A0(n88), .A1(n89), .B0(n90), .Y(n85) );
  XOR2X2 U121 ( .A(n17), .B(n46), .Y(n45) );
  BUFX20 U122 ( .A(B[1]), .Y(n59) );
  DLY1X1 U123 ( .A(n129), .Y(n34) );
  INVX8 U124 ( .A(n70), .Y(n67) );
  BUFX20 U125 ( .A(n190), .Y(SUM[14]) );
  AOI21X4 U126 ( .A0(n185), .A1(n184), .B0(n102), .Y(n181) );
  OR2X4 U127 ( .A(A[11]), .B(B[11]), .Y(n158) );
  NOR2X4 U128 ( .A(A[5]), .B(B[5]), .Y(n35) );
  NOR2X4 U129 ( .A(n54), .B(n36), .Y(n179) );
  NOR2X4 U130 ( .A(B[7]), .B(A[7]), .Y(n54) );
  NAND2BX4 U131 ( .AN(n162), .B(n159), .Y(n139) );
  NAND3BX4 U132 ( .AN(n131), .B(n157), .C(n37), .Y(n156) );
  NOR2X4 U133 ( .A(A[6]), .B(B[6]), .Y(n36) );
  NOR2X4 U134 ( .A(n186), .B(n96), .Y(n184) );
  NOR2BX1 U135 ( .AN(n65), .B(n66), .Y(n64) );
  NAND2X2 U136 ( .A(n80), .B(n35), .Y(n178) );
  OAI2BB1X4 U137 ( .A0N(n153), .A1N(n38), .B0(n127), .Y(n151) );
  BUFX20 U138 ( .A(n195), .Y(SUM[6]) );
  BUFX20 U139 ( .A(n192), .Y(SUM[12]) );
  XOR2X4 U140 ( .A(n113), .B(n112), .Y(n44) );
  NAND2X4 U141 ( .A(A[4]), .B(B[4]), .Y(n81) );
  OAI2BB1X4 U142 ( .A0N(n74), .A1N(n17), .B0(n76), .Y(n71) );
  NAND2X4 U143 ( .A(n111), .B(n110), .Y(n108) );
  BUFX20 U144 ( .A(n191), .Y(SUM[13]) );
  OAI21X4 U145 ( .A0(n85), .A1(n86), .B0(n18), .Y(n84) );
  NAND2X4 U146 ( .A(B[5]), .B(A[5]), .Y(n79) );
  NAND2X4 U147 ( .A(B[6]), .B(A[6]), .Y(n80) );
  OAI2BB1X4 U148 ( .A0N(n87), .A1N(n75), .B0(n81), .Y(n97) );
  NAND2X4 U149 ( .A(n93), .B(n92), .Y(n88) );
  NAND2X4 U150 ( .A(B[8]), .B(A[8]), .Y(n68) );
  NAND3BX4 U151 ( .AN(n31), .B(n60), .C(n11), .Y(n104) );
  AOI2BB1X4 U152 ( .A0N(n59), .A1N(n61), .B0(n96), .Y(n145) );
  OAI21X4 U153 ( .A0(n67), .A1(n172), .B0(n173), .Y(n171) );
  INVX8 U154 ( .A(n51), .Y(SUM[11]) );
  XNOR2X4 U155 ( .A(n114), .B(n49), .Y(SUM[16]) );
  NAND2XL U156 ( .A(B[15]), .B(A[15]), .Y(n121) );
  NOR2BX4 U157 ( .AN(n126), .B(n135), .Y(n152) );
  NOR2BX4 U158 ( .AN(n121), .B(n134), .Y(n150) );
  NOR2XL U159 ( .A(n55), .B(n128), .Y(n124) );
  OR2X4 U160 ( .A(A[15]), .B(B[15]), .Y(n123) );
  OR2X4 U161 ( .A(A[14]), .B(B[14]), .Y(n122) );
  XNOR2X1 U162 ( .A(B[16]), .B(A[16]), .Y(n49) );
  INVX1 U163 ( .A(n65), .Y(n174) );
  NOR2X1 U164 ( .A(n137), .B(n138), .Y(n115) );
  AOI21XL U165 ( .A0(n141), .A1(n24), .B0(n9), .Y(n137) );
  INVX1 U166 ( .A(n122), .Y(n135) );
  AND2X1 U167 ( .A(n2), .B(n170), .Y(n53) );
  NAND2XL U168 ( .A(n22), .B(n101), .Y(n142) );
  INVXL U169 ( .A(n34), .Y(n144) );
  INVX1 U170 ( .A(n123), .Y(n134) );
  NAND2XL U171 ( .A(n126), .B(n127), .Y(n125) );
  NOR2XL U172 ( .A(n134), .B(n135), .Y(n133) );
  NOR2XL U173 ( .A(n55), .B(n136), .Y(n132) );
  NAND2X1 U174 ( .A(n122), .B(n123), .Y(n120) );
  NOR2X1 U175 ( .A(n124), .B(n125), .Y(n119) );
  NOR2X4 U176 ( .A(A[13]), .B(B[13]), .Y(n55) );
  INVX1 U177 ( .A(n96), .Y(n112) );
  AND2X2 U178 ( .A(n96), .B(n183), .Y(SUM[0]) );
  OR2X2 U179 ( .A(A[0]), .B(B[0]), .Y(n183) );
  NAND2X1 U180 ( .A(B[0]), .B(A[0]), .Y(n96) );
  BUFX20 U181 ( .A(A[2]), .Y(n62) );
  NOR2X4 U182 ( .A(n147), .B(n4), .Y(n146) );
  NAND2X2 U183 ( .A(A[3]), .B(B[3]), .Y(n91) );
  XOR2X4 U184 ( .A(n63), .B(n64), .Y(n193) );
  XOR2X4 U185 ( .A(n71), .B(n72), .Y(n194) );
  XOR2X4 U186 ( .A(n84), .B(n8), .Y(n195) );
  XOR2X4 U187 ( .A(n97), .B(n98), .Y(SUM[5]) );
  XOR2X4 U188 ( .A(n105), .B(n106), .Y(SUM[3]) );
  OAI21X4 U189 ( .A0(n11), .A1(n60), .B0(n107), .Y(n109) );
  NAND2X4 U190 ( .A(n60), .B(n62), .Y(n107) );
  XOR2X4 U191 ( .A(n149), .B(n150), .Y(n189) );
  XOR2X4 U192 ( .A(n151), .B(n152), .Y(n190) );
  XOR2X4 U193 ( .A(n153), .B(n154), .Y(n191) );
  NOR2BX4 U194 ( .AN(n127), .B(n55), .Y(n154) );
  NAND2X4 U195 ( .A(B[13]), .B(A[13]), .Y(n127) );
  XOR2X4 U196 ( .A(n160), .B(n161), .Y(n192) );
  OR2X4 U197 ( .A(A[12]), .B(B[12]), .Y(n157) );
  OAI2BB1X4 U198 ( .A0N(n163), .A1N(n164), .B0(n165), .Y(n159) );
  NAND2X4 U199 ( .A(n168), .B(n169), .Y(n131) );
  NOR2X4 U200 ( .A(n167), .B(n162), .Y(n168) );
  OR2X4 U201 ( .A(A[10]), .B(B[10]), .Y(n170) );
  OR2X4 U202 ( .A(A[8]), .B(B[8]), .Y(n69) );
  OAI2BB1X4 U203 ( .A0N(n176), .A1N(n177), .B0(n140), .Y(n70) );
  NAND2X4 U204 ( .A(n187), .B(n188), .Y(n129) );
  NOR2X4 U205 ( .A(n54), .B(n36), .Y(n188) );
  NOR2X4 U206 ( .A(n12), .B(n35), .Y(n187) );
endmodule


module butterfly_DW01_sub_56 ( A, B, DIFF );
  input [16:0] A;
  input [16:0] B;
  output [16:0] DIFF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181;

  INVX1 U3 ( .A(n80), .Y(n77) );
  NAND2BX1 U4 ( .AN(n163), .B(n16), .Y(n160) );
  NAND4BXL U5 ( .AN(n57), .B(n156), .C(n103), .D(n28), .Y(n88) );
  AND2X4 U6 ( .A(n127), .B(n117), .Y(n25) );
  NAND2BX4 U7 ( .AN(A[9]), .B(B[9]), .Y(n153) );
  NAND2X4 U8 ( .A(n1), .B(n29), .Y(n176) );
  NAND2BX4 U9 ( .AN(A[8]), .B(B[8]), .Y(n170) );
  NAND2X4 U10 ( .A(n149), .B(n43), .Y(n175) );
  BUFX20 U11 ( .A(n174), .Y(n29) );
  OR2X4 U12 ( .A(n13), .B(B[10]), .Y(n155) );
  NAND2BX4 U13 ( .AN(A[3]), .B(B[3]), .Y(n180) );
  BUFX20 U14 ( .A(n41), .Y(n15) );
  BUFX16 U15 ( .A(n40), .Y(n1) );
  NAND2BX4 U16 ( .AN(A[15]), .B(B[15]), .Y(n110) );
  INVXL U17 ( .A(A[10]), .Y(n13) );
  NAND2X1 U18 ( .A(n96), .B(n108), .Y(n22) );
  NOR2X2 U19 ( .A(n175), .B(n176), .Y(n171) );
  CLKINVX3 U20 ( .A(n98), .Y(n126) );
  CLKINVX3 U21 ( .A(n7), .Y(n8) );
  NAND2X2 U22 ( .A(n79), .B(n82), .Y(n178) );
  NAND2BX1 U23 ( .AN(B[15]), .B(A[15]), .Y(n94) );
  INVX1 U24 ( .A(n110), .Y(n100) );
  INVX1 U25 ( .A(n76), .Y(n74) );
  OAI21X2 U26 ( .A0(n77), .A1(n78), .B0(n79), .Y(n73) );
  INVX4 U27 ( .A(n72), .Y(n75) );
  INVX1 U28 ( .A(n170), .Y(n35) );
  INVX1 U29 ( .A(n39), .Y(n31) );
  NAND4X2 U30 ( .A(n72), .B(n83), .C(n179), .D(n180), .Y(n57) );
  INVX1 U31 ( .A(n104), .Y(n103) );
  NAND2BX2 U32 ( .AN(B[0]), .B(A[0]), .Y(n82) );
  NOR2X2 U33 ( .A(n61), .B(n62), .Y(n20) );
  NAND3X2 U34 ( .A(n43), .B(n29), .C(n15), .Y(n64) );
  NOR2X2 U35 ( .A(n47), .B(n48), .Y(n46) );
  INVX2 U36 ( .A(n49), .Y(n47) );
  AND2X1 U37 ( .A(n8), .B(n155), .Y(n2) );
  AND2X1 U38 ( .A(n154), .B(n120), .Y(n3) );
  NAND2BX2 U39 ( .AN(B[11]), .B(A[11]), .Y(n120) );
  INVX2 U40 ( .A(n174), .Y(n148) );
  NAND2X1 U41 ( .A(n42), .B(n43), .Y(n166) );
  INVX2 U42 ( .A(n112), .Y(n7) );
  BUFX8 U43 ( .A(n55), .Y(n4) );
  NAND3BX4 U44 ( .AN(n165), .B(n113), .C(n114), .Y(n172) );
  NAND2BX2 U45 ( .AN(B[3]), .B(A[3]), .Y(n59) );
  NAND2XL U46 ( .A(n4), .B(n54), .Y(n63) );
  AND2X4 U47 ( .A(n5), .B(B[7]), .Y(n6) );
  INVX1 U48 ( .A(A[7]), .Y(n5) );
  CLKINVX8 U49 ( .A(n6), .Y(n173) );
  NAND2BX4 U50 ( .AN(A[5]), .B(B[5]), .Y(n174) );
  NAND3X4 U51 ( .A(n153), .B(n112), .C(n154), .Y(n17) );
  AND2X1 U52 ( .A(n116), .B(n117), .Y(n105) );
  INVXL U53 ( .A(n33), .Y(n9) );
  NAND2X2 U54 ( .A(n16), .B(n153), .Y(n144) );
  XNOR2X4 U55 ( .A(n10), .B(n30), .Y(DIFF[9]) );
  AND2X1 U56 ( .A(n153), .B(n36), .Y(n10) );
  OAI21XL U57 ( .A0(n111), .A1(n9), .B0(n28), .Y(n106) );
  NAND2BX2 U58 ( .AN(A[10]), .B(B[10]), .Y(n16) );
  INVX4 U59 ( .A(n17), .Y(n18) );
  AOI21X2 U60 ( .A0(n15), .A1(n171), .B0(n172), .Y(n168) );
  AND2X2 U61 ( .A(n94), .B(n110), .Y(n11) );
  INVX2 U62 ( .A(n155), .Y(n118) );
  NOR2X2 U63 ( .A(n166), .B(n176), .Y(n164) );
  NAND2BX4 U64 ( .AN(A[11]), .B(B[11]), .Y(n154) );
  NAND2BX2 U65 ( .AN(A[11]), .B(B[11]), .Y(n156) );
  AND2X4 U66 ( .A(n15), .B(n142), .Y(n12) );
  NAND2X2 U67 ( .A(n29), .B(n1), .Y(n51) );
  NAND4BX1 U68 ( .AN(n148), .B(n149), .C(n1), .D(n150), .Y(n147) );
  INVX4 U69 ( .A(n1), .Y(n62) );
  CLKINVX3 U70 ( .A(n162), .Y(n14) );
  INVX2 U71 ( .A(n36), .Y(n162) );
  NAND2BX4 U72 ( .AN(A[14]), .B(B[14]), .Y(n102) );
  OAI21X4 U73 ( .A0(n168), .A1(n163), .B0(n14), .Y(n167) );
  INVX8 U74 ( .A(n44), .Y(n33) );
  NAND3X4 U75 ( .A(n113), .B(n49), .C(n114), .Y(n44) );
  OAI21X1 U76 ( .A0(n88), .A1(n89), .B0(n90), .Y(n87) );
  AOI21X2 U77 ( .A0(n91), .A1(n92), .B0(n93), .Y(n90) );
  NAND2BX4 U78 ( .AN(B[13]), .B(A[13]), .Y(n99) );
  NAND2BX4 U79 ( .AN(A[7]), .B(B[7]), .Y(n149) );
  NAND4BX2 U80 ( .AN(n152), .B(n112), .C(n153), .D(n154), .Y(n151) );
  NOR2X2 U81 ( .A(n143), .B(n176), .Y(n142) );
  OAI2BB1X2 U82 ( .A0N(n169), .A1N(B[9]), .B0(n170), .Y(n163) );
  NOR2X4 U83 ( .A(n65), .B(n68), .Y(n67) );
  INVX8 U84 ( .A(n69), .Y(n65) );
  NAND2BX2 U85 ( .AN(B[2]), .B(A[2]), .Y(n76) );
  INVX8 U86 ( .A(n179), .Y(n78) );
  XOR2X2 U87 ( .A(n80), .B(n21), .Y(DIFF[1]) );
  NOR2X4 U88 ( .A(n81), .B(n78), .Y(n21) );
  NAND2BX4 U89 ( .AN(n136), .B(n102), .Y(n122) );
  NAND2BX4 U90 ( .AN(A[13]), .B(B[13]), .Y(n109) );
  NAND2X2 U91 ( .A(n54), .B(n4), .Y(n53) );
  NOR2X2 U92 ( .A(n86), .B(n87), .Y(n84) );
  NAND2X4 U93 ( .A(n39), .B(n49), .Y(n165) );
  OAI21X2 U94 ( .A0(n48), .A1(n52), .B0(n49), .Y(n146) );
  NAND2BX4 U95 ( .AN(B[7]), .B(A[7]), .Y(n49) );
  AOI21X4 U96 ( .A0(n33), .A1(n34), .B0(n35), .Y(n32) );
  NAND2X2 U97 ( .A(n36), .B(n39), .Y(n157) );
  NAND2BX4 U98 ( .AN(B[8]), .B(A[8]), .Y(n39) );
  NAND2BX4 U99 ( .AN(n136), .B(n135), .Y(n133) );
  AOI21X2 U100 ( .A0(n72), .A1(n73), .B0(n74), .Y(n71) );
  NOR2X4 U101 ( .A(n144), .B(n145), .Y(n141) );
  NAND2X2 U102 ( .A(n102), .B(n98), .Y(n132) );
  NAND2BX4 U103 ( .AN(B[14]), .B(A[14]), .Y(n98) );
  INVX8 U104 ( .A(n52), .Y(n61) );
  NAND2BX4 U105 ( .AN(B[6]), .B(A[6]), .Y(n52) );
  XOR2X4 U106 ( .A(n121), .B(n11), .Y(DIFF[15]) );
  OAI21X4 U107 ( .A0(n122), .A1(n123), .B0(n124), .Y(n121) );
  NAND2X4 U108 ( .A(n65), .B(n29), .Y(n54) );
  NAND4BX4 U109 ( .AN(n148), .B(n150), .C(n1), .D(n173), .Y(n114) );
  NOR2X4 U110 ( .A(n31), .B(n32), .Y(n30) );
  AOI21X4 U111 ( .A0(n15), .A1(n43), .B0(n65), .Y(n66) );
  INVX4 U112 ( .A(n149), .Y(n48) );
  XOR2X2 U113 ( .A(n15), .B(n67), .Y(DIFF[4]) );
  AOI21X2 U114 ( .A0(n15), .A1(n164), .B0(n172), .Y(n159) );
  NAND2X1 U115 ( .A(n170), .B(n43), .Y(n143) );
  CLKINVX4 U116 ( .A(n109), .Y(n95) );
  NAND2X2 U117 ( .A(n108), .B(n109), .Y(n136) );
  AND2X2 U118 ( .A(n109), .B(n99), .Y(n24) );
  NAND2X4 U119 ( .A(n61), .B(n42), .Y(n113) );
  AOI21X2 U120 ( .A0(n162), .A1(n16), .B0(n118), .Y(n161) );
  NAND2BX4 U121 ( .AN(A[4]), .B(B[4]), .Y(n43) );
  NAND2BX4 U122 ( .AN(B[4]), .B(A[4]), .Y(n69) );
  XOR2X2 U123 ( .A(n73), .B(n19), .Y(DIFF[2]) );
  NAND2BX4 U124 ( .AN(B[12]), .B(A[12]), .Y(n96) );
  NOR2X4 U125 ( .A(n75), .B(n78), .Y(n177) );
  NAND4BX2 U126 ( .AN(n175), .B(n29), .C(n1), .D(n15), .Y(n34) );
  INVX2 U127 ( .A(n43), .Y(n68) );
  NAND2X4 U128 ( .A(n12), .B(n141), .Y(n128) );
  NAND3X4 U129 ( .A(n27), .B(n140), .C(n128), .Y(n139) );
  NAND2X4 U130 ( .A(n18), .B(n157), .Y(n117) );
  AND2X4 U131 ( .A(n117), .B(n127), .Y(n27) );
  AND2X4 U132 ( .A(n117), .B(n127), .Y(n26) );
  AOI21X2 U133 ( .A0(n181), .A1(B[3]), .B0(n76), .Y(n56) );
  NOR2X2 U134 ( .A(n74), .B(n75), .Y(n19) );
  NAND2X2 U135 ( .A(n33), .B(n34), .Y(n37) );
  AND3X4 U136 ( .A(n140), .B(n128), .C(n25), .Y(n123) );
  NAND4BX2 U137 ( .AN(n100), .B(n102), .C(n108), .D(n109), .Y(n89) );
  NOR2X4 U138 ( .A(n31), .B(n35), .Y(n38) );
  XOR2X4 U139 ( .A(n60), .B(n20), .Y(DIFF[6]) );
  OAI21X4 U140 ( .A0(n95), .A1(n96), .B0(n99), .Y(n125) );
  XNOR2X4 U141 ( .A(n135), .B(n22), .Y(DIFF[12]) );
  XOR2X4 U142 ( .A(n23), .B(n66), .Y(DIFF[5]) );
  NAND2XL U143 ( .A(n29), .B(n55), .Y(n23) );
  XOR2X4 U144 ( .A(n137), .B(n24), .Y(DIFF[13]) );
  NOR2XL U145 ( .A(n100), .B(n101), .Y(n91) );
  AND2X1 U146 ( .A(n99), .B(n98), .Y(n97) );
  NAND2XL U147 ( .A(n82), .B(n83), .Y(DIFF[0]) );
  INVXL U148 ( .A(A[3]), .Y(n181) );
  AOI21X1 U149 ( .A0(n105), .A1(n106), .B0(n107), .Y(n86) );
  INVX1 U150 ( .A(n125), .Y(n134) );
  NAND3X4 U151 ( .A(n26), .B(n140), .C(n128), .Y(n135) );
  AOI21X1 U152 ( .A0(n125), .A1(n102), .B0(n126), .Y(n124) );
  XNOR2X4 U153 ( .A(n131), .B(n132), .Y(DIFF[14]) );
  INVXL U154 ( .A(n102), .Y(n101) );
  INVX1 U155 ( .A(n94), .Y(n93) );
  OAI21XL U156 ( .A0(n95), .A1(n96), .B0(n97), .Y(n92) );
  NAND2X2 U157 ( .A(n156), .B(n42), .Y(n145) );
  NAND2BXL U158 ( .AN(n89), .B(n156), .Y(n107) );
  NAND4BXL U159 ( .AN(n62), .B(n29), .C(n42), .D(n43), .Y(n104) );
  AOI21XL U160 ( .A0(n115), .A1(n58), .B0(n104), .Y(n111) );
  NOR2BX1 U161 ( .AN(n59), .B(n56), .Y(n115) );
  AND3X1 U162 ( .A(n153), .B(n8), .C(n170), .Y(n28) );
  NAND2BX4 U163 ( .AN(n83), .B(n82), .Y(n80) );
  NOR2XL U164 ( .A(n118), .B(n119), .Y(n116) );
  INVXL U165 ( .A(n120), .Y(n119) );
  INVXL U166 ( .A(A[9]), .Y(n169) );
  NAND2BX2 U167 ( .AN(A[12]), .B(B[12]), .Y(n108) );
  OAI2BB1X1 U168 ( .A0N(B[3]), .A1N(n181), .B0(n59), .Y(n70) );
  XOR2X1 U169 ( .A(B[16]), .B(A[16]), .Y(n85) );
  NAND2BX2 U170 ( .AN(B[9]), .B(A[9]), .Y(n36) );
  NOR2BX1 U171 ( .AN(B[8]), .B(A[8]), .Y(n152) );
  NAND2BX2 U172 ( .AN(A[7]), .B(B[7]), .Y(n42) );
  INVX8 U173 ( .A(n151), .Y(n129) );
  XOR2X4 U174 ( .A(n37), .B(n38), .Y(DIFF[8]) );
  XOR2X4 U175 ( .A(n45), .B(n46), .Y(DIFF[7]) );
  OAI21X4 U176 ( .A0(n50), .A1(n51), .B0(n52), .Y(n45) );
  AOI21X4 U177 ( .A0(n15), .A1(n43), .B0(n53), .Y(n50) );
  NAND2BX4 U178 ( .AN(n63), .B(n64), .Y(n60) );
  XOR2X4 U179 ( .A(n70), .B(n71), .Y(DIFF[3]) );
  CLKINVX3 U180 ( .A(n79), .Y(n81) );
  XOR2X4 U181 ( .A(n84), .B(n85), .Y(DIFF[16]) );
  NAND2X4 U182 ( .A(n133), .B(n134), .Y(n131) );
  NAND2X4 U183 ( .A(n138), .B(n96), .Y(n137) );
  NAND2X4 U184 ( .A(n139), .B(n108), .Y(n138) );
  NAND2X4 U185 ( .A(n129), .B(n130), .Y(n140) );
  NAND2BX4 U186 ( .AN(n146), .B(n147), .Y(n130) );
  OAI2BB1X4 U187 ( .A0N(n120), .A1N(n155), .B0(n156), .Y(n127) );
  XOR2X4 U188 ( .A(n158), .B(n3), .Y(DIFF[11]) );
  OAI21X4 U189 ( .A0(n159), .A1(n160), .B0(n161), .Y(n158) );
  XOR2X4 U190 ( .A(n167), .B(n2), .Y(DIFF[10]) );
  NAND2BX4 U191 ( .AN(A[10]), .B(B[10]), .Y(n112) );
  NAND2X4 U192 ( .A(n55), .B(n69), .Y(n150) );
  NAND2BX4 U193 ( .AN(B[5]), .B(A[5]), .Y(n55) );
  NAND2BX4 U194 ( .AN(A[6]), .B(B[6]), .Y(n40) );
  NAND4BX4 U195 ( .AN(n56), .B(n57), .C(n58), .D(n59), .Y(n41) );
  NAND3X4 U196 ( .A(n177), .B(n178), .C(n180), .Y(n58) );
  NAND2BX4 U197 ( .AN(B[1]), .B(A[1]), .Y(n79) );
  NAND2BX4 U198 ( .AN(A[1]), .B(B[1]), .Y(n179) );
  NAND2BX4 U199 ( .AN(A[2]), .B(B[2]), .Y(n72) );
  NAND2BX4 U200 ( .AN(A[0]), .B(B[0]), .Y(n83) );
endmodule


module butterfly_DW01_add_66 ( A, B, SUM );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  wire   n162, n163, n164, n165, n1, n2, n3, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n41,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161;

  CLKBUFX8 U2 ( .A(B[7]), .Y(n15) );
  OAI21X2 U3 ( .A0(n57), .A1(n2), .B0(n58), .Y(n54) );
  INVX1 U4 ( .A(n120), .Y(n122) );
  CLKINVX2 U5 ( .A(n33), .Y(n1) );
  INVX1 U6 ( .A(n1), .Y(n2) );
  INVX8 U7 ( .A(n102), .Y(n8) );
  NOR2BX2 U8 ( .AN(n3), .B(n27), .Y(n141) );
  NAND2X4 U9 ( .A(n147), .B(n53), .Y(n3) );
  INVX2 U10 ( .A(n59), .Y(n57) );
  BUFX3 U11 ( .A(n165), .Y(SUM[4]) );
  BUFX4 U12 ( .A(n164), .Y(SUM[5]) );
  INVX2 U13 ( .A(n66), .Y(n62) );
  INVX1 U14 ( .A(n94), .Y(n25) );
  OR2X2 U15 ( .A(A[4]), .B(B[4]), .Y(n72) );
  INVX1 U16 ( .A(n118), .Y(n123) );
  INVX2 U17 ( .A(n134), .Y(n56) );
  NAND2X1 U18 ( .A(B[0]), .B(A[0]), .Y(n88) );
  INVX1 U19 ( .A(n20), .Y(n21) );
  CLKINVX3 U20 ( .A(n44), .Y(n43) );
  XOR2X1 U21 ( .A(n70), .B(n71), .Y(n165) );
  NOR2BX1 U22 ( .AN(n69), .B(n67), .Y(n71) );
  XOR2X1 U23 ( .A(n64), .B(n65), .Y(n164) );
  XOR2X2 U24 ( .A(n73), .B(n74), .Y(SUM[3]) );
  INVX4 U25 ( .A(n39), .Y(SUM[6]) );
  CLKINVX3 U26 ( .A(n163), .Y(n39) );
  INVX1 U27 ( .A(n152), .Y(n9) );
  AND2X2 U28 ( .A(B[14]), .B(A[14]), .Y(n6) );
  AND2X4 U29 ( .A(n66), .B(n72), .Y(n7) );
  INVX4 U30 ( .A(n22), .Y(n138) );
  OAI21X1 U31 ( .A0(n110), .A1(n111), .B0(n112), .Y(n108) );
  INVX8 U32 ( .A(n101), .Y(n112) );
  NAND3X4 U33 ( .A(n70), .B(n112), .C(n138), .Y(n155) );
  NAND2X4 U34 ( .A(B[10]), .B(A[10]), .Y(n145) );
  OAI2BB1X4 U35 ( .A0N(n109), .A1N(n30), .B0(n8), .Y(n126) );
  OAI2BB1X4 U36 ( .A0N(n13), .A1N(n8), .B0(n125), .Y(n132) );
  XNOR2X4 U37 ( .A(n121), .B(n10), .Y(SUM[14]) );
  OR2X1 U38 ( .A(n99), .B(n6), .Y(n10) );
  BUFX2 U39 ( .A(n132), .Y(n17) );
  CLKINVX4 U40 ( .A(n125), .Y(n31) );
  NOR2BXL U41 ( .AN(n145), .B(n27), .Y(n152) );
  XNOR2X4 U42 ( .A(n150), .B(n9), .Y(SUM[10]) );
  INVX4 U43 ( .A(n64), .Y(n61) );
  XOR2X2 U44 ( .A(n59), .B(n60), .Y(n163) );
  AOI21X2 U45 ( .A0(n118), .A1(n18), .B0(n6), .Y(n117) );
  INVX2 U46 ( .A(n68), .Y(n29) );
  NAND2X2 U47 ( .A(n34), .B(A[4]), .Y(n69) );
  NOR2BX2 U48 ( .AN(n94), .B(n48), .Y(n115) );
  NAND3X2 U49 ( .A(n159), .B(n160), .C(n58), .Y(n12) );
  NAND2X4 U50 ( .A(n145), .B(n149), .Y(n32) );
  NAND2X4 U51 ( .A(n150), .B(n151), .Y(n149) );
  INVX2 U52 ( .A(n23), .Y(n11) );
  OR2X4 U53 ( .A(A[13]), .B(B[13]), .Y(n23) );
  BUFX3 U54 ( .A(n119), .Y(n18) );
  INVXL U55 ( .A(n113), .Y(n111) );
  INVXL U56 ( .A(n27), .Y(n151) );
  NOR2BX2 U57 ( .AN(n18), .B(n120), .Y(n116) );
  NOR2X2 U58 ( .A(n11), .B(n105), .Y(n103) );
  NAND2X4 U59 ( .A(A[9]), .B(B[9]), .Y(n147) );
  NAND2X4 U60 ( .A(n30), .B(n109), .Y(n13) );
  NAND3X4 U61 ( .A(n12), .B(n134), .C(n138), .Y(n154) );
  INVXL U62 ( .A(n139), .Y(n14) );
  BUFX3 U63 ( .A(n51), .Y(n16) );
  OR2XL U64 ( .A(B[9]), .B(A[9]), .Y(n137) );
  NOR2X4 U65 ( .A(A[9]), .B(B[9]), .Y(n148) );
  NAND2X1 U66 ( .A(A[5]), .B(B[5]), .Y(n161) );
  NOR2BX1 U67 ( .AN(n63), .B(n62), .Y(n65) );
  NAND2X1 U68 ( .A(n97), .B(n127), .Y(n131) );
  INVX1 U69 ( .A(n97), .Y(n19) );
  NOR2X4 U70 ( .A(n130), .B(n19), .Y(n129) );
  NAND2X1 U71 ( .A(B[5]), .B(A[5]), .Y(n63) );
  INVX1 U72 ( .A(n53), .Y(n20) );
  NOR2X4 U73 ( .A(n106), .B(n31), .Y(n91) );
  NOR2X4 U74 ( .A(A[8]), .B(B[8]), .Y(n22) );
  NAND2X2 U75 ( .A(n89), .B(n26), .Y(n36) );
  NAND2X2 U76 ( .A(B[3]), .B(A[3]), .Y(n75) );
  AOI2BB1X4 U77 ( .A0N(n93), .A1N(n48), .B0(n25), .Y(n24) );
  XNOR2X4 U78 ( .A(B[16]), .B(A[16]), .Y(n26) );
  NOR2X4 U79 ( .A(B[10]), .B(A[10]), .Y(n27) );
  BUFX8 U80 ( .A(n99), .Y(n28) );
  NOR2X2 U81 ( .A(n139), .B(n148), .Y(n140) );
  NAND2X4 U82 ( .A(n49), .B(n137), .Y(n153) );
  AOI2BB2X4 U83 ( .B0(n15), .B1(A[7]), .A0N(n33), .A1N(n161), .Y(n160) );
  NOR2BX2 U84 ( .AN(n51), .B(n148), .Y(n50) );
  NAND2X4 U85 ( .A(B[15]), .B(A[15]), .Y(n94) );
  XOR2X2 U86 ( .A(n13), .B(n52), .Y(SUM[8]) );
  NAND2X4 U87 ( .A(n29), .B(n112), .Y(n30) );
  INVX4 U88 ( .A(n70), .Y(n68) );
  NAND2X4 U89 ( .A(A[8]), .B(B[8]), .Y(n53) );
  XNOR2X4 U90 ( .A(n32), .B(n43), .Y(SUM[11]) );
  NAND2BX4 U91 ( .AN(n56), .B(n133), .Y(n109) );
  NAND2XL U92 ( .A(B[11]), .B(A[11]), .Y(n143) );
  NAND2X4 U93 ( .A(n98), .B(n97), .Y(n96) );
  NOR2X4 U94 ( .A(n48), .B(n28), .Y(n104) );
  NAND3BX4 U95 ( .AN(n69), .B(n156), .C(n66), .Y(n159) );
  INVX8 U96 ( .A(n146), .Y(n139) );
  NOR2X4 U97 ( .A(n139), .B(n145), .Y(n144) );
  NAND2X2 U98 ( .A(n127), .B(n23), .Y(n120) );
  INVX8 U99 ( .A(n107), .Y(n125) );
  NOR2BX4 U100 ( .AN(n143), .B(n144), .Y(n142) );
  NOR2X4 U101 ( .A(A[6]), .B(B[6]), .Y(n33) );
  BUFX8 U102 ( .A(B[4]), .Y(n34) );
  NAND2X4 U103 ( .A(n104), .B(n103), .Y(n92) );
  OAI21X4 U104 ( .A0(n97), .A1(n100), .B0(n98), .Y(n118) );
  NOR2X4 U105 ( .A(n148), .B(n22), .Y(n136) );
  AOI21X4 U106 ( .A0(n95), .A1(n96), .B0(n6), .Y(n93) );
  NAND3X4 U107 ( .A(n154), .B(n21), .C(n155), .Y(n49) );
  NOR2X4 U108 ( .A(n27), .B(n139), .Y(n135) );
  NOR2X4 U109 ( .A(n99), .B(n100), .Y(n95) );
  INVX8 U110 ( .A(n124), .Y(n100) );
  INVX8 U111 ( .A(n119), .Y(n99) );
  AOI21X2 U112 ( .A0(n108), .A1(n109), .B0(n102), .Y(n106) );
  NAND2X4 U113 ( .A(n135), .B(n136), .Y(n102) );
  NAND2X4 U114 ( .A(B[12]), .B(A[12]), .Y(n97) );
  NAND3X4 U115 ( .A(n7), .B(n46), .C(n156), .Y(n101) );
  NOR2X4 U116 ( .A(A[15]), .B(B[15]), .Y(n48) );
  XOR2X4 U117 ( .A(n54), .B(n55), .Y(SUM[7]) );
  XNOR2X4 U118 ( .A(n131), .B(n17), .Y(SUM[12]) );
  NAND2X4 U119 ( .A(n35), .B(n90), .Y(n37) );
  NAND2X4 U120 ( .A(n37), .B(n36), .Y(SUM[16]) );
  INVX4 U121 ( .A(n89), .Y(n35) );
  OAI21X4 U122 ( .A0(n91), .A1(n92), .B0(n24), .Y(n89) );
  XOR2X4 U123 ( .A(B[16]), .B(A[16]), .Y(n90) );
  NAND2X2 U124 ( .A(B[6]), .B(A[6]), .Y(n58) );
  AND2X4 U125 ( .A(n125), .B(n126), .Y(n38) );
  NOR2X4 U126 ( .A(n38), .B(n105), .Y(n130) );
  INVX4 U127 ( .A(n127), .Y(n105) );
  CLKINVX4 U128 ( .A(n162), .Y(n41) );
  INVX8 U129 ( .A(n41), .Y(SUM[9]) );
  NAND2X2 U130 ( .A(B[13]), .B(A[13]), .Y(n98) );
  OAI21X4 U131 ( .A0(n61), .A1(n62), .B0(n63), .Y(n59) );
  INVXL U132 ( .A(n82), .Y(n78) );
  OAI21X4 U133 ( .A0(n67), .A1(n68), .B0(n69), .Y(n64) );
  NOR2BXL U134 ( .AN(n58), .B(n2), .Y(n60) );
  AND2X1 U135 ( .A(n143), .B(n14), .Y(n44) );
  AND2X4 U136 ( .A(n82), .B(n158), .Y(n47) );
  NAND2X4 U137 ( .A(n47), .B(n157), .Y(n113) );
  OR2X4 U138 ( .A(A[7]), .B(B[7]), .Y(n46) );
  NOR2BX1 U139 ( .AN(n88), .B(n45), .Y(SUM[0]) );
  NOR2XL U140 ( .A(A[0]), .B(B[0]), .Y(n45) );
  OR2X4 U141 ( .A(A[3]), .B(B[3]), .Y(n158) );
  NOR2BX1 U142 ( .AN(n53), .B(n22), .Y(n52) );
  XOR2X1 U143 ( .A(n49), .B(n50), .Y(n162) );
  INVX1 U144 ( .A(n72), .Y(n67) );
  XOR2X1 U145 ( .A(n80), .B(n81), .Y(SUM[2]) );
  NOR2BX1 U146 ( .AN(n79), .B(n78), .Y(n81) );
  XOR2X1 U147 ( .A(n84), .B(n86), .Y(SUM[1]) );
  NOR2BXL U148 ( .AN(n85), .B(n87), .Y(n86) );
  OAI2BB1X1 U149 ( .A0N(n83), .A1N(n84), .B0(n85), .Y(n80) );
  INVX1 U150 ( .A(n88), .Y(n84) );
  AOI21XL U151 ( .A0(n15), .A1(A[7]), .B0(n56), .Y(n55) );
  NAND2X2 U152 ( .A(B[2]), .B(A[2]), .Y(n79) );
  NAND2X1 U153 ( .A(B[1]), .B(A[1]), .Y(n85) );
  INVXL U154 ( .A(n75), .Y(n110) );
  OR2X2 U155 ( .A(A[2]), .B(B[2]), .Y(n82) );
  OAI21XL U156 ( .A0(n77), .A1(n78), .B0(n79), .Y(n73) );
  NOR2BX1 U157 ( .AN(n75), .B(n76), .Y(n74) );
  INVX1 U158 ( .A(n80), .Y(n77) );
  NAND2XL U159 ( .A(A[9]), .B(B[9]), .Y(n51) );
  INVX1 U160 ( .A(n158), .Y(n76) );
  NAND2X4 U161 ( .A(n75), .B(n113), .Y(n70) );
  NAND2XL U162 ( .A(n23), .B(n98), .Y(n128) );
  XOR2X4 U163 ( .A(n114), .B(n115), .Y(SUM[15]) );
  OAI2BB1X4 U164 ( .A0N(n116), .A1N(n132), .B0(n117), .Y(n114) );
  OR2X4 U165 ( .A(B[14]), .B(A[14]), .Y(n119) );
  OAI2BB1X4 U166 ( .A0N(n122), .A1N(n132), .B0(n123), .Y(n121) );
  XOR2X4 U167 ( .A(n129), .B(n128), .Y(SUM[13]) );
  OR2X4 U168 ( .A(B[13]), .B(A[13]), .Y(n124) );
  OAI2BB1X4 U169 ( .A0N(n140), .A1N(n141), .B0(n142), .Y(n107) );
  OR2X4 U170 ( .A(A[12]), .B(B[12]), .Y(n127) );
  OR2X4 U171 ( .A(B[11]), .B(A[11]), .Y(n146) );
  NAND2X4 U172 ( .A(n153), .B(n16), .Y(n150) );
  OAI211X2 U173 ( .A0(n87), .A1(n88), .B0(n85), .C0(n79), .Y(n157) );
  CLKINVX3 U174 ( .A(n83), .Y(n87) );
  OR2X4 U175 ( .A(A[1]), .B(B[1]), .Y(n83) );
  NAND3X4 U176 ( .A(n159), .B(n160), .C(n58), .Y(n133) );
  OR2X4 U177 ( .A(B[6]), .B(A[6]), .Y(n156) );
  OR2X4 U178 ( .A(A[5]), .B(B[5]), .Y(n66) );
  OR2X4 U179 ( .A(A[7]), .B(B[7]), .Y(n134) );
endmodule


module butterfly_DW01_sub_74 ( A, B, DIFF );
  input [16:0] A;
  input [16:0] B;
  output [16:0] DIFF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181;

  AOI21X2 U3 ( .A0(n167), .A1(n157), .B0(n168), .Y(n166) );
  INVX1 U4 ( .A(B[2]), .Y(n179) );
  OAI21X4 U5 ( .A0(A[4]), .A1(n181), .B0(n59), .Y(n156) );
  INVX3 U6 ( .A(n17), .Y(n72) );
  NAND2BX4 U7 ( .AN(n124), .B(n123), .Y(n134) );
  BUFX20 U8 ( .A(B[5]), .Y(n39) );
  NAND2BX2 U9 ( .AN(B[2]), .B(A[2]), .Y(n177) );
  NOR2X4 U10 ( .A(n148), .B(n149), .Y(n158) );
  NAND2X4 U11 ( .A(n1), .B(B[9]), .Y(n48) );
  CLKINVX20 U12 ( .A(A[9]), .Y(n1) );
  OR2XL U13 ( .A(B[9]), .B(n24), .Y(n7) );
  NAND4BX1 U14 ( .AN(n120), .B(n4), .C(n62), .D(n14), .Y(n104) );
  NAND2BX2 U15 ( .AN(B[13]), .B(A[13]), .Y(n112) );
  INVX4 U16 ( .A(n69), .Y(n61) );
  CLKINVX8 U17 ( .A(A[4]), .Y(n37) );
  NAND2BX4 U18 ( .AN(A[4]), .B(B[4]), .Y(n62) );
  INVX1 U19 ( .A(A[7]), .Y(n15) );
  CLKINVX3 U20 ( .A(A[11]), .Y(n25) );
  CLKINVX4 U21 ( .A(n89), .Y(n84) );
  AOI21X1 U22 ( .A0(n113), .A1(n114), .B0(n102), .Y(n94) );
  NOR2X2 U23 ( .A(n68), .B(n61), .Y(n66) );
  INVX1 U24 ( .A(n169), .Y(n33) );
  NAND2X2 U25 ( .A(n178), .B(n89), .Y(n38) );
  AOI31X1 U26 ( .A0(n23), .A1(n4), .A2(n14), .B0(n138), .Y(n136) );
  INVX1 U27 ( .A(A[9]), .Y(n24) );
  BUFX3 U28 ( .A(n59), .Y(n4) );
  INVX1 U29 ( .A(A[6]), .Y(n5) );
  INVX1 U30 ( .A(A[8]), .Y(n13) );
  INVX1 U31 ( .A(n148), .Y(n20) );
  CLKINVX3 U32 ( .A(n62), .Y(n68) );
  OR2X2 U33 ( .A(B[4]), .B(n37), .Y(n16) );
  INVX1 U34 ( .A(n51), .Y(n47) );
  NOR2BX1 U35 ( .AN(n115), .B(n108), .Y(n150) );
  INVX1 U36 ( .A(n85), .Y(n88) );
  NOR2X2 U37 ( .A(n94), .B(n95), .Y(n92) );
  CLKINVX3 U38 ( .A(n46), .Y(n50) );
  AND2X4 U39 ( .A(n115), .B(n109), .Y(n2) );
  INVX1 U40 ( .A(n31), .Y(n27) );
  XOR2X4 U41 ( .A(n125), .B(n3), .Y(DIFF[15]) );
  NAND2X2 U42 ( .A(n98), .B(n107), .Y(n3) );
  NAND3X2 U43 ( .A(n80), .B(n105), .C(n119), .Y(n173) );
  INVX2 U44 ( .A(n63), .Y(n120) );
  NAND2X1 U45 ( .A(n14), .B(n6), .Y(n70) );
  NAND2BX2 U46 ( .AN(A[2]), .B(B[2]), .Y(n76) );
  OR2X4 U47 ( .A(B[6]), .B(n5), .Y(n57) );
  NAND2BX2 U48 ( .AN(A[13]), .B(B[13]), .Y(n109) );
  NAND2XL U49 ( .A(n46), .B(n48), .Y(n169) );
  CLKINVX4 U50 ( .A(n163), .Y(n11) );
  NOR2X1 U51 ( .A(n68), .B(n72), .Y(n73) );
  BUFX12 U52 ( .A(n131), .Y(n22) );
  NAND4BX4 U53 ( .AN(n50), .B(n11), .C(n10), .D(n157), .Y(n103) );
  CLKINVX4 U54 ( .A(n157), .Y(n160) );
  NAND2X2 U55 ( .A(n2), .B(n106), .Y(n132) );
  NOR2XL U56 ( .A(n104), .B(n105), .Y(n100) );
  NAND2X4 U57 ( .A(n5), .B(B[6]), .Y(n59) );
  NAND2X2 U58 ( .A(n121), .B(n64), .Y(n149) );
  NAND2BX1 U59 ( .AN(n39), .B(A[5]), .Y(n6) );
  AND2X2 U60 ( .A(n59), .B(n57), .Y(n26) );
  NAND2X2 U61 ( .A(n25), .B(B[11]), .Y(n153) );
  NAND2BX4 U62 ( .AN(A[1]), .B(B[1]), .Y(n89) );
  AOI21XL U63 ( .A0(n119), .A1(n80), .B0(n104), .Y(n117) );
  NAND2X4 U64 ( .A(n56), .B(n57), .Y(n55) );
  NAND4X4 U65 ( .A(n79), .B(n89), .C(n76), .D(n91), .Y(n105) );
  OAI21X4 U66 ( .A0(n39), .A1(n42), .B0(n17), .Y(n137) );
  INVXL U67 ( .A(n124), .Y(n8) );
  INVX2 U68 ( .A(n8), .Y(n9) );
  INVX1 U69 ( .A(A[14]), .Y(n21) );
  NAND2X2 U70 ( .A(n25), .B(B[11]), .Y(n10) );
  NAND2X2 U71 ( .A(n52), .B(n31), .Y(n29) );
  NAND2XL U72 ( .A(n11), .B(n49), .Y(n43) );
  NAND2X1 U73 ( .A(n157), .B(n48), .Y(n155) );
  OR2X4 U74 ( .A(B[9]), .B(n24), .Y(n49) );
  NAND2X4 U75 ( .A(n58), .B(n4), .Y(n56) );
  NAND3X4 U76 ( .A(n80), .B(n119), .C(n105), .Y(n12) );
  NAND2BX2 U77 ( .AN(B[15]), .B(A[15]), .Y(n98) );
  OR2X4 U78 ( .A(B[8]), .B(n13), .Y(n51) );
  NAND2BX4 U79 ( .AN(A[5]), .B(n39), .Y(n14) );
  OR2X4 U80 ( .A(B[7]), .B(n15), .Y(n64) );
  OR2X4 U81 ( .A(B[4]), .B(n37), .Y(n17) );
  NAND2BX2 U82 ( .AN(n151), .B(n22), .Y(n18) );
  XOR2X4 U83 ( .A(n144), .B(n19), .Y(DIFF[13]) );
  NAND2X1 U84 ( .A(n109), .B(n112), .Y(n19) );
  NAND2BX2 U85 ( .AN(B[12]), .B(A[12]), .Y(n143) );
  NAND2XL U86 ( .A(n111), .B(n112), .Y(n110) );
  AOI21X1 U87 ( .A0(n108), .A1(n109), .B0(n110), .Y(n96) );
  INVX3 U88 ( .A(n122), .Y(n148) );
  NAND2X2 U89 ( .A(n21), .B(B[14]), .Y(n106) );
  OR2X4 U90 ( .A(B[11]), .B(n25), .Y(n123) );
  AOI21X4 U91 ( .A0(n22), .A1(n130), .B0(n132), .Y(n126) );
  NAND2XL U92 ( .A(n62), .B(n59), .Y(n60) );
  NOR2X2 U93 ( .A(n120), .B(n136), .Y(n133) );
  OAI21XL U94 ( .A0(n39), .A1(n42), .B0(n17), .Y(n23) );
  CLKINVX3 U95 ( .A(A[5]), .Y(n42) );
  NAND4BX4 U96 ( .AN(n160), .B(n161), .C(n162), .D(n153), .Y(n135) );
  CLKINVX8 U97 ( .A(n48), .Y(n163) );
  NAND2X2 U98 ( .A(n14), .B(n63), .Y(n180) );
  AOI22X4 U99 ( .A0(B[5]), .A1(n42), .B0(n67), .B1(n16), .Y(n58) );
  XNOR2X4 U100 ( .A(n65), .B(n26), .Y(DIFF[6]) );
  XOR2X4 U101 ( .A(n92), .B(n93), .Y(DIFF[16]) );
  NAND2X2 U102 ( .A(n100), .B(n101), .Y(n99) );
  NAND2X4 U103 ( .A(n28), .B(n27), .Y(n30) );
  NAND2X4 U104 ( .A(n29), .B(n30), .Y(DIFF[7]) );
  INVX4 U105 ( .A(n52), .Y(n28) );
  AOI21X4 U106 ( .A0(n62), .A1(n53), .B0(n72), .Y(n71) );
  AND2X1 U107 ( .A(n63), .B(n64), .Y(n31) );
  NOR2X2 U108 ( .A(n60), .B(n61), .Y(n54) );
  NAND2BX4 U109 ( .AN(A[7]), .B(B[7]), .Y(n63) );
  NAND3BX4 U110 ( .AN(n169), .B(n157), .C(n32), .Y(n165) );
  AOI21X4 U111 ( .A0(n133), .A1(n118), .B0(n134), .Y(n130) );
  NAND3X4 U112 ( .A(n51), .B(n49), .C(n164), .Y(n161) );
  NAND2X2 U113 ( .A(n128), .B(n111), .Y(n127) );
  NAND2BX2 U114 ( .AN(B[14]), .B(A[14]), .Y(n111) );
  NAND2X2 U115 ( .A(n129), .B(n106), .Y(n128) );
  OAI2BB1X4 U116 ( .A0N(n172), .A1N(n173), .B0(n174), .Y(n32) );
  NOR2X4 U117 ( .A(n180), .B(n156), .Y(n172) );
  INVX4 U118 ( .A(n109), .Y(n142) );
  OAI21X4 U119 ( .A0(n83), .A1(n84), .B0(n85), .Y(n77) );
  NAND2BX4 U120 ( .AN(A[15]), .B(B[15]), .Y(n107) );
  OAI21X4 U121 ( .A0(n142), .A1(n143), .B0(n112), .Y(n129) );
  NOR2BX4 U122 ( .AN(n123), .B(n124), .Y(n159) );
  OAI21X4 U123 ( .A0(n158), .A1(n103), .B0(n159), .Y(n151) );
  NAND2X4 U124 ( .A(n163), .B(n164), .Y(n162) );
  OAI2BB1X4 U125 ( .A0N(n45), .A1N(n33), .B0(n171), .Y(n170) );
  XOR2X4 U126 ( .A(n34), .B(n35), .Y(DIFF[11]) );
  NAND2X4 U127 ( .A(n165), .B(n166), .Y(n34) );
  AND2X1 U128 ( .A(n10), .B(n123), .Y(n35) );
  NAND2BX4 U129 ( .AN(A[3]), .B(B[3]), .Y(n79) );
  NOR2BX4 U130 ( .AN(n121), .B(n36), .Y(n174) );
  NAND2X4 U131 ( .A(n122), .B(n64), .Y(n36) );
  OAI21X4 U132 ( .A0(n158), .A1(n103), .B0(n147), .Y(n146) );
  XOR2X2 U133 ( .A(n86), .B(n87), .Y(DIFF[1]) );
  OAI21X2 U134 ( .A0(A[2]), .A1(n179), .B0(n79), .Y(n175) );
  AOI21X4 U135 ( .A0(n45), .A1(n46), .B0(n47), .Y(n44) );
  NAND2BX2 U136 ( .AN(B[3]), .B(A[3]), .Y(n80) );
  INVX8 U137 ( .A(n143), .Y(n108) );
  NOR2BX4 U138 ( .AN(n123), .B(n124), .Y(n147) );
  XOR2X4 U139 ( .A(n44), .B(n43), .Y(DIFF[9]) );
  NAND2BX2 U140 ( .AN(A[12]), .B(B[12]), .Y(n115) );
  NAND3XL U141 ( .A(n121), .B(n64), .C(n20), .Y(n116) );
  NAND3X4 U142 ( .A(n38), .B(n85), .C(n177), .Y(n176) );
  XOR2X4 U143 ( .A(n140), .B(n139), .Y(DIFF[14]) );
  NAND2X4 U144 ( .A(n79), .B(n80), .Y(n74) );
  NAND4X2 U145 ( .A(n107), .B(n106), .C(n115), .D(n109), .Y(n102) );
  AOI21X4 U146 ( .A0(n141), .A1(n2), .B0(n129), .Y(n140) );
  AOI21X4 U147 ( .A0(n12), .A1(n54), .B0(n55), .Y(n52) );
  OAI21X1 U148 ( .A0(n116), .A1(n117), .B0(n118), .Y(n114) );
  INVX4 U149 ( .A(n103), .Y(n118) );
  NOR2X1 U150 ( .A(n102), .B(n103), .Y(n101) );
  NAND2X1 U151 ( .A(n64), .B(n57), .Y(n138) );
  NAND2XL U152 ( .A(n106), .B(n107), .Y(n97) );
  OAI211X2 U153 ( .A0(n96), .A1(n97), .B0(n98), .C0(n99), .Y(n95) );
  NAND2BX4 U154 ( .AN(B[1]), .B(A[1]), .Y(n85) );
  NAND2BX4 U155 ( .AN(n151), .B(n22), .Y(n141) );
  AOI21X4 U156 ( .A0(n66), .A1(n53), .B0(n58), .Y(n65) );
  OAI21X2 U157 ( .A0(n163), .A1(n51), .B0(n7), .Y(n167) );
  XOR2X4 U158 ( .A(n77), .B(n81), .Y(DIFF[2]) );
  NOR2BX2 U159 ( .AN(n177), .B(n82), .Y(n81) );
  XOR2X2 U160 ( .A(n12), .B(n73), .Y(DIFF[4]) );
  NAND2BX4 U161 ( .AN(A[8]), .B(B[8]), .Y(n46) );
  AOI21X2 U162 ( .A0(n76), .A1(n77), .B0(n78), .Y(n75) );
  INVX8 U163 ( .A(n135), .Y(n124) );
  NAND2BX4 U164 ( .AN(n39), .B(A[5]), .Y(n67) );
  NAND2BX4 U165 ( .AN(A[5]), .B(n39), .Y(n69) );
  NOR2X4 U166 ( .A(n126), .B(n127), .Y(n125) );
  NAND4X4 U167 ( .A(n137), .B(n69), .C(n59), .D(n63), .Y(n122) );
  NAND2BX4 U168 ( .AN(n57), .B(n63), .Y(n121) );
  NAND2BX2 U169 ( .AN(n91), .B(n90), .Y(n86) );
  NOR2X2 U170 ( .A(n88), .B(n84), .Y(n87) );
  XNOR2X4 U171 ( .A(n32), .B(n40), .Y(DIFF[8]) );
  OR2X4 U172 ( .A(n50), .B(n47), .Y(n40) );
  INVXL U173 ( .A(n177), .Y(n78) );
  NAND3XL U174 ( .A(n46), .B(n63), .C(n14), .Y(n152) );
  XOR2X4 U175 ( .A(n170), .B(n41), .Y(DIFF[10]) );
  AND2X1 U176 ( .A(n157), .B(n164), .Y(n41) );
  NAND2BXL U177 ( .AN(B[0]), .B(A[0]), .Y(n90) );
  INVX1 U178 ( .A(n167), .Y(n171) );
  NOR2X2 U179 ( .A(n155), .B(n156), .Y(n154) );
  NAND3X4 U180 ( .A(n80), .B(n119), .C(n105), .Y(n53) );
  INVX1 U181 ( .A(n86), .Y(n83) );
  XOR2X2 U182 ( .A(n74), .B(n75), .Y(DIFF[3]) );
  INVXL U183 ( .A(n164), .Y(n168) );
  INVX1 U184 ( .A(n76), .Y(n82) );
  NAND2X1 U185 ( .A(n106), .B(n111), .Y(n139) );
  NAND2XL U186 ( .A(n90), .B(n91), .Y(DIFF[0]) );
  INVX1 U187 ( .A(n90), .Y(n178) );
  INVXL U188 ( .A(B[4]), .Y(n181) );
  XOR2X1 U189 ( .A(B[16]), .B(A[16]), .Y(n93) );
  NOR2BXL U190 ( .AN(n123), .B(n9), .Y(n113) );
  NAND4BX2 U191 ( .AN(n152), .B(n10), .C(n154), .D(n12), .Y(n131) );
  XOR2X4 U192 ( .A(n70), .B(n71), .Y(DIFF[5]) );
  AOI21X4 U193 ( .A0(n145), .A1(n115), .B0(n108), .Y(n144) );
  NAND2BX4 U194 ( .AN(n146), .B(n22), .Y(n145) );
  XOR2X4 U195 ( .A(n18), .B(n150), .Y(DIFF[12]) );
  NAND2BX4 U196 ( .AN(B[10]), .B(A[10]), .Y(n164) );
  NAND2BX4 U197 ( .AN(A[10]), .B(B[10]), .Y(n157) );
  OAI2BB1X4 U198 ( .A0N(n172), .A1N(n173), .B0(n174), .Y(n45) );
  NAND2BX4 U199 ( .AN(n175), .B(n176), .Y(n119) );
  NAND2BX4 U200 ( .AN(A[0]), .B(B[0]), .Y(n91) );
endmodule


module butterfly_DW01_sub_76 ( A, B, DIFF );
  input [16:0] A;
  input [16:0] B;
  output [16:0] DIFF;
  wire   n171, n172, n173, n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n41, n42, n43,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170;

  INVX2 U3 ( .A(n104), .Y(n109) );
  CLKBUFX4 U4 ( .A(n19), .Y(n27) );
  NAND2BX4 U5 ( .AN(A[4]), .B(B[4]), .Y(n71) );
  INVX8 U6 ( .A(n61), .Y(n168) );
  CLKINVX8 U7 ( .A(n157), .Y(n38) );
  NAND4X4 U8 ( .A(n100), .B(n108), .C(n109), .D(n110), .Y(n96) );
  CLKINVX4 U9 ( .A(n101), .Y(n100) );
  INVX8 U10 ( .A(n153), .Y(n17) );
  AND2X4 U11 ( .A(n20), .B(n30), .Y(n60) );
  DLY1X1 U12 ( .A(n56), .Y(n30) );
  BUFX8 U13 ( .A(n112), .Y(n33) );
  NAND2X2 U14 ( .A(n112), .B(n58), .Y(n148) );
  NAND2X4 U15 ( .A(n70), .B(n71), .Y(n68) );
  NOR2XL U16 ( .A(n79), .B(n83), .Y(n82) );
  INVX2 U17 ( .A(n77), .Y(n83) );
  XOR2X2 U18 ( .A(n75), .B(n76), .Y(DIFF[3]) );
  AOI21XL U19 ( .A0(n77), .A1(n78), .B0(n79), .Y(n76) );
  INVX8 U20 ( .A(n69), .Y(n74) );
  NAND2BX4 U21 ( .AN(B[4]), .B(A[4]), .Y(n69) );
  NAND2BX4 U22 ( .AN(A[2]), .B(B[2]), .Y(n77) );
  NAND2BX2 U23 ( .AN(B[2]), .B(A[2]), .Y(n84) );
  BUFX4 U24 ( .A(n84), .Y(n1) );
  INVX4 U25 ( .A(n119), .Y(n127) );
  INVX1 U26 ( .A(n114), .Y(n35) );
  NAND2X2 U27 ( .A(n50), .B(n51), .Y(n151) );
  BUFX2 U28 ( .A(n28), .Y(n29) );
  NAND2BX1 U29 ( .AN(B[3]), .B(A[3]), .Y(n81) );
  OAI21XL U30 ( .A0(n85), .A1(n86), .B0(n87), .Y(n78) );
  NAND2BX2 U31 ( .AN(B[8]), .B(A[8]), .Y(n51) );
  CLKINVX3 U32 ( .A(n144), .Y(n49) );
  NAND2X1 U33 ( .A(n80), .B(n81), .Y(n75) );
  XOR2X2 U34 ( .A(n65), .B(n66), .Y(DIFF[5]) );
  NOR2BX1 U35 ( .AN(n64), .B(n63), .Y(n66) );
  INVX1 U36 ( .A(n168), .Y(n20) );
  CLKINVX3 U37 ( .A(n171), .Y(n43) );
  NAND2X4 U38 ( .A(n145), .B(n146), .Y(n132) );
  BUFX4 U39 ( .A(n113), .Y(n28) );
  XOR2X1 U40 ( .A(n46), .B(n47), .Y(n172) );
  NOR2X4 U41 ( .A(n148), .B(n104), .Y(n131) );
  AOI21X4 U42 ( .A0(n102), .A1(n103), .B0(n104), .Y(n98) );
  BUFX12 U43 ( .A(n172), .Y(DIFF[9]) );
  XNOR2X4 U44 ( .A(n42), .B(n149), .Y(n3) );
  AND2X4 U45 ( .A(n28), .B(n25), .Y(n4) );
  NAND2X2 U46 ( .A(n103), .B(n146), .Y(n53) );
  NAND2BX2 U47 ( .AN(n105), .B(n70), .Y(n146) );
  NAND2BX4 U48 ( .AN(n24), .B(n106), .Y(n102) );
  INVX4 U49 ( .A(A[11]), .Y(n5) );
  NOR2BX4 U50 ( .AN(n80), .B(n83), .Y(n164) );
  NAND2BX4 U51 ( .AN(n152), .B(n154), .Y(n13) );
  NOR2BX4 U52 ( .AN(A[9]), .B(B[9]), .Y(n141) );
  NAND2X4 U53 ( .A(n5), .B(B[11]), .Y(n142) );
  NAND2X4 U54 ( .A(n6), .B(A[13]), .Y(n128) );
  INVX4 U55 ( .A(B[13]), .Y(n6) );
  OAI211X2 U56 ( .A0(n136), .A1(n137), .B0(n138), .C0(n139), .Y(n134) );
  NAND2BX2 U57 ( .AN(B[15]), .B(A[15]), .Y(n123) );
  BUFX3 U58 ( .A(n114), .Y(n7) );
  BUFX1 U59 ( .A(n144), .Y(n8) );
  INVXL U60 ( .A(n121), .Y(n22) );
  INVXL U61 ( .A(n120), .Y(n9) );
  CLKINVX1 U62 ( .A(n17), .Y(n12) );
  INVX4 U63 ( .A(n12), .Y(n152) );
  INVX3 U64 ( .A(n25), .Y(n118) );
  CLKBUFX8 U65 ( .A(n120), .Y(n10) );
  XOR2X2 U66 ( .A(n126), .B(n41), .Y(n11) );
  CLKINVX20 U67 ( .A(n11), .Y(DIFF[13]) );
  NAND2BX4 U68 ( .AN(B[9]), .B(A[9]), .Y(n50) );
  AOI21X4 U69 ( .A0(n30), .A1(n57), .B0(n168), .Y(n55) );
  NAND2X2 U70 ( .A(n126), .B(n29), .Y(n130) );
  NAND4X4 U71 ( .A(n113), .B(n114), .C(n111), .D(n33), .Y(n101) );
  XOR2X4 U72 ( .A(n13), .B(n14), .Y(DIFF[11]) );
  AND2X1 U73 ( .A(n27), .B(n139), .Y(n14) );
  NOR2X4 U74 ( .A(n48), .B(n49), .Y(n47) );
  CLKINVX3 U75 ( .A(A[10]), .Y(n15) );
  CLKINVX4 U76 ( .A(n15), .Y(n16) );
  NAND4BX4 U77 ( .AN(n49), .B(n151), .C(n27), .D(n38), .Y(n150) );
  CLKINVX3 U78 ( .A(n143), .Y(n157) );
  INVXL U79 ( .A(n121), .Y(n18) );
  INVX8 U80 ( .A(n135), .Y(n120) );
  NAND2X4 U81 ( .A(n1), .B(n87), .Y(n163) );
  NAND2BX2 U82 ( .AN(B[1]), .B(A[1]), .Y(n87) );
  NAND2BX4 U83 ( .AN(A[11]), .B(B[11]), .Y(n19) );
  INVX1 U84 ( .A(n147), .Y(n145) );
  NAND2X2 U85 ( .A(n147), .B(n58), .Y(n103) );
  NAND3X4 U86 ( .A(n147), .B(n58), .C(n52), .Y(n159) );
  NAND2BX4 U87 ( .AN(B[11]), .B(n37), .Y(n139) );
  XOR2X1 U88 ( .A(n155), .B(n156), .Y(n171) );
  XNOR2X4 U89 ( .A(n129), .B(n21), .Y(DIFF[14]) );
  OR2X4 U90 ( .A(n118), .B(n127), .Y(n21) );
  AND2X2 U91 ( .A(n138), .B(n139), .Y(n32) );
  INVX4 U92 ( .A(n123), .Y(n116) );
  AOI2BB1X4 U93 ( .A0N(n22), .A1N(n118), .B0(n127), .Y(n124) );
  INVXL U94 ( .A(n121), .Y(n23) );
  INVX8 U95 ( .A(n128), .Y(n121) );
  INVXL U96 ( .A(n108), .Y(n24) );
  NAND2BX4 U97 ( .AN(A[14]), .B(B[14]), .Y(n25) );
  INVX8 U98 ( .A(n3), .Y(DIFF[12]) );
  NAND2X1 U99 ( .A(n28), .B(n18), .Y(n41) );
  BUFX8 U100 ( .A(A[12]), .Y(n34) );
  NAND2X4 U101 ( .A(n126), .B(n4), .Y(n125) );
  XNOR2X4 U102 ( .A(n94), .B(n31), .Y(DIFF[16]) );
  XOR2X4 U103 ( .A(B[16]), .B(A[16]), .Y(n31) );
  OR2X4 U104 ( .A(n35), .B(n116), .Y(n36) );
  NAND2X4 U105 ( .A(n130), .B(n23), .Y(n129) );
  NAND2X4 U106 ( .A(n46), .B(n8), .Y(n158) );
  NAND2BX2 U107 ( .AN(A[7]), .B(B[7]), .Y(n58) );
  NAND2BX2 U108 ( .AN(B[7]), .B(A[7]), .Y(n59) );
  NAND3BX4 U109 ( .AN(B[5]), .B(n56), .C(A[5]), .Y(n169) );
  NAND3X4 U110 ( .A(n56), .B(n67), .C(n74), .Y(n170) );
  NAND3X4 U111 ( .A(n70), .B(n108), .C(n52), .Y(n160) );
  INVX2 U112 ( .A(n50), .Y(n48) );
  NAND2X4 U113 ( .A(n150), .B(n32), .Y(n99) );
  CLKINVX8 U114 ( .A(n105), .Y(n108) );
  NAND2BX4 U115 ( .AN(n117), .B(n25), .Y(n39) );
  NAND2X4 U116 ( .A(n68), .B(n69), .Y(n65) );
  NAND2X4 U117 ( .A(n155), .B(n38), .Y(n154) );
  NAND2BX4 U118 ( .AN(B[14]), .B(A[14]), .Y(n119) );
  BUFX16 U119 ( .A(n173), .Y(DIFF[7]) );
  XOR2X4 U120 ( .A(n55), .B(n54), .Y(n173) );
  INVX4 U121 ( .A(n65), .Y(n62) );
  NAND3X4 U122 ( .A(n159), .B(n160), .C(n51), .Y(n46) );
  XOR2X4 U123 ( .A(n57), .B(n60), .Y(DIFF[6]) );
  NOR2BX4 U124 ( .AN(B[7]), .B(A[7]), .Y(n161) );
  NAND2X4 U125 ( .A(n17), .B(n19), .Y(n138) );
  INVX4 U126 ( .A(n91), .Y(n86) );
  INVX8 U127 ( .A(n43), .Y(DIFF[10]) );
  XNOR2X4 U128 ( .A(n122), .B(n36), .Y(DIFF[15]) );
  NAND2X4 U129 ( .A(n125), .B(n124), .Y(n122) );
  AOI21X4 U130 ( .A0(n120), .A1(n113), .B0(n121), .Y(n117) );
  OAI21X4 U131 ( .A0(n162), .A1(n163), .B0(n164), .Y(n107) );
  AOI21X2 U132 ( .A0(n165), .A1(B[1]), .B0(n92), .Y(n162) );
  OAI21X4 U133 ( .A0(n98), .A1(n99), .B0(n100), .Y(n97) );
  INVX2 U134 ( .A(n5), .Y(n37) );
  AOI21X4 U135 ( .A0(n33), .A1(n134), .B0(n10), .Y(n133) );
  AOI21X4 U136 ( .A0(n115), .A1(n7), .B0(n116), .Y(n95) );
  NAND2X1 U137 ( .A(n81), .B(n107), .Y(n106) );
  XOR2X2 U138 ( .A(n70), .B(n72), .Y(DIFF[4]) );
  NAND2X2 U139 ( .A(n80), .B(n91), .Y(n167) );
  NAND2BX4 U140 ( .AN(A[3]), .B(B[3]), .Y(n80) );
  NAND2X4 U141 ( .A(n158), .B(n50), .Y(n155) );
  NAND2BX4 U142 ( .AN(B[6]), .B(A[6]), .Y(n61) );
  OAI21X4 U143 ( .A0(n140), .A1(n141), .B0(n142), .Y(n137) );
  NAND3X4 U144 ( .A(n95), .B(n96), .C(n97), .Y(n94) );
  NAND2X4 U145 ( .A(n39), .B(n119), .Y(n115) );
  NAND2X4 U146 ( .A(n144), .B(n143), .Y(n136) );
  NAND4BX4 U147 ( .AN(n161), .B(n56), .C(n67), .D(n71), .Y(n105) );
  NOR2BX2 U148 ( .AN(A[8]), .B(B[8]), .Y(n140) );
  NAND4X4 U149 ( .A(n19), .B(n143), .C(n144), .D(n52), .Y(n104) );
  NAND2BX4 U150 ( .AN(A[13]), .B(B[13]), .Y(n113) );
  NAND4BX4 U151 ( .AN(n168), .B(n169), .C(n59), .D(n170), .Y(n147) );
  OAI21X4 U152 ( .A0(n62), .A1(n63), .B0(n64), .Y(n57) );
  XOR2X4 U153 ( .A(n53), .B(n45), .Y(DIFF[8]) );
  NAND2BX2 U154 ( .AN(A[1]), .B(B[1]), .Y(n91) );
  NOR2XL U155 ( .A(n157), .B(n152), .Y(n156) );
  NAND2X1 U156 ( .A(n77), .B(n93), .Y(n166) );
  NAND3BX4 U157 ( .AN(n110), .B(n81), .C(n107), .Y(n70) );
  AND2X1 U158 ( .A(n51), .B(n52), .Y(n45) );
  NAND2XL U159 ( .A(n33), .B(n9), .Y(n42) );
  NOR2XL U160 ( .A(n90), .B(n86), .Y(n89) );
  INVXL U161 ( .A(n87), .Y(n90) );
  INVXL U162 ( .A(n1), .Y(n79) );
  NAND2BXL U163 ( .AN(n93), .B(n92), .Y(n88) );
  NAND2XL U164 ( .A(n92), .B(n93), .Y(DIFF[0]) );
  XOR2X1 U165 ( .A(n78), .B(n82), .Y(DIFF[2]) );
  NAND2X1 U166 ( .A(n58), .B(n59), .Y(n54) );
  NOR2X1 U167 ( .A(n73), .B(n74), .Y(n72) );
  INVX1 U168 ( .A(n71), .Y(n73) );
  XOR2X1 U169 ( .A(n88), .B(n89), .Y(DIFF[1]) );
  INVX1 U170 ( .A(n88), .Y(n85) );
  NAND2BXL U171 ( .AN(B[5]), .B(A[5]), .Y(n64) );
  INVX1 U172 ( .A(A[1]), .Y(n165) );
  NAND2BX1 U173 ( .AN(B[0]), .B(A[0]), .Y(n92) );
  NAND2BX1 U174 ( .AN(A[0]), .B(B[0]), .Y(n93) );
  CLKINVX3 U175 ( .A(n67), .Y(n63) );
  NAND2BX4 U176 ( .AN(A[15]), .B(B[15]), .Y(n114) );
  NAND2BX4 U177 ( .AN(A[14]), .B(B[14]), .Y(n111) );
  OAI2BB1X4 U178 ( .A0N(n131), .A1N(n132), .B0(n133), .Y(n126) );
  AOI21X4 U179 ( .A0(n53), .A1(n109), .B0(n99), .Y(n149) );
  NAND2BX4 U180 ( .AN(A[12]), .B(B[12]), .Y(n112) );
  NAND2BX4 U181 ( .AN(B[12]), .B(n34), .Y(n135) );
  NAND2BX4 U182 ( .AN(B[10]), .B(n16), .Y(n153) );
  NAND2BX4 U183 ( .AN(A[10]), .B(B[10]), .Y(n143) );
  NAND2BX4 U184 ( .AN(A[9]), .B(B[9]), .Y(n144) );
  NOR2X4 U185 ( .A(n166), .B(n167), .Y(n110) );
  NAND2BX4 U186 ( .AN(A[5]), .B(B[5]), .Y(n67) );
  NAND2BX4 U187 ( .AN(A[6]), .B(B[6]), .Y(n56) );
  NAND2BX4 U188 ( .AN(A[8]), .B(B[8]), .Y(n52) );
endmodule


module butterfly_DW01_sub_78 ( A, B, DIFF );
  input [16:0] A;
  input [16:0] B;
  output [16:0] DIFF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218;

  INVX4 U3 ( .A(n196), .Y(n36) );
  CLKINVX3 U4 ( .A(n37), .Y(n38) );
  AND2X2 U5 ( .A(n83), .B(n62), .Y(n17) );
  INVX4 U6 ( .A(n83), .Y(n100) );
  BUFX1 U7 ( .A(A[1]), .Y(n18) );
  INVX4 U8 ( .A(A[1]), .Y(n56) );
  NAND2BXL U9 ( .AN(B[1]), .B(A[1]), .Y(n116) );
  NAND2BX1 U10 ( .AN(A[9]), .B(B[9]), .Y(n183) );
  OAI21X4 U11 ( .A0(n123), .A1(n124), .B0(n125), .Y(n121) );
  NAND4X4 U12 ( .A(n132), .B(n4), .C(n142), .D(n143), .Y(n124) );
  OAI21X2 U13 ( .A0(n115), .A1(n16), .B0(n116), .Y(n109) );
  AND2X4 U14 ( .A(n82), .B(n83), .Y(n58) );
  NAND2X4 U15 ( .A(n157), .B(n156), .Y(n155) );
  NAND2X4 U16 ( .A(n41), .B(n185), .Y(n156) );
  NAND2X4 U17 ( .A(n5), .B(B[4]), .Y(n77) );
  AND2X4 U18 ( .A(n40), .B(n55), .Y(n1) );
  NAND2X2 U19 ( .A(n195), .B(n71), .Y(n191) );
  NAND3X4 U20 ( .A(n20), .B(n77), .C(n54), .Y(n95) );
  BUFX2 U21 ( .A(n111), .Y(n2) );
  NAND4BX4 U22 ( .AN(n31), .B(n62), .C(A[4]), .D(n212), .Y(n211) );
  CLKINVX4 U23 ( .A(B[4]), .Y(n35) );
  OAI21X1 U24 ( .A0(n135), .A1(n136), .B0(n137), .Y(n134) );
  INVX8 U25 ( .A(n143), .Y(n135) );
  AND2X4 U26 ( .A(n130), .B(n132), .Y(n24) );
  NAND2X4 U27 ( .A(n142), .B(n174), .Y(n163) );
  NAND2BX2 U28 ( .AN(n9), .B(n3), .Y(n10) );
  INVX4 U29 ( .A(n91), .Y(n43) );
  INVX1 U30 ( .A(B[1]), .Y(n8) );
  BUFX12 U31 ( .A(n103), .Y(n54) );
  INVX1 U32 ( .A(n120), .Y(n9) );
  BUFX4 U33 ( .A(n66), .Y(n26) );
  CLKINVX3 U34 ( .A(n163), .Y(n25) );
  INVX1 U35 ( .A(n49), .Y(n48) );
  CLKINVX3 U36 ( .A(n169), .Y(n28) );
  CLKINVX3 U37 ( .A(n136), .Y(n169) );
  CLKINVX3 U38 ( .A(n195), .Y(n69) );
  AND2X2 U39 ( .A(n61), .B(n78), .Y(n13) );
  CLKBUFX8 U40 ( .A(n77), .Y(n61) );
  NAND2BX1 U41 ( .AN(A[0]), .B(B[0]), .Y(n120) );
  XOR2X2 U42 ( .A(n117), .B(n118), .Y(DIFF[1]) );
  NAND2X1 U43 ( .A(n54), .B(n2), .Y(n106) );
  INVX3 U44 ( .A(n104), .Y(n39) );
  NAND3X2 U45 ( .A(n98), .B(n97), .C(n96), .Y(n94) );
  CLKINVX8 U46 ( .A(n113), .Y(n30) );
  INVX4 U47 ( .A(n108), .Y(n113) );
  NAND2X4 U48 ( .A(n56), .B(B[1]), .Y(n3) );
  NAND2BX2 U49 ( .AN(B[2]), .B(A[2]), .Y(n114) );
  CLKINVX3 U50 ( .A(n71), .Y(n88) );
  NAND3X4 U51 ( .A(n62), .B(n26), .C(n7), .Y(n53) );
  NAND3X4 U52 ( .A(n60), .B(n218), .C(n217), .Y(n20) );
  NAND2X4 U53 ( .A(n66), .B(n63), .Y(n96) );
  INVX8 U54 ( .A(n64), .Y(n63) );
  BUFX8 U55 ( .A(n131), .Y(n4) );
  INVX2 U56 ( .A(n35), .Y(n31) );
  NAND2BX4 U57 ( .AN(n63), .B(n65), .Y(n212) );
  OAI2BB1X2 U58 ( .A0N(n65), .A1N(n64), .B0(n62), .Y(n93) );
  AOI21X4 U59 ( .A0(n156), .A1(n181), .B0(n182), .Y(n180) );
  INVX4 U60 ( .A(A[4]), .Y(n5) );
  NAND2BX4 U61 ( .AN(B[3]), .B(A[3]), .Y(n111) );
  XOR2X4 U62 ( .A(n179), .B(n6), .Y(DIFF[12]) );
  NAND2XL U63 ( .A(n142), .B(n136), .Y(n6) );
  AND2X4 U64 ( .A(n96), .B(n102), .Y(n46) );
  NAND4BX1 U65 ( .AN(n31), .B(n62), .C(n212), .D(A[4]), .Y(n178) );
  NAND2X4 U66 ( .A(n35), .B(A[4]), .Y(n97) );
  INVX8 U67 ( .A(n141), .Y(n104) );
  INVX8 U68 ( .A(n64), .Y(n7) );
  NOR2X2 U69 ( .A(n79), .B(n188), .Y(n181) );
  NAND3X4 U70 ( .A(n8), .B(n108), .C(n18), .Y(n218) );
  CLKINVX4 U71 ( .A(n89), .Y(n47) );
  NAND3X4 U72 ( .A(n82), .B(n29), .C(n53), .Y(n80) );
  NAND2BX4 U73 ( .AN(B[8]), .B(A[8]), .Y(n71) );
  INVXL U74 ( .A(n55), .Y(n87) );
  BUFX20 U75 ( .A(n76), .Y(n55) );
  AND4X4 U76 ( .A(n15), .B(n47), .C(n48), .D(n140), .Y(n126) );
  NOR2X1 U77 ( .A(n110), .B(n113), .Y(n112) );
  INVX3 U78 ( .A(n114), .Y(n110) );
  NAND3X4 U79 ( .A(n217), .B(n60), .C(n218), .Y(n27) );
  NAND2BX1 U80 ( .AN(B[13]), .B(A[13]), .Y(n137) );
  NAND2BX2 U81 ( .AN(A[7]), .B(B[7]), .Y(n91) );
  NAND3X4 U82 ( .A(n11), .B(n54), .C(n30), .Y(n141) );
  INVX4 U83 ( .A(n10), .Y(n11) );
  NAND2BX4 U84 ( .AN(B[9]), .B(A[9]), .Y(n195) );
  NAND3X4 U85 ( .A(n1), .B(n36), .C(n174), .Y(n146) );
  INVX4 U86 ( .A(n62), .Y(n51) );
  NAND2X4 U87 ( .A(n41), .B(n213), .Y(n205) );
  XOR2X4 U88 ( .A(n50), .B(n12), .Y(DIFF[11]) );
  AND2X1 U89 ( .A(n194), .B(n174), .Y(n12) );
  NAND4X4 U90 ( .A(n13), .B(n14), .C(n62), .D(n41), .Y(n73) );
  AND2X4 U91 ( .A(n44), .B(n55), .Y(n14) );
  NAND3BX4 U92 ( .AN(n88), .B(n72), .C(n73), .Y(n67) );
  INVXL U93 ( .A(n39), .Y(n15) );
  AND2X4 U94 ( .A(n56), .B(B[1]), .Y(n16) );
  NAND2X4 U95 ( .A(n27), .B(n54), .Y(n216) );
  XOR2X4 U96 ( .A(n99), .B(n17), .Y(DIFF[6]) );
  AND2X2 U97 ( .A(n116), .B(n3), .Y(n118) );
  NOR2X4 U98 ( .A(n49), .B(n158), .Y(n153) );
  AOI2BB1X4 U99 ( .A0N(n200), .A1N(n71), .B0(n203), .Y(n197) );
  NAND2BX2 U100 ( .AN(B[14]), .B(A[14]), .Y(n138) );
  AND3X4 U101 ( .A(n27), .B(n77), .C(n54), .Y(n19) );
  AND2X2 U102 ( .A(n22), .B(n25), .Y(n159) );
  INVX4 U103 ( .A(n22), .Y(n162) );
  NAND4BBX4 U104 ( .AN(n89), .BN(n200), .C(n55), .D(n41), .Y(n199) );
  NAND2BX1 U105 ( .AN(n193), .B(n36), .Y(n45) );
  AND2X2 U106 ( .A(n194), .B(n204), .Y(n21) );
  NAND2X1 U107 ( .A(n62), .B(n77), .Y(n187) );
  NAND3X4 U108 ( .A(n166), .B(n165), .C(n164), .Y(n33) );
  OAI2BB1X4 U109 ( .A0N(n190), .A1N(n191), .B0(n21), .Y(n22) );
  AOI21X4 U110 ( .A0(n159), .A1(n154), .B0(n160), .Y(n149) );
  OAI21X4 U111 ( .A0(n79), .A1(n80), .B0(n81), .Y(n72) );
  INVX3 U112 ( .A(n189), .Y(n79) );
  XOR2X4 U113 ( .A(n23), .B(n24), .Y(DIFF[15]) );
  NAND3X4 U114 ( .A(n149), .B(n150), .C(n151), .Y(n23) );
  AOI2BB1X2 U115 ( .A0N(n28), .A1N(n135), .B0(n152), .Y(n164) );
  BUFX4 U116 ( .A(n101), .Y(n32) );
  NAND3X1 U117 ( .A(n25), .B(n143), .C(n168), .Y(n165) );
  AND2X4 U118 ( .A(n194), .B(n204), .Y(n192) );
  CLKINVX4 U119 ( .A(n204), .Y(n193) );
  NAND2BX4 U120 ( .AN(B[10]), .B(A[10]), .Y(n204) );
  AOI21X4 U121 ( .A0(n175), .A1(n156), .B0(n176), .Y(n172) );
  NAND3X2 U122 ( .A(n78), .B(n44), .C(n183), .Y(n215) );
  CLKINVX8 U123 ( .A(n100), .Y(n29) );
  NAND3BX4 U124 ( .AN(n49), .B(n155), .C(n167), .Y(n166) );
  NOR2X1 U125 ( .A(n135), .B(n158), .Y(n167) );
  NAND2X2 U126 ( .A(n82), .B(n83), .Y(n210) );
  NAND2BX4 U127 ( .AN(A[3]), .B(B[3]), .Y(n103) );
  NAND2BX2 U128 ( .AN(B[12]), .B(A[12]), .Y(n136) );
  NAND2X2 U129 ( .A(n184), .B(n40), .Y(n200) );
  XOR2X4 U130 ( .A(n33), .B(n34), .Y(DIFF[14]) );
  AND2X1 U131 ( .A(n131), .B(n138), .Y(n34) );
  OR2X2 U132 ( .A(A[5]), .B(n66), .Y(n102) );
  NAND4X4 U133 ( .A(n35), .B(n62), .C(A[4]), .D(n201), .Y(n189) );
  INVX8 U134 ( .A(A[5]), .Y(n64) );
  NAND2X2 U135 ( .A(n177), .B(n44), .Y(n175) );
  INVX8 U136 ( .A(n139), .Y(n49) );
  CLKINVX2 U137 ( .A(A[6]), .Y(n37) );
  NOR2X2 U138 ( .A(n144), .B(n42), .Y(n123) );
  CLKBUFXL U139 ( .A(n59), .Y(n42) );
  NAND2BX4 U140 ( .AN(A[9]), .B(B[9]), .Y(n40) );
  NAND2X4 U141 ( .A(n147), .B(n44), .Y(n157) );
  INVX8 U142 ( .A(n146), .Y(n139) );
  BUFX20 U143 ( .A(n75), .Y(n41) );
  NAND3BX1 U144 ( .AN(n148), .B(n20), .C(n47), .Y(n145) );
  OAI21X2 U145 ( .A0(n28), .A1(n161), .B0(n138), .Y(n160) );
  NAND2XL U146 ( .A(n88), .B(n40), .Y(n206) );
  INVX8 U147 ( .A(n43), .Y(n44) );
  NAND2X4 U148 ( .A(n139), .B(n44), .Y(n182) );
  INVX2 U149 ( .A(n137), .Y(n152) );
  NOR2X2 U150 ( .A(n69), .B(n70), .Y(n68) );
  NAND3BX2 U151 ( .AN(n200), .B(n147), .C(n81), .Y(n198) );
  XNOR2X4 U152 ( .A(n52), .B(n45), .Y(DIFF[10]) );
  OAI21X2 U153 ( .A0(n128), .A1(n129), .B0(n130), .Y(n127) );
  XOR2X4 U154 ( .A(n32), .B(n46), .Y(DIFF[5]) );
  NOR2X4 U155 ( .A(n70), .B(n202), .Y(n208) );
  NOR2X4 U156 ( .A(n214), .B(n215), .Y(n213) );
  NAND2X4 U157 ( .A(n143), .B(n131), .Y(n161) );
  OAI2BB1X4 U158 ( .A0N(n41), .A1N(n47), .B0(n157), .Y(n85) );
  AND2X2 U159 ( .A(n82), .B(n44), .Y(n57) );
  INVX4 U160 ( .A(n142), .Y(n158) );
  NAND2BX4 U161 ( .AN(A[6]), .B(B[6]), .Y(n74) );
  INVX8 U162 ( .A(n184), .Y(n196) );
  NAND2X2 U163 ( .A(n44), .B(n78), .Y(n186) );
  NAND4BX4 U164 ( .AN(n51), .B(n61), .C(n44), .D(n78), .Y(n89) );
  INVX4 U165 ( .A(n161), .Y(n154) );
  NAND3X4 U166 ( .A(n198), .B(n199), .C(n197), .Y(n50) );
  OAI2BB1X4 U167 ( .A0N(n102), .A1N(n101), .B0(n96), .Y(n99) );
  OAI21X4 U168 ( .A0(n92), .A1(n93), .B0(n29), .Y(n90) );
  NOR2X4 U169 ( .A(n94), .B(n19), .Y(n92) );
  NAND3X2 U170 ( .A(n155), .B(n154), .C(n153), .Y(n150) );
  NOR2X4 U171 ( .A(n70), .B(n196), .Y(n190) );
  BUFX20 U172 ( .A(n74), .Y(n62) );
  AOI21X4 U173 ( .A0(n208), .A1(n209), .B0(n69), .Y(n207) );
  NAND3BX4 U174 ( .AN(n119), .B(n108), .C(n3), .Y(n217) );
  NAND2BX4 U175 ( .AN(A[2]), .B(B[2]), .Y(n108) );
  NAND3X4 U176 ( .A(n207), .B(n206), .C(n205), .Y(n52) );
  NAND3X4 U177 ( .A(n95), .B(n98), .C(n97), .Y(n101) );
  XOR2X4 U178 ( .A(n107), .B(n106), .Y(DIFF[3]) );
  AOI21X2 U179 ( .A0(n30), .A1(n109), .B0(n110), .Y(n107) );
  NAND2BX1 U180 ( .AN(B[15]), .B(A[15]), .Y(n130) );
  OAI21X2 U181 ( .A0(n195), .A1(n196), .B0(n204), .Y(n203) );
  NOR2X4 U182 ( .A(n186), .B(n187), .Y(n185) );
  NAND4BX4 U183 ( .AN(n100), .B(n189), .C(n84), .D(n82), .Y(n147) );
  INVX4 U184 ( .A(n202), .Y(n81) );
  NAND3BX4 U185 ( .AN(n210), .B(n211), .C(n84), .Y(n209) );
  XOR2X4 U186 ( .A(n121), .B(n122), .Y(DIFF[16]) );
  NAND3X2 U187 ( .A(n62), .B(n61), .C(n55), .Y(n214) );
  NOR2X4 U188 ( .A(n180), .B(n59), .Y(n179) );
  NOR2X2 U189 ( .A(n87), .B(n88), .Y(n86) );
  AND2X4 U190 ( .A(n168), .B(n174), .Y(n59) );
  CLKINVX3 U191 ( .A(n124), .Y(n140) );
  NOR2X2 U192 ( .A(n126), .B(n127), .Y(n125) );
  NAND2BX4 U193 ( .AN(A[14]), .B(B[14]), .Y(n131) );
  NAND3X1 U194 ( .A(n58), .B(n178), .C(n53), .Y(n177) );
  NAND2X1 U195 ( .A(n58), .B(n53), .Y(n188) );
  NAND2X4 U196 ( .A(n216), .B(n39), .Y(n75) );
  NAND2X4 U197 ( .A(n104), .B(n77), .Y(n98) );
  XNOR2X4 U198 ( .A(n41), .B(n105), .Y(DIFF[4]) );
  NAND2BX4 U199 ( .AN(A[10]), .B(B[10]), .Y(n184) );
  NAND2BX4 U200 ( .AN(A[8]), .B(B[8]), .Y(n76) );
  OAI21X2 U201 ( .A0(n162), .A1(n163), .B0(n28), .Y(n173) );
  NAND2BX4 U202 ( .AN(A[11]), .B(B[11]), .Y(n174) );
  NAND2BX4 U203 ( .AN(B[11]), .B(A[11]), .Y(n194) );
  NOR2X4 U204 ( .A(n173), .B(n172), .Y(n171) );
  INVX8 U205 ( .A(n66), .Y(n65) );
  INVX8 U206 ( .A(B[5]), .Y(n66) );
  XOR2X4 U207 ( .A(n85), .B(n86), .Y(DIFF[8]) );
  NAND2BX4 U208 ( .AN(B[6]), .B(n38), .Y(n83) );
  NAND2X2 U209 ( .A(n139), .B(n142), .Y(n176) );
  XOR2X4 U210 ( .A(n170), .B(n171), .Y(DIFF[13]) );
  INVX8 U211 ( .A(n40), .Y(n70) );
  NAND3X4 U212 ( .A(n62), .B(n26), .C(n7), .Y(n84) );
  NAND2BX4 U213 ( .AN(n7), .B(n65), .Y(n78) );
  NAND2BX4 U214 ( .AN(n63), .B(n65), .Y(n201) );
  INVXL U215 ( .A(n138), .Y(n133) );
  AND2X4 U216 ( .A(n111), .B(n114), .Y(n60) );
  XOR2X4 U217 ( .A(n90), .B(n57), .Y(DIFF[7]) );
  NAND2XL U218 ( .A(n152), .B(n4), .Y(n151) );
  XOR2X2 U219 ( .A(n109), .B(n112), .Y(DIFF[2]) );
  NAND2XL U220 ( .A(n143), .B(n137), .Y(n170) );
  NOR2X1 U221 ( .A(n133), .B(n134), .Y(n128) );
  NAND2XL U222 ( .A(n4), .B(n132), .Y(n129) );
  INVX1 U223 ( .A(n117), .Y(n115) );
  AOI21XL U224 ( .A0(n145), .A1(n157), .B0(n49), .Y(n144) );
  INVXL U225 ( .A(n54), .Y(n148) );
  XNOR2X1 U226 ( .A(B[16]), .B(A[16]), .Y(n122) );
  NAND2X1 U227 ( .A(n119), .B(n120), .Y(DIFF[0]) );
  NAND2BX1 U228 ( .AN(n120), .B(n119), .Y(n117) );
  NAND2BX1 U229 ( .AN(B[0]), .B(A[0]), .Y(n119) );
  NAND2X2 U230 ( .A(n61), .B(n97), .Y(n105) );
  NAND2X4 U231 ( .A(n55), .B(n44), .Y(n202) );
  XOR2X4 U232 ( .A(n67), .B(n68), .Y(DIFF[9]) );
  NAND2BX4 U233 ( .AN(A[15]), .B(B[15]), .Y(n132) );
  NAND2BX4 U234 ( .AN(A[13]), .B(B[13]), .Y(n143) );
  OAI2BB1X4 U235 ( .A0N(n190), .A1N(n191), .B0(n192), .Y(n168) );
  NAND2BX4 U236 ( .AN(A[12]), .B(B[12]), .Y(n142) );
  NAND2BX4 U237 ( .AN(B[7]), .B(A[7]), .Y(n82) );
endmodule


module butterfly_DW01_sub_84 ( A, B, DIFF );
  input [16:0] A;
  input [16:0] B;
  output [16:0] DIFF;
  wire   n255, n256, n257, n258, n259, n260, n261, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n27, n28, n29, n31, n32, n33, n34, n35, n36, n37,
         n38, n40, n41, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254;

  NAND2X4 U3 ( .A(n15), .B(B[2]), .Y(n22) );
  INVX4 U4 ( .A(A[2]), .Y(n15) );
  AND2X4 U5 ( .A(n124), .B(n22), .Y(n126) );
  INVX4 U6 ( .A(n35), .Y(n127) );
  XOR2X4 U7 ( .A(n92), .B(n1), .Y(n4) );
  NOR2X1 U8 ( .A(n78), .B(n83), .Y(n1) );
  BUFX8 U9 ( .A(n100), .Y(n2) );
  INVX8 U10 ( .A(n253), .Y(n38) );
  CLKINVX3 U11 ( .A(n23), .Y(n24) );
  INVX8 U12 ( .A(n111), .Y(n119) );
  NAND2BX4 U13 ( .AN(B[4]), .B(A[4]), .Y(n111) );
  INVX1 U14 ( .A(n88), .Y(n44) );
  NAND3X4 U15 ( .A(n63), .B(n64), .C(n65), .Y(n217) );
  NOR2X1 U16 ( .A(n114), .B(n223), .Y(n216) );
  CLKINVX4 U17 ( .A(n254), .Y(n36) );
  AND2X4 U18 ( .A(B[1]), .B(n254), .Y(n3) );
  CLKINVX8 U19 ( .A(A[1]), .Y(n254) );
  BUFX3 U20 ( .A(A[12]), .Y(n45) );
  OAI21X4 U21 ( .A0(n47), .A1(n170), .B0(n177), .Y(n175) );
  NAND2BX2 U22 ( .AN(B[13]), .B(A[13]), .Y(n152) );
  INVX4 U23 ( .A(B[1]), .Y(n23) );
  INVX3 U24 ( .A(n253), .Y(n10) );
  INVX20 U25 ( .A(n55), .Y(DIFF[3]) );
  CLKINVX3 U26 ( .A(n46), .Y(n34) );
  XNOR2X1 U27 ( .A(B[16]), .B(A[16]), .Y(n136) );
  OAI21X1 U28 ( .A0(n137), .A1(n138), .B0(n139), .Y(n135) );
  NAND2X2 U29 ( .A(n155), .B(n149), .Y(n172) );
  NAND4X2 U30 ( .A(n65), .B(n64), .C(n63), .D(n62), .Y(n251) );
  INVX4 U31 ( .A(n75), .Y(n84) );
  CLKINVX3 U32 ( .A(n159), .Y(n193) );
  NAND3XL U33 ( .A(n65), .B(n63), .C(n64), .Y(n195) );
  INVX1 U34 ( .A(n146), .Y(n176) );
  INVX1 U35 ( .A(n151), .Y(n169) );
  NOR2BX2 U36 ( .AN(B[9]), .B(A[9]), .Y(n215) );
  AOI21X2 U37 ( .A0(n119), .A1(n64), .B0(n110), .Y(n109) );
  INVX2 U38 ( .A(n124), .Y(n123) );
  CLKINVX3 U39 ( .A(n28), .Y(n29) );
  BUFX16 U40 ( .A(n260), .Y(DIFF[2]) );
  AOI31X1 U41 ( .A0(n140), .A1(n113), .A2(n141), .B0(n142), .Y(n139) );
  NOR2X1 U42 ( .A(n156), .B(n157), .Y(n137) );
  INVX4 U43 ( .A(n102), .Y(n113) );
  AND2X1 U44 ( .A(n27), .B(n214), .Y(n5) );
  AND2X2 U45 ( .A(n64), .B(n98), .Y(n6) );
  OR2X4 U46 ( .A(n113), .B(n112), .Y(n7) );
  AND2X4 U47 ( .A(n65), .B(n11), .Y(n8) );
  OR2XL U48 ( .A(n193), .B(n213), .Y(n9) );
  NOR2X4 U49 ( .A(n171), .B(n178), .Y(n177) );
  NAND2BX4 U50 ( .AN(B[6]), .B(A[6]), .Y(n99) );
  NAND2X4 U51 ( .A(n71), .B(n93), .Y(n243) );
  NOR2BXL U52 ( .AN(n93), .B(n162), .Y(n161) );
  NAND2BX4 U53 ( .AN(A[2]), .B(B[2]), .Y(n121) );
  BUFX12 U54 ( .A(n75), .Y(n11) );
  NAND2X4 U55 ( .A(n2), .B(n20), .Y(n112) );
  NAND3X4 U56 ( .A(n79), .B(n63), .C(n81), .Y(n70) );
  NOR2X2 U57 ( .A(n215), .B(n71), .Y(n209) );
  NAND2X4 U58 ( .A(n25), .B(n93), .Y(n183) );
  BUFX16 U59 ( .A(n166), .Y(n25) );
  NAND2BX2 U60 ( .AN(A[10]), .B(B[10]), .Y(n27) );
  NAND2X1 U61 ( .A(n78), .B(n11), .Y(n72) );
  INVX4 U62 ( .A(n127), .Y(n12) );
  INVXL U63 ( .A(n25), .Y(n165) );
  XOR2X4 U64 ( .A(n53), .B(n9), .Y(n52) );
  INVX8 U65 ( .A(n63), .Y(n97) );
  AND3X4 U66 ( .A(n68), .B(n8), .C(n13), .Y(n51) );
  INVX2 U67 ( .A(n238), .Y(n13) );
  AND2X4 U68 ( .A(B[7]), .B(n43), .Y(n83) );
  INVX8 U69 ( .A(A[7]), .Y(n43) );
  AND2X2 U70 ( .A(n158), .B(n159), .Y(n208) );
  INVX8 U71 ( .A(n33), .Y(DIFF[12]) );
  OAI2BB2X4 U72 ( .B0(n18), .B1(n242), .A0N(n226), .A1N(n44), .Y(n241) );
  NOR2X4 U73 ( .A(n223), .B(n252), .Y(n14) );
  NAND2X4 U74 ( .A(n17), .B(n237), .Y(n228) );
  BUFX20 U75 ( .A(n259), .Y(DIFF[4]) );
  NAND2X4 U76 ( .A(n65), .B(n64), .Y(n108) );
  NOR2X4 U77 ( .A(n18), .B(n234), .Y(n230) );
  NAND2X4 U78 ( .A(n65), .B(n64), .Y(n184) );
  NAND2X4 U79 ( .A(n31), .B(n104), .Y(n114) );
  BUFX20 U80 ( .A(n103), .Y(n31) );
  CLKINVX8 U81 ( .A(n15), .Y(n16) );
  NOR2X4 U82 ( .A(n184), .B(n185), .Y(n181) );
  NAND2X2 U83 ( .A(n62), .B(n63), .Y(n185) );
  INVX8 U84 ( .A(n125), .Y(n253) );
  BUFX8 U85 ( .A(n68), .Y(n17) );
  NOR2X4 U86 ( .A(n240), .B(n241), .Y(n227) );
  NAND2X2 U87 ( .A(n243), .B(n226), .Y(n242) );
  NOR3BX4 U88 ( .AN(n226), .B(n25), .C(n233), .Y(n240) );
  NAND2X4 U89 ( .A(n87), .B(n11), .Y(n233) );
  NAND4BBX4 U90 ( .AN(n74), .BN(n84), .C(n62), .D(n77), .Y(n73) );
  AOI21X4 U91 ( .A0(n158), .A1(n159), .B0(n172), .Y(n178) );
  NOR2X4 U92 ( .A(n183), .B(n162), .Y(n182) );
  NAND2X4 U93 ( .A(n88), .B(n245), .Y(n244) );
  NAND2BX4 U94 ( .AN(B[2]), .B(n16), .Y(n124) );
  NAND2X4 U95 ( .A(n11), .B(n87), .Y(n18) );
  NAND2BX4 U96 ( .AN(A[2]), .B(B[2]), .Y(n21) );
  NAND3BX4 U97 ( .AN(n83), .B(n63), .C(n64), .Y(n238) );
  NAND4X2 U98 ( .A(n23), .B(n38), .C(n121), .D(n36), .Y(n101) );
  NOR2XL U99 ( .A(n153), .B(n154), .Y(n141) );
  AOI21XL U100 ( .A0(n160), .A1(n161), .B0(n153), .Y(n156) );
  NOR2X2 U101 ( .A(n83), .B(n153), .Y(n206) );
  CLKINVX3 U102 ( .A(n153), .Y(n173) );
  NOR3X4 U103 ( .A(n238), .B(n18), .C(n239), .Y(n237) );
  NAND2X4 U104 ( .A(n23), .B(n36), .Y(n129) );
  NOR2X2 U105 ( .A(n200), .B(n201), .Y(n199) );
  NOR2BX1 U106 ( .AN(A[5]), .B(B[5]), .Y(n201) );
  INVX3 U107 ( .A(n98), .Y(n110) );
  NAND4X4 U108 ( .A(n19), .B(n31), .C(n102), .D(n34), .Y(n68) );
  AND2X4 U109 ( .A(n101), .B(n100), .Y(n19) );
  NAND2X4 U110 ( .A(n31), .B(n104), .Y(n252) );
  OAI21X2 U111 ( .A0(n191), .A1(n158), .B0(n192), .Y(n190) );
  NAND4BX4 U112 ( .AN(n24), .B(n35), .C(n38), .D(n36), .Y(n20) );
  NAND4BX2 U113 ( .AN(n82), .B(n250), .C(n63), .D(n62), .Y(n249) );
  INVX8 U114 ( .A(n222), .Y(n82) );
  OAI21X4 U115 ( .A0(n97), .A1(n98), .B0(n99), .Y(n96) );
  CLKINVX2 U116 ( .A(A[3]), .Y(n28) );
  BUFX12 U117 ( .A(n255), .Y(DIFF[15]) );
  BUFX12 U118 ( .A(n132), .Y(n37) );
  NAND2X4 U119 ( .A(B[1]), .B(n254), .Y(n132) );
  BUFX20 U120 ( .A(n256), .Y(DIFF[10]) );
  BUFX20 U121 ( .A(n4), .Y(DIFF[7]) );
  NAND4X4 U122 ( .A(n37), .B(n22), .C(n38), .D(n32), .Y(n103) );
  CLKINVX20 U123 ( .A(n133), .Y(n32) );
  XOR2X4 U124 ( .A(n204), .B(n205), .Y(n33) );
  NAND2X4 U125 ( .A(n27), .B(n65), .Y(n239) );
  XOR2X2 U126 ( .A(n122), .B(n126), .Y(n260) );
  NAND4X1 U127 ( .A(n147), .B(n146), .C(n155), .D(n149), .Y(n138) );
  NAND2BX2 U128 ( .AN(A[14]), .B(B[14]), .Y(n146) );
  NAND2XL U129 ( .A(n31), .B(n104), .Y(n202) );
  NAND2BX4 U130 ( .AN(A[2]), .B(B[2]), .Y(n35) );
  BUFX20 U131 ( .A(n85), .Y(n65) );
  NAND2BX4 U132 ( .AN(A[4]), .B(B[4]), .Y(n85) );
  BUFX20 U133 ( .A(n261), .Y(DIFF[1]) );
  NOR2X4 U134 ( .A(n7), .B(n202), .Y(n194) );
  NOR2X4 U135 ( .A(n118), .B(n119), .Y(n117) );
  NAND3X2 U136 ( .A(n63), .B(n119), .C(n64), .Y(n95) );
  NOR2X4 U137 ( .A(n162), .B(n219), .Y(n218) );
  INVX3 U138 ( .A(n104), .Y(n46) );
  OAI2BB1X4 U139 ( .A0N(n181), .A1N(n68), .B0(n182), .Y(n89) );
  XOR2X4 U140 ( .A(n175), .B(n41), .Y(n40) );
  OR2X4 U141 ( .A(n169), .B(n176), .Y(n41) );
  NAND3BX2 U142 ( .AN(n243), .B(n249), .C(n25), .Y(n247) );
  NAND2X2 U143 ( .A(n236), .B(n235), .Y(n250) );
  NAND3X4 U144 ( .A(n20), .B(n2), .C(n102), .Y(n223) );
  INVX8 U145 ( .A(n40), .Y(DIFF[14]) );
  NAND2X4 U146 ( .A(n88), .B(n214), .Y(n210) );
  NOR2X4 U147 ( .A(n212), .B(n213), .Y(n211) );
  INVX8 U148 ( .A(n220), .Y(n162) );
  NAND4BX4 U149 ( .AN(n82), .B(n221), .C(n63), .D(n62), .Y(n220) );
  AND2X2 U150 ( .A(n38), .B(n104), .Y(n56) );
  NAND2X4 U151 ( .A(n43), .B(B[7]), .Y(n76) );
  AOI21X4 U152 ( .A0(n122), .A1(n12), .B0(n123), .Y(n120) );
  BUFX20 U153 ( .A(n76), .Y(n62) );
  NAND2XL U154 ( .A(n155), .B(n62), .Y(n203) );
  NAND4BX4 U155 ( .AN(n224), .B(n225), .C(n27), .D(n87), .Y(n153) );
  NAND2BX4 U156 ( .AN(B[11]), .B(A[11]), .Y(n159) );
  NAND2BX4 U157 ( .AN(B[8]), .B(A[8]), .Y(n71) );
  NOR2BX2 U158 ( .AN(A[4]), .B(B[4]), .Y(n200) );
  XOR2X4 U159 ( .A(n130), .B(n131), .Y(n261) );
  NOR2BX4 U160 ( .AN(n129), .B(n3), .Y(n131) );
  NAND3X4 U161 ( .A(n228), .B(n227), .C(n229), .Y(n53) );
  NOR2X4 U162 ( .A(n51), .B(n69), .Y(n67) );
  OAI21X2 U163 ( .A0(n47), .A1(n170), .B0(n177), .Y(n168) );
  INVX2 U164 ( .A(n65), .Y(n118) );
  INVX8 U165 ( .A(n89), .Y(n47) );
  NAND2X2 U166 ( .A(n25), .B(n93), .Y(n197) );
  NAND2X2 U167 ( .A(n25), .B(n93), .Y(n219) );
  NOR2X4 U168 ( .A(n14), .B(n251), .Y(n246) );
  BUFX20 U169 ( .A(n86), .Y(n64) );
  NAND2BX4 U170 ( .AN(A[5]), .B(B[5]), .Y(n86) );
  XOR2X4 U171 ( .A(n120), .B(n56), .Y(n55) );
  NOR3X4 U172 ( .A(n114), .B(n113), .C(n112), .Y(n107) );
  NAND4X2 U173 ( .A(n70), .B(n73), .C(n72), .D(n71), .Y(n69) );
  NAND2X2 U174 ( .A(n89), .B(n48), .Y(n49) );
  XOR2X4 U175 ( .A(n17), .B(n117), .Y(n259) );
  OAI21X4 U176 ( .A0(n3), .A1(n128), .B0(n129), .Y(n122) );
  OAI2BB1X4 U177 ( .A0N(n206), .A1N(n207), .B0(n208), .Y(n204) );
  INVX8 U178 ( .A(n52), .Y(DIFF[11]) );
  NAND2X4 U179 ( .A(n47), .B(n90), .Y(n50) );
  NAND2X4 U180 ( .A(n49), .B(n50), .Y(DIFF[8]) );
  INVXL U181 ( .A(n90), .Y(n48) );
  NOR2X4 U182 ( .A(n91), .B(n84), .Y(n90) );
  NAND4BX2 U183 ( .AN(n83), .B(n63), .C(n65), .D(n64), .Y(n154) );
  NOR3X4 U184 ( .A(n97), .B(n83), .C(n212), .Y(n231) );
  NOR2X2 U185 ( .A(n83), .B(n84), .Y(n79) );
  BUFX20 U186 ( .A(n257), .Y(DIFF[9]) );
  NAND2BX4 U187 ( .AN(B[3]), .B(n29), .Y(n104) );
  NAND2BX4 U188 ( .AN(A[12]), .B(B[12]), .Y(n155) );
  NAND3BX4 U189 ( .AN(B[2]), .B(n10), .C(n16), .Y(n100) );
  CLKINVX2 U190 ( .A(n172), .Y(n174) );
  NAND2X2 U191 ( .A(n173), .B(n174), .Y(n170) );
  NAND2XL U192 ( .A(n87), .B(n88), .Y(n66) );
  AOI21X2 U193 ( .A0(n235), .A1(n111), .B0(n82), .Y(n81) );
  AOI21X2 U194 ( .A0(n193), .A1(n155), .B0(n148), .Y(n192) );
  INVXL U195 ( .A(n214), .Y(n232) );
  INVX4 U196 ( .A(n93), .Y(n78) );
  XOR2X4 U197 ( .A(n105), .B(n106), .Y(n258) );
  NOR2X2 U198 ( .A(n203), .B(n153), .Y(n188) );
  XOR2X4 U199 ( .A(n54), .B(n167), .Y(n255) );
  NAND2X2 U200 ( .A(n145), .B(n147), .Y(n54) );
  INVX1 U201 ( .A(n233), .Y(n248) );
  INVX8 U202 ( .A(n226), .Y(n212) );
  AOI21X2 U203 ( .A0(n152), .A1(n179), .B0(n180), .Y(n171) );
  NAND2XL U204 ( .A(n151), .B(n152), .Y(n150) );
  NAND2XL U205 ( .A(n146), .B(n147), .Y(n144) );
  NAND2XL U206 ( .A(n155), .B(n179), .Y(n205) );
  INVX1 U207 ( .A(n155), .Y(n191) );
  NAND2XL U208 ( .A(n149), .B(n152), .Y(n186) );
  INVX1 U209 ( .A(n71), .Y(n91) );
  INVXL U210 ( .A(n149), .Y(n180) );
  INVX1 U211 ( .A(n130), .Y(n128) );
  NAND2X1 U212 ( .A(n221), .B(n222), .Y(n234) );
  INVXL U213 ( .A(B[6]), .Y(n77) );
  INVX1 U214 ( .A(n138), .Y(n140) );
  OAI21XL U215 ( .A0(n143), .A1(n144), .B0(n145), .Y(n142) );
  AOI21X1 U216 ( .A0(n163), .A1(n164), .B0(n165), .Y(n160) );
  INVXL U217 ( .A(n154), .Y(n163) );
  AOI21XL U218 ( .A0(n148), .A1(n149), .B0(n150), .Y(n143) );
  BUFX20 U219 ( .A(n80), .Y(n63) );
  NAND2BX1 U220 ( .AN(A[15]), .B(B[15]), .Y(n147) );
  NAND2BX1 U221 ( .AN(B[15]), .B(A[15]), .Y(n145) );
  NAND2BX1 U222 ( .AN(B[14]), .B(A[14]), .Y(n151) );
  INVXL U223 ( .A(A[6]), .Y(n74) );
  NAND2X1 U224 ( .A(n133), .B(n134), .Y(DIFF[0]) );
  NAND2BX1 U225 ( .AN(n134), .B(n133), .Y(n130) );
  NAND2BX1 U226 ( .AN(A[0]), .B(B[0]), .Y(n134) );
  NAND2BX1 U227 ( .AN(B[0]), .B(A[0]), .Y(n133) );
  BUFX20 U228 ( .A(n258), .Y(DIFF[6]) );
  NAND2BX2 U229 ( .AN(B[5]), .B(A[5]), .Y(n98) );
  NAND3BX4 U230 ( .AN(B[6]), .B(A[6]), .C(n62), .Y(n166) );
  NOR2BX2 U231 ( .AN(n99), .B(n97), .Y(n106) );
  NOR3X2 U232 ( .A(n199), .B(n97), .C(n82), .Y(n198) );
  NAND2XL U233 ( .A(n158), .B(n159), .Y(n157) );
  NOR2BX1 U234 ( .AN(B[8]), .B(A[8]), .Y(n224) );
  NAND2X4 U235 ( .A(n68), .B(n65), .Y(n116) );
  NAND4BXL U236 ( .AN(n46), .B(n31), .C(n2), .D(n20), .Y(n164) );
  XOR2X4 U237 ( .A(n67), .B(n66), .Y(n257) );
  OAI21X4 U238 ( .A0(n217), .A1(n14), .B0(n94), .Y(n92) );
  NOR2BX4 U239 ( .AN(n95), .B(n96), .Y(n94) );
  OAI21X4 U240 ( .A0(n107), .A1(n108), .B0(n109), .Y(n105) );
  XOR2X4 U241 ( .A(n115), .B(n6), .Y(DIFF[5]) );
  NAND2X4 U242 ( .A(n116), .B(n111), .Y(n115) );
  XOR2X4 U243 ( .A(n135), .B(n136), .Y(DIFF[16]) );
  AOI21X4 U244 ( .A0(n168), .A1(n146), .B0(n169), .Y(n167) );
  XOR2X4 U245 ( .A(n187), .B(n186), .Y(DIFF[13]) );
  AOI21X4 U246 ( .A0(n188), .A1(n189), .B0(n190), .Y(n187) );
  CLKINVX3 U247 ( .A(n179), .Y(n148) );
  OAI21X4 U248 ( .A0(n194), .A1(n195), .B0(n196), .Y(n189) );
  NOR2X4 U249 ( .A(n197), .B(n198), .Y(n196) );
  NAND2BX4 U250 ( .AN(A[13]), .B(B[13]), .Y(n149) );
  NAND2BX4 U251 ( .AN(B[12]), .B(n45), .Y(n179) );
  OAI21X4 U252 ( .A0(n209), .A1(n210), .B0(n211), .Y(n158) );
  OAI21X4 U253 ( .A0(n216), .A1(n217), .B0(n218), .Y(n207) );
  CLKINVX3 U254 ( .A(n225), .Y(n213) );
  NAND2BX4 U255 ( .AN(A[11]), .B(B[11]), .Y(n225) );
  AOI21X4 U256 ( .A0(n230), .A1(n231), .B0(n232), .Y(n229) );
  NAND2X4 U257 ( .A(n235), .B(n236), .Y(n221) );
  XOR2X4 U258 ( .A(n244), .B(n5), .Y(n256) );
  NAND2BX4 U259 ( .AN(B[10]), .B(A[10]), .Y(n214) );
  NAND2BX4 U260 ( .AN(A[10]), .B(B[10]), .Y(n226) );
  OAI21X4 U261 ( .A0(n246), .A1(n247), .B0(n248), .Y(n245) );
  NAND2BX4 U262 ( .AN(A[8]), .B(B[8]), .Y(n75) );
  NAND2BX4 U263 ( .AN(A[9]), .B(B[9]), .Y(n87) );
  NAND2BX4 U264 ( .AN(B[5]), .B(A[5]), .Y(n235) );
  NAND2BX4 U265 ( .AN(B[4]), .B(A[4]), .Y(n236) );
  NAND2BX4 U266 ( .AN(A[5]), .B(B[5]), .Y(n222) );
  NAND2BX4 U267 ( .AN(B[7]), .B(A[7]), .Y(n93) );
  NAND2BX4 U268 ( .AN(A[6]), .B(B[6]), .Y(n80) );
  NAND4BX4 U269 ( .AN(n253), .B(n37), .C(n21), .D(n134), .Y(n102) );
  NAND2BX4 U270 ( .AN(A[3]), .B(B[3]), .Y(n125) );
  NAND2BX4 U271 ( .AN(B[9]), .B(A[9]), .Y(n88) );
endmodule


module butterfly_DW01_add_116 ( A, B, SUM );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  wire   n217, n218, n219, n220, n221, n222, n223, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n24, n25, n27, n28, n29, n30, n31, n32, n34, n35, n36, n37, n38,
         n39, n40, n41, n43, n44, n45, n46, n47, n48, n49, n50, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216;

  CLKBUFX3 U2 ( .A(n85), .Y(n10) );
  OR2X4 U3 ( .A(A[6]), .B(B[6]), .Y(n1) );
  BUFX8 U4 ( .A(A[2]), .Y(n25) );
  NAND2XL U5 ( .A(B[10]), .B(A[10]), .Y(n192) );
  AND3X2 U6 ( .A(n215), .B(n17), .C(n20), .Y(n2) );
  NOR2X4 U7 ( .A(n108), .B(n3), .Y(n56) );
  NAND2X4 U8 ( .A(n4), .B(n17), .Y(n3) );
  CLKINVX20 U9 ( .A(n109), .Y(n4) );
  INVX2 U10 ( .A(n12), .Y(n5) );
  NOR2X4 U11 ( .A(B[2]), .B(A[2]), .Y(n12) );
  NAND2X2 U12 ( .A(B[8]), .B(A[8]), .Y(n71) );
  NAND2X2 U13 ( .A(n73), .B(n71), .Y(n166) );
  NOR2X2 U14 ( .A(n16), .B(B[7]), .Y(n211) );
  CLKINVX8 U15 ( .A(n29), .Y(n30) );
  NAND2BX4 U16 ( .AN(n12), .B(n56), .Y(n27) );
  AND2X4 U17 ( .A(n11), .B(n90), .Y(n31) );
  INVX20 U18 ( .A(n47), .Y(SUM[8]) );
  NAND2BX2 U19 ( .AN(n133), .B(n166), .Y(n178) );
  BUFX16 U20 ( .A(n94), .Y(n34) );
  NAND3X2 U21 ( .A(n38), .B(B[6]), .C(n70), .Y(n9) );
  NOR2X4 U22 ( .A(n162), .B(n163), .Y(n161) );
  NOR3X2 U23 ( .A(n164), .B(n48), .C(n165), .Y(n163) );
  AOI21X4 U24 ( .A0(n207), .A1(n208), .B0(n50), .Y(n206) );
  NOR2X4 U25 ( .A(n97), .B(n209), .Y(n208) );
  NAND3X4 U26 ( .A(n38), .B(B[6]), .C(n70), .Y(n145) );
  NAND2X1 U27 ( .A(n179), .B(n127), .Y(n176) );
  NAND2BX4 U28 ( .AN(n127), .B(n170), .Y(n169) );
  NAND2X4 U29 ( .A(B[12]), .B(A[12]), .Y(n127) );
  NOR2X2 U30 ( .A(n164), .B(n178), .Y(n177) );
  OAI21X2 U31 ( .A0(n48), .A1(n191), .B0(n192), .Y(n190) );
  NAND2X1 U32 ( .A(B[13]), .B(A[13]), .Y(n125) );
  INVX8 U33 ( .A(n120), .Y(n132) );
  OR2X4 U34 ( .A(A[14]), .B(B[14]), .Y(n120) );
  OR2X4 U35 ( .A(A[13]), .B(B[13]), .Y(n170) );
  AND2X2 U36 ( .A(A[10]), .B(B[10]), .Y(n49) );
  INVX3 U37 ( .A(n98), .Y(n24) );
  INVX1 U38 ( .A(B[11]), .Y(n18) );
  AOI21X2 U39 ( .A0(n60), .A1(n61), .B0(n62), .Y(n59) );
  NOR3X2 U40 ( .A(n63), .B(n64), .C(n65), .Y(n61) );
  NOR2BX2 U41 ( .AN(n78), .B(n211), .Y(n77) );
  BUFX16 U42 ( .A(n222), .Y(SUM[4]) );
  CLKBUFX8 U43 ( .A(A[6]), .Y(n38) );
  NOR2BX1 U44 ( .AN(n125), .B(n154), .Y(n168) );
  INVX1 U45 ( .A(n169), .Y(n154) );
  NAND2X2 U46 ( .A(n171), .B(n170), .Y(n165) );
  NOR2X1 U47 ( .A(n116), .B(n133), .Y(n174) );
  NOR2BX2 U48 ( .AN(n125), .B(n126), .Y(n173) );
  INVX4 U49 ( .A(n68), .Y(n97) );
  NOR2BX2 U50 ( .AN(n192), .B(n200), .Y(n199) );
  INVX1 U51 ( .A(n184), .Y(n200) );
  NAND2X2 U52 ( .A(B[9]), .B(A[9]), .Y(n73) );
  NAND2X1 U53 ( .A(n85), .B(n210), .Y(n84) );
  NOR2BX1 U54 ( .AN(n156), .B(n116), .Y(n160) );
  OAI2BB1X2 U55 ( .A0N(n156), .A1N(n167), .B0(n168), .Y(n162) );
  INVX4 U56 ( .A(n171), .Y(n133) );
  INVX1 U57 ( .A(n170), .Y(n126) );
  NAND2X1 U58 ( .A(B[15]), .B(A[15]), .Y(n119) );
  CLKINVX3 U59 ( .A(n187), .Y(n62) );
  NOR3BX1 U60 ( .AN(n134), .B(n135), .C(n7), .Y(n112) );
  AOI21X1 U61 ( .A0(n136), .A1(n137), .B0(n116), .Y(n135) );
  INVX3 U62 ( .A(n34), .Y(n29) );
  AND2X2 U63 ( .A(B[8]), .B(A[8]), .Y(n50) );
  INVX4 U64 ( .A(n78), .Y(n65) );
  AND2X2 U65 ( .A(n140), .B(n141), .Y(n6) );
  INVX1 U66 ( .A(n67), .Y(n41) );
  AND2X1 U67 ( .A(B[10]), .B(A[10]), .Y(n7) );
  AND2X4 U68 ( .A(n214), .B(n17), .Y(n8) );
  NAND2X1 U69 ( .A(B[6]), .B(n38), .Y(n81) );
  OAI2BB1X2 U70 ( .A0N(n174), .A1N(n74), .B0(n175), .Y(n172) );
  NAND2X4 U71 ( .A(B[4]), .B(A[4]), .Y(n67) );
  NAND2X2 U72 ( .A(B[4]), .B(A[4]), .Y(n210) );
  NOR2X2 U73 ( .A(n176), .B(n177), .Y(n175) );
  INVX2 U74 ( .A(n157), .Y(n151) );
  NOR2X2 U75 ( .A(n212), .B(n197), .Y(n203) );
  NAND2BX4 U76 ( .AN(n12), .B(n8), .Y(n11) );
  NAND2X2 U77 ( .A(A[2]), .B(B[2]), .Y(n102) );
  NOR2BX2 U78 ( .AN(n85), .B(n97), .Y(n96) );
  BUFX3 U79 ( .A(A[7]), .Y(n16) );
  NOR2BX1 U80 ( .AN(n127), .B(n133), .Y(n180) );
  NAND2X4 U81 ( .A(B[7]), .B(n16), .Y(n78) );
  INVX8 U82 ( .A(n19), .Y(n17) );
  NOR2X4 U83 ( .A(A[6]), .B(B[6]), .Y(n209) );
  NAND2X2 U84 ( .A(n1), .B(n70), .Y(n35) );
  INVX8 U85 ( .A(n145), .Y(n64) );
  OR2X4 U86 ( .A(B[5]), .B(A[5]), .Y(n14) );
  NAND2BX4 U87 ( .AN(n164), .B(n166), .Y(n183) );
  OAI2BB1X4 U88 ( .A0N(n85), .A1N(n67), .B0(n14), .Y(n66) );
  AND2X2 U89 ( .A(n90), .B(n17), .Y(n101) );
  BUFX1 U90 ( .A(n128), .Y(n13) );
  BUFX20 U91 ( .A(n217), .Y(SUM[14]) );
  INVXL U92 ( .A(n87), .Y(n15) );
  OR2X2 U93 ( .A(n97), .B(n209), .Y(n80) );
  NOR2BX4 U94 ( .AN(n146), .B(n144), .Y(n195) );
  NAND2BX4 U95 ( .AN(n144), .B(n146), .Y(n186) );
  NAND2X4 U96 ( .A(n85), .B(n67), .Y(n146) );
  AND2X4 U97 ( .A(B[1]), .B(A[1]), .Y(n20) );
  NOR2X4 U98 ( .A(A[3]), .B(B[3]), .Y(n19) );
  OAI21X2 U99 ( .A0(n138), .A1(n139), .B0(n6), .Y(n137) );
  NAND2X4 U100 ( .A(n83), .B(n68), .Y(n212) );
  NOR2BX2 U101 ( .AN(n21), .B(n108), .Y(n107) );
  NAND2BX4 U102 ( .AN(A[11]), .B(n18), .Y(n128) );
  NAND2BX4 U103 ( .AN(n65), .B(n9), .Y(n185) );
  INVX4 U104 ( .A(n20), .Y(n21) );
  INVXL U105 ( .A(n64), .Y(n22) );
  AOI2BB1X1 U106 ( .A0N(n169), .A1N(n132), .B0(n155), .Y(n153) );
  OAI2BB1X2 U107 ( .A0N(n74), .A1N(n160), .B0(n161), .Y(n158) );
  BUFX16 U108 ( .A(n223), .Y(SUM[1]) );
  INVX3 U109 ( .A(n83), .Y(n98) );
  NAND2X4 U110 ( .A(B[5]), .B(A[5]), .Y(n85) );
  OR2X4 U111 ( .A(n191), .B(n62), .Y(n194) );
  NAND2X2 U112 ( .A(n184), .B(n72), .Y(n191) );
  NAND4X4 U113 ( .A(n187), .B(n72), .C(n128), .D(n184), .Y(n116) );
  NAND2X4 U114 ( .A(n70), .B(n1), .Y(n197) );
  INVX8 U115 ( .A(n45), .Y(SUM[10]) );
  NOR2X4 U116 ( .A(n2), .B(n87), .Y(n86) );
  CLKINVX2 U117 ( .A(n88), .Y(n87) );
  OAI21XL U118 ( .A0(n143), .A1(n144), .B0(n22), .Y(n142) );
  INVX8 U119 ( .A(n105), .Y(n108) );
  XOR2X4 U120 ( .A(n76), .B(n77), .Y(n28) );
  NOR2XL U121 ( .A(n126), .B(n127), .Y(n122) );
  NAND2X4 U122 ( .A(n31), .B(n86), .Y(n82) );
  DLY1X1 U123 ( .A(n11), .Y(n32) );
  BUFX20 U124 ( .A(n28), .Y(SUM[7]) );
  OAI2BB1X2 U125 ( .A0N(n103), .A1N(n5), .B0(n102), .Y(n100) );
  NOR2X4 U126 ( .A(n212), .B(n197), .Y(n196) );
  NAND3X4 U127 ( .A(n69), .B(n70), .C(n14), .Y(n144) );
  OAI2BB1X4 U128 ( .A0N(n24), .A1N(n34), .B0(n67), .Y(n95) );
  AOI21X4 U129 ( .A0(n30), .A1(n203), .B0(n204), .Y(n201) );
  NOR2X4 U130 ( .A(n35), .B(n66), .Y(n63) );
  NAND2X4 U131 ( .A(n89), .B(n88), .Y(n213) );
  OR2X4 U132 ( .A(A[8]), .B(B[8]), .Y(n187) );
  INVXL U133 ( .A(n2), .Y(n36) );
  NOR2X4 U134 ( .A(n37), .B(n194), .Y(n189) );
  AND2X4 U135 ( .A(n60), .B(n193), .Y(n37) );
  INVX8 U136 ( .A(n39), .Y(SUM[13]) );
  XOR2X4 U137 ( .A(n172), .B(n40), .Y(n39) );
  CLKINVX20 U138 ( .A(n173), .Y(n40) );
  OAI2BB1X4 U139 ( .A0N(n106), .A1N(n105), .B0(n21), .Y(n103) );
  XOR2X4 U140 ( .A(n110), .B(n111), .Y(SUM[16]) );
  OAI21X4 U141 ( .A0(n112), .A1(n113), .B0(n114), .Y(n110) );
  NAND2X2 U142 ( .A(n167), .B(n171), .Y(n179) );
  NOR2BX4 U143 ( .AN(n67), .B(n98), .Y(n99) );
  AOI21X4 U144 ( .A0(n82), .A1(n24), .B0(n84), .Y(n79) );
  BUFX20 U145 ( .A(n221), .Y(SUM[5]) );
  BUFX20 U146 ( .A(n220), .Y(SUM[6]) );
  OAI21X4 U147 ( .A0(n151), .A1(n152), .B0(n153), .Y(n149) );
  NAND2X2 U148 ( .A(B[3]), .B(A[3]), .Y(n90) );
  NOR2X4 U149 ( .A(n34), .B(n41), .Y(n93) );
  BUFX20 U150 ( .A(n218), .Y(SUM[12]) );
  NAND2X1 U151 ( .A(n13), .B(n147), .Y(n43) );
  NAND2X1 U152 ( .A(B[11]), .B(A[11]), .Y(n147) );
  XOR2X4 U153 ( .A(n58), .B(n57), .Y(n219) );
  NOR2X4 U154 ( .A(n59), .B(n50), .Y(n58) );
  XOR2X2 U155 ( .A(n34), .B(n99), .Y(n222) );
  NOR2BX4 U156 ( .AN(n81), .B(n209), .Y(n92) );
  NAND2X4 U157 ( .A(n34), .B(n196), .Y(n60) );
  BUFX20 U158 ( .A(n219), .Y(SUM[9]) );
  NOR2X4 U159 ( .A(n65), .B(n64), .Y(n205) );
  OAI2BB1X4 U160 ( .A0N(n181), .A1N(n74), .B0(n182), .Y(n157) );
  NAND3X4 U161 ( .A(B[2]), .B(n17), .C(n25), .Y(n88) );
  NOR2X2 U162 ( .A(n195), .B(n185), .Y(n193) );
  AND2X2 U163 ( .A(n73), .B(n71), .Y(n48) );
  OAI2BB1X4 U164 ( .A0N(n128), .A1N(n49), .B0(n147), .Y(n167) );
  OR2X2 U165 ( .A(A[15]), .B(B[15]), .Y(n121) );
  NOR2XL U166 ( .A(n211), .B(n209), .Y(n141) );
  NAND3X4 U167 ( .A(n184), .B(n72), .C(n128), .Y(n164) );
  INVX8 U168 ( .A(n199), .Y(n46) );
  XOR2X4 U169 ( .A(n188), .B(n43), .Y(SUM[11]) );
  NAND2XL U170 ( .A(n72), .B(n73), .Y(n57) );
  NAND2XL U171 ( .A(n72), .B(n187), .Y(n202) );
  NAND2XL U172 ( .A(n44), .B(n13), .Y(n113) );
  AND2X2 U173 ( .A(n129), .B(n130), .Y(n44) );
  NOR2BX2 U174 ( .AN(n124), .B(n132), .Y(n159) );
  NOR2BX4 U175 ( .AN(n119), .B(n131), .Y(n150) );
  OR2X4 U176 ( .A(A[12]), .B(B[12]), .Y(n171) );
  NAND2XL U177 ( .A(n124), .B(n125), .Y(n123) );
  NAND2XL U178 ( .A(n120), .B(n121), .Y(n118) );
  OR2X4 U179 ( .A(A[1]), .B(B[1]), .Y(n105) );
  XOR2X2 U180 ( .A(B[16]), .B(A[16]), .Y(n111) );
  NOR2XL U181 ( .A(n97), .B(n98), .Y(n140) );
  XOR2X4 U182 ( .A(n198), .B(n46), .Y(n45) );
  INVX1 U183 ( .A(n116), .Y(n181) );
  XNOR2X4 U184 ( .A(n74), .B(n75), .Y(n47) );
  NOR2BXL U185 ( .AN(n147), .B(n148), .Y(n134) );
  NOR2X1 U186 ( .A(n142), .B(n65), .Y(n136) );
  INVXL U187 ( .A(n146), .Y(n143) );
  NOR2XL U188 ( .A(n126), .B(n133), .Y(n129) );
  NOR2X1 U189 ( .A(n131), .B(n132), .Y(n130) );
  NAND2BXL U190 ( .AN(n132), .B(n156), .Y(n152) );
  AOI21X2 U191 ( .A0(n85), .A1(n210), .B0(n211), .Y(n207) );
  NAND2XL U192 ( .A(n32), .B(n90), .Y(n138) );
  OAI21XL U193 ( .A0(n132), .A1(n125), .B0(n124), .Y(n155) );
  INVX1 U194 ( .A(n121), .Y(n131) );
  INVX1 U195 ( .A(n115), .Y(n114) );
  OAI21XL U196 ( .A0(n117), .A1(n118), .B0(n119), .Y(n115) );
  NOR2X1 U197 ( .A(n122), .B(n123), .Y(n117) );
  NAND2X1 U198 ( .A(B[14]), .B(A[14]), .Y(n124) );
  INVX1 U199 ( .A(n109), .Y(n106) );
  AND2X2 U200 ( .A(n109), .B(n216), .Y(SUM[0]) );
  OR2X2 U201 ( .A(A[0]), .B(B[0]), .Y(n216) );
  NAND2X1 U202 ( .A(B[0]), .B(A[0]), .Y(n109) );
  NAND3BX4 U203 ( .AN(n213), .B(n27), .C(n90), .Y(n94) );
  OAI21X4 U204 ( .A0(n93), .A1(n212), .B0(n10), .Y(n91) );
  NAND2XL U205 ( .A(n15), .B(n36), .Y(n139) );
  NOR2BX4 U206 ( .AN(n71), .B(n62), .Y(n75) );
  OAI21X4 U207 ( .A0(n79), .A1(n80), .B0(n81), .Y(n76) );
  XOR2X4 U208 ( .A(n91), .B(n92), .Y(n220) );
  XOR2X4 U209 ( .A(n95), .B(n96), .Y(n221) );
  XOR2X4 U210 ( .A(n100), .B(n101), .Y(SUM[3]) );
  XOR2X4 U211 ( .A(n103), .B(n104), .Y(SUM[2]) );
  NOR2BX4 U212 ( .AN(n102), .B(n12), .Y(n104) );
  XOR2X4 U213 ( .A(n106), .B(n107), .Y(n223) );
  XOR2X4 U214 ( .A(n149), .B(n150), .Y(SUM[15]) );
  XOR2X4 U215 ( .A(n158), .B(n159), .Y(n217) );
  CLKINVX3 U216 ( .A(n165), .Y(n156) );
  XOR2X4 U217 ( .A(n157), .B(n180), .Y(n218) );
  NOR2X4 U218 ( .A(n148), .B(n167), .Y(n182) );
  CLKINVX3 U219 ( .A(n183), .Y(n148) );
  NAND3BX4 U220 ( .AN(n185), .B(n60), .C(n186), .Y(n74) );
  NOR2X4 U221 ( .A(n189), .B(n190), .Y(n188) );
  OR2X4 U222 ( .A(A[10]), .B(B[10]), .Y(n184) );
  OAI21X4 U223 ( .A0(n201), .A1(n202), .B0(n73), .Y(n198) );
  OR2X4 U224 ( .A(A[9]), .B(B[9]), .Y(n72) );
  NAND2X4 U225 ( .A(n206), .B(n205), .Y(n204) );
  OR2X4 U226 ( .A(A[6]), .B(B[6]), .Y(n69) );
  OR2X4 U227 ( .A(A[7]), .B(B[7]), .Y(n70) );
  OR2X4 U228 ( .A(A[5]), .B(B[5]), .Y(n68) );
  OR2X4 U229 ( .A(A[4]), .B(B[4]), .Y(n83) );
  NOR2X4 U230 ( .A(n108), .B(n109), .Y(n214) );
  NAND3X4 U231 ( .A(n215), .B(n17), .C(n20), .Y(n89) );
  OR2X4 U232 ( .A(A[2]), .B(B[2]), .Y(n215) );
endmodule


module butterfly_DW01_add_119 ( A, B, SUM );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182;

  INVX1 U2 ( .A(B[5]), .Y(n1) );
  BUFX4 U3 ( .A(n54), .Y(n26) );
  NAND2X4 U4 ( .A(n57), .B(n56), .Y(n55) );
  INVX8 U5 ( .A(n29), .Y(n28) );
  CLKBUFX8 U6 ( .A(n64), .Y(n29) );
  NOR2XL U7 ( .A(n31), .B(n64), .Y(n2) );
  INVXL U8 ( .A(n81), .Y(n84) );
  CLKBUFX4 U9 ( .A(B[3]), .Y(n5) );
  NOR2X4 U10 ( .A(A[7]), .B(B[7]), .Y(n31) );
  OR2X4 U11 ( .A(A[7]), .B(B[7]), .Y(n153) );
  NAND3X1 U12 ( .A(n6), .B(n24), .C(n51), .Y(n3) );
  XNOR2X2 U13 ( .A(n35), .B(n76), .Y(n4) );
  OR2X2 U14 ( .A(A[13]), .B(B[13]), .Y(n135) );
  OR2X2 U15 ( .A(A[6]), .B(B[6]), .Y(n6) );
  INVX8 U16 ( .A(n145), .Y(n40) );
  NAND2X2 U17 ( .A(A[2]), .B(B[2]), .Y(n49) );
  CLKINVX8 U18 ( .A(n135), .Y(n106) );
  NAND2X1 U19 ( .A(n135), .B(n104), .Y(n17) );
  OAI2BB1X4 U20 ( .A0N(n40), .A1N(n57), .B0(n146), .Y(n20) );
  NAND2X2 U21 ( .A(n124), .B(n125), .Y(n33) );
  OAI21X4 U22 ( .A0(n106), .A1(n21), .B0(n104), .Y(n129) );
  XOR2X4 U23 ( .A(n139), .B(n17), .Y(SUM[13]) );
  NAND2X2 U24 ( .A(n115), .B(n50), .Y(n138) );
  INVX1 U25 ( .A(n129), .Y(n134) );
  INVX1 U26 ( .A(n58), .Y(n178) );
  INVX4 U27 ( .A(n121), .Y(n172) );
  BUFX4 U28 ( .A(n116), .Y(n50) );
  NOR2X2 U29 ( .A(n30), .B(n149), .Y(n148) );
  INVX1 U30 ( .A(n111), .Y(n98) );
  INVX1 U31 ( .A(n30), .Y(n59) );
  NAND2X2 U32 ( .A(B[1]), .B(A[1]), .Y(n87) );
  INVX1 U33 ( .A(n102), .Y(n27) );
  AND2X2 U34 ( .A(n99), .B(n111), .Y(n34) );
  BUFX8 U35 ( .A(n158), .Y(n7) );
  NOR2BX2 U36 ( .AN(n68), .B(n72), .Y(n74) );
  NAND3X4 U37 ( .A(n170), .B(n123), .C(n82), .Y(n43) );
  INVXL U38 ( .A(n70), .Y(n72) );
  AND2X2 U39 ( .A(n162), .B(n11), .Y(n8) );
  AND3X4 U40 ( .A(n13), .B(n123), .C(n82), .Y(n9) );
  AND2X2 U41 ( .A(n32), .B(n127), .Y(n10) );
  OR2X4 U42 ( .A(n52), .B(n150), .Y(n11) );
  INVX8 U43 ( .A(n127), .Y(n105) );
  AOI21X1 U44 ( .A0(n129), .A1(n127), .B0(n102), .Y(n124) );
  OAI21X2 U45 ( .A0(n97), .A1(n98), .B0(n99), .Y(n96) );
  OR2X4 U46 ( .A(n24), .B(n51), .Y(n12) );
  NOR2X4 U47 ( .A(n172), .B(n171), .Y(n13) );
  INVX8 U48 ( .A(n122), .Y(n171) );
  NAND2X2 U49 ( .A(A[3]), .B(n5), .Y(n82) );
  NAND2X2 U50 ( .A(A[4]), .B(B[4]), .Y(n14) );
  NOR2BX4 U51 ( .AN(n23), .B(n14), .Y(n180) );
  NAND2BX4 U52 ( .AN(n15), .B(n176), .Y(n108) );
  NAND2X4 U53 ( .A(n154), .B(n71), .Y(n15) );
  NAND2X1 U54 ( .A(B[13]), .B(A[13]), .Y(n104) );
  INVXL U55 ( .A(n19), .Y(n16) );
  NAND2X2 U56 ( .A(n12), .B(n71), .Y(n19) );
  NAND2X4 U57 ( .A(B[4]), .B(A[4]), .Y(n159) );
  CLKINVX8 U58 ( .A(n4), .Y(SUM[4]) );
  NAND3X4 U59 ( .A(n85), .B(n81), .C(n175), .Y(n123) );
  NAND2X4 U60 ( .A(n3), .B(n179), .Y(n118) );
  AND2X1 U61 ( .A(n52), .B(n53), .Y(n48) );
  BUFX16 U62 ( .A(B[5]), .Y(n24) );
  NAND3BX4 U63 ( .AN(n149), .B(n54), .C(n165), .Y(n164) );
  DLY1X1 U64 ( .A(n65), .Y(n18) );
  NAND4BX4 U65 ( .AN(n19), .B(n35), .C(n28), .D(n153), .Y(n57) );
  INVX8 U66 ( .A(n152), .Y(n64) );
  AOI2BB1X2 U67 ( .A0N(B[3]), .A1N(A[3]), .B0(n90), .Y(n175) );
  INVX1 U68 ( .A(n85), .Y(n89) );
  INVX8 U69 ( .A(n143), .Y(n137) );
  NAND2X4 U70 ( .A(n10), .B(n128), .Y(n125) );
  CLKINVX3 U71 ( .A(n126), .Y(n32) );
  OAI21X1 U72 ( .A0(n5), .A1(A[3]), .B0(n82), .Y(n77) );
  INVX8 U73 ( .A(n9), .Y(n35) );
  INVX8 U74 ( .A(n66), .Y(n63) );
  NAND2X2 U75 ( .A(A[8]), .B(B[8]), .Y(n58) );
  BUFX20 U76 ( .A(A[5]), .Y(n51) );
  OR2X4 U77 ( .A(A[12]), .B(B[12]), .Y(n136) );
  INVX8 U78 ( .A(n107), .Y(n146) );
  BUFX8 U79 ( .A(n103), .Y(n21) );
  NAND2XL U80 ( .A(B[12]), .B(A[12]), .Y(n103) );
  INVX4 U81 ( .A(n174), .Y(n173) );
  AND2X4 U82 ( .A(n78), .B(n79), .Y(n45) );
  NAND2XL U83 ( .A(n123), .B(n82), .Y(n119) );
  AND2X1 U84 ( .A(n2), .B(n16), .Y(n22) );
  OR2X4 U85 ( .A(B[6]), .B(A[6]), .Y(n23) );
  NOR2X2 U86 ( .A(n105), .B(n106), .Y(n100) );
  NOR2XL U87 ( .A(n106), .B(n112), .Y(n109) );
  AND2X1 U88 ( .A(n62), .B(n153), .Y(n61) );
  NAND3X4 U89 ( .A(n43), .B(n70), .C(n71), .Y(n69) );
  AOI21X4 U90 ( .A0(n7), .A1(n157), .B0(n181), .Y(n155) );
  INVX4 U91 ( .A(n71), .Y(n75) );
  NAND2X2 U92 ( .A(n118), .B(n153), .Y(n56) );
  OAI2BB1X4 U93 ( .A0N(n46), .A1N(n47), .B0(n160), .Y(n25) );
  NOR2BX2 U94 ( .AN(n65), .B(n64), .Y(n67) );
  NOR2X4 U95 ( .A(B[3]), .B(A[3]), .Y(n174) );
  INVX3 U96 ( .A(n130), .Y(n102) );
  NAND2X4 U97 ( .A(n62), .B(n65), .Y(n181) );
  AND2X4 U98 ( .A(n50), .B(n161), .Y(n44) );
  NAND2X2 U99 ( .A(A[6]), .B(B[6]), .Y(n65) );
  OR2X4 U100 ( .A(A[11]), .B(B[11]), .Y(n161) );
  NAND2X2 U101 ( .A(B[10]), .B(A[10]), .Y(n162) );
  NOR2BX2 U102 ( .AN(n21), .B(n112), .Y(n144) );
  INVX2 U103 ( .A(n21), .Y(n142) );
  NAND2X4 U104 ( .A(n164), .B(n8), .Y(n163) );
  NAND3X4 U105 ( .A(n20), .B(n115), .C(n50), .Y(n128) );
  OAI21X4 U106 ( .A0(n63), .A1(n29), .B0(n18), .Y(n60) );
  NAND2BX2 U107 ( .AN(n159), .B(n70), .Y(n42) );
  NOR2X4 U108 ( .A(A[8]), .B(B[8]), .Y(n30) );
  OAI21X4 U109 ( .A0(n112), .A1(n25), .B0(n141), .Y(n140) );
  OR2X4 U110 ( .A(A[9]), .B(B[9]), .Y(n53) );
  OR2X2 U111 ( .A(A[14]), .B(B[14]), .Y(n127) );
  NAND2X1 U112 ( .A(n24), .B(n51), .Y(n68) );
  NAND3X4 U113 ( .A(n42), .B(n69), .C(n68), .Y(n66) );
  NOR2X2 U114 ( .A(n31), .B(n30), .Y(n177) );
  AOI21XL U115 ( .A0(n117), .A1(n56), .B0(n107), .Y(n113) );
  NAND2BX4 U116 ( .AN(n51), .B(n1), .Y(n158) );
  OR2X4 U117 ( .A(n174), .B(n49), .Y(n121) );
  NOR2BX2 U118 ( .AN(n87), .B(n89), .Y(n88) );
  XOR2X4 U119 ( .A(n86), .B(n88), .Y(SUM[1]) );
  NAND2XL U120 ( .A(n121), .B(n122), .Y(n120) );
  NAND2X4 U121 ( .A(B[7]), .B(A[7]), .Y(n62) );
  INVX8 U122 ( .A(n136), .Y(n112) );
  OR2X4 U123 ( .A(A[2]), .B(B[2]), .Y(n81) );
  OAI2BB1X4 U124 ( .A0N(n85), .A1N(n86), .B0(n87), .Y(n80) );
  NAND2X1 U125 ( .A(n66), .B(n36), .Y(n37) );
  XOR2X4 U126 ( .A(n33), .B(n34), .Y(SUM[15]) );
  OR2X2 U127 ( .A(A[15]), .B(B[15]), .Y(n111) );
  NAND2X2 U128 ( .A(B[15]), .B(A[15]), .Y(n99) );
  INVX4 U129 ( .A(n161), .Y(n151) );
  NOR2X4 U130 ( .A(n150), .B(n151), .Y(n160) );
  NOR2BX1 U131 ( .AN(n162), .B(n150), .Y(n167) );
  OR2X2 U132 ( .A(A[1]), .B(B[1]), .Y(n85) );
  OAI2BB1X4 U133 ( .A0N(n53), .A1N(n54), .B0(n52), .Y(n166) );
  INVX8 U134 ( .A(n53), .Y(n149) );
  XOR2X2 U135 ( .A(n80), .B(n83), .Y(SUM[2]) );
  XOR2X4 U136 ( .A(n77), .B(n45), .Y(SUM[3]) );
  XOR2X4 U137 ( .A(n91), .B(n92), .Y(SUM[16]) );
  OAI21X4 U138 ( .A0(n93), .A1(n94), .B0(n95), .Y(n91) );
  NAND2X1 U139 ( .A(n25), .B(n50), .Y(n114) );
  NOR2X4 U140 ( .A(n159), .B(n64), .Y(n157) );
  NAND3BX4 U141 ( .AN(n108), .B(n59), .C(n35), .Y(n169) );
  OR2X4 U142 ( .A(n149), .B(n58), .Y(n46) );
  XNOR2X4 U143 ( .A(n41), .B(n55), .Y(SUM[8]) );
  AOI2BB1X4 U144 ( .A0N(n112), .A1N(n50), .B0(n142), .Y(n141) );
  XOR2X4 U145 ( .A(n128), .B(n144), .Y(SUM[12]) );
  AOI21X1 U146 ( .A0(n100), .A1(n101), .B0(n102), .Y(n97) );
  AOI21X4 U147 ( .A0(n118), .A1(n177), .B0(n178), .Y(n168) );
  OAI21X2 U148 ( .A0(n75), .A1(n9), .B0(n159), .Y(n73) );
  NAND3BX4 U149 ( .AN(n87), .B(n173), .C(n81), .Y(n122) );
  NOR2X4 U150 ( .A(n150), .B(n151), .Y(n147) );
  INVX8 U151 ( .A(n165), .Y(n150) );
  OR2X4 U152 ( .A(n24), .B(n51), .Y(n154) );
  XOR2X4 U153 ( .A(n73), .B(n74), .Y(SUM[5]) );
  AOI21X4 U154 ( .A0(n180), .A1(n158), .B0(n181), .Y(n179) );
  XOR2X4 U155 ( .A(n26), .B(n48), .Y(SUM[9]) );
  OR2X4 U156 ( .A(n51), .B(n24), .Y(n70) );
  NAND2X4 U157 ( .A(n147), .B(n148), .Y(n107) );
  NOR2X4 U158 ( .A(n137), .B(n138), .Y(n133) );
  OR2X4 U159 ( .A(B[6]), .B(A[6]), .Y(n152) );
  OR2X4 U160 ( .A(A[4]), .B(B[4]), .Y(n71) );
  NAND2X4 U161 ( .A(n136), .B(n135), .Y(n126) );
  NAND2X2 U162 ( .A(n63), .B(n67), .Y(n38) );
  NAND2X4 U163 ( .A(n37), .B(n38), .Y(SUM[6]) );
  INVXL U164 ( .A(n67), .Y(n36) );
  AOI21X4 U165 ( .A0(n155), .A1(n156), .B0(n31), .Y(n145) );
  NOR2BX2 U166 ( .AN(n159), .B(n75), .Y(n76) );
  NAND2X2 U167 ( .A(B[9]), .B(A[9]), .Y(n52) );
  NAND2X2 U168 ( .A(n80), .B(n81), .Y(n79) );
  OAI2BB1X4 U169 ( .A0N(n57), .A1N(n40), .B0(n146), .Y(n143) );
  OR2X4 U170 ( .A(A[10]), .B(B[10]), .Y(n165) );
  NOR2X4 U171 ( .A(n31), .B(n64), .Y(n176) );
  NOR2BX2 U172 ( .AN(n78), .B(n84), .Y(n83) );
  NAND2XL U173 ( .A(n58), .B(n59), .Y(n41) );
  XOR2X4 U174 ( .A(n163), .B(n44), .Y(SUM[11]) );
  NAND2X1 U175 ( .A(n109), .B(n110), .Y(n94) );
  NOR2X1 U176 ( .A(n98), .B(n105), .Y(n110) );
  OAI2BB1X4 U177 ( .A0N(n46), .A1N(n47), .B0(n160), .Y(n115) );
  AND2X2 U178 ( .A(n52), .B(n162), .Y(n47) );
  NAND3XL U179 ( .A(n152), .B(n24), .C(n51), .Y(n156) );
  INVX1 U180 ( .A(n96), .Y(n95) );
  NAND2XL U181 ( .A(n21), .B(n104), .Y(n101) );
  OAI21XL U182 ( .A0(n119), .A1(n120), .B0(n22), .Y(n117) );
  NAND2XL U183 ( .A(B[14]), .B(A[14]), .Y(n130) );
  NAND2XL U184 ( .A(B[2]), .B(A[2]), .Y(n78) );
  INVX1 U185 ( .A(n90), .Y(n86) );
  XOR2X1 U186 ( .A(B[16]), .B(A[16]), .Y(n92) );
  NOR2X1 U187 ( .A(n113), .B(n114), .Y(n93) );
  AND2X2 U188 ( .A(n90), .B(n182), .Y(SUM[0]) );
  OR2X2 U189 ( .A(A[0]), .B(B[0]), .Y(n182) );
  NAND2X1 U190 ( .A(B[0]), .B(A[0]), .Y(n90) );
  NAND2XL U191 ( .A(B[11]), .B(A[11]), .Y(n116) );
  XOR2X4 U192 ( .A(n60), .B(n61), .Y(SUM[7]) );
  XOR2X4 U193 ( .A(n131), .B(n132), .Y(SUM[14]) );
  NOR2BX4 U194 ( .AN(n27), .B(n105), .Y(n132) );
  OAI21X4 U195 ( .A0(n133), .A1(n126), .B0(n134), .Y(n131) );
  AOI21X4 U196 ( .A0(n137), .A1(n136), .B0(n140), .Y(n139) );
  XOR2X4 U197 ( .A(n166), .B(n167), .Y(SUM[10]) );
  NAND2X4 U198 ( .A(n169), .B(n168), .Y(n54) );
  NOR2X4 U199 ( .A(n171), .B(n172), .Y(n170) );
endmodule


module butterfly_DW01_add_128 ( A, B, SUM );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189;

  NAND2X4 U2 ( .A(B[4]), .B(A[4]), .Y(n158) );
  OR2X4 U3 ( .A(A[6]), .B(B[6]), .Y(n172) );
  NAND2X2 U4 ( .A(B[12]), .B(A[12]), .Y(n110) );
  CLKINVX8 U5 ( .A(n153), .Y(n25) );
  AND2X4 U6 ( .A(n56), .B(n60), .Y(n40) );
  OR2X4 U7 ( .A(A[8]), .B(B[8]), .Y(n1) );
  OR2X2 U8 ( .A(A[8]), .B(B[8]), .Y(n46) );
  NAND2X2 U9 ( .A(n169), .B(n2), .Y(n54) );
  NAND3X4 U10 ( .A(n1), .B(n47), .C(n48), .Y(n167) );
  NAND3X2 U11 ( .A(B[4]), .B(A[4]), .C(n171), .Y(n189) );
  NAND3X4 U12 ( .A(n168), .B(n167), .C(n8), .Y(n164) );
  NOR2X2 U13 ( .A(n173), .B(n11), .Y(n163) );
  NAND3BX4 U14 ( .AN(n53), .B(n1), .C(n48), .Y(n177) );
  CLKINVX8 U15 ( .A(n53), .Y(n47) );
  NOR2BX4 U16 ( .AN(n180), .B(n72), .Y(n79) );
  INVX3 U17 ( .A(n80), .Y(n72) );
  XOR2X2 U18 ( .A(n78), .B(n79), .Y(SUM[2]) );
  NAND3X2 U19 ( .A(n70), .B(n69), .C(n68), .Y(n62) );
  INVX2 U20 ( .A(n32), .Y(n68) );
  OAI21X1 U21 ( .A0(n97), .A1(n4), .B0(n107), .Y(n113) );
  CLKINVX3 U22 ( .A(n49), .Y(n187) );
  INVX4 U23 ( .A(n99), .Y(n144) );
  NAND2BX2 U24 ( .AN(n158), .B(n159), .Y(n156) );
  INVXL U25 ( .A(A[11]), .Y(n27) );
  INVX2 U26 ( .A(n44), .Y(n173) );
  OAI2BB1X2 U27 ( .A0N(n81), .A1N(n82), .B0(n83), .Y(n78) );
  BUFX3 U28 ( .A(n76), .Y(n10) );
  INVX1 U29 ( .A(n11), .Y(n14) );
  CLKINVX3 U30 ( .A(n100), .Y(n109) );
  OAI21X2 U31 ( .A0(n88), .A1(n89), .B0(n90), .Y(n87) );
  INVX1 U32 ( .A(n91), .Y(n90) );
  AOI21X1 U33 ( .A0(n93), .A1(n54), .B0(n23), .Y(n88) );
  NAND2BX1 U34 ( .AN(n117), .B(n118), .Y(n116) );
  XOR2X2 U35 ( .A(n48), .B(n73), .Y(SUM[4]) );
  NOR2BX1 U36 ( .AN(n158), .B(n15), .Y(n73) );
  NOR2BX1 U37 ( .AN(n63), .B(n160), .Y(n67) );
  NAND2X1 U38 ( .A(n61), .B(n17), .Y(n59) );
  INVX4 U39 ( .A(n38), .Y(n8) );
  NAND2X4 U40 ( .A(n132), .B(n5), .Y(n92) );
  NAND2X4 U41 ( .A(A[9]), .B(B[9]), .Y(n153) );
  AOI2BB1X4 U42 ( .A0N(B[9]), .A1N(A[9]), .B0(n152), .Y(n151) );
  OAI21X4 U43 ( .A0(A[14]), .A1(B[14]), .B0(n100), .Y(n117) );
  NAND3X4 U44 ( .A(n40), .B(n156), .C(n157), .Y(n18) );
  BUFX12 U45 ( .A(n57), .Y(n2) );
  INVX8 U46 ( .A(n25), .Y(n3) );
  NAND2X4 U47 ( .A(n40), .B(n188), .Y(n186) );
  BUFX4 U48 ( .A(n108), .Y(n4) );
  NAND2XL U49 ( .A(B[13]), .B(A[13]), .Y(n108) );
  INVX8 U50 ( .A(n143), .Y(n5) );
  INVX8 U51 ( .A(n119), .Y(n143) );
  AND2X2 U52 ( .A(n56), .B(n57), .Y(n13) );
  NAND2BX1 U53 ( .AN(n18), .B(n123), .Y(n121) );
  OR2X2 U54 ( .A(n128), .B(n18), .Y(n6) );
  NOR2X2 U55 ( .A(n160), .B(n184), .Y(n159) );
  NOR2X4 U56 ( .A(A[5]), .B(B[5]), .Y(n160) );
  NAND2X2 U57 ( .A(n129), .B(n6), .Y(n127) );
  OAI2BB1X4 U58 ( .A0N(n61), .A1N(n66), .B0(n63), .Y(n64) );
  NAND2X4 U59 ( .A(A[7]), .B(B[7]), .Y(n56) );
  CLKINVX2 U60 ( .A(A[6]), .Y(n20) );
  NAND2X2 U61 ( .A(n99), .B(n5), .Y(n131) );
  NAND2X4 U62 ( .A(n145), .B(n2), .Y(n150) );
  NAND2X4 U63 ( .A(n145), .B(n146), .Y(n140) );
  NAND3X2 U64 ( .A(A[1]), .B(B[1]), .C(n80), .Y(n181) );
  NAND2X1 U65 ( .A(B[1]), .B(A[1]), .Y(n83) );
  NAND2X2 U66 ( .A(n3), .B(n44), .Y(n43) );
  AND2X2 U67 ( .A(A[5]), .B(B[5]), .Y(n37) );
  NAND2X4 U68 ( .A(n70), .B(n68), .Y(n41) );
  OAI21X4 U69 ( .A0(A[7]), .A1(B[7]), .B0(n69), .Y(n182) );
  OAI211X2 U70 ( .A0(n21), .A1(B[6]), .B0(A[5]), .C0(B[5]), .Y(n157) );
  INVX8 U71 ( .A(B[8]), .Y(n29) );
  INVX8 U72 ( .A(n29), .Y(n30) );
  NOR2X4 U73 ( .A(n143), .B(n144), .Y(n142) );
  OR2X2 U74 ( .A(A[5]), .B(B[5]), .Y(n61) );
  XOR2X4 U75 ( .A(n124), .B(n7), .Y(SUM[14]) );
  AND2X1 U76 ( .A(n107), .B(n104), .Y(n7) );
  NOR2X1 U77 ( .A(n41), .B(n19), .Y(n128) );
  OR2X2 U78 ( .A(A[6]), .B(B[6]), .Y(n12) );
  INVX2 U79 ( .A(n81), .Y(n71) );
  AND2X2 U80 ( .A(n99), .B(n2), .Y(n34) );
  INVX2 U81 ( .A(n78), .Y(n77) );
  NOR2X4 U82 ( .A(n154), .B(n3), .Y(n133) );
  INVXL U83 ( .A(n92), .Y(n89) );
  AND2X2 U84 ( .A(n136), .B(n14), .Y(n24) );
  NOR2X2 U85 ( .A(n94), .B(n31), .Y(n129) );
  AND2X4 U86 ( .A(A[8]), .B(n30), .Y(n38) );
  NAND2XL U87 ( .A(n30), .B(A[8]), .Y(n50) );
  NAND2X1 U88 ( .A(B[14]), .B(A[14]), .Y(n107) );
  NAND4BX2 U89 ( .AN(n113), .B(n115), .C(n114), .D(n116), .Y(n111) );
  NAND2X4 U90 ( .A(n38), .B(n151), .Y(n9) );
  NOR2X4 U91 ( .A(A[10]), .B(B[10]), .Y(n11) );
  NOR2X2 U92 ( .A(B[10]), .B(A[10]), .Y(n154) );
  NAND3BX2 U93 ( .AN(n38), .B(n168), .C(n45), .Y(n42) );
  NAND4X4 U94 ( .A(n10), .B(n179), .C(n180), .D(n181), .Y(n70) );
  NAND2X1 U95 ( .A(B[3]), .B(A[3]), .Y(n76) );
  INVX4 U96 ( .A(n20), .Y(n21) );
  AOI2BB1X2 U97 ( .A0N(n21), .A1N(B[6]), .B0(n189), .Y(n185) );
  NOR2XL U98 ( .A(A[4]), .B(B[4]), .Y(n15) );
  NOR2X4 U99 ( .A(B[10]), .B(A[10]), .Y(n152) );
  DLY1X1 U100 ( .A(n70), .Y(n16) );
  NOR2BX2 U101 ( .AN(n136), .B(n166), .Y(n165) );
  NAND2X4 U102 ( .A(A[10]), .B(B[10]), .Y(n136) );
  NAND3X4 U103 ( .A(n171), .B(n12), .C(n170), .Y(n95) );
  INVX3 U104 ( .A(n184), .Y(n17) );
  NAND2BX2 U105 ( .AN(n182), .B(n183), .Y(n19) );
  NOR2BX2 U106 ( .AN(n25), .B(n11), .Y(n166) );
  OAI21X1 U107 ( .A0(A[12]), .A1(B[12]), .B0(n2), .Y(n130) );
  NOR2X4 U108 ( .A(A[6]), .B(B[6]), .Y(n184) );
  NAND2BX2 U109 ( .AN(n131), .B(n132), .Y(n126) );
  NAND2BX4 U110 ( .AN(n49), .B(n169), .Y(n168) );
  NOR2BX2 U111 ( .AN(n110), .B(n144), .Y(n149) );
  AND2X2 U112 ( .A(n60), .B(n17), .Y(n65) );
  NOR2X4 U113 ( .A(n147), .B(n18), .Y(n139) );
  NOR2X2 U114 ( .A(n94), .B(n117), .Y(n122) );
  CLKINVX8 U115 ( .A(n94), .Y(n145) );
  AND2X1 U116 ( .A(n50), .B(n1), .Y(n52) );
  BUFX8 U117 ( .A(n134), .Y(n22) );
  NAND2XL U118 ( .A(B[11]), .B(A[11]), .Y(n134) );
  INVXL U119 ( .A(n145), .Y(n23) );
  NAND2X2 U120 ( .A(B[2]), .B(A[2]), .Y(n180) );
  NAND4BX4 U121 ( .AN(n133), .B(n9), .C(n22), .D(n136), .Y(n132) );
  AND2X2 U122 ( .A(B[4]), .B(A[4]), .Y(n170) );
  NAND3X4 U123 ( .A(n176), .B(n177), .C(n8), .Y(n175) );
  XOR2X4 U124 ( .A(n74), .B(n75), .Y(SUM[3]) );
  XOR2X4 U125 ( .A(n33), .B(n24), .Y(SUM[10]) );
  NAND3X1 U126 ( .A(n172), .B(B[5]), .C(A[5]), .Y(n188) );
  NAND4X4 U127 ( .A(n95), .B(n26), .C(n60), .D(n56), .Y(n169) );
  NAND2X2 U128 ( .A(n172), .B(n37), .Y(n26) );
  XOR2X4 U129 ( .A(n82), .B(n84), .Y(SUM[1]) );
  NOR2BX4 U130 ( .AN(n83), .B(n71), .Y(n84) );
  OAI21X4 U131 ( .A0(n150), .A1(n139), .B0(n92), .Y(n148) );
  AOI21X4 U132 ( .A0(n120), .A1(n142), .B0(n118), .Y(n141) );
  NAND2X4 U133 ( .A(n175), .B(n44), .Y(n174) );
  AOI21X2 U134 ( .A0(B[11]), .A1(n28), .B0(n143), .Y(n162) );
  NOR2X1 U135 ( .A(n109), .B(n110), .Y(n105) );
  AND2X4 U136 ( .A(n86), .B(n87), .Y(n35) );
  NAND2X1 U137 ( .A(n107), .B(n4), .Y(n106) );
  INVX2 U138 ( .A(n27), .Y(n28) );
  NAND2X4 U139 ( .A(n174), .B(n3), .Y(n33) );
  NAND3X2 U140 ( .A(n122), .B(n121), .C(n34), .Y(n114) );
  OAI21X4 U141 ( .A0(n77), .A1(n72), .B0(n180), .Y(n74) );
  NAND4BX1 U142 ( .AN(n97), .B(n98), .C(n99), .D(n100), .Y(n91) );
  NAND3X2 U143 ( .A(n127), .B(n126), .C(n110), .Y(n125) );
  NAND4BX2 U144 ( .AN(n117), .B(n120), .C(n99), .D(n5), .Y(n115) );
  OAI21X4 U145 ( .A0(n185), .A1(n186), .B0(n187), .Y(n176) );
  INVX4 U146 ( .A(n123), .Y(n147) );
  OAI21X4 U147 ( .A0(n30), .A1(A[8]), .B0(n57), .Y(n49) );
  NAND2X2 U148 ( .A(n103), .B(n98), .Y(n112) );
  OAI21X2 U149 ( .A0(n101), .A1(n102), .B0(n103), .Y(n96) );
  NOR2X2 U150 ( .A(n105), .B(n106), .Y(n101) );
  XNOR2X4 U151 ( .A(n111), .B(n112), .Y(SUM[15]) );
  NAND3X1 U152 ( .A(n46), .B(n47), .C(n48), .Y(n45) );
  NAND3BX2 U153 ( .AN(n85), .B(n80), .C(n81), .Y(n179) );
  NAND2X4 U154 ( .A(n151), .B(n38), .Y(n135) );
  INVX4 U155 ( .A(n104), .Y(n97) );
  NAND2X1 U156 ( .A(n104), .B(n98), .Y(n102) );
  OR2X2 U157 ( .A(A[14]), .B(B[14]), .Y(n104) );
  XOR2X4 U158 ( .A(n148), .B(n149), .Y(SUM[12]) );
  NOR2X4 U159 ( .A(n184), .B(n160), .Y(n183) );
  XOR2X4 U160 ( .A(n161), .B(n162), .Y(SUM[11]) );
  OR2X4 U161 ( .A(B[11]), .B(A[11]), .Y(n119) );
  OAI21X4 U162 ( .A0(n58), .A1(n59), .B0(n60), .Y(n55) );
  NAND2X4 U163 ( .A(B[6]), .B(A[6]), .Y(n60) );
  NAND4BX4 U164 ( .AN(n133), .B(n135), .C(n22), .D(n136), .Y(n120) );
  NOR2X2 U165 ( .A(A[3]), .B(B[3]), .Y(n32) );
  OR2X4 U166 ( .A(B[9]), .B(A[9]), .Y(n44) );
  OAI2BB1X4 U167 ( .A0N(n163), .A1N(n164), .B0(n165), .Y(n161) );
  XOR2X4 U168 ( .A(n64), .B(n65), .Y(SUM[6]) );
  OR2X4 U169 ( .A(A[15]), .B(B[15]), .Y(n98) );
  OR2X4 U170 ( .A(A[5]), .B(B[5]), .Y(n171) );
  NAND4X4 U171 ( .A(n119), .B(n155), .C(n44), .D(n46), .Y(n94) );
  XOR2X4 U172 ( .A(n55), .B(n13), .Y(SUM[7]) );
  NAND2X4 U173 ( .A(B[5]), .B(A[5]), .Y(n63) );
  OR2X4 U174 ( .A(A[10]), .B(B[10]), .Y(n155) );
  OR2X4 U175 ( .A(A[1]), .B(B[1]), .Y(n81) );
  NAND2BX4 U176 ( .AN(n19), .B(n48), .Y(n123) );
  INVX8 U177 ( .A(n41), .Y(n48) );
  OR2X4 U178 ( .A(A[7]), .B(B[7]), .Y(n57) );
  XOR2X4 U179 ( .A(n52), .B(n51), .Y(SUM[8]) );
  OR2X4 U180 ( .A(A[2]), .B(B[2]), .Y(n80) );
  NAND2X2 U181 ( .A(n158), .B(n62), .Y(n66) );
  BUFX4 U182 ( .A(n130), .Y(n31) );
  OR2X4 U183 ( .A(A[4]), .B(B[4]), .Y(n69) );
  OR2X4 U184 ( .A(A[13]), .B(B[13]), .Y(n100) );
  NOR2BX2 U185 ( .AN(n10), .B(n32), .Y(n75) );
  INVX4 U186 ( .A(n110), .Y(n118) );
  OAI21X2 U187 ( .A0(n41), .A1(n19), .B0(n54), .Y(n51) );
  XNOR2X4 U188 ( .A(n42), .B(n43), .Y(SUM[9]) );
  CLKINVX3 U189 ( .A(n31), .Y(n146) );
  NAND2XL U190 ( .A(B[15]), .B(A[15]), .Y(n103) );
  XOR2X2 U191 ( .A(n35), .B(n36), .Y(SUM[16]) );
  XNOR2X1 U192 ( .A(B[16]), .B(A[16]), .Y(n36) );
  XOR2X2 U193 ( .A(n66), .B(n67), .Y(SUM[5]) );
  AND2X2 U194 ( .A(n39), .B(n62), .Y(n58) );
  AND2X2 U195 ( .A(n63), .B(n158), .Y(n39) );
  INVX1 U196 ( .A(n96), .Y(n86) );
  NAND3XL U197 ( .A(n47), .B(n16), .C(n68), .Y(n93) );
  INVX1 U198 ( .A(n85), .Y(n82) );
  AND2X2 U199 ( .A(n85), .B(n178), .Y(SUM[0]) );
  OR2X2 U200 ( .A(A[0]), .B(B[0]), .Y(n178) );
  NAND2X1 U201 ( .A(B[0]), .B(A[0]), .Y(n85) );
  OAI2BB1X4 U202 ( .A0N(n100), .A1N(n125), .B0(n4), .Y(n124) );
  XOR2X4 U203 ( .A(n137), .B(n138), .Y(SUM[13]) );
  NOR2BX4 U204 ( .AN(n4), .B(n109), .Y(n138) );
  OAI21X4 U205 ( .A0(n139), .A1(n140), .B0(n141), .Y(n137) );
  OR2X4 U206 ( .A(A[12]), .B(B[12]), .Y(n99) );
  NAND2BX4 U207 ( .AN(n182), .B(n183), .Y(n53) );
endmodule


module butterfly_DW01_add_129 ( A, B, SUM );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216;

  OAI21X2 U2 ( .A0(n115), .A1(n116), .B0(n117), .Y(n113) );
  NAND2BX4 U3 ( .AN(n1), .B(n186), .Y(n60) );
  CLKINVX20 U4 ( .A(n185), .Y(n1) );
  BUFX16 U5 ( .A(B[5]), .Y(n69) );
  BUFX1 U6 ( .A(n122), .Y(n30) );
  INVXL U7 ( .A(n33), .Y(n2) );
  AND2X2 U8 ( .A(B[4]), .B(A[4]), .Y(n215) );
  NAND2X4 U9 ( .A(B[9]), .B(A[9]), .Y(n184) );
  NAND2BX4 U10 ( .AN(B[3]), .B(n3), .Y(n33) );
  CLKINVX20 U11 ( .A(A[3]), .Y(n3) );
  NAND2X4 U12 ( .A(B[7]), .B(A[7]), .Y(n14) );
  NOR2X4 U13 ( .A(n103), .B(n104), .Y(n207) );
  NAND3X4 U14 ( .A(n72), .B(n7), .C(n73), .Y(n63) );
  NAND2BX4 U15 ( .AN(n75), .B(n15), .Y(n72) );
  XOR2X4 U16 ( .A(n6), .B(n77), .Y(SUM[8]) );
  NOR2X2 U17 ( .A(n136), .B(n142), .Y(n176) );
  INVXL U18 ( .A(A[11]), .Y(n22) );
  INVX4 U19 ( .A(n71), .Y(n8) );
  NAND2X2 U20 ( .A(n137), .B(n138), .Y(n53) );
  NAND2X2 U21 ( .A(n54), .B(n139), .Y(n15) );
  NAND2BX2 U22 ( .AN(n202), .B(n71), .Y(n40) );
  AND2X2 U23 ( .A(n179), .B(n89), .Y(n84) );
  INVX2 U24 ( .A(n90), .Y(n82) );
  NAND2X2 U25 ( .A(n144), .B(n145), .Y(n19) );
  NOR2BX2 U26 ( .AN(n89), .B(n36), .Y(n99) );
  INVX2 U27 ( .A(n97), .Y(n55) );
  NOR2X2 U28 ( .A(A[5]), .B(n69), .Y(n12) );
  INVX4 U29 ( .A(n165), .Y(n158) );
  NOR2X1 U30 ( .A(n127), .B(n128), .Y(n124) );
  INVX1 U31 ( .A(n185), .Y(n35) );
  NAND2X1 U32 ( .A(B[1]), .B(A[1]), .Y(n110) );
  INVX1 U33 ( .A(A[2]), .Y(n5) );
  AND2X2 U34 ( .A(n69), .B(A[5]), .Y(n17) );
  INVX1 U35 ( .A(n170), .Y(n21) );
  NOR2X1 U36 ( .A(n131), .B(n132), .Y(n115) );
  OAI21X1 U37 ( .A0(n140), .A1(n13), .B0(n66), .Y(n135) );
  CLKINVX3 U38 ( .A(n40), .Y(n64) );
  INVX1 U39 ( .A(n34), .Y(n38) );
  NAND2X2 U40 ( .A(n78), .B(n79), .Y(n77) );
  INVX4 U41 ( .A(n208), .Y(n104) );
  OR2X2 U42 ( .A(A[5]), .B(n69), .Y(n144) );
  CLKINVX3 U43 ( .A(n24), .Y(n59) );
  INVX1 U44 ( .A(A[5]), .Y(n70) );
  NAND2X2 U45 ( .A(A[3]), .B(B[3]), .Y(n102) );
  INVX2 U46 ( .A(n96), .Y(n18) );
  OR2X2 U47 ( .A(A[4]), .B(B[4]), .Y(n96) );
  OAI2BB1X4 U48 ( .A0N(n33), .A1N(n4), .B0(n146), .Y(n141) );
  CLKINVX3 U49 ( .A(n105), .Y(n4) );
  NAND2BX4 U50 ( .AN(B[2]), .B(n5), .Y(n208) );
  OAI2BB1X4 U51 ( .A0N(n106), .A1N(n208), .B0(n105), .Y(n100) );
  OAI2BB1X1 U52 ( .A0N(n108), .A1N(n109), .B0(n110), .Y(n106) );
  AOI21X4 U53 ( .A0(n164), .A1(n159), .B0(n158), .Y(n163) );
  AND2X1 U54 ( .A(n73), .B(n80), .Y(n6) );
  INVX8 U55 ( .A(n42), .Y(n26) );
  NAND4BX4 U56 ( .AN(n9), .B(n50), .C(n205), .D(n26), .Y(n7) );
  NAND4BX2 U57 ( .AN(n9), .B(n50), .C(n205), .D(n26), .Y(n74) );
  NAND2X4 U58 ( .A(n91), .B(n25), .Y(n9) );
  NAND2BX4 U59 ( .AN(B[3]), .B(n10), .Y(n209) );
  CLKINVX20 U60 ( .A(A[3]), .Y(n10) );
  XNOR2X4 U61 ( .A(n93), .B(n11), .Y(SUM[6]) );
  AND2X1 U62 ( .A(n52), .B(n90), .Y(n11) );
  INVX2 U63 ( .A(n166), .Y(n127) );
  AND2X1 U64 ( .A(n59), .B(n122), .Y(n39) );
  NAND3X4 U65 ( .A(n33), .B(n208), .C(n210), .Y(n146) );
  NAND3BX4 U66 ( .AN(n12), .B(n52), .C(n215), .Y(n214) );
  OR2X4 U67 ( .A(n189), .B(n35), .Y(n200) );
  NOR2BX4 U68 ( .AN(n71), .B(n189), .Y(n188) );
  INVX4 U69 ( .A(n41), .Y(n71) );
  DLY1X1 U70 ( .A(n141), .Y(n13) );
  AND2X2 U71 ( .A(B[11]), .B(A[11]), .Y(n20) );
  NOR2X4 U72 ( .A(n142), .B(n70), .Y(n198) );
  INVX8 U73 ( .A(n20), .Y(n134) );
  NAND3BX4 U74 ( .AN(n195), .B(n16), .C(n215), .Y(n139) );
  NAND2BX4 U75 ( .AN(n48), .B(n207), .Y(n147) );
  OR2X4 U76 ( .A(A[6]), .B(B[6]), .Y(n16) );
  NOR2BX2 U77 ( .AN(n29), .B(n194), .Y(n193) );
  NAND4BBX4 U78 ( .AN(n19), .BN(n18), .C(n50), .D(n51), .Y(n79) );
  NAND2X2 U79 ( .A(n159), .B(n122), .Y(n23) );
  NAND2X2 U80 ( .A(B[2]), .B(A[2]), .Y(n105) );
  AOI21X4 U81 ( .A0(n198), .A1(n69), .B0(n199), .Y(n197) );
  XNOR2X4 U82 ( .A(n169), .B(n21), .Y(SUM[13]) );
  NAND3X1 U83 ( .A(A[5]), .B(n16), .C(n69), .Y(n137) );
  NAND2BX2 U84 ( .AN(B[11]), .B(n22), .Y(n32) );
  OAI21X4 U85 ( .A0(n195), .A1(n196), .B0(n197), .Y(n192) );
  CLKINVX8 U86 ( .A(n164), .Y(n44) );
  AND2X4 U87 ( .A(B[14]), .B(A[14]), .Y(n24) );
  OR2X4 U88 ( .A(A[8]), .B(B[8]), .Y(n25) );
  NOR2X4 U89 ( .A(A[5]), .B(n69), .Y(n42) );
  AND2X2 U90 ( .A(n38), .B(n28), .Y(n45) );
  NAND2X4 U91 ( .A(n27), .B(n182), .Y(n133) );
  AND2X4 U92 ( .A(n181), .B(n180), .Y(n27) );
  OR2X4 U93 ( .A(A[7]), .B(B[7]), .Y(n28) );
  OR2X4 U94 ( .A(A[7]), .B(B[7]), .Y(n29) );
  NOR2BX2 U95 ( .AN(n126), .B(n127), .Y(n170) );
  NAND2XL U96 ( .A(n59), .B(n126), .Y(n125) );
  NAND2X4 U97 ( .A(B[13]), .B(A[13]), .Y(n126) );
  CLKINVX2 U98 ( .A(n180), .Y(n189) );
  NAND3BX2 U99 ( .AN(n129), .B(n167), .C(n159), .Y(n162) );
  CLKINVX3 U100 ( .A(n29), .Y(n136) );
  AND2X1 U101 ( .A(B[12]), .B(A[12]), .Y(n31) );
  OR2X2 U102 ( .A(B[11]), .B(A[11]), .Y(n181) );
  AND2X4 U103 ( .A(B[7]), .B(A[7]), .Y(n34) );
  NOR2X2 U104 ( .A(A[4]), .B(B[4]), .Y(n36) );
  BUFX12 U105 ( .A(n130), .Y(n37) );
  AND2X2 U106 ( .A(n110), .B(n108), .Y(n111) );
  XOR2X4 U107 ( .A(n160), .B(n39), .Y(SUM[14]) );
  NAND2X1 U108 ( .A(n128), .B(n37), .Y(n174) );
  NOR2BX2 U109 ( .AN(n37), .B(n129), .Y(n171) );
  NAND4BXL U110 ( .AN(n127), .B(n37), .C(n30), .D(n123), .Y(n116) );
  NOR2X4 U111 ( .A(A[5]), .B(n69), .Y(n195) );
  CLKINVX2 U112 ( .A(n184), .Y(n202) );
  OR2X4 U113 ( .A(A[5]), .B(n69), .Y(n87) );
  NOR2X4 U114 ( .A(A[9]), .B(B[9]), .Y(n41) );
  AOI21X4 U115 ( .A0(n85), .A1(n84), .B0(n86), .Y(n83) );
  AND2X4 U116 ( .A(n14), .B(n90), .Y(n138) );
  INVX2 U117 ( .A(n122), .Y(n156) );
  XOR2X2 U118 ( .A(n106), .B(n107), .Y(SUM[2]) );
  AOI21XL U119 ( .A0(n135), .A1(n78), .B0(n129), .Y(n131) );
  AOI21X4 U120 ( .A0(n204), .A1(n74), .B0(n8), .Y(n203) );
  NAND2X2 U121 ( .A(n30), .B(n123), .Y(n120) );
  NOR2BX4 U122 ( .AN(n121), .B(n150), .Y(n149) );
  NOR2X4 U123 ( .A(n44), .B(n23), .Y(n154) );
  INVX1 U124 ( .A(n80), .Y(n194) );
  NAND2X2 U125 ( .A(B[4]), .B(A[4]), .Y(n89) );
  NOR2X4 U126 ( .A(n103), .B(n104), .Y(n43) );
  INVX8 U127 ( .A(n133), .Y(n164) );
  NAND2X4 U128 ( .A(n90), .B(n92), .Y(n199) );
  OR2X4 U129 ( .A(A[14]), .B(B[14]), .Y(n122) );
  NAND2X4 U130 ( .A(n187), .B(n188), .Y(n186) );
  NAND2X4 U131 ( .A(n69), .B(A[5]), .Y(n179) );
  AOI21X4 U132 ( .A0(n176), .A1(n177), .B0(n34), .Y(n175) );
  INVX4 U133 ( .A(n49), .Y(SUM[4]) );
  XNOR2X4 U134 ( .A(n81), .B(n45), .Y(SUM[7]) );
  NAND2X4 U135 ( .A(n25), .B(n28), .Y(n75) );
  AND2X2 U136 ( .A(n32), .B(n134), .Y(n61) );
  NAND2X4 U137 ( .A(n192), .B(n193), .Y(n190) );
  AND3X4 U138 ( .A(n69), .B(n51), .C(A[5]), .Y(n216) );
  NAND3X1 U139 ( .A(B[4]), .B(A[4]), .C(n52), .Y(n196) );
  NAND3X4 U140 ( .A(n7), .B(n190), .C(n191), .Y(n187) );
  NAND2X4 U141 ( .A(n46), .B(n102), .Y(n95) );
  NOR2BX4 U142 ( .AN(n147), .B(n141), .Y(n46) );
  NAND2BX4 U143 ( .AN(n48), .B(n43), .Y(n47) );
  NAND2X2 U144 ( .A(n108), .B(n109), .Y(n48) );
  NAND2X4 U145 ( .A(n47), .B(n102), .Y(n206) );
  NAND2X1 U146 ( .A(A[8]), .B(B[8]), .Y(n183) );
  XNOR2X2 U147 ( .A(n50), .B(n99), .Y(n49) );
  AOI21X4 U148 ( .A0(n213), .A1(n214), .B0(n75), .Y(n212) );
  INVX8 U149 ( .A(n209), .Y(n103) );
  AOI21X4 U150 ( .A0(n95), .A1(n96), .B0(n215), .Y(n98) );
  OAI211X2 U151 ( .A0(n195), .A1(n178), .B0(n179), .C0(n90), .Y(n177) );
  NAND2X2 U152 ( .A(n26), .B(n16), .Y(n86) );
  XOR2X4 U153 ( .A(n63), .B(n64), .Y(SUM[9]) );
  OAI21X2 U154 ( .A0(n151), .A1(n152), .B0(n153), .Y(n148) );
  AOI21X4 U155 ( .A0(n173), .A1(n37), .B0(n31), .Y(n172) );
  NOR2BX1 U156 ( .AN(n105), .B(n104), .Y(n107) );
  OAI2BB1X4 U157 ( .A0N(n171), .A1N(n167), .B0(n172), .Y(n169) );
  NOR2X4 U158 ( .A(n155), .B(n154), .Y(n153) );
  OR2X2 U159 ( .A(A[15]), .B(B[15]), .Y(n123) );
  XOR2X4 U160 ( .A(n113), .B(n114), .Y(SUM[16]) );
  NAND2X2 U161 ( .A(n55), .B(n98), .Y(n58) );
  NAND2X4 U162 ( .A(n89), .B(n85), .Y(n94) );
  NOR2X4 U163 ( .A(n199), .B(n216), .Y(n213) );
  INVX2 U164 ( .A(n123), .Y(n150) );
  NAND2X4 U165 ( .A(B[6]), .B(A[6]), .Y(n90) );
  OR2X4 U166 ( .A(n206), .B(n141), .Y(n50) );
  XOR2X4 U167 ( .A(n148), .B(n149), .Y(SUM[15]) );
  NAND2X4 U168 ( .A(n97), .B(n56), .Y(n57) );
  INVX4 U169 ( .A(n98), .Y(n56) );
  NAND2X4 U170 ( .A(n175), .B(n79), .Y(n167) );
  NOR2X4 U171 ( .A(n203), .B(n202), .Y(n201) );
  OAI2BB1X4 U172 ( .A0N(n128), .A1N(n126), .B0(n166), .Y(n165) );
  NAND2X4 U173 ( .A(B[12]), .B(A[12]), .Y(n128) );
  OAI22X4 U174 ( .A0(n151), .A1(n134), .B0(n156), .B1(n157), .Y(n155) );
  AND3X4 U175 ( .A(n152), .B(n44), .C(n134), .Y(n62) );
  NAND2X4 U176 ( .A(n134), .B(n133), .Y(n173) );
  NOR2X4 U177 ( .A(n83), .B(n82), .Y(n81) );
  CLKINVX3 U178 ( .A(n118), .Y(n117) );
  OAI21X2 U179 ( .A0(n119), .A1(n120), .B0(n121), .Y(n118) );
  NAND2X2 U180 ( .A(B[10]), .B(A[10]), .Y(n185) );
  OR2X4 U181 ( .A(A[6]), .B(B[6]), .Y(n51) );
  OR2X4 U182 ( .A(A[6]), .B(B[6]), .Y(n52) );
  NOR2X4 U183 ( .A(n24), .B(n158), .Y(n157) );
  NAND4BX4 U184 ( .AN(n8), .B(n32), .C(n180), .D(n80), .Y(n129) );
  OR2X4 U185 ( .A(B[10]), .B(A[10]), .Y(n180) );
  NAND2X4 U186 ( .A(n87), .B(n179), .Y(n97) );
  NAND2XL U187 ( .A(n44), .B(n134), .Y(n132) );
  INVX8 U188 ( .A(n88), .Y(n142) );
  NAND2X4 U189 ( .A(B[8]), .B(A[8]), .Y(n73) );
  NOR2X4 U190 ( .A(n212), .B(n211), .Y(n204) );
  XOR2X4 U191 ( .A(n100), .B(n101), .Y(SUM[3]) );
  NAND2X4 U192 ( .A(n159), .B(n122), .Y(n151) );
  INVX8 U193 ( .A(n168), .Y(n159) );
  NAND2X4 U194 ( .A(n95), .B(n96), .Y(n85) );
  NAND2X4 U195 ( .A(n54), .B(n139), .Y(n76) );
  INVX4 U196 ( .A(n53), .Y(n54) );
  NAND2BX4 U197 ( .AN(n136), .B(n76), .Y(n78) );
  NAND2X4 U198 ( .A(n57), .B(n58), .Y(SUM[5]) );
  XOR2X4 U199 ( .A(n201), .B(n200), .Y(SUM[10]) );
  XOR2X4 U200 ( .A(n60), .B(n61), .Y(SUM[11]) );
  OR2XL U201 ( .A(n142), .B(n36), .Y(n68) );
  NAND2XL U202 ( .A(B[0]), .B(A[0]), .Y(n112) );
  NAND2BX4 U203 ( .AN(n129), .B(n167), .Y(n152) );
  NOR2X2 U204 ( .A(n67), .B(n68), .Y(n66) );
  NOR2X4 U205 ( .A(n36), .B(n142), .Y(n205) );
  XOR2X4 U206 ( .A(n174), .B(n62), .Y(SUM[12]) );
  NAND2X4 U207 ( .A(n130), .B(n166), .Y(n168) );
  XOR2X1 U208 ( .A(B[16]), .B(A[16]), .Y(n114) );
  NOR2BX1 U209 ( .AN(n112), .B(n65), .Y(SUM[0]) );
  NOR2XL U210 ( .A(A[0]), .B(B[0]), .Y(n65) );
  OR2X2 U211 ( .A(n143), .B(n42), .Y(n67) );
  XOR2X2 U212 ( .A(n109), .B(n111), .Y(SUM[1]) );
  INVX1 U213 ( .A(n73), .Y(n211) );
  NOR2BX2 U214 ( .AN(n102), .B(n2), .Y(n101) );
  AND2X2 U215 ( .A(n73), .B(n184), .Y(n191) );
  INVXL U216 ( .A(n145), .Y(n143) );
  INVX1 U217 ( .A(n112), .Y(n109) );
  NOR2XL U218 ( .A(n168), .B(n134), .Y(n161) );
  NOR2X1 U219 ( .A(n124), .B(n125), .Y(n119) );
  NAND2XL U220 ( .A(B[15]), .B(A[15]), .Y(n121) );
  NAND2XL U221 ( .A(A[4]), .B(B[4]), .Y(n178) );
  NAND2XL U222 ( .A(n47), .B(n102), .Y(n140) );
  AOI21X4 U223 ( .A0(n94), .A1(n87), .B0(n17), .Y(n93) );
  NAND3BX4 U224 ( .AN(n161), .B(n162), .C(n163), .Y(n160) );
  OR2X4 U225 ( .A(A[13]), .B(B[13]), .Y(n166) );
  OAI211X2 U226 ( .A0(n41), .A1(n183), .B0(n184), .C0(n185), .Y(n182) );
  OR2X4 U227 ( .A(A[12]), .B(B[12]), .Y(n130) );
  OR2X4 U228 ( .A(A[1]), .B(B[1]), .Y(n108) );
  AND2X2 U229 ( .A(B[1]), .B(A[1]), .Y(n210) );
  OR2X4 U230 ( .A(A[7]), .B(B[7]), .Y(n145) );
  OR2X4 U231 ( .A(A[7]), .B(B[7]), .Y(n91) );
  OR2X4 U232 ( .A(A[8]), .B(B[8]), .Y(n80) );
  NAND2X4 U233 ( .A(B[7]), .B(A[7]), .Y(n92) );
  OR2X4 U234 ( .A(A[6]), .B(B[6]), .Y(n88) );
endmodule


module butterfly_DW01_sub_101 ( A, B, DIFF );
  input [16:0] A;
  input [16:0] B;
  output [16:0] DIFF;
  wire   n215, n216, n217, n218, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n37, n39, n40, n41,
         n42, n43, n44, n46, n47, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n60, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214;

  INVX4 U3 ( .A(n103), .Y(n100) );
  INVX2 U4 ( .A(A[8]), .Y(n25) );
  NOR2X4 U5 ( .A(n33), .B(n193), .Y(n197) );
  INVX2 U6 ( .A(n155), .Y(n186) );
  NAND3X4 U7 ( .A(n106), .B(n213), .C(n103), .Y(n4) );
  CLKINVX8 U8 ( .A(n86), .Y(n95) );
  BUFX12 U9 ( .A(n86), .Y(n10) );
  XOR2X4 U10 ( .A(n184), .B(n1), .Y(n216) );
  NOR2X1 U11 ( .A(n156), .B(n160), .Y(n1) );
  DLY1X1 U12 ( .A(n125), .Y(n2) );
  NAND2X1 U13 ( .A(n90), .B(n91), .Y(n28) );
  NAND2BX4 U14 ( .AN(n3), .B(n109), .Y(n18) );
  CLKINVX20 U15 ( .A(n111), .Y(n3) );
  INVX4 U16 ( .A(n106), .Y(n108) );
  NAND3X2 U17 ( .A(n106), .B(n213), .C(n103), .Y(n212) );
  INVX4 U18 ( .A(n109), .Y(n105) );
  XNOR2X4 U19 ( .A(n147), .B(n8), .Y(n57) );
  CLKINVX3 U20 ( .A(n126), .Y(n72) );
  INVX1 U21 ( .A(n136), .Y(n148) );
  NAND2BX2 U22 ( .AN(A[14]), .B(B[14]), .Y(n133) );
  NAND2BX4 U23 ( .AN(B[13]), .B(A[13]), .Y(n139) );
  INVX4 U24 ( .A(B[5]), .Y(n200) );
  INVX4 U25 ( .A(n123), .Y(n141) );
  NAND2X2 U26 ( .A(n114), .B(n115), .Y(n112) );
  INVXL U27 ( .A(n83), .Y(n82) );
  INVX4 U28 ( .A(n192), .Y(n191) );
  INVXL U29 ( .A(n74), .Y(n73) );
  CLKBUFX8 U30 ( .A(A[9]), .Y(n19) );
  CLKINVX3 U31 ( .A(n76), .Y(n174) );
  NAND2BX2 U32 ( .AN(B[11]), .B(A[11]), .Y(n163) );
  INVX1 U33 ( .A(n153), .Y(n160) );
  INVX3 U34 ( .A(n102), .Y(n32) );
  AOI2BB1X1 U35 ( .A0N(n127), .A1N(n128), .B0(n129), .Y(n114) );
  DLY1X1 U36 ( .A(n64), .Y(n5) );
  NAND2X2 U37 ( .A(n7), .B(n81), .Y(n78) );
  NAND2X4 U38 ( .A(n209), .B(n98), .Y(n7) );
  INVX1 U39 ( .A(n52), .Y(n22) );
  NAND2X4 U40 ( .A(n111), .B(n210), .Y(n179) );
  BUFX4 U41 ( .A(A[1]), .Y(n44) );
  NOR3BX4 U42 ( .AN(n125), .B(n198), .C(n172), .Y(n194) );
  AND2X1 U43 ( .A(n88), .B(n89), .Y(n6) );
  NAND2BX2 U44 ( .AN(B[9]), .B(n19), .Y(n69) );
  NAND2X1 U45 ( .A(n139), .B(n136), .Y(n8) );
  INVX8 U46 ( .A(n187), .Y(n166) );
  DLY1X1 U47 ( .A(n124), .Y(n9) );
  NAND2X4 U48 ( .A(n182), .B(n210), .Y(n213) );
  NOR2BX4 U49 ( .AN(A[9]), .B(B[9]), .Y(n167) );
  INVX4 U50 ( .A(B[4]), .Y(n17) );
  CLKBUFX2 U51 ( .A(n81), .Y(n43) );
  AND2X1 U52 ( .A(n83), .B(n76), .Y(n46) );
  NOR2BX4 U53 ( .AN(B[9]), .B(n19), .Y(n164) );
  NAND2BX4 U54 ( .AN(n211), .B(n4), .Y(n34) );
  NOR2X4 U55 ( .A(n11), .B(n205), .Y(n29) );
  NAND2BX4 U56 ( .AN(n206), .B(n203), .Y(n11) );
  INVX8 U57 ( .A(n12), .Y(n178) );
  NAND2X4 U58 ( .A(n42), .B(B[3]), .Y(n12) );
  OAI2BB1X4 U59 ( .A0N(A[5]), .A1N(n200), .B0(n201), .Y(n173) );
  NAND2X4 U60 ( .A(n17), .B(A[4]), .Y(n90) );
  OR2X2 U61 ( .A(n200), .B(A[5]), .Y(n13) );
  INVX4 U62 ( .A(n13), .Y(n205) );
  OR2X4 U63 ( .A(B[3]), .B(n42), .Y(n86) );
  INVX4 U64 ( .A(A[3]), .Y(n42) );
  OAI2BB1X4 U65 ( .A0N(n89), .A1N(n90), .B0(n88), .Y(n81) );
  NOR2X4 U66 ( .A(A[4]), .B(n17), .Y(n14) );
  INVX4 U67 ( .A(n14), .Y(n91) );
  NAND2BX4 U68 ( .AN(A[3]), .B(B[3]), .Y(n16) );
  AND3X4 U69 ( .A(n7), .B(n85), .C(n10), .Y(n15) );
  NOR2X4 U70 ( .A(n15), .B(n190), .Y(n189) );
  NAND2X2 U71 ( .A(n29), .B(n191), .Y(n190) );
  CLKINVX2 U72 ( .A(n80), .Y(n40) );
  INVX4 U73 ( .A(n181), .Y(n47) );
  OAI21X2 U74 ( .A0(n35), .A1(n148), .B0(n139), .Y(n145) );
  DLY1X1 U75 ( .A(n85), .Y(n20) );
  NAND2XL U76 ( .A(n68), .B(n69), .Y(n62) );
  XOR2X4 U77 ( .A(n22), .B(n70), .Y(n21) );
  XOR2X4 U78 ( .A(n104), .B(n60), .Y(n23) );
  NOR2X4 U79 ( .A(n178), .B(n179), .Y(n24) );
  CLKINVX4 U80 ( .A(n25), .Y(n26) );
  NOR3BX4 U81 ( .AN(n177), .B(n18), .C(n178), .Y(n176) );
  NAND2BX4 U82 ( .AN(A[2]), .B(n47), .Y(n177) );
  NAND2BX4 U83 ( .AN(A[9]), .B(B[9]), .Y(n37) );
  NOR3BX4 U84 ( .AN(n125), .B(n198), .C(n172), .Y(n33) );
  OAI2BB1X4 U85 ( .A0N(n31), .A1N(n85), .B0(n202), .Y(n196) );
  AND2X2 U86 ( .A(n84), .B(n10), .Y(n31) );
  NAND2BX2 U87 ( .AN(n178), .B(n86), .Y(n96) );
  NAND2BX4 U88 ( .AN(n95), .B(n85), .Y(n77) );
  OR2X2 U89 ( .A(n166), .B(n186), .Y(n50) );
  NOR2BX2 U90 ( .AN(B[4]), .B(A[4]), .Y(n207) );
  AOI21X4 U91 ( .A0(n173), .A1(n88), .B0(n174), .Y(n171) );
  NOR2BX2 U92 ( .AN(B[6]), .B(A[6]), .Y(n206) );
  NAND2BX4 U93 ( .AN(B[4]), .B(A[4]), .Y(n201) );
  AOI21X4 U94 ( .A0(n80), .A1(n81), .B0(n82), .Y(n79) );
  XOR2X4 U95 ( .A(n27), .B(n28), .Y(DIFF[4]) );
  AND3X2 U96 ( .A(n34), .B(n10), .C(n84), .Y(n27) );
  NOR2BX2 U97 ( .AN(B[7]), .B(A[7]), .Y(n208) );
  NAND2BXL U98 ( .AN(n123), .B(n74), .Y(n122) );
  NOR2X4 U99 ( .A(n205), .B(n206), .Y(n204) );
  BUFX20 U100 ( .A(n215), .Y(DIFF[15]) );
  OAI21X4 U101 ( .A0(n35), .A1(n148), .B0(n139), .Y(n30) );
  INVX8 U102 ( .A(n98), .Y(n102) );
  AOI2BB1X4 U103 ( .A0N(n70), .A1N(n149), .B0(n150), .Y(n35) );
  OAI21X4 U104 ( .A0(n151), .A1(n152), .B0(n140), .Y(n150) );
  NAND2X4 U105 ( .A(n83), .B(n74), .Y(n172) );
  NOR3X4 U106 ( .A(n175), .B(n176), .C(n95), .Y(n168) );
  NOR2BX2 U107 ( .AN(A[1]), .B(B[1]), .Y(n183) );
  BUFX20 U108 ( .A(n21), .Y(DIFF[8]) );
  NAND2X4 U109 ( .A(n181), .B(A[2]), .Y(n103) );
  INVX8 U110 ( .A(B[2]), .Y(n181) );
  NOR3X4 U111 ( .A(n39), .B(n189), .C(n188), .Y(n185) );
  OR2X4 U112 ( .A(n194), .B(n193), .Y(n39) );
  INVX2 U113 ( .A(n69), .Y(n193) );
  NAND2X2 U114 ( .A(n88), .B(n91), .Y(n80) );
  AOI21X2 U115 ( .A0(n180), .A1(n103), .B0(n211), .Y(n175) );
  OAI2BB1X4 U116 ( .A0N(n40), .A1N(n92), .B0(n43), .Y(n87) );
  NAND2X4 U117 ( .A(n154), .B(n155), .Y(n162) );
  NOR2X2 U118 ( .A(n124), .B(n192), .Y(n202) );
  NAND2BX2 U119 ( .AN(B[5]), .B(A[5]), .Y(n89) );
  INVX4 U120 ( .A(n46), .Y(n41) );
  OAI21X4 U121 ( .A0(n164), .A1(n67), .B0(n165), .Y(n154) );
  NAND2BX4 U122 ( .AN(A[1]), .B(B[1]), .Y(n210) );
  NAND2X4 U123 ( .A(n68), .B(n64), .Y(n198) );
  OR2X4 U124 ( .A(n105), .B(n108), .Y(n60) );
  AOI21X2 U125 ( .A0(n133), .A1(n145), .B0(n146), .Y(n144) );
  XOR2X4 U126 ( .A(n87), .B(n41), .Y(n51) );
  NAND2BX4 U127 ( .AN(n160), .B(n161), .Y(n119) );
  NAND2X4 U128 ( .A(n162), .B(n163), .Y(n161) );
  NAND2X4 U129 ( .A(n173), .B(n88), .Y(n199) );
  XOR2X4 U130 ( .A(n99), .B(n101), .Y(n218) );
  BUFX20 U131 ( .A(n218), .Y(DIFF[2]) );
  NOR2X4 U132 ( .A(n171), .B(n172), .Y(n170) );
  BUFX20 U133 ( .A(n23), .Y(DIFF[1]) );
  AOI21X2 U134 ( .A0(n155), .A1(n154), .B0(n156), .Y(n151) );
  AOI21X2 U135 ( .A0(n182), .A1(n109), .B0(n183), .Y(n180) );
  BUFX20 U136 ( .A(n216), .Y(DIFF[11]) );
  INVX8 U137 ( .A(n65), .Y(n70) );
  BUFX20 U138 ( .A(n217), .Y(DIFF[9]) );
  NAND4X2 U139 ( .A(n64), .B(n68), .C(n153), .D(n155), .Y(n123) );
  NAND2X2 U140 ( .A(n64), .B(n37), .Y(n214) );
  INVX8 U141 ( .A(n53), .Y(DIFF[3]) );
  AOI21X2 U142 ( .A0(n141), .A1(n65), .B0(n159), .Y(n158) );
  AOI21X4 U143 ( .A0(n65), .A1(n5), .B0(n66), .Y(n63) );
  NAND2X2 U144 ( .A(n92), .B(n91), .Y(n94) );
  NAND2BX4 U145 ( .AN(B[1]), .B(n44), .Y(n106) );
  OAI21X4 U146 ( .A0(A[2]), .A1(n181), .B0(n16), .Y(n211) );
  NAND2BX2 U147 ( .AN(A[15]), .B(B[15]), .Y(n134) );
  INVXL U148 ( .A(n138), .Y(n146) );
  XNOR2X4 U149 ( .A(n97), .B(n96), .Y(n53) );
  AND2X1 U150 ( .A(n64), .B(n67), .Y(n52) );
  INVX8 U151 ( .A(n55), .Y(DIFF[7]) );
  OR2X2 U152 ( .A(n72), .B(n73), .Y(n56) );
  INVX8 U153 ( .A(n57), .Y(DIFF[13]) );
  INVX8 U154 ( .A(n51), .Y(DIFF[6]) );
  NAND2BX2 U155 ( .AN(B[12]), .B(A[12]), .Y(n140) );
  INVX8 U156 ( .A(n49), .Y(DIFF[10]) );
  INVX4 U157 ( .A(n119), .Y(n159) );
  NAND2XL U158 ( .A(n142), .B(n153), .Y(n152) );
  INVXL U159 ( .A(n118), .Y(n117) );
  NAND2BX4 U160 ( .AN(B[8]), .B(n26), .Y(n67) );
  NAND2X2 U161 ( .A(n132), .B(n134), .Y(n143) );
  NAND2XL U162 ( .A(n138), .B(n139), .Y(n137) );
  NAND2XL U163 ( .A(n133), .B(n134), .Y(n131) );
  OAI21XL U164 ( .A0(n130), .A1(n131), .B0(n132), .Y(n129) );
  XOR2X4 U165 ( .A(n195), .B(n50), .Y(n49) );
  NAND2XL U166 ( .A(n142), .B(n140), .Y(n157) );
  INVX1 U167 ( .A(n163), .Y(n156) );
  INVX1 U168 ( .A(n67), .Y(n66) );
  OAI21X1 U169 ( .A0(n116), .A1(n159), .B0(n117), .Y(n115) );
  AOI21X1 U170 ( .A0(n120), .A1(n121), .B0(n122), .Y(n116) );
  OR2XL U171 ( .A(n54), .B(n9), .Y(n121) );
  AND2X1 U172 ( .A(n20), .B(n10), .Y(n54) );
  XOR2X4 U173 ( .A(n71), .B(n56), .Y(n55) );
  XOR2X4 U174 ( .A(n30), .B(n58), .Y(DIFF[14]) );
  AND2X2 U175 ( .A(n133), .B(n138), .Y(n58) );
  INVX1 U176 ( .A(n107), .Y(n104) );
  NAND4XL U177 ( .A(n134), .B(n133), .C(n142), .D(n136), .Y(n118) );
  AOI21XL U178 ( .A0(n135), .A1(n136), .B0(n137), .Y(n130) );
  INVXL U179 ( .A(n140), .Y(n135) );
  AOI21XL U180 ( .A0(n2), .A1(n83), .B0(n72), .Y(n120) );
  NAND2BXL U181 ( .AN(n118), .B(n141), .Y(n127) );
  XNOR2X1 U182 ( .A(B[16]), .B(A[16]), .Y(n113) );
  NAND2BX1 U183 ( .AN(B[14]), .B(A[14]), .Y(n138) );
  NAND2BX1 U184 ( .AN(B[15]), .B(A[15]), .Y(n132) );
  NAND2X1 U185 ( .A(n110), .B(n111), .Y(DIFF[0]) );
  INVX1 U186 ( .A(n110), .Y(n182) );
  NAND2BX1 U187 ( .AN(n111), .B(n110), .Y(n107) );
  NAND2BX1 U188 ( .AN(A[0]), .B(B[0]), .Y(n111) );
  NAND2BX1 U189 ( .AN(B[0]), .B(A[0]), .Y(n110) );
  NAND2BXL U190 ( .AN(n7), .B(n29), .Y(n128) );
  NAND2BX4 U191 ( .AN(A[1]), .B(B[1]), .Y(n109) );
  NAND2BX4 U192 ( .AN(A[2]), .B(n47), .Y(n98) );
  XOR2X4 U193 ( .A(n63), .B(n62), .Y(n217) );
  NAND2X4 U194 ( .A(n75), .B(n76), .Y(n71) );
  OAI21X4 U195 ( .A0(n77), .A1(n78), .B0(n79), .Y(n75) );
  XOR2X4 U196 ( .A(n93), .B(n6), .Y(DIFF[5]) );
  NAND2X4 U197 ( .A(n94), .B(n90), .Y(n93) );
  NAND3BX4 U198 ( .AN(n95), .B(n34), .C(n84), .Y(n92) );
  AOI21X4 U199 ( .A0(n99), .A1(n32), .B0(n100), .Y(n97) );
  NOR2X4 U200 ( .A(n102), .B(n100), .Y(n101) );
  OAI21X4 U201 ( .A0(n105), .A1(n104), .B0(n106), .Y(n99) );
  XOR2X4 U202 ( .A(n112), .B(n113), .Y(DIFF[16]) );
  XOR2X4 U203 ( .A(n144), .B(n143), .Y(n215) );
  AOI2BB1X4 U204 ( .A0N(n70), .A1N(n149), .B0(n150), .Y(n147) );
  NAND2X4 U205 ( .A(n142), .B(n141), .Y(n149) );
  NAND2BX4 U206 ( .AN(A[13]), .B(B[13]), .Y(n136) );
  XOR2X4 U207 ( .A(n158), .B(n157), .Y(DIFF[12]) );
  NOR2X4 U208 ( .A(n166), .B(n167), .Y(n165) );
  OAI21X4 U209 ( .A0(n168), .A1(n124), .B0(n169), .Y(n65) );
  NOR2X4 U210 ( .A(n72), .B(n170), .Y(n169) );
  NAND2BX4 U211 ( .AN(A[12]), .B(B[12]), .Y(n142) );
  NAND2BX4 U212 ( .AN(A[11]), .B(B[11]), .Y(n153) );
  OAI21X4 U213 ( .A0(n185), .A1(n186), .B0(n187), .Y(n184) );
  NAND2BX4 U214 ( .AN(A[10]), .B(B[10]), .Y(n155) );
  NAND2BX4 U215 ( .AN(B[10]), .B(A[10]), .Y(n187) );
  NAND3BX4 U216 ( .AN(n188), .B(n197), .C(n196), .Y(n195) );
  NAND2BX4 U217 ( .AN(A[7]), .B(B[7]), .Y(n74) );
  NAND2BX4 U218 ( .AN(A[6]), .B(B[6]), .Y(n83) );
  NAND2X4 U219 ( .A(n199), .B(n76), .Y(n125) );
  NAND2BX4 U220 ( .AN(B[6]), .B(A[6]), .Y(n76) );
  NAND2BX4 U221 ( .AN(A[5]), .B(B[5]), .Y(n88) );
  NAND2X4 U222 ( .A(n204), .B(n203), .Y(n124) );
  NOR2X4 U223 ( .A(n207), .B(n208), .Y(n203) );
  NAND2X4 U224 ( .A(n37), .B(n64), .Y(n192) );
  NAND2X4 U225 ( .A(n24), .B(n177), .Y(n84) );
  NOR2X4 U226 ( .A(n178), .B(n18), .Y(n209) );
  NAND2BX4 U227 ( .AN(n211), .B(n212), .Y(n85) );
  AOI21X4 U228 ( .A0(n67), .A1(n126), .B0(n214), .Y(n188) );
  NAND2BX4 U229 ( .AN(A[9]), .B(B[9]), .Y(n68) );
  NAND2BX4 U230 ( .AN(A[8]), .B(B[8]), .Y(n64) );
  NAND2BX4 U231 ( .AN(B[7]), .B(A[7]), .Y(n126) );
endmodule


module butterfly_DW01_sub_96 ( A, B, DIFF );
  input [16:0] A;
  input [16:0] B;
  output [16:0] DIFF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181;

  DLY1X1 U3 ( .A(n29), .Y(n1) );
  INVXL U4 ( .A(B[6]), .Y(n26) );
  CLKINVX4 U5 ( .A(n51), .Y(n4) );
  OAI21X1 U6 ( .A0(n98), .A1(n99), .B0(n100), .Y(n97) );
  AOI21X1 U7 ( .A0(n103), .A1(n33), .B0(n105), .Y(n98) );
  INVX4 U8 ( .A(n118), .Y(n2) );
  INVX8 U9 ( .A(n119), .Y(n118) );
  NAND2BX4 U10 ( .AN(A[4]), .B(B[4]), .Y(n68) );
  INVX8 U11 ( .A(n180), .Y(n8) );
  NAND2BX2 U12 ( .AN(B[14]), .B(A[14]), .Y(n106) );
  NAND2BX2 U13 ( .AN(A[5]), .B(B[5]), .Y(n122) );
  NAND2BX4 U14 ( .AN(B[2]), .B(A[2]), .Y(n80) );
  INVX1 U15 ( .A(n80), .Y(n76) );
  NAND2X4 U16 ( .A(n4), .B(n50), .Y(n5) );
  NAND2X2 U17 ( .A(n3), .B(n51), .Y(n6) );
  NAND2X4 U18 ( .A(n5), .B(n6), .Y(DIFF[7]) );
  CLKINVX2 U19 ( .A(n50), .Y(n3) );
  NAND2X4 U20 ( .A(n15), .B(n34), .Y(n50) );
  NAND4BX4 U21 ( .AN(n18), .B(n8), .C(n31), .D(n35), .Y(n7) );
  NAND4BX2 U22 ( .AN(n18), .B(n8), .C(n31), .D(n35), .Y(n133) );
  NAND3BX4 U23 ( .AN(n29), .B(n78), .C(n28), .Y(n31) );
  NAND2BX1 U24 ( .AN(n180), .B(n60), .Y(n63) );
  CLKBUFX4 U25 ( .A(n31), .Y(n9) );
  NAND3X4 U26 ( .A(n156), .B(A[8]), .C(n45), .Y(n152) );
  NAND2BX2 U27 ( .AN(A[1]), .B(B[1]), .Y(n86) );
  INVX8 U28 ( .A(n57), .Y(n180) );
  NAND4X2 U29 ( .A(n102), .B(n13), .C(n111), .D(n33), .Y(n92) );
  INVX3 U30 ( .A(n61), .Y(n179) );
  AOI21X2 U31 ( .A0(n74), .A1(n75), .B0(n76), .Y(n73) );
  NAND2X2 U32 ( .A(n100), .B(n102), .Y(n123) );
  CLKINVX4 U33 ( .A(n92), .Y(n96) );
  AOI21X2 U34 ( .A0(n127), .A1(n13), .B0(n128), .Y(n126) );
  INVX8 U35 ( .A(n132), .Y(n13) );
  BUFX16 U36 ( .A(n104), .Y(n33) );
  INVX2 U37 ( .A(n74), .Y(n79) );
  AOI21X2 U38 ( .A0(n66), .A1(n67), .B0(n181), .Y(n177) );
  INVX1 U39 ( .A(A[1]), .Y(n176) );
  NOR2X2 U40 ( .A(n135), .B(n134), .Y(n124) );
  NAND2X1 U41 ( .A(n137), .B(n101), .Y(n136) );
  NAND2BX2 U42 ( .AN(A[15]), .B(B[15]), .Y(n102) );
  INVX4 U43 ( .A(n101), .Y(n132) );
  INVX1 U44 ( .A(n106), .Y(n128) );
  INVX1 U45 ( .A(n142), .Y(n103) );
  INVX1 U46 ( .A(n21), .Y(n22) );
  NAND2X1 U47 ( .A(n56), .B(n66), .Y(n69) );
  NOR2X2 U48 ( .A(n44), .B(n48), .Y(n47) );
  NAND2BX1 U49 ( .AN(B[6]), .B(A[6]), .Y(n60) );
  INVX1 U50 ( .A(n111), .Y(n147) );
  NAND3BX4 U51 ( .AN(n29), .B(n78), .C(n120), .Y(n10) );
  NAND2BX1 U52 ( .AN(B[15]), .B(A[15]), .Y(n100) );
  INVXL U53 ( .A(n1), .Y(n109) );
  NOR3X4 U54 ( .A(n48), .B(n154), .C(n168), .Y(n164) );
  BUFX8 U55 ( .A(n7), .Y(n11) );
  XOR2X4 U56 ( .A(n149), .B(n12), .Y(DIFF[12]) );
  AND2X4 U57 ( .A(n111), .B(n142), .Y(n12) );
  NAND2X1 U58 ( .A(n45), .B(n46), .Y(n40) );
  NAND2BX4 U59 ( .AN(B[12]), .B(A[12]), .Y(n142) );
  BUFX4 U60 ( .A(n61), .Y(n15) );
  NOR2X2 U61 ( .A(n48), .B(n168), .Y(n172) );
  INVX8 U62 ( .A(n43), .Y(n48) );
  NAND2X4 U63 ( .A(n111), .B(n33), .Y(n14) );
  NAND2BX4 U64 ( .AN(B[3]), .B(A[3]), .Y(n78) );
  INVX4 U65 ( .A(n45), .Y(n168) );
  AND2X4 U66 ( .A(n178), .B(n177), .Y(n16) );
  BUFX1 U67 ( .A(A[6]), .Y(n17) );
  NAND2BX2 U68 ( .AN(B[13]), .B(A[13]), .Y(n107) );
  NOR2BX2 U69 ( .AN(B[11]), .B(A[11]), .Y(n159) );
  NAND2XL U70 ( .A(n77), .B(n78), .Y(n72) );
  INVX2 U71 ( .A(n46), .Y(n167) );
  NAND2BX2 U72 ( .AN(B[8]), .B(A[8]), .Y(n49) );
  NAND2X4 U73 ( .A(n121), .B(n122), .Y(n18) );
  NAND2BX4 U74 ( .AN(A[10]), .B(B[10]), .Y(n160) );
  NOR2X2 U75 ( .A(n76), .B(n79), .Y(n37) );
  AND2X2 U76 ( .A(n34), .B(n49), .Y(n39) );
  AND2X2 U77 ( .A(n10), .B(n68), .Y(n32) );
  AOI21X4 U78 ( .A0(A[9]), .A1(n157), .B0(n158), .Y(n151) );
  NOR3X4 U79 ( .A(n131), .B(n108), .C(n132), .Y(n130) );
  AND2X4 U80 ( .A(n77), .B(n74), .Y(n175) );
  CLKINVX2 U81 ( .A(n58), .Y(n19) );
  INVX8 U82 ( .A(n67), .Y(n58) );
  BUFX8 U83 ( .A(n114), .Y(n20) );
  AND2X4 U84 ( .A(n27), .B(n20), .Y(n150) );
  NAND2BX2 U85 ( .AN(B[11]), .B(A[11]), .Y(n114) );
  INVXL U86 ( .A(n113), .Y(n21) );
  NAND4X1 U87 ( .A(n56), .B(n15), .C(n68), .D(n8), .Y(n110) );
  XOR2X4 U88 ( .A(n9), .B(n38), .Y(DIFF[4]) );
  INVX8 U89 ( .A(n23), .Y(n119) );
  NAND2XL U90 ( .A(n20), .B(n22), .Y(n144) );
  NAND4BX4 U91 ( .AN(n16), .B(n34), .C(n11), .D(n2), .Y(n129) );
  AND3X4 U92 ( .A(n61), .B(n17), .C(n26), .Y(n23) );
  CLKINVX8 U93 ( .A(n108), .Y(n95) );
  NAND2X1 U94 ( .A(n13), .B(n102), .Y(n99) );
  AOI21X4 U95 ( .A0(n115), .A1(n116), .B0(n108), .Y(n112) );
  XNOR2X4 U96 ( .A(n138), .B(n24), .Y(DIFF[14]) );
  OR2X2 U97 ( .A(n128), .B(n132), .Y(n24) );
  NOR2X2 U98 ( .A(n14), .B(n136), .Y(n134) );
  NOR3X4 U99 ( .A(n27), .B(n132), .C(n131), .Y(n135) );
  NOR2BX4 U100 ( .AN(n60), .B(n52), .Y(n51) );
  XOR2X4 U101 ( .A(n145), .B(n25), .Y(DIFF[13]) );
  AND2X1 U102 ( .A(n107), .B(n33), .Y(n25) );
  OAI2BB1X4 U103 ( .A0N(n151), .A1N(n152), .B0(n153), .Y(n27) );
  OAI21X4 U104 ( .A0(n173), .A1(n174), .B0(n175), .Y(n28) );
  NAND2X4 U105 ( .A(n113), .B(n20), .Y(n148) );
  INVX2 U106 ( .A(n49), .Y(n44) );
  BUFX12 U107 ( .A(n62), .Y(n34) );
  NAND2BX2 U108 ( .AN(B[7]), .B(A[7]), .Y(n62) );
  NAND4BX4 U109 ( .AN(n16), .B(n34), .C(n11), .D(n2), .Y(n143) );
  NAND2X4 U110 ( .A(n80), .B(n83), .Y(n174) );
  INVX2 U111 ( .A(n68), .Y(n71) );
  AND4X4 U112 ( .A(n77), .B(n86), .C(n74), .D(n88), .Y(n29) );
  NAND2BX4 U113 ( .AN(A[2]), .B(B[2]), .Y(n74) );
  NAND2BX4 U114 ( .AN(B[4]), .B(A[4]), .Y(n67) );
  NAND2BX2 U115 ( .AN(B[9]), .B(A[9]), .Y(n46) );
  OAI2BB1X4 U116 ( .A0N(n129), .A1N(n95), .B0(n150), .Y(n149) );
  XNOR2X4 U117 ( .A(n162), .B(n30), .Y(DIFF[11]) );
  OR2X2 U118 ( .A(n137), .B(n155), .Y(n30) );
  OAI21X4 U119 ( .A0(n91), .A1(n92), .B0(n93), .Y(n89) );
  NOR2X2 U120 ( .A(n112), .B(n144), .Y(n91) );
  NOR2XL U121 ( .A(n109), .B(n110), .Y(n94) );
  NOR2X2 U122 ( .A(n117), .B(n118), .Y(n115) );
  NAND2BX2 U123 ( .AN(A[11]), .B(B[11]), .Y(n163) );
  NAND4X4 U124 ( .A(n161), .B(n34), .C(n133), .D(n119), .Y(n42) );
  NAND3X4 U125 ( .A(n124), .B(n125), .C(n126), .Y(n36) );
  OAI21X4 U126 ( .A0(n81), .A1(n82), .B0(n83), .Y(n75) );
  INVX4 U127 ( .A(n86), .Y(n82) );
  NAND2X2 U128 ( .A(n143), .B(n130), .Y(n125) );
  AOI21X1 U129 ( .A0(n28), .A1(n78), .B0(n110), .Y(n117) );
  NAND2BX1 U130 ( .AN(A[4]), .B(B[4]), .Y(n35) );
  INVX4 U131 ( .A(n163), .Y(n155) );
  NAND2BX4 U132 ( .AN(A[13]), .B(B[13]), .Y(n104) );
  INVX4 U133 ( .A(n33), .Y(n141) );
  OAI2BB1X4 U134 ( .A0N(n172), .A1N(n165), .B0(n46), .Y(n169) );
  NAND2BX4 U135 ( .AN(A[5]), .B(B[5]), .Y(n56) );
  NAND2BX2 U136 ( .AN(B[10]), .B(A[10]), .Y(n171) );
  NOR2X2 U137 ( .A(n158), .B(n154), .Y(n170) );
  AOI21X1 U138 ( .A0(n167), .A1(n160), .B0(n158), .Y(n166) );
  XOR2X4 U139 ( .A(n89), .B(n90), .Y(DIFF[16]) );
  NAND4X4 U140 ( .A(n161), .B(n7), .C(n39), .D(n119), .Y(n165) );
  NAND2BX4 U141 ( .AN(A[9]), .B(B[9]), .Y(n45) );
  NAND2X4 U142 ( .A(n10), .B(n68), .Y(n54) );
  AOI31X2 U143 ( .A0(n94), .A1(n95), .A2(n96), .B0(n97), .Y(n93) );
  AOI21X2 U144 ( .A0(n176), .A1(B[1]), .B0(n87), .Y(n173) );
  NAND2BX4 U145 ( .AN(A[7]), .B(B[7]), .Y(n61) );
  NAND2BX4 U146 ( .AN(A[7]), .B(B[7]), .Y(n121) );
  NOR2BX4 U147 ( .AN(n83), .B(n82), .Y(n85) );
  NAND2BX4 U148 ( .AN(B[1]), .B(A[1]), .Y(n83) );
  INVX8 U149 ( .A(n66), .Y(n59) );
  NAND2BX4 U150 ( .AN(B[5]), .B(A[5]), .Y(n66) );
  NAND2BX4 U151 ( .AN(A[8]), .B(B[8]), .Y(n43) );
  INVX8 U152 ( .A(n160), .Y(n154) );
  NOR2X4 U153 ( .A(n32), .B(n58), .Y(n70) );
  AOI21X4 U154 ( .A0(n42), .A1(n43), .B0(n44), .Y(n41) );
  NAND4BX4 U155 ( .AN(n159), .B(n160), .C(n45), .D(n43), .Y(n108) );
  XOR2X2 U156 ( .A(n75), .B(n37), .Y(DIFF[2]) );
  XOR2X4 U157 ( .A(n42), .B(n47), .Y(DIFF[8]) );
  INVX4 U158 ( .A(n114), .Y(n137) );
  XNOR2X4 U159 ( .A(n36), .B(n123), .Y(DIFF[15]) );
  INVX4 U160 ( .A(n171), .Y(n158) );
  AOI21X4 U161 ( .A0(n65), .A1(n56), .B0(n59), .Y(n64) );
  NOR2X4 U162 ( .A(n71), .B(n58), .Y(n38) );
  INVXL U163 ( .A(B[9]), .Y(n157) );
  INVX2 U164 ( .A(n127), .Y(n140) );
  NOR2BXL U165 ( .AN(n34), .B(n16), .Y(n116) );
  NAND2XL U166 ( .A(n106), .B(n107), .Y(n105) );
  INVX1 U167 ( .A(n84), .Y(n81) );
  XNOR2X1 U168 ( .A(B[16]), .B(A[16]), .Y(n90) );
  NAND2X1 U169 ( .A(n87), .B(n88), .Y(DIFF[0]) );
  NAND2BX1 U170 ( .AN(n88), .B(n87), .Y(n84) );
  NAND2BX1 U171 ( .AN(A[0]), .B(B[0]), .Y(n88) );
  NAND2BX1 U172 ( .AN(B[0]), .B(A[0]), .Y(n87) );
  INVXL U173 ( .A(B[8]), .Y(n156) );
  NOR2BX1 U174 ( .AN(B[5]), .B(A[5]), .Y(n181) );
  AOI21X4 U175 ( .A0(n53), .A1(n54), .B0(n55), .Y(n52) );
  NAND2X2 U176 ( .A(n57), .B(n56), .Y(n55) );
  XOR2X4 U177 ( .A(n41), .B(n40), .Y(DIFF[9]) );
  NOR2X4 U178 ( .A(n58), .B(n59), .Y(n53) );
  XOR2X4 U179 ( .A(n63), .B(n64), .Y(DIFF[6]) );
  NAND2X4 U180 ( .A(n19), .B(n54), .Y(n65) );
  XOR2X4 U181 ( .A(n70), .B(n69), .Y(DIFF[5]) );
  XOR2X4 U182 ( .A(n72), .B(n73), .Y(DIFF[3]) );
  XOR2X4 U183 ( .A(n84), .B(n85), .Y(DIFF[1]) );
  NAND2BX4 U184 ( .AN(A[14]), .B(B[14]), .Y(n101) );
  OAI21X4 U185 ( .A0(n139), .A1(n14), .B0(n140), .Y(n138) );
  OAI21X4 U186 ( .A0(n141), .A1(n142), .B0(n107), .Y(n127) );
  NAND2X4 U187 ( .A(n111), .B(n33), .Y(n131) );
  AOI21X4 U188 ( .A0(n129), .A1(n95), .B0(n148), .Y(n139) );
  OAI21X4 U189 ( .A0(n146), .A1(n147), .B0(n142), .Y(n145) );
  AOI21X4 U190 ( .A0(n95), .A1(n143), .B0(n148), .Y(n146) );
  NAND2BX4 U191 ( .AN(A[12]), .B(B[12]), .Y(n111) );
  OAI2BB1X4 U192 ( .A0N(n151), .A1N(n152), .B0(n153), .Y(n113) );
  NOR2X4 U193 ( .A(n154), .B(n155), .Y(n153) );
  OAI2BB1X4 U194 ( .A0N(n164), .A1N(n165), .B0(n166), .Y(n162) );
  XOR2X4 U195 ( .A(n169), .B(n170), .Y(DIFF[10]) );
  OAI21X4 U196 ( .A0(n173), .A1(n174), .B0(n175), .Y(n120) );
  NAND2BX4 U197 ( .AN(A[3]), .B(B[3]), .Y(n77) );
  NAND2X4 U198 ( .A(n177), .B(n178), .Y(n161) );
  NOR2X4 U199 ( .A(n180), .B(n179), .Y(n178) );
  NAND2BX4 U200 ( .AN(A[6]), .B(B[6]), .Y(n57) );
endmodule


module butterfly_DW01_sub_104 ( A, B, DIFF );
  input [16:0] A;
  input [16:0] B;
  output [16:0] DIFF;
  wire   n198, n1, n2, n3, n5, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197;

  NAND2X4 U3 ( .A(n164), .B(n165), .Y(n160) );
  OR2X4 U4 ( .A(B[5]), .B(n1), .Y(n48) );
  CLKINVX20 U5 ( .A(A[5]), .Y(n1) );
  INVX4 U6 ( .A(n180), .Y(n2) );
  INVX4 U7 ( .A(n35), .Y(n180) );
  INVX8 U8 ( .A(n103), .Y(n146) );
  NAND2X4 U9 ( .A(n75), .B(n68), .Y(n193) );
  INVX2 U10 ( .A(n32), .Y(n29) );
  OR2X4 U11 ( .A(B[9]), .B(n19), .Y(n32) );
  NAND2X4 U12 ( .A(n125), .B(n145), .Y(n144) );
  NAND2BX4 U13 ( .AN(A[10]), .B(B[10]), .Y(n163) );
  CLKINVX3 U14 ( .A(n159), .Y(n139) );
  NAND3X4 U15 ( .A(n155), .B(n156), .C(n41), .Y(n159) );
  NAND2BX4 U16 ( .AN(A[6]), .B(B[6]), .Y(n51) );
  INVX8 U17 ( .A(n50), .Y(n58) );
  XOR2X4 U18 ( .A(n21), .B(n3), .Y(DIFF[10]) );
  AND2X1 U19 ( .A(n163), .B(n165), .Y(n3) );
  INVX2 U20 ( .A(n119), .Y(n187) );
  AOI21X2 U21 ( .A0(n184), .A1(n120), .B0(n177), .Y(n182) );
  CLKINVX4 U22 ( .A(n125), .Y(n148) );
  XOR2X4 U23 ( .A(n157), .B(n158), .Y(n198) );
  NOR2X2 U24 ( .A(n154), .B(n148), .Y(n158) );
  XNOR2X2 U25 ( .A(n77), .B(n76), .Y(DIFF[4]) );
  NOR2X2 U26 ( .A(n112), .B(n148), .Y(n147) );
  NAND2BX4 U27 ( .AN(n36), .B(n37), .Y(n34) );
  INVX4 U28 ( .A(n36), .Y(n176) );
  BUFX8 U29 ( .A(n198), .Y(DIFF[12]) );
  NAND2BX4 U30 ( .AN(A[1]), .B(B[1]), .Y(n196) );
  INVX4 U31 ( .A(A[4]), .Y(n18) );
  AOI2BB1X2 U32 ( .A0N(n29), .A1N(n33), .B0(n175), .Y(n172) );
  INVXL U33 ( .A(A[15]), .Y(n14) );
  OAI2BB1X2 U34 ( .A0N(n59), .A1N(n50), .B0(n48), .Y(n55) );
  BUFX3 U35 ( .A(n74), .Y(n17) );
  INVX2 U36 ( .A(n81), .Y(n70) );
  INVX1 U37 ( .A(A[9]), .Y(n19) );
  INVX1 U38 ( .A(n124), .Y(n109) );
  OAI21X1 U39 ( .A0(n112), .A1(n113), .B0(n111), .Y(n143) );
  CLKINVX3 U40 ( .A(n196), .Y(n86) );
  NAND2BX2 U41 ( .AN(B[1]), .B(A[1]), .Y(n87) );
  CLKINVX3 U42 ( .A(n84), .Y(n69) );
  INVX1 U43 ( .A(n33), .Y(n16) );
  INVXL U44 ( .A(n102), .Y(n93) );
  NAND2X2 U45 ( .A(n40), .B(n41), .Y(n39) );
  NAND2BX1 U46 ( .AN(B[0]), .B(A[0]), .Y(n90) );
  NAND2X1 U47 ( .A(n123), .B(n196), .Y(n195) );
  NAND3X1 U48 ( .A(n123), .B(n75), .C(n196), .Y(n65) );
  NAND2X2 U49 ( .A(n195), .B(n84), .Y(n194) );
  NAND2BX4 U50 ( .AN(B[8]), .B(A[8]), .Y(n38) );
  XNOR2X2 U51 ( .A(n85), .B(n89), .Y(DIFF[1]) );
  AND2X4 U52 ( .A(n146), .B(n10), .Y(n5) );
  NAND2X1 U53 ( .A(n50), .B(n51), .Y(n49) );
  NOR2X2 U54 ( .A(n138), .B(n109), .Y(n137) );
  INVX1 U55 ( .A(n110), .Y(n138) );
  NAND2BX2 U56 ( .AN(A[13]), .B(B[13]), .Y(n7) );
  INVX1 U57 ( .A(B[8]), .Y(n183) );
  NAND2XL U58 ( .A(n11), .B(n54), .Y(n43) );
  XOR2X4 U59 ( .A(n171), .B(n8), .Y(DIFF[11]) );
  AND2X2 U60 ( .A(n164), .B(n145), .Y(n8) );
  OAI21X4 U61 ( .A0(n182), .A1(n36), .B0(n16), .Y(n181) );
  AND2X2 U62 ( .A(B[4]), .B(n18), .Y(n67) );
  NAND2BX2 U63 ( .AN(B[3]), .B(A[3]), .Y(n81) );
  NAND2BX1 U64 ( .AN(B[3]), .B(A[3]), .Y(n122) );
  BUFX8 U65 ( .A(n101), .Y(n9) );
  INVX2 U66 ( .A(n51), .Y(n57) );
  NOR2BX4 U67 ( .AN(n51), .B(n190), .Y(n189) );
  NAND2BX4 U68 ( .AN(n177), .B(n25), .Y(n37) );
  INVX1 U69 ( .A(n40), .Y(n118) );
  OAI21X4 U70 ( .A0(n121), .A1(n26), .B0(n11), .Y(n40) );
  OAI21X4 U71 ( .A0(n180), .A1(n181), .B0(n31), .Y(n179) );
  INVX8 U72 ( .A(n126), .Y(n112) );
  INVX1 U73 ( .A(A[14]), .Y(n12) );
  INVX4 U74 ( .A(n148), .Y(n10) );
  NAND2BX4 U75 ( .AN(A[7]), .B(B[7]), .Y(n11) );
  NAND3X2 U76 ( .A(n128), .B(n129), .C(n130), .Y(n23) );
  INVX4 U77 ( .A(n38), .Y(n33) );
  OR2X2 U78 ( .A(B[14]), .B(n12), .Y(n110) );
  OAI21X2 U79 ( .A0(B[1]), .A1(n197), .B0(n90), .Y(n123) );
  BUFX8 U80 ( .A(n42), .Y(n13) );
  OR2X4 U81 ( .A(B[15]), .B(n14), .Y(n97) );
  AND3X4 U82 ( .A(n192), .B(n122), .C(n9), .Y(n15) );
  NAND2BX4 U83 ( .AN(n193), .B(n194), .Y(n192) );
  NAND2BX4 U84 ( .AN(B[7]), .B(A[7]), .Y(n54) );
  OAI21X4 U85 ( .A0(n139), .A1(n140), .B0(n141), .Y(n136) );
  CLKINVX3 U86 ( .A(n88), .Y(n85) );
  NAND3BX4 U87 ( .AN(n58), .B(n42), .C(n17), .Y(n191) );
  NOR2BX2 U88 ( .AN(n87), .B(n86), .Y(n89) );
  AOI21X2 U89 ( .A0(n93), .A1(n94), .B0(n95), .Y(n91) );
  OAI21X1 U90 ( .A0(n114), .A1(n103), .B0(n115), .Y(n94) );
  NAND2X4 U91 ( .A(n163), .B(n31), .Y(n175) );
  NAND3X4 U92 ( .A(n73), .B(n196), .C(n74), .Y(n71) );
  NOR2X1 U93 ( .A(n144), .B(n112), .Y(n142) );
  NAND2X1 U94 ( .A(n74), .B(n50), .Y(n167) );
  NAND2X1 U95 ( .A(n74), .B(n72), .Y(n76) );
  AOI21X2 U96 ( .A0(n133), .A1(n134), .B0(n135), .Y(n129) );
  NAND3BX4 U97 ( .AN(n190), .B(n120), .C(n169), .Y(n155) );
  NAND4BX4 U98 ( .AN(n172), .B(n173), .C(n165), .D(n174), .Y(n171) );
  NAND2BX2 U99 ( .AN(B[11]), .B(A[11]), .Y(n164) );
  NAND3X2 U100 ( .A(n178), .B(n119), .C(n51), .Y(n25) );
  NAND2BX4 U101 ( .AN(A[15]), .B(B[15]), .Y(n127) );
  NOR2X4 U102 ( .A(n151), .B(n112), .Y(n150) );
  NOR2X2 U103 ( .A(n112), .B(n113), .Y(n105) );
  NOR2X2 U104 ( .A(n9), .B(n102), .Y(n100) );
  CLKINVX4 U105 ( .A(n127), .Y(n108) );
  NOR2X4 U106 ( .A(n167), .B(n168), .Y(n166) );
  NAND2X2 U107 ( .A(n11), .B(n51), .Y(n168) );
  OAI21X4 U108 ( .A0(n193), .A1(n71), .B0(n72), .Y(n62) );
  AOI21X4 U109 ( .A0(n47), .A1(n48), .B0(n49), .Y(n46) );
  INVX4 U110 ( .A(n59), .Y(n47) );
  NAND4BX4 U111 ( .AN(n170), .B(n163), .C(n31), .D(n13), .Y(n103) );
  NAND2BX4 U112 ( .AN(B[2]), .B(A[2]), .Y(n84) );
  NAND2BX4 U113 ( .AN(A[2]), .B(B[2]), .Y(n75) );
  NOR2X2 U114 ( .A(n69), .B(n83), .Y(n82) );
  NAND2X4 U115 ( .A(n179), .B(n32), .Y(n21) );
  NAND3X2 U116 ( .A(n96), .B(n97), .C(n98), .Y(n95) );
  NAND2BX4 U117 ( .AN(B[10]), .B(A[10]), .Y(n165) );
  XOR2X4 U118 ( .A(n23), .B(n24), .Y(DIFF[15]) );
  NAND2BX4 U119 ( .AN(A[8]), .B(B[8]), .Y(n42) );
  INVX2 U120 ( .A(n111), .Y(n151) );
  NAND2BX2 U121 ( .AN(A[11]), .B(B[11]), .Y(n145) );
  NAND3BX2 U122 ( .AN(n175), .B(n176), .C(n37), .Y(n173) );
  INVX2 U123 ( .A(n48), .Y(n61) );
  NAND2X4 U124 ( .A(n48), .B(n72), .Y(n120) );
  NOR2X1 U125 ( .A(n144), .B(n132), .Y(n134) );
  NAND2X4 U126 ( .A(n7), .B(n124), .Y(n132) );
  INVX1 U127 ( .A(n132), .Y(n131) );
  NOR2BX2 U128 ( .AN(B[11]), .B(A[11]), .Y(n170) );
  NAND2BX4 U129 ( .AN(A[13]), .B(B[13]), .Y(n126) );
  NOR2X4 U130 ( .A(n29), .B(n30), .Y(n28) );
  NAND2X2 U131 ( .A(n32), .B(n38), .Y(n162) );
  NOR2X4 U132 ( .A(n191), .B(n15), .Y(n188) );
  AOI21X2 U133 ( .A0(n186), .A1(B[6]), .B0(n187), .Y(n184) );
  NAND2X2 U134 ( .A(n48), .B(n72), .Y(n178) );
  AOI21X2 U135 ( .A0(n75), .A1(n80), .B0(n69), .Y(n79) );
  INVX2 U136 ( .A(n53), .Y(n190) );
  NAND2X2 U137 ( .A(n146), .B(n147), .Y(n140) );
  NAND2BX4 U138 ( .AN(A[5]), .B(B[5]), .Y(n50) );
  XOR2X2 U139 ( .A(n59), .B(n60), .Y(DIFF[5]) );
  XOR2X4 U140 ( .A(n22), .B(n39), .Y(DIFF[8]) );
  AND3X4 U141 ( .A(n119), .B(n120), .C(n51), .Y(n26) );
  OAI2BB1X4 U142 ( .A0N(n146), .A1N(n159), .B0(n115), .Y(n157) );
  NAND2BX4 U143 ( .AN(A[0]), .B(B[0]), .Y(n73) );
  OAI21X2 U144 ( .A0(n85), .A1(n86), .B0(n87), .Y(n80) );
  AOI21X2 U145 ( .A0(n133), .A1(n142), .B0(n143), .Y(n141) );
  OAI21X1 U146 ( .A0(n113), .A1(n132), .B0(n110), .Y(n135) );
  NAND4BX1 U147 ( .AN(n103), .B(n131), .C(n10), .D(n159), .Y(n130) );
  NAND4X2 U148 ( .A(n75), .B(n68), .C(n73), .D(n196), .Y(n101) );
  XOR2X2 U149 ( .A(n78), .B(n79), .Y(DIFF[3]) );
  OAI21X2 U150 ( .A0(B[6]), .A1(n186), .B0(n54), .Y(n121) );
  NAND2BX4 U151 ( .AN(A[4]), .B(B[4]), .Y(n74) );
  XOR2X4 U152 ( .A(n55), .B(n56), .Y(DIFF[6]) );
  OR2X4 U153 ( .A(n35), .B(n175), .Y(n174) );
  NAND3X4 U154 ( .A(n192), .B(n122), .C(n9), .Y(n77) );
  AOI21X2 U155 ( .A0(n153), .A1(n133), .B0(n154), .Y(n152) );
  INVXL U156 ( .A(n144), .Y(n153) );
  NAND2X4 U157 ( .A(n77), .B(n166), .Y(n41) );
  NAND2BX4 U158 ( .AN(A[14]), .B(B[14]), .Y(n124) );
  XOR2X4 U159 ( .A(n91), .B(n92), .Y(DIFF[16]) );
  XOR2X4 U160 ( .A(n136), .B(n137), .Y(DIFF[14]) );
  NAND2BX4 U161 ( .AN(A[3]), .B(B[3]), .Y(n68) );
  OAI2BB1X4 U162 ( .A0N(n185), .A1N(A[6]), .B0(n54), .Y(n177) );
  NAND2BX4 U163 ( .AN(A[7]), .B(B[7]), .Y(n53) );
  NAND2X2 U164 ( .A(n121), .B(n11), .Y(n156) );
  NAND3X2 U165 ( .A(n162), .B(n31), .C(n163), .Y(n161) );
  NAND3BX2 U166 ( .AN(n33), .B(n34), .C(n2), .Y(n27) );
  NAND2BX4 U167 ( .AN(B[13]), .B(A[13]), .Y(n111) );
  NAND2BX4 U168 ( .AN(A[9]), .B(B[9]), .Y(n31) );
  NAND4BX2 U169 ( .AN(n108), .B(n124), .C(n10), .D(n7), .Y(n102) );
  NAND2X4 U170 ( .A(n159), .B(n5), .Y(n20) );
  NAND2X4 U171 ( .A(n20), .B(n152), .Y(n149) );
  XOR2X4 U172 ( .A(n149), .B(n150), .Y(DIFF[13]) );
  NOR2BX4 U173 ( .AN(n52), .B(n57), .Y(n56) );
  AND2X1 U174 ( .A(n119), .B(n51), .Y(n169) );
  NAND2XL U175 ( .A(n110), .B(n111), .Y(n106) );
  INVXL U176 ( .A(B[6]), .Y(n185) );
  INVXL U177 ( .A(n75), .Y(n83) );
  AND2X1 U178 ( .A(n13), .B(n38), .Y(n22) );
  INVXL U179 ( .A(n52), .Y(n45) );
  AND2X1 U180 ( .A(n97), .B(n127), .Y(n24) );
  NOR2XL U181 ( .A(n103), .B(n104), .Y(n99) );
  NAND2BXL U182 ( .AN(n111), .B(n124), .Y(n128) );
  OAI21X1 U183 ( .A0(n105), .A1(n106), .B0(n107), .Y(n96) );
  NOR2BX2 U184 ( .AN(n68), .B(n67), .Y(n66) );
  AOI31X1 U185 ( .A0(n116), .A1(n68), .A2(n117), .B0(n118), .Y(n114) );
  NAND3X1 U186 ( .A(n122), .B(n84), .C(n65), .Y(n116) );
  INVX1 U187 ( .A(n104), .Y(n117) );
  INVX1 U188 ( .A(n31), .Y(n30) );
  NOR2X2 U189 ( .A(n61), .B(n58), .Y(n60) );
  NAND2X2 U190 ( .A(n145), .B(n133), .Y(n115) );
  OAI2BB1X2 U191 ( .A0N(n64), .A1N(n65), .B0(n66), .Y(n63) );
  NOR2X2 U192 ( .A(n69), .B(n70), .Y(n64) );
  NAND2X1 U193 ( .A(n99), .B(n100), .Y(n98) );
  NAND4BXL U194 ( .AN(n190), .B(n51), .C(n17), .D(n50), .Y(n104) );
  NAND2X1 U195 ( .A(n90), .B(n73), .Y(DIFF[0]) );
  XOR2X2 U196 ( .A(n80), .B(n82), .Y(DIFF[2]) );
  NOR2XL U197 ( .A(n108), .B(n109), .Y(n107) );
  NAND2BX1 U198 ( .AN(n73), .B(n90), .Y(n88) );
  INVXL U199 ( .A(A[6]), .Y(n186) );
  INVX2 U200 ( .A(A[1]), .Y(n197) );
  NAND2BX2 U201 ( .AN(A[5]), .B(B[5]), .Y(n119) );
  NAND2XL U202 ( .A(n68), .B(n81), .Y(n78) );
  XOR2X1 U203 ( .A(B[16]), .B(A[16]), .Y(n92) );
  NAND2BX1 U204 ( .AN(B[6]), .B(A[6]), .Y(n52) );
  XOR2X4 U205 ( .A(n27), .B(n28), .Y(DIFF[9]) );
  XOR2X4 U206 ( .A(n43), .B(n44), .Y(DIFF[7]) );
  NOR2X4 U207 ( .A(n45), .B(n46), .Y(n44) );
  NAND2BX4 U208 ( .AN(n62), .B(n63), .Y(n59) );
  NAND2BX4 U209 ( .AN(A[12]), .B(B[12]), .Y(n125) );
  CLKINVX3 U210 ( .A(n113), .Y(n154) );
  NAND2BX4 U211 ( .AN(B[12]), .B(A[12]), .Y(n113) );
  NAND2BX4 U212 ( .AN(n160), .B(n161), .Y(n133) );
  OAI21X4 U213 ( .A0(n183), .A1(A[8]), .B0(n53), .Y(n36) );
  NAND2BX4 U214 ( .AN(B[4]), .B(A[4]), .Y(n72) );
  NAND2X4 U215 ( .A(n188), .B(n189), .Y(n35) );
endmodule


module butterfly_DW01_add_151 ( A, B, SUM );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  wire   n212, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211;

  BUFX3 U2 ( .A(n6), .Y(n12) );
  NAND3X4 U3 ( .A(A[12]), .B(B[12]), .C(n142), .Y(n164) );
  AND2X2 U4 ( .A(B[10]), .B(A[10]), .Y(n25) );
  AOI21X2 U5 ( .A0(n143), .A1(n144), .B0(n145), .Y(n122) );
  NAND2X4 U6 ( .A(n207), .B(n209), .Y(n1) );
  NAND2X4 U7 ( .A(n2), .B(n38), .Y(n99) );
  INVX4 U8 ( .A(n1), .Y(n2) );
  NAND3BX4 U9 ( .AN(n126), .B(n172), .C(n45), .Y(n3) );
  CLKINVX3 U10 ( .A(n80), .Y(n172) );
  NAND2XL U11 ( .A(n133), .B(n134), .Y(n131) );
  INVX20 U12 ( .A(n53), .Y(n7) );
  INVX2 U13 ( .A(n25), .Y(n4) );
  NAND2BX4 U14 ( .AN(B[11]), .B(n46), .Y(n36) );
  NAND2X4 U15 ( .A(n206), .B(n205), .Y(n5) );
  NOR2BX4 U16 ( .AN(n115), .B(n119), .Y(n205) );
  NAND2BXL U17 ( .AN(n4), .B(n36), .Y(n6) );
  CLKINVX3 U18 ( .A(n200), .Y(n9) );
  AND2X2 U19 ( .A(B[4]), .B(A[4]), .Y(n200) );
  AND2X2 U20 ( .A(B[0]), .B(A[0]), .Y(n31) );
  NAND2X4 U21 ( .A(n89), .B(n87), .Y(n151) );
  NAND2X2 U22 ( .A(B[4]), .B(A[4]), .Y(n102) );
  NAND2X4 U23 ( .A(n169), .B(n7), .Y(n62) );
  INVX4 U24 ( .A(n40), .Y(n16) );
  OR2X4 U25 ( .A(B[8]), .B(A[8]), .Y(n185) );
  INVX4 U26 ( .A(n22), .Y(n183) );
  AND2X4 U27 ( .A(n146), .B(n147), .Y(n8) );
  BUFX12 U28 ( .A(n212), .Y(SUM[12]) );
  NAND2X1 U29 ( .A(n141), .B(n142), .Y(n165) );
  OR2X4 U30 ( .A(A[12]), .B(B[12]), .Y(n141) );
  NOR2X1 U31 ( .A(n150), .B(n40), .Y(n193) );
  NOR2BX2 U32 ( .AN(n112), .B(n111), .Y(n114) );
  CLKINVX8 U33 ( .A(n207), .Y(n111) );
  INVX8 U34 ( .A(A[11]), .Y(n46) );
  NOR4X4 U35 ( .A(n91), .B(n54), .C(n21), .D(n175), .Y(n43) );
  INVX2 U36 ( .A(n133), .Y(n53) );
  NAND2X1 U37 ( .A(B[12]), .B(A[12]), .Y(n133) );
  XOR2X2 U38 ( .A(n114), .B(n113), .Y(SUM[2]) );
  NOR4BX2 U39 ( .AN(n84), .B(n175), .C(n54), .D(n21), .Y(n22) );
  INVXL U40 ( .A(A[5]), .Y(n15) );
  INVX1 U41 ( .A(n48), .Y(n19) );
  INVX1 U42 ( .A(A[4]), .Y(n54) );
  CLKINVX3 U43 ( .A(n57), .Y(n58) );
  INVX1 U44 ( .A(n94), .Y(n60) );
  INVX1 U45 ( .A(A[6]), .Y(n32) );
  NAND2XL U46 ( .A(n164), .B(n134), .Y(n167) );
  NAND2X1 U47 ( .A(B[15]), .B(A[15]), .Y(n129) );
  OR2X2 U48 ( .A(A[15]), .B(B[15]), .Y(n139) );
  CLKINVX3 U49 ( .A(n31), .Y(n119) );
  BUFX3 U50 ( .A(n73), .Y(n41) );
  INVX1 U51 ( .A(n47), .Y(n52) );
  NAND2X1 U52 ( .A(n137), .B(n138), .Y(n123) );
  INVX2 U53 ( .A(n89), .Y(n184) );
  NAND2X1 U54 ( .A(n42), .B(n89), .Y(n82) );
  NOR2BX2 U55 ( .AN(n9), .B(n105), .Y(n107) );
  AND2X4 U56 ( .A(n102), .B(n101), .Y(n10) );
  NAND2X1 U57 ( .A(n129), .B(n139), .Y(n11) );
  INVX1 U58 ( .A(B[4]), .Y(n21) );
  INVXL U59 ( .A(n91), .Y(n13) );
  NAND3X2 U60 ( .A(n74), .B(n41), .C(n72), .Y(n69) );
  INVX4 U61 ( .A(n79), .Y(n45) );
  NAND4X4 U62 ( .A(n67), .B(n16), .C(n34), .D(n20), .Y(n14) );
  NAND3BX4 U63 ( .AN(n15), .B(n58), .C(n84), .Y(n152) );
  NOR2X4 U64 ( .A(B[8]), .B(A[8]), .Y(n40) );
  AND2X2 U65 ( .A(n163), .B(n161), .Y(n65) );
  OR2X2 U66 ( .A(B[7]), .B(A[7]), .Y(n17) );
  AOI21X2 U67 ( .A0(n72), .A1(n191), .B0(n192), .Y(n190) );
  OAI21X2 U68 ( .A0(n193), .A1(n194), .B0(n195), .Y(n192) );
  OR2X4 U69 ( .A(n60), .B(n59), .Y(n18) );
  NOR2X4 U70 ( .A(n92), .B(n93), .Y(n59) );
  NOR2X2 U71 ( .A(n56), .B(n47), .Y(n195) );
  NAND2X4 U72 ( .A(n201), .B(n19), .Y(n50) );
  INVX2 U73 ( .A(n71), .Y(n48) );
  NAND2BX2 U74 ( .AN(n75), .B(n76), .Y(n74) );
  NAND2X4 U75 ( .A(n24), .B(n23), .Y(n20) );
  OAI21X4 U76 ( .A0(n118), .A1(n119), .B0(n116), .Y(n113) );
  NAND2X1 U77 ( .A(B[1]), .B(A[1]), .Y(n116) );
  INVX2 U78 ( .A(n25), .Y(n33) );
  OR2X4 U79 ( .A(B[10]), .B(A[10]), .Y(n27) );
  NAND2BX4 U80 ( .AN(n151), .B(n152), .Y(n210) );
  NAND2X4 U81 ( .A(n23), .B(n24), .Y(n186) );
  INVX4 U82 ( .A(B[9]), .Y(n23) );
  INVX1 U83 ( .A(A[9]), .Y(n24) );
  NAND2X2 U84 ( .A(n99), .B(n100), .Y(n98) );
  NAND2X4 U85 ( .A(n99), .B(n100), .Y(n155) );
  NAND2BX4 U86 ( .AN(n112), .B(n38), .Y(n100) );
  DLY1X1 U87 ( .A(n148), .Y(n37) );
  XNOR2X4 U88 ( .A(n62), .B(n26), .Y(SUM[13]) );
  NAND2XL U89 ( .A(n142), .B(n134), .Y(n26) );
  NAND2X2 U90 ( .A(n170), .B(n171), .Y(n49) );
  NAND3X2 U91 ( .A(n200), .B(n96), .C(n84), .Y(n153) );
  NAND2BX4 U92 ( .AN(B[11]), .B(n46), .Y(n180) );
  INVX1 U93 ( .A(B[5]), .Y(n57) );
  NAND2X4 U94 ( .A(n10), .B(n103), .Y(n97) );
  NAND2XL U95 ( .A(n5), .B(n101), .Y(n154) );
  NOR2XL U96 ( .A(n154), .B(n155), .Y(n149) );
  OR2X4 U97 ( .A(B[5]), .B(A[5]), .Y(n28) );
  AND3X2 U98 ( .A(A[5]), .B(n58), .C(n84), .Y(n55) );
  AND2X2 U99 ( .A(n119), .B(n29), .Y(SUM[0]) );
  OR2XL U100 ( .A(A[0]), .B(B[0]), .Y(n29) );
  INVXL U101 ( .A(n56), .Y(n30) );
  NOR2BX4 U102 ( .AN(n32), .B(B[6]), .Y(n68) );
  NAND4X4 U103 ( .A(n67), .B(n16), .C(n34), .D(n20), .Y(n126) );
  OR2X4 U104 ( .A(B[11]), .B(A[11]), .Y(n34) );
  DLY1X1 U105 ( .A(n126), .Y(n35) );
  INVX1 U106 ( .A(n33), .Y(n189) );
  OR2X4 U107 ( .A(A[1]), .B(B[1]), .Y(n115) );
  XNOR2X4 U108 ( .A(n158), .B(n64), .Y(n212) );
  INVX4 U109 ( .A(n115), .Y(n118) );
  OR2X4 U110 ( .A(A[3]), .B(B[3]), .Y(n38) );
  AND2X1 U111 ( .A(B[8]), .B(A[8]), .Y(n39) );
  INVX8 U112 ( .A(n150), .Y(n42) );
  AND2X2 U113 ( .A(n52), .B(n33), .Y(n51) );
  NOR2X4 U114 ( .A(n110), .B(n111), .Y(n206) );
  INVX8 U115 ( .A(n208), .Y(n110) );
  INVX8 U116 ( .A(n84), .Y(n91) );
  INVX8 U117 ( .A(n28), .Y(n175) );
  NAND2BX1 U118 ( .AN(n199), .B(n84), .Y(n198) );
  XOR2X4 U119 ( .A(n45), .B(n107), .Y(SUM[4]) );
  NOR2BX2 U120 ( .AN(n116), .B(n118), .Y(n117) );
  INVX8 U121 ( .A(n106), .Y(n79) );
  OAI2BB1X4 U122 ( .A0N(n113), .A1N(n207), .B0(n112), .Y(n108) );
  INVXL U123 ( .A(n35), .Y(n144) );
  NOR2BX2 U124 ( .AN(n71), .B(n56), .Y(n70) );
  NAND2X1 U125 ( .A(n28), .B(n200), .Y(n197) );
  INVX8 U126 ( .A(n186), .Y(n56) );
  NOR2BX2 U127 ( .AN(n41), .B(n40), .Y(n78) );
  NAND2X4 U128 ( .A(n202), .B(n30), .Y(n201) );
  OR2X2 U129 ( .A(B[4]), .B(A[4]), .Y(n95) );
  XOR2X4 U130 ( .A(n120), .B(n121), .Y(SUM[16]) );
  AOI21X2 U131 ( .A0(n130), .A1(n131), .B0(n132), .Y(n127) );
  NAND2X1 U132 ( .A(B[5]), .B(A[5]), .Y(n94) );
  NOR2X2 U133 ( .A(B[10]), .B(A[10]), .Y(n47) );
  AOI21X4 U134 ( .A0(n158), .A1(n157), .B0(n159), .Y(n156) );
  NAND2X4 U135 ( .A(n71), .B(n73), .Y(n194) );
  XOR2X4 U136 ( .A(n50), .B(n51), .Y(SUM[10]) );
  NAND2X2 U137 ( .A(B[11]), .B(A[11]), .Y(n147) );
  NAND3XL U138 ( .A(n37), .B(n12), .C(n147), .Y(n145) );
  NAND2XL U139 ( .A(n147), .B(n36), .Y(n187) );
  XOR2X4 U140 ( .A(n108), .B(n109), .Y(SUM[3]) );
  NAND2X4 U141 ( .A(n49), .B(n141), .Y(n169) );
  NAND2X4 U142 ( .A(B[10]), .B(A[10]), .Y(n181) );
  INVX8 U143 ( .A(n88), .Y(n150) );
  AND2X4 U144 ( .A(n17), .B(n84), .Y(n61) );
  NAND2X2 U145 ( .A(n95), .B(n96), .Y(n93) );
  NAND3BX4 U146 ( .AN(n39), .B(n203), .C(n72), .Y(n202) );
  OR2X4 U147 ( .A(n179), .B(n151), .Y(n66) );
  NAND3BX4 U148 ( .AN(n55), .B(n182), .C(n183), .Y(n177) );
  OAI21X4 U149 ( .A0(n43), .A1(n210), .B0(n211), .Y(n203) );
  NOR2X4 U150 ( .A(n175), .B(n105), .Y(n204) );
  XOR2X4 U151 ( .A(n156), .B(n11), .Y(SUM[15]) );
  NOR2X4 U152 ( .A(n66), .B(n196), .Y(n191) );
  OAI2BB1X4 U153 ( .A0N(n160), .A1N(n161), .B0(n162), .Y(n159) );
  NAND2X4 U154 ( .A(A[7]), .B(B[7]), .Y(n89) );
  INVX4 U155 ( .A(n75), .Y(n211) );
  NAND2X4 U156 ( .A(n42), .B(n185), .Y(n75) );
  OAI21X2 U157 ( .A0(n197), .A1(n91), .B0(n198), .Y(n196) );
  NAND3BX4 U158 ( .AN(n126), .B(n172), .C(n45), .Y(n171) );
  NAND2X4 U159 ( .A(n148), .B(n8), .Y(n178) );
  NOR2X4 U160 ( .A(n14), .B(n150), .Y(n176) );
  AOI2BB1X4 U161 ( .A0N(n135), .A1N(n134), .B0(n132), .Y(n162) );
  NOR2X2 U162 ( .A(n128), .B(n135), .Y(n138) );
  NOR2X1 U163 ( .A(n135), .B(n136), .Y(n130) );
  OAI21X2 U164 ( .A0(n127), .A1(n128), .B0(n129), .Y(n125) );
  NAND4X4 U165 ( .A(n106), .B(n61), .C(n185), .D(n204), .Y(n72) );
  NOR2BX2 U166 ( .AN(n101), .B(n110), .Y(n109) );
  NAND2X2 U167 ( .A(B[3]), .B(A[3]), .Y(n101) );
  NOR2X4 U168 ( .A(n97), .B(n98), .Y(n92) );
  XOR2X2 U169 ( .A(n31), .B(n117), .Y(SUM[1]) );
  NOR2X4 U170 ( .A(n190), .B(n189), .Y(n188) );
  NOR2BX2 U171 ( .AN(n87), .B(n91), .Y(n90) );
  NAND2X4 U172 ( .A(B[6]), .B(A[6]), .Y(n87) );
  CLKINVX8 U173 ( .A(n161), .Y(n135) );
  INVX2 U174 ( .A(n164), .Y(n160) );
  NAND2BX4 U175 ( .AN(n181), .B(n180), .Y(n146) );
  INVX8 U176 ( .A(n68), .Y(n84) );
  NAND4BX4 U177 ( .AN(n56), .B(n36), .C(n27), .D(n194), .Y(n148) );
  INVX8 U178 ( .A(n95), .Y(n105) );
  INVX2 U179 ( .A(n125), .Y(n124) );
  NAND2X2 U180 ( .A(B[13]), .B(A[13]), .Y(n134) );
  NAND2X2 U181 ( .A(n133), .B(n141), .Y(n64) );
  XOR2X4 U182 ( .A(n188), .B(n187), .Y(SUM[11]) );
  OAI21X2 U183 ( .A0(n79), .A1(n80), .B0(n81), .Y(n77) );
  XOR2X4 U184 ( .A(n104), .B(n63), .Y(SUM[5]) );
  OAI21X4 U185 ( .A0(n79), .A1(n105), .B0(n9), .Y(n104) );
  AOI21X4 U186 ( .A0(n176), .A1(n177), .B0(n178), .Y(n170) );
  XOR2X4 U187 ( .A(n18), .B(n90), .Y(SUM[6]) );
  NOR2X4 U188 ( .A(n150), .B(n91), .Y(n174) );
  NAND2X4 U189 ( .A(A[9]), .B(B[9]), .Y(n71) );
  OAI21X4 U190 ( .A0(n122), .A1(n123), .B0(n124), .Y(n120) );
  XOR2X4 U191 ( .A(n83), .B(n82), .Y(SUM[7]) );
  AOI21X4 U192 ( .A0(n13), .A1(n85), .B0(n86), .Y(n83) );
  NAND2BX4 U193 ( .AN(n150), .B(n76), .Y(n81) );
  NAND3BX4 U194 ( .AN(n151), .B(n152), .C(n153), .Y(n76) );
  OR2X4 U195 ( .A(A[13]), .B(B[13]), .Y(n142) );
  OR2X4 U196 ( .A(n59), .B(n60), .Y(n85) );
  OR2X4 U197 ( .A(B[10]), .B(A[10]), .Y(n67) );
  NOR2X2 U198 ( .A(n175), .B(n105), .Y(n173) );
  NAND2X2 U199 ( .A(B[2]), .B(A[2]), .Y(n112) );
  NAND2BX2 U200 ( .AN(n165), .B(n158), .Y(n168) );
  AND2X1 U201 ( .A(n94), .B(n96), .Y(n63) );
  INVX4 U202 ( .A(n163), .Y(n132) );
  XOR2X4 U203 ( .A(n166), .B(n65), .Y(SUM[14]) );
  INVXL U204 ( .A(n142), .Y(n136) );
  NOR2XL U205 ( .A(n136), .B(n140), .Y(n137) );
  NAND2X2 U206 ( .A(n71), .B(n73), .Y(n179) );
  INVX1 U207 ( .A(n139), .Y(n128) );
  INVX1 U208 ( .A(n141), .Y(n140) );
  NOR2X2 U209 ( .A(n86), .B(n184), .Y(n182) );
  XOR2X1 U210 ( .A(B[16]), .B(A[16]), .Y(n121) );
  NAND3BX4 U211 ( .AN(n155), .B(n5), .C(n101), .Y(n106) );
  NOR2X2 U212 ( .A(n165), .B(n135), .Y(n157) );
  OAI21XL U213 ( .A0(n149), .A1(n80), .B0(n81), .Y(n143) );
  NAND2X1 U214 ( .A(B[14]), .B(A[14]), .Y(n163) );
  NAND2XL U215 ( .A(A[5]), .B(B[5]), .Y(n199) );
  XOR2X4 U216 ( .A(n69), .B(n70), .Y(SUM[9]) );
  XOR2X4 U217 ( .A(n77), .B(n78), .Y(SUM[8]) );
  CLKINVX3 U218 ( .A(n87), .Y(n86) );
  OR2X4 U219 ( .A(A[14]), .B(B[14]), .Y(n161) );
  NAND2BX4 U220 ( .AN(n167), .B(n168), .Y(n166) );
  NAND2X4 U221 ( .A(n170), .B(n3), .Y(n158) );
  NAND2X4 U222 ( .A(n173), .B(n174), .Y(n80) );
  NAND2X4 U223 ( .A(n206), .B(n205), .Y(n103) );
  AND2X2 U224 ( .A(B[1]), .B(A[1]), .Y(n209) );
  OR2X4 U225 ( .A(A[2]), .B(B[2]), .Y(n207) );
  OR2X4 U226 ( .A(A[3]), .B(B[3]), .Y(n208) );
  OR2X4 U227 ( .A(B[7]), .B(A[7]), .Y(n88) );
  OR2X4 U228 ( .A(B[5]), .B(A[5]), .Y(n96) );
  NAND2X4 U229 ( .A(A[8]), .B(B[8]), .Y(n73) );
endmodule


module butterfly_DW01_add_141 ( A, B, SUM );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  wire   n187, n188, n189, n190, n1, n2, n3, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n40, n41, n43,
         n44, n45, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186;

  NOR2X4 U2 ( .A(n185), .B(n186), .Y(n184) );
  BUFX3 U3 ( .A(n158), .Y(n8) );
  NAND2X1 U4 ( .A(n27), .B(n118), .Y(n158) );
  NAND2X4 U5 ( .A(n119), .B(n118), .Y(n117) );
  NOR2BX1 U6 ( .AN(n85), .B(n2), .Y(n87) );
  NAND2X4 U7 ( .A(n51), .B(n1), .Y(n106) );
  AND2X4 U8 ( .A(n52), .B(n18), .Y(n1) );
  INVX1 U9 ( .A(n114), .Y(n24) );
  CLKBUFX3 U10 ( .A(n65), .Y(n30) );
  NOR2X4 U11 ( .A(A[4]), .B(B[4]), .Y(n2) );
  INVX4 U12 ( .A(n67), .Y(n66) );
  OAI2BB1X4 U13 ( .A0N(n17), .A1N(n66), .B0(n178), .Y(n14) );
  OR2X2 U14 ( .A(A[14]), .B(B[14]), .Y(n27) );
  OR2X4 U15 ( .A(B[10]), .B(A[10]), .Y(n3) );
  INVX8 U16 ( .A(n152), .Y(n168) );
  NAND2X2 U17 ( .A(n27), .B(n115), .Y(n112) );
  BUFX3 U18 ( .A(n190), .Y(SUM[4]) );
  AOI2BB1X2 U19 ( .A0N(n50), .A1N(n109), .B0(n151), .Y(n146) );
  XOR2X2 U20 ( .A(n88), .B(n89), .Y(SUM[3]) );
  NOR2BX1 U21 ( .AN(n90), .B(n91), .Y(n89) );
  NOR3X2 U22 ( .A(n186), .B(n78), .C(n85), .Y(n156) );
  INVX3 U23 ( .A(n16), .Y(n78) );
  NAND3X1 U24 ( .A(A[1]), .B(B[1]), .C(n97), .Y(n183) );
  CLKINVX3 U25 ( .A(n65), .Y(n73) );
  OAI21X2 U26 ( .A0(n79), .A1(n80), .B0(n81), .Y(n75) );
  INVX1 U27 ( .A(n177), .Y(n17) );
  INVX4 U28 ( .A(n73), .Y(n19) );
  INVX1 U29 ( .A(n163), .Y(n20) );
  INVX1 U30 ( .A(n120), .Y(n37) );
  INVX1 U31 ( .A(n31), .Y(n32) );
  NAND2X1 U32 ( .A(B[0]), .B(A[0]), .Y(n103) );
  XOR2X1 U33 ( .A(n21), .B(n87), .Y(n190) );
  INVX1 U34 ( .A(n71), .Y(n23) );
  NOR2BX1 U35 ( .AN(n127), .B(n176), .Y(n175) );
  NOR2BX2 U36 ( .AN(n63), .B(n61), .Y(n69) );
  OR2X4 U37 ( .A(A[13]), .B(B[13]), .Y(n123) );
  CLKINVX3 U38 ( .A(n137), .Y(n91) );
  XOR2X4 U39 ( .A(n57), .B(n58), .Y(n5) );
  NOR2X4 U40 ( .A(n33), .B(n120), .Y(n116) );
  NAND2XL U41 ( .A(n113), .B(n115), .Y(n145) );
  NAND2X4 U42 ( .A(A[13]), .B(B[13]), .Y(n119) );
  NOR2X1 U43 ( .A(B[6]), .B(A[6]), .Y(n185) );
  BUFX8 U44 ( .A(n16), .Y(n6) );
  NOR2BXL U45 ( .AN(n76), .B(n78), .Y(n77) );
  NOR2X2 U46 ( .A(n163), .B(n33), .Y(n160) );
  INVX2 U47 ( .A(n122), .Y(n163) );
  NOR2X4 U48 ( .A(n7), .B(n2), .Y(n26) );
  NOR2X2 U49 ( .A(B[7]), .B(A[7]), .Y(n7) );
  INVX4 U50 ( .A(n64), .Y(n11) );
  CLKBUFX8 U51 ( .A(n72), .Y(n29) );
  NOR2BX4 U52 ( .AN(n19), .B(n177), .Y(n179) );
  OAI2BB1X2 U53 ( .A0N(n6), .A1N(n75), .B0(n76), .Y(n70) );
  OR2X2 U54 ( .A(B[11]), .B(A[11]), .Y(n43) );
  NAND2X1 U55 ( .A(n18), .B(n142), .Y(n53) );
  OR2X4 U56 ( .A(A[13]), .B(B[13]), .Y(n9) );
  XOR2X2 U57 ( .A(n75), .B(n77), .Y(SUM[6]) );
  OR2X4 U58 ( .A(A[11]), .B(B[11]), .Y(n10) );
  NOR2BX2 U59 ( .AN(n142), .B(n143), .Y(n124) );
  BUFX3 U60 ( .A(n10), .Y(n18) );
  NAND3X1 U61 ( .A(n114), .B(n9), .C(n122), .Y(n147) );
  OAI2BB1X4 U62 ( .A0N(n120), .A1N(n119), .B0(n9), .Y(n162) );
  OAI2BB1X2 U63 ( .A0N(B[5]), .A1N(A[5]), .B0(n76), .Y(n173) );
  OR2X2 U64 ( .A(A[5]), .B(B[5]), .Y(n141) );
  NOR2X4 U65 ( .A(n11), .B(n12), .Y(n13) );
  NOR2X2 U66 ( .A(n13), .B(n66), .Y(n62) );
  INVX1 U67 ( .A(n30), .Y(n12) );
  BUFX20 U68 ( .A(n187), .Y(SUM[15]) );
  INVX12 U69 ( .A(n132), .Y(n61) );
  BUFX4 U70 ( .A(B[5]), .Y(n25) );
  INVXL U71 ( .A(n34), .Y(n15) );
  INVX2 U72 ( .A(n162), .Y(n149) );
  OR2X4 U73 ( .A(A[6]), .B(B[6]), .Y(n16) );
  NOR2X2 U74 ( .A(n110), .B(n84), .Y(n44) );
  NAND2X4 U75 ( .A(n59), .B(n63), .Y(n169) );
  NOR2BX4 U76 ( .AN(n140), .B(n91), .Y(n21) );
  NAND2X4 U77 ( .A(n132), .B(n60), .Y(n177) );
  INVX8 U78 ( .A(n5), .Y(SUM[9]) );
  NOR2X4 U79 ( .A(B[9]), .B(A[9]), .Y(n34) );
  NAND3X4 U80 ( .A(n28), .B(n43), .C(n131), .Y(n109) );
  XNOR2X4 U81 ( .A(n70), .B(n23), .Y(SUM[7]) );
  AOI2BB1X4 U82 ( .A0N(n162), .A1N(n24), .B0(n150), .Y(n148) );
  NOR2X2 U83 ( .A(n186), .B(n85), .Y(n172) );
  OR2X4 U84 ( .A(n143), .B(n168), .Y(n151) );
  NOR2BX1 U85 ( .AN(n81), .B(n80), .Y(n83) );
  NAND2X4 U86 ( .A(n26), .B(n184), .Y(n110) );
  AND2X4 U87 ( .A(n60), .B(n132), .Y(n28) );
  INVXL U88 ( .A(n3), .Y(n176) );
  INVXL U89 ( .A(n129), .Y(n31) );
  NAND2X2 U90 ( .A(A[15]), .B(B[15]), .Y(n113) );
  NOR2X2 U91 ( .A(B[13]), .B(A[13]), .Y(n33) );
  NAND2X4 U92 ( .A(A[9]), .B(B[9]), .Y(n59) );
  NAND2X4 U93 ( .A(A[11]), .B(B[11]), .Y(n142) );
  NAND2X2 U94 ( .A(n74), .B(n141), .Y(n138) );
  XOR2X2 U95 ( .A(n14), .B(n175), .Y(SUM[10]) );
  AND2X4 U96 ( .A(n123), .B(n122), .Y(n52) );
  NAND2X4 U97 ( .A(A[10]), .B(B[10]), .Y(n127) );
  NOR2X4 U98 ( .A(n116), .B(n117), .Y(n111) );
  NAND2BX4 U99 ( .AN(n110), .B(n21), .Y(n155) );
  INVXL U100 ( .A(n141), .Y(n80) );
  NOR2X4 U101 ( .A(A[5]), .B(B[5]), .Y(n186) );
  NAND2X4 U102 ( .A(n35), .B(n36), .Y(n45) );
  AND2X4 U103 ( .A(n6), .B(n65), .Y(n35) );
  OR2X4 U104 ( .A(n172), .B(n173), .Y(n36) );
  NAND2BX4 U105 ( .AN(n37), .B(n165), .Y(n49) );
  BUFX20 U106 ( .A(n188), .Y(SUM[13]) );
  XNOR2X2 U107 ( .A(n161), .B(n38), .Y(n189) );
  NAND2XL U108 ( .A(n120), .B(n122), .Y(n38) );
  OAI2BB1X2 U109 ( .A0N(n19), .A1N(n64), .B0(n67), .Y(n68) );
  OR2X4 U110 ( .A(A[10]), .B(B[10]), .Y(n131) );
  NAND2X4 U111 ( .A(n181), .B(n6), .Y(n136) );
  NOR2X2 U112 ( .A(n85), .B(n186), .Y(n181) );
  NAND2X4 U113 ( .A(A[6]), .B(B[6]), .Y(n76) );
  OAI21X4 U114 ( .A0(n111), .A1(n112), .B0(n113), .Y(n108) );
  AOI21X4 U115 ( .A0(n64), .A1(n179), .B0(n180), .Y(n178) );
  OAI21X2 U116 ( .A0(n157), .A1(n156), .B0(n30), .Y(n154) );
  AOI21X4 U117 ( .A0(n128), .A1(n32), .B0(n130), .Y(n125) );
  NAND2X4 U118 ( .A(B[2]), .B(A[2]), .Y(n94) );
  XOR2X4 U119 ( .A(n104), .B(n41), .Y(n40) );
  XNOR2X4 U120 ( .A(B[16]), .B(A[16]), .Y(n41) );
  INVX4 U121 ( .A(n108), .Y(n107) );
  NAND4BX2 U122 ( .AN(n34), .B(n131), .C(n132), .D(n19), .Y(n130) );
  NAND3X2 U123 ( .A(n72), .B(n76), .C(n136), .Y(n135) );
  OR2X4 U124 ( .A(A[8]), .B(B[8]), .Y(n132) );
  INVX8 U125 ( .A(n153), .Y(n143) );
  AND2X4 U126 ( .A(n115), .B(n114), .Y(n51) );
  NAND3X4 U127 ( .A(n54), .B(n182), .C(n183), .Y(n140) );
  AND2X4 U128 ( .A(n94), .B(n90), .Y(n54) );
  NAND2XL U129 ( .A(n9), .B(n119), .Y(n164) );
  INVX2 U130 ( .A(n69), .Y(n48) );
  OAI21X1 U131 ( .A0(n34), .A1(n63), .B0(n59), .Y(n180) );
  NAND3X4 U132 ( .A(n74), .B(n25), .C(A[5]), .Y(n129) );
  AOI21X4 U133 ( .A0(n133), .A1(n134), .B0(n135), .Y(n128) );
  NAND4BX4 U134 ( .AN(n34), .B(n121), .C(n170), .D(n169), .Y(n153) );
  OAI2BB1X4 U135 ( .A0N(n127), .A1N(n142), .B0(n10), .Y(n152) );
  BUFX12 U136 ( .A(n189), .Y(SUM[12]) );
  AND3X4 U137 ( .A(n154), .B(n155), .C(n29), .Y(n50) );
  NAND2X1 U138 ( .A(n76), .B(n129), .Y(n157) );
  NAND2X4 U139 ( .A(n20), .B(n161), .Y(n165) );
  NOR3BX4 U140 ( .AN(n124), .B(n125), .C(n126), .Y(n105) );
  NOR2X4 U141 ( .A(n44), .B(n171), .Y(n166) );
  NAND2X4 U142 ( .A(n45), .B(n29), .Y(n171) );
  NAND2X2 U143 ( .A(A[7]), .B(B[7]), .Y(n72) );
  INVX8 U144 ( .A(n40), .Y(SUM[16]) );
  XNOR2X4 U145 ( .A(n68), .B(n48), .Y(SUM[8]) );
  NAND2X4 U146 ( .A(B[8]), .B(A[8]), .Y(n63) );
  OR2X1 U147 ( .A(A[3]), .B(B[3]), .Y(n137) );
  XOR2X4 U148 ( .A(n174), .B(n53), .Y(SUM[11]) );
  NAND2X2 U149 ( .A(B[14]), .B(A[14]), .Y(n118) );
  OAI21X4 U150 ( .A0(n2), .A1(n84), .B0(n85), .Y(n82) );
  INVX4 U151 ( .A(n86), .Y(n84) );
  XNOR2X4 U152 ( .A(n49), .B(n164), .Y(n188) );
  NAND2X4 U153 ( .A(B[4]), .B(A[4]), .Y(n85) );
  NAND2XL U154 ( .A(n59), .B(n15), .Y(n58) );
  INVXL U155 ( .A(n97), .Y(n93) );
  NOR2BX1 U156 ( .AN(n103), .B(n55), .Y(SUM[0]) );
  NOR2XL U157 ( .A(A[0]), .B(B[0]), .Y(n55) );
  NOR2BX1 U158 ( .AN(n29), .B(n73), .Y(n71) );
  XOR2X1 U159 ( .A(n82), .B(n83), .Y(SUM[5]) );
  INVX1 U160 ( .A(n127), .Y(n126) );
  XNOR2X4 U161 ( .A(n144), .B(n145), .Y(n187) );
  NAND2X4 U162 ( .A(n56), .B(n136), .Y(n64) );
  AND3X4 U163 ( .A(n129), .B(n76), .C(n72), .Y(n56) );
  INVX1 U164 ( .A(n118), .Y(n150) );
  NOR2X2 U165 ( .A(n91), .B(n2), .Y(n134) );
  NOR2X1 U166 ( .A(n138), .B(n139), .Y(n133) );
  NOR2BX4 U167 ( .AN(n140), .B(n91), .Y(n86) );
  OAI21XL U168 ( .A0(n92), .A1(n93), .B0(n94), .Y(n88) );
  INVX1 U169 ( .A(n95), .Y(n92) );
  XOR2X1 U170 ( .A(n95), .B(n96), .Y(SUM[2]) );
  NOR2BX1 U171 ( .AN(n94), .B(n93), .Y(n96) );
  XOR2X1 U172 ( .A(n99), .B(n101), .Y(SUM[1]) );
  NOR2BX1 U173 ( .AN(n100), .B(n102), .Y(n101) );
  INVX1 U174 ( .A(n98), .Y(n102) );
  OAI2BB1X1 U175 ( .A0N(n98), .A1N(n99), .B0(n100), .Y(n95) );
  INVX1 U176 ( .A(n140), .Y(n139) );
  INVX1 U177 ( .A(n103), .Y(n99) );
  NAND2XL U178 ( .A(n25), .B(A[5]), .Y(n81) );
  NAND3BX1 U179 ( .AN(n103), .B(n97), .C(n98), .Y(n182) );
  NAND2X2 U180 ( .A(B[3]), .B(A[3]), .Y(n90) );
  NAND2XL U181 ( .A(B[1]), .B(A[1]), .Y(n100) );
  OAI21X4 U182 ( .A0(n61), .A1(n62), .B0(n63), .Y(n57) );
  CLKINVX3 U183 ( .A(n82), .Y(n79) );
  OAI21X4 U184 ( .A0(n106), .A1(n105), .B0(n107), .Y(n104) );
  OR2X4 U185 ( .A(B[15]), .B(A[15]), .Y(n115) );
  OAI21X4 U186 ( .A0(n146), .A1(n147), .B0(n148), .Y(n144) );
  XOR2X4 U187 ( .A(n159), .B(n8), .Y(SUM[14]) );
  AOI21X4 U188 ( .A0(n161), .A1(n160), .B0(n149), .Y(n159) );
  OR2X4 U189 ( .A(A[14]), .B(B[14]), .Y(n114) );
  OR2X4 U190 ( .A(B[12]), .B(A[12]), .Y(n122) );
  NAND2X4 U191 ( .A(A[12]), .B(B[12]), .Y(n120) );
  OAI21X4 U192 ( .A0(n109), .A1(n166), .B0(n167), .Y(n161) );
  NOR2X4 U193 ( .A(n143), .B(n168), .Y(n167) );
  AOI21X4 U194 ( .A0(n14), .A1(n3), .B0(n126), .Y(n174) );
  OR2X4 U195 ( .A(B[11]), .B(A[11]), .Y(n121) );
  OR2X4 U196 ( .A(B[10]), .B(A[10]), .Y(n170) );
  OR2X4 U197 ( .A(B[6]), .B(A[6]), .Y(n74) );
  OR2X4 U198 ( .A(B[7]), .B(A[7]), .Y(n65) );
  NAND2BX4 U199 ( .AN(n110), .B(n21), .Y(n67) );
  OR2X4 U200 ( .A(A[1]), .B(B[1]), .Y(n98) );
  OR2X4 U201 ( .A(A[2]), .B(B[2]), .Y(n97) );
  OR2X4 U202 ( .A(B[9]), .B(A[9]), .Y(n60) );
endmodule


module butterfly_DW01_sub_115 ( A, B, DIFF );
  input [16:0] A;
  input [16:0] B;
  output [16:0] DIFF;
  wire   n251, n252, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n18, n19, n20, n21, n22, n24, n25, n26, n28, n29, n30,
         n31, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250;

  BUFX8 U3 ( .A(n69), .Y(n29) );
  INVX4 U4 ( .A(A[6]), .Y(n16) );
  INVX8 U5 ( .A(n90), .Y(n139) );
  NAND2BX4 U6 ( .AN(A[7]), .B(B[7]), .Y(n106) );
  NAND2BX4 U7 ( .AN(A[7]), .B(B[7]), .Y(n247) );
  INVX8 U8 ( .A(B[7]), .Y(n9) );
  NOR2BX4 U9 ( .AN(n53), .B(n52), .Y(n121) );
  NAND2BX4 U10 ( .AN(n53), .B(n52), .Y(n132) );
  NOR2X4 U11 ( .A(n249), .B(n250), .Y(n246) );
  NOR2BX4 U12 ( .AN(n52), .B(n53), .Y(n116) );
  NAND2BX4 U13 ( .AN(B[1]), .B(A[1]), .Y(n145) );
  INVX8 U14 ( .A(B[1]), .Y(n240) );
  NAND3X4 U15 ( .A(n74), .B(n72), .C(n18), .Y(n77) );
  INVX1 U16 ( .A(n85), .Y(n26) );
  OAI2BB1X4 U17 ( .A0N(n76), .A1N(n77), .B0(n78), .Y(n75) );
  NAND4X1 U18 ( .A(n170), .B(n166), .C(n183), .D(n168), .Y(n160) );
  INVX4 U19 ( .A(n183), .Y(n195) );
  AND2X1 U20 ( .A(n183), .B(n199), .Y(n39) );
  OAI22X4 U21 ( .A0(n241), .A1(n52), .B0(n98), .B1(n99), .Y(n237) );
  INVX8 U22 ( .A(n99), .Y(n31) );
  AOI21X4 U23 ( .A0(n207), .A1(n174), .B0(n208), .Y(n206) );
  INVX4 U24 ( .A(n173), .Y(n208) );
  NAND3BX4 U25 ( .AN(n194), .B(n24), .C(n231), .Y(n235) );
  NAND4BX4 U26 ( .AN(n246), .B(n218), .C(n248), .D(n247), .Y(n194) );
  INVX8 U27 ( .A(n68), .Y(n85) );
  NAND2BX2 U28 ( .AN(B[14]), .B(A[14]), .Y(n165) );
  NAND2BX4 U29 ( .AN(A[14]), .B(B[14]), .Y(n166) );
  NAND2X4 U30 ( .A(n215), .B(n216), .Y(n214) );
  NAND2BX4 U31 ( .AN(B[10]), .B(A[10]), .Y(n216) );
  NOR2X2 U32 ( .A(n84), .B(n139), .Y(n138) );
  NAND2X2 U33 ( .A(n156), .B(n170), .Y(n185) );
  NAND3X2 U34 ( .A(n187), .B(n186), .C(n165), .Y(n184) );
  CLKINVX3 U35 ( .A(n145), .Y(n148) );
  INVX2 U36 ( .A(n60), .Y(n213) );
  CLKINVX3 U37 ( .A(n199), .Y(n167) );
  INVX1 U38 ( .A(n200), .Y(n169) );
  NAND2BX2 U39 ( .AN(B[11]), .B(A[11]), .Y(n215) );
  CLKINVX3 U40 ( .A(n83), .Y(n89) );
  BUFX16 U41 ( .A(n67), .Y(n50) );
  INVX4 U42 ( .A(n230), .Y(n56) );
  INVX2 U43 ( .A(n231), .Y(n57) );
  NAND2BX2 U44 ( .AN(A[15]), .B(B[15]), .Y(n170) );
  NOR2XL U45 ( .A(n142), .B(n102), .Y(n180) );
  OAI21X2 U46 ( .A0(n82), .A1(n83), .B0(n50), .Y(n81) );
  NOR2X2 U47 ( .A(n84), .B(n85), .Y(n82) );
  BUFX16 U48 ( .A(n66), .Y(n51) );
  CLKINVX8 U49 ( .A(n19), .Y(n217) );
  XNOR2X4 U50 ( .A(n224), .B(n41), .Y(n1) );
  XNOR2X4 U51 ( .A(n206), .B(n39), .Y(n2) );
  XNOR2X4 U52 ( .A(n188), .B(n201), .Y(n3) );
  AND2X1 U53 ( .A(n24), .B(n60), .Y(n4) );
  NAND2X1 U54 ( .A(n15), .B(n216), .Y(n5) );
  OAI21X4 U55 ( .A0(n227), .A1(n22), .B0(n228), .Y(n226) );
  NAND4BX4 U56 ( .AN(n245), .B(n12), .C(n247), .D(n91), .Y(n6) );
  NAND4BX2 U57 ( .AN(n245), .B(n12), .C(n106), .D(n91), .Y(n71) );
  NOR2BX4 U58 ( .AN(B[6]), .B(A[6]), .Y(n245) );
  CLKINVX4 U59 ( .A(n76), .Y(n25) );
  NAND3BX2 U60 ( .AN(n121), .B(n100), .C(n122), .Y(n117) );
  XOR2X4 U61 ( .A(n7), .B(n5), .Y(n38) );
  NAND3X4 U62 ( .A(n235), .B(n236), .C(n234), .Y(n7) );
  NOR2BX4 U63 ( .AN(n52), .B(n53), .Y(n97) );
  NAND4X4 U64 ( .A(n120), .B(n50), .C(B[5]), .D(n51), .Y(n218) );
  NAND2X4 U65 ( .A(n9), .B(A[7]), .Y(n66) );
  AOI2BB1X4 U66 ( .A0N(A[0]), .A1N(n8), .B0(n115), .Y(n112) );
  INVX1 U67 ( .A(B[0]), .Y(n8) );
  AOI2BB2X4 U68 ( .B0(A[7]), .B1(n9), .A0N(n16), .A1N(B[6]), .Y(n10) );
  INVX8 U69 ( .A(n10), .Y(n250) );
  AOI21X2 U70 ( .A0(n243), .A1(n101), .B0(n102), .Y(n86) );
  AOI21X1 U71 ( .A0(n168), .A1(n167), .B0(n169), .Y(n11) );
  NAND2BX2 U72 ( .AN(A[13]), .B(B[13]), .Y(n168) );
  NAND2BX1 U73 ( .AN(B[12]), .B(A[12]), .Y(n199) );
  NAND2BX1 U74 ( .AN(B[13]), .B(A[13]), .Y(n200) );
  OAI21XL U75 ( .A0(n43), .A1(n177), .B0(n178), .Y(n176) );
  NAND3X2 U76 ( .A(n219), .B(n61), .C(n62), .Y(n59) );
  INVXL U77 ( .A(n106), .Y(n222) );
  NOR2X2 U78 ( .A(n221), .B(n63), .Y(n62) );
  AOI2BB1X4 U79 ( .A0N(n99), .A1N(n98), .B0(n124), .Y(n122) );
  NAND2X4 U80 ( .A(n28), .B(n73), .Y(n30) );
  CLKINVX8 U81 ( .A(n96), .Y(n28) );
  INVXL U82 ( .A(n31), .Y(n21) );
  CLKINVX4 U83 ( .A(n161), .Y(n174) );
  NAND2X4 U84 ( .A(n19), .B(n203), .Y(n193) );
  BUFX16 U85 ( .A(n137), .Y(n19) );
  NAND4BX1 U86 ( .AN(n195), .B(n196), .C(n168), .D(n197), .Y(n190) );
  AND2X4 U87 ( .A(n118), .B(n14), .Y(n243) );
  NAND2X4 U88 ( .A(n104), .B(n53), .Y(n144) );
  OAI21X2 U89 ( .A0(n99), .A1(B[1]), .B0(n100), .Y(n238) );
  NAND2X4 U90 ( .A(n131), .B(n18), .Y(n130) );
  NAND4X4 U91 ( .A(n76), .B(n19), .C(n24), .D(n231), .Y(n236) );
  NAND4X4 U92 ( .A(n11), .B(n190), .C(n191), .D(n192), .Y(n189) );
  CLKINVX8 U93 ( .A(n71), .Y(n76) );
  INVX8 U94 ( .A(n52), .Y(n104) );
  AOI2BB1X4 U95 ( .A0N(n53), .A1N(n104), .B0(n115), .Y(n119) );
  NAND3X4 U96 ( .A(n16), .B(B[6]), .C(n51), .Y(n248) );
  NAND2BX4 U97 ( .AN(A[1]), .B(B[1]), .Y(n14) );
  OAI2BB1X4 U98 ( .A0N(n241), .A1N(n52), .B0(n28), .Y(n135) );
  CLKINVX8 U99 ( .A(n139), .Y(n12) );
  AOI21X4 U100 ( .A0(n56), .A1(n15), .B0(n214), .Y(n209) );
  NAND3X4 U101 ( .A(n15), .B(n24), .C(n231), .Y(n227) );
  NAND2BX4 U102 ( .AN(A[10]), .B(B[10]), .Y(n15) );
  NAND3X2 U103 ( .A(n211), .B(n213), .C(n212), .Y(n210) );
  NAND2X2 U104 ( .A(n229), .B(n15), .Y(n228) );
  INVXL U105 ( .A(n174), .Y(n13) );
  INVX8 U106 ( .A(n22), .Y(n205) );
  AOI2BB1X4 U107 ( .A0N(n104), .A1N(n53), .B0(n96), .Y(n239) );
  NAND4X2 U108 ( .A(n205), .B(n168), .C(n174), .D(n183), .Y(n191) );
  AOI21X4 U109 ( .A0(n241), .A1(n52), .B0(n105), .Y(n242) );
  INVX8 U110 ( .A(n53), .Y(n241) );
  NOR2BX1 U111 ( .AN(B[9]), .B(A[9]), .Y(n223) );
  NAND2X4 U112 ( .A(n204), .B(n205), .Y(n202) );
  NOR2X2 U113 ( .A(n195), .B(n161), .Y(n204) );
  BUFX20 U114 ( .A(n2), .Y(DIFF[12]) );
  CLKINVX3 U115 ( .A(n102), .Y(n18) );
  AOI21X2 U116 ( .A0(n241), .A1(n52), .B0(n105), .Y(n101) );
  CLKINVX1 U117 ( .A(n56), .Y(n20) );
  OAI21X4 U118 ( .A0(n217), .A1(n232), .B0(n216), .Y(n225) );
  INVX8 U119 ( .A(A[1]), .Y(n99) );
  OAI21X4 U120 ( .A0(n217), .A1(n25), .B0(n78), .Y(n207) );
  NAND2BX4 U121 ( .AN(n193), .B(n168), .Y(n192) );
  NOR3X4 U122 ( .A(n161), .B(n195), .C(n6), .Y(n203) );
  NAND4BX4 U123 ( .AN(n246), .B(n218), .C(n248), .D(n247), .Y(n22) );
  BUFX20 U124 ( .A(n1), .Y(DIFF[11]) );
  OAI2BB1X4 U125 ( .A0N(n146), .A1N(n14), .B0(n145), .Y(n141) );
  BUFX20 U126 ( .A(n64), .Y(n24) );
  NOR2X4 U127 ( .A(n96), .B(n103), .Y(n133) );
  NOR3X4 U128 ( .A(n94), .B(n136), .C(n121), .Y(n134) );
  NOR2X4 U129 ( .A(n148), .B(n103), .Y(n147) );
  AOI2BB1X4 U130 ( .A0N(n102), .A1N(n84), .B0(n115), .Y(n114) );
  INVX8 U131 ( .A(n3), .Y(DIFF[13]) );
  OAI21X2 U132 ( .A0(n57), .A1(n60), .B0(n20), .Y(n229) );
  NOR2XL U133 ( .A(n160), .B(n13), .Y(n158) );
  NAND3X2 U134 ( .A(n117), .B(n28), .C(n119), .Y(n110) );
  OAI2BB1X4 U135 ( .A0N(n52), .A1N(n241), .B0(n144), .Y(n143) );
  NAND3X1 U136 ( .A(n166), .B(n168), .C(n188), .Y(n187) );
  NAND2X2 U137 ( .A(n89), .B(n12), .Y(n88) );
  NOR2X4 U138 ( .A(n226), .B(n225), .Y(n224) );
  NAND2X4 U139 ( .A(n29), .B(n68), .Y(n249) );
  NAND2BX1 U140 ( .AN(A[9]), .B(B[9]), .Y(n211) );
  NAND2BX2 U141 ( .AN(B[9]), .B(A[9]), .Y(n230) );
  NOR2X4 U142 ( .A(n134), .B(n135), .Y(n129) );
  INVX2 U143 ( .A(n100), .Y(n136) );
  NAND2BX4 U144 ( .AN(n6), .B(n24), .Y(n70) );
  NAND4BX4 U145 ( .AN(n167), .B(n193), .C(n202), .D(n35), .Y(n188) );
  NAND4X2 U146 ( .A(n68), .B(n50), .C(n51), .D(n29), .Y(n219) );
  INVX4 U147 ( .A(A[5]), .Y(n120) );
  INVX4 U148 ( .A(n65), .Y(n221) );
  AOI21X2 U149 ( .A0(n213), .A1(n231), .B0(n56), .Y(n234) );
  INVX8 U150 ( .A(n69), .Y(n84) );
  OAI22X4 U151 ( .A0(n98), .A1(n99), .B0(n99), .B1(B[1]), .Y(n94) );
  NAND3X4 U152 ( .A(n220), .B(n219), .C(n218), .Y(n78) );
  NOR2X4 U153 ( .A(n221), .B(n222), .Y(n220) );
  AND2X4 U154 ( .A(n31), .B(n240), .Y(n124) );
  OAI21X4 U155 ( .A0(n130), .A1(n129), .B0(n12), .Y(n128) );
  XOR2X4 U156 ( .A(n140), .B(n30), .Y(n36) );
  INVXL U157 ( .A(n92), .Y(n109) );
  AND2X1 U158 ( .A(n165), .B(n166), .Y(n37) );
  NAND2X4 U159 ( .A(n128), .B(n29), .Y(n125) );
  NAND2X4 U160 ( .A(n209), .B(n210), .Y(n197) );
  BUFX20 U161 ( .A(n252), .Y(DIFF[2]) );
  NOR2X2 U162 ( .A(n96), .B(n97), .Y(n95) );
  AOI21X4 U163 ( .A0(n112), .A1(n113), .B0(n114), .Y(n111) );
  NAND3X2 U164 ( .A(n196), .B(n183), .C(n197), .Y(n35) );
  INVX8 U165 ( .A(n73), .Y(n102) );
  AND2X1 U166 ( .A(n26), .B(n29), .Y(n43) );
  NOR3X2 U167 ( .A(n96), .B(n116), .C(n103), .Y(n113) );
  NAND2X2 U168 ( .A(n247), .B(n24), .Y(n63) );
  CLKINVX3 U169 ( .A(n227), .Y(n233) );
  AOI21XL U170 ( .A0(n180), .A1(n181), .B0(n25), .Y(n175) );
  XNOR2X4 U171 ( .A(n141), .B(n143), .Y(n252) );
  INVX20 U172 ( .A(n44), .Y(DIFF[6]) );
  BUFX20 U173 ( .A(n36), .Y(DIFF[3]) );
  AOI21X2 U174 ( .A0(n152), .A1(n153), .B0(n154), .Y(n150) );
  OAI21X2 U175 ( .A0(n52), .A1(n241), .B0(n100), .Y(n93) );
  NAND3BX2 U176 ( .AN(A[6]), .B(B[6]), .C(n51), .Y(n65) );
  INVX8 U177 ( .A(n47), .Y(DIFF[1]) );
  XNOR2X4 U178 ( .A(n146), .B(n147), .Y(n47) );
  NAND2BX4 U179 ( .AN(A[8]), .B(B[8]), .Y(n64) );
  NAND2X2 U180 ( .A(n196), .B(n197), .Y(n173) );
  NAND2X2 U181 ( .A(n76), .B(n233), .Y(n232) );
  NAND2BX4 U182 ( .AN(A[9]), .B(B[9]), .Y(n231) );
  BUFX20 U183 ( .A(n251), .Y(DIFF[4]) );
  INVX4 U184 ( .A(n168), .Y(n198) );
  INVX4 U185 ( .A(n144), .Y(n142) );
  NAND2X4 U186 ( .A(n123), .B(n240), .Y(n100) );
  INVX8 U187 ( .A(n38), .Y(DIFF[10]) );
  XOR2X4 U188 ( .A(n19), .B(n138), .Y(n251) );
  NAND2BX4 U189 ( .AN(B[5]), .B(A[5]), .Y(n68) );
  OAI2BB1X4 U190 ( .A0N(n120), .A1N(B[5]), .B0(n90), .Y(n115) );
  AND3X4 U191 ( .A(n111), .B(n110), .C(n26), .Y(n45) );
  NAND2BX4 U192 ( .AN(B[8]), .B(A[8]), .Y(n60) );
  NAND2X4 U193 ( .A(n91), .B(n92), .Y(n83) );
  INVX8 U194 ( .A(n42), .Y(DIFF[5]) );
  NAND2BX4 U195 ( .AN(A[6]), .B(B[6]), .Y(n92) );
  NAND3X1 U196 ( .A(n155), .B(n156), .C(n157), .Y(n154) );
  XOR2X4 U197 ( .A(n34), .B(n79), .Y(DIFF[7]) );
  NAND2XL U198 ( .A(n106), .B(n51), .Y(n34) );
  INVXL U199 ( .A(n50), .Y(n108) );
  INVXL U200 ( .A(n160), .Y(n152) );
  AND2X1 U201 ( .A(n50), .B(n51), .Y(n178) );
  NAND2BX4 U202 ( .AN(B[4]), .B(A[4]), .Y(n69) );
  INVX8 U203 ( .A(n46), .Y(DIFF[15]) );
  OAI21XL U204 ( .A0(n163), .A1(n164), .B0(n165), .Y(n162) );
  INVXL U205 ( .A(n166), .Y(n164) );
  NAND2XL U206 ( .A(n170), .B(n162), .Y(n155) );
  XNOR2X4 U207 ( .A(n54), .B(n55), .Y(n40) );
  INVX8 U208 ( .A(n40), .Y(DIFF[9]) );
  INVXL U209 ( .A(n91), .Y(n127) );
  AND2X1 U210 ( .A(n196), .B(n215), .Y(n41) );
  XNOR2X4 U211 ( .A(n125), .B(n126), .Y(n42) );
  INVXL U212 ( .A(n72), .Y(n159) );
  XOR2X4 U213 ( .A(n45), .B(n107), .Y(n44) );
  XOR2X4 U214 ( .A(n184), .B(n185), .Y(n46) );
  OAI21XL U215 ( .A0(n179), .A1(A[5]), .B0(n92), .Y(n177) );
  INVXL U216 ( .A(B[5]), .Y(n179) );
  OAI21XL U217 ( .A0(n171), .A1(n172), .B0(n173), .Y(n153) );
  NAND2XL U218 ( .A(n174), .B(n106), .Y(n172) );
  AOI21XL U219 ( .A0(n175), .A1(n28), .B0(n176), .Y(n171) );
  AOI21XL U220 ( .A0(n167), .A1(n168), .B0(n169), .Y(n163) );
  NAND2XL U221 ( .A(n169), .B(n166), .Y(n186) );
  BUFX20 U222 ( .A(A[2]), .Y(n53) );
  XOR2X1 U223 ( .A(B[16]), .B(A[16]), .Y(n151) );
  OAI21XL U224 ( .A0(n148), .A1(n182), .B0(n132), .Y(n181) );
  NAND2BX1 U225 ( .AN(B[15]), .B(A[15]), .Y(n156) );
  NAND2X1 U226 ( .A(n98), .B(n149), .Y(DIFF[0]) );
  INVX1 U227 ( .A(n149), .Y(n105) );
  INVX1 U228 ( .A(n98), .Y(n123) );
  NAND2BX1 U229 ( .AN(n149), .B(n98), .Y(n146) );
  NAND2BX1 U230 ( .AN(B[0]), .B(A[0]), .Y(n98) );
  NAND2BX1 U231 ( .AN(A[0]), .B(B[0]), .Y(n149) );
  NOR2BX4 U232 ( .AN(n77), .B(n70), .Y(n58) );
  NAND4BXL U233 ( .AN(A[5]), .B(n50), .C(n51), .D(B[5]), .Y(n61) );
  BUFX20 U234 ( .A(B[2]), .Y(n52) );
  OAI21X2 U235 ( .A0(n93), .A1(n94), .B0(n95), .Y(n87) );
  NAND3XL U236 ( .A(n76), .B(n158), .C(n159), .Y(n157) );
  INVX8 U237 ( .A(n244), .Y(n103) );
  NAND2BX4 U238 ( .AN(A[1]), .B(B[1]), .Y(n244) );
  INVX8 U239 ( .A(n118), .Y(n96) );
  OAI21XL U240 ( .A0(n98), .A1(n21), .B0(n100), .Y(n182) );
  NOR2X4 U241 ( .A(n56), .B(n57), .Y(n55) );
  NAND3BX4 U242 ( .AN(n58), .B(n59), .C(n60), .Y(n54) );
  XOR2X4 U243 ( .A(n75), .B(n4), .Y(DIFF[8]) );
  NOR2X4 U244 ( .A(n80), .B(n81), .Y(n79) );
  AOI21X4 U245 ( .A0(n87), .A1(n86), .B0(n88), .Y(n80) );
  NOR2X4 U246 ( .A(n108), .B(n109), .Y(n107) );
  NOR2X4 U247 ( .A(n85), .B(n127), .Y(n126) );
  NAND3X4 U248 ( .A(n133), .B(n132), .C(n149), .Y(n131) );
  AOI21X4 U249 ( .A0(n141), .A1(n132), .B0(n142), .Y(n140) );
  XOR2X4 U250 ( .A(n150), .B(n151), .Y(DIFF[16]) );
  XOR2X4 U251 ( .A(n189), .B(n37), .Y(DIFF[14]) );
  NOR2X4 U252 ( .A(n198), .B(n169), .Y(n201) );
  NAND4BX4 U253 ( .AN(n223), .B(n196), .C(n212), .D(n24), .Y(n161) );
  NAND2BX4 U254 ( .AN(A[12]), .B(B[12]), .Y(n183) );
  NAND2BX4 U255 ( .AN(A[11]), .B(B[11]), .Y(n196) );
  NAND2BX4 U256 ( .AN(A[10]), .B(B[10]), .Y(n212) );
  NAND3BX4 U257 ( .AN(n102), .B(n74), .C(n72), .Y(n137) );
  OAI21X4 U258 ( .A0(n237), .A1(n238), .B0(n239), .Y(n74) );
  NAND2X4 U259 ( .A(n242), .B(n243), .Y(n72) );
  NAND2BX4 U260 ( .AN(A[3]), .B(B[3]), .Y(n118) );
  NAND2BX4 U261 ( .AN(B[3]), .B(A[3]), .Y(n73) );
  NAND2BX4 U262 ( .AN(A[5]), .B(B[5]), .Y(n91) );
  NAND2BX4 U263 ( .AN(A[4]), .B(B[4]), .Y(n90) );
  NAND2BX4 U264 ( .AN(B[6]), .B(A[6]), .Y(n67) );
endmodule


module butterfly_DW01_add_158 ( A, B, SUM );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  wire   n186, n187, n188, n189, n190, n191, n192, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n29, n30, n31, n33, n34, n35, n36, n37,
         n38, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185;

  INVX8 U2 ( .A(n122), .Y(n120) );
  OAI21X1 U3 ( .A0(n141), .A1(n113), .B0(n17), .Y(n149) );
  NAND2X2 U4 ( .A(B[15]), .B(A[15]), .Y(n111) );
  AOI2BB1X4 U5 ( .A0N(n109), .A1N(n110), .B0(n2), .Y(n1) );
  CLKINVX20 U6 ( .A(n111), .Y(n2) );
  NAND2X1 U7 ( .A(B[1]), .B(A[1]), .Y(n101) );
  CLKINVX3 U8 ( .A(n141), .Y(n139) );
  NAND2X4 U9 ( .A(A[12]), .B(B[12]), .Y(n141) );
  NOR2X4 U10 ( .A(A[13]), .B(B[13]), .Y(n113) );
  NAND2X4 U11 ( .A(n17), .B(n115), .Y(n114) );
  NOR2BX4 U12 ( .AN(n59), .B(n6), .Y(n58) );
  INVX2 U13 ( .A(n6), .Y(n7) );
  CLKINVX2 U14 ( .A(n12), .Y(n6) );
  NAND3BX2 U15 ( .AN(n63), .B(n86), .C(n183), .Y(n5) );
  INVX4 U16 ( .A(n181), .Y(n129) );
  OR2X2 U17 ( .A(A[1]), .B(B[1]), .Y(n99) );
  INVX1 U18 ( .A(n150), .Y(n30) );
  NOR2BX2 U19 ( .AN(n141), .B(n9), .Y(n159) );
  NAND2X1 U20 ( .A(B[0]), .B(A[0]), .Y(n104) );
  INVX2 U21 ( .A(n99), .Y(n103) );
  BUFX3 U22 ( .A(n191), .Y(SUM[5]) );
  NOR2BX1 U23 ( .AN(n79), .B(n78), .Y(n81) );
  XOR2X2 U24 ( .A(n89), .B(n90), .Y(SUM[3]) );
  INVX4 U25 ( .A(n10), .Y(SUM[4]) );
  BUFX8 U26 ( .A(n189), .Y(SUM[8]) );
  XOR2X2 U27 ( .A(n60), .B(n61), .Y(n189) );
  NOR2BX1 U28 ( .AN(n62), .B(n63), .Y(n61) );
  OAI21X4 U29 ( .A0(n142), .A1(n17), .B0(n115), .Y(n140) );
  CLKINVX3 U30 ( .A(n118), .Y(n183) );
  OR2X4 U31 ( .A(n152), .B(n153), .Y(n3) );
  AND2X4 U32 ( .A(A[13]), .B(B[13]), .Y(n4) );
  NAND4X4 U33 ( .A(n51), .B(n21), .C(n19), .D(n137), .Y(n136) );
  AND2X4 U34 ( .A(n21), .B(n65), .Y(n15) );
  INVX8 U35 ( .A(n86), .Y(n84) );
  NAND4X4 U36 ( .A(n127), .B(n181), .C(n18), .D(n69), .Y(n64) );
  INVX2 U37 ( .A(A[9]), .Y(n13) );
  NAND2X1 U38 ( .A(n30), .B(n22), .Y(n160) );
  NAND3BX4 U39 ( .AN(n13), .B(n36), .C(n38), .Y(n163) );
  BUFX20 U40 ( .A(n186), .Y(SUM[12]) );
  OAI21X4 U41 ( .A0(n146), .A1(n145), .B0(n147), .Y(n143) );
  AND2X2 U42 ( .A(n127), .B(n128), .Y(n50) );
  NOR2X1 U43 ( .A(n129), .B(n130), .Y(n128) );
  OR2X4 U44 ( .A(A[9]), .B(B[9]), .Y(n165) );
  INVX2 U45 ( .A(B[9]), .Y(n35) );
  NAND2X2 U46 ( .A(B[9]), .B(A[9]), .Y(n59) );
  NAND3X2 U47 ( .A(n175), .B(n176), .C(n62), .Y(n8) );
  CLKINVX4 U48 ( .A(n35), .Y(n36) );
  BUFX4 U49 ( .A(n121), .Y(n37) );
  NOR2X4 U50 ( .A(A[12]), .B(B[12]), .Y(n9) );
  INVX2 U51 ( .A(n142), .Y(n29) );
  XOR2X1 U52 ( .A(n84), .B(n87), .Y(n10) );
  NAND2XL U53 ( .A(n115), .B(n112), .Y(n144) );
  NAND2X2 U54 ( .A(B[8]), .B(A[8]), .Y(n62) );
  OAI2BB1X2 U55 ( .A0N(n65), .A1N(n64), .B0(n66), .Y(n60) );
  INVX4 U56 ( .A(n66), .Y(n152) );
  NAND2X4 U57 ( .A(n54), .B(n119), .Y(n108) );
  NAND2X2 U58 ( .A(n166), .B(n167), .Y(n161) );
  NAND2XL U59 ( .A(A[8]), .B(B[8]), .Y(n27) );
  AND3X4 U60 ( .A(n20), .B(n19), .C(n65), .Y(n11) );
  NAND2X1 U61 ( .A(n124), .B(n112), .Y(n110) );
  CLKINVX8 U62 ( .A(n23), .Y(n12) );
  NOR2X4 U63 ( .A(B[9]), .B(A[9]), .Y(n23) );
  AND3X4 U64 ( .A(n175), .B(n176), .C(n45), .Y(n173) );
  NAND4X4 U65 ( .A(n24), .B(n29), .C(n19), .D(n22), .Y(n134) );
  OAI21X4 U66 ( .A0(n71), .A1(n72), .B0(n18), .Y(n67) );
  INVX4 U67 ( .A(n112), .Y(n142) );
  NAND4BBX2 U68 ( .AN(n70), .BN(n113), .C(n20), .D(n19), .Y(n146) );
  NAND3BX4 U69 ( .AN(n161), .B(n162), .C(n163), .Y(n22) );
  OR2X4 U70 ( .A(B[6]), .B(A[6]), .Y(n14) );
  INVX4 U71 ( .A(n172), .Y(n34) );
  NAND2BX2 U72 ( .AN(n56), .B(A[6]), .Y(n73) );
  INVX2 U73 ( .A(B[6]), .Y(n56) );
  INVX8 U74 ( .A(n125), .Y(n124) );
  AOI21X4 U75 ( .A0(n138), .A1(n139), .B0(n140), .Y(n135) );
  NOR2BX2 U76 ( .AN(n18), .B(n72), .Y(n75) );
  OAI2BB1X4 U77 ( .A0N(n15), .A1N(n3), .B0(n160), .Y(n158) );
  NAND3X4 U78 ( .A(n135), .B(n134), .C(n136), .Y(n132) );
  CLKBUFX2 U79 ( .A(n166), .Y(n16) );
  INVX8 U80 ( .A(n4), .Y(n17) );
  INVX3 U81 ( .A(n82), .Y(n78) );
  NAND2BX4 U82 ( .AN(n56), .B(A[6]), .Y(n18) );
  INVX1 U83 ( .A(n65), .Y(n70) );
  NAND4BX2 U84 ( .AN(n129), .B(n127), .C(n69), .D(n18), .Y(n153) );
  AOI21X4 U85 ( .A0(n119), .A1(n157), .B0(n139), .Y(n156) );
  AOI21X4 U86 ( .A0(n119), .A1(n148), .B0(n149), .Y(n147) );
  INVX8 U87 ( .A(n9), .Y(n19) );
  NOR2X4 U88 ( .A(n169), .B(n168), .Y(n20) );
  NOR2X4 U89 ( .A(n169), .B(n168), .Y(n21) );
  AND2X2 U90 ( .A(n117), .B(n37), .Y(n24) );
  INVX4 U91 ( .A(n80), .Y(n77) );
  NAND2X4 U92 ( .A(n3), .B(n11), .Y(n25) );
  NAND2X4 U93 ( .A(n25), .B(n156), .Y(n154) );
  NOR2X2 U94 ( .A(n152), .B(n153), .Y(n145) );
  AND2X4 U95 ( .A(B[4]), .B(A[4]), .Y(n180) );
  OAI22X2 U96 ( .A0(B[13]), .A1(A[13]), .B0(B[14]), .B1(A[14]), .Y(n123) );
  INVX12 U97 ( .A(n121), .Y(n150) );
  XNOR2X4 U98 ( .A(n105), .B(n26), .Y(SUM[16]) );
  XNOR2X4 U99 ( .A(B[16]), .B(A[16]), .Y(n26) );
  NAND3BX4 U100 ( .AN(n27), .B(n164), .C(n165), .Y(n162) );
  NOR2X2 U101 ( .A(n142), .B(n113), .Y(n138) );
  NOR2BX2 U102 ( .AN(n167), .B(n150), .Y(n172) );
  XOR2X4 U103 ( .A(n8), .B(n58), .Y(n188) );
  NAND2X2 U104 ( .A(n69), .B(n73), .Y(n130) );
  AOI21X4 U105 ( .A0(n57), .A1(n7), .B0(n179), .Y(n178) );
  NAND2X2 U106 ( .A(A[5]), .B(B[5]), .Y(n182) );
  NAND2X4 U107 ( .A(B[5]), .B(A[5]), .Y(n79) );
  INVX1 U108 ( .A(n59), .Y(n179) );
  NAND2X2 U109 ( .A(n117), .B(n116), .Y(n151) );
  OAI2BB1X2 U110 ( .A0N(n49), .A1N(n50), .B0(n65), .Y(n106) );
  INVX3 U111 ( .A(n170), .Y(n63) );
  AND2X2 U112 ( .A(n59), .B(n62), .Y(n45) );
  NAND3BX4 U113 ( .AN(n63), .B(n86), .C(n183), .Y(n176) );
  NAND2X2 U114 ( .A(B[10]), .B(A[10]), .Y(n166) );
  OR2X4 U115 ( .A(A[4]), .B(B[4]), .Y(n88) );
  NAND2BX4 U116 ( .AN(n64), .B(n66), .Y(n137) );
  AOI21X2 U117 ( .A0(n131), .A1(n91), .B0(n118), .Y(n126) );
  NAND2X2 U118 ( .A(A[11]), .B(B[11]), .Y(n167) );
  BUFX20 U119 ( .A(n190), .Y(SUM[6]) );
  XOR2X4 U120 ( .A(n74), .B(n75), .Y(n190) );
  CLKINVX8 U121 ( .A(n187), .Y(n31) );
  INVX8 U122 ( .A(n31), .Y(SUM[11]) );
  XNOR2X4 U123 ( .A(n158), .B(n33), .Y(n186) );
  CLKINVX20 U124 ( .A(n159), .Y(n33) );
  XNOR2X4 U125 ( .A(n171), .B(n34), .Y(n187) );
  NAND3X4 U126 ( .A(n175), .B(n5), .C(n62), .Y(n57) );
  BUFX20 U127 ( .A(n188), .Y(SUM[9]) );
  NAND2X4 U128 ( .A(n12), .B(n170), .Y(n168) );
  NAND2X4 U129 ( .A(n121), .B(n164), .Y(n169) );
  AND3X4 U130 ( .A(n112), .B(n117), .C(n65), .Y(n51) );
  NAND2X4 U131 ( .A(B[2]), .B(A[2]), .Y(n95) );
  OR2X4 U132 ( .A(A[10]), .B(B[10]), .Y(n38) );
  NAND2BX4 U133 ( .AN(n118), .B(n86), .Y(n66) );
  NOR2X2 U134 ( .A(n150), .B(n9), .Y(n157) );
  OAI21X4 U135 ( .A0(n173), .A1(n174), .B0(n16), .Y(n171) );
  NAND4X4 U136 ( .A(n55), .B(n88), .C(n82), .D(n76), .Y(n118) );
  NAND2X4 U137 ( .A(n64), .B(n52), .Y(n175) );
  XOR2X4 U138 ( .A(n67), .B(n68), .Y(SUM[7]) );
  BUFX3 U139 ( .A(n192), .Y(SUM[0]) );
  AND2X2 U140 ( .A(n170), .B(n65), .Y(n52) );
  NOR2XL U141 ( .A(A[0]), .B(B[0]), .Y(n44) );
  NAND2X4 U142 ( .A(n91), .B(n131), .Y(n86) );
  NAND2X1 U143 ( .A(n111), .B(n124), .Y(n133) );
  INVX4 U144 ( .A(n74), .Y(n71) );
  INVX2 U145 ( .A(n126), .Y(n49) );
  INVXL U146 ( .A(n104), .Y(n100) );
  NOR2BX1 U147 ( .AN(n104), .B(n44), .Y(n192) );
  INVX1 U148 ( .A(n96), .Y(n93) );
  XOR2X4 U149 ( .A(n132), .B(n133), .Y(n46) );
  INVX8 U150 ( .A(n46), .Y(SUM[15]) );
  XOR2X4 U151 ( .A(n143), .B(n144), .Y(n47) );
  INVX8 U152 ( .A(n47), .Y(SUM[14]) );
  XOR2X4 U153 ( .A(n154), .B(n155), .Y(n48) );
  INVX8 U154 ( .A(n48), .Y(SUM[13]) );
  NAND2XL U155 ( .A(n17), .B(n117), .Y(n155) );
  XOR2X1 U156 ( .A(n80), .B(n81), .Y(n191) );
  NOR2BX1 U157 ( .AN(n91), .B(n92), .Y(n90) );
  OAI21XL U158 ( .A0(n93), .A1(n94), .B0(n95), .Y(n89) );
  INVX1 U159 ( .A(n185), .Y(n92) );
  XOR2X1 U160 ( .A(n96), .B(n97), .Y(SUM[2]) );
  NOR2BX1 U161 ( .AN(n95), .B(n94), .Y(n97) );
  XOR2X1 U162 ( .A(n100), .B(n102), .Y(SUM[1]) );
  NOR2BXL U163 ( .AN(n101), .B(n103), .Y(n102) );
  NOR2BXL U164 ( .AN(n85), .B(n83), .Y(n87) );
  OAI2BB1X1 U165 ( .A0N(n99), .A1N(n100), .B0(n101), .Y(n96) );
  NAND2X4 U166 ( .A(n53), .B(n184), .Y(n131) );
  AND2X4 U167 ( .A(n98), .B(n185), .Y(n53) );
  AND2X4 U168 ( .A(n120), .B(n37), .Y(n54) );
  NAND2XL U169 ( .A(B[4]), .B(A[4]), .Y(n85) );
  NAND2X1 U170 ( .A(B[3]), .B(A[3]), .Y(n91) );
  OR2X4 U171 ( .A(A[7]), .B(B[7]), .Y(n55) );
  NAND2X2 U172 ( .A(n120), .B(n21), .Y(n107) );
  NOR2X2 U173 ( .A(n150), .B(n151), .Y(n148) );
  NOR2BX1 U174 ( .AN(n69), .B(n70), .Y(n68) );
  NAND2XL U175 ( .A(n166), .B(n164), .Y(n177) );
  INVXL U176 ( .A(n14), .Y(n72) );
  NAND2XL U177 ( .A(n38), .B(n12), .Y(n174) );
  NAND2X2 U178 ( .A(B[14]), .B(A[14]), .Y(n115) );
  OAI21X4 U179 ( .A0(n77), .A1(n78), .B0(n79), .Y(n74) );
  OAI21X4 U180 ( .A0(n83), .A1(n84), .B0(n85), .Y(n80) );
  CLKINVX3 U181 ( .A(n88), .Y(n83) );
  CLKINVX3 U182 ( .A(n98), .Y(n94) );
  OAI211X2 U183 ( .A0(n107), .A1(n106), .B0(n108), .C0(n1), .Y(n105) );
  AOI2BB1X4 U184 ( .A0N(n113), .A1N(n141), .B0(n114), .Y(n109) );
  NAND3BX4 U185 ( .AN(n123), .B(n116), .C(n124), .Y(n122) );
  NOR2X4 U186 ( .A(B[15]), .B(A[15]), .Y(n125) );
  OR2X4 U187 ( .A(B[14]), .B(A[14]), .Y(n112) );
  OR2X4 U188 ( .A(A[13]), .B(B[13]), .Y(n117) );
  OR2X4 U189 ( .A(A[12]), .B(B[12]), .Y(n116) );
  NAND3BX4 U190 ( .AN(n161), .B(n162), .C(n163), .Y(n119) );
  OR2X4 U191 ( .A(A[11]), .B(B[11]), .Y(n121) );
  XOR2X4 U192 ( .A(n178), .B(n177), .Y(SUM[10]) );
  NAND3X4 U193 ( .A(n82), .B(n76), .C(n180), .Y(n127) );
  NAND2X4 U194 ( .A(B[7]), .B(A[7]), .Y(n69) );
  NAND2BX4 U195 ( .AN(n182), .B(n14), .Y(n181) );
  OR2X4 U196 ( .A(A[7]), .B(B[7]), .Y(n65) );
  OR2X4 U197 ( .A(B[6]), .B(A[6]), .Y(n76) );
  OR2X4 U198 ( .A(B[5]), .B(A[5]), .Y(n82) );
  OAI211X2 U199 ( .A0(n103), .A1(n104), .B0(n101), .C0(n95), .Y(n184) );
  OR2X4 U200 ( .A(A[2]), .B(B[2]), .Y(n98) );
  OR2X4 U201 ( .A(A[3]), .B(B[3]), .Y(n185) );
  OR2X4 U202 ( .A(B[8]), .B(A[8]), .Y(n170) );
  OR2X4 U203 ( .A(B[10]), .B(A[10]), .Y(n164) );
endmodule


module butterfly_DW01_sub_118 ( A, B, DIFF );
  input [16:0] A;
  input [16:0] B;
  output [16:0] DIFF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216;

  NAND2BX4 U3 ( .AN(A[3]), .B(B[3]), .Y(n194) );
  NAND2BX4 U4 ( .AN(A[12]), .B(n30), .Y(n152) );
  NAND2BX4 U5 ( .AN(A[12]), .B(n30), .Y(n20) );
  CLKINVX3 U6 ( .A(n146), .Y(n142) );
  NAND2X4 U7 ( .A(n94), .B(n95), .Y(n93) );
  NOR2X4 U8 ( .A(n74), .B(n81), .Y(n210) );
  INVX4 U9 ( .A(n216), .Y(n81) );
  INVX8 U10 ( .A(n47), .Y(n31) );
  NOR2BX2 U11 ( .AN(B[9]), .B(A[9]), .Y(n173) );
  OAI21X4 U12 ( .A0(n52), .A1(n56), .B0(n53), .Y(n185) );
  INVX4 U13 ( .A(n32), .Y(n56) );
  INVX2 U14 ( .A(n113), .Y(n10) );
  NAND2X2 U15 ( .A(n43), .B(n68), .Y(n198) );
  NAND2BX4 U16 ( .AN(A[1]), .B(B[1]), .Y(n216) );
  XOR2X4 U17 ( .A(n114), .B(n115), .Y(DIFF[1]) );
  INVX3 U18 ( .A(A[4]), .Y(n16) );
  XOR2X4 U19 ( .A(n109), .B(n111), .Y(DIFF[2]) );
  INVX1 U20 ( .A(n25), .Y(n8) );
  AND2X2 U21 ( .A(n179), .B(n84), .Y(n43) );
  INVX4 U22 ( .A(n29), .Y(n30) );
  NOR2X1 U23 ( .A(n80), .B(n81), .Y(n75) );
  NAND2BX2 U24 ( .AN(A[3]), .B(B[3]), .Y(n72) );
  NAND2X2 U25 ( .A(n202), .B(n203), .Y(n201) );
  INVX4 U26 ( .A(n184), .Y(n175) );
  INVX4 U27 ( .A(n150), .Y(n130) );
  NAND2X1 U28 ( .A(n185), .B(n170), .Y(n183) );
  INVX4 U29 ( .A(n136), .Y(n124) );
  NAND2X1 U30 ( .A(n134), .B(n159), .Y(n158) );
  NAND2X1 U31 ( .A(n130), .B(n21), .Y(n159) );
  NAND2BX2 U32 ( .AN(A[15]), .B(B[15]), .Y(n129) );
  NAND2BX1 U33 ( .AN(B[15]), .B(A[15]), .Y(n127) );
  NOR2X1 U34 ( .A(n54), .B(n32), .Y(n83) );
  NOR2X1 U35 ( .A(n136), .B(n168), .Y(n162) );
  NOR2BX1 U36 ( .AN(n53), .B(n52), .Y(n51) );
  NAND2BX1 U37 ( .AN(B[0]), .B(A[0]), .Y(n116) );
  NOR2X2 U38 ( .A(n110), .B(n74), .Y(n111) );
  NAND2X1 U39 ( .A(n72), .B(n78), .Y(n107) );
  AND2X2 U40 ( .A(n190), .B(n87), .Y(n1) );
  AND2X4 U41 ( .A(n89), .B(n205), .Y(n2) );
  AND2X4 U42 ( .A(n165), .B(n166), .Y(n3) );
  NOR2X2 U43 ( .A(n196), .B(n175), .Y(n4) );
  INVX1 U44 ( .A(A[9]), .Y(n14) );
  XNOR2X4 U45 ( .A(n5), .B(n98), .Y(DIFF[6]) );
  OR2X2 U46 ( .A(n19), .B(n64), .Y(n5) );
  AOI21X4 U47 ( .A0(n92), .A1(n104), .B0(n105), .Y(n103) );
  AND2X2 U48 ( .A(n127), .B(n129), .Y(n41) );
  AND2X4 U49 ( .A(n142), .B(n129), .Y(n42) );
  NAND2BX1 U50 ( .AN(A[5]), .B(n48), .Y(n6) );
  NAND2BX2 U51 ( .AN(A[5]), .B(n48), .Y(n205) );
  NAND2BX2 U52 ( .AN(A[6]), .B(B[6]), .Y(n89) );
  NAND2X2 U53 ( .A(n92), .B(n89), .Y(n192) );
  INVX8 U54 ( .A(n92), .Y(n67) );
  AND3X4 U55 ( .A(n89), .B(n91), .C(n92), .Y(n35) );
  AND3X2 U56 ( .A(n73), .B(n76), .C(n213), .Y(n7) );
  NOR2X2 U57 ( .A(n7), .B(n214), .Y(n206) );
  NOR2X2 U58 ( .A(n81), .B(n215), .Y(n213) );
  NOR2BX1 U59 ( .AN(n194), .B(n79), .Y(n214) );
  NAND2XL U60 ( .A(n210), .B(n73), .Y(n70) );
  AND2X4 U61 ( .A(n11), .B(n216), .Y(n115) );
  NAND2X4 U62 ( .A(n164), .B(n150), .Y(n163) );
  AND2X1 U63 ( .A(n97), .B(n78), .Y(n17) );
  NAND2X2 U64 ( .A(n2), .B(n204), .Y(n202) );
  AOI21X2 U65 ( .A0(n76), .A1(n109), .B0(n110), .Y(n108) );
  XOR2X4 U66 ( .A(n169), .B(n8), .Y(DIFF[12]) );
  OAI21X1 U67 ( .A0(n125), .A1(n126), .B0(n127), .Y(n122) );
  OR2X4 U68 ( .A(B[9]), .B(n14), .Y(n53) );
  OR2X4 U69 ( .A(B[4]), .B(n16), .Y(n9) );
  CLKINVX8 U70 ( .A(n10), .Y(n11) );
  INVX8 U71 ( .A(n37), .Y(n26) );
  AND2X4 U72 ( .A(n206), .B(n207), .Y(n28) );
  AOI21X2 U73 ( .A0(n209), .A1(n210), .B0(n211), .Y(n207) );
  INVX1 U74 ( .A(n185), .Y(n199) );
  NAND2X4 U75 ( .A(n14), .B(B[9]), .Y(n179) );
  BUFX8 U76 ( .A(n61), .Y(n15) );
  NAND2BX4 U77 ( .AN(B[10]), .B(A[10]), .Y(n184) );
  NAND3BX4 U78 ( .AN(n60), .B(n15), .C(n62), .Y(n59) );
  BUFX16 U79 ( .A(B[5]), .Y(n48) );
  INVX8 U80 ( .A(n82), .Y(n37) );
  AND2X4 U81 ( .A(B[6]), .B(n12), .Y(n64) );
  INVX1 U82 ( .A(A[6]), .Y(n12) );
  XOR2X2 U83 ( .A(n104), .B(n106), .Y(DIFF[4]) );
  NOR2X1 U84 ( .A(n149), .B(n150), .Y(n147) );
  NAND4X4 U85 ( .A(n216), .B(n194), .C(n76), .D(n73), .Y(n97) );
  DLY1X1 U86 ( .A(n97), .Y(n13) );
  NAND2X2 U87 ( .A(n53), .B(n56), .Y(n171) );
  XOR2X4 U88 ( .A(n195), .B(n4), .Y(DIFF[10]) );
  NAND3BX4 U89 ( .AN(n63), .B(n204), .C(n189), .Y(n62) );
  NAND2X4 U90 ( .A(n3), .B(n167), .Y(n151) );
  NAND2BX2 U91 ( .AN(n146), .B(n151), .Y(n143) );
  NAND2X2 U92 ( .A(n151), .B(n20), .Y(n164) );
  NAND2BX2 U93 ( .AN(B[13]), .B(A[13]), .Y(n134) );
  OR2X4 U94 ( .A(B[4]), .B(n16), .Y(n96) );
  INVX3 U95 ( .A(n178), .Y(n27) );
  NAND2BX2 U96 ( .AN(A[11]), .B(B[11]), .Y(n176) );
  NAND2BX2 U97 ( .AN(B[11]), .B(A[11]), .Y(n165) );
  BUFX12 U98 ( .A(n131), .Y(n21) );
  NAND2BX2 U99 ( .AN(A[13]), .B(B[13]), .Y(n131) );
  OAI2BB1X4 U100 ( .A0N(n34), .A1N(n35), .B0(n88), .Y(n85) );
  INVX2 U101 ( .A(n96), .Y(n105) );
  OAI2BB1X4 U102 ( .A0N(n17), .A1N(n18), .B0(n191), .Y(n157) );
  AND2X1 U103 ( .A(n95), .B(n94), .Y(n18) );
  CLKINVX2 U104 ( .A(B[3]), .Y(n212) );
  NOR2BX1 U105 ( .AN(B[3]), .B(A[3]), .Y(n215) );
  AND3X2 U106 ( .A(n27), .B(n87), .C(n15), .Y(n39) );
  NAND2BX4 U107 ( .AN(B[12]), .B(A[12]), .Y(n150) );
  NAND4X4 U108 ( .A(n97), .B(n95), .C(n94), .D(n78), .Y(n104) );
  OAI21X4 U109 ( .A0(n48), .A1(n49), .B0(n9), .Y(n204) );
  NOR2X4 U110 ( .A(B[6]), .B(n12), .Y(n19) );
  NAND2BX4 U111 ( .AN(A[7]), .B(B[7]), .Y(n190) );
  NOR2X4 U112 ( .A(n105), .B(n67), .Y(n106) );
  NOR2BX2 U113 ( .AN(n152), .B(n130), .Y(n25) );
  NAND3X4 U114 ( .A(n21), .B(n152), .C(n128), .Y(n146) );
  XNOR2X4 U115 ( .A(n22), .B(n180), .Y(DIFF[11]) );
  AND2X2 U116 ( .A(n165), .B(n176), .Y(n22) );
  XOR2X4 U117 ( .A(n23), .B(n24), .Y(DIFF[14]) );
  NAND2X4 U118 ( .A(n154), .B(n153), .Y(n23) );
  AND2X1 U119 ( .A(n128), .B(n133), .Y(n24) );
  NAND2X2 U120 ( .A(n91), .B(n90), .Y(n102) );
  NAND3X4 U121 ( .A(n96), .B(n97), .C(n78), .Y(n101) );
  NAND2X2 U122 ( .A(n43), .B(n170), .Y(n187) );
  AOI21X4 U123 ( .A0(n57), .A1(n58), .B0(n59), .Y(n55) );
  AOI2BB1X2 U124 ( .A0N(n90), .A1N(n64), .B0(n19), .Y(n88) );
  NAND2BXL U125 ( .AN(A[7]), .B(B[7]), .Y(n68) );
  INVX2 U126 ( .A(n86), .Y(n66) );
  NAND2BX4 U127 ( .AN(A[7]), .B(B[7]), .Y(n86) );
  NOR2BX4 U128 ( .AN(B[11]), .B(A[11]), .Y(n174) );
  NOR2X2 U129 ( .A(n19), .B(n60), .Y(n203) );
  NAND3X4 U130 ( .A(n145), .B(n143), .C(n144), .Y(n40) );
  NAND3BX2 U131 ( .AN(n136), .B(n142), .C(n26), .Y(n145) );
  AOI21X4 U132 ( .A0(n70), .A1(n69), .B0(n71), .Y(n57) );
  INVX4 U133 ( .A(n76), .Y(n74) );
  NAND2X2 U134 ( .A(n72), .B(n91), .Y(n71) );
  NOR2X4 U135 ( .A(n178), .B(n31), .Y(n186) );
  NAND2X2 U136 ( .A(n91), .B(n92), .Y(n100) );
  NAND2BX4 U137 ( .AN(B[3]), .B(A[3]), .Y(n78) );
  AOI21X4 U138 ( .A0(n42), .A1(n120), .B0(n121), .Y(n118) );
  NAND2BX4 U139 ( .AN(n122), .B(n123), .Y(n121) );
  NAND2BX4 U140 ( .AN(A[14]), .B(B[14]), .Y(n128) );
  NOR2X4 U141 ( .A(n64), .B(n65), .Y(n189) );
  INVX2 U142 ( .A(B[12]), .Y(n29) );
  AOI21X4 U143 ( .A0(n157), .A1(n186), .B0(n187), .Y(n181) );
  OAI21X4 U144 ( .A0(n99), .A1(n100), .B0(n90), .Y(n98) );
  NAND2XL U145 ( .A(n47), .B(n27), .Y(n140) );
  NOR2BX4 U146 ( .AN(n48), .B(A[5]), .Y(n188) );
  INVX8 U147 ( .A(n141), .Y(n178) );
  NOR2X4 U148 ( .A(n192), .B(n193), .Y(n191) );
  NAND2X2 U149 ( .A(n86), .B(n205), .Y(n193) );
  NAND2BX4 U150 ( .AN(A[5]), .B(n48), .Y(n91) );
  OAI2BB1X2 U151 ( .A0N(n39), .A1N(n157), .B0(n155), .Y(n154) );
  AOI21X2 U152 ( .A0(n44), .A1(n151), .B0(n158), .Y(n153) );
  AND2X2 U153 ( .A(n48), .B(n49), .Y(n63) );
  NOR2X4 U154 ( .A(n28), .B(n208), .Y(n200) );
  NAND2X2 U155 ( .A(n183), .B(n184), .Y(n182) );
  XOR2X4 U156 ( .A(n118), .B(n119), .Y(DIFF[16]) );
  AOI21X4 U157 ( .A0(n162), .A1(n26), .B0(n163), .Y(n161) );
  NAND2BX4 U158 ( .AN(n48), .B(A[5]), .Y(n90) );
  NAND2XL U159 ( .A(n128), .B(n129), .Y(n126) );
  NAND2BX2 U160 ( .AN(B[14]), .B(A[14]), .Y(n133) );
  AOI21X2 U161 ( .A0(n147), .A1(n21), .B0(n148), .Y(n144) );
  AND2X4 U162 ( .A(n61), .B(n87), .Y(n47) );
  NOR2X4 U163 ( .A(B[8]), .B(n33), .Y(n32) );
  CLKINVX20 U164 ( .A(A[8]), .Y(n33) );
  NOR2X4 U165 ( .A(n178), .B(n31), .Y(n177) );
  XOR2X4 U166 ( .A(n103), .B(n102), .Y(DIFF[5]) );
  NAND3X1 U167 ( .A(n92), .B(n89), .C(n6), .Y(n208) );
  XOR2X4 U168 ( .A(n26), .B(n83), .Y(DIFF[8]) );
  OR2X4 U169 ( .A(n93), .B(n101), .Y(n34) );
  INVX4 U170 ( .A(n128), .Y(n149) );
  NAND3X2 U171 ( .A(n165), .B(n166), .C(n167), .Y(n138) );
  NAND3X4 U172 ( .A(n170), .B(n171), .C(n172), .Y(n167) );
  NOR2X1 U173 ( .A(n156), .B(n136), .Y(n155) );
  OAI21X1 U174 ( .A0(n135), .A1(n136), .B0(n137), .Y(n120) );
  INVX4 U175 ( .A(n124), .Y(n36) );
  INVX8 U176 ( .A(n84), .Y(n54) );
  NAND2BX4 U177 ( .AN(A[8]), .B(B[8]), .Y(n84) );
  AOI21X1 U178 ( .A0(n130), .A1(n21), .B0(n132), .Y(n125) );
  XOR2X4 U179 ( .A(n85), .B(n1), .Y(DIFF[7]) );
  NAND2X1 U180 ( .A(n78), .B(n79), .Y(n77) );
  AND2X2 U181 ( .A(n94), .B(n78), .Y(n46) );
  INVX2 U182 ( .A(n78), .Y(n211) );
  AOI21X1 U183 ( .A0(n75), .A1(n76), .B0(n77), .Y(n69) );
  INVX4 U184 ( .A(n87), .Y(n60) );
  NOR2X4 U185 ( .A(n200), .B(n201), .Y(n197) );
  NAND2X4 U186 ( .A(n175), .B(n176), .Y(n166) );
  NAND2BX4 U187 ( .AN(A[10]), .B(B[10]), .Y(n170) );
  NOR2X4 U188 ( .A(n181), .B(n182), .Y(n180) );
  NAND2X1 U189 ( .A(n133), .B(n134), .Y(n132) );
  OAI21X1 U190 ( .A0(n149), .A1(n134), .B0(n133), .Y(n148) );
  INVX4 U191 ( .A(n179), .Y(n52) );
  OAI21X4 U192 ( .A0(n197), .A1(n198), .B0(n199), .Y(n195) );
  NOR2X2 U193 ( .A(n173), .B(n174), .Y(n172) );
  INVX4 U194 ( .A(n190), .Y(n65) );
  OAI21X4 U195 ( .A0(n55), .A1(n54), .B0(n56), .Y(n50) );
  NAND4BX4 U196 ( .AN(n80), .B(n72), .C(n216), .D(n76), .Y(n95) );
  NAND4BX1 U197 ( .AN(n95), .B(n45), .C(n124), .D(n42), .Y(n123) );
  NOR2X2 U198 ( .A(n101), .B(n93), .Y(n99) );
  XOR2X4 U199 ( .A(n40), .B(n41), .Y(DIFF[15]) );
  XOR2X4 U200 ( .A(n161), .B(n160), .Y(DIFF[13]) );
  OAI21X4 U201 ( .A0(n112), .A1(n81), .B0(n11), .Y(n109) );
  NAND3BX4 U202 ( .AN(n188), .B(n204), .C(n189), .Y(n141) );
  NOR2X4 U203 ( .A(n36), .B(n37), .Y(n38) );
  NOR2X4 U204 ( .A(n38), .B(n138), .Y(n169) );
  NAND2X4 U205 ( .A(n113), .B(n116), .Y(n73) );
  NAND2X4 U206 ( .A(n110), .B(n194), .Y(n94) );
  AND2X2 U207 ( .A(n20), .B(n21), .Y(n44) );
  NAND2BX2 U208 ( .AN(A[0]), .B(B[0]), .Y(n117) );
  AOI2BB1XL U209 ( .A0N(A[3]), .A1N(n212), .B0(n80), .Y(n209) );
  INVX2 U210 ( .A(n114), .Y(n112) );
  NAND2XL U211 ( .A(n21), .B(n134), .Y(n160) );
  NAND2XL U212 ( .A(n46), .B(n13), .Y(n139) );
  INVXL U213 ( .A(A[5]), .Y(n49) );
  INVX1 U214 ( .A(n138), .Y(n137) );
  INVX1 U215 ( .A(n170), .Y(n196) );
  XOR2X2 U216 ( .A(n107), .B(n108), .Y(DIFF[3]) );
  AOI21X1 U217 ( .A0(n45), .A1(n139), .B0(n140), .Y(n135) );
  INVX1 U218 ( .A(n152), .Y(n168) );
  NAND2X1 U219 ( .A(n21), .B(n20), .Y(n156) );
  INVX4 U220 ( .A(n79), .Y(n110) );
  AND4X1 U221 ( .A(n91), .B(n68), .C(n92), .D(n89), .Y(n45) );
  INVX1 U222 ( .A(n117), .Y(n80) );
  NAND2X1 U223 ( .A(n117), .B(n116), .Y(DIFF[0]) );
  NAND2BX1 U224 ( .AN(n117), .B(n116), .Y(n114) );
  XOR2X1 U225 ( .A(B[16]), .B(A[16]), .Y(n119) );
  NOR3X2 U226 ( .A(n66), .B(n64), .C(n67), .Y(n58) );
  XOR2X4 U227 ( .A(n50), .B(n51), .Y(DIFF[9]) );
  NAND2X4 U228 ( .A(n157), .B(n177), .Y(n82) );
  NAND4BX4 U229 ( .AN(n174), .B(n170), .C(n179), .D(n84), .Y(n136) );
  NAND2X4 U230 ( .A(n19), .B(n86), .Y(n61) );
  NAND2BX4 U231 ( .AN(B[7]), .B(A[7]), .Y(n87) );
  NAND2BX4 U232 ( .AN(A[4]), .B(B[4]), .Y(n92) );
  NAND2BX4 U233 ( .AN(B[2]), .B(A[2]), .Y(n79) );
  NAND2BX4 U234 ( .AN(A[2]), .B(B[2]), .Y(n76) );
  NAND2BX4 U235 ( .AN(B[1]), .B(A[1]), .Y(n113) );
endmodule


module butterfly_DW01_add_164 ( A, B, SUM );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220;

  AOI2BB1X2 U2 ( .A0N(A[1]), .A1N(B[1]), .B0(n64), .Y(n214) );
  CLKINVX3 U3 ( .A(n46), .Y(n1) );
  CLKINVX8 U4 ( .A(n38), .Y(n131) );
  INVX2 U5 ( .A(B[10]), .Y(n14) );
  NAND2X1 U6 ( .A(n149), .B(n173), .Y(n144) );
  NAND2X4 U7 ( .A(n54), .B(n85), .Y(n177) );
  INVX4 U8 ( .A(n201), .Y(n12) );
  NOR2BX2 U9 ( .AN(n131), .B(n151), .Y(n146) );
  CLKINVX3 U10 ( .A(n182), .Y(n33) );
  BUFX3 U11 ( .A(n152), .Y(n25) );
  INVX8 U12 ( .A(n154), .Y(n182) );
  NAND2X1 U13 ( .A(n127), .B(n128), .Y(n150) );
  OR2X4 U14 ( .A(B[13]), .B(A[13]), .Y(n132) );
  NOR2X4 U15 ( .A(n164), .B(n42), .Y(n163) );
  BUFX12 U16 ( .A(n19), .Y(n2) );
  OAI21XL U17 ( .A0(n119), .A1(n120), .B0(n121), .Y(n118) );
  OAI21X2 U18 ( .A0(n83), .A1(n84), .B0(n85), .Y(n79) );
  CLKINVX3 U19 ( .A(n26), .Y(n68) );
  INVX4 U20 ( .A(n27), .Y(n11) );
  INVX1 U21 ( .A(n36), .Y(n157) );
  INVX1 U22 ( .A(n127), .Y(n42) );
  XOR2X1 U23 ( .A(B[16]), .B(A[16]), .Y(n114) );
  INVX1 U24 ( .A(n118), .Y(n117) );
  NAND3BX4 U25 ( .AN(n3), .B(n214), .C(n211), .Y(n141) );
  NAND2X2 U26 ( .A(n212), .B(n213), .Y(n3) );
  NAND2X1 U27 ( .A(n30), .B(n127), .Y(n4) );
  NAND2X2 U28 ( .A(A[10]), .B(B[10]), .Y(n192) );
  NAND3BX4 U29 ( .AN(n5), .B(n59), .C(n218), .Y(n216) );
  NOR2X2 U30 ( .A(n39), .B(n200), .Y(n5) );
  NAND2XL U31 ( .A(B[3]), .B(A[3]), .Y(n101) );
  NAND2X1 U32 ( .A(n13), .B(n14), .Y(n6) );
  NAND3BX4 U33 ( .AN(n2), .B(n17), .C(n131), .Y(n166) );
  INVX4 U34 ( .A(n2), .Y(n30) );
  NOR3X2 U35 ( .A(n176), .B(n45), .C(n177), .Y(n193) );
  BUFX8 U36 ( .A(n78), .Y(n7) );
  CLKINVX8 U37 ( .A(n37), .Y(n85) );
  NAND4X4 U38 ( .A(n8), .B(n209), .C(n7), .D(n35), .Y(n34) );
  AND2X4 U39 ( .A(n136), .B(n40), .Y(n8) );
  NAND2X2 U40 ( .A(B[13]), .B(A[13]), .Y(n127) );
  OAI21XL U41 ( .A0(n137), .A1(n138), .B0(n61), .Y(n135) );
  NOR2X2 U42 ( .A(n62), .B(n63), .Y(n61) );
  OR2X2 U43 ( .A(n82), .B(n11), .Y(n63) );
  NAND2X2 U44 ( .A(n86), .B(n27), .Y(n84) );
  CLKINVX8 U45 ( .A(n190), .Y(n9) );
  CLKINVX3 U46 ( .A(n190), .Y(n23) );
  NAND3X4 U47 ( .A(n33), .B(n25), .C(n153), .Y(n134) );
  AOI21X2 U48 ( .A0(n87), .A1(n88), .B0(n89), .Y(n83) );
  OAI21X1 U49 ( .A0(n69), .A1(n190), .B0(n192), .Y(n199) );
  NAND3X2 U50 ( .A(n72), .B(n34), .C(n71), .Y(n67) );
  CLKINVX8 U51 ( .A(n129), .Y(n173) );
  OR2X2 U52 ( .A(B[9]), .B(A[9]), .Y(n10) );
  NAND3XL U53 ( .A(n29), .B(n27), .C(n87), .Y(n156) );
  NOR2X4 U54 ( .A(n94), .B(n196), .Y(n195) );
  AND2X4 U55 ( .A(B[6]), .B(A[6]), .Y(n37) );
  INVX12 U56 ( .A(n60), .Y(n27) );
  BUFX12 U57 ( .A(A[5]), .Y(n66) );
  AOI31X2 U58 ( .A0(n74), .A1(n12), .A2(n215), .B0(n199), .Y(n198) );
  NAND2X4 U59 ( .A(n13), .B(n14), .Y(n167) );
  INVX8 U60 ( .A(A[10]), .Y(n13) );
  AOI21X4 U61 ( .A0(n52), .A1(n171), .B0(n172), .Y(n170) );
  INVX8 U62 ( .A(n31), .Y(n210) );
  NAND2X4 U63 ( .A(n173), .B(n186), .Y(n185) );
  INVXL U64 ( .A(n10), .Y(n47) );
  NAND3X4 U65 ( .A(n15), .B(n40), .C(n219), .Y(n218) );
  OR2X4 U66 ( .A(n66), .B(n65), .Y(n15) );
  BUFX12 U67 ( .A(B[5]), .Y(n65) );
  INVX4 U68 ( .A(n22), .Y(n16) );
  CLKINVX8 U69 ( .A(n16), .Y(n17) );
  DLY1X1 U70 ( .A(n141), .Y(n18) );
  NOR2X4 U71 ( .A(n82), .B(n175), .Y(n186) );
  INVX8 U72 ( .A(n44), .Y(n22) );
  CLKINVX8 U73 ( .A(n50), .Y(n39) );
  INVX3 U74 ( .A(n35), .Y(n20) );
  NAND2X4 U75 ( .A(n66), .B(n65), .Y(n200) );
  OR2XL U76 ( .A(n1), .B(n206), .Y(n26) );
  OAI21X2 U77 ( .A0(n155), .A1(n53), .B0(n186), .Y(n143) );
  NAND2XL U78 ( .A(n140), .B(n31), .Y(n138) );
  NAND2X1 U79 ( .A(n66), .B(n65), .Y(n32) );
  INVX8 U80 ( .A(n49), .Y(n136) );
  INVX8 U81 ( .A(n39), .Y(n40) );
  NAND3BX2 U82 ( .AN(n210), .B(n140), .C(n141), .Y(n36) );
  AOI21X4 U83 ( .A0(n184), .A1(n52), .B0(n185), .Y(n179) );
  NOR2X4 U84 ( .A(B[13]), .B(A[13]), .Y(n19) );
  NAND2BX2 U85 ( .AN(n94), .B(n21), .Y(n77) );
  NOR2X1 U86 ( .A(n196), .B(n20), .Y(n21) );
  NAND2BX4 U87 ( .AN(n192), .B(n22), .Y(n152) );
  INVX8 U88 ( .A(n167), .Y(n190) );
  NAND2X1 U89 ( .A(A[9]), .B(B[9]), .Y(n69) );
  NAND4BX2 U90 ( .AN(n60), .B(n15), .C(B[4]), .D(A[4]), .Y(n24) );
  NOR2X2 U91 ( .A(B[6]), .B(A[6]), .Y(n60) );
  INVX4 U92 ( .A(n69), .Y(n206) );
  INVX8 U93 ( .A(n24), .Y(n176) );
  OR2X4 U94 ( .A(n66), .B(n65), .Y(n43) );
  NOR3X4 U95 ( .A(n176), .B(n45), .C(n177), .Y(n184) );
  NOR2X2 U96 ( .A(n210), .B(n102), .Y(n100) );
  OAI2BB1X2 U97 ( .A0N(n107), .A1N(n108), .B0(n109), .Y(n105) );
  INVX8 U98 ( .A(n73), .Y(n215) );
  NAND3X1 U99 ( .A(n23), .B(n46), .C(n169), .Y(n165) );
  NOR2X2 U100 ( .A(n2), .B(n128), .Y(n124) );
  CLKBUFXL U101 ( .A(n173), .Y(n28) );
  AND2X1 U102 ( .A(B[4]), .B(A[4]), .Y(n219) );
  NAND2X2 U103 ( .A(B[4]), .B(A[4]), .Y(n90) );
  NOR3BX4 U104 ( .AN(n131), .B(n2), .C(n82), .Y(n174) );
  CLKINVX8 U105 ( .A(n131), .Y(n175) );
  NAND4BX4 U106 ( .AN(n60), .B(n29), .C(B[4]), .D(A[4]), .Y(n159) );
  OR2X4 U107 ( .A(n66), .B(n65), .Y(n29) );
  NAND2BX2 U108 ( .AN(n73), .B(n74), .Y(n72) );
  NOR3X4 U109 ( .A(n176), .B(n45), .C(n177), .Y(n171) );
  BUFX8 U110 ( .A(n158), .Y(n45) );
  OR2X4 U111 ( .A(B[6]), .B(A[6]), .Y(n50) );
  BUFX4 U112 ( .A(n101), .Y(n31) );
  INVX1 U113 ( .A(n28), .Y(n51) );
  NAND2X2 U114 ( .A(n173), .B(n136), .Y(n194) );
  NAND2X4 U115 ( .A(n136), .B(n40), .Y(n196) );
  NOR2X2 U116 ( .A(n156), .B(n157), .Y(n155) );
  AND2X4 U117 ( .A(n32), .B(n43), .Y(n56) );
  OAI21X2 U118 ( .A0(n103), .A1(n64), .B0(n104), .Y(n99) );
  INVX2 U119 ( .A(n105), .Y(n103) );
  NAND3BX4 U120 ( .AN(n210), .B(n140), .C(n141), .Y(n35) );
  NAND2BX2 U121 ( .AN(A[1]), .B(n112), .Y(n212) );
  NOR2X4 U122 ( .A(B[12]), .B(A[12]), .Y(n38) );
  OAI2BB1X2 U123 ( .A0N(B[9]), .A1N(A[9]), .B0(n191), .Y(n169) );
  NAND2BX4 U124 ( .AN(B[1]), .B(n112), .Y(n213) );
  INVX8 U125 ( .A(n70), .Y(n46) );
  INVX2 U126 ( .A(n123), .Y(n58) );
  NAND2X1 U127 ( .A(B[15]), .B(A[15]), .Y(n121) );
  NAND2X2 U128 ( .A(n6), .B(n10), .Y(n201) );
  XOR2X4 U129 ( .A(n41), .B(n75), .Y(SUM[8]) );
  AND2X1 U130 ( .A(n7), .B(n71), .Y(n41) );
  NOR2X2 U131 ( .A(n133), .B(n134), .Y(n115) );
  AOI21XL U132 ( .A0(n135), .A1(n76), .B0(n51), .Y(n133) );
  BUFX20 U133 ( .A(n81), .Y(n54) );
  NAND2X4 U134 ( .A(B[7]), .B(A[7]), .Y(n81) );
  OAI2BB1X4 U135 ( .A0N(n149), .A1N(n150), .B0(n126), .Y(n148) );
  NOR2X4 U136 ( .A(B[11]), .B(A[11]), .Y(n44) );
  NAND3X4 U137 ( .A(A[2]), .B(n211), .C(B[2]), .Y(n140) );
  INVX2 U138 ( .A(n211), .Y(n102) );
  NOR2BX2 U139 ( .AN(n85), .B(n11), .Y(n92) );
  XOR2X4 U140 ( .A(n178), .B(n4), .Y(SUM[13]) );
  XOR2X1 U141 ( .A(n35), .B(n97), .Y(SUM[4]) );
  OR2X2 U142 ( .A(A[14]), .B(B[14]), .Y(n122) );
  INVXL U143 ( .A(n18), .Y(n137) );
  OAI21X4 U144 ( .A0(A[14]), .A1(B[14]), .B0(n132), .Y(n151) );
  NAND2X4 U145 ( .A(n87), .B(n86), .Y(n94) );
  XOR2X4 U146 ( .A(n55), .B(n48), .Y(SUM[11]) );
  AND2X1 U147 ( .A(n17), .B(n153), .Y(n48) );
  NAND2XL U148 ( .A(n126), .B(n127), .Y(n125) );
  NAND2X2 U149 ( .A(n36), .B(n87), .Y(n96) );
  NOR2X4 U150 ( .A(A[7]), .B(B[7]), .Y(n49) );
  NAND2X2 U151 ( .A(n90), .B(n96), .Y(n95) );
  NAND2XL U152 ( .A(n192), .B(n23), .Y(n204) );
  XOR2X2 U153 ( .A(n105), .B(n106), .Y(SUM[2]) );
  NOR2BX2 U154 ( .AN(n104), .B(n64), .Y(n106) );
  NAND4BBX4 U155 ( .AN(n158), .BN(n37), .C(n159), .D(n54), .Y(n74) );
  XOR2X4 U156 ( .A(n95), .B(n56), .Y(SUM[5]) );
  NOR2X4 U157 ( .A(n202), .B(n203), .Y(n197) );
  NOR2BX2 U158 ( .AN(n54), .B(n82), .Y(n80) );
  AND2X4 U159 ( .A(n54), .B(n85), .Y(n59) );
  INVX4 U160 ( .A(n151), .Y(n149) );
  NOR2X2 U161 ( .A(n201), .B(n71), .Y(n203) );
  NOR2X4 U162 ( .A(n34), .B(n201), .Y(n202) );
  OAI21X4 U163 ( .A0(n93), .A1(n94), .B0(n32), .Y(n91) );
  AOI21X4 U164 ( .A0(n208), .A1(n34), .B0(n47), .Y(n207) );
  OAI21X4 U165 ( .A0(n181), .A1(n175), .B0(n128), .Y(n180) );
  NAND2X2 U166 ( .A(B[14]), .B(A[14]), .Y(n126) );
  NAND3X1 U167 ( .A(n153), .B(n154), .C(n152), .Y(n147) );
  NAND2X2 U168 ( .A(B[8]), .B(A[8]), .Y(n191) );
  OR2X4 U169 ( .A(B[3]), .B(A[3]), .Y(n211) );
  NAND2X4 U170 ( .A(n173), .B(n174), .Y(n172) );
  NAND2X2 U171 ( .A(B[11]), .B(A[11]), .Y(n153) );
  INVX8 U172 ( .A(n168), .Y(n70) );
  AOI21X4 U173 ( .A0(n216), .A1(n215), .B0(n217), .Y(n208) );
  NAND2X4 U174 ( .A(n76), .B(n52), .Y(n75) );
  NAND2XL U175 ( .A(n122), .B(n123), .Y(n120) );
  INVX2 U176 ( .A(n122), .Y(n130) );
  NAND2X2 U177 ( .A(B[12]), .B(A[12]), .Y(n128) );
  NOR2BX4 U178 ( .AN(n90), .B(n88), .Y(n93) );
  NAND2X4 U179 ( .A(n195), .B(n88), .Y(n52) );
  NAND4BX4 U180 ( .AN(n158), .B(n159), .C(n54), .D(n85), .Y(n53) );
  NAND2X1 U181 ( .A(n131), .B(n128), .Y(n187) );
  NAND2X4 U182 ( .A(n197), .B(n198), .Y(n55) );
  NOR2X4 U183 ( .A(n170), .B(n124), .Y(n162) );
  OR2X4 U184 ( .A(A[15]), .B(B[15]), .Y(n123) );
  INVX4 U185 ( .A(n43), .Y(n139) );
  NOR2X4 U186 ( .A(n139), .B(n98), .Y(n209) );
  NAND2X1 U187 ( .A(n200), .B(n90), .Y(n89) );
  NOR2X4 U188 ( .A(A[2]), .B(B[2]), .Y(n64) );
  XOR2X4 U189 ( .A(n205), .B(n204), .Y(SUM[10]) );
  NOR2X4 U190 ( .A(n207), .B(n206), .Y(n205) );
  NAND2X4 U191 ( .A(n78), .B(n136), .Y(n73) );
  INVX8 U192 ( .A(n136), .Y(n82) );
  OR2X4 U193 ( .A(A[9]), .B(B[9]), .Y(n168) );
  OR2X2 U194 ( .A(A[1]), .B(B[1]), .Y(n107) );
  XOR2X4 U195 ( .A(n108), .B(n110), .Y(SUM[1]) );
  NOR2BX4 U196 ( .AN(n109), .B(n111), .Y(n110) );
  NOR2BX2 U197 ( .AN(n90), .B(n98), .Y(n97) );
  NAND2X2 U198 ( .A(B[8]), .B(A[8]), .Y(n71) );
  NOR2X4 U199 ( .A(n200), .B(n39), .Y(n158) );
  OR2X4 U200 ( .A(n66), .B(n65), .Y(n86) );
  NAND4BX4 U201 ( .AN(n190), .B(n22), .C(n46), .D(n169), .Y(n154) );
  NAND2X4 U202 ( .A(n53), .B(n136), .Y(n76) );
  NOR2BX4 U203 ( .AN(n121), .B(n58), .Y(n57) );
  NOR2BX4 U204 ( .AN(n126), .B(n130), .Y(n161) );
  NAND2XL U205 ( .A(B[1]), .B(A[1]), .Y(n109) );
  OAI21X4 U206 ( .A0(n115), .A1(n116), .B0(n117), .Y(n113) );
  OR2X2 U207 ( .A(n139), .B(n98), .Y(n62) );
  INVX1 U208 ( .A(n71), .Y(n217) );
  INVX1 U209 ( .A(n107), .Y(n111) );
  NOR2X1 U210 ( .A(n124), .B(n125), .Y(n119) );
  NAND2XL U211 ( .A(B[2]), .B(A[2]), .Y(n104) );
  INVX1 U212 ( .A(n112), .Y(n108) );
  NAND2X1 U213 ( .A(B[0]), .B(A[0]), .Y(n112) );
  AND2X2 U214 ( .A(n112), .B(n220), .Y(SUM[0]) );
  OR2X2 U215 ( .A(A[0]), .B(B[0]), .Y(n220) );
  NAND3BX4 U216 ( .AN(n210), .B(n141), .C(n140), .Y(n88) );
  NAND4BXL U217 ( .AN(n130), .B(n123), .C(n131), .D(n30), .Y(n116) );
  INVX8 U218 ( .A(n87), .Y(n98) );
  XOR2X4 U219 ( .A(n67), .B(n68), .Y(SUM[9]) );
  XOR2X4 U220 ( .A(n79), .B(n80), .Y(SUM[7]) );
  XOR2X4 U221 ( .A(n91), .B(n92), .Y(SUM[6]) );
  XOR2X4 U222 ( .A(n99), .B(n100), .Y(SUM[3]) );
  XOR2X4 U223 ( .A(n113), .B(n114), .Y(SUM[16]) );
  XOR2X4 U224 ( .A(n142), .B(n57), .Y(SUM[15]) );
  OAI21X4 U225 ( .A0(n143), .A1(n144), .B0(n145), .Y(n142) );
  AOI21X4 U226 ( .A0(n147), .A1(n146), .B0(n148), .Y(n145) );
  XOR2X4 U227 ( .A(n160), .B(n161), .Y(SUM[14]) );
  NAND2X4 U228 ( .A(n162), .B(n163), .Y(n160) );
  AOI31X2 U229 ( .A0(n165), .A1(n153), .A2(n152), .B0(n166), .Y(n164) );
  NOR2X4 U230 ( .A(n180), .B(n179), .Y(n178) );
  NOR2X4 U231 ( .A(n183), .B(n182), .Y(n181) );
  NAND2X4 U232 ( .A(n153), .B(n152), .Y(n183) );
  XOR2X4 U233 ( .A(n188), .B(n187), .Y(SUM[12]) );
  NOR2X4 U234 ( .A(n189), .B(n134), .Y(n188) );
  AOI21X4 U235 ( .A0(n77), .A1(n193), .B0(n194), .Y(n189) );
  NAND4BX4 U236 ( .AN(n70), .B(n22), .C(n9), .D(n78), .Y(n129) );
  OR2X4 U237 ( .A(A[4]), .B(B[4]), .Y(n87) );
  OR2X4 U238 ( .A(A[8]), .B(B[8]), .Y(n78) );
endmodule


module butterfly_DW01_add_170 ( A, B, SUM );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  wire   n186, n187, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185;

  INVX4 U2 ( .A(n19), .Y(n56) );
  AND2X4 U3 ( .A(B[7]), .B(A[7]), .Y(n21) );
  INVX8 U4 ( .A(n72), .Y(n63) );
  NAND2X1 U5 ( .A(B[15]), .B(A[15]), .Y(n102) );
  NOR2X4 U6 ( .A(A[13]), .B(B[13]), .Y(n1) );
  NOR2BX2 U7 ( .AN(n155), .B(n150), .Y(n167) );
  NOR2X4 U8 ( .A(B[3]), .B(A[3]), .Y(n183) );
  INVX8 U9 ( .A(n8), .Y(n170) );
  NAND3X2 U10 ( .A(n24), .B(n50), .C(n51), .Y(n164) );
  OAI2BB1X4 U11 ( .A0N(n46), .A1N(n47), .B0(n48), .Y(n43) );
  CLKINVX3 U12 ( .A(n90), .Y(n12) );
  INVX4 U13 ( .A(n21), .Y(n50) );
  NOR2BX2 U14 ( .AN(n81), .B(n87), .Y(n86) );
  INVXL U15 ( .A(B[5]), .Y(n23) );
  INVX1 U16 ( .A(A[5]), .Y(n22) );
  NAND2X2 U17 ( .A(B[11]), .B(A[11]), .Y(n154) );
  OR2X2 U18 ( .A(n130), .B(n25), .Y(n36) );
  NAND2X1 U19 ( .A(n107), .B(n108), .Y(n106) );
  NAND2X2 U20 ( .A(B[8]), .B(A[8]), .Y(n48) );
  BUFX16 U21 ( .A(n186), .Y(SUM[10]) );
  INVX1 U22 ( .A(n64), .Y(n70) );
  NOR2BX2 U23 ( .AN(n108), .B(n1), .Y(n140) );
  OR2X2 U24 ( .A(A[12]), .B(B[12]), .Y(n111) );
  AOI21X1 U25 ( .A0(n53), .A1(n116), .B0(n14), .Y(n113) );
  INVXL U26 ( .A(n118), .Y(n53) );
  NOR2BX2 U27 ( .AN(n50), .B(n56), .Y(n55) );
  OAI21X2 U28 ( .A0(n57), .A1(n58), .B0(n59), .Y(n54) );
  AOI21X2 U29 ( .A0(n60), .A1(n31), .B0(n62), .Y(n57) );
  INVX1 U30 ( .A(n85), .Y(n74) );
  OR2X4 U31 ( .A(A[11]), .B(B[11]), .Y(n2) );
  NAND2X1 U32 ( .A(n48), .B(n47), .Y(n3) );
  NOR2BXL U33 ( .AN(n20), .B(B[10]), .Y(n157) );
  AND2X1 U34 ( .A(B[9]), .B(A[9]), .Y(n33) );
  NAND2X4 U35 ( .A(n42), .B(n164), .Y(n158) );
  XOR2X4 U36 ( .A(n4), .B(n121), .Y(SUM[15]) );
  NAND3X4 U37 ( .A(n123), .B(n125), .C(n124), .Y(n4) );
  OAI21X2 U38 ( .A0(n63), .A1(n64), .B0(n65), .Y(n62) );
  AND2X2 U39 ( .A(n109), .B(n111), .Y(n10) );
  NAND2X4 U40 ( .A(B[3]), .B(A[3]), .Y(n85) );
  INVX4 U41 ( .A(n51), .Y(n145) );
  NAND4BX4 U42 ( .AN(n157), .B(n2), .C(n47), .D(n30), .Y(n110) );
  INVX1 U43 ( .A(A[10]), .Y(n20) );
  OAI2BB2X4 U44 ( .B0(A[14]), .B1(B[14]), .A0N(n5), .A1N(n6), .Y(n129) );
  INVX1 U45 ( .A(A[13]), .Y(n5) );
  CLKINVX2 U46 ( .A(B[13]), .Y(n6) );
  NAND2BX4 U47 ( .AN(n6), .B(A[13]), .Y(n108) );
  NOR3BX2 U48 ( .AN(n111), .B(n1), .C(n110), .Y(n135) );
  AOI2BB1X2 U49 ( .A0N(B[3]), .A1N(A[3]), .B0(n93), .Y(n184) );
  XOR2X4 U50 ( .A(n3), .B(n7), .Y(SUM[8]) );
  NOR2X4 U51 ( .A(n118), .B(n170), .Y(n7) );
  AND2X2 U52 ( .A(n107), .B(n103), .Y(n134) );
  OR2X4 U53 ( .A(B[9]), .B(A[9]), .Y(n45) );
  INVX4 U54 ( .A(n69), .Y(n66) );
  INVXL U55 ( .A(n129), .Y(n112) );
  NOR3X2 U56 ( .A(n129), .B(n25), .C(n110), .Y(n132) );
  NAND2X4 U57 ( .A(n48), .B(n50), .Y(n173) );
  NAND2XL U58 ( .A(B[2]), .B(A[2]), .Y(n81) );
  OAI21X4 U59 ( .A0(n178), .A1(n179), .B0(n180), .Y(n8) );
  INVXL U60 ( .A(n115), .Y(n114) );
  NAND2BX4 U61 ( .AN(B[10]), .B(n20), .Y(n165) );
  NAND2X4 U62 ( .A(n11), .B(n155), .Y(n163) );
  NAND2X4 U63 ( .A(n149), .B(n148), .Y(n9) );
  XOR2X4 U64 ( .A(n146), .B(n10), .Y(SUM[12]) );
  OR2X4 U65 ( .A(n162), .B(n48), .Y(n11) );
  AOI2BB1X4 U66 ( .A0N(n15), .A1N(n44), .B0(n163), .Y(n159) );
  NOR2BX1 U67 ( .AN(n90), .B(n92), .Y(n91) );
  NAND2X4 U68 ( .A(n51), .B(n172), .Y(n171) );
  INVX8 U69 ( .A(n165), .Y(n150) );
  OAI21X2 U70 ( .A0(n71), .A1(n63), .B0(n65), .Y(n67) );
  NAND2X2 U71 ( .A(B[1]), .B(A[1]), .Y(n90) );
  NOR2X4 U72 ( .A(n87), .B(n92), .Y(n185) );
  NAND2X2 U73 ( .A(B[0]), .B(A[0]), .Y(n93) );
  OR2X4 U74 ( .A(A[9]), .B(B[9]), .Y(n30) );
  NAND2X4 U75 ( .A(n13), .B(n12), .Y(n78) );
  NOR2X4 U76 ( .A(n87), .B(n183), .Y(n13) );
  INVX1 U77 ( .A(n147), .Y(n14) );
  INVX2 U78 ( .A(n110), .Y(n147) );
  NAND2X4 U79 ( .A(n81), .B(n82), .Y(n80) );
  OAI21X2 U80 ( .A0(n1), .A1(n109), .B0(n108), .Y(n138) );
  INVX4 U81 ( .A(n17), .Y(n109) );
  CLKINVX2 U82 ( .A(n161), .Y(n15) );
  INVX8 U83 ( .A(n162), .Y(n161) );
  NOR2BX4 U84 ( .AN(n78), .B(n77), .Y(n18) );
  AND2X2 U85 ( .A(B[12]), .B(A[12]), .Y(n17) );
  NAND3BX4 U86 ( .AN(n74), .B(n18), .C(n75), .Y(n31) );
  OR2X4 U87 ( .A(A[7]), .B(B[7]), .Y(n19) );
  OR2X2 U88 ( .A(A[7]), .B(B[7]), .Y(n174) );
  OAI2BB1X4 U89 ( .A0N(n22), .A1N(n23), .B0(n177), .Y(n181) );
  CLKINVX3 U90 ( .A(n120), .Y(n24) );
  INVX8 U91 ( .A(n49), .Y(n120) );
  NOR2X4 U92 ( .A(A[12]), .B(B[12]), .Y(n25) );
  NAND2X2 U93 ( .A(B[14]), .B(A[14]), .Y(n107) );
  INVX4 U94 ( .A(n33), .Y(n44) );
  NOR2BX4 U95 ( .AN(n26), .B(n145), .Y(n144) );
  AND2X2 U96 ( .A(n49), .B(n50), .Y(n26) );
  NAND3BX2 U97 ( .AN(n52), .B(n47), .C(n161), .Y(n160) );
  AOI21X4 U98 ( .A0(n9), .A1(n143), .B0(n17), .Y(n142) );
  XOR2X4 U99 ( .A(n27), .B(n28), .Y(SUM[11]) );
  NAND3X4 U100 ( .A(n159), .B(n158), .C(n160), .Y(n27) );
  AND2X1 U101 ( .A(n154), .B(n156), .Y(n28) );
  NOR2X4 U102 ( .A(n56), .B(n58), .Y(n29) );
  NOR2X2 U103 ( .A(n66), .B(n63), .Y(n60) );
  OAI2BB1X4 U104 ( .A0N(n135), .A1N(n131), .B0(n136), .Y(n133) );
  NOR2X2 U105 ( .A(n130), .B(n25), .Y(n143) );
  BUFX8 U106 ( .A(n187), .Y(SUM[5]) );
  OAI21X4 U107 ( .A0(n168), .A1(n169), .B0(n44), .Y(n166) );
  NOR2X4 U108 ( .A(n170), .B(n171), .Y(n168) );
  NAND2X4 U109 ( .A(n175), .B(n29), .Y(n34) );
  NAND4X4 U110 ( .A(n52), .B(n34), .C(n24), .D(n50), .Y(n46) );
  XNOR2X4 U111 ( .A(n79), .B(n80), .Y(SUM[3]) );
  NOR2X2 U112 ( .A(n25), .B(n110), .Y(n141) );
  AND2X2 U113 ( .A(n44), .B(n30), .Y(n37) );
  NAND3BX4 U114 ( .AN(n150), .B(n30), .C(n151), .Y(n149) );
  INVX4 U115 ( .A(n84), .Y(n87) );
  AOI21X4 U116 ( .A0(n61), .A1(n69), .B0(n70), .Y(n71) );
  NAND2BX2 U117 ( .AN(n77), .B(n78), .Y(n179) );
  INVX8 U118 ( .A(n177), .Y(n58) );
  NAND2X4 U119 ( .A(n144), .B(n8), .Y(n131) );
  OAI21XL U120 ( .A0(B[3]), .A1(A[3]), .B0(n85), .Y(n79) );
  NAND2X4 U121 ( .A(n69), .B(n174), .Y(n182) );
  NAND2X4 U122 ( .A(n119), .B(n34), .Y(n118) );
  OAI2BB1X4 U123 ( .A0N(n141), .A1N(n131), .B0(n142), .Y(n139) );
  NOR2X4 U124 ( .A(n181), .B(n182), .Y(n180) );
  NOR2BX1 U125 ( .AN(n59), .B(n58), .Y(n68) );
  NOR2BX4 U126 ( .AN(n50), .B(n120), .Y(n119) );
  XOR2X2 U127 ( .A(n31), .B(n73), .Y(SUM[4]) );
  AOI21X2 U128 ( .A0(n137), .A1(n127), .B0(n138), .Y(n136) );
  NAND2X2 U129 ( .A(n131), .B(n132), .Y(n124) );
  NAND2X2 U130 ( .A(B[10]), .B(A[10]), .Y(n155) );
  OAI21X2 U131 ( .A0(n109), .A1(n129), .B0(n107), .Y(n128) );
  NAND2X1 U132 ( .A(n75), .B(n85), .Y(n117) );
  NAND2BX4 U133 ( .AN(n74), .B(n75), .Y(n178) );
  NOR3X2 U134 ( .A(n1), .B(n25), .C(n130), .Y(n137) );
  INVX8 U135 ( .A(n156), .Y(n130) );
  XOR2X4 U136 ( .A(n67), .B(n68), .Y(SUM[6]) );
  AOI21X2 U137 ( .A0(n126), .A1(n127), .B0(n128), .Y(n125) );
  NOR2X2 U138 ( .A(n36), .B(n129), .Y(n126) );
  NOR2X4 U139 ( .A(n39), .B(n183), .Y(n77) );
  OAI2BB1X4 U140 ( .A0N(n88), .A1N(n89), .B0(n90), .Y(n83) );
  NAND2X2 U141 ( .A(n154), .B(n155), .Y(n153) );
  AOI2BB1X4 U142 ( .A0N(n150), .A1N(n152), .B0(n153), .Y(n148) );
  INVX4 U143 ( .A(n88), .Y(n92) );
  NAND2BX4 U144 ( .AN(n130), .B(n9), .Y(n115) );
  OR2X4 U145 ( .A(B[5]), .B(A[5]), .Y(n72) );
  NAND2X4 U146 ( .A(B[5]), .B(A[5]), .Y(n65) );
  NAND2X4 U147 ( .A(B[4]), .B(A[4]), .Y(n64) );
  OR2X4 U148 ( .A(B[2]), .B(A[2]), .Y(n84) );
  NAND2X1 U149 ( .A(n83), .B(n84), .Y(n82) );
  NOR2X2 U150 ( .A(n120), .B(n173), .Y(n172) );
  NAND2BX4 U151 ( .AN(n59), .B(n19), .Y(n49) );
  OR2X4 U152 ( .A(B[6]), .B(A[6]), .Y(n177) );
  XOR2X4 U153 ( .A(n94), .B(n95), .Y(SUM[16]) );
  XNOR2X2 U154 ( .A(n71), .B(n38), .Y(n187) );
  AND2X2 U155 ( .A(n35), .B(n176), .Y(n41) );
  NOR2XL U156 ( .A(n63), .B(n66), .Y(n35) );
  NAND2X4 U157 ( .A(n165), .B(n45), .Y(n162) );
  NAND2XL U158 ( .A(n30), .B(n47), .Y(n169) );
  NOR2X1 U159 ( .A(n113), .B(n114), .Y(n96) );
  AND2X2 U160 ( .A(n47), .B(n161), .Y(n42) );
  XOR2X4 U161 ( .A(n43), .B(n37), .Y(SUM[9]) );
  AND2X1 U162 ( .A(n72), .B(n65), .Y(n38) );
  NOR2BX4 U163 ( .AN(n78), .B(n77), .Y(n76) );
  NOR2BX1 U164 ( .AN(n64), .B(n66), .Y(n73) );
  OAI21X1 U165 ( .A0(n100), .A1(n101), .B0(n102), .Y(n99) );
  NAND2X4 U166 ( .A(B[6]), .B(A[6]), .Y(n59) );
  NAND2XL U167 ( .A(A[2]), .B(B[2]), .Y(n39) );
  NOR2BX1 U168 ( .AN(n93), .B(n40), .Y(SUM[0]) );
  NOR2XL U169 ( .A(A[0]), .B(B[0]), .Y(n40) );
  OAI21X2 U170 ( .A0(n96), .A1(n97), .B0(n98), .Y(n94) );
  INVX1 U171 ( .A(n99), .Y(n98) );
  OAI21X1 U172 ( .A0(n117), .A1(n179), .B0(n41), .Y(n116) );
  NOR2BX2 U173 ( .AN(n102), .B(n122), .Y(n121) );
  NAND2BXL U174 ( .AN(n108), .B(n103), .Y(n123) );
  XOR2X2 U175 ( .A(n83), .B(n86), .Y(SUM[2]) );
  XOR2X2 U176 ( .A(n89), .B(n91), .Y(SUM[1]) );
  NOR2XL U177 ( .A(n1), .B(n109), .Y(n105) );
  NAND2XL U178 ( .A(n103), .B(n104), .Y(n101) );
  NOR2X1 U179 ( .A(n105), .B(n106), .Y(n100) );
  INVX1 U180 ( .A(n93), .Y(n89) );
  XOR2X1 U181 ( .A(B[16]), .B(A[16]), .Y(n95) );
  NAND3BX4 U182 ( .AN(n74), .B(n76), .C(n75), .Y(n61) );
  AND2X1 U183 ( .A(B[8]), .B(A[8]), .Y(n151) );
  OR2X2 U184 ( .A(A[14]), .B(B[14]), .Y(n103) );
  NAND3XL U185 ( .A(n111), .B(n104), .C(n112), .Y(n97) );
  NAND2XL U186 ( .A(A[9]), .B(B[9]), .Y(n152) );
  OR2X2 U187 ( .A(A[1]), .B(B[1]), .Y(n88) );
  XOR2X4 U188 ( .A(n54), .B(n55), .Y(SUM[7]) );
  CLKINVX3 U189 ( .A(n104), .Y(n122) );
  OR2X4 U190 ( .A(A[15]), .B(B[15]), .Y(n104) );
  XOR2X4 U191 ( .A(n133), .B(n134), .Y(SUM[14]) );
  XOR2X4 U192 ( .A(n139), .B(n140), .Y(SUM[13]) );
  OAI2BB1X4 U193 ( .A0N(n147), .A1N(n46), .B0(n115), .Y(n146) );
  NAND2X4 U194 ( .A(n148), .B(n149), .Y(n127) );
  OR2X4 U195 ( .A(A[11]), .B(B[11]), .Y(n156) );
  XOR2X4 U196 ( .A(n166), .B(n167), .Y(n186) );
  OR2X4 U197 ( .A(A[8]), .B(B[8]), .Y(n47) );
  NAND2X4 U198 ( .A(n176), .B(n175), .Y(n51) );
  NOR2X4 U199 ( .A(n56), .B(n58), .Y(n176) );
  AOI21X4 U200 ( .A0(n65), .A1(n64), .B0(n63), .Y(n175) );
  OAI21X4 U201 ( .A0(n178), .A1(n179), .B0(n180), .Y(n52) );
  OR2X4 U202 ( .A(A[4]), .B(B[4]), .Y(n69) );
  NAND2X4 U203 ( .A(n184), .B(n185), .Y(n75) );
endmodule


module butterfly_DW01_sub_121 ( A, B, DIFF );
  input [16:0] A;
  input [16:0] B;
  output [16:0] DIFF;
  wire   n223, n224, n225, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222;

  NAND2X1 U3 ( .A(n133), .B(n186), .Y(n185) );
  AND2X4 U4 ( .A(n32), .B(n202), .Y(n1) );
  NAND2BX4 U5 ( .AN(A[7]), .B(B[7]), .Y(n218) );
  CLKINVX3 U6 ( .A(n164), .Y(n2) );
  CLKINVX3 U7 ( .A(n132), .Y(n164) );
  NAND2BX4 U8 ( .AN(A[13]), .B(B[13]), .Y(n130) );
  NAND3BX4 U9 ( .AN(n194), .B(n168), .C(n21), .Y(n188) );
  NAND2BX4 U10 ( .AN(n194), .B(n168), .Y(n3) );
  NAND4X4 U11 ( .A(n213), .B(n17), .C(n87), .D(n84), .Y(n28) );
  XOR2X2 U12 ( .A(n100), .B(n101), .Y(DIFF[3]) );
  AOI21X1 U13 ( .A0(n102), .A1(n103), .B0(n104), .Y(n101) );
  INVX8 U14 ( .A(B[11]), .Y(n67) );
  INVX8 U15 ( .A(n171), .Y(n194) );
  INVX3 U16 ( .A(n172), .Y(n34) );
  CLKINVX4 U17 ( .A(n28), .Y(n172) );
  CLKINVX3 U18 ( .A(n145), .Y(n41) );
  INVX1 U19 ( .A(A[10]), .Y(n14) );
  NAND3BX2 U20 ( .AN(n94), .B(n80), .C(n153), .Y(n17) );
  NAND2X2 U21 ( .A(n65), .B(n141), .Y(n11) );
  INVX4 U22 ( .A(n65), .Y(n199) );
  CLKINVX2 U23 ( .A(n70), .Y(n27) );
  NAND4X2 U24 ( .A(n45), .B(n170), .C(n168), .D(n38), .Y(n160) );
  NAND2X2 U25 ( .A(n49), .B(n50), .Y(n147) );
  INVX4 U26 ( .A(n18), .Y(n89) );
  NAND2BX2 U27 ( .AN(A[5]), .B(B[5]), .Y(n18) );
  INVX4 U28 ( .A(n86), .Y(n46) );
  INVX1 U29 ( .A(n87), .Y(n82) );
  INVXL U30 ( .A(n94), .Y(n99) );
  AND2X2 U31 ( .A(n181), .B(n76), .Y(n60) );
  XNOR2X1 U32 ( .A(n112), .B(n63), .Y(DIFF[1]) );
  NOR2BX1 U33 ( .AN(n90), .B(n89), .Y(n92) );
  NAND2BX1 U34 ( .AN(B[5]), .B(A[5]), .Y(n90) );
  XNOR2X4 U35 ( .A(n78), .B(n79), .Y(n4) );
  INVX4 U36 ( .A(n23), .Y(n52) );
  AND3X4 U37 ( .A(n177), .B(n203), .C(n77), .Y(n5) );
  NOR2X2 U38 ( .A(n183), .B(n136), .Y(n182) );
  NOR2X4 U39 ( .A(n48), .B(n166), .Y(n170) );
  NAND4X4 U40 ( .A(n213), .B(n214), .C(n84), .D(n87), .Y(n10) );
  NAND4X4 U41 ( .A(n128), .B(n7), .C(n21), .D(n47), .Y(n6) );
  INVX3 U42 ( .A(n199), .Y(n33) );
  BUFX8 U43 ( .A(n127), .Y(n7) );
  NOR2X4 U44 ( .A(n98), .B(n152), .Y(n202) );
  BUFX16 U45 ( .A(n130), .Y(n47) );
  XNOR2X4 U46 ( .A(n8), .B(n204), .Y(DIFF[11]) );
  NOR2X4 U47 ( .A(n51), .B(n52), .Y(n8) );
  NAND2BX4 U48 ( .AN(A[13]), .B(B[13]), .Y(n9) );
  INVX8 U49 ( .A(n20), .Y(n86) );
  INVX2 U50 ( .A(A[13]), .Y(n16) );
  NAND2BX4 U51 ( .AN(n48), .B(n38), .Y(n187) );
  INVX4 U52 ( .A(n141), .Y(n176) );
  NAND2BX4 U53 ( .AN(n11), .B(n38), .Y(n193) );
  INVX8 U54 ( .A(A[9]), .Y(n151) );
  NAND2BX2 U55 ( .AN(n199), .B(n38), .Y(n197) );
  BUFX1 U56 ( .A(n72), .Y(n12) );
  NOR2X4 U57 ( .A(n197), .B(n198), .Y(n196) );
  NOR2X2 U58 ( .A(n136), .B(n137), .Y(n121) );
  BUFX4 U59 ( .A(n144), .Y(n66) );
  INVX2 U60 ( .A(n203), .Y(n175) );
  NAND2BX4 U61 ( .AN(n149), .B(n181), .Y(n148) );
  BUFX12 U62 ( .A(A[8]), .Y(n13) );
  NAND2X4 U63 ( .A(n132), .B(n133), .Y(n131) );
  NAND2BX2 U64 ( .AN(A[7]), .B(B[7]), .Y(n83) );
  INVX1 U65 ( .A(n114), .Y(n110) );
  BUFX12 U66 ( .A(n141), .Y(n21) );
  AND3X1 U67 ( .A(n77), .B(n83), .C(n177), .Y(n25) );
  AND2X2 U68 ( .A(n24), .B(n128), .Y(n44) );
  CLKINVX4 U69 ( .A(n135), .Y(n140) );
  NAND3X4 U70 ( .A(n41), .B(n14), .C(n144), .Y(n171) );
  NAND2BX2 U71 ( .AN(B[15]), .B(A[15]), .Y(n126) );
  NAND3X2 U72 ( .A(n72), .B(n66), .C(n23), .Y(n149) );
  XNOR2X4 U73 ( .A(n189), .B(n15), .Y(DIFF[13]) );
  AND2X1 U74 ( .A(n47), .B(n133), .Y(n15) );
  OR2X4 U75 ( .A(B[13]), .B(n16), .Y(n133) );
  NAND2BX4 U76 ( .AN(A[6]), .B(B[6]), .Y(n80) );
  NAND4BBX4 U77 ( .AN(n152), .BN(n98), .C(n153), .D(n46), .Y(n137) );
  CLKINVX4 U78 ( .A(n218), .Y(n152) );
  INVX8 U79 ( .A(n96), .Y(n98) );
  OR2X1 U80 ( .A(n69), .B(n70), .Y(n29) );
  NAND2BXL U81 ( .AN(n74), .B(n10), .Y(n73) );
  OR2X2 U82 ( .A(n31), .B(n151), .Y(n50) );
  NAND2X4 U83 ( .A(n151), .B(B[9]), .Y(n177) );
  NAND2X4 U84 ( .A(n145), .B(A[10]), .Y(n23) );
  INVX4 U85 ( .A(B[10]), .Y(n145) );
  OAI21X2 U86 ( .A0(A[10]), .A1(n145), .B0(n65), .Y(n143) );
  CLKINVX8 U87 ( .A(n177), .Y(n70) );
  BUFX3 U88 ( .A(n225), .Y(DIFF[4]) );
  INVX4 U89 ( .A(A[7]), .Y(n215) );
  NAND2BX4 U90 ( .AN(A[6]), .B(B[6]), .Y(n20) );
  OR2X4 U91 ( .A(B[7]), .B(n215), .Y(n84) );
  INVX4 U92 ( .A(n200), .Y(n69) );
  NAND3XL U93 ( .A(n12), .B(n71), .C(n73), .Y(n68) );
  AND2X2 U94 ( .A(B[9]), .B(n151), .Y(n22) );
  NAND2BX4 U95 ( .AN(n166), .B(n128), .Y(n125) );
  NOR2X2 U96 ( .A(n52), .B(n69), .Y(n142) );
  BUFX8 U97 ( .A(n126), .Y(n24) );
  NAND3BX4 U98 ( .AN(n94), .B(n20), .C(n153), .Y(n214) );
  NAND4X4 U99 ( .A(n25), .B(n40), .C(n174), .D(n33), .Y(n173) );
  CLKINVX8 U100 ( .A(n69), .Y(n26) );
  NAND2X1 U101 ( .A(n203), .B(n23), .Y(n209) );
  XNOR2X4 U102 ( .A(n68), .B(n29), .Y(DIFF[9]) );
  AND2X2 U103 ( .A(n66), .B(n33), .Y(n204) );
  AND2X4 U104 ( .A(n1), .B(n61), .Y(n30) );
  NOR2X2 U105 ( .A(n89), .B(n86), .Y(n61) );
  DLY1X1 U106 ( .A(B[9]), .Y(n31) );
  BUFX8 U107 ( .A(n95), .Y(n32) );
  NAND2BX1 U108 ( .AN(n166), .B(n2), .Y(n39) );
  OAI21X4 U109 ( .A0(n124), .A1(n125), .B0(n24), .Y(n123) );
  NAND2BX4 U110 ( .AN(n176), .B(n47), .Y(n183) );
  NAND2X2 U111 ( .A(n28), .B(n83), .Y(n181) );
  NAND2BX4 U112 ( .AN(B[6]), .B(A[6]), .Y(n87) );
  NAND2XL U113 ( .A(n12), .B(n77), .Y(n75) );
  NAND2X4 U114 ( .A(n9), .B(n65), .Y(n48) );
  NAND2XL U115 ( .A(n83), .B(n84), .Y(n78) );
  NOR2X4 U116 ( .A(n6), .B(n134), .Y(n122) );
  NAND4X4 U117 ( .A(n128), .B(n7), .C(n21), .D(n47), .Y(n135) );
  INVX4 U118 ( .A(n91), .Y(n88) );
  NAND3X4 U119 ( .A(n22), .B(n144), .C(n146), .Y(n168) );
  NAND2X4 U120 ( .A(n209), .B(n57), .Y(n58) );
  NAND4X4 U121 ( .A(n144), .B(n146), .C(n200), .D(n72), .Y(n169) );
  OAI21X4 U122 ( .A0(n142), .A1(n143), .B0(n66), .Y(n139) );
  AOI21X2 U123 ( .A0(n27), .A1(n206), .B0(n211), .Y(n210) );
  CLKINVX3 U124 ( .A(n9), .Y(n167) );
  OAI2BB1X4 U125 ( .A0N(n215), .A1N(B[7]), .B0(n77), .Y(n74) );
  NOR2X4 U126 ( .A(n34), .B(n30), .Y(n35) );
  NOR2X4 U127 ( .A(n173), .B(n35), .Y(n158) );
  NAND2X2 U128 ( .A(n129), .B(n47), .Y(n186) );
  INVX4 U129 ( .A(n165), .Y(n129) );
  NAND2X1 U130 ( .A(n26), .B(n208), .Y(n211) );
  XNOR2X4 U131 ( .A(n195), .B(n36), .Y(DIFF[12]) );
  AND2X1 U132 ( .A(n21), .B(n165), .Y(n36) );
  NOR2X4 U133 ( .A(n205), .B(n175), .Y(n51) );
  OR2X4 U134 ( .A(n150), .B(n137), .Y(n49) );
  AOI21X4 U135 ( .A0(n129), .A1(n47), .B0(n131), .Y(n124) );
  AOI21X4 U136 ( .A0(n162), .A1(n163), .B0(n164), .Y(n161) );
  CLKINVX8 U137 ( .A(n169), .Y(n37) );
  INVX8 U138 ( .A(n37), .Y(n38) );
  NOR2X2 U139 ( .A(n166), .B(n167), .Y(n162) );
  NOR2X4 U140 ( .A(n175), .B(n176), .Y(n174) );
  XNOR2X4 U141 ( .A(n178), .B(n39), .Y(DIFF[14]) );
  NOR2X4 U142 ( .A(n166), .B(n167), .Y(n40) );
  OAI21X2 U143 ( .A0(n109), .A1(n110), .B0(n111), .Y(n103) );
  NOR2X4 U144 ( .A(n74), .B(n70), .Y(n212) );
  XNOR2X4 U145 ( .A(n117), .B(n42), .Y(n223) );
  XOR2X4 U146 ( .A(B[16]), .B(A[16]), .Y(n42) );
  NAND2X4 U147 ( .A(n67), .B(A[11]), .Y(n144) );
  NOR2X4 U148 ( .A(n188), .B(n187), .Y(n184) );
  INVX8 U149 ( .A(n127), .Y(n166) );
  AOI21X4 U150 ( .A0(n121), .A1(n122), .B0(n123), .Y(n120) );
  NOR2X2 U151 ( .A(n194), .B(n176), .Y(n45) );
  NAND3X4 U152 ( .A(n217), .B(n32), .C(n216), .Y(n71) );
  NOR2X4 U153 ( .A(n89), .B(n86), .Y(n216) );
  NAND2BX4 U154 ( .AN(n194), .B(n168), .Y(n198) );
  NAND2X4 U155 ( .A(n93), .B(n94), .Y(n91) );
  NAND2X4 U156 ( .A(n95), .B(n96), .Y(n93) );
  BUFX20 U157 ( .A(n223), .Y(DIFF[16]) );
  NOR2BX4 U158 ( .AN(B[8]), .B(n13), .Y(n219) );
  NOR3BX4 U159 ( .AN(n218), .B(n98), .C(n219), .Y(n217) );
  NAND2BX4 U160 ( .AN(B[9]), .B(A[9]), .Y(n200) );
  XNOR2X4 U161 ( .A(n157), .B(n44), .Y(DIFF[15]) );
  NAND2X4 U162 ( .A(n208), .B(n26), .Y(n207) );
  NOR2X4 U163 ( .A(n147), .B(n148), .Y(n118) );
  NOR2X1 U164 ( .A(n98), .B(n99), .Y(n97) );
  AOI21X4 U165 ( .A0(n206), .A1(n27), .B0(n207), .Y(n205) );
  AOI21X4 U166 ( .A0(n46), .A1(n81), .B0(n82), .Y(n79) );
  NOR2X2 U167 ( .A(n136), .B(n176), .Y(n190) );
  NAND2BX4 U168 ( .AN(A[2]), .B(B[2]), .Y(n102) );
  NAND2BX4 U169 ( .AN(B[3]), .B(A[3]), .Y(n106) );
  NAND3X2 U170 ( .A(n221), .B(n111), .C(n108), .Y(n220) );
  OAI21X4 U171 ( .A0(n3), .A1(n193), .B0(n165), .Y(n192) );
  NAND2X4 U172 ( .A(n10), .B(n212), .Y(n208) );
  NAND2X4 U173 ( .A(n64), .B(n220), .Y(n156) );
  OAI21X4 U174 ( .A0(n138), .A1(n139), .B0(n140), .Y(n119) );
  NAND2X4 U175 ( .A(n160), .B(n161), .Y(n159) );
  NAND2X2 U176 ( .A(n133), .B(n165), .Y(n163) );
  INVX4 U177 ( .A(n136), .Y(n138) );
  NAND3BX4 U178 ( .AN(B[5]), .B(A[5]), .C(n80), .Y(n213) );
  AOI21X4 U179 ( .A0(n190), .A1(n191), .B0(n192), .Y(n189) );
  NOR2X1 U180 ( .A(n154), .B(n155), .Y(n150) );
  NAND2X4 U181 ( .A(n1), .B(n61), .Y(n76) );
  OAI2BB1X4 U182 ( .A0N(n181), .A1N(n76), .B0(n182), .Y(n180) );
  CLKINVX4 U183 ( .A(n224), .Y(n53) );
  INVX8 U184 ( .A(n53), .Y(DIFF[5]) );
  NAND2X4 U185 ( .A(n222), .B(n114), .Y(n221) );
  NAND4X2 U186 ( .A(n102), .B(n114), .C(n105), .D(n116), .Y(n134) );
  NAND2BX4 U187 ( .AN(A[1]), .B(B[1]), .Y(n114) );
  XOR2X2 U188 ( .A(n81), .B(n85), .Y(DIFF[6]) );
  OAI21X4 U189 ( .A0(n88), .A1(n89), .B0(n90), .Y(n81) );
  OAI21X4 U190 ( .A0(n201), .A1(n172), .B0(n76), .Y(n191) );
  INVX2 U191 ( .A(n83), .Y(n201) );
  INVX8 U192 ( .A(n4), .Y(DIFF[7]) );
  NAND2BX4 U193 ( .AN(A[8]), .B(B[8]), .Y(n77) );
  NAND2X2 U194 ( .A(n56), .B(n210), .Y(n59) );
  NAND2X4 U195 ( .A(n58), .B(n59), .Y(DIFF[10]) );
  INVXL U196 ( .A(n209), .Y(n56) );
  INVX4 U197 ( .A(n210), .Y(n57) );
  NAND2BX4 U198 ( .AN(B[1]), .B(A[1]), .Y(n111) );
  NAND2X4 U199 ( .A(n5), .B(n65), .Y(n136) );
  OR2XL U200 ( .A(n104), .B(n107), .Y(n62) );
  XNOR2X1 U201 ( .A(n103), .B(n62), .Y(DIFF[2]) );
  OR2XL U202 ( .A(n113), .B(n110), .Y(n63) );
  XOR2X4 U203 ( .A(n75), .B(n60), .Y(DIFF[8]) );
  NAND2X4 U204 ( .A(n71), .B(n72), .Y(n206) );
  NAND3X4 U205 ( .A(n134), .B(n106), .C(n156), .Y(n95) );
  NAND2BX2 U206 ( .AN(B[2]), .B(A[2]), .Y(n108) );
  AND2X2 U207 ( .A(n102), .B(n105), .Y(n64) );
  NAND2BX4 U208 ( .AN(B[4]), .B(A[4]), .Y(n94) );
  OR2X4 U209 ( .A(n67), .B(A[11]), .Y(n65) );
  NAND2XL U210 ( .A(n105), .B(n106), .Y(n100) );
  INVXL U211 ( .A(n106), .Y(n154) );
  NAND2BXL U212 ( .AN(n116), .B(n115), .Y(n112) );
  NAND2XL U213 ( .A(n115), .B(n116), .Y(DIFF[0]) );
  NOR2X1 U214 ( .A(n82), .B(n86), .Y(n85) );
  XOR2X1 U215 ( .A(n32), .B(n97), .Y(n225) );
  INVX1 U216 ( .A(n102), .Y(n107) );
  INVX1 U217 ( .A(n111), .Y(n113) );
  XOR2X1 U218 ( .A(n91), .B(n92), .Y(n224) );
  INVX1 U219 ( .A(n112), .Y(n109) );
  INVX1 U220 ( .A(n108), .Y(n104) );
  INVX1 U221 ( .A(n156), .Y(n155) );
  INVX1 U222 ( .A(n115), .Y(n222) );
  NAND2BX1 U223 ( .AN(A[0]), .B(B[0]), .Y(n116) );
  NAND2BX1 U224 ( .AN(B[0]), .B(A[0]), .Y(n115) );
  AOI21X4 U225 ( .A0(n138), .A1(n191), .B0(n196), .Y(n195) );
  OAI21X4 U226 ( .A0(n118), .A1(n119), .B0(n120), .Y(n117) );
  NOR2X4 U227 ( .A(n159), .B(n158), .Y(n157) );
  NAND2BX4 U228 ( .AN(A[15]), .B(B[15]), .Y(n128) );
  NAND2BX4 U229 ( .AN(B[14]), .B(A[14]), .Y(n132) );
  NAND2BX4 U230 ( .AN(A[14]), .B(B[14]), .Y(n127) );
  NAND2X4 U231 ( .A(n179), .B(n180), .Y(n178) );
  NOR2X4 U232 ( .A(n184), .B(n185), .Y(n179) );
  NAND2BX4 U233 ( .AN(B[12]), .B(A[12]), .Y(n165) );
  NAND2BX4 U234 ( .AN(A[12]), .B(B[12]), .Y(n141) );
  NAND2BX4 U235 ( .AN(B[8]), .B(n13), .Y(n72) );
  NAND2BX4 U236 ( .AN(A[4]), .B(B[4]), .Y(n96) );
  NAND2BX4 U237 ( .AN(A[3]), .B(B[3]), .Y(n105) );
  NAND2BX4 U238 ( .AN(A[5]), .B(B[5]), .Y(n153) );
  NAND2BX4 U239 ( .AN(B[10]), .B(A[10]), .Y(n146) );
  NAND2BX4 U240 ( .AN(A[10]), .B(B[10]), .Y(n203) );
endmodule


module butterfly_DW01_sub_123 ( A, B, DIFF );
  input [16:0] A;
  input [16:0] B;
  output [16:0] DIFF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187;

  INVX2 U3 ( .A(n30), .Y(n1) );
  BUFX16 U4 ( .A(n43), .Y(n30) );
  BUFX20 U5 ( .A(n68), .Y(n32) );
  INVX4 U6 ( .A(n23), .Y(n24) );
  INVX3 U7 ( .A(n42), .Y(n23) );
  BUFX3 U8 ( .A(n105), .Y(n28) );
  OAI2BB1X2 U9 ( .A0N(n105), .A1N(n144), .B0(n110), .Y(n131) );
  NAND2BX4 U10 ( .AN(A[1]), .B(B[1]), .Y(n87) );
  NAND2BX4 U11 ( .AN(B[1]), .B(A[1]), .Y(n120) );
  NAND2BX4 U12 ( .AN(A[9]), .B(B[9]), .Y(n164) );
  INVX8 U13 ( .A(n161), .Y(n7) );
  AOI21X2 U14 ( .A0(n1), .A1(n24), .B0(n177), .Y(n176) );
  NOR2X4 U15 ( .A(n64), .B(n177), .Y(n63) );
  AND4X4 U16 ( .A(n33), .B(n37), .C(n7), .D(n69), .Y(n11) );
  NOR2BX4 U17 ( .AN(B[11]), .B(A[11]), .Y(n157) );
  NAND2BX4 U18 ( .AN(B[7]), .B(A[7]), .Y(n174) );
  AND2X4 U19 ( .A(n72), .B(n32), .Y(n25) );
  NAND3X4 U20 ( .A(n67), .B(n66), .C(n72), .Y(n62) );
  AND2X2 U21 ( .A(n175), .B(n174), .Y(n173) );
  NOR2X2 U22 ( .A(n104), .B(n136), .Y(n17) );
  INVX1 U23 ( .A(n111), .Y(n144) );
  INVX4 U24 ( .A(n60), .Y(n19) );
  NOR2X1 U25 ( .A(n103), .B(n29), .Y(n99) );
  NAND2X1 U26 ( .A(n110), .B(n111), .Y(n109) );
  BUFX8 U27 ( .A(n158), .Y(n41) );
  CLKINVX3 U28 ( .A(n121), .Y(n79) );
  NAND3BX2 U29 ( .AN(n107), .B(n151), .C(n152), .Y(n34) );
  NAND2X2 U30 ( .A(n17), .B(n153), .Y(n152) );
  INVX1 U31 ( .A(n164), .Y(n46) );
  AND2X2 U32 ( .A(n39), .B(n69), .Y(n74) );
  BUFX4 U33 ( .A(n37), .Y(n4) );
  NOR2BX2 U34 ( .AN(n120), .B(n84), .Y(n86) );
  AOI21X2 U35 ( .A0(n92), .A1(n93), .B0(n94), .Y(n90) );
  INVX4 U36 ( .A(n73), .Y(n71) );
  NAND2BX2 U37 ( .AN(A[15]), .B(B[15]), .Y(n106) );
  CLKINVX3 U38 ( .A(n61), .Y(n64) );
  CLKINVX3 U39 ( .A(n80), .Y(n2) );
  CLKINVX3 U40 ( .A(n2), .Y(n3) );
  NAND2BX4 U41 ( .AN(n87), .B(n121), .Y(n187) );
  AOI21X2 U42 ( .A0(n107), .A1(n108), .B0(n144), .Y(n143) );
  AND2X1 U43 ( .A(n108), .B(n111), .Y(n35) );
  INVX4 U44 ( .A(n108), .Y(n150) );
  AOI21X4 U45 ( .A0(n71), .A1(n176), .B0(n64), .Y(n172) );
  NAND3X1 U46 ( .A(n108), .B(n19), .C(n105), .Y(n137) );
  INVX8 U47 ( .A(A[8]), .Y(n6) );
  NAND2X4 U48 ( .A(n77), .B(n80), .Y(n185) );
  NAND2X4 U49 ( .A(n5), .B(n163), .Y(n21) );
  INVX2 U50 ( .A(n162), .Y(n5) );
  NAND2X4 U51 ( .A(n6), .B(B[8]), .Y(n56) );
  NAND2X4 U52 ( .A(n116), .B(n20), .Y(n161) );
  INVX4 U53 ( .A(n134), .Y(n142) );
  INVX2 U54 ( .A(n148), .Y(n29) );
  INVX1 U55 ( .A(n47), .Y(n45) );
  XNOR2X4 U56 ( .A(n8), .B(n138), .Y(DIFF[14]) );
  AND2X1 U57 ( .A(n28), .B(n110), .Y(n8) );
  CLKINVX4 U58 ( .A(n115), .Y(n9) );
  INVX3 U59 ( .A(n146), .Y(n115) );
  NAND2BX2 U60 ( .AN(B[3]), .B(A[3]), .Y(n81) );
  BUFX20 U61 ( .A(B[5]), .Y(n42) );
  NOR2XL U62 ( .A(n101), .B(n102), .Y(n100) );
  NAND2BX4 U63 ( .AN(A[6]), .B(B[6]), .Y(n10) );
  AOI21X1 U64 ( .A0(n114), .A1(n3), .B0(n115), .Y(n112) );
  INVX8 U65 ( .A(n52), .Y(n181) );
  NAND3BX4 U66 ( .AN(n179), .B(n50), .C(n49), .Y(n13) );
  INVXL U67 ( .A(A[7]), .Y(n59) );
  XNOR2X4 U68 ( .A(n168), .B(n12), .Y(DIFF[11]) );
  NAND2XL U69 ( .A(n133), .B(n166), .Y(n12) );
  OAI21XL U70 ( .A0(n29), .A1(n112), .B0(n113), .Y(n93) );
  XOR2X4 U71 ( .A(n13), .B(n14), .Y(DIFF[9]) );
  NOR2X2 U72 ( .A(n45), .B(n46), .Y(n14) );
  XOR2X4 U73 ( .A(n4), .B(n74), .Y(DIFF[4]) );
  XNOR2X4 U74 ( .A(n36), .B(n15), .Y(DIFF[10]) );
  NAND2XL U75 ( .A(n41), .B(n167), .Y(n15) );
  XNOR2X4 U76 ( .A(n78), .B(n16), .Y(DIFF[2]) );
  OR2X4 U77 ( .A(n79), .B(n82), .Y(n16) );
  XNOR2X4 U78 ( .A(n154), .B(n18), .Y(DIFF[12]) );
  AND2X1 U79 ( .A(n122), .B(n145), .Y(n18) );
  BUFX3 U80 ( .A(n133), .Y(n22) );
  NAND2X4 U81 ( .A(n129), .B(n130), .Y(n128) );
  NAND2BX4 U82 ( .AN(B[6]), .B(A[6]), .Y(n61) );
  AOI21X4 U83 ( .A0(n172), .A1(n173), .B0(n51), .Y(n171) );
  INVX4 U84 ( .A(n116), .Y(n60) );
  NAND2X4 U85 ( .A(n44), .B(n42), .Y(n68) );
  NAND2BX4 U86 ( .AN(B[2]), .B(A[2]), .Y(n121) );
  AOI2BB1X2 U87 ( .A0N(B[7]), .A1N(n59), .B0(n60), .Y(n58) );
  NAND2BX2 U88 ( .AN(A[10]), .B(B[10]), .Y(n158) );
  NAND3BX4 U89 ( .AN(n73), .B(n10), .C(n183), .Y(n182) );
  OAI2BB1X2 U90 ( .A0N(n69), .A1N(n70), .B0(n39), .Y(n38) );
  INVX4 U91 ( .A(n55), .Y(n26) );
  INVX8 U92 ( .A(n177), .Y(n20) );
  INVX8 U93 ( .A(n65), .Y(n177) );
  INVX4 U94 ( .A(n71), .Y(n39) );
  CLKINVX8 U95 ( .A(n104), .Y(n148) );
  NAND2X4 U96 ( .A(n166), .B(n167), .Y(n162) );
  AOI21X4 U97 ( .A0(n9), .A1(n27), .B0(n147), .Y(n139) );
  NAND2BX4 U98 ( .AN(B[4]), .B(A[4]), .Y(n73) );
  NAND2X2 U99 ( .A(n97), .B(n106), .Y(n124) );
  NAND3X2 U100 ( .A(n21), .B(n122), .C(n22), .Y(n151) );
  NAND3X2 U101 ( .A(n21), .B(n22), .C(n135), .Y(n129) );
  NAND2X4 U102 ( .A(n47), .B(n49), .Y(n165) );
  NAND2XL U103 ( .A(n41), .B(n164), .Y(n169) );
  XOR2X4 U104 ( .A(n25), .B(n38), .Y(DIFF[5]) );
  NAND2X2 U105 ( .A(n55), .B(n146), .Y(n54) );
  INVX8 U106 ( .A(n26), .Y(n27) );
  INVX8 U107 ( .A(n48), .Y(n179) );
  NAND2BX4 U108 ( .AN(B[11]), .B(A[11]), .Y(n166) );
  NOR3X4 U109 ( .A(n11), .B(n171), .C(n165), .Y(n170) );
  NOR2X4 U110 ( .A(n136), .B(n132), .Y(n135) );
  NOR2X1 U111 ( .A(n136), .B(n104), .Y(n127) );
  NAND2BX4 U112 ( .AN(B[13]), .B(A[13]), .Y(n111) );
  OAI21X4 U113 ( .A0(n141), .A1(n142), .B0(n143), .Y(n140) );
  AOI21X4 U114 ( .A0(n31), .A1(n27), .B0(n156), .Y(n155) );
  NAND2BX2 U115 ( .AN(B[14]), .B(A[14]), .Y(n110) );
  INVX8 U116 ( .A(n145), .Y(n107) );
  OAI21X4 U117 ( .A0(n83), .A1(n84), .B0(n120), .Y(n78) );
  NAND2X2 U118 ( .A(n146), .B(n55), .Y(n153) );
  NAND3X1 U119 ( .A(n122), .B(n108), .C(n133), .Y(n141) );
  NAND2X4 U120 ( .A(n108), .B(n105), .Y(n132) );
  NAND2BX4 U121 ( .AN(B[10]), .B(A[10]), .Y(n167) );
  NAND2BX4 U122 ( .AN(A[3]), .B(B[3]), .Y(n80) );
  NOR2X2 U123 ( .A(n150), .B(n136), .Y(n149) );
  NAND2BX4 U124 ( .AN(B[9]), .B(A[9]), .Y(n47) );
  INVX2 U125 ( .A(n40), .Y(n31) );
  NAND4X4 U126 ( .A(n33), .B(n37), .C(n7), .D(n69), .Y(n48) );
  AND2X4 U127 ( .A(n32), .B(n56), .Y(n33) );
  OAI2BB1X4 U128 ( .A0N(n20), .A1N(n62), .B0(n61), .Y(n57) );
  AOI21X4 U129 ( .A0(n123), .A1(n107), .B0(n131), .Y(n130) );
  NAND2BX2 U130 ( .AN(n42), .B(n30), .Y(n72) );
  INVX4 U131 ( .A(n132), .Y(n123) );
  NAND4BX2 U132 ( .AN(n60), .B(n20), .C(n69), .D(n32), .Y(n102) );
  AOI21X2 U133 ( .A0(n117), .A1(n118), .B0(n102), .Y(n114) );
  XOR2X4 U134 ( .A(n34), .B(n35), .Y(DIFF[13]) );
  AOI21X2 U135 ( .A0(n31), .A1(n27), .B0(n137), .Y(n126) );
  BUFX8 U136 ( .A(n70), .Y(n37) );
  NAND3BX4 U137 ( .AN(n42), .B(n10), .C(n30), .Y(n175) );
  NAND3X2 U138 ( .A(n121), .B(n88), .C(n120), .Y(n186) );
  XOR2X2 U139 ( .A(n85), .B(n86), .Y(DIFF[1]) );
  NAND2X4 U140 ( .A(n56), .B(n116), .Y(n51) );
  INVX8 U141 ( .A(A[5]), .Y(n44) );
  NAND2X4 U142 ( .A(n178), .B(n47), .Y(n36) );
  NAND2X2 U143 ( .A(n148), .B(n19), .Y(n156) );
  XOR2X2 U144 ( .A(n75), .B(n76), .Y(DIFF[3]) );
  AOI21X2 U145 ( .A0(n77), .A1(n78), .B0(n79), .Y(n76) );
  NAND2X2 U146 ( .A(n148), .B(n149), .Y(n147) );
  INVX8 U147 ( .A(n122), .Y(n136) );
  NAND3X4 U148 ( .A(n164), .B(n165), .C(n41), .Y(n163) );
  NAND4X2 U149 ( .A(n77), .B(n80), .C(n89), .D(n87), .Y(n101) );
  NAND2BX1 U150 ( .AN(B[15]), .B(A[15]), .Y(n97) );
  INVX8 U151 ( .A(n181), .Y(n40) );
  NAND2X4 U152 ( .A(n71), .B(n32), .Y(n66) );
  NAND3X4 U153 ( .A(n32), .B(n70), .C(n69), .Y(n67) );
  NAND2BX4 U154 ( .AN(A[2]), .B(B[2]), .Y(n77) );
  INVX8 U155 ( .A(n44), .Y(n43) );
  NAND2BX2 U156 ( .AN(B[12]), .B(A[12]), .Y(n145) );
  OAI21X4 U157 ( .A0(n180), .A1(n179), .B0(n164), .Y(n178) );
  OAI21X4 U158 ( .A0(n51), .A1(n181), .B0(n49), .Y(n180) );
  NOR2X4 U159 ( .A(n139), .B(n140), .Y(n138) );
  NAND2BX4 U160 ( .AN(n51), .B(n40), .Y(n50) );
  NAND2X2 U161 ( .A(n22), .B(n134), .Y(n113) );
  NAND2BX2 U162 ( .AN(A[11]), .B(B[11]), .Y(n133) );
  NAND2X4 U163 ( .A(n69), .B(n32), .Y(n160) );
  NAND2BX4 U164 ( .AN(A[13]), .B(B[13]), .Y(n108) );
  XNOR2X4 U165 ( .A(n54), .B(n53), .Y(DIFF[8]) );
  NAND3BX4 U166 ( .AN(n185), .B(n186), .C(n187), .Y(n184) );
  XOR2X4 U167 ( .A(n125), .B(n124), .Y(DIFF[15]) );
  AOI21X4 U168 ( .A0(n127), .A1(n126), .B0(n128), .Y(n125) );
  NAND4X4 U169 ( .A(n182), .B(n175), .C(n174), .D(n61), .Y(n52) );
  XOR2X4 U170 ( .A(n90), .B(n91), .Y(DIFF[16]) );
  OAI211X2 U171 ( .A0(n95), .A1(n96), .B0(n97), .C0(n98), .Y(n94) );
  NAND2X2 U172 ( .A(n99), .B(n100), .Y(n98) );
  NAND2BX4 U173 ( .AN(B[8]), .B(A[8]), .Y(n49) );
  NAND3X2 U174 ( .A(n106), .B(n122), .C(n123), .Y(n103) );
  NAND2X4 U175 ( .A(n19), .B(n52), .Y(n146) );
  NAND4BX4 U176 ( .AN(n157), .B(n41), .C(n164), .D(n56), .Y(n104) );
  NAND2BX4 U177 ( .AN(A[4]), .B(B[4]), .Y(n69) );
  INVX4 U178 ( .A(n87), .Y(n84) );
  AOI21XL U179 ( .A0(n107), .A1(n108), .B0(n109), .Y(n95) );
  NAND3XL U180 ( .A(n77), .B(n87), .C(n119), .Y(n118) );
  NAND2XL U181 ( .A(n28), .B(n106), .Y(n96) );
  NAND2XL U182 ( .A(n49), .B(n56), .Y(n53) );
  INVX1 U183 ( .A(n77), .Y(n82) );
  NOR2BXL U184 ( .AN(n81), .B(n79), .Y(n117) );
  INVX1 U185 ( .A(n85), .Y(n83) );
  XOR2X1 U186 ( .A(B[16]), .B(A[16]), .Y(n91) );
  INVXL U187 ( .A(n103), .Y(n92) );
  NAND2XL U188 ( .A(n88), .B(n120), .Y(n119) );
  NAND2X1 U189 ( .A(n88), .B(n89), .Y(DIFF[0]) );
  NAND2BX1 U190 ( .AN(n89), .B(n88), .Y(n85) );
  NAND2BX1 U191 ( .AN(B[0]), .B(A[0]), .Y(n88) );
  NAND2BX1 U192 ( .AN(A[0]), .B(B[0]), .Y(n89) );
  NAND2XL U193 ( .A(n3), .B(n81), .Y(n75) );
  XOR2X4 U194 ( .A(n57), .B(n58), .Y(DIFF[7]) );
  XOR2X4 U195 ( .A(n62), .B(n63), .Y(DIFF[6]) );
  NAND2BX4 U196 ( .AN(A[14]), .B(B[14]), .Y(n105) );
  NOR2BX4 U197 ( .AN(n113), .B(n155), .Y(n154) );
  NAND2X4 U198 ( .A(n37), .B(n159), .Y(n55) );
  NOR2X4 U199 ( .A(n160), .B(n161), .Y(n159) );
  NAND2BX4 U200 ( .AN(n162), .B(n163), .Y(n134) );
  NAND2BX4 U201 ( .AN(A[12]), .B(B[12]), .Y(n122) );
  OAI21X4 U202 ( .A0(n170), .A1(n169), .B0(n167), .Y(n168) );
  NAND2BX4 U203 ( .AN(n43), .B(n42), .Y(n183) );
  NAND3X4 U204 ( .A(n101), .B(n184), .C(n81), .Y(n70) );
  NAND2BX4 U205 ( .AN(A[6]), .B(B[6]), .Y(n65) );
  NAND2BX4 U206 ( .AN(A[7]), .B(B[7]), .Y(n116) );
endmodule


module butterfly_DW01_add_184 ( A, B, SUM );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  wire   n221, n222, n223, n224, n225, n226, n227, n228, n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n70, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220;

  BUFX8 U2 ( .A(n112), .Y(n23) );
  NAND2X2 U3 ( .A(n41), .B(n30), .Y(n1) );
  INVX2 U4 ( .A(n88), .Y(n166) );
  NAND3BXL U5 ( .AN(n26), .B(n88), .C(n89), .Y(n183) );
  NAND3BX2 U6 ( .AN(n60), .B(B[6]), .C(n88), .Y(n165) );
  NOR2X2 U7 ( .A(n40), .B(n93), .Y(n91) );
  INVX4 U8 ( .A(n40), .Y(n39) );
  NAND2X4 U9 ( .A(n50), .B(n107), .Y(n120) );
  XOR2X4 U10 ( .A(n50), .B(n122), .Y(n70) );
  OAI2BB1X2 U11 ( .A0N(n130), .A1N(n129), .B0(n9), .Y(n2) );
  OAI2BB1X2 U12 ( .A0N(n130), .A1N(n129), .B0(n9), .Y(n127) );
  BUFX8 U13 ( .A(n131), .Y(n9) );
  NOR2BX1 U14 ( .AN(n197), .B(n209), .Y(n204) );
  CLKINVX4 U15 ( .A(n111), .Y(n93) );
  NAND2X1 U16 ( .A(B[1]), .B(A[1]), .Y(n131) );
  AND2X2 U17 ( .A(A[1]), .B(B[1]), .Y(n217) );
  NAND2X1 U18 ( .A(n76), .B(n34), .Y(n75) );
  NAND2X4 U19 ( .A(n45), .B(n47), .Y(n117) );
  NAND2X4 U20 ( .A(n41), .B(n30), .Y(n17) );
  BUFX2 U21 ( .A(B[2]), .Y(n57) );
  NAND2X4 U22 ( .A(n90), .B(n108), .Y(n213) );
  INVXL U23 ( .A(n94), .Y(n3) );
  INVX2 U24 ( .A(n3), .Y(n4) );
  NOR2X4 U25 ( .A(n26), .B(n166), .Y(n214) );
  INVXL U26 ( .A(B[6]), .Y(n5) );
  INVX1 U27 ( .A(n5), .Y(n6) );
  NOR2X4 U28 ( .A(n133), .B(n134), .Y(n7) );
  NOR2BX2 U29 ( .AN(n80), .B(n79), .Y(n97) );
  INVX2 U30 ( .A(A[4]), .Y(n27) );
  NAND2X2 U31 ( .A(n159), .B(n158), .Y(n192) );
  INVX4 U32 ( .A(n107), .Y(n105) );
  INVX2 U33 ( .A(n72), .Y(n73) );
  NAND2X1 U34 ( .A(n59), .B(B[2]), .Y(n125) );
  NAND3X4 U35 ( .A(n94), .B(n58), .C(n47), .Y(n121) );
  OAI2BB1X4 U36 ( .A0N(n173), .A1N(n176), .B0(n148), .Y(n174) );
  CLKINVX1 U37 ( .A(n125), .Y(n51) );
  NAND2X2 U38 ( .A(n6), .B(n56), .Y(n102) );
  CLKINVX3 U39 ( .A(n92), .Y(n40) );
  INVX12 U40 ( .A(B[4]), .Y(n41) );
  NOR2BX4 U41 ( .AN(n182), .B(n190), .Y(n188) );
  NAND2X2 U42 ( .A(n34), .B(n198), .Y(n209) );
  INVX4 U43 ( .A(n61), .Y(n34) );
  BUFX4 U44 ( .A(n99), .Y(n8) );
  BUFX20 U45 ( .A(n221), .Y(SUM[15]) );
  NAND2XL U46 ( .A(A[8]), .B(B[8]), .Y(n62) );
  BUFX4 U47 ( .A(n164), .Y(n29) );
  NOR2BX1 U48 ( .AN(n148), .B(n146), .Y(n177) );
  NOR2BX2 U49 ( .AN(n159), .B(n203), .Y(n202) );
  NAND2X2 U50 ( .A(n196), .B(n197), .Y(n190) );
  NOR2X2 U51 ( .A(n61), .B(n62), .Y(n199) );
  NAND2X2 U52 ( .A(A[9]), .B(B[9]), .Y(n76) );
  INVX1 U53 ( .A(n209), .Y(n212) );
  INVX1 U54 ( .A(n38), .Y(n207) );
  INVX4 U55 ( .A(n154), .Y(n35) );
  NAND2X1 U56 ( .A(B[8]), .B(A[8]), .Y(n80) );
  NAND2X1 U57 ( .A(B[12]), .B(A[12]), .Y(n147) );
  NAND2X1 U58 ( .A(B[13]), .B(A[13]), .Y(n148) );
  NAND2BX2 U59 ( .AN(n190), .B(n189), .Y(n158) );
  AOI21XL U60 ( .A0(n163), .A1(n162), .B0(n29), .Y(n161) );
  INVX1 U61 ( .A(n27), .Y(n28) );
  INVX2 U62 ( .A(n143), .Y(n153) );
  NOR2X1 U63 ( .A(A[15]), .B(B[15]), .Y(n64) );
  NAND2XL U64 ( .A(B[7]), .B(A[7]), .Y(n99) );
  INVX1 U65 ( .A(n60), .Y(n56) );
  NAND4BX2 U66 ( .AN(n164), .B(n195), .C(n84), .D(n80), .Y(n205) );
  INVX20 U67 ( .A(n70), .Y(SUM[4]) );
  AND2X1 U68 ( .A(n8), .B(n43), .Y(n10) );
  AND2X2 U69 ( .A(n147), .B(n35), .Y(n11) );
  BUFX20 U70 ( .A(n227), .Y(SUM[6]) );
  NAND3X1 U71 ( .A(n13), .B(n4), .C(n47), .Y(n20) );
  CLKINVX3 U72 ( .A(n12), .Y(n13) );
  NOR2BX2 U73 ( .AN(n200), .B(n207), .Y(n211) );
  AOI2BB1X2 U74 ( .A0N(n207), .A1N(n76), .B0(n208), .Y(n206) );
  CLKINVX2 U75 ( .A(n58), .Y(n12) );
  BUFX8 U76 ( .A(A[2]), .Y(n59) );
  AND2X2 U77 ( .A(n178), .B(n179), .Y(n14) );
  CLKINVX3 U78 ( .A(n195), .Y(n32) );
  INVX2 U79 ( .A(n93), .Y(n24) );
  NOR2X4 U80 ( .A(n185), .B(n15), .Y(n178) );
  AND3X4 U81 ( .A(n49), .B(n35), .C(n155), .Y(n15) );
  XOR2X4 U82 ( .A(n201), .B(n202), .Y(n224) );
  NAND2X2 U83 ( .A(n90), .B(n23), .Y(n122) );
  INVX3 U84 ( .A(n89), .Y(n31) );
  XNOR2X4 U85 ( .A(n36), .B(n2), .Y(n16) );
  INVX8 U86 ( .A(n16), .Y(SUM[2]) );
  AND2X2 U87 ( .A(n124), .B(n95), .Y(n54) );
  NAND2X1 U88 ( .A(n89), .B(n90), .Y(n85) );
  BUFX20 U89 ( .A(n106), .Y(n30) );
  INVX3 U90 ( .A(n18), .Y(n19) );
  INVX1 U91 ( .A(n128), .Y(n18) );
  NAND2X4 U92 ( .A(n19), .B(n127), .Y(n126) );
  INVX8 U93 ( .A(n129), .Y(n133) );
  NAND2X4 U94 ( .A(n105), .B(n30), .Y(n104) );
  INVX8 U95 ( .A(n63), .Y(SUM[1]) );
  NOR2X4 U96 ( .A(n49), .B(n164), .Y(n194) );
  INVX1 U97 ( .A(B[3]), .Y(n21) );
  INVX8 U98 ( .A(n149), .Y(n155) );
  NAND2X2 U99 ( .A(n107), .B(n89), .Y(n116) );
  BUFX16 U100 ( .A(n223), .Y(SUM[13]) );
  XOR2X2 U101 ( .A(n176), .B(n177), .Y(n223) );
  NOR2X4 U102 ( .A(n109), .B(n110), .Y(n100) );
  NAND3X2 U103 ( .A(n94), .B(n47), .C(n30), .Y(n109) );
  NAND3X4 U104 ( .A(n39), .B(n23), .C(n24), .Y(n110) );
  INVX2 U105 ( .A(n21), .Y(n22) );
  AND2X2 U106 ( .A(n30), .B(n89), .Y(n53) );
  INVXL U107 ( .A(A[3]), .Y(n72) );
  OR2X4 U108 ( .A(B[4]), .B(A[4]), .Y(n90) );
  NOR2X4 U109 ( .A(A[6]), .B(B[6]), .Y(n26) );
  NAND3X4 U110 ( .A(n45), .B(n58), .C(n47), .Y(n50) );
  OR2X4 U111 ( .A(B[5]), .B(A[5]), .Y(n89) );
  NAND2X2 U112 ( .A(n106), .B(n27), .Y(n218) );
  OR2X2 U113 ( .A(A[13]), .B(B[13]), .Y(n173) );
  INVX2 U114 ( .A(A[6]), .Y(n60) );
  AOI21X4 U115 ( .A0(n20), .A1(n180), .B0(n181), .Y(n179) );
  NAND2BX4 U116 ( .AN(n117), .B(n91), .Y(n81) );
  AND2X4 U117 ( .A(n128), .B(n124), .Y(n216) );
  NOR2X4 U118 ( .A(n117), .B(n118), .Y(n115) );
  NAND2X4 U119 ( .A(n119), .B(n39), .Y(n118) );
  INVXL U120 ( .A(n41), .Y(n42) );
  INVX4 U121 ( .A(n32), .Y(n33) );
  NOR3X4 U122 ( .A(n184), .B(n44), .C(n183), .Y(n180) );
  NAND2X1 U123 ( .A(n182), .B(n107), .Y(n184) );
  OAI2BB1X1 U124 ( .A0N(n42), .A1N(n28), .B0(n30), .Y(n163) );
  NOR2X4 U125 ( .A(A[9]), .B(B[9]), .Y(n61) );
  INVX8 U126 ( .A(n182), .Y(n154) );
  AND2X2 U127 ( .A(n128), .B(n125), .Y(n36) );
  NOR2BX4 U128 ( .AN(n108), .B(n219), .Y(n37) );
  NAND4BXL U129 ( .AN(n166), .B(n55), .C(n89), .D(n107), .Y(n150) );
  OR2X4 U130 ( .A(A[10]), .B(B[10]), .Y(n38) );
  OR2X4 U131 ( .A(B[7]), .B(A[7]), .Y(n43) );
  NAND4BX4 U132 ( .AN(n79), .B(n77), .C(n196), .D(n38), .Y(n44) );
  OAI21X2 U133 ( .A0(n137), .A1(n138), .B0(n139), .Y(n135) );
  NAND2X4 U134 ( .A(n215), .B(n216), .Y(n45) );
  NOR2BX4 U135 ( .AN(n102), .B(n26), .Y(n114) );
  INVX4 U136 ( .A(n95), .Y(n46) );
  INVX8 U137 ( .A(n46), .Y(n47) );
  NAND2X2 U138 ( .A(n73), .B(n22), .Y(n95) );
  NAND2X4 U139 ( .A(A[4]), .B(B[4]), .Y(n112) );
  AND3X4 U140 ( .A(n162), .B(n1), .C(n218), .Y(n49) );
  INVX8 U141 ( .A(n167), .Y(n58) );
  NAND2X2 U142 ( .A(B[10]), .B(A[10]), .Y(n200) );
  NAND2X4 U143 ( .A(n165), .B(n8), .Y(n164) );
  NAND2BX4 U144 ( .AN(n192), .B(n193), .Y(n191) );
  NAND2BX2 U145 ( .AN(n44), .B(n96), .Y(n193) );
  INVX8 U146 ( .A(n198), .Y(n79) );
  OAI21X4 U147 ( .A0(n14), .A1(n170), .B0(n171), .Y(n168) );
  NAND2BX4 U148 ( .AN(n51), .B(n126), .Y(n123) );
  XOR2X4 U149 ( .A(n52), .B(n53), .Y(n228) );
  NAND2X4 U150 ( .A(n120), .B(n23), .Y(n52) );
  XOR2X4 U151 ( .A(n123), .B(n54), .Y(SUM[3]) );
  INVXL U152 ( .A(n26), .Y(n55) );
  NAND3X4 U153 ( .A(n29), .B(n35), .C(n155), .Y(n186) );
  XOR2X4 U154 ( .A(n135), .B(n136), .Y(SUM[16]) );
  NAND2XL U155 ( .A(n87), .B(n43), .Y(n86) );
  XOR2X4 U156 ( .A(n134), .B(n132), .Y(n63) );
  NOR2BX4 U157 ( .AN(n9), .B(n133), .Y(n132) );
  NOR2XL U158 ( .A(n117), .B(n12), .Y(n160) );
  NAND2BX4 U159 ( .AN(n164), .B(n84), .Y(n83) );
  NAND2X4 U160 ( .A(n194), .B(n33), .Y(n96) );
  NAND3X4 U161 ( .A(n124), .B(n59), .C(n57), .Y(n111) );
  NAND2X4 U162 ( .A(n92), .B(n111), .Y(n167) );
  OAI21X4 U163 ( .A0(n115), .A1(n116), .B0(n30), .Y(n113) );
  BUFX20 U164 ( .A(n224), .Y(SUM[11]) );
  NOR2BX4 U165 ( .AN(n112), .B(n93), .Y(n119) );
  OR2X4 U166 ( .A(A[12]), .B(B[12]), .Y(n182) );
  OAI21X1 U167 ( .A0(n154), .A1(n159), .B0(n147), .Y(n181) );
  NAND3X4 U168 ( .A(n128), .B(n124), .C(n217), .Y(n92) );
  BUFX20 U169 ( .A(n222), .Y(SUM[14]) );
  BUFX20 U170 ( .A(n228), .Y(SUM[5]) );
  BUFX20 U171 ( .A(n226), .Y(SUM[9]) );
  BUFX20 U172 ( .A(n225), .Y(SUM[10]) );
  NAND2XL U173 ( .A(B[15]), .B(A[15]), .Y(n142) );
  NAND2X4 U174 ( .A(B[5]), .B(A[5]), .Y(n106) );
  OAI2BB1X4 U175 ( .A0N(n204), .A1N(n205), .B0(n206), .Y(n201) );
  AOI2BB1X1 U176 ( .A0N(n153), .A1N(n148), .B0(n145), .Y(n171) );
  NAND2XL U177 ( .A(n143), .B(n173), .Y(n170) );
  NOR2X4 U178 ( .A(n86), .B(n85), .Y(n82) );
  XOR2X4 U179 ( .A(n174), .B(n175), .Y(n222) );
  INVXL U180 ( .A(n172), .Y(n145) );
  NAND2X2 U181 ( .A(B[11]), .B(A[11]), .Y(n159) );
  NOR2BX1 U182 ( .AN(n142), .B(n64), .Y(n169) );
  XNOR2X4 U183 ( .A(n74), .B(n75), .Y(n226) );
  NOR2BX4 U184 ( .AN(n108), .B(n219), .Y(n162) );
  INVX1 U185 ( .A(n200), .Y(n208) );
  AOI21XL U186 ( .A0(n155), .A1(n156), .B0(n157), .Y(n137) );
  NAND2XL U187 ( .A(n158), .B(n159), .Y(n157) );
  OAI21XL U188 ( .A0(n160), .A1(n150), .B0(n161), .Y(n156) );
  INVXL U189 ( .A(n196), .Y(n203) );
  NAND2X1 U190 ( .A(n151), .B(n152), .Y(n138) );
  NOR2XL U191 ( .A(n64), .B(n153), .Y(n152) );
  NOR2XL U192 ( .A(n146), .B(n154), .Y(n151) );
  INVX1 U193 ( .A(n140), .Y(n139) );
  OAI21XL U194 ( .A0(n141), .A1(n64), .B0(n142), .Y(n140) );
  AOI21XL U195 ( .A0(n143), .A1(n144), .B0(n145), .Y(n141) );
  OAI21XL U196 ( .A0(n146), .A1(n147), .B0(n148), .Y(n144) );
  XOR2X1 U197 ( .A(B[16]), .B(A[16]), .Y(n136) );
  OR2X2 U198 ( .A(A[14]), .B(B[14]), .Y(n143) );
  NAND2X1 U199 ( .A(B[14]), .B(A[14]), .Y(n172) );
  INVX1 U200 ( .A(n134), .Y(n130) );
  AND2X2 U201 ( .A(n134), .B(n220), .Y(SUM[0]) );
  OR2X2 U202 ( .A(A[0]), .B(B[0]), .Y(n220) );
  NAND2X1 U203 ( .A(B[0]), .B(A[0]), .Y(n134) );
  NAND3BX4 U204 ( .AN(n213), .B(n121), .C(n214), .Y(n195) );
  OAI21X4 U205 ( .A0(n78), .A1(n79), .B0(n80), .Y(n74) );
  AOI21X4 U206 ( .A0(n81), .A1(n82), .B0(n83), .Y(n78) );
  XOR2X4 U207 ( .A(n96), .B(n97), .Y(SUM[8]) );
  XOR2X4 U208 ( .A(n98), .B(n10), .Y(SUM[7]) );
  OAI21X4 U209 ( .A0(n100), .A1(n101), .B0(n102), .Y(n98) );
  NAND2X4 U210 ( .A(n104), .B(n103), .Y(n101) );
  NOR2X4 U211 ( .A(n26), .B(n31), .Y(n103) );
  XOR2X4 U212 ( .A(n113), .B(n114), .Y(n227) );
  XOR2X4 U213 ( .A(n168), .B(n169), .Y(n221) );
  NOR2BX4 U214 ( .AN(n172), .B(n153), .Y(n175) );
  CLKINVX3 U215 ( .A(n173), .Y(n146) );
  NAND2X4 U216 ( .A(n178), .B(n179), .Y(n176) );
  OR2X4 U217 ( .A(B[4]), .B(A[4]), .Y(n107) );
  NAND2X4 U218 ( .A(n186), .B(n187), .Y(n185) );
  NAND2X4 U219 ( .A(n188), .B(n189), .Y(n187) );
  XOR2X4 U220 ( .A(n191), .B(n11), .Y(SUM[12]) );
  NAND4BX4 U221 ( .AN(n79), .B(n77), .C(n196), .D(n197), .Y(n149) );
  NAND3BX4 U222 ( .AN(n199), .B(n200), .C(n76), .Y(n189) );
  OR2X4 U223 ( .A(A[11]), .B(B[11]), .Y(n196) );
  XOR2X4 U224 ( .A(n210), .B(n211), .Y(n225) );
  OR2X4 U225 ( .A(B[10]), .B(A[10]), .Y(n197) );
  OAI2BB1X4 U226 ( .A0N(n212), .A1N(n205), .B0(n76), .Y(n210) );
  NAND2X4 U227 ( .A(n216), .B(n7), .Y(n94) );
  NOR2X4 U228 ( .A(n133), .B(n134), .Y(n215) );
  OR2X4 U229 ( .A(B[1]), .B(A[1]), .Y(n129) );
  OR2X4 U230 ( .A(B[2]), .B(A[2]), .Y(n128) );
  OR2X4 U231 ( .A(A[3]), .B(B[3]), .Y(n124) );
  NAND3X4 U232 ( .A(n37), .B(n17), .C(n218), .Y(n84) );
  NAND2X4 U233 ( .A(n87), .B(n43), .Y(n219) );
  OR2X4 U234 ( .A(B[6]), .B(A[6]), .Y(n87) );
  OR2X4 U235 ( .A(B[5]), .B(A[5]), .Y(n108) );
  OR2X4 U236 ( .A(B[7]), .B(A[7]), .Y(n88) );
  OR2X4 U237 ( .A(B[8]), .B(A[8]), .Y(n198) );
  OR2X4 U238 ( .A(B[9]), .B(A[9]), .Y(n77) );
endmodule


module butterfly_DW01_sub_124 ( A, B, DIFF );
  input [16:0] A;
  input [16:0] B;
  output [16:0] DIFF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206;

  NAND2BX2 U3 ( .AN(A[6]), .B(B[6]), .Y(n1) );
  CLKBUFX3 U4 ( .A(n196), .Y(n17) );
  NOR2BX2 U5 ( .AN(B[1]), .B(A[1]), .Y(n146) );
  NAND2BX4 U6 ( .AN(B[2]), .B(A[2]), .Y(n200) );
  NAND2X4 U7 ( .A(n66), .B(n180), .Y(n5) );
  AND3X4 U8 ( .A(n103), .B(n101), .C(n100), .Y(n60) );
  NOR2BX2 U9 ( .AN(A[1]), .B(B[1]), .Y(n147) );
  NAND2BX2 U10 ( .AN(B[3]), .B(A[3]), .Y(n83) );
  NAND3BX4 U11 ( .AN(n128), .B(n84), .C(n129), .Y(n127) );
  NAND2X2 U12 ( .A(n64), .B(n62), .Y(n186) );
  NAND4BX4 U13 ( .AN(n7), .B(n30), .C(n26), .D(n205), .Y(n22) );
  AND2X2 U14 ( .A(n180), .B(n62), .Y(n40) );
  OAI21X4 U15 ( .A0(n195), .A1(n61), .B0(n196), .Y(n194) );
  NAND2X2 U16 ( .A(n135), .B(n137), .Y(n156) );
  NAND2BX2 U17 ( .AN(B[14]), .B(A[14]), .Y(n135) );
  BUFX12 U18 ( .A(n1), .Y(n26) );
  INVX4 U19 ( .A(n195), .Y(n28) );
  INVX4 U20 ( .A(n102), .Y(n116) );
  AOI31X1 U21 ( .A0(n67), .A1(n69), .A2(n22), .B0(n5), .Y(n189) );
  NOR2X1 U22 ( .A(n158), .B(n136), .Y(n155) );
  NAND2X1 U23 ( .A(n149), .B(n161), .Y(n165) );
  INVX1 U24 ( .A(n137), .Y(n167) );
  INVX1 U25 ( .A(n149), .Y(n46) );
  INVX2 U26 ( .A(n13), .Y(n14) );
  INVX2 U27 ( .A(n55), .Y(n109) );
  OAI21X2 U28 ( .A0(n115), .A1(n116), .B0(n201), .Y(n112) );
  CLKINVX3 U29 ( .A(n71), .Y(n33) );
  BUFX3 U30 ( .A(n66), .Y(n8) );
  BUFX8 U31 ( .A(n179), .Y(n23) );
  AOI21X2 U32 ( .A0(n197), .A1(n198), .B0(n199), .Y(n191) );
  INVX1 U33 ( .A(n171), .Y(n48) );
  NAND2X1 U34 ( .A(n103), .B(n83), .Y(n110) );
  NAND3X2 U35 ( .A(n101), .B(n102), .C(n103), .Y(n99) );
  NAND4X4 U36 ( .A(n100), .B(n94), .C(n95), .D(n96), .Y(n91) );
  NAND3X2 U37 ( .A(n2), .B(n47), .C(n91), .Y(n74) );
  AOI21X2 U38 ( .A0(n90), .A1(n91), .B0(n92), .Y(n89) );
  NAND3X4 U39 ( .A(n15), .B(n83), .C(n91), .Y(n107) );
  INVX4 U40 ( .A(n100), .Y(n93) );
  AND2X2 U41 ( .A(n83), .B(n15), .Y(n2) );
  AND2X4 U42 ( .A(n159), .B(n35), .Y(n3) );
  CLKINVX3 U43 ( .A(n161), .Y(n158) );
  INVXL U44 ( .A(n15), .Y(n84) );
  AOI21X2 U45 ( .A0(n61), .A1(n195), .B0(n206), .Y(n7) );
  INVX4 U46 ( .A(n83), .Y(n199) );
  AOI21X2 U47 ( .A0(n146), .A1(n200), .B0(n93), .Y(n197) );
  AND2X2 U48 ( .A(A[10]), .B(n4), .Y(n177) );
  INVX4 U49 ( .A(B[10]), .Y(n4) );
  OAI21X4 U50 ( .A0(n174), .A1(n12), .B0(n19), .Y(n159) );
  OR2X4 U51 ( .A(n61), .B(n195), .Y(n204) );
  NAND4BX2 U52 ( .AN(n138), .B(n16), .C(n35), .D(n6), .Y(n151) );
  INVX1 U53 ( .A(n169), .Y(n6) );
  AND2X2 U54 ( .A(n205), .B(n73), .Y(n21) );
  NOR2BX4 U55 ( .AN(n23), .B(n5), .Y(n184) );
  NAND3X4 U56 ( .A(n159), .B(n16), .C(n35), .Y(n58) );
  INVX8 U57 ( .A(B[5]), .Y(n195) );
  INVX8 U58 ( .A(n32), .Y(n169) );
  NAND3BX2 U59 ( .AN(n147), .B(n119), .C(n200), .Y(n94) );
  NAND2BX2 U60 ( .AN(B[13]), .B(A[13]), .Y(n137) );
  INVXL U61 ( .A(n76), .Y(n144) );
  NAND2X4 U62 ( .A(n82), .B(n80), .Y(n92) );
  CLKINVX4 U63 ( .A(n34), .Y(n9) );
  INVX3 U64 ( .A(n34), .Y(n35) );
  XOR2X4 U65 ( .A(n10), .B(n11), .Y(DIFF[10]) );
  OR2X4 U66 ( .A(n189), .B(n190), .Y(n10) );
  AND2X2 U67 ( .A(n23), .B(n188), .Y(n11) );
  NAND2BX4 U68 ( .AN(A[1]), .B(B[1]), .Y(n102) );
  XOR2X2 U69 ( .A(n117), .B(n118), .Y(DIFF[1]) );
  NAND3X4 U70 ( .A(n9), .B(n161), .C(n149), .Y(n168) );
  NAND2BX2 U71 ( .AN(B[1]), .B(A[1]), .Y(n201) );
  NOR2X4 U72 ( .A(n71), .B(n181), .Y(n12) );
  NOR2BX4 U73 ( .AN(A[9]), .B(B[9]), .Y(n181) );
  CLKINVX8 U74 ( .A(n160), .Y(n34) );
  CLKINVX2 U75 ( .A(n138), .Y(n13) );
  NAND2BX4 U76 ( .AN(n116), .B(n60), .Y(n15) );
  BUFX20 U77 ( .A(A[5]), .Y(n61) );
  INVX8 U78 ( .A(n86), .Y(n81) );
  NAND2BX4 U79 ( .AN(A[3]), .B(B[3]), .Y(n103) );
  NAND2BX4 U80 ( .AN(B[7]), .B(A[7]), .Y(n73) );
  NAND2BX4 U81 ( .AN(A[12]), .B(B[12]), .Y(n16) );
  CLKINVX3 U82 ( .A(n36), .Y(n18) );
  NOR2X2 U83 ( .A(n130), .B(n138), .Y(n154) );
  INVX2 U84 ( .A(n17), .Y(n27) );
  NAND2BX2 U85 ( .AN(A[4]), .B(B[4]), .Y(n82) );
  NAND3XL U86 ( .A(n200), .B(n201), .C(n119), .Y(n198) );
  AOI21X2 U87 ( .A0(n100), .A1(n112), .B0(n113), .Y(n111) );
  NOR2X2 U88 ( .A(n99), .B(n93), .Y(n98) );
  OAI2BB1X1 U89 ( .A0N(n145), .A1N(A[2]), .B0(n146), .Y(n95) );
  NOR2X4 U90 ( .A(n176), .B(n177), .Y(n19) );
  INVX2 U91 ( .A(n141), .Y(n20) );
  CLKINVX3 U92 ( .A(n130), .Y(n141) );
  NOR2X2 U93 ( .A(n176), .B(n34), .Y(n38) );
  INVX8 U94 ( .A(n178), .Y(n176) );
  XOR2X4 U95 ( .A(n72), .B(n21), .Y(DIFF[7]) );
  NAND2X2 U96 ( .A(n125), .B(n134), .Y(n150) );
  NAND2BX4 U97 ( .AN(A[7]), .B(B[7]), .Y(n205) );
  NAND2BX4 U98 ( .AN(A[7]), .B(B[7]), .Y(n196) );
  NOR2X2 U99 ( .A(n113), .B(n93), .Y(n114) );
  INVX1 U100 ( .A(n200), .Y(n113) );
  NAND2X2 U101 ( .A(n30), .B(n86), .Y(n105) );
  INVX2 U102 ( .A(n188), .Y(n187) );
  NOR2X1 U103 ( .A(n20), .B(n131), .Y(n129) );
  AND2X4 U104 ( .A(n26), .B(n76), .Y(n24) );
  INVX20 U105 ( .A(n24), .Y(n87) );
  INVXL U106 ( .A(n3), .Y(n25) );
  NAND2BX4 U107 ( .AN(n27), .B(n122), .Y(n128) );
  XOR2X4 U108 ( .A(n107), .B(n108), .Y(DIFF[4]) );
  NOR2X2 U109 ( .A(n130), .B(n46), .Y(n57) );
  INVX4 U110 ( .A(n109), .Y(n29) );
  NOR2X2 U111 ( .A(n81), .B(n82), .Y(n77) );
  NOR2X4 U112 ( .A(n85), .B(n109), .Y(n108) );
  INVX12 U113 ( .A(n104), .Y(n85) );
  NAND2BX4 U114 ( .AN(n61), .B(n28), .Y(n30) );
  BUFX3 U115 ( .A(n180), .Y(n31) );
  NAND2BX4 U116 ( .AN(B[6]), .B(A[6]), .Y(n76) );
  NAND2X4 U117 ( .A(n65), .B(n8), .Y(n63) );
  AND2X2 U118 ( .A(n33), .B(n8), .Y(n70) );
  OAI21X4 U119 ( .A0(n173), .A1(n174), .B0(n175), .Y(n32) );
  OAI2BB1X4 U120 ( .A0N(n74), .A1N(n75), .B0(n76), .Y(n72) );
  NAND2X2 U121 ( .A(n104), .B(n83), .Y(n97) );
  XOR2X4 U122 ( .A(n110), .B(n111), .Y(DIFF[3]) );
  AOI21XL U123 ( .A0(n91), .A1(n83), .B0(n131), .Y(n143) );
  XOR2X2 U124 ( .A(n112), .B(n114), .Y(DIFF[2]) );
  NAND3XL U125 ( .A(n82), .B(n26), .C(n30), .Y(n131) );
  NAND2BX4 U126 ( .AN(A[14]), .B(B[14]), .Y(n157) );
  AND2X2 U127 ( .A(n135), .B(n157), .Y(n45) );
  OAI2BB1X4 U128 ( .A0N(n122), .A1N(n123), .B0(n124), .Y(n120) );
  CLKINVX8 U129 ( .A(n43), .Y(n36) );
  INVX8 U130 ( .A(n36), .Y(n37) );
  INVX4 U131 ( .A(n172), .Y(n49) );
  OAI21X1 U132 ( .A0(n139), .A1(n140), .B0(n25), .Y(n123) );
  XOR2X4 U133 ( .A(n183), .B(n38), .Y(DIFF[11]) );
  NAND2BX2 U134 ( .AN(B[9]), .B(A[9]), .Y(n62) );
  NAND2BX2 U135 ( .AN(A[3]), .B(B[3]), .Y(n96) );
  NAND2X4 U136 ( .A(n63), .B(n33), .Y(n39) );
  NAND2X2 U137 ( .A(n26), .B(n204), .Y(n78) );
  NOR2X4 U138 ( .A(n177), .B(n176), .Y(n175) );
  NOR2BX2 U139 ( .AN(B[9]), .B(A[9]), .Y(n182) );
  XOR2X4 U140 ( .A(n39), .B(n40), .Y(DIFF[9]) );
  AOI31X2 U141 ( .A0(n23), .A1(n186), .A2(n31), .B0(n187), .Y(n185) );
  AND3X4 U142 ( .A(n125), .B(n126), .C(n127), .Y(n124) );
  NOR2X4 U143 ( .A(n166), .B(n167), .Y(n162) );
  OAI22X4 U144 ( .A0(n169), .A1(n168), .B0(n158), .B1(n136), .Y(n166) );
  NOR2X4 U145 ( .A(n42), .B(n41), .Y(n56) );
  NAND2X4 U146 ( .A(n58), .B(n136), .Y(n41) );
  AND2X4 U147 ( .A(n57), .B(n37), .Y(n42) );
  NAND3X4 U148 ( .A(n69), .B(n68), .C(n67), .Y(n43) );
  NAND2X1 U149 ( .A(n161), .B(n137), .Y(n170) );
  NAND2X4 U150 ( .A(n16), .B(n136), .Y(n171) );
  NAND2BX4 U151 ( .AN(B[12]), .B(A[12]), .Y(n136) );
  XOR2X4 U152 ( .A(n44), .B(n45), .Y(DIFF[14]) );
  NAND2X4 U153 ( .A(n162), .B(n163), .Y(n44) );
  INVX4 U154 ( .A(n104), .Y(n206) );
  NOR2X4 U155 ( .A(n81), .B(n85), .Y(n47) );
  NAND2BX1 U156 ( .AN(B[10]), .B(A[10]), .Y(n188) );
  NAND2X4 U157 ( .A(n76), .B(n73), .Y(n202) );
  AOI21X4 U158 ( .A0(n61), .A1(n195), .B0(n206), .Y(n203) );
  AOI21X4 U159 ( .A0(n141), .A1(n18), .B0(n3), .Y(n172) );
  NAND3X4 U160 ( .A(n69), .B(n68), .C(n67), .Y(n65) );
  NAND3X4 U161 ( .A(n79), .B(n96), .C(n55), .Y(n193) );
  NAND2X4 U162 ( .A(n171), .B(n49), .Y(n50) );
  NAND2X4 U163 ( .A(n48), .B(n172), .Y(n51) );
  NAND2X4 U164 ( .A(n50), .B(n51), .Y(DIFF[12]) );
  CLKINVX8 U165 ( .A(n64), .Y(n71) );
  NAND2BX4 U166 ( .AN(A[6]), .B(B[6]), .Y(n79) );
  NAND2BX4 U167 ( .AN(A[9]), .B(B[9]), .Y(n180) );
  NOR2BX2 U168 ( .AN(n201), .B(n116), .Y(n118) );
  NAND2BX4 U169 ( .AN(B[8]), .B(A[8]), .Y(n64) );
  NAND2X4 U170 ( .A(n180), .B(n179), .Y(n174) );
  NOR2X4 U171 ( .A(n98), .B(n97), .Y(n90) );
  XOR2X4 U172 ( .A(n70), .B(n37), .Y(DIFF[8]) );
  OAI2BB1X4 U173 ( .A0N(n65), .A1N(n184), .B0(n185), .Y(n183) );
  OAI21X2 U174 ( .A0(n155), .A1(n156), .B0(n157), .Y(n152) );
  NAND2BX4 U175 ( .AN(A[2]), .B(B[2]), .Y(n100) );
  NAND2BX4 U176 ( .AN(A[4]), .B(B[4]), .Y(n55) );
  XOR2X4 U177 ( .A(n120), .B(n121), .Y(DIFF[16]) );
  AND3X4 U178 ( .A(n151), .B(n152), .C(n153), .Y(n59) );
  NAND2X2 U179 ( .A(n134), .B(n16), .Y(n148) );
  NOR2X2 U180 ( .A(n130), .B(n165), .Y(n164) );
  NAND4BX4 U181 ( .AN(n182), .B(n160), .C(n179), .D(n66), .Y(n130) );
  NAND2X2 U182 ( .A(n164), .B(n18), .Y(n163) );
  NAND2BX4 U183 ( .AN(B[11]), .B(A[11]), .Y(n178) );
  XOR2X4 U184 ( .A(n106), .B(n105), .Y(DIFF[5]) );
  AOI21X4 U185 ( .A0(n107), .A1(n29), .B0(n85), .Y(n106) );
  NAND2BX4 U186 ( .AN(A[13]), .B(B[13]), .Y(n161) );
  XOR2X4 U187 ( .A(n59), .B(n150), .Y(DIFF[15]) );
  NAND2BX4 U188 ( .AN(B[4]), .B(A[4]), .Y(n104) );
  NAND2BX4 U189 ( .AN(B[5]), .B(n61), .Y(n86) );
  XOR2X4 U190 ( .A(n56), .B(n170), .Y(DIFF[13]) );
  NAND2BX4 U191 ( .AN(A[10]), .B(B[10]), .Y(n179) );
  NOR2BX4 U192 ( .AN(n86), .B(n89), .Y(n88) );
  NAND2BX4 U193 ( .AN(n61), .B(n28), .Y(n80) );
  NAND2X4 U194 ( .A(n87), .B(n52), .Y(n53) );
  NAND2X2 U195 ( .A(n88), .B(n24), .Y(n54) );
  NAND2X4 U196 ( .A(n53), .B(n54), .Y(DIFF[6]) );
  INVX4 U197 ( .A(n88), .Y(n52) );
  NAND2BX4 U198 ( .AN(A[8]), .B(B[8]), .Y(n66) );
  NAND2BX4 U199 ( .AN(A[11]), .B(B[11]), .Y(n160) );
  NOR2X4 U200 ( .A(n14), .B(n148), .Y(n122) );
  NAND2X4 U201 ( .A(n161), .B(n157), .Y(n138) );
  NAND3X1 U202 ( .A(n65), .B(n16), .C(n154), .Y(n153) );
  NAND2BX4 U203 ( .AN(A[15]), .B(B[15]), .Y(n134) );
  NOR2X2 U204 ( .A(n77), .B(n78), .Y(n75) );
  NOR3X1 U205 ( .A(n142), .B(n143), .C(n144), .Y(n139) );
  OAI21X1 U206 ( .A0(n5), .A1(n64), .B0(n62), .Y(n190) );
  AOI21XL U207 ( .A0(n136), .A1(n137), .B0(n138), .Y(n132) );
  INVX1 U208 ( .A(n117), .Y(n115) );
  NAND2BXL U209 ( .AN(B[15]), .B(A[15]), .Y(n125) );
  OAI21XL U210 ( .A0(n132), .A1(n133), .B0(n134), .Y(n126) );
  INVXL U211 ( .A(n135), .Y(n133) );
  INVXL U212 ( .A(B[2]), .Y(n145) );
  XNOR2X1 U213 ( .A(B[16]), .B(A[16]), .Y(n121) );
  NAND2X1 U214 ( .A(n119), .B(n101), .Y(DIFF[0]) );
  NAND2BX1 U215 ( .AN(n101), .B(n119), .Y(n117) );
  NAND2BX1 U216 ( .AN(B[0]), .B(A[0]), .Y(n119) );
  NAND2BX1 U217 ( .AN(A[0]), .B(B[0]), .Y(n101) );
  NAND2XL U218 ( .A(n141), .B(n205), .Y(n140) );
  NOR2X4 U219 ( .A(n71), .B(n181), .Y(n173) );
  NAND2XL U220 ( .A(n73), .B(n22), .Y(n142) );
  NAND2BX4 U221 ( .AN(A[12]), .B(B[12]), .Y(n149) );
  OAI2BB1X4 U222 ( .A0N(n191), .A1N(n15), .B0(n192), .Y(n69) );
  NOR2X4 U223 ( .A(n194), .B(n193), .Y(n192) );
  NAND2X4 U224 ( .A(n202), .B(n205), .Y(n67) );
  NAND4BX4 U225 ( .AN(n203), .B(n204), .C(n26), .D(n205), .Y(n68) );
endmodule


module butterfly_DW01_add_185 ( A, B, SUM );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208;

  CLKINVX3 U2 ( .A(n92), .Y(n90) );
  NAND2X2 U3 ( .A(n166), .B(n167), .Y(n165) );
  NAND2X2 U4 ( .A(B[2]), .B(A[2]), .Y(n201) );
  NAND4BBX4 U5 ( .AN(n125), .BN(n1), .C(n16), .D(n158), .Y(n131) );
  NAND2X2 U6 ( .A(n25), .B(n19), .Y(n1) );
  OR2X2 U7 ( .A(B[5]), .B(A[5]), .Y(n2) );
  CLKINVX3 U8 ( .A(n49), .Y(n28) );
  NOR2X4 U9 ( .A(B[8]), .B(A[8]), .Y(n181) );
  NOR2X4 U10 ( .A(A[12]), .B(B[12]), .Y(n14) );
  NAND2X2 U11 ( .A(n126), .B(n45), .Y(n125) );
  INVX8 U12 ( .A(n23), .Y(n158) );
  BUFX1 U13 ( .A(n164), .Y(n17) );
  CLKINVX4 U14 ( .A(n136), .Y(n9) );
  NAND3X2 U15 ( .A(n75), .B(n74), .C(n63), .Y(n71) );
  NOR2X4 U16 ( .A(B[7]), .B(A[7]), .Y(n204) );
  AND2X2 U17 ( .A(n168), .B(n166), .Y(n36) );
  NOR2X4 U18 ( .A(n49), .B(n187), .Y(n189) );
  AND2X2 U19 ( .A(n11), .B(n32), .Y(n39) );
  NOR2X4 U20 ( .A(n134), .B(n121), .Y(n133) );
  NAND4X2 U21 ( .A(n53), .B(n52), .C(n54), .D(n32), .Y(n198) );
  NAND3X2 U22 ( .A(A[1]), .B(n31), .C(n94), .Y(n202) );
  BUFX16 U23 ( .A(n48), .Y(n32) );
  INVX1 U24 ( .A(n6), .Y(n7) );
  INVX1 U25 ( .A(n88), .Y(n199) );
  INVX2 U26 ( .A(B[5]), .Y(n6) );
  NOR2X2 U27 ( .A(n139), .B(n140), .Y(n135) );
  CLKINVX3 U28 ( .A(n15), .Y(n12) );
  CLKBUFXL U29 ( .A(n168), .Y(n24) );
  INVX1 U30 ( .A(n94), .Y(n91) );
  NAND2BX1 U31 ( .AN(n122), .B(n54), .Y(n69) );
  NAND2X1 U32 ( .A(n121), .B(n45), .Y(n154) );
  INVX1 U33 ( .A(n28), .Y(n13) );
  XOR2X2 U34 ( .A(n96), .B(n98), .Y(SUM[1]) );
  NAND2X1 U35 ( .A(n18), .B(n61), .Y(n5) );
  XOR2X1 U36 ( .A(B[16]), .B(A[16]), .Y(n102) );
  AOI21X1 U37 ( .A0(n112), .A1(n113), .B0(n114), .Y(n103) );
  AOI21X2 U38 ( .A0(n63), .A1(n75), .B0(n73), .Y(n78) );
  NAND2X2 U39 ( .A(n81), .B(n83), .Y(n44) );
  XOR2X4 U40 ( .A(n3), .B(n80), .Y(SUM[5]) );
  NAND2X2 U41 ( .A(n63), .B(n75), .Y(n3) );
  INVXL U42 ( .A(n82), .Y(n85) );
  OR2X2 U43 ( .A(A[11]), .B(B[11]), .Y(n168) );
  AOI21X2 U44 ( .A0(n189), .A1(n190), .B0(n191), .Y(n183) );
  NAND2X2 U45 ( .A(B[3]), .B(A[3]), .Y(n88) );
  NAND2BX4 U46 ( .AN(n6), .B(A[5]), .Y(n74) );
  NAND3BX4 U47 ( .AN(n151), .B(n54), .C(n152), .Y(n145) );
  NAND2X1 U48 ( .A(n45), .B(n126), .Y(n151) );
  NAND3X4 U49 ( .A(n4), .B(n150), .C(n16), .Y(n146) );
  AND2X2 U50 ( .A(n45), .B(n19), .Y(n4) );
  XNOR2X4 U51 ( .A(n40), .B(n5), .Y(SUM[7]) );
  AND2X2 U52 ( .A(n167), .B(n163), .Y(n173) );
  NAND2X2 U53 ( .A(B[13]), .B(A[13]), .Y(n121) );
  NAND2X2 U54 ( .A(n70), .B(n62), .Y(n40) );
  NOR2BX4 U55 ( .AN(n45), .B(n139), .Y(n148) );
  INVX8 U56 ( .A(n190), .Y(n188) );
  NOR2X2 U57 ( .A(n29), .B(n111), .Y(n152) );
  NOR2X1 U58 ( .A(A[10]), .B(B[10]), .Y(n174) );
  NOR2X2 U59 ( .A(B[11]), .B(A[11]), .Y(n180) );
  NAND2X2 U60 ( .A(B[11]), .B(A[11]), .Y(n166) );
  AND2X4 U61 ( .A(n52), .B(n19), .Y(n57) );
  NOR2X4 U62 ( .A(n120), .B(n138), .Y(n137) );
  NAND2X4 U63 ( .A(n45), .B(n25), .Y(n140) );
  BUFX12 U64 ( .A(n68), .Y(n22) );
  NOR2X2 U65 ( .A(n193), .B(n194), .Y(n192) );
  INVX8 U66 ( .A(n18), .Y(n194) );
  NAND4X4 U67 ( .A(n130), .B(n8), .C(n131), .D(n132), .Y(n128) );
  OR2X4 U68 ( .A(n141), .B(n142), .Y(n8) );
  INVX4 U69 ( .A(n9), .Y(n10) );
  BUFX8 U70 ( .A(n47), .Y(n11) );
  INVX8 U71 ( .A(n22), .Y(n15) );
  CLKINVX4 U72 ( .A(n111), .Y(n123) );
  NAND3X4 U73 ( .A(n50), .B(n13), .C(n51), .Y(n46) );
  INVX8 U74 ( .A(n15), .Y(n16) );
  NAND2BX4 U75 ( .AN(n27), .B(n22), .Y(n182) );
  NOR2BX2 U76 ( .AN(n49), .B(n181), .Y(n67) );
  NAND2X2 U77 ( .A(A[9]), .B(B[9]), .Y(n47) );
  XNOR2X2 U78 ( .A(n90), .B(n93), .Y(SUM[2]) );
  BUFX8 U79 ( .A(n41), .Y(n18) );
  OR2X4 U80 ( .A(n174), .B(n47), .Y(n163) );
  BUFX12 U81 ( .A(n18), .Y(n19) );
  OR2X2 U82 ( .A(B[7]), .B(A[7]), .Y(n41) );
  OAI22X2 U83 ( .A0(A[9]), .A1(B[9]), .B0(A[10]), .B1(B[10]), .Y(n164) );
  AND2X2 U84 ( .A(n167), .B(n190), .Y(n38) );
  NOR2BX4 U85 ( .AN(n32), .B(n181), .Y(n186) );
  INVX8 U86 ( .A(n32), .Y(n187) );
  NAND2X4 U87 ( .A(n52), .B(n32), .Y(n207) );
  BUFX1 U88 ( .A(n159), .Y(n20) );
  BUFX4 U89 ( .A(n118), .Y(n21) );
  NAND3BX4 U90 ( .AN(n44), .B(n186), .C(n185), .Y(n184) );
  NAND4X4 U91 ( .A(n145), .B(n147), .C(n146), .D(n121), .Y(n143) );
  NAND2XL U92 ( .A(n60), .B(n2), .Y(n64) );
  NAND3BX4 U93 ( .AN(n89), .B(n82), .C(n83), .Y(n75) );
  OR2X2 U94 ( .A(A[3]), .B(B[3]), .Y(n81) );
  INVX2 U95 ( .A(n81), .Y(n89) );
  NAND2X1 U96 ( .A(A[5]), .B(B[5]), .Y(n26) );
  NOR2BX2 U97 ( .AN(n126), .B(n111), .Y(n150) );
  NAND4X2 U98 ( .A(n159), .B(n62), .C(n61), .D(n177), .Y(n68) );
  NAND2X4 U99 ( .A(n43), .B(n42), .Y(n23) );
  NOR2BX4 U100 ( .AN(n60), .B(n73), .Y(n72) );
  BUFX16 U101 ( .A(n116), .Y(n25) );
  NAND3X1 U102 ( .A(n25), .B(n45), .C(n54), .Y(n142) );
  OR2X4 U103 ( .A(n205), .B(n26), .Y(n177) );
  OAI22X1 U104 ( .A0(A[10]), .A1(B[10]), .B0(B[9]), .B1(A[9]), .Y(n193) );
  OAI2BB1X2 U105 ( .A0N(n28), .A1N(n32), .B0(n11), .Y(n196) );
  NAND2X1 U106 ( .A(B[1]), .B(A[1]), .Y(n97) );
  AOI21X4 U107 ( .A0(n136), .A1(n148), .B0(n149), .Y(n147) );
  NOR2X4 U108 ( .A(n205), .B(n204), .Y(n203) );
  NAND2BX2 U109 ( .AN(n58), .B(n59), .Y(n56) );
  NAND3XL U110 ( .A(A[5]), .B(n7), .C(n60), .Y(n59) );
  OAI21X4 U111 ( .A0(n55), .A1(n56), .B0(n57), .Y(n50) );
  NOR2X2 U112 ( .A(n63), .B(n64), .Y(n55) );
  NAND3X4 U113 ( .A(n156), .B(n155), .C(n157), .Y(n153) );
  NAND4BBX2 U114 ( .AN(n23), .BN(n14), .C(n19), .D(n22), .Y(n156) );
  OAI2BB1X4 U115 ( .A0N(n33), .A1N(n20), .B0(n206), .Y(n197) );
  NOR2X4 U116 ( .A(n194), .B(n207), .Y(n206) );
  NAND2X2 U117 ( .A(n52), .B(n192), .Y(n27) );
  INVX8 U118 ( .A(n14), .Y(n126) );
  OR2X4 U119 ( .A(A[10]), .B(B[10]), .Y(n190) );
  AOI21X4 U120 ( .A0(n135), .A1(n10), .B0(n137), .Y(n130) );
  NAND2X2 U121 ( .A(B[7]), .B(A[7]), .Y(n61) );
  NAND3X4 U122 ( .A(n203), .B(n65), .C(n82), .Y(n122) );
  INVX2 U123 ( .A(B[1]), .Y(n30) );
  OR2X4 U124 ( .A(A[1]), .B(B[1]), .Y(n95) );
  INVX4 U125 ( .A(n74), .Y(n77) );
  INVX4 U126 ( .A(n2), .Y(n73) );
  NOR2X4 U127 ( .A(B[6]), .B(A[6]), .Y(n205) );
  NAND2X2 U128 ( .A(n61), .B(n62), .Y(n58) );
  NAND3BX4 U129 ( .AN(n196), .B(n198), .C(n197), .Y(n195) );
  NAND3BX4 U130 ( .AN(n205), .B(n65), .C(n79), .Y(n159) );
  NOR2BX2 U131 ( .AN(n63), .B(n85), .Y(n84) );
  OAI21X2 U132 ( .A0(n105), .A1(n106), .B0(n107), .Y(n104) );
  XOR2X4 U133 ( .A(n101), .B(n102), .Y(SUM[16]) );
  NAND2XL U134 ( .A(B[15]), .B(A[15]), .Y(n115) );
  INVX4 U135 ( .A(n45), .Y(n119) );
  BUFX20 U136 ( .A(n127), .Y(n45) );
  NOR2X2 U137 ( .A(A[10]), .B(B[10]), .Y(n178) );
  NAND4BX2 U138 ( .AN(n29), .B(n158), .C(n54), .D(n126), .Y(n157) );
  NOR2X2 U139 ( .A(A[9]), .B(B[9]), .Y(n179) );
  OR2X4 U140 ( .A(A[9]), .B(B[9]), .Y(n48) );
  NOR2X4 U141 ( .A(n179), .B(n178), .Y(n43) );
  NAND2X2 U142 ( .A(n25), .B(n45), .Y(n138) );
  INVX4 U143 ( .A(n25), .Y(n134) );
  OAI21X1 U144 ( .A0(n119), .A1(n120), .B0(n121), .Y(n117) );
  NOR2BX4 U145 ( .AN(n21), .B(n133), .Y(n132) );
  OAI21X2 U146 ( .A0(n188), .A1(n11), .B0(n167), .Y(n191) );
  NAND2XL U147 ( .A(n12), .B(n19), .Y(n110) );
  INVX8 U148 ( .A(n44), .Y(n54) );
  NAND2X1 U149 ( .A(n60), .B(n62), .Y(n37) );
  NAND2X2 U150 ( .A(n103), .B(n104), .Y(n101) );
  NOR2X4 U151 ( .A(n188), .B(n29), .Y(n185) );
  NOR2X4 U152 ( .A(n180), .B(n181), .Y(n42) );
  AND3X2 U153 ( .A(n61), .B(n62), .C(n177), .Y(n33) );
  OAI2BB1X4 U154 ( .A0N(n22), .A1N(n19), .B0(n69), .Y(n66) );
  AOI21X4 U155 ( .A0(n160), .A1(n136), .B0(n161), .Y(n155) );
  NAND2X4 U156 ( .A(n72), .B(n71), .Y(n70) );
  OR2X4 U157 ( .A(B[13]), .B(A[13]), .Y(n127) );
  INVX4 U158 ( .A(n63), .Y(n79) );
  NOR2BX2 U159 ( .AN(n97), .B(n99), .Y(n98) );
  NAND2X4 U160 ( .A(B[8]), .B(A[8]), .Y(n49) );
  INVX8 U161 ( .A(n53), .Y(n29) );
  NAND2X4 U162 ( .A(n126), .B(n168), .Y(n139) );
  XOR2X4 U163 ( .A(n86), .B(n87), .Y(SUM[3]) );
  OAI21X2 U164 ( .A0(n90), .A1(n91), .B0(n201), .Y(n86) );
  CLKINVX8 U165 ( .A(n122), .Y(n53) );
  OR2X4 U166 ( .A(A[15]), .B(B[15]), .Y(n112) );
  NOR2X2 U167 ( .A(n119), .B(n120), .Y(n149) );
  NAND2X2 U168 ( .A(B[12]), .B(A[12]), .Y(n120) );
  CLKINVX3 U169 ( .A(n30), .Y(n31) );
  AOI2BB1X4 U170 ( .A0N(n164), .A1N(n49), .B0(n165), .Y(n162) );
  NAND3X4 U171 ( .A(n182), .B(n183), .C(n184), .Y(n35) );
  NAND3X1 U172 ( .A(n61), .B(n175), .C(n69), .Y(n170) );
  XOR2X4 U173 ( .A(n143), .B(n144), .Y(SUM[14]) );
  NAND3XL U174 ( .A(n62), .B(n159), .C(n177), .Y(n176) );
  NAND3X1 U175 ( .A(n126), .B(n123), .C(n53), .Y(n141) );
  OR2X4 U176 ( .A(A[2]), .B(B[2]), .Y(n94) );
  OR2X4 U177 ( .A(A[14]), .B(B[14]), .Y(n116) );
  XNOR2X4 U178 ( .A(n153), .B(n154), .Y(SUM[13]) );
  INVX1 U179 ( .A(n120), .Y(n161) );
  OR2X4 U180 ( .A(A[4]), .B(B[4]), .Y(n82) );
  NAND3X1 U181 ( .A(n53), .B(n54), .C(n52), .Y(n51) );
  NOR2BX2 U182 ( .AN(n201), .B(n91), .Y(n93) );
  OAI2BB1X4 U183 ( .A0N(n123), .A1N(n170), .B0(n108), .Y(n169) );
  AND2X2 U184 ( .A(n120), .B(n126), .Y(n34) );
  XOR2X2 U185 ( .A(n54), .B(n84), .Y(SUM[4]) );
  INVX2 U186 ( .A(n139), .Y(n160) );
  XNOR2X4 U187 ( .A(n128), .B(n129), .Y(SUM[15]) );
  XOR2X4 U188 ( .A(n35), .B(n36), .Y(SUM[11]) );
  XOR2X4 U189 ( .A(n37), .B(n76), .Y(SUM[6]) );
  XOR2X4 U190 ( .A(n195), .B(n38), .Y(SUM[10]) );
  XOR2X4 U191 ( .A(n46), .B(n39), .Y(SUM[9]) );
  NAND2X4 U192 ( .A(n42), .B(n43), .Y(n111) );
  INVXL U193 ( .A(n95), .Y(n99) );
  NOR2BX2 U194 ( .AN(n88), .B(n89), .Y(n87) );
  NAND2X1 U195 ( .A(n176), .B(n19), .Y(n175) );
  NOR2X1 U196 ( .A(n124), .B(n125), .Y(n107) );
  NAND2X1 U197 ( .A(n115), .B(n112), .Y(n129) );
  INVXL U198 ( .A(n108), .Y(n106) );
  INVX1 U199 ( .A(n115), .Y(n114) );
  OAI2BB1X2 U200 ( .A0N(n95), .A1N(n96), .B0(n97), .Y(n92) );
  AOI21XL U201 ( .A0(n109), .A1(n110), .B0(n23), .Y(n105) );
  NAND3XL U202 ( .A(n83), .B(n53), .C(n81), .Y(n109) );
  NAND3BX2 U203 ( .AN(n100), .B(n94), .C(n95), .Y(n200) );
  INVX1 U204 ( .A(n100), .Y(n96) );
  AND2X2 U205 ( .A(n100), .B(n208), .Y(SUM[0]) );
  OR2X2 U206 ( .A(A[0]), .B(B[0]), .Y(n208) );
  NAND2X1 U207 ( .A(B[0]), .B(A[0]), .Y(n100) );
  NAND2XL U208 ( .A(A[8]), .B(B[8]), .Y(n172) );
  NAND2X2 U209 ( .A(B[6]), .B(A[6]), .Y(n62) );
  OAI2BB1X1 U210 ( .A0N(n25), .A1N(n117), .B0(n21), .Y(n113) );
  NAND2XL U211 ( .A(n25), .B(n112), .Y(n124) );
  NAND2XL U212 ( .A(B[14]), .B(A[14]), .Y(n118) );
  NAND2X2 U213 ( .A(B[10]), .B(A[10]), .Y(n167) );
  XOR2X4 U214 ( .A(n66), .B(n67), .Y(SUM[8]) );
  NOR2X4 U215 ( .A(n78), .B(n77), .Y(n76) );
  NOR2BX4 U216 ( .AN(n74), .B(n73), .Y(n80) );
  NOR2BX4 U217 ( .AN(n21), .B(n134), .Y(n144) );
  NAND2X4 U218 ( .A(n162), .B(n163), .Y(n136) );
  XOR2X4 U219 ( .A(n169), .B(n34), .Y(SUM[12]) );
  NAND2X4 U220 ( .A(n24), .B(n171), .Y(n108) );
  OAI211X2 U221 ( .A0(n17), .A1(n172), .B0(n166), .C0(n173), .Y(n171) );
  NAND4BX4 U222 ( .AN(n199), .B(n200), .C(n201), .D(n202), .Y(n83) );
  OR2X4 U223 ( .A(B[8]), .B(A[8]), .Y(n52) );
  NAND2X4 U224 ( .A(B[4]), .B(A[4]), .Y(n63) );
  OR2X4 U225 ( .A(B[5]), .B(A[5]), .Y(n65) );
  OR2X4 U226 ( .A(B[6]), .B(A[6]), .Y(n60) );
endmodule


module butterfly ( calc_in, rotation, calc_out );
  input [135:0] calc_in;
  input [2:0] rotation;
  output [135:0] calc_out;
  wire   n135, n136, n137, n138, n139, n140, n141, n142, n143, N6, N9, N42,
         N43, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296,
         N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285,
         N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274,
         N273, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229,
         N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218,
         N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207,
         N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196,
         N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185,
         N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174,
         N173, N172, N171, N136, N135, N134, N133, N132, N131, N130, N129,
         N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118,
         N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107,
         N106, N105, N104, N103, N340, N339, N338, N337, N336, N335, N334,
         N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323,
         N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312,
         N311, N310, N309, N308, N307, N272, N271, N270, N269, N268, N267,
         N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256,
         N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245,
         N244, N243, N242, N241, N240, N239, N170, N169, N168, N167, N166,
         N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155,
         N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144,
         N143, N142, N141, N140, N139, N138, N137, N99, N98, N97, N96, N95,
         N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81,
         N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N102,
         N101, N100, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n22, n23, n24, n25, n26, n27, n28, n29, n30, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n62, n63,
         n64, n65, n66, n68, n69, n71, n73, n75, n76, n78, n79, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110;
  wire   [16:0] temp_2_1_real;
  wire   [16:0] temp_2_2_real;
  wire   [16:0] temp_2_1_imag;
  wire   [16:0] temp_2_2_imag;
  wire   [16:0] temp_3_1_real;
  wire   [16:0] temp_3_2_real;
  wire   [16:0] temp_3_1_imag;
  wire   [16:0] temp_3_2_imag;
  wire   [16:0] temp_4_1_real;
  wire   [16:0] temp_4_2_real;
  wire   [16:0] temp_4_1_imag;
  wire   [16:0] temp_4_2_imag;
  wire   [16:0] temp_1_real;
  wire   [16:0] temp_1_imag;
  wire   [16:0] temp_2_real;
  wire   [16:0] temp_2_imag;
  wire   [16:0] temp_3_real;
  wire   [16:0] temp_3_imag;

  multi16_0 multiBRR ( .in_17bit({n106, calc_in[66:51]}), .in_8bit({1'b0, n12, 
        n17, 1'b1, n82, n102, n12, n99}), .out(temp_2_1_real) );
  multi16_11 multiBII ( .in_17bit(calc_in[50:34]), .in_8bit({n89, n91, n88, 
        1'b0, n92, n100, n89, n90}), .out(temp_2_2_real) );
  multi16_10 multiBRI ( .in_17bit({n106, calc_in[66:51]}), .in_8bit({n89, n91, 
        n88, 1'b0, n92, n100, n89, n90}), .out(temp_2_1_imag) );
  multi16_9 multiBIR ( .in_17bit(calc_in[50:34]), .in_8bit({1'b0, n12, n18, 
        1'b1, n82, n102, n12, N9}), .out(temp_2_2_imag) );
  multi16_8 multiCRR ( .in_17bit({n108, calc_in[100:85]}), .in_8bit({n96, n102, 
        N9, n102, n102, n97, n19, n41}), .out(temp_3_1_real) );
  multi16_7 multiCII ( .in_17bit({n107, calc_in[83:68]}), .in_8bit({n89, 1'b0, 
        n92, 1'b0, 1'b0, n92, n92, n88}), .out(temp_3_2_real) );
  multi16_6 multiCRI ( .in_17bit({n108, calc_in[100:85]}), .in_8bit({n89, 1'b0, 
        n92, 1'b0, 1'b0, n92, n92, n88}), .out(temp_3_1_imag) );
  multi16_5 multiCIR ( .in_17bit({n107, calc_in[83:68]}), .in_8bit({n96, n102, 
        N9, n102, n102, n98, n20, n41}), .out(temp_3_2_imag) );
  multi16_4 multiDRR ( .in_17bit(calc_in[135:119]), .in_8bit({n103, n16, n12, 
        n102, n98, n83, n11, n102}), .out(temp_4_1_real) );
  multi16_3 multiDII ( .in_17bit({n109, calc_in[117:102]}), .in_8bit({n101, 
        1'b0, n104, n14, n90, n88, n100, n13}), .out(temp_4_2_real) );
  multi16_2 multiDRI ( .in_17bit(calc_in[135:119]), .in_8bit({n44, 1'b0, n104, 
        n13, n90, n88, n100, n14}), .out(temp_4_1_imag) );
  multi16_1 multiDIR ( .in_17bit({n109, calc_in[117:102]}), .in_8bit({n103, 
        n16, n12, n102, n97, n83, n11, n102}), .out(temp_4_2_imag) );
  butterfly_DW01_add_18 add_0_root_sub_0_root_add_301 ( .A({N340, N339, N338, 
        N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, 
        N325, N324}), .B({N323, N322, N321, N320, N319, N318, N317, N316, N315, 
        N314, N313, N312, N311, n57, N309, N308, N307}), .SUM({calc_out[50:49], 
        n139, calc_out[47:34]}) );
  butterfly_DW01_add_49 add_2_root_add_0_root_add_292_3 ( .A({calc_in[33:21], 
        n9, calc_in[19:18], n26}), .B({temp_2_real[16:15], n79, 
        temp_2_real[13:9], n32, n75, temp_2_real[6], n54, temp_2_real[4:0]}), 
        .SUM({N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, 
        N90, N89, N88, N87, N86}) );
  butterfly_DW01_add_50 add_0_root_add_0_root_add_293_3 ( .A({N136, N135, N134, 
        N133, n86, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, 
        N121, N120}), .B({N119, N118, N117, N116, N115, N114, N113, N112, N111, 
        N110, N109, N108, N107, N106, N105, N104, N103}), .SUM({
        calc_out[16:14], n142, calc_out[12:10], n143, calc_out[8:0]}) );
  butterfly_DW01_add_52 add_0_root_sub_0_root_add_298 ( .A({N238, N237, N236, 
        N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, 
        N223, N222}), .B({N221, N220, N219, N218, N217, N216, N215, N214, N213, 
        N212, N211, N210, N209, N208, N207, N206, N205}), .SUM(
        calc_out[135:119]) );
  butterfly_DW01_add_56 add_279 ( .A(temp_3_1_imag), .B(temp_3_2_imag), .SUM(
        temp_2_imag) );
  butterfly_DW01_sub_56 sub_2_root_sub_0_root_add_298 ( .A({calc_in[33:21], n9, 
        calc_in[19:18], n26}), .B({temp_1_imag[16:13], n40, temp_1_imag[11:9], 
        n68, n63, temp_1_imag[6:4], n62, temp_1_imag[2:0]}), .DIFF({N238, N237, 
        N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, 
        N224, N223, N222}) );
  butterfly_DW01_add_66 add_0_root_sub_0_root_sub_296_2 ( .A({N204, N203, N202, 
        N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, 
        N189, N188}), .B({N187, N186, N185, N184, N183, N182, N181, N180, N179, 
        N178, N177, N176, N175, N174, N173, N172, N171}), .SUM({
        calc_out[84:82], n137, calc_out[80:68]}) );
  butterfly_DW01_sub_74 sub_2_root_sub_0_root_sub_299_2 ( .A({calc_in[16:6], 
        n105, calc_in[4:0]}), .B({temp_3_real[16:15], n55, temp_3_real[13], 
        n64, temp_3_real[11:6], n93, n87, temp_3_real[3:0]}), .DIFF({N272, 
        N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, 
        N259, N258, N257, N256}) );
  butterfly_DW01_sub_76 sub_0_root_sub_0_root_sub_300_2 ( .A({N306, N305, N304, 
        N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, 
        N291, N290}), .B({N289, N288, N287, N286, N285, N284, N283, N282, N281, 
        N280, N279, N278, N277, N276, N275, N274, N273}), .DIFF({
        calc_out[67:63], n138, calc_out[61:51]}) );
  butterfly_DW01_sub_78 sub_1_root_sub_0_root_add_301 ( .A({temp_3_real[16:15], 
        n55, temp_3_real[13], n64, temp_3_real[11], n49, temp_3_real[9:6], n93, 
        n87, temp_3_real[3:0]}), .B({temp_2_imag[16:6], n94, temp_2_imag[4], 
        n78, temp_2_imag[2:0]}), .DIFF({N323, N322, N321, N320, N319, N318, 
        N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307}) );
  butterfly_DW01_sub_84 sub_275 ( .A(temp_2_1_real), .B({temp_2_2_real[16:3], 
        n51, n30, temp_2_2_real[0]}), .DIFF(temp_1_real) );
  butterfly_DW01_add_116 add_282 ( .A(temp_4_1_imag), .B(temp_4_2_imag), .SUM(
        temp_3_imag) );
  butterfly_DW01_add_119 add_1_root_sub_0_root_sub_295_2 ( .A({
        temp_1_real[16:14], n36, temp_1_real[12:9], n53, temp_1_real[7:6], n95, 
        temp_1_real[4:0]}), .B({temp_3_real[16:15], n55, temp_3_real[13], n64, 
        temp_3_real[11], n49, temp_3_real[9:8], n47, temp_3_real[6], n93, n87, 
        temp_3_real[3:0]}), .SUM({N153, N152, N151, N150, N149, N148, N147, 
        N146, N145, N144, N143, N142, N141, N140, N139, N138, N137}) );
  butterfly_DW01_add_128 add_1_root_sub_0_root_sub_300_2 ( .A({temp_3_imag[16], 
        n37, temp_3_imag[14:12], n65, n29, temp_3_imag[9:4], n56, n38, 
        temp_3_imag[1:0]}), .B({temp_2_real[16:15], n79, temp_2_real[13:11], 
        n35, temp_2_real[9], n32, n75, temp_2_real[6], n28, temp_2_real[4:0]}), 
        .SUM({N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, 
        N278, N277, N276, N275, N274, N273}) );
  butterfly_DW01_add_129 add_2_root_add_0_root_add_293_3 ( .A({calc_in[16:6], 
        n105, calc_in[4:0]}), .B({temp_2_imag[16:8], n39, temp_2_imag[6], n94, 
        temp_2_imag[4], n78, temp_2_imag[2:0]}), .SUM({N136, N135, N134, N133, 
        N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, 
        N120}) );
  butterfly_DW01_sub_101 sub_281 ( .A({temp_4_1_real[16:6], n27, 
        temp_4_1_real[4:0]}), .B(temp_4_2_real), .DIFF(temp_3_real) );
  butterfly_DW01_sub_96 sub_1_root_sub_0_root_add_298 ( .A({temp_3_imag[16], 
        n37, temp_3_imag[14:12], n65, temp_3_imag[10:4], n56, n7, 
        temp_3_imag[1:0]}), .B({temp_2_real[16:15], n79, n24, 
        temp_2_real[12:9], n32, n75, temp_2_real[6], n54, temp_2_real[4:0]}), 
        .DIFF({N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, 
        N211, N210, N209, N208, N207, N206, N205}) );
  butterfly_DW01_sub_104 sub_2_root_sub_0_root_sub_296_2 ( .A({calc_in[16:6], 
        n105, calc_in[4:0]}), .B({temp_1_imag[16:13], n40, temp_1_imag[11:9], 
        n68, n63, temp_1_imag[6:4], n62, temp_1_imag[2:0]}), .DIFF({N204, N203, 
        N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, 
        N190, N189, N188}) );
  butterfly_DW01_add_151 add_2_root_sub_0_root_sub_300_2 ( .A({calc_in[33:21], 
        n9, calc_in[19:18], n26}), .B({temp_1_imag[16:13], n40, 
        temp_1_imag[11:9], n68, n63, temp_1_imag[6:4], n62, temp_1_imag[2:0]}), 
        .SUM({N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, 
        N295, N294, N293, N292, N291, N290}) );
  butterfly_DW01_add_141 add_0_root_sub_0_root_sub_299_2 ( .A({N272, N271, 
        N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, 
        N258, N257, N256}), .B({N255, N254, N253, N252, N251, N250, N249, N248, 
        N247, N246, N245, N244, N243, N242, N241, N240, N239}), .SUM({
        calc_out[118:117], n135, calc_out[115:114], n136, calc_out[112:102]})
         );
  butterfly_DW01_sub_115 sub_278 ( .A({temp_3_1_real[16:5], n52, 
        temp_3_1_real[3:0]}), .B(temp_3_2_real), .DIFF(temp_2_real) );
  butterfly_DW01_add_158 add_0_root_add_0_root_add_292_3 ( .A({N102, N101, 
        N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, 
        N86}), .B({N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, 
        n46, N72, N71, N70, N69}), .SUM({n140, calc_out[32:28], n141, 
        calc_out[26:17]}) );
  butterfly_DW01_sub_118 sub_2_root_sub_0_root_add_301 ( .A({calc_in[16:6], 
        n105, calc_in[4:0]}), .B({temp_1_real[16:14], n36, temp_1_real[12:9], 
        n53, temp_1_real[7:6], n95, temp_1_real[4:0]}), .DIFF({N340, N339, 
        N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, 
        N326, N325, N324}) );
  butterfly_DW01_add_164 add_1_root_add_0_root_add_292_3 ( .A({
        temp_1_real[16:14], n36, temp_1_real[12:9], n53, temp_1_real[7:6], n95, 
        temp_1_real[4:0]}), .B({temp_3_real[16:15], n55, temp_3_real[13], n64, 
        temp_3_real[11:8], n47, temp_3_real[6], n93, n87, temp_3_real[3:0]}), 
        .SUM({N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, 
        N72, N71, N70, N69}) );
  butterfly_DW01_add_170 add_2_root_sub_0_root_sub_295_2 ( .A({calc_in[33:21], 
        n9, calc_in[19:18], n26}), .B({temp_2_real[16:15], n79, 
        temp_2_real[13:9], n32, n75, temp_2_real[6], n28, temp_2_real[4:0]}), 
        .SUM({N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, 
        N159, N158, N157, N156, N155, N154}) );
  butterfly_DW01_sub_121 sub_0_root_sub_0_root_sub_295_2 ( .A({N170, N169, 
        N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, 
        N156, N155, N154}), .B({N153, N152, N151, N150, N149, N148, N147, N146, 
        N145, n50, N143, N142, N141, N140, N139, N138, N137}), .DIFF(
        calc_out[101:85]) );
  butterfly_DW01_sub_123 sub_1_root_sub_0_root_sub_299_2 ( .A({
        temp_1_real[16:14], n36, temp_1_real[12:9], n53, temp_1_real[7:6], n95, 
        temp_1_real[4:0]}), .B({temp_2_imag[16:8], n43, temp_2_imag[6], n94, 
        temp_2_imag[4], n78, temp_2_imag[2:0]}), .DIFF({N255, N254, N253, N252, 
        N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, 
        N239}) );
  butterfly_DW01_add_184 add_276 ( .A(temp_2_1_imag), .B({temp_2_2_imag[16:6], 
        n45, temp_2_2_imag[4:0]}), .SUM(temp_1_imag) );
  butterfly_DW01_sub_124 sub_1_root_sub_0_root_sub_296_2 ( .A({
        temp_2_imag[16:6], n94, temp_2_imag[4], n78, temp_2_imag[2:0]}), .B({
        temp_3_imag[16], n37, temp_3_imag[14:12], n65, temp_3_imag[10:4], n56, 
        n7, temp_3_imag[1:0]}), .DIFF({N187, N186, N185, N184, N183, N182, 
        N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171}) );
  butterfly_DW01_add_185 add_1_root_add_0_root_add_293_3 ( .A({
        temp_1_imag[16:13], n40, temp_1_imag[11:10], n25, n68, n63, 
        temp_1_imag[6:5], n59, n62, temp_1_imag[2:0]}), .B({temp_3_imag[16:12], 
        n65, temp_3_imag[10:4], n56, n38, temp_3_imag[1:0]}), .SUM({N119, N118, 
        N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, 
        N105, N104, N103}) );
  BUFX16 U9 ( .A(calc_in[67]), .Y(n106) );
  NAND2X4 U10 ( .A(rotation[1]), .B(rotation[2]), .Y(N6) );
  BUFX20 U11 ( .A(calc_in[84]), .Y(n107) );
  CLKINVX4 U12 ( .A(temp_2_real[13]), .Y(n23) );
  BUFX20 U13 ( .A(N144), .Y(n50) );
  INVX4 U14 ( .A(N42), .Y(n22) );
  BUFX8 U15 ( .A(temp_3_imag[2]), .Y(n7) );
  CLKBUFX8 U16 ( .A(temp_3_imag[2]), .Y(n38) );
  INVX2 U17 ( .A(rotation[0]), .Y(n110) );
  CLKINVX4 U18 ( .A(temp_1_imag[4]), .Y(n58) );
  BUFX20 U19 ( .A(calc_in[101]), .Y(n108) );
  BUFX20 U20 ( .A(temp_1_imag[12]), .Y(n40) );
  BUFX12 U21 ( .A(temp_2_2_real[2]), .Y(n51) );
  INVX4 U22 ( .A(n110), .Y(n33) );
  INVX4 U23 ( .A(calc_in[20]), .Y(n8) );
  INVX8 U24 ( .A(n8), .Y(n9) );
  INVX4 U25 ( .A(n23), .Y(n24) );
  BUFX20 U26 ( .A(temp_3_real[4]), .Y(n87) );
  BUFX12 U27 ( .A(temp_2_imag[7]), .Y(n43) );
  BUFX3 U28 ( .A(N43), .Y(n12) );
  AND2X1 U29 ( .A(n103), .B(n110), .Y(n10) );
  CLKBUFX8 U30 ( .A(calc_in[5]), .Y(n105) );
  INVX8 U31 ( .A(N43), .Y(n96) );
  OR2X2 U32 ( .A(n82), .B(n42), .Y(n11) );
  INVXL U33 ( .A(n100), .Y(n98) );
  INVXL U34 ( .A(n12), .Y(n13) );
  INVXL U35 ( .A(n12), .Y(n14) );
  BUFX16 U36 ( .A(n143), .Y(calc_out[9]) );
  XOR2X4 U37 ( .A(rotation[1]), .B(rotation[0]), .Y(n84) );
  INVX8 U38 ( .A(n99), .Y(n101) );
  INVX8 U39 ( .A(N6), .Y(n103) );
  BUFX20 U40 ( .A(temp_3_real[7]), .Y(n47) );
  INVXL U41 ( .A(n41), .Y(n15) );
  INVXL U42 ( .A(n15), .Y(n16) );
  INVXL U43 ( .A(n10), .Y(n17) );
  INVXL U44 ( .A(n10), .Y(n18) );
  INVXL U45 ( .A(n10), .Y(n19) );
  INVXL U46 ( .A(n10), .Y(n20) );
  BUFX20 U47 ( .A(n142), .Y(calc_out[13]) );
  BUFX20 U48 ( .A(temp_2_real[5]), .Y(n54) );
  BUFX20 U49 ( .A(temp_3_imag[10]), .Y(n29) );
  INVX8 U50 ( .A(n139), .Y(n60) );
  BUFX16 U51 ( .A(temp_2_real[5]), .Y(n28) );
  BUFX20 U52 ( .A(temp_2_real[8]), .Y(n32) );
  BUFX20 U53 ( .A(temp_1_imag[9]), .Y(n25) );
  BUFX16 U54 ( .A(calc_in[17]), .Y(n26) );
  INVX8 U55 ( .A(n44), .Y(n99) );
  BUFX8 U56 ( .A(temp_4_1_real[5]), .Y(n27) );
  INVX4 U57 ( .A(temp_2_real[10]), .Y(n34) );
  INVX8 U58 ( .A(temp_3_real[10]), .Y(n48) );
  BUFX20 U59 ( .A(temp_2_imag[7]), .Y(n39) );
  AND2X2 U60 ( .A(rotation[1]), .B(rotation[2]), .Y(n85) );
  BUFX20 U61 ( .A(temp_1_real[13]), .Y(n36) );
  BUFX8 U62 ( .A(temp_2_2_real[1]), .Y(n30) );
  INVXL U63 ( .A(n101), .Y(N9) );
  INVXL U64 ( .A(N9), .Y(n100) );
  INVX8 U65 ( .A(n58), .Y(n59) );
  BUFX20 U66 ( .A(calc_in[118]), .Y(n109) );
  INVX8 U67 ( .A(n34), .Y(n35) );
  NAND2X4 U68 ( .A(n85), .B(n33), .Y(N43) );
  BUFX12 U69 ( .A(temp_3_imag[15]), .Y(n37) );
  BUFX16 U70 ( .A(N132), .Y(n86) );
  BUFX20 U71 ( .A(temp_3_imag[3]), .Y(n56) );
  BUFX8 U72 ( .A(N73), .Y(n46) );
  INVXL U73 ( .A(n89), .Y(n41) );
  DLY1X1 U74 ( .A(rotation[1]), .Y(n42) );
  INVX8 U75 ( .A(n137), .Y(n71) );
  AND2X4 U76 ( .A(n84), .B(rotation[2]), .Y(n44) );
  BUFX8 U77 ( .A(temp_2_2_imag[5]), .Y(n45) );
  BUFX20 U78 ( .A(n140), .Y(calc_out[33]) );
  BUFX8 U79 ( .A(temp_3_1_real[4]), .Y(n52) );
  BUFX20 U80 ( .A(temp_2_real[7]), .Y(n75) );
  BUFX20 U81 ( .A(temp_2_imag[5]), .Y(n94) );
  BUFX20 U82 ( .A(temp_2_imag[3]), .Y(n78) );
  INVX8 U83 ( .A(n48), .Y(n49) );
  BUFX20 U84 ( .A(temp_3_real[12]), .Y(n64) );
  BUFX20 U85 ( .A(temp_1_imag[3]), .Y(n62) );
  BUFX20 U86 ( .A(temp_1_imag[8]), .Y(n68) );
  BUFX20 U87 ( .A(temp_1_imag[7]), .Y(n63) );
  BUFX20 U88 ( .A(temp_3_real[14]), .Y(n55) );
  BUFX20 U89 ( .A(temp_3_imag[11]), .Y(n65) );
  BUFX20 U90 ( .A(temp_1_real[8]), .Y(n53) );
  BUFX8 U91 ( .A(N310), .Y(n57) );
  INVX8 U92 ( .A(n60), .Y(calc_out[48]) );
  CLKINVX8 U93 ( .A(n141), .Y(n66) );
  INVX8 U94 ( .A(n66), .Y(calc_out[27]) );
  CLKINVX8 U95 ( .A(n136), .Y(n69) );
  INVX8 U96 ( .A(n69), .Y(calc_out[113]) );
  INVX8 U97 ( .A(n71), .Y(calc_out[81]) );
  CLKINVX8 U98 ( .A(n138), .Y(n73) );
  INVX8 U99 ( .A(n73), .Y(calc_out[62]) );
  CLKINVX8 U100 ( .A(n135), .Y(n76) );
  INVX8 U101 ( .A(n76), .Y(calc_out[116]) );
  BUFX20 U102 ( .A(temp_2_real[14]), .Y(n79) );
  BUFX20 U103 ( .A(temp_3_real[5]), .Y(n93) );
  OAI21X2 U104 ( .A0(rotation[0]), .A1(rotation[1]), .B0(rotation[2]), .Y(N42)
         );
  BUFX20 U105 ( .A(temp_1_real[5]), .Y(n95) );
  AND2X1 U106 ( .A(n33), .B(rotation[2]), .Y(n81) );
  INVX1 U107 ( .A(n81), .Y(n82) );
  INVX1 U108 ( .A(n81), .Y(n83) );
  CLKINVX3 U109 ( .A(n104), .Y(n102) );
  INVX1 U110 ( .A(n100), .Y(n97) );
  INVX1 U111 ( .A(n11), .Y(n90) );
  INVX1 U112 ( .A(n11), .Y(n91) );
  BUFX3 U113 ( .A(n81), .Y(n92) );
  BUFX3 U114 ( .A(n10), .Y(n88) );
  INVXL U115 ( .A(N6), .Y(n104) );
  BUFX20 U116 ( .A(n22), .Y(n89) );
endmodule


module reg1 ( clk, rst_n, data_in_2, reg_datain_flag, data_out_2 );
  input [135:0] data_in_2;
  output [135:0] data_out_2;
  input clk, rst_n, reg_datain_flag;
  wire   reg_flag_mux, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62,
         N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76,
         N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90,
         N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, N124, N125,
         N126, N127, N128, N129, N130, N131, N132, N133, N134, N135, N136,
         N137, N138, N139, N140, N141, N142, N143, N144, N145, N146, N147,
         N148, N149, N150, N151, N152, N153, N154, N155, N156, N157, N158,
         N159, N160, N161, N162, N163, N164, N165, N166, N167, N168, N169,
         N170, N171, N172, N173, N174, N175, N176, N177, N178, N179, N180,
         N181, N182, N183, N184, N185, N186, N187, n146, n148, n149, n150,
         n151, n152, n153, n165, n169, n182, n184, n185, n186, n187, n199,
         n200, n202, n204, n282, n284, n285, n286, n287, n288, n289, n301,
         n305, n318, n320, n321, n322, n323, n335, n336, n338, n340, n418,
         n420, n421, n422, n423, n424, n437, n441, n454, n458, n471, n472,
         n474, n476, n522, n525, n526, n539, n540, n542, n554, n557, n558,
         n559, n560, n573, n577, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n961, n962, n963, n964, n965, n966, n967, n969, n971, n973,
         n974, n975, n976, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
         n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
         n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
         n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
         n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
         n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
         n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
         n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
         n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
         n6, n7, n14, n15, n16, n17, n18, n19, n20, n30, n31, n32, n33, n38,
         n39, n43, n44, n61, n63, n68, n69, n70, n71, n72, n73, n75, n77, n83,
         n84, n85, n86, n87, n89, n90, n91, n92, n93, n95, n96, n97, n98, n100,
         n102, n104, n105, n109, n195, n196, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n958, n959,
         n960, n968, n970, n972, n977, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1235, n1236,
         n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
         n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
         n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
         n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
         n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
         n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
         n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
         n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
         n1317, n1318, n1319, n1320, n1321, n1322, n1323;
  wire   [1:0] counter1;
  wire   [32:0] R0;
  wire   [30:0] R1;
  wire   [32:0] R4;
  wire   [32:0] R5;
  wire   [32:0] R8;
  wire   [32:0] R9;
  wire   [33:0] R12;
  wire   [32:0] R13;
  wire   [1:0] counter2;

  CLKINVX4 U302 ( .A(rst_n), .Y(n961) );
  EDFFXL R11_reg_30_ ( .D(data_in_2[132]), .E(n1248), .CK(clk), .QN(n689) );
  EDFFXL R15_reg_30_ ( .D(data_in_2[132]), .E(n1273), .CK(clk), .QN(n791) );
  EDFFXL R3_reg_30_ ( .D(data_in_2[132]), .E(n1260), .CK(clk), .QN(n859) );
  EDFFXL R7_reg_30_ ( .D(data_in_2[132]), .E(n1288), .CK(clk), .QN(n927) );
  EDFFXL data_out_2_reg_33_ ( .D(N85), .E(n1317), .CK(clk), .Q(data_out_2[33])
         );
  DFFHQXL R12_reg_11_ ( .D(n1221), .CK(clk), .Q(R12[11]) );
  DFFHQXL R8_reg_11_ ( .D(n1220), .CK(clk), .Q(R8[11]) );
  DFFHQXL R4_reg_11_ ( .D(n1219), .CK(clk), .Q(R4[11]) );
  DFFHQXL R0_reg_11_ ( .D(n1218), .CK(clk), .Q(R0[11]) );
  DFFHQXL R13_reg_13_ ( .D(n1217), .CK(clk), .Q(R13[13]) );
  DFFHQXL R9_reg_13_ ( .D(n1216), .CK(clk), .Q(R9[13]) );
  DFFHQXL R5_reg_13_ ( .D(n1215), .CK(clk), .Q(R5[13]) );
  DFFHQXL R1_reg_13_ ( .D(n1214), .CK(clk), .Q(R1[13]) );
  DFFHQXL R12_reg_14_ ( .D(n1213), .CK(clk), .Q(R12[14]) );
  DFFHQXL R8_reg_14_ ( .D(n1212), .CK(clk), .Q(R8[14]) );
  DFFHQXL R4_reg_14_ ( .D(n1211), .CK(clk), .Q(R4[14]) );
  DFFHQXL R0_reg_14_ ( .D(n1210), .CK(clk), .Q(R0[14]) );
  DFFHQXL R13_reg_29_ ( .D(n1209), .CK(clk), .Q(R13[29]) );
  DFFHQXL R9_reg_29_ ( .D(n1208), .CK(clk), .Q(R9[29]) );
  DFFHQXL R5_reg_29_ ( .D(n1207), .CK(clk), .Q(R5[29]) );
  DFFHQXL R1_reg_29_ ( .D(n1206), .CK(clk), .Q(R1[29]) );
  DFFHQXL R13_reg_28_ ( .D(n1204), .CK(clk), .Q(R13[28]) );
  DFFHQXL R9_reg_28_ ( .D(n1203), .CK(clk), .Q(R9[28]) );
  DFFHQXL R5_reg_28_ ( .D(n1202), .CK(clk), .Q(R5[28]) );
  DFFHQXL R1_reg_28_ ( .D(n1201), .CK(clk), .Q(R1[28]) );
  MX2X1 R12_reg_28__U3 ( .A(R12[28]), .B(data_in_2[28]), .S0(n105), .Y(n1200)
         );
  DFFHQXL R12_reg_28_ ( .D(n1200), .CK(clk), .Q(R12[28]) );
  MX2X1 R8_reg_28__U3 ( .A(R8[28]), .B(data_in_2[28]), .S0(n1250), .Y(n1199)
         );
  DFFHQXL R8_reg_28_ ( .D(n1199), .CK(clk), .Q(R8[28]) );
  MX2X1 R4_reg_28__U3 ( .A(R4[28]), .B(data_in_2[28]), .S0(n1283), .Y(n1198)
         );
  DFFHQXL R4_reg_28_ ( .D(n1198), .CK(clk), .Q(R4[28]) );
  MX2X1 R0_reg_28__U3 ( .A(R0[28]), .B(data_in_2[28]), .S0(n1256), .Y(n1197)
         );
  DFFHQXL R0_reg_28_ ( .D(n1197), .CK(clk), .Q(R0[28]) );
  DFFHQXL R12_reg_15_ ( .D(n1196), .CK(clk), .Q(R12[15]) );
  DFFHQXL R8_reg_15_ ( .D(n1195), .CK(clk), .Q(R8[15]) );
  DFFHQXL R4_reg_15_ ( .D(n1194), .CK(clk), .Q(R4[15]) );
  DFFHQXL R0_reg_15_ ( .D(n1193), .CK(clk), .Q(R0[15]) );
  DFFHQXL R13_reg_16_ ( .D(n1192), .CK(clk), .Q(R13[16]) );
  DFFHQXL R9_reg_16_ ( .D(n1191), .CK(clk), .Q(R9[16]) );
  DFFHQXL R5_reg_16_ ( .D(n1190), .CK(clk), .Q(R5[16]) );
  DFFHQXL R1_reg_16_ ( .D(n1189), .CK(clk), .Q(R1[16]) );
  DFFHQXL R12_reg_10_ ( .D(n1185), .CK(clk), .Q(R12[10]) );
  DFFHQXL R4_reg_10_ ( .D(n1184), .CK(clk), .Q(R4[10]) );
  DFFHQXL R12_reg_30_ ( .D(n1183), .CK(clk), .Q(R12[30]) );
  DFFHQXL R8_reg_30_ ( .D(n1182), .CK(clk), .Q(R8[30]) );
  DFFHQXL R4_reg_30_ ( .D(n1181), .CK(clk), .Q(R4[30]) );
  DFFHQXL R0_reg_30_ ( .D(n1180), .CK(clk), .Q(R0[30]) );
  DFFHQXL R12_reg_13_ ( .D(n1179), .CK(clk), .Q(R12[13]) );
  DFFHQXL R8_reg_13_ ( .D(n1178), .CK(clk), .Q(R8[13]) );
  DFFHQXL R4_reg_13_ ( .D(n1177), .CK(clk), .Q(R4[13]) );
  DFFHQXL R0_reg_13_ ( .D(n1176), .CK(clk), .Q(R0[13]) );
  MX2X1 R8_reg_31__U3 ( .A(n77), .B(data_in_2[31]), .S0(n1251), .Y(n1174) );
  DFFHQXL R4_reg_31_ ( .D(n1173), .CK(clk), .Q(R4[31]) );
  DFFHQXL R0_reg_31_ ( .D(n1172), .CK(clk), .Q(R0[31]) );
  DFFHQXL R12_reg_32_ ( .D(n1171), .CK(clk), .Q(R12[32]) );
  DFFHQXL R8_reg_32_ ( .D(n1170), .CK(clk), .Q(R8[32]) );
  DFFHQXL R4_reg_32_ ( .D(n1169), .CK(clk), .Q(R4[32]) );
  DFFHQXL R0_reg_32_ ( .D(n1168), .CK(clk), .Q(R0[32]) );
  DFFHQXL R13_reg_11_ ( .D(n1167), .CK(clk), .Q(R13[11]) );
  DFFHQXL R9_reg_11_ ( .D(n1166), .CK(clk), .Q(R9[11]) );
  DFFHQXL R5_reg_11_ ( .D(n1165), .CK(clk), .Q(R5[11]) );
  MX2X1 R12_reg_27__U3 ( .A(R12[27]), .B(data_in_2[27]), .S0(n105), .Y(n1159)
         );
  DFFHQXL R12_reg_27_ ( .D(n1159), .CK(clk), .Q(R12[27]) );
  MX2X1 R4_reg_27__U3 ( .A(R4[27]), .B(data_in_2[27]), .S0(n1283), .Y(n1158)
         );
  DFFHQXL R4_reg_27_ ( .D(n1158), .CK(clk), .Q(R4[27]) );
  MX2X1 R0_reg_27__U3 ( .A(R0[27]), .B(data_in_2[27]), .S0(n1256), .Y(n1157)
         );
  DFFHQXL R0_reg_27_ ( .D(n1157), .CK(clk), .Q(R0[27]) );
  DFFHQXL R12_reg_29_ ( .D(n1156), .CK(clk), .Q(R12[29]) );
  DFFHQXL R8_reg_29_ ( .D(n1155), .CK(clk), .Q(R8[29]) );
  DFFHQXL R4_reg_29_ ( .D(n1154), .CK(clk), .Q(R4[29]) );
  DFFHQXL R0_reg_29_ ( .D(n1153), .CK(clk), .Q(R0[29]) );
  DFFHQXL R13_reg_14_ ( .D(n1152), .CK(clk), .Q(R13[14]) );
  DFFHQXL R9_reg_14_ ( .D(n1151), .CK(clk), .Q(R9[14]) );
  DFFHQXL R5_reg_14_ ( .D(n1150), .CK(clk), .Q(R5[14]) );
  DFFHQXL R1_reg_14_ ( .D(n1149), .CK(clk), .Q(R1[14]) );
  DFFXL R15_reg_33_ ( .D(n1141), .CK(clk), .Q(n1228), .QN(n788) );
  DFFXL R11_reg_33_ ( .D(n1140), .CK(clk), .Q(n1227), .QN(n686) );
  DFFXL R7_reg_33_ ( .D(n1139), .CK(clk), .Q(n1230), .QN(n924) );
  DFFXL R3_reg_33_ ( .D(n1138), .CK(clk), .Q(n1229), .QN(n856) );
  MX2X1 R15_reg_9__U3 ( .A(n418), .B(data_in_2[111]), .S0(n1271), .Y(n1137) );
  DFFXL R15_reg_9_ ( .D(n1137), .CK(clk), .Q(n418), .QN(n812) );
  MX2X1 R11_reg_9__U3 ( .A(n554), .B(data_in_2[111]), .S0(n1247), .Y(n1136) );
  DFFXL R11_reg_9_ ( .D(n1136), .CK(clk), .Q(n554), .QN(n710) );
  MX2X1 R7_reg_9__U3 ( .A(n146), .B(data_in_2[111]), .S0(n1286), .Y(n1135) );
  DFFXL R7_reg_9_ ( .D(n1135), .CK(clk), .Q(n146), .QN(n948) );
  MX2X1 R3_reg_9__U3 ( .A(n282), .B(data_in_2[111]), .S0(n1261), .Y(n1134) );
  DFFXL R3_reg_9_ ( .D(n1134), .CK(clk), .Q(n282), .QN(n880) );
  MX2X1 R15_reg_12__U3 ( .A(n421), .B(data_in_2[114]), .S0(n1272), .Y(n1133)
         );
  DFFXL R15_reg_12_ ( .D(n1133), .CK(clk), .Q(n421), .QN(n809) );
  MX2X1 R11_reg_12__U3 ( .A(n557), .B(data_in_2[114]), .S0(n1247), .Y(n1132)
         );
  DFFXL R11_reg_12_ ( .D(n1132), .CK(clk), .Q(n557), .QN(n707) );
  MX2X1 R7_reg_12__U3 ( .A(n149), .B(data_in_2[114]), .S0(n1288), .Y(n1131) );
  DFFXL R7_reg_12_ ( .D(n1131), .CK(clk), .Q(n149), .QN(n945) );
  MX2X1 R3_reg_12__U3 ( .A(n285), .B(data_in_2[114]), .S0(n1261), .Y(n1130) );
  DFFXL R3_reg_12_ ( .D(n1130), .CK(clk), .Q(n285), .QN(n877) );
  DFFXL R14_reg_11_ ( .D(n1129), .CK(clk), .Q(n454), .QN(n776) );
  MX2X1 R10_reg_11__U3 ( .A(n522), .B(data_in_2[79]), .S0(n1244), .Y(n1128) );
  DFFXL R10_reg_11_ ( .D(n1128), .CK(clk), .Q(n522), .QN(n742) );
  MX2X1 R6_reg_11__U3 ( .A(n182), .B(data_in_2[79]), .S0(n1287), .Y(n1127) );
  DFFXL R6_reg_11_ ( .D(n1127), .CK(clk), .Q(n182), .QN(n912) );
  MX2X1 R2_reg_11__U3 ( .A(n318), .B(data_in_2[79]), .S0(n1260), .Y(n1126) );
  DFFXL R2_reg_11_ ( .D(n1126), .CK(clk), .Q(n318), .QN(n844) );
  DFFXL R15_reg_31_ ( .D(n1125), .CK(clk), .Q(n1236), .QN(n790) );
  DFFXL R11_reg_31_ ( .D(n1124), .CK(clk), .Q(n1235), .QN(n688) );
  DFFXL R7_reg_31_ ( .D(n1123), .CK(clk), .Q(n1238), .QN(n926) );
  DFFXL R3_reg_31_ ( .D(n1122), .CK(clk), .Q(n1237), .QN(n858) );
  DFFXL R14_reg_28_ ( .D(n1121), .CK(clk), .Q(n471), .QN(n759) );
  MX2X1 R10_reg_28__U3 ( .A(n539), .B(data_in_2[96]), .S0(n1246), .Y(n1120) );
  DFFXL R10_reg_28_ ( .D(n1120), .CK(clk), .Q(n539), .QN(n725) );
  MX2X1 R6_reg_28__U3 ( .A(n199), .B(data_in_2[96]), .S0(n1286), .Y(n1119) );
  DFFXL R6_reg_28_ ( .D(n1119), .CK(clk), .Q(n199), .QN(n895) );
  MX2X1 R2_reg_28__U3 ( .A(n335), .B(data_in_2[96]), .S0(n1259), .Y(n1118) );
  DFFXL R2_reg_28_ ( .D(n1118), .CK(clk), .Q(n335), .QN(n827) );
  DFFXL R15_reg_28_ ( .D(n1117), .CK(clk), .Q(n437), .QN(n793) );
  DFFXL R11_reg_28_ ( .D(n977), .CK(clk), .Q(n573), .QN(n691) );
  DFFXL R7_reg_28_ ( .D(n972), .CK(clk), .Q(n165), .QN(n929) );
  DFFXL R3_reg_28_ ( .D(n970), .CK(clk), .Q(n301), .QN(n861) );
  MX2X1 R15_reg_15__U3 ( .A(n424), .B(data_in_2[117]), .S0(n1272), .Y(n968) );
  DFFXL R15_reg_15_ ( .D(n968), .CK(clk), .Q(n424), .QN(n806) );
  MX2X1 R11_reg_15__U3 ( .A(n560), .B(data_in_2[117]), .S0(n1247), .Y(n960) );
  DFFXL R11_reg_15_ ( .D(n960), .CK(clk), .Q(n560), .QN(n704) );
  MX2X1 R7_reg_15__U3 ( .A(n152), .B(data_in_2[117]), .S0(n1288), .Y(n959) );
  DFFXL R7_reg_15_ ( .D(n959), .CK(clk), .Q(n152), .QN(n942) );
  MX2X1 R3_reg_15__U3 ( .A(n288), .B(data_in_2[117]), .S0(n1261), .Y(n958) );
  DFFXL R3_reg_15_ ( .D(n958), .CK(clk), .Q(n288), .QN(n874) );
  DFFXL R6_reg_16_ ( .D(n685), .CK(clk), .Q(n187), .QN(n907) );
  DFFXL R2_reg_16_ ( .D(n684), .CK(clk), .Q(n323), .QN(n839) );
  DFFXL R6_reg_13_ ( .D(n683), .CK(clk), .Q(n184), .QN(n910) );
  DFFXL R2_reg_13_ ( .D(n682), .CK(clk), .Q(n320), .QN(n842) );
  MX2X1 R14_reg_30__U3 ( .A(n1224), .B(data_in_2[98]), .S0(n1275), .Y(n681) );
  DFFXL R14_reg_30_ ( .D(n681), .CK(clk), .Q(n1224), .QN(n757) );
  MX2X1 R10_reg_30__U3 ( .A(n1223), .B(data_in_2[98]), .S0(n1246), .Y(n680) );
  DFFXL R10_reg_30_ ( .D(n680), .CK(clk), .Q(n1223), .QN(n723) );
  MX2X1 R6_reg_30__U3 ( .A(n1226), .B(data_in_2[98]), .S0(n1286), .Y(n679) );
  DFFXL R6_reg_30_ ( .D(n679), .CK(clk), .Q(n1226), .QN(n893) );
  MX2X1 R2_reg_30__U3 ( .A(n1225), .B(data_in_2[98]), .S0(n1259), .Y(n678) );
  DFFXL R2_reg_30_ ( .D(n678), .CK(clk), .Q(n1225), .QN(n825) );
  DFFXL R14_reg_32_ ( .D(n677), .CK(clk), .Q(n1240), .QN(n755) );
  DFFXL R10_reg_32_ ( .D(n676), .CK(clk), .Q(n1239), .QN(n721) );
  DFFXL R6_reg_32_ ( .D(n675), .CK(clk), .Q(n1242), .QN(n891) );
  DFFXL R2_reg_32_ ( .D(n674), .CK(clk), .Q(n1241), .QN(n823) );
  DFFXL R15_reg_13_ ( .D(n673), .CK(clk), .Q(n422), .QN(n808) );
  DFFXL R11_reg_13_ ( .D(n672), .CK(clk), .Q(n558), .QN(n706) );
  DFFXL R7_reg_13_ ( .D(n671), .CK(clk), .Q(n150), .QN(n944) );
  DFFXL R3_reg_13_ ( .D(n670), .CK(clk), .Q(n286), .QN(n876) );
  DFFXL R14_reg_15_ ( .D(n669), .CK(clk), .Q(n458), .QN(n772) );
  MX2X1 R10_reg_15__U3 ( .A(n526), .B(data_in_2[83]), .S0(n1245), .Y(n668) );
  DFFXL R10_reg_15_ ( .D(n668), .CK(clk), .Q(n526), .QN(n738) );
  MX2X1 R6_reg_15__U3 ( .A(n186), .B(data_in_2[83]), .S0(n1287), .Y(n667) );
  DFFXL R6_reg_15_ ( .D(n667), .CK(clk), .Q(n186), .QN(n908) );
  MX2X1 R2_reg_15__U3 ( .A(n322), .B(data_in_2[83]), .S0(n1260), .Y(n666) );
  DFFXL R2_reg_15_ ( .D(n666), .CK(clk), .Q(n322), .QN(n840) );
  MX2X1 R10_reg_14__U3 ( .A(n525), .B(data_in_2[82]), .S0(n1245), .Y(n665) );
  DFFXL R10_reg_14_ ( .D(n665), .CK(clk), .Q(n525), .QN(n739) );
  MX2X1 R6_reg_14__U3 ( .A(n185), .B(data_in_2[82]), .S0(n1287), .Y(n664) );
  DFFXL R6_reg_14_ ( .D(n664), .CK(clk), .Q(n185), .QN(n909) );
  MX2X1 R2_reg_14__U3 ( .A(n321), .B(data_in_2[82]), .S0(n1260), .Y(n663) );
  DFFXL R2_reg_14_ ( .D(n663), .CK(clk), .Q(n321), .QN(n841) );
  DFFXL R14_reg_31_ ( .D(n662), .CK(clk), .Q(n474), .QN(n756) );
  DFFXL R10_reg_31_ ( .D(n661), .CK(clk), .Q(n542), .QN(n722) );
  DFFXL R6_reg_31_ ( .D(n660), .CK(clk), .Q(n202), .QN(n892) );
  DFFXL R2_reg_31_ ( .D(n659), .CK(clk), .Q(n338), .QN(n824) );
  MX2X1 R14_reg_29__U3 ( .A(n472), .B(data_in_2[97]), .S0(n1275), .Y(n658) );
  DFFXL R14_reg_29_ ( .D(n658), .CK(clk), .Q(n472), .QN(n758) );
  MX2X1 R10_reg_29__U3 ( .A(n540), .B(data_in_2[97]), .S0(n1246), .Y(n657) );
  DFFXL R10_reg_29_ ( .D(n657), .CK(clk), .Q(n540), .QN(n724) );
  MX2X1 R6_reg_29__U3 ( .A(n200), .B(data_in_2[97]), .S0(n1286), .Y(n656) );
  DFFXL R6_reg_29_ ( .D(n656), .CK(clk), .Q(n200), .QN(n894) );
  MX2X1 R2_reg_29__U3 ( .A(n336), .B(data_in_2[97]), .S0(n1259), .Y(n655) );
  DFFXL R2_reg_29_ ( .D(n655), .CK(clk), .Q(n336), .QN(n826) );
  DFFXL R15_reg_32_ ( .D(n654), .CK(clk), .Q(n441), .QN(n789) );
  DFFXL R11_reg_32_ ( .D(n653), .CK(clk), .Q(n577), .QN(n687) );
  DFFXL R7_reg_32_ ( .D(n652), .CK(clk), .Q(n169), .QN(n925) );
  DFFXL R3_reg_32_ ( .D(n651), .CK(clk), .Q(n305), .QN(n857) );
  DFFXL R7_reg_16_ ( .D(n650), .CK(clk), .Q(n153), .QN(n941) );
  DFFXL R3_reg_16_ ( .D(n649), .CK(clk), .Q(n289), .QN(n873) );
  DFFXL R14_reg_33_ ( .D(n648), .CK(clk), .Q(n476), .QN(n754) );
  DFFXL R6_reg_33_ ( .D(n647), .CK(clk), .Q(n204), .QN(n890) );
  DFFXL R2_reg_33_ ( .D(n646), .CK(clk), .Q(n340), .QN(n822) );
  MX2X1 R15_reg_11__U3 ( .A(n420), .B(data_in_2[113]), .S0(n1271), .Y(n645) );
  DFFXL R15_reg_11_ ( .D(n645), .CK(clk), .Q(n420), .QN(n810) );
  MX2X1 R7_reg_11__U3 ( .A(n148), .B(data_in_2[113]), .S0(n1288), .Y(n644) );
  DFFXL R7_reg_11_ ( .D(n644), .CK(clk), .Q(n148), .QN(n946) );
  MX2X1 R3_reg_11__U3 ( .A(n284), .B(data_in_2[113]), .S0(n1261), .Y(n643) );
  DFFXL R3_reg_11_ ( .D(n643), .CK(clk), .Q(n284), .QN(n878) );
  MX2X1 R15_reg_14__U3 ( .A(n423), .B(data_in_2[116]), .S0(n1272), .Y(n642) );
  DFFXL R15_reg_14_ ( .D(n642), .CK(clk), .Q(n423), .QN(n807) );
  MX2X1 R11_reg_14__U3 ( .A(n559), .B(data_in_2[116]), .S0(n1247), .Y(n641) );
  DFFXL R11_reg_14_ ( .D(n641), .CK(clk), .Q(n559), .QN(n705) );
  MX2X1 R7_reg_14__U3 ( .A(n151), .B(data_in_2[116]), .S0(n1288), .Y(n640) );
  DFFXL R7_reg_14_ ( .D(n640), .CK(clk), .Q(n151), .QN(n943) );
  MX2X1 R3_reg_14__U3 ( .A(n287), .B(data_in_2[116]), .S0(n1261), .Y(n639) );
  DFFXL R3_reg_14_ ( .D(n639), .CK(clk), .Q(n287), .QN(n875) );
  EDFFX1 data_out_2_reg_134_ ( .D(N186), .E(n1315), .CK(clk), .Q(
        data_out_2[134]) );
  EDFFX1 data_out_2_reg_133_ ( .D(N185), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[133]) );
  EDFFX1 data_out_2_reg_132_ ( .D(N184), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[132]) );
  EDFFX1 data_out_2_reg_131_ ( .D(N183), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[131]) );
  EDFFX1 data_out_2_reg_130_ ( .D(N182), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[130]) );
  EDFFX1 data_out_2_reg_129_ ( .D(N181), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[129]) );
  EDFFX1 data_out_2_reg_128_ ( .D(N180), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[128]) );
  EDFFX1 data_out_2_reg_127_ ( .D(N179), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[127]) );
  EDFFX1 data_out_2_reg_126_ ( .D(N178), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[126]) );
  EDFFX1 data_out_2_reg_125_ ( .D(N177), .E(n1317), .CK(clk), .Q(
        data_out_2[125]) );
  EDFFX1 data_out_2_reg_124_ ( .D(N176), .E(n1315), .CK(clk), .Q(
        data_out_2[124]) );
  EDFFX1 data_out_2_reg_123_ ( .D(N175), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[123]) );
  EDFFX1 data_out_2_reg_122_ ( .D(N174), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[122]) );
  EDFFX1 data_out_2_reg_121_ ( .D(N173), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[121]) );
  EDFFX1 data_out_2_reg_120_ ( .D(N172), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[120]) );
  EDFFX1 data_out_2_reg_117_ ( .D(N169), .E(n1317), .CK(clk), .Q(
        data_out_2[117]) );
  EDFFX1 data_out_2_reg_116_ ( .D(N168), .E(n1315), .CK(clk), .Q(
        data_out_2[116]) );
  EDFFX1 data_out_2_reg_115_ ( .D(N167), .E(n1317), .CK(clk), .Q(
        data_out_2[115]) );
  EDFFX1 data_out_2_reg_114_ ( .D(N166), .E(n1316), .CK(clk), .Q(
        data_out_2[114]) );
  EDFFX1 data_out_2_reg_113_ ( .D(N165), .E(n1317), .CK(clk), .Q(
        data_out_2[113]) );
  EDFFX1 data_out_2_reg_112_ ( .D(N164), .E(n1315), .CK(clk), .Q(
        data_out_2[112]) );
  EDFFX1 data_out_2_reg_111_ ( .D(N163), .E(n1316), .CK(clk), .Q(
        data_out_2[111]) );
  EDFFX1 data_out_2_reg_110_ ( .D(N162), .E(n1316), .CK(clk), .Q(
        data_out_2[110]) );
  EDFFX1 data_out_2_reg_109_ ( .D(N161), .E(n1317), .CK(clk), .Q(
        data_out_2[109]) );
  EDFFX1 data_out_2_reg_108_ ( .D(N160), .E(n1315), .CK(clk), .Q(
        data_out_2[108]) );
  EDFFX1 data_out_2_reg_107_ ( .D(N159), .E(n1315), .CK(clk), .Q(
        data_out_2[107]) );
  EDFFX1 data_out_2_reg_106_ ( .D(N158), .E(n1316), .CK(clk), .Q(
        data_out_2[106]) );
  EDFFX1 data_out_2_reg_105_ ( .D(N157), .E(n1317), .CK(clk), .Q(
        data_out_2[105]) );
  EDFFX1 data_out_2_reg_104_ ( .D(N156), .E(n1315), .CK(clk), .Q(
        data_out_2[104]) );
  EDFFX1 data_out_2_reg_103_ ( .D(N155), .E(n1316), .CK(clk), .Q(
        data_out_2[103]) );
  EDFFX1 data_out_2_reg_100_ ( .D(N152), .E(n1317), .CK(clk), .Q(
        data_out_2[100]) );
  EDFFX1 data_out_2_reg_99_ ( .D(N151), .E(n1316), .CK(clk), .Q(data_out_2[99]) );
  EDFFX1 data_out_2_reg_98_ ( .D(N150), .E(n1315), .CK(clk), .Q(data_out_2[98]) );
  EDFFX1 data_out_2_reg_97_ ( .D(N149), .E(n1315), .CK(clk), .Q(data_out_2[97]) );
  EDFFX1 data_out_2_reg_96_ ( .D(N148), .E(n1315), .CK(clk), .Q(data_out_2[96]) );
  EDFFX1 data_out_2_reg_95_ ( .D(N147), .E(n1315), .CK(clk), .Q(data_out_2[95]) );
  EDFFX1 data_out_2_reg_94_ ( .D(N146), .E(n1315), .CK(clk), .Q(data_out_2[94]) );
  EDFFX1 data_out_2_reg_93_ ( .D(N145), .E(n1315), .CK(clk), .Q(data_out_2[93]) );
  EDFFX1 data_out_2_reg_92_ ( .D(N144), .E(n1315), .CK(clk), .Q(data_out_2[92]) );
  EDFFX1 data_out_2_reg_91_ ( .D(N143), .E(n1315), .CK(clk), .Q(data_out_2[91]) );
  EDFFX1 data_out_2_reg_90_ ( .D(N142), .E(n1315), .CK(clk), .Q(data_out_2[90]) );
  EDFFX1 data_out_2_reg_89_ ( .D(N141), .E(n1315), .CK(clk), .Q(data_out_2[89]) );
  EDFFX1 data_out_2_reg_88_ ( .D(N140), .E(n1315), .CK(clk), .Q(data_out_2[88]) );
  EDFFX1 data_out_2_reg_87_ ( .D(N139), .E(n1315), .CK(clk), .Q(data_out_2[87]) );
  EDFFX1 data_out_2_reg_86_ ( .D(N138), .E(n1315), .CK(clk), .Q(data_out_2[86]) );
  EDFFX1 data_out_2_reg_83_ ( .D(N135), .E(n1315), .CK(clk), .Q(data_out_2[83]) );
  EDFFX1 data_out_2_reg_82_ ( .D(N134), .E(n1315), .CK(clk), .Q(data_out_2[82]) );
  EDFFX1 data_out_2_reg_81_ ( .D(N133), .E(n1315), .CK(clk), .Q(data_out_2[81]) );
  EDFFX1 data_out_2_reg_80_ ( .D(N132), .E(n1315), .CK(clk), .Q(data_out_2[80]) );
  EDFFX1 data_out_2_reg_79_ ( .D(N131), .E(n1315), .CK(clk), .Q(data_out_2[79]) );
  EDFFX1 data_out_2_reg_78_ ( .D(N130), .E(n1315), .CK(clk), .Q(data_out_2[78]) );
  EDFFX1 data_out_2_reg_77_ ( .D(N129), .E(n1317), .CK(clk), .Q(data_out_2[77]) );
  EDFFX1 data_out_2_reg_76_ ( .D(N128), .E(n1316), .CK(clk), .Q(data_out_2[76]) );
  EDFFX1 data_out_2_reg_75_ ( .D(N127), .E(n1315), .CK(clk), .Q(data_out_2[75]) );
  EDFFX1 data_out_2_reg_74_ ( .D(N126), .E(n1317), .CK(clk), .Q(data_out_2[74]) );
  EDFFX1 data_out_2_reg_73_ ( .D(N125), .E(n1317), .CK(clk), .Q(data_out_2[73]) );
  EDFFX1 data_out_2_reg_72_ ( .D(N124), .E(n1315), .CK(clk), .Q(data_out_2[72]) );
  EDFFX1 data_out_2_reg_71_ ( .D(N123), .E(n1317), .CK(clk), .Q(data_out_2[71]) );
  EDFFX1 data_out_2_reg_70_ ( .D(N122), .E(n1315), .CK(clk), .Q(data_out_2[70]) );
  EDFFX1 data_out_2_reg_69_ ( .D(N121), .E(n1316), .CK(clk), .Q(data_out_2[69]) );
  EDFFX1 data_out_2_reg_66_ ( .D(N118), .E(n1315), .CK(clk), .Q(data_out_2[66]) );
  EDFFX1 data_out_2_reg_65_ ( .D(N117), .E(n1316), .CK(clk), .Q(data_out_2[65]) );
  EDFFX1 data_out_2_reg_64_ ( .D(N116), .E(n1316), .CK(clk), .Q(data_out_2[64]) );
  EDFFX1 data_out_2_reg_63_ ( .D(N115), .E(n1317), .CK(clk), .Q(data_out_2[63]) );
  EDFFX1 data_out_2_reg_62_ ( .D(N114), .E(n1315), .CK(clk), .Q(data_out_2[62]) );
  EDFFX1 data_out_2_reg_61_ ( .D(N113), .E(n1316), .CK(clk), .Q(data_out_2[61]) );
  EDFFX1 data_out_2_reg_60_ ( .D(N112), .E(n1316), .CK(clk), .Q(data_out_2[60]) );
  EDFFX1 data_out_2_reg_59_ ( .D(N111), .E(n1316), .CK(clk), .Q(data_out_2[59]) );
  EDFFX1 data_out_2_reg_58_ ( .D(N110), .E(n1316), .CK(clk), .Q(data_out_2[58]) );
  EDFFX1 data_out_2_reg_57_ ( .D(N109), .E(n1316), .CK(clk), .Q(data_out_2[57]) );
  EDFFX1 data_out_2_reg_56_ ( .D(N108), .E(n1316), .CK(clk), .Q(data_out_2[56]) );
  EDFFX1 data_out_2_reg_55_ ( .D(N107), .E(n1316), .CK(clk), .Q(data_out_2[55]) );
  EDFFX1 data_out_2_reg_54_ ( .D(N106), .E(n1316), .CK(clk), .Q(data_out_2[54]) );
  EDFFX1 data_out_2_reg_53_ ( .D(N105), .E(n1316), .CK(clk), .Q(data_out_2[53]) );
  EDFFX1 data_out_2_reg_52_ ( .D(N104), .E(n1316), .CK(clk), .Q(data_out_2[52]) );
  EDFFX1 data_out_2_reg_49_ ( .D(N101), .E(n1316), .CK(clk), .Q(data_out_2[49]) );
  EDFFX1 data_out_2_reg_48_ ( .D(N100), .E(n1316), .CK(clk), .Q(data_out_2[48]) );
  EDFFX1 data_out_2_reg_47_ ( .D(N99), .E(n1316), .CK(clk), .Q(data_out_2[47])
         );
  EDFFX1 data_out_2_reg_46_ ( .D(N98), .E(n1316), .CK(clk), .Q(data_out_2[46])
         );
  EDFFX1 data_out_2_reg_45_ ( .D(N97), .E(n1316), .CK(clk), .Q(data_out_2[45])
         );
  EDFFX1 data_out_2_reg_44_ ( .D(N96), .E(n1316), .CK(clk), .Q(data_out_2[44])
         );
  EDFFX1 data_out_2_reg_43_ ( .D(N95), .E(n1316), .CK(clk), .Q(data_out_2[43])
         );
  EDFFX1 data_out_2_reg_42_ ( .D(N94), .E(n1316), .CK(clk), .Q(data_out_2[42])
         );
  EDFFX1 data_out_2_reg_41_ ( .D(N93), .E(n1316), .CK(clk), .Q(data_out_2[41])
         );
  EDFFX1 data_out_2_reg_40_ ( .D(N92), .E(n1316), .CK(clk), .Q(data_out_2[40])
         );
  EDFFX1 data_out_2_reg_39_ ( .D(N91), .E(n1317), .CK(clk), .Q(data_out_2[39])
         );
  EDFFX1 data_out_2_reg_38_ ( .D(N90), .E(n1317), .CK(clk), .Q(data_out_2[38])
         );
  EDFFX1 data_out_2_reg_37_ ( .D(N89), .E(n1317), .CK(clk), .Q(data_out_2[37])
         );
  EDFFX1 data_out_2_reg_36_ ( .D(N88), .E(n1317), .CK(clk), .Q(data_out_2[36])
         );
  EDFFX1 data_out_2_reg_35_ ( .D(N87), .E(n1317), .CK(clk), .Q(data_out_2[35])
         );
  EDFFX1 data_out_2_reg_119_ ( .D(N171), .E(n1317), .CK(clk), .Q(
        data_out_2[119]) );
  EDFFX1 data_out_2_reg_102_ ( .D(N154), .E(n1315), .CK(clk), .Q(
        data_out_2[102]) );
  EDFFX1 data_out_2_reg_85_ ( .D(N137), .E(n1315), .CK(clk), .Q(data_out_2[85]) );
  EDFFX1 data_out_2_reg_68_ ( .D(N120), .E(n1317), .CK(clk), .Q(data_out_2[68]) );
  EDFFX1 data_out_2_reg_51_ ( .D(N103), .E(n1316), .CK(clk), .Q(data_out_2[51]) );
  EDFFX1 data_out_2_reg_34_ ( .D(N86), .E(n1317), .CK(clk), .Q(data_out_2[34])
         );
  EDFFX1 R10_reg_24_ ( .D(data_in_2[92]), .E(n1245), .CK(clk), .QN(n729) );
  EDFFX1 R10_reg_22_ ( .D(data_in_2[90]), .E(n1245), .CK(clk), .QN(n731) );
  EDFFX1 R10_reg_20_ ( .D(data_in_2[88]), .E(n1245), .CK(clk), .QN(n733) );
  EDFFXL R10_reg_19_ ( .D(data_in_2[87]), .E(n1245), .CK(clk), .QN(n734) );
  EDFFXL R10_reg_18_ ( .D(data_in_2[86]), .E(n1245), .CK(clk), .QN(n735) );
  EDFFX1 R10_reg_10_ ( .D(data_in_2[78]), .E(n1244), .CK(clk), .QN(n743) );
  EDFFX1 R10_reg_9_ ( .D(data_in_2[77]), .E(n1244), .CK(clk), .QN(n744) );
  EDFFX1 R10_reg_6_ ( .D(data_in_2[74]), .E(n1244), .CK(clk), .QN(n747) );
  EDFFX1 R10_reg_3_ ( .D(data_in_2[71]), .E(n1244), .CK(clk), .QN(n750) );
  EDFFX1 R10_reg_2_ ( .D(data_in_2[70]), .E(n1244), .CK(clk), .QN(n751) );
  EDFFXL R10_reg_1_ ( .D(data_in_2[69]), .E(n1243), .CK(clk), .QN(n752) );
  EDFFX1 R10_reg_0_ ( .D(data_in_2[68]), .E(n1243), .CK(clk), .QN(n753) );
  EDFFX1 R14_reg_24_ ( .D(data_in_2[92]), .E(n1275), .CK(clk), .QN(n763) );
  EDFFX1 R14_reg_20_ ( .D(data_in_2[88]), .E(n1278), .CK(clk), .QN(n767) );
  EDFFXL R14_reg_19_ ( .D(data_in_2[87]), .E(n1278), .CK(clk), .QN(n768) );
  EDFFXL R14_reg_18_ ( .D(data_in_2[86]), .E(n1272), .CK(clk), .QN(n769) );
  EDFFX1 R14_reg_17_ ( .D(data_in_2[85]), .E(n1276), .CK(clk), .QN(n770) );
  EDFFX1 R14_reg_10_ ( .D(data_in_2[78]), .E(n1274), .CK(clk), .QN(n777) );
  EDFFX1 R14_reg_9_ ( .D(data_in_2[77]), .E(n1274), .CK(clk), .QN(n778) );
  EDFFX1 R14_reg_6_ ( .D(data_in_2[74]), .E(n1274), .CK(clk), .QN(n781) );
  EDFFX1 R14_reg_3_ ( .D(data_in_2[71]), .E(n1274), .CK(clk), .QN(n784) );
  EDFFX1 R14_reg_2_ ( .D(data_in_2[70]), .E(n1274), .CK(clk), .QN(n785) );
  EDFFXL R14_reg_1_ ( .D(data_in_2[69]), .E(n1273), .CK(clk), .QN(n786) );
  EDFFX1 R14_reg_0_ ( .D(data_in_2[68]), .E(n1273), .CK(clk), .QN(n787) );
  EDFFX1 R2_reg_24_ ( .D(data_in_2[92]), .E(n1259), .CK(clk), .QN(n831) );
  EDFFX1 R2_reg_22_ ( .D(data_in_2[90]), .E(n1259), .CK(clk), .QN(n833) );
  EDFFX1 R2_reg_20_ ( .D(data_in_2[88]), .E(n1259), .CK(clk), .QN(n835) );
  EDFFXL R2_reg_19_ ( .D(data_in_2[87]), .E(n1259), .CK(clk), .QN(n836) );
  EDFFXL R2_reg_18_ ( .D(data_in_2[86]), .E(n1259), .CK(clk), .QN(n837) );
  EDFFX1 R2_reg_17_ ( .D(data_in_2[85]), .E(n1259), .CK(clk), .QN(n838) );
  EDFFX1 R2_reg_10_ ( .D(data_in_2[78]), .E(n1260), .CK(clk), .QN(n845) );
  EDFFX1 R2_reg_9_ ( .D(data_in_2[77]), .E(n1260), .CK(clk), .QN(n846) );
  EDFFX1 R2_reg_6_ ( .D(data_in_2[74]), .E(n1260), .CK(clk), .QN(n849) );
  EDFFX1 R2_reg_3_ ( .D(data_in_2[71]), .E(n1260), .CK(clk), .QN(n852) );
  EDFFX1 R2_reg_2_ ( .D(data_in_2[70]), .E(n1260), .CK(clk), .QN(n853) );
  EDFFXL R2_reg_1_ ( .D(data_in_2[69]), .E(n1260), .CK(clk), .QN(n854) );
  EDFFX1 R2_reg_0_ ( .D(data_in_2[68]), .E(n1260), .CK(clk), .QN(n855) );
  EDFFXL R6_reg_27_ ( .D(data_in_2[95]), .E(n1286), .CK(clk), .QN(n896) );
  EDFFXL R6_reg_26_ ( .D(data_in_2[94]), .E(n1286), .CK(clk), .QN(n897) );
  EDFFXL R6_reg_25_ ( .D(data_in_2[93]), .E(n1286), .CK(clk), .QN(n898) );
  EDFFXL R6_reg_24_ ( .D(data_in_2[92]), .E(n1286), .CK(clk), .QN(n899) );
  EDFFXL R6_reg_23_ ( .D(data_in_2[91]), .E(n1286), .CK(clk), .QN(n900) );
  EDFFXL R6_reg_22_ ( .D(data_in_2[90]), .E(n1286), .CK(clk), .QN(n901) );
  EDFFXL R6_reg_21_ ( .D(data_in_2[89]), .E(n1286), .CK(clk), .QN(n902) );
  EDFFXL R6_reg_20_ ( .D(data_in_2[88]), .E(n1286), .CK(clk), .QN(n903) );
  EDFFXL R6_reg_19_ ( .D(data_in_2[87]), .E(n1286), .CK(clk), .QN(n904) );
  EDFFX1 R6_reg_18_ ( .D(data_in_2[86]), .E(n1287), .CK(clk), .QN(n905) );
  EDFFX1 R6_reg_17_ ( .D(data_in_2[85]), .E(n1287), .CK(clk), .QN(n906) );
  EDFFXL R6_reg_12_ ( .D(data_in_2[80]), .E(n1287), .CK(clk), .QN(n911) );
  EDFFXL R6_reg_10_ ( .D(data_in_2[78]), .E(n1287), .CK(clk), .QN(n913) );
  EDFFXL R6_reg_9_ ( .D(data_in_2[77]), .E(n1287), .CK(clk), .QN(n914) );
  EDFFXL R6_reg_8_ ( .D(data_in_2[76]), .E(n1287), .CK(clk), .QN(n915) );
  EDFFXL R6_reg_7_ ( .D(data_in_2[75]), .E(n1287), .CK(clk), .QN(n916) );
  EDFFXL R6_reg_6_ ( .D(data_in_2[74]), .E(n1287), .CK(clk), .QN(n917) );
  EDFFXL R6_reg_5_ ( .D(data_in_2[73]), .E(n1287), .CK(clk), .QN(n918) );
  EDFFXL R6_reg_4_ ( .D(data_in_2[72]), .E(n1287), .CK(clk), .QN(n919) );
  EDFFXL R6_reg_3_ ( .D(data_in_2[71]), .E(n1287), .CK(clk), .QN(n920) );
  EDFFXL R6_reg_2_ ( .D(data_in_2[70]), .E(n1287), .CK(clk), .QN(n921) );
  EDFFXL R6_reg_1_ ( .D(data_in_2[69]), .E(n1287), .CK(clk), .QN(n922) );
  EDFFX1 R6_reg_0_ ( .D(data_in_2[68]), .E(n1287), .CK(clk), .QN(n923) );
  EDFFX1 R11_reg_25_ ( .D(data_in_2[127]), .E(n109), .CK(clk), .QN(n694) );
  EDFFX1 R11_reg_24_ ( .D(data_in_2[126]), .E(n109), .CK(clk), .QN(n695) );
  EDFFX1 R11_reg_22_ ( .D(data_in_2[124]), .E(n109), .CK(clk), .QN(n697) );
  EDFFXL R11_reg_19_ ( .D(data_in_2[121]), .E(n109), .CK(clk), .QN(n700) );
  EDFFXL R11_reg_18_ ( .D(data_in_2[120]), .E(n109), .CK(clk), .QN(n701) );
  EDFFX1 R11_reg_8_ ( .D(data_in_2[110]), .E(n1247), .CK(clk), .QN(n711) );
  EDFFXL R11_reg_3_ ( .D(data_in_2[105]), .E(n1246), .CK(clk), .QN(n716) );
  EDFFXL R11_reg_2_ ( .D(data_in_2[104]), .E(n1246), .CK(clk), .QN(n717) );
  EDFFX1 R15_reg_25_ ( .D(data_in_2[127]), .E(n1273), .CK(clk), .QN(n796) );
  EDFFX1 R15_reg_24_ ( .D(data_in_2[126]), .E(n1273), .CK(clk), .QN(n797) );
  EDFFX1 R15_reg_22_ ( .D(data_in_2[124]), .E(n1272), .CK(clk), .QN(n799) );
  EDFFXL R15_reg_19_ ( .D(data_in_2[121]), .E(n1272), .CK(clk), .QN(n802) );
  EDFFXL R15_reg_18_ ( .D(data_in_2[120]), .E(n1272), .CK(clk), .QN(n803) );
  EDFFX1 R15_reg_17_ ( .D(data_in_2[119]), .E(n1272), .CK(clk), .QN(n804) );
  EDFFX1 R15_reg_8_ ( .D(data_in_2[110]), .E(n1271), .CK(clk), .QN(n813) );
  EDFFXL R15_reg_3_ ( .D(data_in_2[105]), .E(n1271), .CK(clk), .QN(n818) );
  EDFFXL R15_reg_2_ ( .D(data_in_2[104]), .E(n1271), .CK(clk), .QN(n819) );
  EDFFX1 R15_reg_1_ ( .D(data_in_2[103]), .E(n1271), .CK(clk), .QN(n820) );
  EDFFX1 R15_reg_0_ ( .D(data_in_2[102]), .E(n1271), .CK(clk), .QN(n821) );
  EDFFX1 R3_reg_25_ ( .D(data_in_2[127]), .E(n1261), .CK(clk), .QN(n864) );
  EDFFX1 R3_reg_24_ ( .D(data_in_2[126]), .E(n1261), .CK(clk), .QN(n865) );
  EDFFX1 R3_reg_22_ ( .D(data_in_2[124]), .E(n1261), .CK(clk), .QN(n867) );
  EDFFXL R3_reg_19_ ( .D(data_in_2[121]), .E(n1261), .CK(clk), .QN(n870) );
  EDFFXL R3_reg_18_ ( .D(data_in_2[120]), .E(n1261), .CK(clk), .QN(n871) );
  EDFFX1 R3_reg_17_ ( .D(data_in_2[119]), .E(n1261), .CK(clk), .QN(n872) );
  EDFFX1 R3_reg_8_ ( .D(data_in_2[110]), .E(n1261), .CK(clk), .QN(n881) );
  EDFFXL R3_reg_3_ ( .D(data_in_2[105]), .E(n1261), .CK(clk), .QN(n886) );
  EDFFXL R3_reg_2_ ( .D(data_in_2[104]), .E(n1261), .CK(clk), .QN(n887) );
  EDFFX1 R3_reg_1_ ( .D(data_in_2[103]), .E(n1261), .CK(clk), .QN(n888) );
  EDFFX1 R3_reg_0_ ( .D(data_in_2[102]), .E(n1260), .CK(clk), .QN(n889) );
  EDFFXL R7_reg_29_ ( .D(data_in_2[131]), .E(n1288), .CK(clk), .QN(n928) );
  EDFFXL R7_reg_27_ ( .D(data_in_2[129]), .E(n1288), .CK(clk), .QN(n930) );
  EDFFXL R7_reg_26_ ( .D(data_in_2[128]), .E(n1288), .CK(clk), .QN(n931) );
  EDFFXL R7_reg_25_ ( .D(data_in_2[127]), .E(n1288), .CK(clk), .QN(n932) );
  EDFFXL R7_reg_24_ ( .D(data_in_2[126]), .E(n1288), .CK(clk), .QN(n933) );
  EDFFXL R7_reg_23_ ( .D(data_in_2[125]), .E(n1288), .CK(clk), .QN(n934) );
  EDFFXL R7_reg_22_ ( .D(data_in_2[124]), .E(n1288), .CK(clk), .QN(n935) );
  EDFFXL R7_reg_21_ ( .D(data_in_2[123]), .E(n1288), .CK(clk), .QN(n936) );
  EDFFXL R7_reg_20_ ( .D(data_in_2[122]), .E(n1288), .CK(clk), .QN(n937) );
  EDFFXL R7_reg_19_ ( .D(data_in_2[121]), .E(n1288), .CK(clk), .QN(n938) );
  EDFFXL R7_reg_18_ ( .D(data_in_2[120]), .E(n1288), .CK(clk), .QN(n939) );
  EDFFX1 R7_reg_17_ ( .D(data_in_2[119]), .E(n1288), .CK(clk), .QN(n940) );
  EDFFXL R7_reg_10_ ( .D(data_in_2[112]), .E(n1288), .CK(clk), .QN(n947) );
  EDFFXL R7_reg_8_ ( .D(data_in_2[110]), .E(n1285), .CK(clk), .QN(n949) );
  EDFFXL R7_reg_7_ ( .D(data_in_2[109]), .E(n1286), .CK(clk), .QN(n950) );
  EDFFXL R7_reg_6_ ( .D(data_in_2[108]), .E(n1288), .CK(clk), .QN(n951) );
  EDFFXL R7_reg_5_ ( .D(data_in_2[107]), .E(n1286), .CK(clk), .QN(n952) );
  EDFFXL R7_reg_4_ ( .D(data_in_2[106]), .E(n1288), .CK(clk), .QN(n953) );
  EDFFXL R7_reg_3_ ( .D(data_in_2[105]), .E(n1285), .CK(clk), .QN(n954) );
  EDFFXL R7_reg_2_ ( .D(data_in_2[104]), .E(n1287), .CK(clk), .QN(n955) );
  EDFFX1 R7_reg_1_ ( .D(data_in_2[103]), .E(n1285), .CK(clk), .QN(n956) );
  EDFFX1 R7_reg_0_ ( .D(data_in_2[102]), .E(n1285), .CK(clk), .QN(n957) );
  EDFFX1 R8_reg_26_ ( .D(data_in_2[26]), .E(n1250), .CK(clk), .Q(R8[26]) );
  EDFFX1 R8_reg_25_ ( .D(data_in_2[25]), .E(n1250), .CK(clk), .Q(R8[25]) );
  EDFFX1 R8_reg_23_ ( .D(data_in_2[23]), .E(n1250), .CK(clk), .Q(R8[23]) );
  EDFFX1 R8_reg_22_ ( .D(data_in_2[22]), .E(n1250), .CK(clk), .Q(R8[22]) );
  EDFFXL R8_reg_20_ ( .D(data_in_2[20]), .E(n1250), .CK(clk), .Q(R8[20]) );
  EDFFXL R8_reg_19_ ( .D(n14), .E(n1250), .CK(clk), .Q(R8[19]) );
  EDFFX1 R8_reg_17_ ( .D(data_in_2[17]), .E(n1249), .CK(clk), .Q(R8[17]) );
  EDFFX1 R8_reg_9_ ( .D(data_in_2[9]), .E(n1249), .CK(clk), .Q(R8[9]) );
  EDFFX1 R8_reg_6_ ( .D(data_in_2[6]), .E(n1249), .CK(clk), .Q(R8[6]) );
  EDFFX1 R8_reg_5_ ( .D(data_in_2[5]), .E(n1248), .CK(clk), .Q(R8[5]) );
  EDFFX1 R8_reg_3_ ( .D(data_in_2[3]), .E(n1248), .CK(clk), .Q(R8[3]) );
  EDFFXL R8_reg_2_ ( .D(data_in_2[2]), .E(n1248), .CK(clk), .Q(R8[2]) );
  EDFFX1 R8_reg_1_ ( .D(data_in_2[1]), .E(n1248), .CK(clk), .Q(R8[1]) );
  EDFFX1 R8_reg_0_ ( .D(data_in_2[0]), .E(n1248), .CK(clk), .Q(R8[0]) );
  EDFFX1 R12_reg_26_ ( .D(data_in_2[26]), .E(n1271), .CK(clk), .Q(R12[26]) );
  EDFFX1 R12_reg_23_ ( .D(data_in_2[23]), .E(n1272), .CK(clk), .Q(R12[23]) );
  EDFFX1 R12_reg_22_ ( .D(data_in_2[22]), .E(n1275), .CK(clk), .Q(R12[22]) );
  EDFFXL R12_reg_20_ ( .D(data_in_2[20]), .E(n1275), .CK(clk), .Q(R12[20]) );
  EDFFXL R12_reg_19_ ( .D(n14), .E(n1276), .CK(clk), .Q(R12[19]) );
  EDFFX1 R12_reg_17_ ( .D(data_in_2[17]), .E(n1272), .CK(clk), .Q(R12[17]) );
  EDFFX1 R12_reg_9_ ( .D(data_in_2[9]), .E(n1276), .CK(clk), .Q(R12[9]) );
  EDFFX1 R12_reg_5_ ( .D(data_in_2[5]), .E(n1276), .CK(clk), .Q(R12[5]) );
  EDFFX1 R12_reg_3_ ( .D(data_in_2[3]), .E(n1275), .CK(clk), .Q(R12[3]) );
  EDFFXL R12_reg_2_ ( .D(data_in_2[2]), .E(n1275), .CK(clk), .Q(R12[2]) );
  EDFFX1 R12_reg_1_ ( .D(data_in_2[1]), .E(n1275), .CK(clk), .Q(R12[1]) );
  EDFFX1 R12_reg_0_ ( .D(data_in_2[0]), .E(n1275), .CK(clk), .Q(R12[0]) );
  EDFFX1 R0_reg_26_ ( .D(data_in_2[26]), .E(n1256), .CK(clk), .Q(R0[26]) );
  EDFFX1 R0_reg_25_ ( .D(data_in_2[25]), .E(n1256), .CK(clk), .Q(R0[25]) );
  EDFFX1 R0_reg_23_ ( .D(data_in_2[23]), .E(n1256), .CK(clk), .Q(R0[23]) );
  EDFFX1 R0_reg_22_ ( .D(data_in_2[22]), .E(n1256), .CK(clk), .Q(R0[22]) );
  EDFFXL R0_reg_20_ ( .D(data_in_2[20]), .E(n1256), .CK(clk), .Q(R0[20]) );
  EDFFXL R0_reg_19_ ( .D(n14), .E(n1256), .CK(clk), .Q(R0[19]) );
  EDFFX1 R0_reg_17_ ( .D(data_in_2[17]), .E(n1256), .CK(clk), .Q(R0[17]) );
  EDFFX1 R0_reg_9_ ( .D(data_in_2[9]), .E(n1257), .CK(clk), .Q(R0[9]) );
  EDFFX1 R0_reg_6_ ( .D(data_in_2[6]), .E(n1257), .CK(clk), .Q(R0[6]) );
  EDFFX1 R0_reg_5_ ( .D(data_in_2[5]), .E(n1257), .CK(clk), .Q(R0[5]) );
  EDFFX1 R0_reg_3_ ( .D(data_in_2[3]), .E(n1257), .CK(clk), .Q(R0[3]) );
  EDFFXL R0_reg_2_ ( .D(data_in_2[2]), .E(n1257), .CK(clk), .Q(R0[2]) );
  EDFFX1 R0_reg_1_ ( .D(data_in_2[1]), .E(n1257), .CK(clk), .Q(R0[1]) );
  EDFFX1 R0_reg_0_ ( .D(data_in_2[0]), .E(n1257), .CK(clk), .Q(R0[0]) );
  EDFFXL R4_reg_26_ ( .D(data_in_2[26]), .E(n1283), .CK(clk), .Q(R4[26]) );
  EDFFXL R4_reg_25_ ( .D(data_in_2[25]), .E(n1283), .CK(clk), .Q(R4[25]) );
  EDFFXL R4_reg_24_ ( .D(data_in_2[24]), .E(n1283), .CK(clk), .Q(R4[24]) );
  EDFFXL R4_reg_23_ ( .D(data_in_2[23]), .E(n1283), .CK(clk), .Q(R4[23]) );
  EDFFXL R4_reg_22_ ( .D(data_in_2[22]), .E(n1283), .CK(clk), .Q(R4[22]) );
  EDFFXL R4_reg_21_ ( .D(data_in_2[21]), .E(n1283), .CK(clk), .Q(R4[21]) );
  EDFFXL R4_reg_20_ ( .D(data_in_2[20]), .E(n1283), .CK(clk), .Q(R4[20]) );
  EDFFXL R4_reg_19_ ( .D(n14), .E(n1283), .CK(clk), .Q(R4[19]) );
  EDFFX1 R4_reg_17_ ( .D(data_in_2[17]), .E(n1283), .CK(clk), .Q(R4[17]) );
  EDFFXL R4_reg_12_ ( .D(data_in_2[12]), .E(n1284), .CK(clk), .Q(R4[12]) );
  EDFFXL R4_reg_8_ ( .D(data_in_2[8]), .E(n1284), .CK(clk), .Q(R4[8]) );
  EDFFXL R4_reg_7_ ( .D(data_in_2[7]), .E(n1284), .CK(clk), .Q(R4[7]) );
  EDFFXL R4_reg_6_ ( .D(data_in_2[6]), .E(n1284), .CK(clk), .Q(R4[6]) );
  EDFFXL R4_reg_5_ ( .D(data_in_2[5]), .E(n1284), .CK(clk), .Q(R4[5]) );
  EDFFXL R4_reg_4_ ( .D(data_in_2[4]), .E(n1284), .CK(clk), .Q(R4[4]) );
  EDFFXL R4_reg_3_ ( .D(data_in_2[3]), .E(n1284), .CK(clk), .Q(R4[3]) );
  EDFFXL R4_reg_2_ ( .D(data_in_2[2]), .E(n1284), .CK(clk), .Q(R4[2]) );
  EDFFX1 R4_reg_1_ ( .D(data_in_2[1]), .E(n1284), .CK(clk), .Q(R4[1]) );
  EDFFX1 R4_reg_0_ ( .D(data_in_2[0]), .E(n1284), .CK(clk), .Q(R4[0]) );
  EDFFXL R13_reg_30_ ( .D(data_in_2[64]), .E(n105), .CK(clk), .Q(R13[30]) );
  EDFFXL R13_reg_27_ ( .D(data_in_2[61]), .E(n1278), .CK(clk), .Q(R13[27]) );
  EDFFXL R13_reg_26_ ( .D(data_in_2[60]), .E(n1278), .CK(clk), .Q(R13[26]) );
  EDFFXL R13_reg_25_ ( .D(data_in_2[59]), .E(n1278), .CK(clk), .Q(R13[25]) );
  EDFFXL R13_reg_24_ ( .D(data_in_2[58]), .E(n1278), .CK(clk), .Q(R13[24]) );
  EDFFXL R13_reg_23_ ( .D(data_in_2[57]), .E(n1278), .CK(clk), .Q(R13[23]) );
  EDFFXL R13_reg_22_ ( .D(data_in_2[56]), .E(n1278), .CK(clk), .Q(R13[22]) );
  EDFFXL R13_reg_21_ ( .D(data_in_2[55]), .E(n1278), .CK(clk), .Q(R13[21]) );
  EDFFXL R13_reg_20_ ( .D(data_in_2[54]), .E(n1278), .CK(clk), .Q(R13[20]) );
  EDFFXL R13_reg_19_ ( .D(data_in_2[53]), .E(n1278), .CK(clk), .Q(R13[19]) );
  EDFFX1 R13_reg_18_ ( .D(data_in_2[52]), .E(n1278), .CK(clk), .Q(R13[18]) );
  EDFFX1 R13_reg_17_ ( .D(data_in_2[51]), .E(n1277), .CK(clk), .Q(R13[17]) );
  EDFFXL R13_reg_12_ ( .D(data_in_2[46]), .E(n1277), .CK(clk), .Q(R13[12]) );
  EDFFXL R13_reg_10_ ( .D(data_in_2[44]), .E(n1277), .CK(clk), .Q(R13[10]) );
  EDFFXL R13_reg_8_ ( .D(data_in_2[42]), .E(n1277), .CK(clk), .Q(R13[8]) );
  EDFFXL R13_reg_7_ ( .D(data_in_2[41]), .E(n1277), .CK(clk), .Q(R13[7]) );
  EDFFXL R13_reg_6_ ( .D(data_in_2[40]), .E(n1277), .CK(clk), .Q(R13[6]) );
  EDFFXL R13_reg_5_ ( .D(data_in_2[39]), .E(n1275), .CK(clk), .Q(R13[5]) );
  EDFFXL R13_reg_4_ ( .D(data_in_2[38]), .E(n105), .CK(clk), .Q(R13[4]) );
  EDFFXL R13_reg_3_ ( .D(data_in_2[37]), .E(n1276), .CK(clk), .Q(R13[3]) );
  EDFFXL R13_reg_2_ ( .D(data_in_2[36]), .E(n1276), .CK(clk), .Q(R13[2]) );
  EDFFX1 R13_reg_1_ ( .D(data_in_2[35]), .E(n105), .CK(clk), .Q(R13[1]) );
  EDFFX1 R13_reg_0_ ( .D(data_in_2[34]), .E(n105), .CK(clk), .Q(R13[0]) );
  EDFFXL R9_reg_30_ ( .D(data_in_2[64]), .E(n1243), .CK(clk), .Q(R9[30]) );
  EDFFXL R9_reg_27_ ( .D(data_in_2[61]), .E(n1243), .CK(clk), .Q(R9[27]) );
  EDFFXL R9_reg_26_ ( .D(data_in_2[60]), .E(n1243), .CK(clk), .Q(R9[26]) );
  EDFFXL R9_reg_25_ ( .D(data_in_2[59]), .E(n1243), .CK(clk), .Q(R9[25]) );
  EDFFXL R9_reg_24_ ( .D(data_in_2[58]), .E(n1243), .CK(clk), .Q(R9[24]) );
  EDFFXL R9_reg_23_ ( .D(data_in_2[57]), .E(n1247), .CK(clk), .Q(R9[23]) );
  EDFFXL R9_reg_22_ ( .D(data_in_2[56]), .E(n1246), .CK(clk), .Q(R9[22]) );
  EDFFXL R9_reg_21_ ( .D(data_in_2[55]), .E(n1245), .CK(clk), .Q(R9[21]) );
  EDFFXL R9_reg_20_ ( .D(data_in_2[54]), .E(n1243), .CK(clk), .Q(R9[20]) );
  EDFFXL R9_reg_19_ ( .D(data_in_2[53]), .E(n1249), .CK(clk), .Q(R9[19]) );
  EDFFX1 R9_reg_18_ ( .D(data_in_2[52]), .E(n1243), .CK(clk), .Q(R9[18]) );
  EDFFX1 R9_reg_17_ ( .D(data_in_2[51]), .E(n1251), .CK(clk), .Q(R9[17]) );
  EDFFXL R9_reg_12_ ( .D(data_in_2[46]), .E(n1251), .CK(clk), .Q(R9[12]) );
  EDFFXL R9_reg_10_ ( .D(data_in_2[44]), .E(n1249), .CK(clk), .Q(R9[10]) );
  EDFFXL R9_reg_8_ ( .D(data_in_2[42]), .E(n1244), .CK(clk), .Q(R9[8]) );
  EDFFXL R9_reg_7_ ( .D(data_in_2[41]), .E(n1251), .CK(clk), .Q(R9[7]) );
  EDFFXL R9_reg_6_ ( .D(data_in_2[40]), .E(n1249), .CK(clk), .Q(R9[6]) );
  EDFFXL R9_reg_5_ ( .D(data_in_2[39]), .E(n1251), .CK(clk), .Q(R9[5]) );
  EDFFXL R9_reg_4_ ( .D(data_in_2[38]), .E(n1249), .CK(clk), .Q(R9[4]) );
  EDFFXL R9_reg_3_ ( .D(data_in_2[37]), .E(n1243), .CK(clk), .Q(R9[3]) );
  EDFFXL R9_reg_2_ ( .D(data_in_2[36]), .E(n1243), .CK(clk), .Q(R9[2]) );
  EDFFX1 R9_reg_1_ ( .D(data_in_2[35]), .E(n1251), .CK(clk), .Q(R9[1]) );
  EDFFX1 R9_reg_0_ ( .D(data_in_2[34]), .E(n1251), .CK(clk), .Q(R9[0]) );
  EDFFXL R1_reg_30_ ( .D(data_in_2[64]), .E(n1257), .CK(clk), .Q(R1[30]) );
  EDFFXL R1_reg_27_ ( .D(data_in_2[61]), .E(n1257), .CK(clk), .Q(R1[27]) );
  EDFFXL R1_reg_26_ ( .D(data_in_2[60]), .E(n1257), .CK(clk), .Q(R1[26]) );
  EDFFXL R1_reg_25_ ( .D(data_in_2[59]), .E(n1258), .CK(clk), .Q(R1[25]) );
  EDFFXL R1_reg_24_ ( .D(data_in_2[58]), .E(n1258), .CK(clk), .Q(R1[24]) );
  EDFFXL R1_reg_23_ ( .D(data_in_2[57]), .E(n1258), .CK(clk), .Q(R1[23]) );
  EDFFXL R1_reg_22_ ( .D(data_in_2[56]), .E(n1258), .CK(clk), .Q(R1[22]) );
  EDFFXL R1_reg_21_ ( .D(data_in_2[55]), .E(n1258), .CK(clk), .Q(R1[21]) );
  EDFFXL R1_reg_20_ ( .D(data_in_2[54]), .E(n1258), .CK(clk), .Q(R1[20]) );
  EDFFXL R1_reg_19_ ( .D(data_in_2[53]), .E(n1258), .CK(clk), .Q(R1[19]) );
  EDFFX1 R1_reg_18_ ( .D(data_in_2[52]), .E(n1258), .CK(clk), .Q(R1[18]) );
  EDFFX1 R1_reg_17_ ( .D(data_in_2[51]), .E(n1258), .CK(clk), .Q(R1[17]) );
  EDFFXL R1_reg_12_ ( .D(data_in_2[46]), .E(n1258), .CK(clk), .Q(R1[12]) );
  EDFFXL R1_reg_10_ ( .D(data_in_2[44]), .E(n1258), .CK(clk), .Q(R1[10]) );
  EDFFXL R1_reg_8_ ( .D(data_in_2[42]), .E(n1258), .CK(clk), .Q(R1[8]) );
  EDFFXL R1_reg_7_ ( .D(data_in_2[41]), .E(n1258), .CK(clk), .Q(R1[7]) );
  EDFFXL R1_reg_6_ ( .D(data_in_2[40]), .E(n1258), .CK(clk), .Q(R1[6]) );
  EDFFXL R1_reg_5_ ( .D(data_in_2[39]), .E(n1258), .CK(clk), .Q(R1[5]) );
  EDFFXL R1_reg_4_ ( .D(data_in_2[38]), .E(n1258), .CK(clk), .Q(R1[4]) );
  EDFFXL R1_reg_3_ ( .D(data_in_2[37]), .E(n1259), .CK(clk), .Q(R1[3]) );
  EDFFXL R1_reg_2_ ( .D(data_in_2[36]), .E(n1259), .CK(clk), .Q(R1[2]) );
  EDFFX1 R1_reg_1_ ( .D(data_in_2[35]), .E(n1259), .CK(clk), .Q(R1[1]) );
  EDFFX1 R1_reg_0_ ( .D(data_in_2[34]), .E(n1259), .CK(clk), .Q(R1[0]) );
  EDFFXL R5_reg_30_ ( .D(data_in_2[64]), .E(n1284), .CK(clk), .Q(R5[30]) );
  EDFFXL R5_reg_27_ ( .D(data_in_2[61]), .E(n1284), .CK(clk), .Q(R5[27]) );
  EDFFXL R5_reg_26_ ( .D(data_in_2[60]), .E(n1285), .CK(clk), .Q(R5[26]) );
  EDFFXL R5_reg_25_ ( .D(data_in_2[59]), .E(n1285), .CK(clk), .Q(R5[25]) );
  EDFFXL R5_reg_24_ ( .D(data_in_2[58]), .E(n1285), .CK(clk), .Q(R5[24]) );
  EDFFXL R5_reg_23_ ( .D(data_in_2[57]), .E(n1285), .CK(clk), .Q(R5[23]) );
  EDFFXL R5_reg_22_ ( .D(data_in_2[56]), .E(n1285), .CK(clk), .Q(R5[22]) );
  EDFFXL R5_reg_21_ ( .D(data_in_2[55]), .E(n1285), .CK(clk), .Q(R5[21]) );
  EDFFXL R5_reg_20_ ( .D(data_in_2[54]), .E(n1285), .CK(clk), .Q(R5[20]) );
  EDFFXL R5_reg_19_ ( .D(data_in_2[53]), .E(n1285), .CK(clk), .Q(R5[19]) );
  EDFFX1 R5_reg_18_ ( .D(data_in_2[52]), .E(n1285), .CK(clk), .Q(R5[18]) );
  EDFFX1 R5_reg_17_ ( .D(data_in_2[51]), .E(n1285), .CK(clk), .Q(R5[17]) );
  EDFFXL R5_reg_12_ ( .D(data_in_2[46]), .E(n1285), .CK(clk), .Q(R5[12]) );
  EDFFXL R5_reg_10_ ( .D(data_in_2[44]), .E(n1285), .CK(clk), .Q(R5[10]) );
  EDFFXL R5_reg_8_ ( .D(data_in_2[42]), .E(n1285), .CK(clk), .Q(R5[8]) );
  EDFFXL R5_reg_7_ ( .D(data_in_2[41]), .E(n1285), .CK(clk), .Q(R5[7]) );
  EDFFXL R5_reg_6_ ( .D(data_in_2[40]), .E(n1285), .CK(clk), .Q(R5[6]) );
  EDFFXL R5_reg_5_ ( .D(data_in_2[39]), .E(n1286), .CK(clk), .Q(R5[5]) );
  EDFFXL R5_reg_4_ ( .D(data_in_2[38]), .E(n1286), .CK(clk), .Q(R5[4]) );
  EDFFXL R5_reg_3_ ( .D(data_in_2[37]), .E(n1286), .CK(clk), .Q(R5[3]) );
  EDFFXL R5_reg_2_ ( .D(data_in_2[36]), .E(n1286), .CK(clk), .Q(R5[2]) );
  EDFFX1 R5_reg_1_ ( .D(data_in_2[35]), .E(n1286), .CK(clk), .Q(R5[1]) );
  EDFFX1 R5_reg_0_ ( .D(data_in_2[34]), .E(n1286), .CK(clk), .Q(R5[0]) );
  DFFHQX1 reg_flag_mux_reg ( .D(n1319), .CK(clk), .Q(reg_flag_mux) );
  DFFHQX1 counter1_reg_1_ ( .D(n1115), .CK(clk), .Q(counter1[1]) );
  EDFFX1 data_out_2_reg_16_ ( .D(N68), .E(n1315), .CK(clk), .Q(data_out_2[16])
         );
  DFFHQX1 counter2_reg_0_ ( .D(n1114), .CK(clk), .Q(counter2[0]) );
  DFFHQX1 counter2_reg_1_ ( .D(n1113), .CK(clk), .Q(counter2[1]) );
  EDFFX1 data_out_2_reg_32_ ( .D(N84), .E(n1317), .CK(clk), .Q(data_out_2[32])
         );
  EDFFX1 data_out_2_reg_15_ ( .D(N67), .E(n1315), .CK(clk), .Q(data_out_2[15])
         );
  EDFFX1 data_out_2_reg_31_ ( .D(N83), .E(n1317), .CK(clk), .Q(data_out_2[31])
         );
  EDFFX1 data_out_2_reg_30_ ( .D(N82), .E(n1317), .CK(clk), .Q(data_out_2[30])
         );
  EDFFX1 data_out_2_reg_29_ ( .D(N81), .E(n1317), .CK(clk), .Q(data_out_2[29])
         );
  EDFFX1 data_out_2_reg_28_ ( .D(N80), .E(n1317), .CK(clk), .Q(data_out_2[28])
         );
  EDFFX1 data_out_2_reg_27_ ( .D(N79), .E(n1317), .CK(clk), .Q(data_out_2[27])
         );
  EDFFX1 data_out_2_reg_26_ ( .D(N78), .E(n1317), .CK(clk), .Q(data_out_2[26])
         );
  EDFFX1 data_out_2_reg_25_ ( .D(N77), .E(n1317), .CK(clk), .Q(data_out_2[25])
         );
  EDFFX1 data_out_2_reg_14_ ( .D(N66), .E(n1317), .CK(clk), .Q(data_out_2[14])
         );
  EDFFX1 data_out_2_reg_13_ ( .D(N65), .E(n1316), .CK(clk), .Q(data_out_2[13])
         );
  EDFFX1 data_out_2_reg_12_ ( .D(N64), .E(n1315), .CK(clk), .Q(data_out_2[12])
         );
  EDFFX1 data_out_2_reg_11_ ( .D(N63), .E(n1315), .CK(clk), .Q(data_out_2[11])
         );
  EDFFX1 data_out_2_reg_10_ ( .D(N62), .E(n1317), .CK(clk), .Q(data_out_2[10])
         );
  EDFFX1 data_out_2_reg_5_ ( .D(N57), .E(n1316), .CK(clk), .Q(data_out_2[5])
         );
  EDFFX1 data_out_2_reg_24_ ( .D(N76), .E(n1317), .CK(clk), .Q(data_out_2[24])
         );
  EDFFX1 data_out_2_reg_23_ ( .D(N75), .E(n1317), .CK(clk), .Q(data_out_2[23])
         );
  EDFFX1 data_out_2_reg_22_ ( .D(N74), .E(n1317), .CK(clk), .Q(data_out_2[22])
         );
  EDFFX1 data_out_2_reg_21_ ( .D(N73), .E(n1317), .CK(clk), .Q(data_out_2[21])
         );
  EDFFX1 data_out_2_reg_20_ ( .D(N72), .E(n1317), .CK(clk), .Q(data_out_2[20])
         );
  EDFFX1 data_out_2_reg_19_ ( .D(N71), .E(n1316), .CK(clk), .Q(data_out_2[19])
         );
  EDFFX1 data_out_2_reg_18_ ( .D(N70), .E(n1317), .CK(clk), .Q(data_out_2[18])
         );
  EDFFX1 data_out_2_reg_17_ ( .D(N69), .E(n1316), .CK(clk), .Q(data_out_2[17])
         );
  EDFFX1 data_out_2_reg_9_ ( .D(N61), .E(n1317), .CK(clk), .Q(data_out_2[9])
         );
  EDFFX1 data_out_2_reg_8_ ( .D(N60), .E(n1316), .CK(clk), .Q(data_out_2[8])
         );
  EDFFX1 data_out_2_reg_7_ ( .D(N59), .E(n1316), .CK(clk), .Q(data_out_2[7])
         );
  EDFFX1 data_out_2_reg_6_ ( .D(N58), .E(n1315), .CK(clk), .Q(data_out_2[6])
         );
  EDFFX1 data_out_2_reg_4_ ( .D(N56), .E(n1317), .CK(clk), .Q(data_out_2[4])
         );
  EDFFX1 data_out_2_reg_3_ ( .D(N55), .E(n1316), .CK(clk), .Q(data_out_2[3])
         );
  EDFFX1 data_out_2_reg_2_ ( .D(N54), .E(n1317), .CK(clk), .Q(data_out_2[2])
         );
  EDFFX1 data_out_2_reg_1_ ( .D(N53), .E(n1315), .CK(clk), .Q(data_out_2[1])
         );
  EDFFX1 data_out_2_reg_0_ ( .D(N52), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[0]) );
  EDFFX1 data_out_2_reg_135_ ( .D(N187), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[135]) );
  EDFFXL R8_reg_18_ ( .D(data_in_2[18]), .E(n1250), .CK(clk), .Q(R8[18]) );
  EDFFXL R12_reg_18_ ( .D(data_in_2[18]), .E(n1272), .CK(clk), .Q(R12[18]) );
  EDFFXL R0_reg_18_ ( .D(data_in_2[18]), .E(n1256), .CK(clk), .Q(R0[18]) );
  EDFFXL R4_reg_18_ ( .D(data_in_2[18]), .E(n1283), .CK(clk), .Q(R4[18]) );
  EDFFX1 R10_reg_17_ ( .D(data_in_2[85]), .E(n1245), .CK(clk), .QN(n736) );
  EDFFX1 R11_reg_17_ ( .D(data_in_2[119]), .E(n109), .CK(clk), .QN(n702) );
  EDFFX1 R11_reg_1_ ( .D(data_in_2[103]), .E(n1246), .CK(clk), .QN(n718) );
  EDFFX1 R11_reg_0_ ( .D(data_in_2[102]), .E(n1246), .CK(clk), .QN(n719) );
  EDFFXL R10_reg_27_ ( .D(data_in_2[95]), .E(n1246), .CK(clk), .QN(n726) );
  EDFFXL R2_reg_27_ ( .D(data_in_2[95]), .E(n1259), .CK(clk), .QN(n828) );
  EDFFXL R14_reg_27_ ( .D(data_in_2[95]), .E(n1275), .CK(clk), .QN(n760) );
  EDFFXL R8_reg_8_ ( .D(data_in_2[8]), .E(n1249), .CK(clk), .Q(R8[8]) );
  EDFFXL R12_reg_8_ ( .D(data_in_2[8]), .E(n1276), .CK(clk), .Q(R12[8]) );
  EDFFXL R0_reg_8_ ( .D(data_in_2[8]), .E(n1257), .CK(clk), .Q(R0[8]) );
  EDFFXL R8_reg_4_ ( .D(data_in_2[4]), .E(n1248), .CK(clk), .Q(R8[4]) );
  EDFFXL R12_reg_4_ ( .D(data_in_2[4]), .E(n1276), .CK(clk), .Q(R12[4]) );
  EDFFXL R0_reg_4_ ( .D(data_in_2[4]), .E(n1257), .CK(clk), .Q(R0[4]) );
  EDFFXL R3_reg_5_ ( .D(data_in_2[107]), .E(n1260), .CK(clk), .QN(n884) );
  EDFFXL R15_reg_5_ ( .D(data_in_2[107]), .E(n1271), .CK(clk), .QN(n816) );
  EDFFXL R11_reg_5_ ( .D(data_in_2[107]), .E(n1247), .CK(clk), .QN(n714) );
  EDFFXL R11_reg_7_ ( .D(data_in_2[109]), .E(n1247), .CK(clk), .QN(n712) );
  EDFFXL R15_reg_7_ ( .D(data_in_2[109]), .E(n1271), .CK(clk), .QN(n814) );
  EDFFXL R3_reg_7_ ( .D(data_in_2[109]), .E(n1261), .CK(clk), .QN(n882) );
  EDFFXL R15_reg_23_ ( .D(data_in_2[125]), .E(n1272), .CK(clk), .QN(n798) );
  EDFFXL R3_reg_23_ ( .D(data_in_2[125]), .E(n1261), .CK(clk), .QN(n866) );
  EDFFXL R11_reg_23_ ( .D(data_in_2[125]), .E(n109), .CK(clk), .QN(n696) );
  EDFFXL R11_reg_6_ ( .D(data_in_2[108]), .E(n1247), .CK(clk), .QN(n713) );
  EDFFXL R15_reg_6_ ( .D(data_in_2[108]), .E(n1271), .CK(clk), .QN(n815) );
  EDFFXL R3_reg_6_ ( .D(data_in_2[108]), .E(n1261), .CK(clk), .QN(n883) );
  EDFFXL R8_reg_24_ ( .D(data_in_2[24]), .E(n1250), .CK(clk), .Q(R8[24]) );
  EDFFXL R12_reg_24_ ( .D(data_in_2[24]), .E(n105), .CK(clk), .Q(R12[24]) );
  EDFFXL R0_reg_24_ ( .D(data_in_2[24]), .E(n1256), .CK(clk), .Q(R0[24]) );
  EDFFXL R10_reg_23_ ( .D(data_in_2[91]), .E(n1245), .CK(clk), .QN(n730) );
  EDFFXL R14_reg_23_ ( .D(data_in_2[91]), .E(n1275), .CK(clk), .QN(n764) );
  EDFFXL R2_reg_23_ ( .D(data_in_2[91]), .E(n1259), .CK(clk), .QN(n832) );
  EDFFXL R10_reg_7_ ( .D(data_in_2[75]), .E(n1244), .CK(clk), .QN(n746) );
  EDFFXL R14_reg_7_ ( .D(data_in_2[75]), .E(n1274), .CK(clk), .QN(n780) );
  EDFFXL R2_reg_7_ ( .D(data_in_2[75]), .E(n1260), .CK(clk), .QN(n848) );
  EDFFXL R8_reg_7_ ( .D(data_in_2[7]), .E(n1249), .CK(clk), .Q(R8[7]) );
  EDFFXL R12_reg_7_ ( .D(data_in_2[7]), .E(n1276), .CK(clk), .Q(R12[7]) );
  EDFFXL R0_reg_7_ ( .D(data_in_2[7]), .E(n1257), .CK(clk), .Q(R0[7]) );
  EDFFXL R10_reg_25_ ( .D(data_in_2[93]), .E(n1245), .CK(clk), .QN(n728) );
  EDFFXL R14_reg_25_ ( .D(data_in_2[93]), .E(n105), .CK(clk), .QN(n762) );
  EDFFXL R2_reg_25_ ( .D(data_in_2[93]), .E(n1259), .CK(clk), .QN(n830) );
  EDFFXL R10_reg_4_ ( .D(data_in_2[72]), .E(n1244), .CK(clk), .QN(n749) );
  EDFFXL R14_reg_4_ ( .D(data_in_2[72]), .E(n1274), .CK(clk), .QN(n783) );
  EDFFXL R2_reg_4_ ( .D(data_in_2[72]), .E(n1260), .CK(clk), .QN(n851) );
  EDFFXL R2_reg_21_ ( .D(data_in_2[89]), .E(n1259), .CK(clk), .QN(n834) );
  EDFFXL R14_reg_21_ ( .D(data_in_2[89]), .E(n1277), .CK(clk), .QN(n766) );
  EDFFXL R10_reg_21_ ( .D(data_in_2[89]), .E(n1245), .CK(clk), .QN(n732) );
  EDFFXL R2_reg_5_ ( .D(data_in_2[73]), .E(n1260), .CK(clk), .QN(n850) );
  EDFFXL R14_reg_5_ ( .D(data_in_2[73]), .E(n1274), .CK(clk), .QN(n782) );
  EDFFXL R10_reg_5_ ( .D(data_in_2[73]), .E(n1244), .CK(clk), .QN(n748) );
  EDFFXL R8_reg_21_ ( .D(data_in_2[21]), .E(n1250), .CK(clk), .Q(R8[21]) );
  EDFFXL R12_reg_21_ ( .D(data_in_2[21]), .E(n1274), .CK(clk), .Q(R12[21]) );
  EDFFXL R0_reg_21_ ( .D(data_in_2[21]), .E(n1256), .CK(clk), .Q(R0[21]) );
  EDFFXL R10_reg_12_ ( .D(data_in_2[80]), .E(n1244), .CK(clk), .QN(n741) );
  EDFFXL R14_reg_12_ ( .D(data_in_2[80]), .E(n1274), .CK(clk), .QN(n775) );
  EDFFXL R2_reg_12_ ( .D(data_in_2[80]), .E(n1260), .CK(clk), .QN(n843) );
  EDFFXL R15_reg_4_ ( .D(data_in_2[106]), .E(n1271), .CK(clk), .QN(n817) );
  EDFFXL R3_reg_4_ ( .D(data_in_2[106]), .E(n1260), .CK(clk), .QN(n885) );
  EDFFXL R11_reg_4_ ( .D(data_in_2[106]), .E(n1247), .CK(clk), .QN(n715) );
  EDFFXL R11_reg_10_ ( .D(data_in_2[112]), .E(n1247), .CK(clk), .QN(n709) );
  EDFFXL R15_reg_10_ ( .D(data_in_2[112]), .E(n1271), .CK(clk), .QN(n811) );
  EDFFXL R3_reg_10_ ( .D(data_in_2[112]), .E(n1261), .CK(clk), .QN(n879) );
  EDFFXL R11_reg_26_ ( .D(data_in_2[128]), .E(n109), .CK(clk), .QN(n693) );
  EDFFXL R15_reg_26_ ( .D(data_in_2[128]), .E(n1273), .CK(clk), .QN(n795) );
  EDFFXL R3_reg_26_ ( .D(data_in_2[128]), .E(n1261), .CK(clk), .QN(n863) );
  EDFFXL R11_reg_29_ ( .D(data_in_2[131]), .E(n1248), .CK(clk), .QN(n690) );
  EDFFXL R15_reg_29_ ( .D(data_in_2[131]), .E(n1273), .CK(clk), .QN(n792) );
  EDFFXL R3_reg_29_ ( .D(data_in_2[131]), .E(n1260), .CK(clk), .QN(n860) );
  EDFFXL R8_reg_12_ ( .D(data_in_2[12]), .E(n1249), .CK(clk), .Q(R8[12]) );
  EDFFXL R12_reg_12_ ( .D(data_in_2[12]), .E(n1276), .CK(clk), .Q(R12[12]) );
  EDFFXL R0_reg_12_ ( .D(data_in_2[12]), .E(n1257), .CK(clk), .Q(R0[12]) );
  DFFXL R4_reg_33_ ( .D(n1187), .CK(clk), .Q(n102) );
  DFFXL R8_reg_33_ ( .D(n1188), .CK(clk), .Q(n100) );
  DFFXL R1_reg_33_ ( .D(n1142), .CK(clk), .Q(n97) );
  DFFXL R9_reg_33_ ( .D(n1144), .CK(clk), .Q(n93) );
  DFFXL R13_reg_33_ ( .D(n1145), .CK(clk), .Q(n92) );
  DFFXL R5_reg_33_ ( .D(n1143), .CK(clk), .Q(n91) );
  DFFXL R4_reg_16_ ( .D(n1205), .CK(clk), .Q(n87) );
  EDFFX1 R4_reg_9_ ( .D(data_in_2[9]), .E(n1284), .CK(clk), .Q(R4[9]) );
  EDFFXL R10_reg_26_ ( .D(data_in_2[94]), .E(n1246), .CK(clk), .QN(n727) );
  EDFFXL R14_reg_26_ ( .D(data_in_2[94]), .E(n1275), .CK(clk), .QN(n761) );
  EDFFXL R2_reg_26_ ( .D(data_in_2[94]), .E(n1259), .CK(clk), .QN(n829) );
  DFFXL R8_reg_31_ ( .D(n1174), .CK(clk), .Q(n77) );
  DFFXL R12_reg_31_ ( .D(n1175), .CK(clk), .Q(n75) );
  DFFXL R13_reg_31_ ( .D(n1163), .CK(clk), .Q(n73) );
  DFFXL R9_reg_31_ ( .D(n1162), .CK(clk), .Q(n71), .QN(n70) );
  DFFXL R5_reg_31_ ( .D(n1161), .CK(clk), .Q(n69) );
  DFFXL R1_reg_31_ ( .D(n1160), .CK(clk), .Q(n68) );
  EDFFXL R3_reg_27_ ( .D(data_in_2[129]), .E(n1261), .CK(clk), .QN(n862) );
  EDFFXL R15_reg_27_ ( .D(data_in_2[129]), .E(n1273), .CK(clk), .QN(n794) );
  EDFFXL R11_reg_27_ ( .D(data_in_2[129]), .E(n109), .CK(clk), .QN(n692) );
  DFFXL R1_reg_11_ ( .D(n1164), .CK(clk), .Q(n63) );
  DFFXL R0_reg_33_ ( .D(n1186), .CK(clk), .Q(n61) );
  EDFFX1 R13_reg_9_ ( .D(data_in_2[43]), .E(n1277), .CK(clk), .Q(R13[9]) );
  EDFFXL R9_reg_32_ ( .D(data_in_2[66]), .E(n195), .CK(clk), .Q(R9[32]) );
  EDFFXL R12_reg_33_ ( .D(data_in_2[33]), .E(n971), .CK(clk), .Q(R12[33]) );
  EDFFXL R13_reg_15_ ( .D(data_in_2[49]), .E(n971), .CK(clk), .Q(R13[15]) );
  EDFFXL R8_reg_16_ ( .D(data_in_2[16]), .E(n195), .CK(clk), .Q(n90) );
  EDFFXL R15_reg_16_ ( .D(data_in_2[118]), .E(n971), .CK(clk), .QN(n805) );
  EDFFXL R14_reg_16_ ( .D(data_in_2[84]), .E(n1274), .CK(clk), .QN(n771) );
  EDFFXL R10_reg_16_ ( .D(data_in_2[84]), .E(n195), .CK(clk), .QN(n737) );
  EDFFXL R14_reg_13_ ( .D(data_in_2[81]), .E(n1274), .CK(clk), .QN(n774) );
  EDFFXL R9_reg_15_ ( .D(data_in_2[49]), .E(n195), .CK(clk), .Q(R9[15]) );
  EDFFXL R11_reg_16_ ( .D(data_in_2[118]), .E(n195), .CK(clk), .QN(n703) );
  DFFXL R13_reg_32_ ( .D(n1148), .CK(clk), .Q(R13[32]) );
  EDFFXL R5_reg_32_ ( .D(data_in_2[66]), .E(n969), .CK(clk), .Q(R5[32]) );
  EDFFXL R10_reg_13_ ( .D(data_in_2[81]), .E(n195), .CK(clk), .QN(n740) );
  EDFFXL R8_reg_10_ ( .D(data_in_2[10]), .E(n195), .CK(clk), .Q(n98) );
  EDFFXL R12_reg_16_ ( .D(data_in_2[16]), .E(n1278), .CK(clk), .Q(n89) );
  EDFFX1 R5_reg_9_ ( .D(data_in_2[43]), .E(n1285), .CK(clk), .Q(R5[9]) );
  EDFFX1 R1_reg_9_ ( .D(data_in_2[43]), .E(n1258), .CK(clk), .Q(R1[9]) );
  EDFFX1 R9_reg_9_ ( .D(data_in_2[43]), .E(n1251), .CK(clk), .Q(R9[9]) );
  DFFXL R1_reg_32_ ( .D(n1147), .CK(clk), .Q(n39) );
  EDFFXL R10_reg_33_ ( .D(data_in_2[101]), .E(n195), .CK(clk), .QN(n720) );
  EDFFXL R10_reg_8_ ( .D(data_in_2[76]), .E(n1244), .CK(clk), .QN(n745) );
  EDFFXL R14_reg_8_ ( .D(data_in_2[76]), .E(n1274), .CK(clk), .QN(n779) );
  EDFFXL R2_reg_8_ ( .D(data_in_2[76]), .E(n1260), .CK(clk), .QN(n847) );
  DFFXL R1_reg_15_ ( .D(n1146), .CK(clk), .Q(n31), .QN(n30) );
  EDFFXL R11_reg_11_ ( .D(data_in_2[113]), .E(n195), .CK(clk), .QN(n708) );
  EDFFXL R8_reg_27_ ( .D(data_in_2[27]), .E(n195), .CK(clk), .Q(R8[27]) );
  EDFFXL R0_reg_16_ ( .D(data_in_2[16]), .E(n1256), .CK(clk), .Q(R0[16]) );
  DFFXL counter1_reg_0_ ( .D(n1116), .CK(clk), .Q(counter1[0]), .QN(n1320) );
  EDFFXL R0_reg_10_ ( .D(data_in_2[10]), .E(n196), .CK(clk), .Q(n96) );
  EDFFXL R12_reg_25_ ( .D(data_in_2[25]), .E(n1271), .CK(clk), .Q(R12[25]) );
  EDFFXL R14_reg_22_ ( .D(data_in_2[90]), .E(n1271), .CK(clk), .QN(n765) );
  EDFFXL R14_reg_14_ ( .D(data_in_2[82]), .E(n1273), .CK(clk), .QN(n773) );
  EDFFXL R5_reg_15_ ( .D(data_in_2[49]), .E(n1285), .CK(clk), .Q(n33) );
  EDFFXL R12_reg_6_ ( .D(data_in_2[6]), .E(n1276), .CK(clk), .Q(R12[6]) );
  EDFFXL R3_reg_21_ ( .D(data_in_2[123]), .E(n1261), .CK(clk), .QN(n868) );
  EDFFXL R11_reg_21_ ( .D(data_in_2[123]), .E(n109), .CK(clk), .QN(n698) );
  EDFFXL R15_reg_21_ ( .D(data_in_2[123]), .E(n1272), .CK(clk), .QN(n800) );
  EDFFXL R3_reg_20_ ( .D(data_in_2[122]), .E(n1261), .CK(clk), .QN(n869) );
  EDFFXL R11_reg_20_ ( .D(data_in_2[122]), .E(n109), .CK(clk), .QN(n699) );
  EDFFXL R15_reg_20_ ( .D(data_in_2[122]), .E(n1272), .CK(clk), .QN(n801) );
  EDFFX2 data_out_2_reg_118_ ( .D(N170), .E(n1316), .CK(clk), .Q(
        data_out_2[118]) );
  EDFFX2 data_out_2_reg_84_ ( .D(N136), .E(n1315), .CK(clk), .Q(data_out_2[84]) );
  EDFFX1 data_out_2_reg_67_ ( .D(N119), .E(n1315), .CK(clk), .Q(data_out_2[67]) );
  EDFFX2 data_out_2_reg_101_ ( .D(N153), .E(n1317), .CK(clk), .Q(
        data_out_2[101]) );
  EDFFX2 data_out_2_reg_50_ ( .D(N102), .E(n1316), .CK(clk), .Q(data_out_2[50]) );
  MX2X2 U3 ( .A(data_in_2[135]), .B(n1227), .S0(n1255), .Y(n1140) );
  MX2X2 U4 ( .A(data_in_2[135]), .B(n1228), .S0(n1279), .Y(n1141) );
  MX2X2 U5 ( .A(data_in_2[11]), .B(R0[11]), .S0(n16), .Y(n1218) );
  MX2X2 U6 ( .A(data_in_2[16]), .B(n87), .S0(n17), .Y(n1205) );
  INVX1 U7 ( .A(n1257), .Y(n85) );
  INVX1 U8 ( .A(n105), .Y(n38) );
  INVX1 U9 ( .A(n1287), .Y(n18) );
  INVX1 U10 ( .A(n1259), .Y(n44) );
  NAND2X1 U11 ( .A(n471), .B(n104), .Y(n19) );
  MX2X2 U12 ( .A(data_in_2[79]), .B(n454), .S0(n43), .Y(n1129) );
  INVX1 U13 ( .A(n1274), .Y(n43) );
  INVX1 U14 ( .A(n1277), .Y(n84) );
  AOI22XL U15 ( .A0(R5[11]), .A1(n1305), .B0(n1270), .B1(R4[11]), .Y(n979) );
  AOI22XL U16 ( .A0(R9[11]), .A1(n1300), .B0(n1264), .B1(R8[11]), .Y(n1081) );
  AOI22XL U17 ( .A0(R13[11]), .A1(n1302), .B0(n1267), .B1(R12[11]), .Y(n1047)
         );
  MX2X1 U18 ( .A(n63), .B(data_in_2[45]), .S0(n1258), .Y(n1164) );
  AND2X2 U19 ( .A(counter2[1]), .B(n1322), .Y(n6) );
  OR2X2 U20 ( .A(counter2[0]), .B(counter2[1]), .Y(n7) );
  INVX1 U21 ( .A(n1252), .Y(n109) );
  INVX1 U22 ( .A(n1256), .Y(n95) );
  INVX1 U23 ( .A(n1283), .Y(n17) );
  INVX1 U24 ( .A(n1283), .Y(n86) );
  INVX1 U25 ( .A(n1281), .Y(n105) );
  INVX1 U26 ( .A(n1281), .Y(n1275) );
  INVX1 U27 ( .A(n105), .Y(n104) );
  INVX1 U28 ( .A(n1284), .Y(n83) );
  INVX1 U29 ( .A(n196), .Y(n16) );
  MX2X2 U30 ( .A(R4[11]), .B(data_in_2[11]), .S0(n1284), .Y(n1219) );
  MX2X1 U31 ( .A(data_in_2[11]), .B(R8[11]), .S0(n1253), .Y(n1220) );
  MX2X1 U32 ( .A(data_in_2[11]), .B(R12[11]), .S0(n104), .Y(n1221) );
  BUFX3 U33 ( .A(data_in_2[19]), .Y(n14) );
  MX2X2 U34 ( .A(data_in_2[67]), .B(n97), .S0(n15), .Y(n1142) );
  CLKINVX20 U35 ( .A(n1257), .Y(n15) );
  MX2X2 U36 ( .A(data_in_2[81]), .B(n320), .S0(n16), .Y(n682) );
  MX2X2 U37 ( .A(data_in_2[33]), .B(n102), .S0(n17), .Y(n1187) );
  MX2X2 U38 ( .A(data_in_2[81]), .B(n184), .S0(n18), .Y(n683) );
  NAND2X1 U39 ( .A(data_in_2[96]), .B(n1275), .Y(n20) );
  NAND2X2 U40 ( .A(n19), .B(n20), .Y(n1121) );
  MX2X2 U41 ( .A(data_in_2[66]), .B(n39), .S0(n85), .Y(n1147) );
  MX2X4 U42 ( .A(data_in_2[66]), .B(R13[32]), .S0(n1279), .Y(n1148) );
  MX2X2 U43 ( .A(n474), .B(data_in_2[99]), .S0(n1275), .Y(n662) );
  MX2X2 U44 ( .A(n542), .B(data_in_2[99]), .S0(n1246), .Y(n661) );
  MX2X2 U45 ( .A(n338), .B(data_in_2[99]), .S0(n1259), .Y(n659) );
  MX2X2 U46 ( .A(n202), .B(data_in_2[99]), .S0(n1286), .Y(n660) );
  MX2X2 U47 ( .A(n1229), .B(data_in_2[135]), .S0(n1260), .Y(n1138) );
  MX2X2 U48 ( .A(n1230), .B(data_in_2[135]), .S0(n1287), .Y(n1139) );
  INVX1 U49 ( .A(n30), .Y(n32) );
  MX2X2 U50 ( .A(data_in_2[15]), .B(R8[15]), .S0(n1253), .Y(n1195) );
  MX2X2 U51 ( .A(data_in_2[15]), .B(R12[15]), .S0(n104), .Y(n1196) );
  MX2X2 U52 ( .A(data_in_2[15]), .B(R0[15]), .S0(n16), .Y(n1193) );
  MX2X2 U53 ( .A(data_in_2[15]), .B(R4[15]), .S0(n83), .Y(n1194) );
  MX2X2 U54 ( .A(R12[13]), .B(data_in_2[13]), .S0(n1276), .Y(n1179) );
  MX2X2 U55 ( .A(R8[13]), .B(data_in_2[13]), .S0(n1249), .Y(n1178) );
  MX2X2 U56 ( .A(R0[13]), .B(data_in_2[13]), .S0(n1257), .Y(n1176) );
  MX2X2 U57 ( .A(R4[13]), .B(data_in_2[13]), .S0(n1284), .Y(n1177) );
  AOI22XL U58 ( .A0(n68), .A1(n1305), .B0(n1270), .B1(R0[31]), .Y(n993) );
  AOI22XL U59 ( .A0(n69), .A1(n1299), .B0(n1269), .B1(R4[31]), .Y(n1095) );
  AOI22XL U60 ( .A0(n33), .A1(n1298), .B0(n1263), .B1(R4[15]), .Y(n1111) );
  AOI22XL U61 ( .A0(n31), .A1(n1303), .B0(n1263), .B1(R0[15]), .Y(n1009) );
  MX2X4 U62 ( .A(data_in_2[49]), .B(n32), .S0(n16), .Y(n1146) );
  MX2X2 U63 ( .A(n1236), .B(data_in_2[133]), .S0(n1273), .Y(n1125) );
  MX2X2 U64 ( .A(n1235), .B(data_in_2[133]), .S0(n1248), .Y(n1124) );
  MX2X2 U65 ( .A(n1237), .B(data_in_2[133]), .S0(n1260), .Y(n1122) );
  MX2X2 U66 ( .A(n1238), .B(data_in_2[133]), .S0(n1288), .Y(n1123) );
  MX2X2 U67 ( .A(R4[14]), .B(data_in_2[14]), .S0(n1283), .Y(n1211) );
  MX2X2 U68 ( .A(R0[14]), .B(data_in_2[14]), .S0(n1256), .Y(n1210) );
  MX2X2 U69 ( .A(data_in_2[14]), .B(R8[14]), .S0(n1253), .Y(n1212) );
  MX2X2 U70 ( .A(data_in_2[84]), .B(n323), .S0(n44), .Y(n684) );
  MX2X2 U71 ( .A(data_in_2[62]), .B(R9[28]), .S0(n1254), .Y(n1203) );
  MX2X4 U72 ( .A(data_in_2[10]), .B(R12[10]), .S0(n1281), .Y(n1185) );
  MX2X4 U73 ( .A(data_in_2[10]), .B(R4[10]), .S0(n1289), .Y(n1184) );
  MX2X1 U74 ( .A(data_in_2[83]), .B(n458), .S0(n38), .Y(n669) );
  AOI22XL U75 ( .A0(n39), .A1(n1305), .B0(n1270), .B1(R0[32]), .Y(n992) );
  MX2X2 U76 ( .A(n100), .B(data_in_2[33]), .S0(n1251), .Y(n1188) );
  MX2X2 U77 ( .A(n61), .B(data_in_2[33]), .S0(n196), .Y(n1186) );
  MX2X2 U78 ( .A(n437), .B(data_in_2[130]), .S0(n1273), .Y(n1117) );
  MX2X2 U79 ( .A(n573), .B(data_in_2[130]), .S0(n1248), .Y(n977) );
  MX2X2 U80 ( .A(n301), .B(data_in_2[130]), .S0(n1260), .Y(n970) );
  MX2X2 U81 ( .A(n165), .B(data_in_2[130]), .S0(n1288), .Y(n972) );
  MX2X2 U82 ( .A(R12[14]), .B(data_in_2[14]), .S0(n1276), .Y(n1213) );
  MX2X4 U83 ( .A(data_in_2[45]), .B(R5[11]), .S0(n83), .Y(n1165) );
  MX2X4 U84 ( .A(data_in_2[45]), .B(R9[11]), .S0(n1255), .Y(n1166) );
  MX2X4 U85 ( .A(data_in_2[45]), .B(R13[11]), .S0(n84), .Y(n1167) );
  MX2X2 U86 ( .A(n289), .B(data_in_2[118]), .S0(n1261), .Y(n649) );
  MX2X2 U87 ( .A(n153), .B(data_in_2[118]), .S0(n1288), .Y(n650) );
  MX2X2 U88 ( .A(n1240), .B(data_in_2[100]), .S0(n105), .Y(n677) );
  MX2X2 U89 ( .A(n1239), .B(data_in_2[100]), .S0(n109), .Y(n676) );
  MX2X2 U90 ( .A(n1241), .B(data_in_2[100]), .S0(n1259), .Y(n674) );
  MX2X2 U91 ( .A(n1242), .B(data_in_2[100]), .S0(n1286), .Y(n675) );
  MX2X2 U92 ( .A(data_in_2[62]), .B(R13[28]), .S0(n1279), .Y(n1204) );
  MX2X2 U93 ( .A(n187), .B(data_in_2[84]), .S0(n1287), .Y(n685) );
  INVX1 U94 ( .A(n70), .Y(n72) );
  MX2X2 U95 ( .A(data_in_2[65]), .B(n73), .S0(n38), .Y(n1163) );
  MX2X2 U96 ( .A(data_in_2[65]), .B(n69), .S0(n17), .Y(n1161) );
  MX2X2 U97 ( .A(data_in_2[65]), .B(n68), .S0(n95), .Y(n1160) );
  MX2X4 U98 ( .A(data_in_2[31]), .B(R0[31]), .S0(n95), .Y(n1172) );
  MX2X4 U99 ( .A(data_in_2[31]), .B(R4[31]), .S0(n83), .Y(n1173) );
  MX2X2 U100 ( .A(data_in_2[65]), .B(n72), .S0(n1255), .Y(n1162) );
  MX2X2 U101 ( .A(data_in_2[30]), .B(R12[30]), .S0(n1280), .Y(n1183) );
  MX2X2 U102 ( .A(data_in_2[30]), .B(R0[30]), .S0(n1262), .Y(n1180) );
  MX2X2 U103 ( .A(data_in_2[30]), .B(R4[30]), .S0(n86), .Y(n1181) );
  MX2X2 U104 ( .A(data_in_2[67]), .B(n91), .S0(n86), .Y(n1143) );
  MX2X2 U105 ( .A(data_in_2[67]), .B(n92), .S0(n1282), .Y(n1145) );
  MX2X2 U106 ( .A(R8[30]), .B(data_in_2[30]), .S0(n1251), .Y(n1182) );
  MX2X2 U107 ( .A(data_in_2[67]), .B(n93), .S0(n1254), .Y(n1144) );
  AOI22XL U108 ( .A0(n91), .A1(n1299), .B0(n1268), .B1(n102), .Y(n1093) );
  AOI22XL U109 ( .A0(n92), .A1(n1303), .B0(n1269), .B1(R12[33]), .Y(n1025) );
  MX2X2 U110 ( .A(R13[29]), .B(data_in_2[63]), .S0(n1278), .Y(n1209) );
  MX2X2 U111 ( .A(R9[29]), .B(data_in_2[63]), .S0(n1243), .Y(n1208) );
  MX2X2 U112 ( .A(R1[29]), .B(data_in_2[63]), .S0(n1257), .Y(n1206) );
  MX2X2 U113 ( .A(R5[29]), .B(data_in_2[63]), .S0(n1284), .Y(n1207) );
  MX2X1 U114 ( .A(data_in_2[31]), .B(n75), .S0(n1280), .Y(n1175) );
  MX2X2 U115 ( .A(R4[29]), .B(data_in_2[29]), .S0(n1283), .Y(n1154) );
  MX2X2 U116 ( .A(R0[29]), .B(data_in_2[29]), .S0(n1256), .Y(n1153) );
  MX2X2 U117 ( .A(data_in_2[29]), .B(R12[29]), .S0(n104), .Y(n1156) );
  MX2X2 U118 ( .A(data_in_2[29]), .B(R8[29]), .S0(n1252), .Y(n1155) );
  MX2X2 U119 ( .A(data_in_2[32]), .B(R12[32]), .S0(n1280), .Y(n1171) );
  MX2X2 U120 ( .A(R4[32]), .B(data_in_2[32]), .S0(n1283), .Y(n1169) );
  MX2X1 U121 ( .A(n150), .B(data_in_2[115]), .S0(n1288), .Y(n671) );
  MX2X1 U122 ( .A(n286), .B(data_in_2[115]), .S0(n1261), .Y(n670) );
  MX2X1 U123 ( .A(n422), .B(data_in_2[115]), .S0(n1272), .Y(n673) );
  MX2X1 U124 ( .A(n558), .B(data_in_2[115]), .S0(n1247), .Y(n672) );
  MX2X1 U125 ( .A(n169), .B(data_in_2[134]), .S0(n1287), .Y(n652) );
  MX2X1 U126 ( .A(n305), .B(data_in_2[134]), .S0(n1260), .Y(n651) );
  MX2X1 U127 ( .A(n441), .B(data_in_2[134]), .S0(n1273), .Y(n654) );
  MX2X1 U128 ( .A(n577), .B(data_in_2[134]), .S0(n1248), .Y(n653) );
  MX2X2 U129 ( .A(n476), .B(data_in_2[101]), .S0(n1275), .Y(n648) );
  MX2X2 U130 ( .A(n204), .B(data_in_2[101]), .S0(n1286), .Y(n647) );
  MX2X2 U131 ( .A(n340), .B(data_in_2[101]), .S0(n1259), .Y(n646) );
  MX2X2 U132 ( .A(R8[32]), .B(data_in_2[32]), .S0(n1251), .Y(n1170) );
  MX2X2 U133 ( .A(R0[32]), .B(data_in_2[32]), .S0(n1256), .Y(n1168) );
  MX2X2 U134 ( .A(R13[13]), .B(data_in_2[47]), .S0(n1277), .Y(n1217) );
  MX2X2 U135 ( .A(R9[13]), .B(data_in_2[47]), .S0(n1246), .Y(n1216) );
  MX2X2 U136 ( .A(R1[13]), .B(data_in_2[47]), .S0(n1258), .Y(n1214) );
  MX2X2 U137 ( .A(R5[13]), .B(data_in_2[47]), .S0(n1285), .Y(n1215) );
  MX2X2 U138 ( .A(R1[28]), .B(data_in_2[62]), .S0(n1257), .Y(n1201) );
  MX2X2 U139 ( .A(R5[28]), .B(data_in_2[62]), .S0(n1284), .Y(n1202) );
  MX2X2 U140 ( .A(R13[14]), .B(data_in_2[48]), .S0(n1277), .Y(n1152) );
  MX2X2 U141 ( .A(R9[14]), .B(data_in_2[48]), .S0(n1249), .Y(n1151) );
  MX2X2 U142 ( .A(R1[14]), .B(data_in_2[48]), .S0(n1258), .Y(n1149) );
  MX2X2 U143 ( .A(R5[14]), .B(data_in_2[48]), .S0(n1285), .Y(n1150) );
  MX2X2 U144 ( .A(R13[16]), .B(data_in_2[50]), .S0(n1277), .Y(n1192) );
  MX2X2 U145 ( .A(R9[16]), .B(data_in_2[50]), .S0(n1250), .Y(n1191) );
  MX2X2 U146 ( .A(R1[16]), .B(data_in_2[50]), .S0(n1258), .Y(n1189) );
  MX2X2 U147 ( .A(R5[16]), .B(data_in_2[50]), .S0(n1285), .Y(n1190) );
  CLKINVX3 U148 ( .A(n1289), .Y(n1285) );
  CLKINVX3 U149 ( .A(n1289), .Y(n1286) );
  CLKINVX3 U150 ( .A(n1289), .Y(n1287) );
  CLKINVX3 U151 ( .A(n1289), .Y(n1284) );
  CLKINVX3 U152 ( .A(n1289), .Y(n1288) );
  INVX1 U153 ( .A(n1306), .Y(n1303) );
  INVX1 U154 ( .A(n1306), .Y(n1304) );
  INVX1 U155 ( .A(n1306), .Y(n1305) );
  INVX1 U156 ( .A(n1306), .Y(n1299) );
  INVX1 U157 ( .A(n1306), .Y(n1300) );
  INVX1 U158 ( .A(n1306), .Y(n1301) );
  INVX1 U159 ( .A(n1306), .Y(n1302) );
  CLKINVX3 U160 ( .A(n16), .Y(n1258) );
  CLKINVX3 U161 ( .A(n1262), .Y(n1261) );
  CLKINVX3 U162 ( .A(n1262), .Y(n1259) );
  CLKINVX3 U163 ( .A(n16), .Y(n1257) );
  CLKINVX3 U164 ( .A(n1262), .Y(n1260) );
  INVX1 U165 ( .A(n7), .Y(n1270) );
  INVX1 U166 ( .A(n7), .Y(n1263) );
  INVX1 U167 ( .A(n7), .Y(n1264) );
  INVX1 U168 ( .A(n7), .Y(n1265) );
  INVX1 U169 ( .A(n7), .Y(n1266) );
  INVX1 U170 ( .A(n7), .Y(n1267) );
  INVX1 U171 ( .A(n7), .Y(n1268) );
  INVX1 U172 ( .A(n7), .Y(n1269) );
  INVX1 U173 ( .A(n1314), .Y(n1312) );
  INVX1 U174 ( .A(n1314), .Y(n1311) );
  INVX1 U175 ( .A(n1314), .Y(n1309) );
  INVX1 U176 ( .A(n1314), .Y(n1308) );
  INVX1 U177 ( .A(n1314), .Y(n1313) );
  INVX1 U178 ( .A(n1314), .Y(n1310) );
  INVX1 U179 ( .A(n6), .Y(n1296) );
  INVX1 U180 ( .A(n6), .Y(n1297) );
  INVX1 U181 ( .A(n6), .Y(n1290) );
  INVX1 U182 ( .A(n6), .Y(n1291) );
  INVX1 U183 ( .A(n6), .Y(n1292) );
  INVX1 U184 ( .A(n6), .Y(n1294) );
  INVX1 U185 ( .A(n6), .Y(n1295) );
  INVX1 U186 ( .A(n6), .Y(n1293) );
  INVX1 U187 ( .A(n1282), .Y(n1271) );
  INVX1 U188 ( .A(n1282), .Y(n1274) );
  INVX1 U189 ( .A(n1254), .Y(n1244) );
  INVX1 U190 ( .A(n1279), .Y(n1278) );
  INVX1 U191 ( .A(n1252), .Y(n1245) );
  INVX1 U192 ( .A(n1252), .Y(n1250) );
  INVX1 U193 ( .A(n1282), .Y(n1272) );
  INVX1 U194 ( .A(n1254), .Y(n1243) );
  INVX1 U195 ( .A(n1279), .Y(n1276) );
  INVX1 U196 ( .A(n1280), .Y(n1277) );
  INVX1 U197 ( .A(n1254), .Y(n1246) );
  INVX1 U198 ( .A(n1252), .Y(n1247) );
  INVX1 U199 ( .A(n1253), .Y(n1249) );
  INVX1 U200 ( .A(n1279), .Y(n1273) );
  INVX1 U201 ( .A(n1253), .Y(n1248) );
  INVX1 U202 ( .A(n1252), .Y(n1251) );
  CLKINVX3 U203 ( .A(n1289), .Y(n1283) );
  INVX1 U204 ( .A(n969), .Y(n1289) );
  INVX1 U205 ( .A(n966), .Y(n1323) );
  NOR2X1 U206 ( .A(n973), .B(n1321), .Y(n969) );
  NOR2X1 U207 ( .A(n1321), .B(n1320), .Y(n964) );
  INVX1 U208 ( .A(n1306), .Y(n1298) );
  INVX1 U209 ( .A(n1314), .Y(n1307) );
  INVX1 U210 ( .A(n195), .Y(n1252) );
  INVX1 U211 ( .A(n195), .Y(n1255) );
  INVX1 U212 ( .A(n195), .Y(n1254) );
  INVX1 U213 ( .A(n195), .Y(n1253) );
  INVX1 U214 ( .A(n963), .Y(n1314) );
  INVX1 U215 ( .A(n967), .Y(n1306) );
  INVX1 U216 ( .A(n971), .Y(n1282) );
  INVX1 U217 ( .A(n971), .Y(n1281) );
  INVX1 U218 ( .A(n971), .Y(n1280) );
  INVX1 U219 ( .A(n971), .Y(n1279) );
  CLKINVX3 U220 ( .A(n1262), .Y(n1256) );
  INVX1 U221 ( .A(n196), .Y(n1262) );
  CLKINVX3 U222 ( .A(n1318), .Y(n1316) );
  CLKINVX3 U223 ( .A(n1318), .Y(n1315) );
  CLKINVX3 U224 ( .A(n1318), .Y(n1317) );
  OAI32X1 U225 ( .A0(n961), .A1(counter2[0]), .A2(n966), .B0(n1322), .B1(n1323), .Y(n1114) );
  NOR2X1 U226 ( .A(n961), .B(reg_flag_mux), .Y(n966) );
  OAI22X1 U227 ( .A0(n1320), .A1(n974), .B0(n961), .B1(n973), .Y(n1116) );
  NAND2BX1 U228 ( .AN(reg_datain_flag), .B(rst_n), .Y(n974) );
  OAI21XL U229 ( .A0(n1321), .A1(n974), .B0(n975), .Y(n1115) );
  OAI21XL U230 ( .A0(n1256), .A1(n1283), .B0(rst_n), .Y(n975) );
  OAI2BB2X1 U231 ( .B0(n965), .B1(n961), .A0N(counter2[1]), .A1N(n966), .Y(
        n1113) );
  AOI21X1 U232 ( .A0(n1303), .A1(n1323), .B0(n6), .Y(n965) );
  INVX1 U233 ( .A(n962), .Y(n1319) );
  AOI32X1 U234 ( .A0(reg_flag_mux), .A1(n1307), .A2(rst_n), .B0(n964), .B1(
        rst_n), .Y(n962) );
  AOI22X1 U235 ( .A0(n93), .A1(n1302), .B0(n1266), .B1(n100), .Y(n1059) );
  AOI22X1 U236 ( .A0(n97), .A1(n1305), .B0(n1270), .B1(n61), .Y(n991) );
  NOR2X1 U237 ( .A(n973), .B(counter1[1]), .Y(n971) );
  NOR2X1 U238 ( .A(n1322), .B(counter2[1]), .Y(n967) );
  NAND2X1 U239 ( .A(reg_datain_flag), .B(n1320), .Y(n973) );
  NAND2X1 U240 ( .A(counter2[1]), .B(counter2[0]), .Y(n963) );
  OAI221XL U241 ( .A0(n878), .A1(n1309), .B0(n844), .B1(n1296), .C0(n1013), 
        .Y(N63) );
  AOI22X1 U242 ( .A0(n63), .A1(n1303), .B0(n1263), .B1(R0[11]), .Y(n1013) );
  OAI221XL U243 ( .A0(n876), .A1(n1310), .B0(n842), .B1(n1296), .C0(n1011), 
        .Y(N65) );
  AOI22X1 U244 ( .A0(R1[13]), .A1(n1303), .B0(n1269), .B1(R0[13]), .Y(n1011)
         );
  OAI221XL U245 ( .A0(n875), .A1(n1311), .B0(n841), .B1(n1296), .C0(n1010), 
        .Y(N66) );
  AOI22X1 U246 ( .A0(R1[14]), .A1(n1303), .B0(n1270), .B1(R0[14]), .Y(n1010)
         );
  OAI221XL U247 ( .A0(n874), .A1(n1307), .B0(n840), .B1(n1296), .C0(n1009), 
        .Y(N67) );
  OAI221XL U248 ( .A0(n873), .A1(n1308), .B0(n839), .B1(n1296), .C0(n1008), 
        .Y(N68) );
  AOI22X1 U249 ( .A0(R1[16]), .A1(n1304), .B0(n1264), .B1(R0[16]), .Y(n1008)
         );
  OAI221XL U250 ( .A0(n861), .A1(n1310), .B0(n827), .B1(n1297), .C0(n996), .Y(
        N80) );
  AOI22X1 U251 ( .A0(R1[28]), .A1(n1304), .B0(n1265), .B1(R0[28]), .Y(n996) );
  OAI221XL U252 ( .A0(n860), .A1(n1311), .B0(n826), .B1(n1297), .C0(n995), .Y(
        N81) );
  AOI22X1 U253 ( .A0(R1[29]), .A1(n1305), .B0(n1269), .B1(R0[29]), .Y(n995) );
  OAI221XL U254 ( .A0(n859), .A1(n1308), .B0(n825), .B1(n1297), .C0(n994), .Y(
        N82) );
  AOI22X1 U255 ( .A0(R1[30]), .A1(n1305), .B0(n1265), .B1(R0[30]), .Y(n994) );
  OAI221XL U256 ( .A0(n858), .A1(n1312), .B0(n824), .B1(n1297), .C0(n993), .Y(
        N83) );
  OAI221XL U257 ( .A0(n857), .A1(n963), .B0(n823), .B1(n1297), .C0(n992), .Y(
        N84) );
  OAI221XL U258 ( .A0(n946), .A1(n1307), .B0(n912), .B1(n1291), .C0(n979), .Y(
        N97) );
  OAI221XL U259 ( .A0(n944), .A1(n1307), .B0(n910), .B1(n1292), .C0(n976), .Y(
        N99) );
  AOI22X1 U260 ( .A0(R5[13]), .A1(n1304), .B0(n1270), .B1(R4[13]), .Y(n976) );
  OAI221XL U261 ( .A0(n943), .A1(n1313), .B0(n909), .B1(n1290), .C0(n1112), 
        .Y(N100) );
  AOI22X1 U262 ( .A0(R5[14]), .A1(n1298), .B0(n1263), .B1(R4[14]), .Y(n1112)
         );
  OAI221XL U263 ( .A0(n942), .A1(n1307), .B0(n908), .B1(n1290), .C0(n1111), 
        .Y(N101) );
  OAI221XL U264 ( .A0(n941), .A1(n963), .B0(n907), .B1(n1290), .C0(n1110), .Y(
        N102) );
  AOI22X1 U265 ( .A0(R5[16]), .A1(n1298), .B0(n1263), .B1(n87), .Y(n1110) );
  OAI221XL U266 ( .A0(n929), .A1(n1313), .B0(n895), .B1(n1293), .C0(n1098), 
        .Y(N114) );
  AOI22X1 U267 ( .A0(R5[28]), .A1(n1299), .B0(n1265), .B1(R4[28]), .Y(n1098)
         );
  OAI221XL U268 ( .A0(n928), .A1(n1313), .B0(n894), .B1(n1294), .C0(n1097), 
        .Y(N115) );
  AOI22X1 U269 ( .A0(R5[29]), .A1(n1299), .B0(n1266), .B1(R4[29]), .Y(n1097)
         );
  OAI221XL U270 ( .A0(n927), .A1(n1313), .B0(n893), .B1(n1292), .C0(n1096), 
        .Y(N116) );
  AOI22X1 U271 ( .A0(R5[30]), .A1(n1299), .B0(n1267), .B1(R4[30]), .Y(n1096)
         );
  OAI221XL U272 ( .A0(n926), .A1(n1313), .B0(n892), .B1(n1293), .C0(n1095), 
        .Y(N117) );
  OAI221XL U273 ( .A0(n925), .A1(n1313), .B0(n891), .B1(n1294), .C0(n1094), 
        .Y(N118) );
  AOI22X1 U274 ( .A0(R5[32]), .A1(n1299), .B0(n1265), .B1(R4[32]), .Y(n1094)
         );
  OAI221XL U275 ( .A0(n708), .A1(n1312), .B0(n742), .B1(n1291), .C0(n1081), 
        .Y(N131) );
  OAI221XL U276 ( .A0(n706), .A1(n1311), .B0(n740), .B1(n1291), .C0(n1079), 
        .Y(N133) );
  AOI22X1 U277 ( .A0(R9[13]), .A1(n1300), .B0(n1264), .B1(R8[13]), .Y(n1079)
         );
  OAI221XL U278 ( .A0(n705), .A1(n1311), .B0(n739), .B1(n1291), .C0(n1078), 
        .Y(N134) );
  AOI22X1 U279 ( .A0(R9[14]), .A1(n1300), .B0(n1264), .B1(R8[14]), .Y(n1078)
         );
  OAI221XL U280 ( .A0(n704), .A1(n1311), .B0(n738), .B1(n1291), .C0(n1077), 
        .Y(N135) );
  AOI22X1 U281 ( .A0(R9[15]), .A1(n1300), .B0(n1264), .B1(R8[15]), .Y(n1077)
         );
  OAI221XL U282 ( .A0(n703), .A1(n1311), .B0(n737), .B1(n1292), .C0(n1076), 
        .Y(N136) );
  AOI22X1 U283 ( .A0(R9[16]), .A1(n1300), .B0(n1265), .B1(n90), .Y(n1076) );
  OAI221XL U284 ( .A0(n691), .A1(n1310), .B0(n725), .B1(n1293), .C0(n1064), 
        .Y(N148) );
  AOI22X1 U285 ( .A0(R9[28]), .A1(n1301), .B0(n1266), .B1(R8[28]), .Y(n1064)
         );
  OAI221XL U286 ( .A0(n690), .A1(n1310), .B0(n724), .B1(n1293), .C0(n1063), 
        .Y(N149) );
  AOI22X1 U287 ( .A0(R9[29]), .A1(n1301), .B0(n1266), .B1(R8[29]), .Y(n1063)
         );
  OAI221XL U288 ( .A0(n689), .A1(n1310), .B0(n723), .B1(n1293), .C0(n1062), 
        .Y(N150) );
  AOI22X1 U289 ( .A0(R9[30]), .A1(n1301), .B0(n1266), .B1(R8[30]), .Y(n1062)
         );
  OAI221XL U290 ( .A0(n688), .A1(n1310), .B0(n722), .B1(n1293), .C0(n1061), 
        .Y(N151) );
  AOI22X1 U291 ( .A0(n71), .A1(n1301), .B0(n1266), .B1(n77), .Y(n1061) );
  OAI221XL U292 ( .A0(n687), .A1(n1310), .B0(n721), .B1(n1293), .C0(n1060), 
        .Y(N152) );
  AOI22X1 U293 ( .A0(R9[32]), .A1(n1302), .B0(n1266), .B1(R8[32]), .Y(n1060)
         );
  OAI221XL U294 ( .A0(n810), .A1(n1309), .B0(n776), .B1(n1294), .C0(n1047), 
        .Y(N165) );
  OAI221XL U295 ( .A0(n808), .A1(n1309), .B0(n774), .B1(n1294), .C0(n1045), 
        .Y(N167) );
  AOI22X1 U296 ( .A0(R13[13]), .A1(n1301), .B0(n1267), .B1(R12[13]), .Y(n1045)
         );
  OAI221XL U297 ( .A0(n807), .A1(n1309), .B0(n773), .B1(n1294), .C0(n1044), 
        .Y(N168) );
  AOI22X1 U298 ( .A0(R13[14]), .A1(n1302), .B0(n1267), .B1(R12[14]), .Y(n1044)
         );
  OAI221XL U299 ( .A0(n806), .A1(n1309), .B0(n772), .B1(n1294), .C0(n1043), 
        .Y(N169) );
  AOI22X1 U300 ( .A0(R13[15]), .A1(n1301), .B0(n1267), .B1(R12[15]), .Y(n1043)
         );
  OAI221XL U301 ( .A0(n805), .A1(n1309), .B0(n771), .B1(n1294), .C0(n1042), 
        .Y(N170) );
  AOI22X1 U303 ( .A0(R13[16]), .A1(n1302), .B0(n1267), .B1(n89), .Y(n1042) );
  OAI221XL U304 ( .A0(n793), .A1(n1308), .B0(n759), .B1(n1295), .C0(n1030), 
        .Y(N182) );
  AOI22X1 U305 ( .A0(R13[28]), .A1(n1301), .B0(n1268), .B1(R12[28]), .Y(n1030)
         );
  OAI221XL U306 ( .A0(n792), .A1(n1308), .B0(n758), .B1(n1295), .C0(n1029), 
        .Y(N183) );
  AOI22X1 U307 ( .A0(R13[29]), .A1(n1300), .B0(n1268), .B1(R12[29]), .Y(n1029)
         );
  OAI221XL U308 ( .A0(n791), .A1(n1308), .B0(n757), .B1(n1297), .C0(n1028), 
        .Y(N184) );
  AOI22X1 U309 ( .A0(R13[30]), .A1(n1304), .B0(n1269), .B1(R12[30]), .Y(n1028)
         );
  OAI221XL U310 ( .A0(n790), .A1(n1309), .B0(n756), .B1(n1295), .C0(n1027), 
        .Y(N185) );
  AOI22X1 U311 ( .A0(n73), .A1(n1303), .B0(n1269), .B1(n75), .Y(n1027) );
  OAI221XL U312 ( .A0(n789), .A1(n1310), .B0(n755), .B1(n1296), .C0(n1026), 
        .Y(N186) );
  AOI22X1 U313 ( .A0(R13[32]), .A1(n1298), .B0(n1269), .B1(R12[32]), .Y(n1026)
         );
  OAI221XL U314 ( .A0(n889), .A1(n1311), .B0(n855), .B1(n1291), .C0(n1024), 
        .Y(N52) );
  AOI22X1 U315 ( .A0(R1[0]), .A1(n1299), .B0(n1269), .B1(R0[0]), .Y(n1024) );
  OAI221XL U316 ( .A0(n888), .A1(n1312), .B0(n854), .B1(n1294), .C0(n1023), 
        .Y(N53) );
  AOI22X1 U317 ( .A0(R1[1]), .A1(n1305), .B0(n1269), .B1(R0[1]), .Y(n1023) );
  OAI221XL U318 ( .A0(n887), .A1(n1313), .B0(n853), .B1(n1294), .C0(n1022), 
        .Y(N54) );
  AOI22X1 U319 ( .A0(R1[2]), .A1(n1303), .B0(n1269), .B1(R0[2]), .Y(n1022) );
  OAI221XL U320 ( .A0(n886), .A1(n1308), .B0(n852), .B1(n1292), .C0(n1021), 
        .Y(N55) );
  AOI22X1 U321 ( .A0(R1[3]), .A1(n1303), .B0(n1269), .B1(R0[3]), .Y(n1021) );
  OAI221XL U322 ( .A0(n885), .A1(n1313), .B0(n851), .B1(n1292), .C0(n1020), 
        .Y(N56) );
  AOI22X1 U323 ( .A0(R1[4]), .A1(n1303), .B0(n1269), .B1(R0[4]), .Y(n1020) );
  OAI221XL U324 ( .A0(n884), .A1(n1309), .B0(n850), .B1(n1293), .C0(n1019), 
        .Y(N57) );
  AOI22X1 U325 ( .A0(R1[5]), .A1(n1303), .B0(n1269), .B1(R0[5]), .Y(n1019) );
  OAI221XL U326 ( .A0(n883), .A1(n1310), .B0(n849), .B1(n1290), .C0(n1018), 
        .Y(N58) );
  AOI22X1 U327 ( .A0(R1[6]), .A1(n1303), .B0(n1269), .B1(R0[6]), .Y(n1018) );
  OAI221XL U328 ( .A0(n882), .A1(n1311), .B0(n848), .B1(n1297), .C0(n1017), 
        .Y(N59) );
  AOI22X1 U329 ( .A0(R1[7]), .A1(n1303), .B0(n1269), .B1(R0[7]), .Y(n1017) );
  OAI221XL U330 ( .A0(n881), .A1(n1312), .B0(n847), .B1(n1296), .C0(n1016), 
        .Y(N60) );
  AOI22X1 U331 ( .A0(R1[8]), .A1(n1303), .B0(n1263), .B1(R0[8]), .Y(n1016) );
  OAI221XL U332 ( .A0(n880), .A1(n1309), .B0(n846), .B1(n1296), .C0(n1015), 
        .Y(N61) );
  AOI22X1 U333 ( .A0(R1[9]), .A1(n1303), .B0(n1269), .B1(R0[9]), .Y(n1015) );
  OAI221XL U334 ( .A0(n879), .A1(n1312), .B0(n845), .B1(n1296), .C0(n1014), 
        .Y(N62) );
  AOI22X1 U335 ( .A0(R1[10]), .A1(n1303), .B0(n1270), .B1(n96), .Y(n1014) );
  OAI221XL U336 ( .A0(n877), .A1(n963), .B0(n843), .B1(n1296), .C0(n1012), .Y(
        N64) );
  AOI22X1 U337 ( .A0(R1[12]), .A1(n1303), .B0(n1267), .B1(R0[12]), .Y(n1012)
         );
  OAI221XL U338 ( .A0(n872), .A1(n963), .B0(n838), .B1(n1296), .C0(n1007), .Y(
        N69) );
  AOI22X1 U339 ( .A0(R1[17]), .A1(n1304), .B0(n1268), .B1(R0[17]), .Y(n1007)
         );
  OAI221XL U340 ( .A0(n871), .A1(n963), .B0(n837), .B1(n1296), .C0(n1006), .Y(
        N70) );
  AOI22X1 U341 ( .A0(R1[18]), .A1(n1304), .B0(n1265), .B1(R0[18]), .Y(n1006)
         );
  OAI221XL U342 ( .A0(n870), .A1(n963), .B0(n836), .B1(n1296), .C0(n1005), .Y(
        N71) );
  AOI22X1 U343 ( .A0(R1[19]), .A1(n1304), .B0(n1266), .B1(R0[19]), .Y(n1005)
         );
  OAI221XL U344 ( .A0(n869), .A1(n963), .B0(n835), .B1(n1297), .C0(n1004), .Y(
        N72) );
  AOI22X1 U345 ( .A0(R1[20]), .A1(n1304), .B0(n1266), .B1(R0[20]), .Y(n1004)
         );
  OAI221XL U346 ( .A0(n868), .A1(n963), .B0(n834), .B1(n1297), .C0(n1003), .Y(
        N73) );
  AOI22X1 U347 ( .A0(R1[21]), .A1(n1304), .B0(n1267), .B1(R0[21]), .Y(n1003)
         );
  OAI221XL U348 ( .A0(n867), .A1(n963), .B0(n833), .B1(n1297), .C0(n1002), .Y(
        N74) );
  AOI22X1 U349 ( .A0(R1[22]), .A1(n1304), .B0(n1264), .B1(R0[22]), .Y(n1002)
         );
  OAI221XL U350 ( .A0(n866), .A1(n963), .B0(n832), .B1(n1297), .C0(n1001), .Y(
        N75) );
  AOI22X1 U351 ( .A0(R1[23]), .A1(n1304), .B0(n1266), .B1(R0[23]), .Y(n1001)
         );
  OAI221XL U352 ( .A0(n865), .A1(n963), .B0(n831), .B1(n1297), .C0(n1000), .Y(
        N76) );
  AOI22X1 U353 ( .A0(R1[24]), .A1(n1304), .B0(n1267), .B1(R0[24]), .Y(n1000)
         );
  OAI221XL U354 ( .A0(n864), .A1(n963), .B0(n830), .B1(n1297), .C0(n999), .Y(
        N77) );
  AOI22X1 U355 ( .A0(R1[25]), .A1(n1304), .B0(n1264), .B1(R0[25]), .Y(n999) );
  OAI221XL U356 ( .A0(n863), .A1(n963), .B0(n829), .B1(n1297), .C0(n998), .Y(
        N78) );
  AOI22X1 U357 ( .A0(R1[26]), .A1(n1304), .B0(n1268), .B1(R0[26]), .Y(n998) );
  OAI221XL U358 ( .A0(n862), .A1(n963), .B0(n828), .B1(n1297), .C0(n997), .Y(
        N79) );
  AOI22X1 U359 ( .A0(R1[27]), .A1(n1304), .B0(n1263), .B1(R0[27]), .Y(n997) );
  OAI221XL U360 ( .A0(n957), .A1(n963), .B0(n923), .B1(n1295), .C0(n990), .Y(
        N86) );
  AOI22X1 U361 ( .A0(R5[0]), .A1(n1305), .B0(n1270), .B1(R4[0]), .Y(n990) );
  OAI221XL U362 ( .A0(n956), .A1(n1307), .B0(n922), .B1(n1296), .C0(n989), .Y(
        N87) );
  AOI22X1 U363 ( .A0(R5[1]), .A1(n1305), .B0(n1270), .B1(R4[1]), .Y(n989) );
  OAI221XL U364 ( .A0(n955), .A1(n1307), .B0(n921), .B1(n1290), .C0(n988), .Y(
        N88) );
  AOI22X1 U365 ( .A0(R5[2]), .A1(n1305), .B0(n1270), .B1(R4[2]), .Y(n988) );
  OAI221XL U366 ( .A0(n954), .A1(n1307), .B0(n920), .B1(n1291), .C0(n987), .Y(
        N89) );
  AOI22X1 U367 ( .A0(R5[3]), .A1(n1305), .B0(n1270), .B1(R4[3]), .Y(n987) );
  OAI221XL U368 ( .A0(n953), .A1(n1307), .B0(n919), .B1(n1297), .C0(n986), .Y(
        N90) );
  AOI22X1 U369 ( .A0(R5[4]), .A1(n1305), .B0(n1270), .B1(R4[4]), .Y(n986) );
  OAI221XL U370 ( .A0(n952), .A1(n1307), .B0(n918), .B1(n1295), .C0(n985), .Y(
        N91) );
  AOI22X1 U371 ( .A0(R5[5]), .A1(n1305), .B0(n1270), .B1(R4[5]), .Y(n985) );
  OAI221XL U372 ( .A0(n951), .A1(n1307), .B0(n917), .B1(n1296), .C0(n984), .Y(
        N92) );
  AOI22X1 U373 ( .A0(R5[6]), .A1(n1305), .B0(n1270), .B1(R4[6]), .Y(n984) );
  OAI221XL U374 ( .A0(n950), .A1(n1307), .B0(n916), .B1(n1290), .C0(n983), .Y(
        N93) );
  AOI22X1 U375 ( .A0(R5[7]), .A1(n1305), .B0(n1270), .B1(R4[7]), .Y(n983) );
  OAI221XL U376 ( .A0(n949), .A1(n1307), .B0(n915), .B1(n1290), .C0(n982), .Y(
        N94) );
  AOI22X1 U377 ( .A0(R5[8]), .A1(n1305), .B0(n1270), .B1(R4[8]), .Y(n982) );
  OAI221XL U378 ( .A0(n948), .A1(n1307), .B0(n914), .B1(n1291), .C0(n981), .Y(
        N95) );
  AOI22X1 U379 ( .A0(R5[9]), .A1(n1300), .B0(n1270), .B1(R4[9]), .Y(n981) );
  OAI221XL U380 ( .A0(n947), .A1(n1307), .B0(n913), .B1(n1293), .C0(n980), .Y(
        N96) );
  AOI22X1 U381 ( .A0(R5[10]), .A1(n1298), .B0(n1264), .B1(R4[10]), .Y(n980) );
  OAI221XL U382 ( .A0(n945), .A1(n1307), .B0(n911), .B1(n1294), .C0(n978), .Y(
        N98) );
  AOI22X1 U383 ( .A0(R5[12]), .A1(n1298), .B0(n1268), .B1(R4[12]), .Y(n978) );
  OAI221XL U384 ( .A0(n940), .A1(n1313), .B0(n906), .B1(n1290), .C0(n1109), 
        .Y(N103) );
  AOI22X1 U385 ( .A0(R5[17]), .A1(n1298), .B0(n1263), .B1(R4[17]), .Y(n1109)
         );
  OAI221XL U386 ( .A0(n939), .A1(n1307), .B0(n905), .B1(n1290), .C0(n1108), 
        .Y(N104) );
  AOI22X1 U387 ( .A0(R5[18]), .A1(n1298), .B0(n1263), .B1(R4[18]), .Y(n1108)
         );
  OAI221XL U388 ( .A0(n938), .A1(n963), .B0(n904), .B1(n1290), .C0(n1107), .Y(
        N105) );
  AOI22X1 U389 ( .A0(R5[19]), .A1(n1298), .B0(n1263), .B1(R4[19]), .Y(n1107)
         );
  OAI221XL U390 ( .A0(n937), .A1(n963), .B0(n903), .B1(n1290), .C0(n1106), .Y(
        N106) );
  AOI22X1 U391 ( .A0(R5[20]), .A1(n1298), .B0(n1263), .B1(R4[20]), .Y(n1106)
         );
  OAI221XL U392 ( .A0(n936), .A1(n1313), .B0(n902), .B1(n1290), .C0(n1105), 
        .Y(N107) );
  AOI22X1 U393 ( .A0(R5[21]), .A1(n1298), .B0(n1263), .B1(R4[21]), .Y(n1105)
         );
  OAI221XL U394 ( .A0(n935), .A1(n1313), .B0(n901), .B1(n1290), .C0(n1104), 
        .Y(N108) );
  AOI22X1 U395 ( .A0(R5[22]), .A1(n1298), .B0(n1263), .B1(R4[22]), .Y(n1104)
         );
  OAI221XL U396 ( .A0(n934), .A1(n1313), .B0(n900), .B1(n1290), .C0(n1103), 
        .Y(N109) );
  AOI22X1 U397 ( .A0(R5[23]), .A1(n1298), .B0(n1263), .B1(R4[23]), .Y(n1103)
         );
  OAI221XL U398 ( .A0(n933), .A1(n1313), .B0(n899), .B1(n1290), .C0(n1102), 
        .Y(N110) );
  AOI22X1 U399 ( .A0(R5[24]), .A1(n1298), .B0(n1263), .B1(R4[24]), .Y(n1102)
         );
  OAI221XL U400 ( .A0(n932), .A1(n1313), .B0(n898), .B1(n1290), .C0(n1101), 
        .Y(N111) );
  AOI22X1 U401 ( .A0(R5[25]), .A1(n1298), .B0(n1263), .B1(R4[25]), .Y(n1101)
         );
  OAI221XL U402 ( .A0(n931), .A1(n1313), .B0(n897), .B1(n1292), .C0(n1100), 
        .Y(N112) );
  AOI22X1 U403 ( .A0(R5[26]), .A1(n1298), .B0(n1263), .B1(R4[26]), .Y(n1100)
         );
  OAI221XL U404 ( .A0(n930), .A1(n1313), .B0(n896), .B1(n1290), .C0(n1099), 
        .Y(N113) );
  AOI22X1 U405 ( .A0(R5[27]), .A1(n1299), .B0(n1266), .B1(R4[27]), .Y(n1099)
         );
  OAI221XL U406 ( .A0(n719), .A1(n1312), .B0(n753), .B1(n1291), .C0(n1092), 
        .Y(N120) );
  AOI22X1 U407 ( .A0(R9[0]), .A1(n1299), .B0(n1267), .B1(R8[0]), .Y(n1092) );
  OAI221XL U408 ( .A0(n718), .A1(n1312), .B0(n752), .B1(n1297), .C0(n1091), 
        .Y(N121) );
  AOI22X1 U409 ( .A0(R9[1]), .A1(n1299), .B0(n1264), .B1(R8[1]), .Y(n1091) );
  OAI221XL U410 ( .A0(n717), .A1(n1312), .B0(n751), .B1(n1295), .C0(n1090), 
        .Y(N122) );
  AOI22X1 U411 ( .A0(R9[2]), .A1(n1299), .B0(n1268), .B1(R8[2]), .Y(n1090) );
  OAI221XL U412 ( .A0(n716), .A1(n1312), .B0(n750), .B1(n1296), .C0(n1089), 
        .Y(N123) );
  AOI22X1 U413 ( .A0(R9[3]), .A1(n1299), .B0(n1269), .B1(R8[3]), .Y(n1089) );
  OAI221XL U414 ( .A0(n715), .A1(n1312), .B0(n749), .B1(n1291), .C0(n1088), 
        .Y(N124) );
  AOI22X1 U415 ( .A0(R9[4]), .A1(n1299), .B0(n1264), .B1(R8[4]), .Y(n1088) );
  OAI221XL U416 ( .A0(n714), .A1(n1312), .B0(n748), .B1(n1291), .C0(n1087), 
        .Y(N125) );
  AOI22X1 U417 ( .A0(R9[5]), .A1(n1299), .B0(n1264), .B1(R8[5]), .Y(n1087) );
  OAI221XL U418 ( .A0(n713), .A1(n1312), .B0(n747), .B1(n1291), .C0(n1086), 
        .Y(N126) );
  AOI22X1 U419 ( .A0(R9[6]), .A1(n1300), .B0(n1264), .B1(R8[6]), .Y(n1086) );
  OAI221XL U420 ( .A0(n712), .A1(n1312), .B0(n746), .B1(n1291), .C0(n1085), 
        .Y(N127) );
  AOI22X1 U421 ( .A0(R9[7]), .A1(n1300), .B0(n1264), .B1(R8[7]), .Y(n1085) );
  OAI221XL U422 ( .A0(n711), .A1(n1312), .B0(n745), .B1(n1291), .C0(n1084), 
        .Y(N128) );
  AOI22X1 U423 ( .A0(R9[8]), .A1(n1300), .B0(n1264), .B1(R8[8]), .Y(n1084) );
  OAI221XL U424 ( .A0(n710), .A1(n1312), .B0(n744), .B1(n1291), .C0(n1083), 
        .Y(N129) );
  AOI22X1 U425 ( .A0(R9[9]), .A1(n1300), .B0(n1264), .B1(R8[9]), .Y(n1083) );
  OAI221XL U426 ( .A0(n709), .A1(n1312), .B0(n743), .B1(n1291), .C0(n1082), 
        .Y(N130) );
  AOI22X1 U427 ( .A0(R9[10]), .A1(n1300), .B0(n1264), .B1(n98), .Y(n1082) );
  OAI221XL U428 ( .A0(n707), .A1(n1312), .B0(n741), .B1(n1291), .C0(n1080), 
        .Y(N132) );
  AOI22X1 U429 ( .A0(R9[12]), .A1(n1300), .B0(n1264), .B1(R8[12]), .Y(n1080)
         );
  OAI221XL U430 ( .A0(n702), .A1(n1311), .B0(n736), .B1(n1292), .C0(n1075), 
        .Y(N137) );
  AOI22X1 U431 ( .A0(R9[17]), .A1(n1300), .B0(n1265), .B1(R8[17]), .Y(n1075)
         );
  OAI221XL U432 ( .A0(n701), .A1(n1311), .B0(n735), .B1(n1292), .C0(n1074), 
        .Y(N138) );
  AOI22X1 U433 ( .A0(R9[18]), .A1(n1300), .B0(n1265), .B1(R8[18]), .Y(n1074)
         );
  OAI221XL U434 ( .A0(n700), .A1(n1311), .B0(n734), .B1(n1292), .C0(n1073), 
        .Y(N139) );
  AOI22X1 U435 ( .A0(R9[19]), .A1(n1301), .B0(n1265), .B1(R8[19]), .Y(n1073)
         );
  OAI221XL U436 ( .A0(n699), .A1(n1311), .B0(n733), .B1(n1292), .C0(n1072), 
        .Y(N140) );
  AOI22X1 U437 ( .A0(R9[20]), .A1(n1301), .B0(n1265), .B1(R8[20]), .Y(n1072)
         );
  OAI221XL U438 ( .A0(n698), .A1(n1311), .B0(n732), .B1(n1292), .C0(n1071), 
        .Y(N141) );
  AOI22X1 U439 ( .A0(R9[21]), .A1(n1301), .B0(n1265), .B1(R8[21]), .Y(n1071)
         );
  OAI221XL U440 ( .A0(n697), .A1(n1311), .B0(n731), .B1(n1292), .C0(n1070), 
        .Y(N142) );
  AOI22X1 U441 ( .A0(R9[22]), .A1(n1301), .B0(n1265), .B1(R8[22]), .Y(n1070)
         );
  OAI221XL U442 ( .A0(n696), .A1(n1311), .B0(n730), .B1(n1292), .C0(n1069), 
        .Y(N143) );
  AOI22X1 U443 ( .A0(R9[23]), .A1(n1301), .B0(n1265), .B1(R8[23]), .Y(n1069)
         );
  OAI221XL U444 ( .A0(n695), .A1(n1311), .B0(n729), .B1(n1292), .C0(n1068), 
        .Y(N144) );
  AOI22X1 U445 ( .A0(R9[24]), .A1(n1301), .B0(n1265), .B1(R8[24]), .Y(n1068)
         );
  OAI221XL U446 ( .A0(n694), .A1(n1311), .B0(n728), .B1(n1292), .C0(n1067), 
        .Y(N145) );
  AOI22X1 U447 ( .A0(R9[25]), .A1(n1301), .B0(n1265), .B1(R8[25]), .Y(n1067)
         );
  OAI221XL U448 ( .A0(n693), .A1(n1310), .B0(n727), .B1(n1292), .C0(n1066), 
        .Y(N146) );
  AOI22X1 U449 ( .A0(R9[26]), .A1(n1301), .B0(n1265), .B1(R8[26]), .Y(n1066)
         );
  OAI221XL U450 ( .A0(n692), .A1(n1310), .B0(n726), .B1(n1292), .C0(n1065), 
        .Y(N147) );
  AOI22X1 U451 ( .A0(R9[27]), .A1(n1301), .B0(n1265), .B1(R8[27]), .Y(n1065)
         );
  OAI221XL U452 ( .A0(n821), .A1(n1310), .B0(n787), .B1(n1293), .C0(n1058), 
        .Y(N154) );
  AOI22X1 U453 ( .A0(R13[0]), .A1(n1302), .B0(n1266), .B1(R12[0]), .Y(n1058)
         );
  OAI221XL U454 ( .A0(n820), .A1(n1310), .B0(n786), .B1(n1293), .C0(n1057), 
        .Y(N155) );
  AOI22X1 U455 ( .A0(R13[1]), .A1(n1302), .B0(n1266), .B1(R12[1]), .Y(n1057)
         );
  OAI221XL U456 ( .A0(n819), .A1(n1310), .B0(n785), .B1(n1293), .C0(n1056), 
        .Y(N156) );
  AOI22X1 U457 ( .A0(R13[2]), .A1(n1302), .B0(n1266), .B1(R12[2]), .Y(n1056)
         );
  OAI221XL U458 ( .A0(n818), .A1(n1310), .B0(n784), .B1(n1293), .C0(n1055), 
        .Y(N157) );
  AOI22X1 U459 ( .A0(R13[3]), .A1(n1302), .B0(n1266), .B1(R12[3]), .Y(n1055)
         );
  OAI221XL U460 ( .A0(n817), .A1(n1310), .B0(n783), .B1(n1293), .C0(n1054), 
        .Y(N158) );
  AOI22X1 U461 ( .A0(R13[4]), .A1(n1302), .B0(n1266), .B1(R12[4]), .Y(n1054)
         );
  OAI221XL U462 ( .A0(n816), .A1(n1309), .B0(n782), .B1(n1293), .C0(n1053), 
        .Y(N159) );
  AOI22X1 U463 ( .A0(R13[5]), .A1(n1302), .B0(n1266), .B1(R12[5]), .Y(n1053)
         );
  OAI221XL U464 ( .A0(n815), .A1(n1309), .B0(n781), .B1(n1294), .C0(n1052), 
        .Y(N160) );
  AOI22X1 U465 ( .A0(R13[6]), .A1(n1302), .B0(n1267), .B1(R12[6]), .Y(n1052)
         );
  OAI221XL U466 ( .A0(n814), .A1(n1309), .B0(n780), .B1(n1294), .C0(n1051), 
        .Y(N161) );
  AOI22X1 U467 ( .A0(R13[7]), .A1(n1302), .B0(n1267), .B1(R12[7]), .Y(n1051)
         );
  OAI221XL U468 ( .A0(n813), .A1(n1309), .B0(n779), .B1(n1294), .C0(n1050), 
        .Y(N162) );
  AOI22X1 U469 ( .A0(R13[8]), .A1(n1302), .B0(n1267), .B1(R12[8]), .Y(n1050)
         );
  OAI221XL U470 ( .A0(n812), .A1(n1309), .B0(n778), .B1(n1294), .C0(n1049), 
        .Y(N163) );
  AOI22X1 U471 ( .A0(R13[9]), .A1(n1302), .B0(n1267), .B1(R12[9]), .Y(n1049)
         );
  OAI221XL U472 ( .A0(n811), .A1(n1309), .B0(n777), .B1(n1294), .C0(n1048), 
        .Y(N164) );
  AOI22X1 U473 ( .A0(R13[10]), .A1(n1302), .B0(n1267), .B1(R12[10]), .Y(n1048)
         );
  OAI221XL U474 ( .A0(n809), .A1(n1309), .B0(n775), .B1(n1294), .C0(n1046), 
        .Y(N166) );
  AOI22X1 U475 ( .A0(R13[12]), .A1(n1300), .B0(n1267), .B1(R12[12]), .Y(n1046)
         );
  OAI221XL U476 ( .A0(n804), .A1(n1309), .B0(n770), .B1(n1294), .C0(n1041), 
        .Y(N171) );
  AOI22X1 U477 ( .A0(R13[17]), .A1(n1304), .B0(n1267), .B1(R12[17]), .Y(n1041)
         );
  OAI221XL U478 ( .A0(n803), .A1(n1308), .B0(n769), .B1(n1295), .C0(n1040), 
        .Y(N172) );
  AOI22X1 U479 ( .A0(R13[18]), .A1(n1299), .B0(n1268), .B1(R12[18]), .Y(n1040)
         );
  OAI221XL U480 ( .A0(n802), .A1(n1308), .B0(n768), .B1(n1295), .C0(n1039), 
        .Y(N173) );
  AOI22X1 U481 ( .A0(R13[19]), .A1(n1302), .B0(n1268), .B1(R12[19]), .Y(n1039)
         );
  OAI221XL U482 ( .A0(n801), .A1(n1308), .B0(n767), .B1(n1295), .C0(n1038), 
        .Y(N174) );
  AOI22X1 U483 ( .A0(R13[20]), .A1(n1301), .B0(n1268), .B1(R12[20]), .Y(n1038)
         );
  OAI221XL U484 ( .A0(n800), .A1(n1308), .B0(n766), .B1(n1295), .C0(n1037), 
        .Y(N175) );
  AOI22X1 U485 ( .A0(R13[21]), .A1(n1300), .B0(n1268), .B1(R12[21]), .Y(n1037)
         );
  OAI221XL U486 ( .A0(n799), .A1(n1308), .B0(n765), .B1(n1295), .C0(n1036), 
        .Y(N176) );
  AOI22X1 U487 ( .A0(R13[22]), .A1(n1304), .B0(n1268), .B1(R12[22]), .Y(n1036)
         );
  OAI221XL U488 ( .A0(n798), .A1(n1308), .B0(n764), .B1(n1295), .C0(n1035), 
        .Y(N177) );
  AOI22X1 U489 ( .A0(R13[23]), .A1(n1299), .B0(n1268), .B1(R12[23]), .Y(n1035)
         );
  OAI221XL U490 ( .A0(n797), .A1(n1308), .B0(n763), .B1(n1295), .C0(n1034), 
        .Y(N178) );
  AOI22X1 U491 ( .A0(R13[24]), .A1(n1298), .B0(n1268), .B1(R12[24]), .Y(n1034)
         );
  OAI221XL U492 ( .A0(n796), .A1(n1308), .B0(n762), .B1(n1295), .C0(n1033), 
        .Y(N179) );
  AOI22X1 U493 ( .A0(R13[25]), .A1(n1299), .B0(n1268), .B1(R12[25]), .Y(n1033)
         );
  OAI221XL U494 ( .A0(n795), .A1(n1308), .B0(n761), .B1(n1295), .C0(n1032), 
        .Y(N180) );
  AOI22X1 U495 ( .A0(R13[26]), .A1(n1305), .B0(n1268), .B1(R12[26]), .Y(n1032)
         );
  OAI221XL U496 ( .A0(n794), .A1(n1308), .B0(n760), .B1(n1295), .C0(n1031), 
        .Y(N181) );
  AOI22X1 U497 ( .A0(R13[27]), .A1(n967), .B0(n1268), .B1(R12[27]), .Y(n1031)
         );
  AND2X2 U498 ( .A(reg_datain_flag), .B(n964), .Y(n195) );
  INVX1 U499 ( .A(counter1[1]), .Y(n1321) );
  INVX1 U500 ( .A(counter2[0]), .Y(n1322) );
  AND3X2 U501 ( .A(counter1[0]), .B(n1321), .C(reg_datain_flag), .Y(n196) );
  INVX1 U502 ( .A(reg_flag_mux), .Y(n1318) );
  OAI221XL U503 ( .A0(n686), .A1(n1310), .B0(n720), .B1(n1293), .C0(n1059), 
        .Y(N153) );
  OAI221XL U504 ( .A0(n788), .A1(n1308), .B0(n754), .B1(n1295), .C0(n1025), 
        .Y(N187) );
  OAI221XL U505 ( .A0(n856), .A1(n1313), .B0(n822), .B1(n1296), .C0(n991), .Y(
        N85) );
  OAI221XL U506 ( .A0(n924), .A1(n1313), .B0(n890), .B1(n1293), .C0(n1093), 
        .Y(N119) );
endmodule


module p_s ( clk, rst_n, data_in_3, p_s_flag_in, data_out_3 );
  input [135:0] data_in_3;
  output [33:0] data_out_3;
  input clk, rst_n, p_s_flag_in;
  wire   N26, N50, N52, N119, N120, N121, N122, N123, N124, N125, N126, N127,
         N128, N129, N130, N131, N132, N133, N134, N135, N136, N137, N138,
         N139, N140, N141, N142, N143, N144, N145, N146, N147, N148, N149,
         N150, N151, N152, n83, n86, n87, n100, n101, n105, n117, n119, n120,
         n121, n122, n134, n135, n138, n219, n222, n223, n236, n237, n239,
         n241, n253, n255, n256, n257, n258, n270, n271, n274, n355, n358,
         n359, n360, n372, n373, n375, n377, n389, n391, n392, n393, n394,
         n406, n407, n410, n411, n423, n426, n427, n440, n441, n445, n525,
         n527, n528, n529, n530, n542, n543, n546, n547, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n861, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n879, n882, n884, n886, n888,
         n889, n894, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n34, n40, n42, n43, n49, n50, n51,
         n53, n75, n76, n77, n78, n88, n89, n90, n91, n93, n95, n96, n97, n103,
         n104, n108, n109, n110, n111, n114, n116, n123, n125, n131, n133,
         n136, n137, n139, n141, n142, n143, n145, n146, n147, n149, n150,
         n151, n155, n156, n157, n158, n161, n162, n163, n225, n226, n227,
         n891, n892, n893, n895, n1165, n1166, n1167, n1168, n1169, n1170,
         n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
         n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
         n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
         n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
         n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
         n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
         n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
         n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
         n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
         n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
         n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
         n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
         n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
         n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406;
  wire   [1:0] counter_1;
  wire   [32:0] R0;
  wire   [30:0] R12;
  wire   [32:0] R1;
  wire   [30:0] R13;
  wire   [32:0] R2;
  wire   [32:0] R14;
  wire   [32:0] R3;
  wire   [30:0] R15;
  wire   [3:0] counter_2;

  AND2X2 U321 ( .A(n1157), .B(n869), .Y(n886) );
  AND2X2 U324 ( .A(counter_2[3]), .B(n861), .Y(n1157) );
  AND2X2 U326 ( .A(counter_2[3]), .B(counter_2[0]), .Y(n1158) );
  EDFFXL R12_reg_30_ ( .D(data_in_3[132]), .E(n1361), .CK(clk), .Q(R12[30]) );
  EDFFXL R13_reg_30_ ( .D(data_in_3[132]), .E(n1374), .CK(clk), .Q(R13[30]) );
  DFFHQXL R3_reg_11_ ( .D(n1304), .CK(clk), .Q(R3[11]) );
  DFFHQXL R2_reg_11_ ( .D(n1303), .CK(clk), .Q(R2[11]) );
  DFFHQXL R1_reg_11_ ( .D(n1302), .CK(clk), .Q(R1[11]) );
  DFFHQXL R0_reg_11_ ( .D(n1301), .CK(clk), .Q(R0[11]) );
  DFFHQXL R15_reg_9_ ( .D(n1298), .CK(clk), .Q(R15[9]) );
  DFFHQXL R14_reg_9_ ( .D(n1297), .CK(clk), .Q(R14[9]) );
  DFFHQXL R13_reg_9_ ( .D(n1296), .CK(clk), .Q(R13[9]) );
  DFFHQXL R12_reg_9_ ( .D(n1295), .CK(clk), .Q(R12[9]) );
  DFFHQXL R3_reg_14_ ( .D(n1294), .CK(clk), .Q(R3[14]) );
  DFFHQXL R2_reg_14_ ( .D(n1293), .CK(clk), .Q(R2[14]) );
  DFFHQXL R1_reg_14_ ( .D(n1292), .CK(clk), .Q(R1[14]) );
  DFFHQXL R0_reg_14_ ( .D(n1291), .CK(clk), .Q(R0[14]) );
  MX2X1 R15_reg_12__U3 ( .A(R15[12]), .B(data_in_3[114]), .S0(n1347), .Y(n1290) );
  DFFHQXL R15_reg_12_ ( .D(n1290), .CK(clk), .Q(R15[12]) );
  MX2X1 R13_reg_12__U3 ( .A(R13[12]), .B(data_in_3[114]), .S0(n1373), .Y(n1289) );
  DFFHQXL R13_reg_12_ ( .D(n1289), .CK(clk), .Q(R13[12]) );
  MX2X1 R12_reg_12__U3 ( .A(R12[12]), .B(data_in_3[114]), .S0(n1360), .Y(n1288) );
  DFFHQXL R12_reg_12_ ( .D(n1288), .CK(clk), .Q(R12[12]) );
  MX2X1 R3_reg_28__U3 ( .A(R3[28]), .B(data_in_3[28]), .S0(n1353), .Y(n1283)
         );
  DFFHQXL R3_reg_28_ ( .D(n1283), .CK(clk), .Q(R3[28]) );
  MX2X1 R2_reg_28__U3 ( .A(R2[28]), .B(data_in_3[28]), .S0(n1393), .Y(n1282)
         );
  DFFHQXL R2_reg_28_ ( .D(n1282), .CK(clk), .Q(R2[28]) );
  MX2X1 R1_reg_28__U3 ( .A(R1[28]), .B(data_in_3[28]), .S0(n1382), .Y(n1281)
         );
  DFFHQXL R1_reg_28_ ( .D(n1281), .CK(clk), .Q(R1[28]) );
  MX2X1 R0_reg_28__U3 ( .A(R0[28]), .B(data_in_3[28]), .S0(n1369), .Y(n1280)
         );
  DFFHQXL R0_reg_28_ ( .D(n1280), .CK(clk), .Q(R0[28]) );
  DFFHQXL R1_reg_15_ ( .D(n1279), .CK(clk), .Q(R1[15]) );
  DFFHQXL R14_reg_15_ ( .D(n1274), .CK(clk), .Q(R14[15]) );
  DFFHQXL R12_reg_15_ ( .D(n1272), .CK(clk), .Q(R12[15]) );
  DFFHQXL R15_reg_30_ ( .D(n1267), .CK(clk), .Q(R15[30]) );
  DFFHQXL R2_reg_10_ ( .D(n1266), .CK(clk), .Q(R2[10]) );
  DFFHQXL R3_reg_30_ ( .D(n1265), .CK(clk), .Q(R3[30]) );
  DFFHQXL R2_reg_30_ ( .D(n1264), .CK(clk), .Q(R2[30]) );
  DFFHQXL R1_reg_30_ ( .D(n1263), .CK(clk), .Q(R1[30]) );
  DFFHQXL R0_reg_30_ ( .D(n1262), .CK(clk), .Q(R0[30]) );
  DFFHQXL R2_reg_13_ ( .D(n1261), .CK(clk), .Q(R2[13]) );
  DFFHQXL R0_reg_13_ ( .D(n1260), .CK(clk), .Q(R0[13]) );
  MX2X1 R2_reg_31__U3 ( .A(n97), .B(data_in_3[31]), .S0(n1394), .Y(n1259) );
  MX2X1 R1_reg_31__U3 ( .A(n96), .B(data_in_3[31]), .S0(n1383), .Y(n1258) );
  MX2X1 R0_reg_31__U3 ( .A(n95), .B(data_in_3[31]), .S0(n1370), .Y(n1257) );
  DFFHQXL R3_reg_32_ ( .D(n1256), .CK(clk), .Q(R3[32]) );
  DFFHQXL R2_reg_32_ ( .D(n1255), .CK(clk), .Q(R2[32]) );
  DFFHQXL R1_reg_32_ ( .D(n1254), .CK(clk), .Q(R1[32]) );
  DFFHQXL R0_reg_32_ ( .D(n1253), .CK(clk), .Q(R0[32]) );
  MX2X1 R3_reg_27__U3 ( .A(R3[27]), .B(data_in_3[27]), .S0(n1352), .Y(n1252)
         );
  DFFHQXL R3_reg_27_ ( .D(n1252), .CK(clk), .Q(R3[27]) );
  MX2X1 R2_reg_27__U3 ( .A(R2[27]), .B(data_in_3[27]), .S0(n1393), .Y(n1251)
         );
  DFFHQXL R2_reg_27_ ( .D(n1251), .CK(clk), .Q(R2[27]) );
  MX2X1 R1_reg_27__U3 ( .A(R1[27]), .B(data_in_3[27]), .S0(n1382), .Y(n1250)
         );
  DFFHQXL R1_reg_27_ ( .D(n1250), .CK(clk), .Q(R1[27]) );
  MX2X1 R0_reg_27__U3 ( .A(R0[27]), .B(data_in_3[27]), .S0(n1369), .Y(n1249)
         );
  DFFHQXL R0_reg_27_ ( .D(n1249), .CK(clk), .Q(R0[27]) );
  DFFHQXL R3_reg_29_ ( .D(n1248), .CK(clk), .Q(R3[29]) );
  DFFHQXL R14_reg_13_ ( .D(n1244), .CK(clk), .Q(R14[13]) );
  DFFHQXL R14_reg_32_ ( .D(n1240), .CK(clk), .Q(R14[32]) );
  DFFHQXL R15_reg_11_ ( .D(n1236), .CK(clk), .Q(R15[11]) );
  DFFHQXL R14_reg_11_ ( .D(n1235), .CK(clk), .Q(R14[11]) );
  DFFHQXL R13_reg_11_ ( .D(n1234), .CK(clk), .Q(R13[11]) );
  DFFHQXL R12_reg_11_ ( .D(n1233), .CK(clk), .Q(R12[11]) );
  DFFHQXL R14_reg_14_ ( .D(n1231), .CK(clk), .Q(R14[14]) );
  MX2X1 R7_reg_13__U3 ( .A(n527), .B(data_in_3[47]), .S0(n1354), .Y(n1228) );
  DFFXL R7_reg_13_ ( .D(n1228), .CK(clk), .Q(n527), .QN(n605) );
  MX2X1 R6_reg_13__U3 ( .A(n391), .B(data_in_3[47]), .S0(n1386), .Y(n1227) );
  DFFXL R6_reg_13_ ( .D(n1227), .CK(clk), .Q(n391), .QN(n673) );
  MX2X1 R5_reg_13__U3 ( .A(n119), .B(data_in_3[47]), .S0(n1378), .Y(n1226) );
  DFFXL R5_reg_13_ ( .D(n1226), .CK(clk), .Q(n119), .QN(n809) );
  MX2X1 R4_reg_13__U3 ( .A(n255), .B(data_in_3[47]), .S0(n1365), .Y(n1225) );
  DFFXL R4_reg_13_ ( .D(n1225), .CK(clk), .Q(n255), .QN(n741) );
  MX2X1 R7_reg_29__U3 ( .A(n543), .B(data_in_3[63]), .S0(n1355), .Y(n1224) );
  DFFXL R7_reg_29_ ( .D(n1224), .CK(clk), .Q(n543), .QN(n589) );
  MX2X1 R6_reg_29__U3 ( .A(n407), .B(data_in_3[63]), .S0(n1387), .Y(n1223) );
  DFFXL R6_reg_29_ ( .D(n1223), .CK(clk), .Q(n407), .QN(n657) );
  MX2X1 R5_reg_29__U3 ( .A(n135), .B(data_in_3[63]), .S0(n1380), .Y(n1222) );
  DFFXL R5_reg_29_ ( .D(n1222), .CK(clk), .Q(n135), .QN(n793) );
  MX2X1 R4_reg_29__U3 ( .A(n271), .B(data_in_3[63]), .S0(n1367), .Y(n1221) );
  DFFXL R4_reg_29_ ( .D(n1221), .CK(clk), .Q(n271), .QN(n725) );
  MX2X1 R11_reg_11__U3 ( .A(n355), .B(data_in_3[79]), .S0(n1348), .Y(n1220) );
  DFFXL R11_reg_11_ ( .D(n1220), .CK(clk), .Q(n355), .QN(n709) );
  MX2X1 R10_reg_11__U3 ( .A(n423), .B(data_in_3[79]), .S0(n1388), .Y(n1219) );
  DFFXL R10_reg_11_ ( .D(n1219), .CK(clk), .Q(n423), .QN(n641) );
  MX2X1 R9_reg_11__U3 ( .A(n83), .B(data_in_3[79]), .S0(n1375), .Y(n1218) );
  DFFXL R9_reg_11_ ( .D(n1218), .CK(clk), .Q(n83), .QN(n845) );
  MX2X1 R8_reg_11__U3 ( .A(n219), .B(data_in_3[79]), .S0(n1362), .Y(n1217) );
  DFFXL R8_reg_11_ ( .D(n1217), .CK(clk), .Q(n219), .QN(n777) );
  MX2X1 R7_reg_28__U3 ( .A(n542), .B(data_in_3[62]), .S0(n1355), .Y(n1216) );
  DFFXL R7_reg_28_ ( .D(n1216), .CK(clk), .Q(n542), .QN(n590) );
  MX2X1 R6_reg_28__U3 ( .A(n406), .B(data_in_3[62]), .S0(n1387), .Y(n1215) );
  DFFXL R6_reg_28_ ( .D(n1215), .CK(clk), .Q(n406), .QN(n658) );
  MX2X1 R5_reg_28__U3 ( .A(n134), .B(data_in_3[62]), .S0(n1380), .Y(n1214) );
  DFFXL R5_reg_28_ ( .D(n1214), .CK(clk), .Q(n134), .QN(n794) );
  MX2X1 R4_reg_28__U3 ( .A(n270), .B(data_in_3[62]), .S0(n1367), .Y(n1213) );
  DFFXL R4_reg_28_ ( .D(n1213), .CK(clk), .Q(n270), .QN(n726) );
  DFFXL R11_reg_28_ ( .D(n1212), .CK(clk), .Q(n372), .QN(n692) );
  MX2X1 R10_reg_28__U3 ( .A(n440), .B(data_in_3[96]), .S0(n1390), .Y(n1211) );
  DFFXL R10_reg_28_ ( .D(n1211), .CK(clk), .Q(n440), .QN(n624) );
  MX2X1 R9_reg_28__U3 ( .A(n100), .B(data_in_3[96]), .S0(n1377), .Y(n1210) );
  DFFXL R9_reg_28_ ( .D(n1210), .CK(clk), .Q(n100), .QN(n828) );
  DFFXL R8_reg_28_ ( .D(n1209), .CK(clk), .Q(n236), .QN(n760) );
  MX2X1 R7_reg_16__U3 ( .A(n530), .B(data_in_3[50]), .S0(n1354), .Y(n1208) );
  DFFXL R7_reg_16_ ( .D(n1208), .CK(clk), .Q(n530), .QN(n602) );
  MX2X1 R6_reg_16__U3 ( .A(n394), .B(data_in_3[50]), .S0(n1386), .Y(n1207) );
  DFFXL R6_reg_16_ ( .D(n1207), .CK(clk), .Q(n394), .QN(n670) );
  MX2X1 R5_reg_16__U3 ( .A(n122), .B(data_in_3[50]), .S0(n1379), .Y(n1206) );
  DFFXL R5_reg_16_ ( .D(n1206), .CK(clk), .Q(n122), .QN(n806) );
  MX2X1 R4_reg_16__U3 ( .A(n258), .B(data_in_3[50]), .S0(n1366), .Y(n1205) );
  DFFXL R4_reg_16_ ( .D(n1205), .CK(clk), .Q(n258), .QN(n738) );
  DFFXL R11_reg_16_ ( .D(n1204), .CK(clk), .Q(n360), .QN(n704) );
  DFFXL R11_reg_30_ ( .D(n1203), .CK(clk), .Q(n1306), .QN(n690) );
  MX2X1 R10_reg_30__U3 ( .A(n1305), .B(data_in_3[98]), .S0(n1390), .Y(n1202)
         );
  DFFXL R10_reg_30_ ( .D(n1202), .CK(clk), .Q(n1305), .QN(n622) );
  MX2X1 R9_reg_30__U3 ( .A(n1308), .B(data_in_3[98]), .S0(n1377), .Y(n1201) );
  DFFXL R9_reg_30_ ( .D(n1201), .CK(clk), .Q(n1308), .QN(n826) );
  MX2X1 R8_reg_30__U3 ( .A(n1307), .B(data_in_3[98]), .S0(n1364), .Y(n1200) );
  DFFXL R8_reg_30_ ( .D(n1200), .CK(clk), .Q(n1307), .QN(n758) );
  DFFXL R7_reg_11_ ( .D(n1199), .CK(clk), .Q(n525), .QN(n607) );
  DFFXL R6_reg_11_ ( .D(n1198), .CK(clk), .Q(n389), .QN(n675) );
  DFFXL R5_reg_11_ ( .D(n1197), .CK(clk), .Q(n117), .QN(n811) );
  DFFXL R4_reg_11_ ( .D(n1196), .CK(clk), .Q(n253), .QN(n743) );
  DFFXL R10_reg_32_ ( .D(n1195), .CK(clk), .Q(n1311), .QN(n620) );
  DFFXL R9_reg_32_ ( .D(n1194), .CK(clk), .Q(n1313), .QN(n824) );
  DFFXL R8_reg_32_ ( .D(n1193), .CK(clk), .Q(n1312), .QN(n756) );
  MX2X1 R7_reg_14__U3 ( .A(n528), .B(data_in_3[48]), .S0(n1354), .Y(n1192) );
  DFFXL R7_reg_14_ ( .D(n1192), .CK(clk), .Q(n528), .QN(n604) );
  MX2X1 R6_reg_14__U3 ( .A(n392), .B(data_in_3[48]), .S0(n1386), .Y(n1191) );
  DFFXL R6_reg_14_ ( .D(n1191), .CK(clk), .Q(n392), .QN(n672) );
  MX2X1 R5_reg_14__U3 ( .A(n120), .B(data_in_3[48]), .S0(n1378), .Y(n1190) );
  DFFXL R5_reg_14_ ( .D(n1190), .CK(clk), .Q(n120), .QN(n808) );
  MX2X1 R4_reg_14__U3 ( .A(n256), .B(data_in_3[48]), .S0(n1365), .Y(n1189) );
  DFFXL R4_reg_14_ ( .D(n1189), .CK(clk), .Q(n256), .QN(n740) );
  MX2X1 R7_reg_32__U3 ( .A(n546), .B(data_in_3[66]), .S0(n1356), .Y(n1188) );
  DFFXL R7_reg_32_ ( .D(n1188), .CK(clk), .Q(n546), .QN(n586) );
  MX2X1 R6_reg_32__U3 ( .A(n410), .B(data_in_3[66]), .S0(n1387), .Y(n1187) );
  DFFXL R6_reg_32_ ( .D(n1187), .CK(clk), .Q(n410), .QN(n654) );
  MX2X1 R5_reg_32__U3 ( .A(n138), .B(data_in_3[66]), .S0(n1380), .Y(n1186) );
  DFFXL R5_reg_32_ ( .D(n1186), .CK(clk), .Q(n138), .QN(n790) );
  MX2X1 R4_reg_32__U3 ( .A(n274), .B(data_in_3[66]), .S0(n1367), .Y(n1185) );
  DFFXL R4_reg_32_ ( .D(n1185), .CK(clk), .Q(n274), .QN(n722) );
  DFFXL R11_reg_15_ ( .D(n1184), .CK(clk), .Q(n359), .QN(n705) );
  MX2X1 R10_reg_15__U3 ( .A(n427), .B(data_in_3[83]), .S0(n1389), .Y(n1183) );
  DFFXL R10_reg_15_ ( .D(n1183), .CK(clk), .Q(n427), .QN(n637) );
  MX2X1 R9_reg_15__U3 ( .A(n87), .B(data_in_3[83]), .S0(n1376), .Y(n1182) );
  DFFXL R9_reg_15_ ( .D(n1182), .CK(clk), .Q(n87), .QN(n841) );
  MX2X1 R8_reg_15__U3 ( .A(n223), .B(data_in_3[83]), .S0(n1363), .Y(n1181) );
  DFFXL R8_reg_15_ ( .D(n1181), .CK(clk), .Q(n223), .QN(n773) );
  MX2X1 R11_reg_14__U3 ( .A(n358), .B(data_in_3[82]), .S0(n1349), .Y(n1180) );
  DFFXL R11_reg_14_ ( .D(n1180), .CK(clk), .Q(n358), .QN(n706) );
  MX2X1 R10_reg_14__U3 ( .A(n426), .B(data_in_3[82]), .S0(n1389), .Y(n1179) );
  DFFXL R10_reg_14_ ( .D(n1179), .CK(clk), .Q(n426), .QN(n638) );
  MX2X1 R9_reg_14__U3 ( .A(n86), .B(data_in_3[82]), .S0(n1376), .Y(n1178) );
  DFFXL R9_reg_14_ ( .D(n1178), .CK(clk), .Q(n86), .QN(n842) );
  MX2X1 R8_reg_14__U3 ( .A(n222), .B(data_in_3[82]), .S0(n1363), .Y(n1177) );
  DFFXL R8_reg_14_ ( .D(n1177), .CK(clk), .Q(n222), .QN(n774) );
  DFFXL R7_reg_15_ ( .D(n1176), .CK(clk), .Q(n529), .QN(n603) );
  DFFXL R6_reg_15_ ( .D(n1175), .CK(clk), .Q(n393), .QN(n671) );
  DFFXL R5_reg_15_ ( .D(n1174), .CK(clk), .Q(n121), .QN(n807) );
  DFFXL R4_reg_15_ ( .D(n1173), .CK(clk), .Q(n257), .QN(n739) );
  DFFXL R7_reg_33_ ( .D(n1172), .CK(clk), .Q(n547), .QN(n585) );
  DFFXL R6_reg_33_ ( .D(n1171), .CK(clk), .Q(n411), .QN(n653) );
  DFFXL R11_reg_31_ ( .D(n1170), .CK(clk), .Q(n375), .QN(n689) );
  DFFXL R8_reg_31_ ( .D(n1169), .CK(clk), .Q(n239), .QN(n757) );
  DFFXL R11_reg_29_ ( .D(n1168), .CK(clk), .Q(n373), .QN(n691) );
  MX2X1 R10_reg_29__U3 ( .A(n441), .B(data_in_3[97]), .S0(n1390), .Y(n1167) );
  DFFXL R10_reg_29_ ( .D(n1167), .CK(clk), .Q(n441), .QN(n623) );
  MX2X1 R9_reg_29__U3 ( .A(n101), .B(data_in_3[97]), .S0(n1377), .Y(n1166) );
  DFFXL R9_reg_29_ ( .D(n1166), .CK(clk), .Q(n101), .QN(n827) );
  MX2X1 R8_reg_29__U3 ( .A(n237), .B(data_in_3[97]), .S0(n1364), .Y(n1165) );
  DFFXL R8_reg_29_ ( .D(n1165), .CK(clk), .Q(n237), .QN(n759) );
  DFFXL R11_reg_33_ ( .D(n895), .CK(clk), .Q(n377), .QN(n687) );
  DFFXL R10_reg_33_ ( .D(n893), .CK(clk), .Q(n445), .QN(n619) );
  DFFXL R9_reg_33_ ( .D(n892), .CK(clk), .Q(n105), .QN(n823) );
  DFFXL R8_reg_33_ ( .D(n891), .CK(clk), .Q(n241), .QN(n755) );
  EDFFX1 R7_reg_26_ ( .D(data_in_3[60]), .E(n1355), .CK(clk), .QN(n592) );
  EDFFX1 R7_reg_25_ ( .D(data_in_3[59]), .E(n1355), .CK(clk), .QN(n593) );
  EDFFX1 R7_reg_24_ ( .D(data_in_3[58]), .E(n1355), .CK(clk), .QN(n594) );
  EDFFX1 R7_reg_21_ ( .D(data_in_3[55]), .E(n1355), .CK(clk), .QN(n597) );
  EDFFXL R7_reg_20_ ( .D(data_in_3[54]), .E(n1355), .CK(clk), .QN(n598) );
  EDFFXL R7_reg_19_ ( .D(data_in_3[53]), .E(n1355), .CK(clk), .QN(n599) );
  EDFFX1 R7_reg_18_ ( .D(data_in_3[52]), .E(n1355), .CK(clk), .QN(n600) );
  EDFFX1 R7_reg_17_ ( .D(data_in_3[51]), .E(n1354), .CK(clk), .QN(n601) );
  EDFFX1 R7_reg_9_ ( .D(data_in_3[43]), .E(n1354), .CK(clk), .QN(n609) );
  EDFFX1 R7_reg_8_ ( .D(data_in_3[42]), .E(n1354), .CK(clk), .QN(n610) );
  EDFFX1 R7_reg_6_ ( .D(data_in_3[40]), .E(n1354), .CK(clk), .QN(n612) );
  EDFFX1 R7_reg_5_ ( .D(data_in_3[39]), .E(n1353), .CK(clk), .QN(n613) );
  EDFFX1 R7_reg_4_ ( .D(data_in_3[38]), .E(n1353), .CK(clk), .QN(n614) );
  EDFFX1 R7_reg_3_ ( .D(data_in_3[37]), .E(n1353), .CK(clk), .QN(n615) );
  EDFFXL R7_reg_2_ ( .D(data_in_3[36]), .E(n1353), .CK(clk), .QN(n616) );
  EDFFX1 R7_reg_1_ ( .D(data_in_3[35]), .E(n1353), .CK(clk), .QN(n617) );
  EDFFX1 R7_reg_0_ ( .D(data_in_3[34]), .E(n1353), .CK(clk), .QN(n618) );
  EDFFX1 R6_reg_26_ ( .D(data_in_3[60]), .E(n1387), .CK(clk), .QN(n660) );
  EDFFX1 R6_reg_25_ ( .D(data_in_3[59]), .E(n1387), .CK(clk), .QN(n661) );
  EDFFX1 R6_reg_24_ ( .D(data_in_3[58]), .E(n1387), .CK(clk), .QN(n662) );
  EDFFX1 R6_reg_23_ ( .D(data_in_3[57]), .E(n1386), .CK(clk), .QN(n663) );
  EDFFX1 R6_reg_21_ ( .D(data_in_3[55]), .E(n1386), .CK(clk), .QN(n665) );
  EDFFXL R6_reg_20_ ( .D(data_in_3[54]), .E(n1386), .CK(clk), .QN(n666) );
  EDFFXL R6_reg_19_ ( .D(data_in_3[53]), .E(n1386), .CK(clk), .QN(n667) );
  EDFFX1 R6_reg_18_ ( .D(data_in_3[52]), .E(n1386), .CK(clk), .QN(n668) );
  EDFFX1 R6_reg_17_ ( .D(data_in_3[51]), .E(n1386), .CK(clk), .QN(n669) );
  EDFFX1 R6_reg_9_ ( .D(data_in_3[43]), .E(n1385), .CK(clk), .QN(n677) );
  EDFFX1 R6_reg_8_ ( .D(data_in_3[42]), .E(n1385), .CK(clk), .QN(n678) );
  EDFFX1 R6_reg_6_ ( .D(data_in_3[40]), .E(n1385), .CK(clk), .QN(n680) );
  EDFFX1 R6_reg_5_ ( .D(data_in_3[39]), .E(n1385), .CK(clk), .QN(n681) );
  EDFFX1 R6_reg_4_ ( .D(data_in_3[38]), .E(n1385), .CK(clk), .QN(n682) );
  EDFFX1 R6_reg_3_ ( .D(data_in_3[37]), .E(n1385), .CK(clk), .QN(n683) );
  EDFFXL R6_reg_2_ ( .D(data_in_3[36]), .E(n1385), .CK(clk), .QN(n684) );
  EDFFX1 R6_reg_1_ ( .D(data_in_3[35]), .E(n1385), .CK(clk), .QN(n685) );
  EDFFX1 R6_reg_0_ ( .D(data_in_3[34]), .E(n1385), .CK(clk), .QN(n686) );
  EDFFX1 R4_reg_26_ ( .D(data_in_3[60]), .E(n1366), .CK(clk), .QN(n728) );
  EDFFX1 R4_reg_25_ ( .D(data_in_3[59]), .E(n1366), .CK(clk), .QN(n729) );
  EDFFX1 R4_reg_24_ ( .D(data_in_3[58]), .E(n1366), .CK(clk), .QN(n730) );
  EDFFX1 R4_reg_23_ ( .D(data_in_3[57]), .E(n1366), .CK(clk), .QN(n731) );
  EDFFX1 R4_reg_21_ ( .D(data_in_3[55]), .E(n1366), .CK(clk), .QN(n733) );
  EDFFXL R4_reg_20_ ( .D(data_in_3[54]), .E(n1366), .CK(clk), .QN(n734) );
  EDFFXL R4_reg_19_ ( .D(data_in_3[53]), .E(n1366), .CK(clk), .QN(n735) );
  EDFFX1 R4_reg_18_ ( .D(data_in_3[52]), .E(n1366), .CK(clk), .QN(n736) );
  EDFFX1 R4_reg_17_ ( .D(data_in_3[51]), .E(n1366), .CK(clk), .QN(n737) );
  EDFFX1 R4_reg_9_ ( .D(data_in_3[43]), .E(n1365), .CK(clk), .QN(n745) );
  EDFFX1 R4_reg_8_ ( .D(data_in_3[42]), .E(n1365), .CK(clk), .QN(n746) );
  EDFFX1 R4_reg_6_ ( .D(data_in_3[40]), .E(n1365), .CK(clk), .QN(n748) );
  EDFFX1 R4_reg_5_ ( .D(data_in_3[39]), .E(n1365), .CK(clk), .QN(n749) );
  EDFFX1 R4_reg_4_ ( .D(data_in_3[38]), .E(n1365), .CK(clk), .QN(n750) );
  EDFFX1 R4_reg_3_ ( .D(data_in_3[37]), .E(n1364), .CK(clk), .QN(n751) );
  EDFFXL R4_reg_2_ ( .D(data_in_3[36]), .E(n1364), .CK(clk), .QN(n752) );
  EDFFX1 R4_reg_1_ ( .D(data_in_3[35]), .E(n1364), .CK(clk), .QN(n753) );
  EDFFX1 R4_reg_0_ ( .D(data_in_3[34]), .E(n1364), .CK(clk), .QN(n754) );
  EDFFXL R5_reg_30_ ( .D(data_in_3[64]), .E(n1380), .CK(clk), .QN(n792) );
  EDFFXL R5_reg_27_ ( .D(data_in_3[61]), .E(n1379), .CK(clk), .QN(n795) );
  EDFFXL R5_reg_26_ ( .D(data_in_3[60]), .E(n1379), .CK(clk), .QN(n796) );
  EDFFXL R5_reg_25_ ( .D(data_in_3[59]), .E(n1379), .CK(clk), .QN(n797) );
  EDFFXL R5_reg_24_ ( .D(data_in_3[58]), .E(n1379), .CK(clk), .QN(n798) );
  EDFFXL R5_reg_23_ ( .D(data_in_3[57]), .E(n1379), .CK(clk), .QN(n799) );
  EDFFXL R5_reg_22_ ( .D(data_in_3[56]), .E(n1379), .CK(clk), .QN(n800) );
  EDFFXL R5_reg_21_ ( .D(data_in_3[55]), .E(n1379), .CK(clk), .QN(n801) );
  EDFFXL R5_reg_20_ ( .D(data_in_3[54]), .E(n1379), .CK(clk), .QN(n802) );
  EDFFXL R5_reg_19_ ( .D(data_in_3[53]), .E(n1379), .CK(clk), .QN(n803) );
  EDFFXL R5_reg_12_ ( .D(data_in_3[46]), .E(n1378), .CK(clk), .QN(n810) );
  EDFFXL R5_reg_10_ ( .D(data_in_3[44]), .E(n1378), .CK(clk), .QN(n812) );
  EDFFXL R5_reg_9_ ( .D(n53), .E(n1378), .CK(clk), .QN(n813) );
  EDFFXL R5_reg_8_ ( .D(data_in_3[42]), .E(n1378), .CK(clk), .QN(n814) );
  EDFFXL R5_reg_7_ ( .D(data_in_3[41]), .E(n1378), .CK(clk), .QN(n815) );
  EDFFXL R5_reg_6_ ( .D(data_in_3[40]), .E(n1378), .CK(clk), .QN(n816) );
  EDFFXL R5_reg_5_ ( .D(data_in_3[39]), .E(n1378), .CK(clk), .QN(n817) );
  EDFFXL R5_reg_4_ ( .D(data_in_3[38]), .E(n1378), .CK(clk), .QN(n818) );
  EDFFXL R5_reg_3_ ( .D(data_in_3[37]), .E(n1377), .CK(clk), .QN(n819) );
  EDFFXL R5_reg_2_ ( .D(data_in_3[36]), .E(n1377), .CK(clk), .QN(n820) );
  EDFFXL R10_reg_27_ ( .D(data_in_3[95]), .E(n1390), .CK(clk), .QN(n625) );
  EDFFXL R10_reg_26_ ( .D(data_in_3[94]), .E(n1390), .CK(clk), .QN(n626) );
  EDFFXL R10_reg_25_ ( .D(data_in_3[93]), .E(n1389), .CK(clk), .QN(n627) );
  EDFFXL R10_reg_24_ ( .D(data_in_3[92]), .E(n1389), .CK(clk), .QN(n628) );
  EDFFXL R10_reg_23_ ( .D(data_in_3[91]), .E(n1389), .CK(clk), .QN(n629) );
  EDFFXL R10_reg_22_ ( .D(data_in_3[90]), .E(n1389), .CK(clk), .QN(n630) );
  EDFFXL R10_reg_21_ ( .D(data_in_3[89]), .E(n1389), .CK(clk), .QN(n631) );
  EDFFXL R10_reg_20_ ( .D(data_in_3[88]), .E(n1389), .CK(clk), .QN(n632) );
  EDFFXL R10_reg_19_ ( .D(data_in_3[87]), .E(n1389), .CK(clk), .QN(n633) );
  EDFFX1 R10_reg_18_ ( .D(data_in_3[86]), .E(n1389), .CK(clk), .QN(n634) );
  EDFFX1 R10_reg_17_ ( .D(data_in_3[85]), .E(n1389), .CK(clk), .QN(n635) );
  EDFFXL R10_reg_12_ ( .D(data_in_3[80]), .E(n1388), .CK(clk), .QN(n640) );
  EDFFXL R10_reg_10_ ( .D(data_in_3[78]), .E(n1388), .CK(clk), .QN(n642) );
  EDFFXL R10_reg_9_ ( .D(data_in_3[77]), .E(n1388), .CK(clk), .QN(n643) );
  EDFFXL R10_reg_8_ ( .D(data_in_3[76]), .E(n1388), .CK(clk), .QN(n644) );
  EDFFXL R10_reg_7_ ( .D(data_in_3[75]), .E(n1388), .CK(clk), .QN(n645) );
  EDFFXL R10_reg_6_ ( .D(data_in_3[74]), .E(n1388), .CK(clk), .QN(n646) );
  EDFFXL R10_reg_5_ ( .D(data_in_3[73]), .E(n1388), .CK(clk), .QN(n647) );
  EDFFXL R10_reg_4_ ( .D(data_in_3[72]), .E(n1388), .CK(clk), .QN(n648) );
  EDFFXL R10_reg_3_ ( .D(data_in_3[71]), .E(n1388), .CK(clk), .QN(n649) );
  EDFFXL R10_reg_2_ ( .D(data_in_3[70]), .E(n1388), .CK(clk), .QN(n650) );
  EDFFXL R10_reg_1_ ( .D(data_in_3[69]), .E(n1387), .CK(clk), .QN(n651) );
  EDFFX1 R10_reg_0_ ( .D(data_in_3[68]), .E(n1387), .CK(clk), .QN(n652) );
  EDFFXL R11_reg_27_ ( .D(data_in_3[95]), .E(n1350), .CK(clk), .QN(n693) );
  EDFFXL R11_reg_26_ ( .D(data_in_3[94]), .E(n1350), .CK(clk), .QN(n694) );
  EDFFXL R11_reg_25_ ( .D(data_in_3[93]), .E(n1349), .CK(clk), .QN(n695) );
  EDFFXL R11_reg_24_ ( .D(data_in_3[92]), .E(n1349), .CK(clk), .QN(n696) );
  EDFFXL R11_reg_23_ ( .D(data_in_3[91]), .E(n1349), .CK(clk), .QN(n697) );
  EDFFXL R11_reg_22_ ( .D(data_in_3[90]), .E(n1349), .CK(clk), .QN(n698) );
  EDFFXL R11_reg_21_ ( .D(data_in_3[89]), .E(n1349), .CK(clk), .QN(n699) );
  EDFFXL R11_reg_20_ ( .D(data_in_3[88]), .E(n1349), .CK(clk), .QN(n700) );
  EDFFXL R11_reg_19_ ( .D(data_in_3[87]), .E(n1349), .CK(clk), .QN(n701) );
  EDFFX1 R11_reg_18_ ( .D(data_in_3[86]), .E(n1349), .CK(clk), .QN(n702) );
  EDFFX1 R11_reg_17_ ( .D(data_in_3[85]), .E(n1349), .CK(clk), .QN(n703) );
  EDFFXL R11_reg_12_ ( .D(data_in_3[80]), .E(n1348), .CK(clk), .QN(n708) );
  EDFFXL R11_reg_10_ ( .D(data_in_3[78]), .E(n1348), .CK(clk), .QN(n710) );
  EDFFXL R11_reg_9_ ( .D(data_in_3[77]), .E(n1348), .CK(clk), .QN(n711) );
  EDFFXL R11_reg_8_ ( .D(data_in_3[76]), .E(n1348), .CK(clk), .QN(n712) );
  EDFFXL R11_reg_7_ ( .D(data_in_3[75]), .E(n1348), .CK(clk), .QN(n713) );
  EDFFXL R11_reg_6_ ( .D(data_in_3[74]), .E(n1348), .CK(clk), .QN(n714) );
  EDFFXL R11_reg_5_ ( .D(data_in_3[73]), .E(n1348), .CK(clk), .QN(n715) );
  EDFFXL R11_reg_4_ ( .D(data_in_3[72]), .E(n1348), .CK(clk), .QN(n716) );
  EDFFXL R11_reg_3_ ( .D(data_in_3[71]), .E(n1348), .CK(clk), .QN(n717) );
  EDFFXL R11_reg_2_ ( .D(data_in_3[70]), .E(n1348), .CK(clk), .QN(n718) );
  EDFFXL R11_reg_1_ ( .D(data_in_3[69]), .E(n1347), .CK(clk), .QN(n719) );
  EDFFX1 R11_reg_0_ ( .D(data_in_3[68]), .E(n1351), .CK(clk), .QN(n720) );
  EDFFXL R8_reg_27_ ( .D(data_in_3[95]), .E(n1364), .CK(clk), .QN(n761) );
  EDFFXL R8_reg_26_ ( .D(data_in_3[94]), .E(n1364), .CK(clk), .QN(n762) );
  EDFFXL R8_reg_25_ ( .D(data_in_3[93]), .E(n1363), .CK(clk), .QN(n763) );
  EDFFXL R8_reg_24_ ( .D(data_in_3[92]), .E(n1363), .CK(clk), .QN(n764) );
  EDFFXL R8_reg_23_ ( .D(data_in_3[91]), .E(n1363), .CK(clk), .QN(n765) );
  EDFFXL R8_reg_22_ ( .D(data_in_3[90]), .E(n1363), .CK(clk), .QN(n766) );
  EDFFXL R8_reg_21_ ( .D(data_in_3[89]), .E(n1363), .CK(clk), .QN(n767) );
  EDFFXL R8_reg_20_ ( .D(data_in_3[88]), .E(n1363), .CK(clk), .QN(n768) );
  EDFFXL R8_reg_19_ ( .D(data_in_3[87]), .E(n1363), .CK(clk), .QN(n769) );
  EDFFX1 R8_reg_18_ ( .D(data_in_3[86]), .E(n1363), .CK(clk), .QN(n770) );
  EDFFX1 R8_reg_17_ ( .D(data_in_3[85]), .E(n1363), .CK(clk), .QN(n771) );
  EDFFXL R8_reg_12_ ( .D(data_in_3[80]), .E(n1362), .CK(clk), .QN(n776) );
  EDFFXL R8_reg_10_ ( .D(data_in_3[78]), .E(n1362), .CK(clk), .QN(n778) );
  EDFFXL R8_reg_9_ ( .D(data_in_3[77]), .E(n1362), .CK(clk), .QN(n779) );
  EDFFXL R8_reg_8_ ( .D(data_in_3[76]), .E(n1362), .CK(clk), .QN(n780) );
  EDFFXL R8_reg_7_ ( .D(data_in_3[75]), .E(n1362), .CK(clk), .QN(n781) );
  EDFFXL R8_reg_6_ ( .D(data_in_3[74]), .E(n1362), .CK(clk), .QN(n782) );
  EDFFXL R8_reg_5_ ( .D(data_in_3[73]), .E(n1362), .CK(clk), .QN(n783) );
  EDFFXL R8_reg_4_ ( .D(data_in_3[72]), .E(n1362), .CK(clk), .QN(n784) );
  EDFFXL R8_reg_3_ ( .D(data_in_3[71]), .E(n1362), .CK(clk), .QN(n785) );
  EDFFXL R8_reg_2_ ( .D(data_in_3[70]), .E(n1362), .CK(clk), .QN(n786) );
  EDFFXL R8_reg_1_ ( .D(data_in_3[69]), .E(n1361), .CK(clk), .QN(n787) );
  EDFFX1 R8_reg_0_ ( .D(data_in_3[68]), .E(n1361), .CK(clk), .QN(n788) );
  EDFFXL R9_reg_27_ ( .D(data_in_3[95]), .E(n1377), .CK(clk), .QN(n829) );
  EDFFXL R9_reg_26_ ( .D(data_in_3[94]), .E(n1377), .CK(clk), .QN(n830) );
  EDFFXL R9_reg_25_ ( .D(data_in_3[93]), .E(n1376), .CK(clk), .QN(n831) );
  EDFFXL R9_reg_24_ ( .D(data_in_3[92]), .E(n1376), .CK(clk), .QN(n832) );
  EDFFXL R9_reg_23_ ( .D(data_in_3[91]), .E(n1376), .CK(clk), .QN(n833) );
  EDFFXL R9_reg_22_ ( .D(data_in_3[90]), .E(n1376), .CK(clk), .QN(n834) );
  EDFFXL R9_reg_21_ ( .D(data_in_3[89]), .E(n1376), .CK(clk), .QN(n835) );
  EDFFXL R9_reg_20_ ( .D(data_in_3[88]), .E(n1376), .CK(clk), .QN(n836) );
  EDFFXL R9_reg_19_ ( .D(data_in_3[87]), .E(n1376), .CK(clk), .QN(n837) );
  EDFFX1 R9_reg_18_ ( .D(data_in_3[86]), .E(n1376), .CK(clk), .QN(n838) );
  EDFFX1 R9_reg_17_ ( .D(data_in_3[85]), .E(n1376), .CK(clk), .QN(n839) );
  EDFFXL R9_reg_12_ ( .D(data_in_3[80]), .E(n1375), .CK(clk), .QN(n844) );
  EDFFXL R9_reg_10_ ( .D(data_in_3[78]), .E(n1375), .CK(clk), .QN(n846) );
  EDFFXL R9_reg_9_ ( .D(data_in_3[77]), .E(n1375), .CK(clk), .QN(n847) );
  EDFFXL R9_reg_8_ ( .D(data_in_3[76]), .E(n1375), .CK(clk), .QN(n848) );
  EDFFXL R9_reg_7_ ( .D(data_in_3[75]), .E(n1375), .CK(clk), .QN(n849) );
  EDFFXL R9_reg_6_ ( .D(data_in_3[74]), .E(n1375), .CK(clk), .QN(n850) );
  EDFFXL R9_reg_5_ ( .D(data_in_3[73]), .E(n1375), .CK(clk), .QN(n851) );
  EDFFXL R9_reg_4_ ( .D(data_in_3[72]), .E(n1375), .CK(clk), .QN(n852) );
  EDFFXL R9_reg_3_ ( .D(data_in_3[71]), .E(n1375), .CK(clk), .QN(n853) );
  EDFFXL R9_reg_2_ ( .D(data_in_3[70]), .E(n1375), .CK(clk), .QN(n854) );
  EDFFXL R9_reg_1_ ( .D(data_in_3[69]), .E(n1374), .CK(clk), .QN(n855) );
  EDFFX1 R9_reg_0_ ( .D(data_in_3[68]), .E(n1374), .CK(clk), .QN(n856) );
  EDFFXL R14_reg_29_ ( .D(data_in_3[131]), .E(n1391), .CK(clk), .Q(R14[29]) );
  EDFFXL R14_reg_27_ ( .D(data_in_3[129]), .E(n1394), .CK(clk), .Q(R14[27]) );
  EDFFXL R14_reg_26_ ( .D(data_in_3[128]), .E(n1394), .CK(clk), .Q(R14[26]) );
  EDFFXL R14_reg_25_ ( .D(data_in_3[127]), .E(n1389), .CK(clk), .Q(R14[25]) );
  EDFFXL R14_reg_24_ ( .D(data_in_3[126]), .E(n1392), .CK(clk), .Q(R14[24]) );
  EDFFXL R14_reg_23_ ( .D(data_in_3[125]), .E(n163), .CK(clk), .Q(R14[23]) );
  EDFFXL R14_reg_22_ ( .D(data_in_3[124]), .E(n1394), .CK(clk), .Q(R14[22]) );
  EDFFXL R14_reg_21_ ( .D(data_in_3[123]), .E(n1390), .CK(clk), .Q(R14[21]) );
  EDFFXL R14_reg_20_ ( .D(data_in_3[122]), .E(n163), .CK(clk), .Q(R14[20]) );
  EDFFXL R14_reg_19_ ( .D(data_in_3[121]), .E(n1394), .CK(clk), .Q(R14[19]) );
  EDFFXL R14_reg_18_ ( .D(data_in_3[120]), .E(n163), .CK(clk), .Q(R14[18]) );
  EDFFX1 R14_reg_17_ ( .D(data_in_3[119]), .E(n163), .CK(clk), .Q(R14[17]) );
  EDFFXL R14_reg_10_ ( .D(data_in_3[112]), .E(n1394), .CK(clk), .Q(R14[10]) );
  EDFFXL R14_reg_8_ ( .D(data_in_3[110]), .E(n163), .CK(clk), .Q(R14[8]) );
  EDFFXL R14_reg_7_ ( .D(data_in_3[109]), .E(n163), .CK(clk), .Q(R14[7]) );
  EDFFXL R14_reg_6_ ( .D(data_in_3[108]), .E(n1394), .CK(clk), .Q(R14[6]) );
  EDFFXL R14_reg_5_ ( .D(data_in_3[107]), .E(n163), .CK(clk), .Q(R14[5]) );
  EDFFXL R14_reg_4_ ( .D(data_in_3[106]), .E(n1394), .CK(clk), .Q(R14[4]) );
  EDFFXL R14_reg_3_ ( .D(data_in_3[105]), .E(n1390), .CK(clk), .Q(R14[3]) );
  EDFFXL R14_reg_2_ ( .D(data_in_3[104]), .E(n1390), .CK(clk), .Q(R14[2]) );
  EDFFX1 R14_reg_1_ ( .D(data_in_3[103]), .E(n1390), .CK(clk), .Q(R14[1]) );
  EDFFX1 R14_reg_0_ ( .D(data_in_3[102]), .E(n1390), .CK(clk), .Q(R14[0]) );
  EDFFXL R15_reg_29_ ( .D(data_in_3[131]), .E(n1352), .CK(clk), .Q(R15[29]) );
  EDFFXL R15_reg_27_ ( .D(data_in_3[129]), .E(n1351), .CK(clk), .Q(R15[27]) );
  EDFFXL R15_reg_26_ ( .D(data_in_3[128]), .E(n1356), .CK(clk), .Q(R15[26]) );
  EDFFXL R15_reg_25_ ( .D(data_in_3[127]), .E(n1351), .CK(clk), .Q(R15[25]) );
  EDFFXL R15_reg_24_ ( .D(data_in_3[126]), .E(n1356), .CK(clk), .Q(R15[24]) );
  EDFFXL R15_reg_23_ ( .D(data_in_3[125]), .E(n1347), .CK(clk), .Q(R15[23]) );
  EDFFXL R15_reg_22_ ( .D(data_in_3[124]), .E(n1347), .CK(clk), .Q(R15[22]) );
  EDFFXL R15_reg_21_ ( .D(data_in_3[123]), .E(n1347), .CK(clk), .Q(R15[21]) );
  EDFFXL R15_reg_20_ ( .D(data_in_3[122]), .E(n1347), .CK(clk), .Q(R15[20]) );
  EDFFXL R15_reg_19_ ( .D(data_in_3[121]), .E(n1347), .CK(clk), .Q(R15[19]) );
  EDFFXL R15_reg_18_ ( .D(data_in_3[120]), .E(n1347), .CK(clk), .Q(R15[18]) );
  EDFFX1 R15_reg_17_ ( .D(data_in_3[119]), .E(n1347), .CK(clk), .Q(R15[17]) );
  EDFFXL R15_reg_8_ ( .D(data_in_3[110]), .E(n1346), .CK(clk), .Q(R15[8]) );
  EDFFXL R15_reg_7_ ( .D(data_in_3[109]), .E(n1346), .CK(clk), .Q(R15[7]) );
  EDFFXL R15_reg_6_ ( .D(data_in_3[108]), .E(n1346), .CK(clk), .Q(R15[6]) );
  EDFFXL R15_reg_5_ ( .D(data_in_3[107]), .E(n1346), .CK(clk), .Q(R15[5]) );
  EDFFXL R15_reg_4_ ( .D(data_in_3[106]), .E(n1346), .CK(clk), .Q(R15[4]) );
  EDFFXL R15_reg_3_ ( .D(data_in_3[105]), .E(n1346), .CK(clk), .Q(R15[3]) );
  EDFFXL R15_reg_2_ ( .D(data_in_3[104]), .E(n1346), .CK(clk), .Q(R15[2]) );
  EDFFX1 R15_reg_1_ ( .D(data_in_3[103]), .E(n1346), .CK(clk), .Q(R15[1]) );
  EDFFX1 R15_reg_0_ ( .D(data_in_3[102]), .E(n1346), .CK(clk), .Q(R15[0]) );
  EDFFXL R12_reg_29_ ( .D(data_in_3[131]), .E(n1361), .CK(clk), .Q(R12[29]) );
  EDFFXL R12_reg_27_ ( .D(data_in_3[129]), .E(n1361), .CK(clk), .Q(R12[27]) );
  EDFFXL R12_reg_26_ ( .D(data_in_3[128]), .E(n1361), .CK(clk), .Q(R12[26]) );
  EDFFXL R12_reg_25_ ( .D(data_in_3[127]), .E(n1361), .CK(clk), .Q(R12[25]) );
  EDFFXL R12_reg_24_ ( .D(data_in_3[126]), .E(n1361), .CK(clk), .Q(R12[24]) );
  EDFFXL R12_reg_23_ ( .D(data_in_3[125]), .E(n1360), .CK(clk), .Q(R12[23]) );
  EDFFXL R12_reg_22_ ( .D(data_in_3[124]), .E(n1360), .CK(clk), .Q(R12[22]) );
  EDFFXL R12_reg_21_ ( .D(data_in_3[123]), .E(n1360), .CK(clk), .Q(R12[21]) );
  EDFFXL R12_reg_20_ ( .D(data_in_3[122]), .E(n1360), .CK(clk), .Q(R12[20]) );
  EDFFXL R12_reg_19_ ( .D(data_in_3[121]), .E(n1360), .CK(clk), .Q(R12[19]) );
  EDFFXL R12_reg_18_ ( .D(data_in_3[120]), .E(n1360), .CK(clk), .Q(R12[18]) );
  EDFFX1 R12_reg_17_ ( .D(data_in_3[119]), .E(n1360), .CK(clk), .Q(R12[17]) );
  EDFFXL R12_reg_10_ ( .D(data_in_3[112]), .E(n1359), .CK(clk), .Q(R12[10]) );
  EDFFXL R12_reg_8_ ( .D(data_in_3[110]), .E(n1359), .CK(clk), .Q(R12[8]) );
  EDFFXL R12_reg_7_ ( .D(data_in_3[109]), .E(n1359), .CK(clk), .Q(R12[7]) );
  EDFFXL R12_reg_6_ ( .D(data_in_3[108]), .E(n1359), .CK(clk), .Q(R12[6]) );
  EDFFXL R12_reg_5_ ( .D(data_in_3[107]), .E(n1359), .CK(clk), .Q(R12[5]) );
  EDFFXL R12_reg_4_ ( .D(data_in_3[106]), .E(n1359), .CK(clk), .Q(R12[4]) );
  EDFFXL R12_reg_3_ ( .D(data_in_3[105]), .E(n1359), .CK(clk), .Q(R12[3]) );
  EDFFXL R12_reg_2_ ( .D(data_in_3[104]), .E(n1359), .CK(clk), .Q(R12[2]) );
  EDFFX1 R12_reg_1_ ( .D(data_in_3[103]), .E(n1359), .CK(clk), .Q(R12[1]) );
  EDFFX1 R12_reg_0_ ( .D(data_in_3[102]), .E(n1359), .CK(clk), .Q(R12[0]) );
  EDFFXL R13_reg_29_ ( .D(data_in_3[131]), .E(n1374), .CK(clk), .Q(R13[29]) );
  EDFFXL R13_reg_27_ ( .D(data_in_3[129]), .E(n1374), .CK(clk), .Q(R13[27]) );
  EDFFXL R13_reg_26_ ( .D(data_in_3[128]), .E(n1374), .CK(clk), .Q(R13[26]) );
  EDFFXL R13_reg_25_ ( .D(data_in_3[127]), .E(n1374), .CK(clk), .Q(R13[25]) );
  EDFFXL R13_reg_24_ ( .D(data_in_3[126]), .E(n1374), .CK(clk), .Q(R13[24]) );
  EDFFXL R13_reg_23_ ( .D(data_in_3[125]), .E(n1373), .CK(clk), .Q(R13[23]) );
  EDFFXL R13_reg_22_ ( .D(data_in_3[124]), .E(n1373), .CK(clk), .Q(R13[22]) );
  EDFFXL R13_reg_21_ ( .D(data_in_3[123]), .E(n1373), .CK(clk), .Q(R13[21]) );
  EDFFXL R13_reg_20_ ( .D(data_in_3[122]), .E(n1373), .CK(clk), .Q(R13[20]) );
  EDFFXL R13_reg_19_ ( .D(data_in_3[121]), .E(n1373), .CK(clk), .Q(R13[19]) );
  EDFFXL R13_reg_18_ ( .D(data_in_3[120]), .E(n1373), .CK(clk), .Q(R13[18]) );
  EDFFX1 R13_reg_17_ ( .D(data_in_3[119]), .E(n1373), .CK(clk), .Q(R13[17]) );
  EDFFXL R13_reg_10_ ( .D(data_in_3[112]), .E(n1372), .CK(clk), .Q(R13[10]) );
  EDFFXL R13_reg_8_ ( .D(data_in_3[110]), .E(n1372), .CK(clk), .Q(R13[8]) );
  EDFFXL R13_reg_7_ ( .D(data_in_3[109]), .E(n1372), .CK(clk), .Q(R13[7]) );
  EDFFXL R13_reg_6_ ( .D(data_in_3[108]), .E(n1372), .CK(clk), .Q(R13[6]) );
  EDFFXL R13_reg_5_ ( .D(data_in_3[107]), .E(n1372), .CK(clk), .Q(R13[5]) );
  EDFFXL R13_reg_4_ ( .D(data_in_3[106]), .E(n1372), .CK(clk), .Q(R13[4]) );
  EDFFXL R13_reg_3_ ( .D(data_in_3[105]), .E(n1372), .CK(clk), .Q(R13[3]) );
  EDFFXL R13_reg_2_ ( .D(data_in_3[104]), .E(n1372), .CK(clk), .Q(R13[2]) );
  EDFFX1 R13_reg_1_ ( .D(data_in_3[103]), .E(n1372), .CK(clk), .Q(R13[1]) );
  EDFFX1 R13_reg_0_ ( .D(data_in_3[102]), .E(n1372), .CK(clk), .Q(R13[0]) );
  EDFFXL R2_reg_26_ ( .D(data_in_3[26]), .E(n1393), .CK(clk), .Q(R2[26]) );
  EDFFXL R2_reg_25_ ( .D(data_in_3[25]), .E(n1393), .CK(clk), .Q(R2[25]) );
  EDFFXL R2_reg_24_ ( .D(data_in_3[24]), .E(n1393), .CK(clk), .Q(R2[24]) );
  EDFFXL R2_reg_23_ ( .D(data_in_3[23]), .E(n1393), .CK(clk), .Q(R2[23]) );
  EDFFXL R2_reg_22_ ( .D(data_in_3[22]), .E(n1393), .CK(clk), .Q(R2[22]) );
  EDFFXL R2_reg_21_ ( .D(data_in_3[21]), .E(n1393), .CK(clk), .Q(R2[21]) );
  EDFFXL R2_reg_20_ ( .D(data_in_3[20]), .E(n1393), .CK(clk), .Q(R2[20]) );
  EDFFXL R2_reg_19_ ( .D(data_in_3[19]), .E(n1393), .CK(clk), .Q(R2[19]) );
  EDFFX1 R2_reg_17_ ( .D(data_in_3[17]), .E(n1392), .CK(clk), .Q(R2[17]) );
  EDFFXL R2_reg_12_ ( .D(data_in_3[12]), .E(n1392), .CK(clk), .Q(R2[12]) );
  EDFFXL R2_reg_8_ ( .D(data_in_3[8]), .E(n1392), .CK(clk), .Q(R2[8]) );
  EDFFXL R2_reg_7_ ( .D(data_in_3[7]), .E(n1392), .CK(clk), .Q(R2[7]) );
  EDFFXL R2_reg_6_ ( .D(data_in_3[6]), .E(n1392), .CK(clk), .Q(R2[6]) );
  EDFFXL R2_reg_5_ ( .D(data_in_3[5]), .E(n1391), .CK(clk), .Q(R2[5]) );
  EDFFXL R2_reg_4_ ( .D(data_in_3[4]), .E(n1391), .CK(clk), .Q(R2[4]) );
  EDFFXL R2_reg_3_ ( .D(data_in_3[3]), .E(n1391), .CK(clk), .Q(R2[3]) );
  EDFFXL R2_reg_2_ ( .D(data_in_3[2]), .E(n1391), .CK(clk), .Q(R2[2]) );
  EDFFX1 R2_reg_1_ ( .D(data_in_3[1]), .E(n1391), .CK(clk), .Q(R2[1]) );
  EDFFX1 R2_reg_0_ ( .D(data_in_3[0]), .E(n1391), .CK(clk), .Q(R2[0]) );
  EDFFXL R3_reg_26_ ( .D(data_in_3[26]), .E(n1352), .CK(clk), .Q(R3[26]) );
  EDFFXL R3_reg_25_ ( .D(data_in_3[25]), .E(n1352), .CK(clk), .Q(R3[25]) );
  EDFFXL R3_reg_24_ ( .D(data_in_3[24]), .E(n1352), .CK(clk), .Q(R3[24]) );
  EDFFXL R3_reg_23_ ( .D(data_in_3[23]), .E(n1352), .CK(clk), .Q(R3[23]) );
  EDFFXL R3_reg_22_ ( .D(data_in_3[22]), .E(n1352), .CK(clk), .Q(R3[22]) );
  EDFFXL R3_reg_21_ ( .D(data_in_3[21]), .E(n1352), .CK(clk), .Q(R3[21]) );
  EDFFXL R3_reg_20_ ( .D(data_in_3[20]), .E(n1352), .CK(clk), .Q(R3[20]) );
  EDFFXL R3_reg_19_ ( .D(data_in_3[19]), .E(n1352), .CK(clk), .Q(R3[19]) );
  EDFFX1 R3_reg_17_ ( .D(data_in_3[17]), .E(n1352), .CK(clk), .Q(R3[17]) );
  EDFFXL R3_reg_12_ ( .D(data_in_3[12]), .E(n1351), .CK(clk), .Q(R3[12]) );
  EDFFXL R3_reg_8_ ( .D(data_in_3[8]), .E(n1351), .CK(clk), .Q(R3[8]) );
  EDFFXL R3_reg_7_ ( .D(data_in_3[7]), .E(n1351), .CK(clk), .Q(R3[7]) );
  EDFFXL R3_reg_6_ ( .D(data_in_3[6]), .E(n1351), .CK(clk), .Q(R3[6]) );
  EDFFXL R3_reg_5_ ( .D(data_in_3[5]), .E(n1351), .CK(clk), .Q(R3[5]) );
  EDFFXL R3_reg_4_ ( .D(data_in_3[4]), .E(n1351), .CK(clk), .Q(R3[4]) );
  EDFFXL R3_reg_3_ ( .D(data_in_3[3]), .E(n1350), .CK(clk), .Q(R3[3]) );
  EDFFXL R3_reg_2_ ( .D(data_in_3[2]), .E(n1350), .CK(clk), .Q(R3[2]) );
  EDFFX1 R3_reg_1_ ( .D(data_in_3[1]), .E(n1350), .CK(clk), .Q(R3[1]) );
  EDFFX1 R3_reg_0_ ( .D(data_in_3[0]), .E(n1350), .CK(clk), .Q(R3[0]) );
  EDFFXL R0_reg_26_ ( .D(data_in_3[26]), .E(n1369), .CK(clk), .Q(R0[26]) );
  EDFFXL R0_reg_25_ ( .D(data_in_3[25]), .E(n1369), .CK(clk), .Q(R0[25]) );
  EDFFXL R0_reg_24_ ( .D(data_in_3[24]), .E(n1369), .CK(clk), .Q(R0[24]) );
  EDFFXL R0_reg_23_ ( .D(data_in_3[23]), .E(n1369), .CK(clk), .Q(R0[23]) );
  EDFFXL R0_reg_22_ ( .D(data_in_3[22]), .E(n1369), .CK(clk), .Q(R0[22]) );
  EDFFXL R0_reg_21_ ( .D(data_in_3[21]), .E(n1369), .CK(clk), .Q(R0[21]) );
  EDFFXL R0_reg_20_ ( .D(data_in_3[20]), .E(n1369), .CK(clk), .Q(R0[20]) );
  EDFFXL R0_reg_19_ ( .D(data_in_3[19]), .E(n1369), .CK(clk), .Q(R0[19]) );
  EDFFX1 R0_reg_17_ ( .D(data_in_3[17]), .E(n1368), .CK(clk), .Q(R0[17]) );
  EDFFXL R0_reg_12_ ( .D(data_in_3[12]), .E(n1368), .CK(clk), .Q(R0[12]) );
  EDFFXL R0_reg_8_ ( .D(data_in_3[8]), .E(n1368), .CK(clk), .Q(R0[8]) );
  EDFFXL R0_reg_7_ ( .D(data_in_3[7]), .E(n1368), .CK(clk), .Q(R0[7]) );
  EDFFXL R0_reg_6_ ( .D(data_in_3[6]), .E(n1368), .CK(clk), .Q(R0[6]) );
  EDFFXL R0_reg_5_ ( .D(data_in_3[5]), .E(n1367), .CK(clk), .Q(R0[5]) );
  EDFFXL R0_reg_4_ ( .D(data_in_3[4]), .E(n1367), .CK(clk), .Q(R0[4]) );
  EDFFXL R0_reg_3_ ( .D(data_in_3[3]), .E(n1367), .CK(clk), .Q(R0[3]) );
  EDFFXL R0_reg_2_ ( .D(data_in_3[2]), .E(n1367), .CK(clk), .Q(R0[2]) );
  EDFFX1 R0_reg_1_ ( .D(data_in_3[1]), .E(n1367), .CK(clk), .Q(R0[1]) );
  EDFFX1 R0_reg_0_ ( .D(data_in_3[0]), .E(n1367), .CK(clk), .Q(R0[0]) );
  EDFFXL R1_reg_26_ ( .D(data_in_3[26]), .E(n1382), .CK(clk), .Q(R1[26]) );
  EDFFXL R1_reg_25_ ( .D(data_in_3[25]), .E(n1382), .CK(clk), .Q(R1[25]) );
  EDFFXL R1_reg_24_ ( .D(data_in_3[24]), .E(n1382), .CK(clk), .Q(R1[24]) );
  EDFFXL R1_reg_23_ ( .D(data_in_3[23]), .E(n1382), .CK(clk), .Q(R1[23]) );
  EDFFXL R1_reg_22_ ( .D(data_in_3[22]), .E(n1382), .CK(clk), .Q(R1[22]) );
  EDFFXL R1_reg_21_ ( .D(data_in_3[21]), .E(n1382), .CK(clk), .Q(R1[21]) );
  EDFFXL R1_reg_20_ ( .D(data_in_3[20]), .E(n1382), .CK(clk), .Q(R1[20]) );
  EDFFXL R1_reg_19_ ( .D(data_in_3[19]), .E(n1382), .CK(clk), .Q(R1[19]) );
  EDFFX1 R1_reg_17_ ( .D(data_in_3[17]), .E(n1381), .CK(clk), .Q(R1[17]) );
  EDFFXL R1_reg_12_ ( .D(data_in_3[12]), .E(n1381), .CK(clk), .Q(R1[12]) );
  EDFFXL R1_reg_8_ ( .D(data_in_3[8]), .E(n1381), .CK(clk), .Q(R1[8]) );
  EDFFXL R1_reg_7_ ( .D(data_in_3[7]), .E(n1381), .CK(clk), .Q(R1[7]) );
  EDFFXL R1_reg_6_ ( .D(data_in_3[6]), .E(n1381), .CK(clk), .Q(R1[6]) );
  EDFFXL R1_reg_5_ ( .D(data_in_3[5]), .E(n1380), .CK(clk), .Q(R1[5]) );
  EDFFXL R1_reg_4_ ( .D(data_in_3[4]), .E(n1380), .CK(clk), .Q(R1[4]) );
  EDFFXL R1_reg_3_ ( .D(data_in_3[3]), .E(n1380), .CK(clk), .Q(R1[3]) );
  EDFFXL R1_reg_2_ ( .D(data_in_3[2]), .E(n1380), .CK(clk), .Q(R1[2]) );
  EDFFX1 R1_reg_1_ ( .D(data_in_3[1]), .E(n1380), .CK(clk), .Q(R1[1]) );
  EDFFX1 R1_reg_0_ ( .D(data_in_3[0]), .E(n1380), .CK(clk), .Q(R1[0]) );
  JKFFRXL counter_1_reg_0_ ( .J(1'b1), .K(1'b1), .CK(clk), .RN(rst_n), .Q(
        counter_1[0]), .QN(n584) );
  DFFRHQX1 counter_1_reg_1_ ( .D(N26), .CK(clk), .RN(rst_n), .Q(counter_1[1])
         );
  JKFFRXL counter_2_reg_0_ ( .J(1'b1), .K(1'b1), .CK(clk), .RN(rst_n), .Q(
        counter_2[0]), .QN(n861) );
  DFFRHQX1 counter_2_reg_1_ ( .D(N50), .CK(clk), .RN(rst_n), .Q(counter_2[1])
         );
  DFFRHQX1 counter_2_reg_2_ ( .D(n1403), .CK(clk), .RN(rst_n), .Q(counter_2[2]) );
  DFFRHQX1 counter_2_reg_3_ ( .D(N52), .CK(clk), .RN(rst_n), .Q(counter_2[3])
         );
  EDFFX1 data_out_3_reg_33_ ( .D(N152), .E(n1400), .CK(clk), .Q(data_out_3[33]) );
  EDFFX1 data_out_3_reg_32_ ( .D(N151), .E(n1400), .CK(clk), .Q(data_out_3[32]) );
  EDFFX1 data_out_3_reg_31_ ( .D(N150), .E(n1400), .CK(clk), .Q(data_out_3[31]) );
  EDFFX1 data_out_3_reg_30_ ( .D(N149), .E(n1400), .CK(clk), .Q(data_out_3[30]) );
  EDFFX1 data_out_3_reg_29_ ( .D(N148), .E(n1400), .CK(clk), .Q(data_out_3[29]) );
  EDFFX1 data_out_3_reg_28_ ( .D(N147), .E(n1400), .CK(clk), .Q(data_out_3[28]) );
  EDFFX1 data_out_3_reg_27_ ( .D(N146), .E(n1400), .CK(clk), .Q(data_out_3[27]) );
  EDFFX1 data_out_3_reg_26_ ( .D(N145), .E(n1400), .CK(clk), .Q(data_out_3[26]) );
  EDFFX1 data_out_3_reg_25_ ( .D(N144), .E(n1400), .CK(clk), .Q(data_out_3[25]) );
  EDFFX1 data_out_3_reg_24_ ( .D(N143), .E(n1400), .CK(clk), .Q(data_out_3[24]) );
  EDFFX1 data_out_3_reg_23_ ( .D(N142), .E(n1400), .CK(clk), .Q(data_out_3[23]) );
  EDFFX1 data_out_3_reg_22_ ( .D(N141), .E(n1400), .CK(clk), .Q(data_out_3[22]) );
  EDFFX1 data_out_3_reg_21_ ( .D(N140), .E(n1400), .CK(clk), .Q(data_out_3[21]) );
  EDFFX1 data_out_3_reg_20_ ( .D(N139), .E(n1400), .CK(clk), .Q(data_out_3[20]) );
  EDFFX1 data_out_3_reg_19_ ( .D(N138), .E(n1400), .CK(clk), .Q(data_out_3[19]) );
  EDFFX1 data_out_3_reg_18_ ( .D(N137), .E(n1400), .CK(clk), .Q(data_out_3[18]) );
  EDFFX1 data_out_3_reg_17_ ( .D(N136), .E(n1400), .CK(clk), .Q(data_out_3[17]) );
  EDFFX1 data_out_3_reg_16_ ( .D(N135), .E(n1400), .CK(clk), .Q(data_out_3[16]) );
  EDFFX1 data_out_3_reg_15_ ( .D(N134), .E(n1400), .CK(clk), .Q(data_out_3[15]) );
  EDFFX1 data_out_3_reg_14_ ( .D(N133), .E(n1400), .CK(clk), .Q(data_out_3[14]) );
  EDFFX1 data_out_3_reg_13_ ( .D(N132), .E(n1400), .CK(clk), .Q(data_out_3[13]) );
  EDFFX1 data_out_3_reg_12_ ( .D(N131), .E(n1400), .CK(clk), .Q(data_out_3[12]) );
  EDFFX1 data_out_3_reg_11_ ( .D(N130), .E(n1400), .CK(clk), .Q(data_out_3[11]) );
  EDFFX1 data_out_3_reg_10_ ( .D(N129), .E(n1400), .CK(clk), .Q(data_out_3[10]) );
  EDFFX1 data_out_3_reg_9_ ( .D(N128), .E(n1400), .CK(clk), .Q(data_out_3[9])
         );
  EDFFX1 data_out_3_reg_8_ ( .D(N127), .E(n1400), .CK(clk), .Q(data_out_3[8])
         );
  EDFFX1 data_out_3_reg_7_ ( .D(N126), .E(n1400), .CK(clk), .Q(data_out_3[7])
         );
  EDFFX1 data_out_3_reg_6_ ( .D(N125), .E(n1400), .CK(clk), .Q(data_out_3[6])
         );
  EDFFX1 data_out_3_reg_5_ ( .D(N124), .E(n1400), .CK(clk), .Q(data_out_3[5])
         );
  EDFFX1 data_out_3_reg_4_ ( .D(N123), .E(n1400), .CK(clk), .Q(data_out_3[4])
         );
  EDFFX1 data_out_3_reg_3_ ( .D(N122), .E(n1400), .CK(clk), .Q(data_out_3[3])
         );
  EDFFX1 data_out_3_reg_2_ ( .D(N121), .E(n1400), .CK(clk), .Q(data_out_3[2])
         );
  EDFFX1 data_out_3_reg_1_ ( .D(N120), .E(n1400), .CK(clk), .Q(data_out_3[1])
         );
  EDFFX1 data_out_3_reg_0_ ( .D(N119), .E(n1400), .CK(clk), .Q(data_out_3[0])
         );
  EDFFXL R2_reg_18_ ( .D(data_in_3[18]), .E(n1393), .CK(clk), .Q(R2[18]) );
  EDFFXL R3_reg_18_ ( .D(data_in_3[18]), .E(n1352), .CK(clk), .Q(R3[18]) );
  EDFFXL R0_reg_18_ ( .D(data_in_3[18]), .E(n1369), .CK(clk), .Q(R0[18]) );
  EDFFXL R1_reg_18_ ( .D(data_in_3[18]), .E(n1382), .CK(clk), .Q(R1[18]) );
  EDFFX1 R5_reg_18_ ( .D(data_in_3[52]), .E(n1379), .CK(clk), .QN(n804) );
  EDFFX1 R5_reg_17_ ( .D(data_in_3[51]), .E(n1379), .CK(clk), .QN(n805) );
  EDFFX1 R5_reg_1_ ( .D(data_in_3[35]), .E(n1377), .CK(clk), .QN(n821) );
  EDFFX1 R5_reg_0_ ( .D(data_in_3[34]), .E(n1377), .CK(clk), .QN(n822) );
  EDFFXL R7_reg_7_ ( .D(data_in_3[41]), .E(n1354), .CK(clk), .QN(n611) );
  EDFFXL R4_reg_7_ ( .D(data_in_3[41]), .E(n1365), .CK(clk), .QN(n747) );
  EDFFXL R6_reg_7_ ( .D(data_in_3[41]), .E(n1385), .CK(clk), .QN(n679) );
  EDFFXL R7_reg_30_ ( .D(data_in_3[64]), .E(n1356), .CK(clk), .QN(n588) );
  EDFFXL R6_reg_30_ ( .D(data_in_3[64]), .E(n1387), .CK(clk), .QN(n656) );
  EDFFXL R4_reg_30_ ( .D(data_in_3[64]), .E(n1367), .CK(clk), .QN(n724) );
  EDFFXL R7_reg_12_ ( .D(data_in_3[46]), .E(n1354), .CK(clk), .QN(n606) );
  EDFFXL R6_reg_12_ ( .D(data_in_3[46]), .E(n1386), .CK(clk), .QN(n674) );
  EDFFXL R4_reg_12_ ( .D(data_in_3[46]), .E(n1365), .CK(clk), .QN(n742) );
  EDFFXL R7_reg_22_ ( .D(data_in_3[56]), .E(n1355), .CK(clk), .QN(n596) );
  EDFFXL R6_reg_22_ ( .D(data_in_3[56]), .E(n1386), .CK(clk), .QN(n664) );
  EDFFXL R4_reg_22_ ( .D(data_in_3[56]), .E(n1366), .CK(clk), .QN(n732) );
  EDFFXL R7_reg_10_ ( .D(data_in_3[44]), .E(n1354), .CK(clk), .QN(n608) );
  EDFFXL R6_reg_10_ ( .D(data_in_3[44]), .E(n1385), .CK(clk), .QN(n676) );
  EDFFXL R4_reg_10_ ( .D(data_in_3[44]), .E(n1365), .CK(clk), .QN(n744) );
  EDFFXL R15_reg_10_ ( .D(data_in_3[112]), .E(n1346), .CK(clk), .Q(R15[10]) );
  DFFXL R1_reg_29_ ( .D(n1247), .CK(clk), .Q(n157) );
  DFFXL R0_reg_29_ ( .D(n1246), .CK(clk), .Q(n156) );
  DFFXL R2_reg_33_ ( .D(n1270), .CK(clk), .Q(n151) );
  DFFXL R1_reg_33_ ( .D(n1269), .CK(clk), .Q(n150) );
  DFFXL R0_reg_33_ ( .D(n1268), .CK(clk), .Q(n149) );
  DFFXL R3_reg_33_ ( .D(n1271), .CK(clk), .Q(n147) );
  DFFXL R1_reg_16_ ( .D(n1286), .CK(clk), .Q(n143) );
  DFFXL R2_reg_16_ ( .D(n1287), .CK(clk), .Q(n139) );
  DFFXL R12_reg_14_ ( .D(n1229), .CK(clk), .Q(n131) );
  EDFFX1 R1_reg_9_ ( .D(data_in_3[9]), .E(n1381), .CK(clk), .Q(R1[9]) );
  EDFFX1 R0_reg_9_ ( .D(data_in_3[9]), .E(n1368), .CK(clk), .Q(R0[9]) );
  EDFFX1 R3_reg_9_ ( .D(data_in_3[9]), .E(n1351), .CK(clk), .Q(R3[9]) );
  EDFFX1 R2_reg_9_ ( .D(data_in_3[9]), .E(n1392), .CK(clk), .Q(R2[9]) );
  DFFXL R15_reg_14_ ( .D(n1232), .CK(clk), .Q(n125) );
  DFFXL R13_reg_14_ ( .D(n1230), .CK(clk), .Q(n123) );
  DFFXL R15_reg_28_ ( .D(n1278), .CK(clk), .Q(n116) );
  DFFXL R14_reg_28_ ( .D(n1277), .CK(clk), .Q(n114) );
  DFFXL R13_reg_28_ ( .D(n1276), .CK(clk), .Q(n111) );
  DFFXL R12_reg_28_ ( .D(n1275), .CK(clk), .Q(n110) );
  DFFXL R13_reg_31_ ( .D(n1285), .CK(clk), .Q(n104) );
  DFFXL R12_reg_31_ ( .D(n1284), .CK(clk), .Q(n103) );
  DFFXL R2_reg_31_ ( .D(n1259), .CK(clk), .Q(n97) );
  DFFXL R1_reg_31_ ( .D(n1258), .CK(clk), .Q(n96) );
  DFFXL R0_reg_31_ ( .D(n1257), .CK(clk), .Q(n95) );
  DFFXL R15_reg_33_ ( .D(n1300), .CK(clk), .Q(n93) );
  DFFXL R14_reg_33_ ( .D(n1299), .CK(clk), .Q(n91) );
  EDFFXL R7_reg_27_ ( .D(data_in_3[61]), .E(n1355), .CK(clk), .QN(n591) );
  EDFFXL R6_reg_27_ ( .D(data_in_3[61]), .E(n1387), .CK(clk), .QN(n659) );
  EDFFXL R4_reg_27_ ( .D(data_in_3[61]), .E(n1366), .CK(clk), .QN(n727) );
  DFFXL R15_reg_13_ ( .D(n1245), .CK(clk), .Q(n78) );
  DFFXL R13_reg_13_ ( .D(n1243), .CK(clk), .Q(n77) );
  DFFXL R12_reg_13_ ( .D(n1242), .CK(clk), .Q(n76) );
  DFFXL R14_reg_16_ ( .D(n1237), .CK(clk), .Q(n75) );
  EDFFXL R11_reg_13_ ( .D(data_in_3[81]), .E(n1352), .CK(clk), .QN(n707) );
  EDFFXL R13_reg_16_ ( .D(data_in_3[118]), .E(n1376), .CK(clk), .Q(n136) );
  EDFFXL R10_reg_13_ ( .D(data_in_3[81]), .E(n6), .CK(clk), .QN(n639) );
  EDFFXL R3_reg_10_ ( .D(data_in_3[10]), .E(n1356), .CK(clk), .Q(n155) );
  EDFFXL R12_reg_16_ ( .D(data_in_3[118]), .E(n1369), .CK(clk), .Q(n133) );
  EDFFXL R0_reg_16_ ( .D(data_in_3[16]), .E(n1365), .CK(clk), .Q(n142) );
  EDFFXL R9_reg_13_ ( .D(data_in_3[81]), .E(n1375), .CK(clk), .QN(n843) );
  EDFFXL R15_reg_16_ ( .D(data_in_3[118]), .E(n1351), .CK(clk), .Q(n88) );
  EDFFXL R10_reg_16_ ( .D(data_in_3[84]), .E(n6), .CK(clk), .QN(n636) );
  EDFFXL R5_reg_31_ ( .D(data_in_3[65]), .E(n1378), .CK(clk), .QN(n791) );
  EDFFXL R1_reg_10_ ( .D(data_in_3[10]), .E(n1374), .CK(clk), .Q(n146) );
  EDFFXL R9_reg_16_ ( .D(data_in_3[84]), .E(n1376), .CK(clk), .QN(n840) );
  EDFFXL R4_reg_31_ ( .D(data_in_3[65]), .E(n1359), .CK(clk), .QN(n723) );
  EDFFXL R8_reg_13_ ( .D(data_in_3[81]), .E(n1366), .CK(clk), .QN(n775) );
  EDFFXL R8_reg_16_ ( .D(data_in_3[84]), .E(n1365), .CK(clk), .QN(n772) );
  EDFFXL R6_reg_31_ ( .D(data_in_3[65]), .E(n6), .CK(clk), .QN(n655) );
  EDFFXL R5_reg_33_ ( .D(data_in_3[67]), .E(n1374), .CK(clk), .QN(n789) );
  EDFFXL R15_reg_15_ ( .D(data_in_3[117]), .E(n1352), .CK(clk), .Q(R15[15]) );
  EDFFXL R0_reg_10_ ( .D(data_in_3[10]), .E(n1366), .CK(clk), .Q(n145) );
  EDFFXL R3_reg_16_ ( .D(data_in_3[16]), .E(n1347), .CK(clk), .Q(n141) );
  EDFFXL R3_reg_15_ ( .D(data_in_3[15]), .E(n1347), .CK(clk), .Q(R3[15]) );
  DFFXL R13_reg_15_ ( .D(n1273), .CK(clk), .Q(n51) );
  EDFFXL R15_reg_31_ ( .D(data_in_3[133]), .E(n1352), .CK(clk), .Q(n109) );
  EDFFXL R14_reg_31_ ( .D(data_in_3[133]), .E(n6), .CK(clk), .Q(n108) );
  EDFFXL R11_reg_32_ ( .D(data_in_3[100]), .E(n1347), .CK(clk), .QN(n688) );
  DFFXL R13_reg_32_ ( .D(n1239), .CK(clk), .Q(n43) );
  DFFXL R12_reg_32_ ( .D(n1238), .CK(clk), .Q(n42) );
  DFFXL R15_reg_32_ ( .D(n1241), .CK(clk), .Q(n40) );
  EDFFXL R1_reg_13_ ( .D(data_in_3[13]), .E(n1379), .CK(clk), .Q(R1[13]) );
  EDFFXL R3_reg_31_ ( .D(data_in_3[31]), .E(n1347), .CK(clk), .Q(R3[31]) );
  EDFFXL R3_reg_13_ ( .D(data_in_3[13]), .E(n1351), .CK(clk), .Q(R3[13]) );
  EDFFXL R10_reg_31_ ( .D(data_in_3[99]), .E(n6), .CK(clk), .QN(n621) );
  EDFFXL R12_reg_33_ ( .D(data_in_3[135]), .E(n1366), .CK(clk), .Q(n89) );
  EDFFXL R4_reg_33_ ( .D(data_in_3[67]), .E(n1359), .CK(clk), .QN(n721) );
  EDFFXL R13_reg_33_ ( .D(data_in_3[135]), .E(n1373), .CK(clk), .Q(n90) );
  EDFFXL R9_reg_31_ ( .D(data_in_3[99]), .E(n1375), .CK(clk), .QN(n825) );
  EDFFXL R7_reg_31_ ( .D(data_in_3[65]), .E(n1352), .CK(clk), .QN(n587) );
  EDFFXL R0_reg_15_ ( .D(data_in_3[15]), .E(n1368), .CK(clk), .Q(n49) );
  EDFFXL R2_reg_15_ ( .D(data_in_3[15]), .E(n1392), .CK(clk), .Q(n50) );
  EDFFXL R14_reg_12_ ( .D(data_in_3[114]), .E(n163), .CK(clk), .Q(R14[12]) );
  EDFFXL R7_reg_23_ ( .D(data_in_3[57]), .E(n1355), .CK(clk), .QN(n595) );
  EDFFXL R14_reg_30_ ( .D(data_in_3[132]), .E(n1391), .CK(clk), .Q(R14[30]) );
  EDFFXL R2_reg_29_ ( .D(data_in_3[29]), .E(n1393), .CK(clk), .Q(n158) );
  JKFFRX2 p_s_flag_out_reg ( .J(n1406), .K(1'b0), .CK(clk), .RN(rst_n), .Q(
        n1400) );
  MX2X2 U3 ( .A(data_in_3[135]), .B(n93), .S0(n227), .Y(n1300) );
  MX2X2 U6 ( .A(data_in_3[16]), .B(n143), .S0(n1), .Y(n1286) );
  CLKINVX20 U7 ( .A(n1381), .Y(n1) );
  MX2X2 U8 ( .A(data_in_3[16]), .B(n139), .S0(n1396), .Y(n1287) );
  BUFX1 U9 ( .A(data_in_3[43]), .Y(n53) );
  NAND2X2 U10 ( .A(data_in_3[134]), .B(n2), .Y(n3) );
  NAND2X4 U11 ( .A(R14[32]), .B(n1396), .Y(n4) );
  NAND2X2 U12 ( .A(n3), .B(n4), .Y(n1240) );
  INVX20 U13 ( .A(n1396), .Y(n2) );
  INVX4 U14 ( .A(n6), .Y(n1396) );
  INVX1 U15 ( .A(n1347), .Y(n5) );
  MX2X4 U16 ( .A(data_in_3[130]), .B(n116), .S0(n5), .Y(n1278) );
  INVX1 U17 ( .A(n226), .Y(n161) );
  INVX1 U18 ( .A(n1364), .Y(n21) );
  NOR3X2 U19 ( .A(counter_1[1]), .B(p_s_flag_in), .C(counter_1[0]), .Y(n6) );
  AND2X2 U20 ( .A(n1162), .B(n872), .Y(n7) );
  NAND2X1 U21 ( .A(n1162), .B(n869), .Y(n8) );
  NAND2X1 U22 ( .A(n1162), .B(n871), .Y(n9) );
  AND2X2 U23 ( .A(n872), .B(n1157), .Y(n10) );
  AND2X2 U24 ( .A(n872), .B(n1163), .Y(n11) );
  AND2X2 U25 ( .A(n1159), .B(n1163), .Y(n12) );
  AND2X2 U26 ( .A(n1159), .B(n1158), .Y(n13) );
  AND2X2 U27 ( .A(n1159), .B(n1157), .Y(n14) );
  NAND2X1 U28 ( .A(n1158), .B(n871), .Y(n15) );
  NAND2X1 U29 ( .A(n1158), .B(n869), .Y(n16) );
  NAND2X1 U30 ( .A(n871), .B(n1163), .Y(n17) );
  NAND2X1 U31 ( .A(n1157), .B(n871), .Y(n18) );
  INVX1 U32 ( .A(n1353), .Y(n137) );
  INVX1 U33 ( .A(n1399), .Y(n163) );
  INVX1 U34 ( .A(n1356), .Y(n19) );
  MX2X1 U35 ( .A(data_in_3[11]), .B(R3[11]), .S0(n19), .Y(n1304) );
  MX2X1 U36 ( .A(data_in_3[11]), .B(R1[11]), .S0(n1384), .Y(n1302) );
  MX2X1 U37 ( .A(data_in_3[11]), .B(R2[11]), .S0(n1397), .Y(n1303) );
  MX2X2 U38 ( .A(data_in_3[67]), .B(n547), .S0(n19), .Y(n1172) );
  MX2X2 U39 ( .A(data_in_3[67]), .B(n411), .S0(n20), .Y(n1171) );
  CLKINVX20 U40 ( .A(n1387), .Y(n20) );
  AOI22XL U41 ( .A0(n1333), .A1(R3[15]), .B0(n886), .B1(R14[15]), .Y(n1037) );
  AOI22XL U42 ( .A0(n1314), .A1(R1[15]), .B0(n1316), .B1(R12[15]), .Y(n1039)
         );
  MX2X4 U43 ( .A(data_in_3[117]), .B(R14[15]), .S0(n1395), .Y(n1274) );
  MX2X4 U44 ( .A(data_in_3[117]), .B(R12[15]), .S0(n1371), .Y(n1272) );
  MX2X1 U45 ( .A(n373), .B(data_in_3[97]), .S0(n1350), .Y(n1168) );
  MX2X1 U46 ( .A(data_in_3[96]), .B(n236), .S0(n21), .Y(n1209) );
  INVXL U47 ( .A(p_s_flag_in), .Y(n1406) );
  MX2X2 U49 ( .A(n239), .B(data_in_3[99]), .S0(n1364), .Y(n1169) );
  MX2X2 U50 ( .A(n375), .B(data_in_3[99]), .S0(n1350), .Y(n1170) );
  MX2X1 U51 ( .A(data_in_3[11]), .B(R0[11]), .S0(n1371), .Y(n1301) );
  MX2X2 U52 ( .A(n91), .B(data_in_3[135]), .S0(n1391), .Y(n1299) );
  MX2X1 U53 ( .A(n42), .B(data_in_3[134]), .S0(n1361), .Y(n1238) );
  MX2X1 U54 ( .A(n43), .B(data_in_3[134]), .S0(n1374), .Y(n1239) );
  MX2X1 U55 ( .A(n40), .B(data_in_3[134]), .S0(n1351), .Y(n1241) );
  MX2X2 U56 ( .A(data_in_3[33]), .B(n147), .S0(n1357), .Y(n1271) );
  MX2X1 U57 ( .A(n359), .B(data_in_3[83]), .S0(n1349), .Y(n1184) );
  MX2X2 U58 ( .A(n121), .B(data_in_3[49]), .S0(n1378), .Y(n1174) );
  MX2X2 U59 ( .A(n529), .B(data_in_3[49]), .S0(n1354), .Y(n1176) );
  MX2X2 U60 ( .A(n393), .B(data_in_3[49]), .S0(n1386), .Y(n1175) );
  MX2X2 U61 ( .A(n257), .B(data_in_3[49]), .S0(n1365), .Y(n1173) );
  MX2X2 U62 ( .A(data_in_3[15]), .B(R1[15]), .S0(n1384), .Y(n1279) );
  MX2X1 U63 ( .A(n1306), .B(data_in_3[98]), .S0(n34), .Y(n1203) );
  CLKINVX20 U64 ( .A(n1358), .Y(n34) );
  MX2X2 U65 ( .A(R2[13]), .B(data_in_3[13]), .S0(n1392), .Y(n1261) );
  MX2X2 U66 ( .A(R0[13]), .B(data_in_3[13]), .S0(n1368), .Y(n1260) );
  AOI22XL U67 ( .A0(n1332), .A1(R3[31]), .B0(n886), .B1(n108), .Y(n909) );
  MX2X2 U68 ( .A(n103), .B(data_in_3[133]), .S0(n1361), .Y(n1284) );
  MX2X2 U69 ( .A(n104), .B(data_in_3[133]), .S0(n1374), .Y(n1285) );
  MX2X2 U70 ( .A(data_in_3[14]), .B(R2[14]), .S0(n1396), .Y(n1293) );
  MX2X2 U71 ( .A(data_in_3[84]), .B(n360), .S0(n1358), .Y(n1204) );
  MX2X4 U72 ( .A(data_in_3[10]), .B(R2[10]), .S0(n1399), .Y(n1266) );
  MX2X1 U73 ( .A(n51), .B(data_in_3[117]), .S0(n1373), .Y(n1273) );
  MX2X2 U74 ( .A(data_in_3[118]), .B(n75), .S0(n1395), .Y(n1237) );
  MX2X2 U75 ( .A(n151), .B(data_in_3[33]), .S0(n1394), .Y(n1270) );
  MX2X2 U76 ( .A(n149), .B(data_in_3[33]), .S0(n1370), .Y(n1268) );
  MX2X2 U77 ( .A(n150), .B(data_in_3[33]), .S0(n1383), .Y(n1269) );
  MX2X2 U78 ( .A(R12[9]), .B(data_in_3[111]), .S0(n1359), .Y(n1295) );
  MX2X2 U79 ( .A(R13[9]), .B(data_in_3[111]), .S0(n1372), .Y(n1296) );
  MX2X2 U80 ( .A(R15[9]), .B(data_in_3[111]), .S0(n1346), .Y(n1298) );
  MX2X2 U81 ( .A(R14[9]), .B(data_in_3[111]), .S0(n163), .Y(n1297) );
  MX2X2 U82 ( .A(n1312), .B(data_in_3[100]), .S0(n161), .Y(n1193) );
  MX2X2 U83 ( .A(n1313), .B(data_in_3[100]), .S0(n162), .Y(n1194) );
  MX2X2 U84 ( .A(n1311), .B(data_in_3[100]), .S0(n163), .Y(n1195) );
  MX2X4 U85 ( .A(data_in_3[115]), .B(R14[13]), .S0(n1397), .Y(n1244) );
  MX2X1 U86 ( .A(n76), .B(data_in_3[115]), .S0(n1360), .Y(n1242) );
  MX2X1 U87 ( .A(n77), .B(data_in_3[115]), .S0(n1373), .Y(n1243) );
  MX2X1 U88 ( .A(n78), .B(data_in_3[115]), .S0(n1347), .Y(n1245) );
  AOI22XL U89 ( .A0(n1333), .A1(n141), .B0(n886), .B1(n75), .Y(n1029) );
  MX2X1 U90 ( .A(n525), .B(data_in_3[45]), .S0(n1354), .Y(n1199) );
  MX2X1 U91 ( .A(n389), .B(data_in_3[45]), .S0(n1385), .Y(n1198) );
  MX2X1 U92 ( .A(n117), .B(data_in_3[45]), .S0(n1378), .Y(n1197) );
  MX2X1 U93 ( .A(n253), .B(data_in_3[45]), .S0(n1365), .Y(n1196) );
  MX2X1 U94 ( .A(n123), .B(data_in_3[116]), .S0(n1373), .Y(n1230) );
  MX2X1 U95 ( .A(n125), .B(data_in_3[116]), .S0(n1347), .Y(n1232) );
  MX2X2 U96 ( .A(data_in_3[30]), .B(R3[30]), .S0(n137), .Y(n1265) );
  MX2X2 U97 ( .A(data_in_3[116]), .B(R14[14]), .S0(n1398), .Y(n1231) );
  MX2X1 U98 ( .A(n131), .B(data_in_3[116]), .S0(n1360), .Y(n1229) );
  MX2X2 U99 ( .A(R3[14]), .B(data_in_3[14]), .S0(n1351), .Y(n1294) );
  MX2X2 U100 ( .A(R0[14]), .B(data_in_3[14]), .S0(n1368), .Y(n1291) );
  MX2X2 U101 ( .A(R1[14]), .B(data_in_3[14]), .S0(n1381), .Y(n1292) );
  MX2X2 U102 ( .A(R0[30]), .B(data_in_3[30]), .S0(n1370), .Y(n1262) );
  MX2X2 U103 ( .A(R1[30]), .B(data_in_3[30]), .S0(n1383), .Y(n1263) );
  MX2X2 U104 ( .A(R2[30]), .B(data_in_3[30]), .S0(n1394), .Y(n1264) );
  MX2X2 U105 ( .A(data_in_3[32]), .B(R3[32]), .S0(n137), .Y(n1256) );
  MX2X2 U106 ( .A(data_in_3[29]), .B(R3[29]), .S0(n19), .Y(n1248) );
  MX2X2 U107 ( .A(R0[32]), .B(data_in_3[32]), .S0(n1370), .Y(n1253) );
  MX2X2 U108 ( .A(R1[32]), .B(data_in_3[32]), .S0(n1383), .Y(n1254) );
  MX2X2 U109 ( .A(R2[32]), .B(data_in_3[32]), .S0(n1394), .Y(n1255) );
  CLKINVX20 U110 ( .A(n1384), .Y(n162) );
  MX2X2 U111 ( .A(n445), .B(data_in_3[101]), .S0(n1390), .Y(n893) );
  MX2X2 U112 ( .A(n241), .B(data_in_3[101]), .S0(n1364), .Y(n891) );
  MX2X2 U113 ( .A(n105), .B(data_in_3[101]), .S0(n1377), .Y(n892) );
  MX2X1 U114 ( .A(data_in_3[96]), .B(n372), .S0(n137), .Y(n1212) );
  MX2X2 U115 ( .A(n377), .B(data_in_3[101]), .S0(n1350), .Y(n895) );
  MX2X1 U116 ( .A(n156), .B(data_in_3[29]), .S0(n1369), .Y(n1246) );
  MX2X1 U117 ( .A(n157), .B(data_in_3[29]), .S0(n1382), .Y(n1247) );
  MX2X2 U118 ( .A(R14[11]), .B(data_in_3[113]), .S0(n163), .Y(n1235) );
  MX2X2 U119 ( .A(R12[11]), .B(data_in_3[113]), .S0(n1359), .Y(n1233) );
  MX2X2 U120 ( .A(R13[11]), .B(data_in_3[113]), .S0(n1372), .Y(n1234) );
  MX2X2 U121 ( .A(R15[11]), .B(data_in_3[113]), .S0(n1346), .Y(n1236) );
  MX2X2 U122 ( .A(R15[30]), .B(data_in_3[132]), .S0(n1356), .Y(n1267) );
  MX2X2 U123 ( .A(n110), .B(data_in_3[130]), .S0(n1361), .Y(n1275) );
  MX2X2 U124 ( .A(n111), .B(data_in_3[130]), .S0(n1374), .Y(n1276) );
  MX2X2 U125 ( .A(n114), .B(data_in_3[130]), .S0(n1391), .Y(n1277) );
  INVX1 U126 ( .A(n867), .Y(n1314) );
  INVX1 U127 ( .A(n16), .Y(n1333) );
  INVX1 U128 ( .A(n18), .Y(n1339) );
  INVX1 U129 ( .A(n9), .Y(n1321) );
  INVX1 U130 ( .A(n8), .Y(n1316) );
  INVX1 U131 ( .A(n15), .Y(n1341) );
  INVX1 U132 ( .A(n9), .Y(n1322) );
  INVX1 U133 ( .A(n17), .Y(n1324) );
  INVX1 U134 ( .A(n13), .Y(n1345) );
  INVX1 U135 ( .A(n12), .Y(n1329) );
  INVX1 U136 ( .A(n11), .Y(n1320) );
  INVX1 U137 ( .A(n14), .Y(n1342) );
  INVX1 U138 ( .A(n10), .Y(n1335) );
  INVX1 U139 ( .A(n1327), .Y(n1325) );
  INVX1 U140 ( .A(n7), .Y(n1317) );
  INVX1 U141 ( .A(n14), .Y(n1343) );
  INVX1 U142 ( .A(n1327), .Y(n1326) );
  INVX1 U143 ( .A(n7), .Y(n1318) );
  INVX1 U144 ( .A(n225), .Y(n1379) );
  INVX1 U145 ( .A(n226), .Y(n1366) );
  INVX1 U146 ( .A(n1399), .Y(n1385) );
  INVX1 U147 ( .A(n225), .Y(n1372) );
  INVX1 U148 ( .A(n225), .Y(n1375) );
  INVX1 U149 ( .A(n226), .Y(n1359) );
  INVX1 U150 ( .A(n21), .Y(n1362) );
  INVX1 U151 ( .A(n1357), .Y(n1348) );
  INVX1 U152 ( .A(n1396), .Y(n1388) );
  INVX1 U153 ( .A(n227), .Y(n1352) );
  INVX1 U154 ( .A(n1358), .Y(n1355) );
  INVX1 U155 ( .A(n225), .Y(n1376) );
  INVX1 U156 ( .A(n225), .Y(n1382) );
  INVX1 U157 ( .A(n1371), .Y(n1363) );
  INVX1 U158 ( .A(n226), .Y(n1369) );
  INVX1 U159 ( .A(n1358), .Y(n1349) );
  INVX1 U160 ( .A(n1398), .Y(n1389) );
  INVX1 U161 ( .A(n1395), .Y(n1393) );
  INVX1 U162 ( .A(n225), .Y(n1378) );
  INVX1 U163 ( .A(n226), .Y(n1365) );
  INVX1 U164 ( .A(n1399), .Y(n1386) );
  INVX1 U165 ( .A(n225), .Y(n1373) );
  INVX1 U166 ( .A(n1384), .Y(n1380) );
  INVX1 U167 ( .A(n21), .Y(n1360) );
  INVX1 U168 ( .A(n1371), .Y(n1367) );
  INVX1 U169 ( .A(n227), .Y(n1347) );
  INVX1 U170 ( .A(n1398), .Y(n1387) );
  INVX1 U171 ( .A(n227), .Y(n1351) );
  INVX1 U172 ( .A(n1357), .Y(n1354) );
  INVX1 U173 ( .A(n1396), .Y(n1391) );
  INVX1 U174 ( .A(n225), .Y(n1377) );
  INVX1 U175 ( .A(n1384), .Y(n1381) );
  INVX1 U176 ( .A(n226), .Y(n1364) );
  INVX1 U177 ( .A(n1371), .Y(n1368) );
  INVX1 U178 ( .A(n1398), .Y(n1390) );
  INVX1 U179 ( .A(n1358), .Y(n1350) );
  INVX1 U180 ( .A(n1357), .Y(n1353) );
  INVX1 U181 ( .A(n1396), .Y(n1392) );
  INVX1 U182 ( .A(n1357), .Y(n1346) );
  INVX1 U183 ( .A(n225), .Y(n1374) );
  INVX1 U184 ( .A(n21), .Y(n1361) );
  INVX1 U185 ( .A(n1337), .Y(n1336) );
  INVX1 U186 ( .A(n227), .Y(n1356) );
  INVX1 U187 ( .A(n1371), .Y(n1370) );
  INVX1 U188 ( .A(n1384), .Y(n1383) );
  INVX1 U189 ( .A(n1395), .Y(n1394) );
  INVX1 U190 ( .A(n15), .Y(n1340) );
  INVX1 U191 ( .A(n16), .Y(n1332) );
  INVX1 U192 ( .A(n18), .Y(n1338) );
  INVX1 U193 ( .A(n1331), .Y(n1330) );
  INVX1 U194 ( .A(n886), .Y(n1331) );
  INVX1 U195 ( .A(n8), .Y(n1315) );
  INVX1 U196 ( .A(n17), .Y(n1323) );
  INVX1 U197 ( .A(n867), .Y(n1402) );
  INVX1 U198 ( .A(n13), .Y(n1344) );
  INVX1 U199 ( .A(n12), .Y(n1328) );
  INVX1 U200 ( .A(n11), .Y(n1319) );
  INVX1 U201 ( .A(n10), .Y(n1334) );
  INVX1 U202 ( .A(n6), .Y(n1395) );
  INVX1 U203 ( .A(n1377), .Y(n1384) );
  INVX1 U204 ( .A(n161), .Y(n1371) );
  INVX1 U205 ( .A(n6), .Y(n1399) );
  INVX1 U206 ( .A(n6), .Y(n1398) );
  INVX1 U207 ( .A(n6), .Y(n1397) );
  INVX1 U208 ( .A(n1356), .Y(n1358) );
  INVX1 U209 ( .A(n1356), .Y(n1357) );
  INVX1 U210 ( .A(n882), .Y(n1337) );
  INVX1 U211 ( .A(n888), .Y(n1327) );
  NOR2X1 U212 ( .A(n1405), .B(n1404), .Y(n869) );
  NAND2X1 U213 ( .A(n1163), .B(n869), .Y(n867) );
  NAND2X1 U214 ( .A(n872), .B(n1158), .Y(n882) );
  NAND2X1 U215 ( .A(n1162), .B(n1159), .Y(n888) );
  NOR2X1 U216 ( .A(n861), .B(counter_2[3]), .Y(n1163) );
  OAI221XL U217 ( .A0(n856), .A1(n1345), .B0(n822), .B1(n1343), .C0(n1156), 
        .Y(n1155) );
  AOI22X1 U218 ( .A0(n1340), .A1(R2[0]), .B0(n1338), .B1(R13[0]), .Y(n1156) );
  OAI221XL U219 ( .A0(n855), .A1(n1344), .B0(n821), .B1(n1343), .C0(n1148), 
        .Y(n1147) );
  AOI22X1 U220 ( .A0(n1340), .A1(R2[1]), .B0(n1338), .B1(R13[1]), .Y(n1148) );
  OAI221XL U221 ( .A0(n854), .A1(n1345), .B0(n820), .B1(n1343), .C0(n1140), 
        .Y(n1139) );
  AOI22X1 U222 ( .A0(n1340), .A1(R2[2]), .B0(n1338), .B1(R13[2]), .Y(n1140) );
  OAI221XL U223 ( .A0(n853), .A1(n1344), .B0(n819), .B1(n1343), .C0(n1132), 
        .Y(n1131) );
  AOI22X1 U224 ( .A0(n1340), .A1(R2[3]), .B0(n1338), .B1(R13[3]), .Y(n1132) );
  OAI221XL U225 ( .A0(n852), .A1(n1345), .B0(n818), .B1(n1343), .C0(n1124), 
        .Y(n1123) );
  AOI22X1 U226 ( .A0(n1340), .A1(R2[4]), .B0(n1338), .B1(R13[4]), .Y(n1124) );
  OAI221XL U227 ( .A0(n851), .A1(n1344), .B0(n817), .B1(n1343), .C0(n1116), 
        .Y(n1115) );
  AOI22X1 U228 ( .A0(n1340), .A1(R2[5]), .B0(n1338), .B1(R13[5]), .Y(n1116) );
  OAI221XL U229 ( .A0(n850), .A1(n1345), .B0(n816), .B1(n1343), .C0(n1108), 
        .Y(n1107) );
  AOI22X1 U230 ( .A0(n1340), .A1(R2[6]), .B0(n1338), .B1(R13[6]), .Y(n1108) );
  OAI221XL U231 ( .A0(n849), .A1(n1344), .B0(n815), .B1(n1343), .C0(n1100), 
        .Y(n1099) );
  AOI22X1 U232 ( .A0(n1340), .A1(R2[7]), .B0(n1338), .B1(R13[7]), .Y(n1100) );
  OAI221XL U233 ( .A0(n848), .A1(n1345), .B0(n814), .B1(n1343), .C0(n1092), 
        .Y(n1091) );
  AOI22X1 U234 ( .A0(n1340), .A1(R2[8]), .B0(n1338), .B1(R13[8]), .Y(n1092) );
  OAI221XL U235 ( .A0(n839), .A1(n1345), .B0(n805), .B1(n1342), .C0(n1020), 
        .Y(n1019) );
  AOI22X1 U236 ( .A0(n1341), .A1(R2[17]), .B0(n1339), .B1(R13[17]), .Y(n1020)
         );
  OAI221XL U237 ( .A0(n838), .A1(n1345), .B0(n804), .B1(n1342), .C0(n1012), 
        .Y(n1011) );
  AOI22X1 U238 ( .A0(n1341), .A1(R2[18]), .B0(n1339), .B1(R13[18]), .Y(n1012)
         );
  OAI221XL U239 ( .A0(n837), .A1(n1345), .B0(n803), .B1(n1342), .C0(n1004), 
        .Y(n1003) );
  AOI22X1 U240 ( .A0(n1340), .A1(R2[19]), .B0(n1339), .B1(R13[19]), .Y(n1004)
         );
  OAI221XL U241 ( .A0(n836), .A1(n1345), .B0(n802), .B1(n1342), .C0(n996), .Y(
        n995) );
  AOI22X1 U242 ( .A0(n1341), .A1(R2[20]), .B0(n1339), .B1(R13[20]), .Y(n996)
         );
  OAI221XL U243 ( .A0(n835), .A1(n1344), .B0(n801), .B1(n1342), .C0(n988), .Y(
        n987) );
  AOI22X1 U244 ( .A0(n1340), .A1(R2[21]), .B0(n1339), .B1(R13[21]), .Y(n988)
         );
  OAI221XL U245 ( .A0(n834), .A1(n1344), .B0(n800), .B1(n1343), .C0(n980), .Y(
        n979) );
  AOI22X1 U246 ( .A0(n1341), .A1(R2[22]), .B0(n1339), .B1(R13[22]), .Y(n980)
         );
  OAI221XL U247 ( .A0(n833), .A1(n1344), .B0(n799), .B1(n1343), .C0(n972), .Y(
        n971) );
  AOI22X1 U248 ( .A0(n1340), .A1(R2[23]), .B0(n1339), .B1(R13[23]), .Y(n972)
         );
  OAI221XL U249 ( .A0(n832), .A1(n1344), .B0(n798), .B1(n1342), .C0(n964), .Y(
        n963) );
  AOI22X1 U250 ( .A0(n1341), .A1(R2[24]), .B0(n1339), .B1(R13[24]), .Y(n964)
         );
  OAI221XL U251 ( .A0(n831), .A1(n1344), .B0(n797), .B1(n1343), .C0(n956), .Y(
        n955) );
  AOI22X1 U252 ( .A0(n1341), .A1(R2[25]), .B0(n1338), .B1(R13[25]), .Y(n956)
         );
  OAI221XL U253 ( .A0(n830), .A1(n1344), .B0(n796), .B1(n1342), .C0(n948), .Y(
        n947) );
  AOI22X1 U254 ( .A0(n1341), .A1(R2[26]), .B0(n1339), .B1(R13[26]), .Y(n948)
         );
  OAI221XL U255 ( .A0(n710), .A1(n1329), .B0(n608), .B1(n1325), .C0(n1078), 
        .Y(n1073) );
  NOR2X1 U256 ( .A(counter_2[3]), .B(counter_2[0]), .Y(n1162) );
  NOR2X1 U257 ( .A(n1404), .B(counter_2[2]), .Y(n871) );
  INVX1 U258 ( .A(counter_2[1]), .Y(n1404) );
  AOI22X1 U259 ( .A0(n1340), .A1(R2[10]), .B0(n1338), .B1(R13[10]), .Y(n1076)
         );
  AOI22X1 U260 ( .A0(n1332), .A1(n155), .B0(n1330), .B1(R14[10]), .Y(n1077) );
  AOI22X1 U261 ( .A0(n1314), .A1(n146), .B0(n1315), .B1(R12[10]), .Y(n1079) );
  AOI22X1 U262 ( .A0(n1332), .A1(R3[11]), .B0(n1330), .B1(R14[11]), .Y(n1069)
         );
  AOI22X1 U263 ( .A0(n1323), .A1(R0[11]), .B0(n1322), .B1(R15[11]), .Y(n1070)
         );
  AOI22X1 U264 ( .A0(n1314), .A1(R1[11]), .B0(n1315), .B1(R12[11]), .Y(n1071)
         );
  AOI22X1 U265 ( .A0(n1333), .A1(R3[13]), .B0(n886), .B1(R14[13]), .Y(n1053)
         );
  AOI22X1 U266 ( .A0(n1324), .A1(R0[13]), .B0(n1321), .B1(n78), .Y(n1054) );
  AOI22X1 U267 ( .A0(n1314), .A1(R1[13]), .B0(n1316), .B1(n76), .Y(n1055) );
  AOI22X1 U268 ( .A0(n1333), .A1(R3[14]), .B0(n886), .B1(R14[14]), .Y(n1045)
         );
  AOI22X1 U269 ( .A0(n1324), .A1(R0[14]), .B0(n1321), .B1(n125), .Y(n1046) );
  AOI22X1 U270 ( .A0(n1314), .A1(R1[14]), .B0(n1316), .B1(n131), .Y(n1047) );
  AOI22X1 U271 ( .A0(n1324), .A1(n49), .B0(n1321), .B1(R15[15]), .Y(n1038) );
  AOI22X1 U272 ( .A0(n1324), .A1(n142), .B0(n1321), .B1(n88), .Y(n1030) );
  AOI22X1 U273 ( .A0(n1314), .A1(n143), .B0(n1316), .B1(n133), .Y(n1031) );
  AOI22X1 U274 ( .A0(n1332), .A1(R3[27]), .B0(n886), .B1(R14[27]), .Y(n941) );
  AOI22X1 U275 ( .A0(n1324), .A1(R0[27]), .B0(n1322), .B1(R15[27]), .Y(n942)
         );
  AOI22X1 U276 ( .A0(n1402), .A1(R1[27]), .B0(n1315), .B1(R12[27]), .Y(n943)
         );
  AOI22X1 U277 ( .A0(n1333), .A1(R3[28]), .B0(n886), .B1(n114), .Y(n933) );
  AOI22X1 U278 ( .A0(n1323), .A1(R0[28]), .B0(n1322), .B1(n116), .Y(n934) );
  AOI22X1 U279 ( .A0(n1402), .A1(R1[28]), .B0(n1315), .B1(n110), .Y(n935) );
  AOI22X1 U280 ( .A0(n1332), .A1(R3[29]), .B0(n886), .B1(R14[29]), .Y(n925) );
  AOI22X1 U281 ( .A0(n1324), .A1(n156), .B0(n1322), .B1(R15[29]), .Y(n926) );
  AOI22X1 U282 ( .A0(n1402), .A1(n157), .B0(n1316), .B1(R12[29]), .Y(n927) );
  AOI22X1 U283 ( .A0(n1333), .A1(R3[30]), .B0(n886), .B1(R14[30]), .Y(n917) );
  AOI22X1 U284 ( .A0(n1323), .A1(R0[30]), .B0(n1322), .B1(R15[30]), .Y(n918)
         );
  AOI22X1 U285 ( .A0(n1402), .A1(R1[30]), .B0(n1315), .B1(R12[30]), .Y(n919)
         );
  AOI22X1 U286 ( .A0(n1324), .A1(n95), .B0(n1322), .B1(n109), .Y(n910) );
  AOI22X1 U287 ( .A0(n1402), .A1(n96), .B0(n1316), .B1(n103), .Y(n911) );
  AOI22X1 U288 ( .A0(n1333), .A1(R3[32]), .B0(n1330), .B1(R14[32]), .Y(n901)
         );
  AOI22X1 U289 ( .A0(n1323), .A1(R0[32]), .B0(n1322), .B1(n40), .Y(n902) );
  AOI22X1 U290 ( .A0(n1402), .A1(R1[32]), .B0(n1315), .B1(n42), .Y(n903) );
  OAI221XL U291 ( .A0(n845), .A1(n1345), .B0(n811), .B1(n1342), .C0(n1068), 
        .Y(n1067) );
  AOI22X1 U292 ( .A0(n1340), .A1(R2[11]), .B0(n1338), .B1(R13[11]), .Y(n1068)
         );
  OAI221XL U293 ( .A0(n843), .A1(n1345), .B0(n809), .B1(n1342), .C0(n1052), 
        .Y(n1051) );
  AOI22X1 U294 ( .A0(n1341), .A1(R2[13]), .B0(n1339), .B1(n77), .Y(n1052) );
  OAI221XL U295 ( .A0(n842), .A1(n1345), .B0(n808), .B1(n1342), .C0(n1044), 
        .Y(n1043) );
  AOI22X1 U296 ( .A0(n1340), .A1(R2[14]), .B0(n1339), .B1(n123), .Y(n1044) );
  OAI221XL U297 ( .A0(n841), .A1(n1345), .B0(n807), .B1(n1342), .C0(n1036), 
        .Y(n1035) );
  AOI22X1 U298 ( .A0(n1341), .A1(n50), .B0(n1339), .B1(n51), .Y(n1036) );
  OAI221XL U299 ( .A0(n840), .A1(n1345), .B0(n806), .B1(n1342), .C0(n1028), 
        .Y(n1027) );
  AOI22X1 U300 ( .A0(n1340), .A1(n139), .B0(n1339), .B1(n136), .Y(n1028) );
  OAI221XL U301 ( .A0(n829), .A1(n1344), .B0(n795), .B1(n1343), .C0(n940), .Y(
        n939) );
  AOI22X1 U302 ( .A0(n1341), .A1(R2[27]), .B0(n1338), .B1(R13[27]), .Y(n940)
         );
  OAI221XL U303 ( .A0(n828), .A1(n1344), .B0(n794), .B1(n1342), .C0(n932), .Y(
        n931) );
  AOI22X1 U304 ( .A0(n1341), .A1(R2[28]), .B0(n1339), .B1(n111), .Y(n932) );
  OAI221XL U305 ( .A0(n827), .A1(n1344), .B0(n793), .B1(n1343), .C0(n924), .Y(
        n923) );
  AOI22X1 U306 ( .A0(n1341), .A1(n158), .B0(n1338), .B1(R13[29]), .Y(n924) );
  OAI221XL U307 ( .A0(n826), .A1(n1344), .B0(n792), .B1(n1342), .C0(n916), .Y(
        n915) );
  AOI22X1 U308 ( .A0(n1341), .A1(R2[30]), .B0(n1339), .B1(R13[30]), .Y(n916)
         );
  OAI221XL U309 ( .A0(n825), .A1(n1344), .B0(n791), .B1(n1343), .C0(n908), .Y(
        n907) );
  AOI22X1 U310 ( .A0(n1341), .A1(n97), .B0(n1338), .B1(n104), .Y(n908) );
  OAI221XL U311 ( .A0(n824), .A1(n1344), .B0(n790), .B1(n1342), .C0(n900), .Y(
        n899) );
  AOI22X1 U312 ( .A0(n1341), .A1(R2[32]), .B0(n1339), .B1(n43), .Y(n900) );
  AOI22X1 U313 ( .A0(n1332), .A1(R3[9]), .B0(n1330), .B1(R14[9]), .Y(n1085) );
  AOI22X1 U314 ( .A0(n1323), .A1(R0[9]), .B0(n1322), .B1(R15[9]), .Y(n1086) );
  AOI22X1 U315 ( .A0(n1314), .A1(R1[9]), .B0(n1315), .B1(R12[9]), .Y(n1087) );
  AOI22X1 U316 ( .A0(n1333), .A1(R3[12]), .B0(n886), .B1(R14[12]), .Y(n1061)
         );
  AOI22X1 U317 ( .A0(n1324), .A1(R0[12]), .B0(n1321), .B1(R15[12]), .Y(n1062)
         );
  AOI22X1 U318 ( .A0(n1314), .A1(R1[12]), .B0(n1316), .B1(R12[12]), .Y(n1063)
         );
  OAI221XL U319 ( .A0(n847), .A1(n1345), .B0(n813), .B1(n1343), .C0(n1084), 
        .Y(n1083) );
  AOI22X1 U320 ( .A0(n1340), .A1(R2[9]), .B0(n1338), .B1(R13[9]), .Y(n1084) );
  OAI221XL U322 ( .A0(n844), .A1(n1345), .B0(n810), .B1(n1342), .C0(n1060), 
        .Y(n1059) );
  AOI22X1 U323 ( .A0(n1341), .A1(R2[12]), .B0(n1339), .B1(R13[12]), .Y(n1060)
         );
  INVX1 U325 ( .A(counter_2[2]), .Y(n1405) );
  AOI22X1 U327 ( .A0(n1332), .A1(R3[0]), .B0(n1330), .B1(R14[0]), .Y(n1160) );
  AOI22X1 U328 ( .A0(n1323), .A1(R0[0]), .B0(n1321), .B1(R15[0]), .Y(n1161) );
  AOI22X1 U329 ( .A0(n1402), .A1(R1[0]), .B0(n1315), .B1(R12[0]), .Y(n1164) );
  AOI22X1 U330 ( .A0(n1332), .A1(R3[1]), .B0(n1330), .B1(R14[1]), .Y(n1149) );
  AOI22X1 U331 ( .A0(n1323), .A1(R0[1]), .B0(n1322), .B1(R15[1]), .Y(n1150) );
  AOI22X1 U332 ( .A0(n1402), .A1(R1[1]), .B0(n1315), .B1(R12[1]), .Y(n1151) );
  AOI22X1 U333 ( .A0(n1332), .A1(R3[2]), .B0(n1330), .B1(R14[2]), .Y(n1141) );
  AOI22X1 U334 ( .A0(n1323), .A1(R0[2]), .B0(n1321), .B1(R15[2]), .Y(n1142) );
  AOI22X1 U335 ( .A0(n1314), .A1(R1[2]), .B0(n1315), .B1(R12[2]), .Y(n1143) );
  AOI22X1 U336 ( .A0(n1332), .A1(R3[3]), .B0(n1330), .B1(R14[3]), .Y(n1133) );
  AOI22X1 U337 ( .A0(n1323), .A1(R0[3]), .B0(n1322), .B1(R15[3]), .Y(n1134) );
  AOI22X1 U338 ( .A0(n1402), .A1(R1[3]), .B0(n1315), .B1(R12[3]), .Y(n1135) );
  AOI22X1 U339 ( .A0(n1332), .A1(R3[4]), .B0(n1330), .B1(R14[4]), .Y(n1125) );
  AOI22X1 U340 ( .A0(n1323), .A1(R0[4]), .B0(n1321), .B1(R15[4]), .Y(n1126) );
  AOI22X1 U341 ( .A0(n1314), .A1(R1[4]), .B0(n1315), .B1(R12[4]), .Y(n1127) );
  AOI22X1 U342 ( .A0(n1332), .A1(R3[5]), .B0(n1330), .B1(R14[5]), .Y(n1117) );
  AOI22X1 U343 ( .A0(n1323), .A1(R0[5]), .B0(n1322), .B1(R15[5]), .Y(n1118) );
  AOI22X1 U344 ( .A0(n1402), .A1(R1[5]), .B0(n1315), .B1(R12[5]), .Y(n1119) );
  AOI22X1 U345 ( .A0(n1332), .A1(R3[6]), .B0(n1330), .B1(R14[6]), .Y(n1109) );
  AOI22X1 U346 ( .A0(n1323), .A1(R0[6]), .B0(n1321), .B1(R15[6]), .Y(n1110) );
  AOI22X1 U347 ( .A0(n1314), .A1(R1[6]), .B0(n1315), .B1(R12[6]), .Y(n1111) );
  AOI22X1 U348 ( .A0(n1332), .A1(R3[7]), .B0(n1330), .B1(R14[7]), .Y(n1101) );
  AOI22X1 U349 ( .A0(n1323), .A1(R0[7]), .B0(n1322), .B1(R15[7]), .Y(n1102) );
  AOI22X1 U350 ( .A0(n1402), .A1(R1[7]), .B0(n1315), .B1(R12[7]), .Y(n1103) );
  AOI22X1 U351 ( .A0(n1332), .A1(R3[8]), .B0(n1330), .B1(R14[8]), .Y(n1093) );
  AOI22X1 U352 ( .A0(n1323), .A1(R0[8]), .B0(n1321), .B1(R15[8]), .Y(n1094) );
  AOI22X1 U353 ( .A0(n1314), .A1(R1[8]), .B0(n1315), .B1(R12[8]), .Y(n1095) );
  AOI22X1 U354 ( .A0(n1333), .A1(R3[17]), .B0(n886), .B1(R14[17]), .Y(n1021)
         );
  AOI22X1 U355 ( .A0(n1324), .A1(R0[17]), .B0(n1321), .B1(R15[17]), .Y(n1022)
         );
  AOI22X1 U356 ( .A0(n1314), .A1(R1[17]), .B0(n1316), .B1(R12[17]), .Y(n1023)
         );
  AOI22X1 U357 ( .A0(n1333), .A1(R3[18]), .B0(n886), .B1(R14[18]), .Y(n1013)
         );
  AOI22X1 U358 ( .A0(n1324), .A1(R0[18]), .B0(n1321), .B1(R15[18]), .Y(n1014)
         );
  AOI22X1 U359 ( .A0(n1314), .A1(R1[18]), .B0(n1316), .B1(R12[18]), .Y(n1015)
         );
  AOI22X1 U360 ( .A0(n1333), .A1(R3[19]), .B0(n886), .B1(R14[19]), .Y(n1005)
         );
  AOI22X1 U361 ( .A0(n1324), .A1(R0[19]), .B0(n1321), .B1(R15[19]), .Y(n1006)
         );
  AOI22X1 U362 ( .A0(n1314), .A1(R1[19]), .B0(n1316), .B1(R12[19]), .Y(n1007)
         );
  AOI22X1 U363 ( .A0(n1333), .A1(R3[20]), .B0(n886), .B1(R14[20]), .Y(n997) );
  AOI22X1 U364 ( .A0(n1324), .A1(R0[20]), .B0(n1321), .B1(R15[20]), .Y(n998)
         );
  AOI22X1 U365 ( .A0(n1314), .A1(R1[20]), .B0(n1316), .B1(R12[20]), .Y(n999)
         );
  AOI22X1 U366 ( .A0(n1333), .A1(R3[21]), .B0(n886), .B1(R14[21]), .Y(n989) );
  AOI22X1 U367 ( .A0(n1324), .A1(R0[21]), .B0(n1321), .B1(R15[21]), .Y(n990)
         );
  AOI22X1 U368 ( .A0(n1314), .A1(R1[21]), .B0(n1316), .B1(R12[21]), .Y(n991)
         );
  AOI22X1 U369 ( .A0(n1333), .A1(R3[22]), .B0(n886), .B1(R14[22]), .Y(n981) );
  AOI22X1 U370 ( .A0(n1324), .A1(R0[22]), .B0(n1321), .B1(R15[22]), .Y(n982)
         );
  AOI22X1 U371 ( .A0(n1402), .A1(R1[22]), .B0(n1316), .B1(R12[22]), .Y(n983)
         );
  AOI22X1 U372 ( .A0(n1333), .A1(R3[23]), .B0(n886), .B1(R14[23]), .Y(n973) );
  AOI22X1 U373 ( .A0(n1324), .A1(R0[23]), .B0(n1321), .B1(R15[23]), .Y(n974)
         );
  AOI22X1 U374 ( .A0(n1402), .A1(R1[23]), .B0(n1316), .B1(R12[23]), .Y(n975)
         );
  AOI22X1 U375 ( .A0(n1332), .A1(R3[24]), .B0(n886), .B1(R14[24]), .Y(n965) );
  AOI22X1 U376 ( .A0(n1324), .A1(R0[24]), .B0(n1322), .B1(R15[24]), .Y(n966)
         );
  AOI22X1 U377 ( .A0(n1402), .A1(R1[24]), .B0(n1316), .B1(R12[24]), .Y(n967)
         );
  AOI22X1 U378 ( .A0(n1333), .A1(R3[25]), .B0(n886), .B1(R14[25]), .Y(n957) );
  AOI22X1 U379 ( .A0(n1323), .A1(R0[25]), .B0(n1322), .B1(R15[25]), .Y(n958)
         );
  AOI22X1 U380 ( .A0(n1402), .A1(R1[25]), .B0(n1315), .B1(R12[25]), .Y(n959)
         );
  AOI22X1 U381 ( .A0(n1332), .A1(R3[26]), .B0(n886), .B1(R14[26]), .Y(n949) );
  AOI22X1 U382 ( .A0(n1324), .A1(R0[26]), .B0(n1322), .B1(R15[26]), .Y(n950)
         );
  AOI22X1 U383 ( .A0(n1402), .A1(R1[26]), .B0(n1316), .B1(R12[26]), .Y(n951)
         );
  OR4X2 U384 ( .A(n873), .B(n874), .C(n875), .D(n876), .Y(N152) );
  OR4X2 U385 ( .A(n1072), .B(n1073), .C(n1074), .D(n1075), .Y(N129) );
  OAI221XL U386 ( .A0(n778), .A1(n1320), .B0(n744), .B1(n1317), .C0(n1079), 
        .Y(n1072) );
  OAI221XL U387 ( .A0(n642), .A1(n882), .B0(n676), .B1(n1335), .C0(n1077), .Y(
        n1074) );
  OAI221XL U388 ( .A0(n846), .A1(n1345), .B0(n812), .B1(n1342), .C0(n1076), 
        .Y(n1075) );
  OR4X2 U389 ( .A(n1064), .B(n1065), .C(n1066), .D(n1067), .Y(N130) );
  OAI221XL U390 ( .A0(n777), .A1(n1320), .B0(n743), .B1(n1317), .C0(n1071), 
        .Y(n1064) );
  OAI221XL U391 ( .A0(n709), .A1(n1329), .B0(n607), .B1(n1325), .C0(n1070), 
        .Y(n1065) );
  OAI221XL U392 ( .A0(n641), .A1(n882), .B0(n675), .B1(n1335), .C0(n1069), .Y(
        n1066) );
  OR4X2 U393 ( .A(n1048), .B(n1049), .C(n1050), .D(n1051), .Y(N132) );
  OAI221XL U394 ( .A0(n775), .A1(n1320), .B0(n741), .B1(n1317), .C0(n1055), 
        .Y(n1048) );
  OAI221XL U395 ( .A0(n707), .A1(n1329), .B0(n605), .B1(n1325), .C0(n1054), 
        .Y(n1049) );
  OAI221XL U396 ( .A0(n639), .A1(n882), .B0(n673), .B1(n1335), .C0(n1053), .Y(
        n1050) );
  OR4X2 U397 ( .A(n1040), .B(n1041), .C(n1042), .D(n1043), .Y(N133) );
  OAI221XL U398 ( .A0(n774), .A1(n1320), .B0(n740), .B1(n1317), .C0(n1047), 
        .Y(n1040) );
  OAI221XL U399 ( .A0(n706), .A1(n1329), .B0(n604), .B1(n1325), .C0(n1046), 
        .Y(n1041) );
  OAI221XL U400 ( .A0(n638), .A1(n882), .B0(n672), .B1(n1335), .C0(n1045), .Y(
        n1042) );
  OR4X2 U401 ( .A(n1032), .B(n1033), .C(n1034), .D(n1035), .Y(N134) );
  OAI221XL U402 ( .A0(n773), .A1(n1320), .B0(n739), .B1(n1317), .C0(n1039), 
        .Y(n1032) );
  OAI221XL U403 ( .A0(n705), .A1(n1329), .B0(n603), .B1(n1325), .C0(n1038), 
        .Y(n1033) );
  OAI221XL U404 ( .A0(n637), .A1(n882), .B0(n671), .B1(n1335), .C0(n1037), .Y(
        n1034) );
  OR4X2 U405 ( .A(n1024), .B(n1025), .C(n1026), .D(n1027), .Y(N135) );
  OAI221XL U406 ( .A0(n772), .A1(n1320), .B0(n738), .B1(n1317), .C0(n1031), 
        .Y(n1024) );
  OAI221XL U407 ( .A0(n704), .A1(n1329), .B0(n602), .B1(n1325), .C0(n1030), 
        .Y(n1025) );
  OAI221XL U408 ( .A0(n636), .A1(n882), .B0(n670), .B1(n1335), .C0(n1029), .Y(
        n1026) );
  OR4X2 U409 ( .A(n936), .B(n937), .C(n938), .D(n939), .Y(N146) );
  OAI221XL U410 ( .A0(n761), .A1(n1319), .B0(n727), .B1(n1318), .C0(n943), .Y(
        n936) );
  OAI221XL U411 ( .A0(n693), .A1(n1328), .B0(n591), .B1(n1326), .C0(n942), .Y(
        n937) );
  OAI221XL U412 ( .A0(n625), .A1(n1336), .B0(n659), .B1(n1334), .C0(n941), .Y(
        n938) );
  OR4X2 U413 ( .A(n928), .B(n929), .C(n930), .D(n931), .Y(N147) );
  OAI221XL U414 ( .A0(n760), .A1(n1319), .B0(n726), .B1(n1318), .C0(n935), .Y(
        n928) );
  OAI221XL U415 ( .A0(n692), .A1(n1328), .B0(n590), .B1(n1326), .C0(n934), .Y(
        n929) );
  OAI221XL U416 ( .A0(n624), .A1(n1336), .B0(n658), .B1(n1334), .C0(n933), .Y(
        n930) );
  OR4X2 U417 ( .A(n920), .B(n921), .C(n922), .D(n923), .Y(N148) );
  OAI221XL U418 ( .A0(n759), .A1(n1319), .B0(n725), .B1(n1317), .C0(n927), .Y(
        n920) );
  OAI221XL U419 ( .A0(n691), .A1(n1328), .B0(n589), .B1(n1325), .C0(n926), .Y(
        n921) );
  OAI221XL U420 ( .A0(n623), .A1(n1336), .B0(n657), .B1(n1334), .C0(n925), .Y(
        n922) );
  OR4X2 U421 ( .A(n912), .B(n913), .C(n914), .D(n915), .Y(N149) );
  OAI221XL U422 ( .A0(n758), .A1(n1319), .B0(n724), .B1(n1318), .C0(n919), .Y(
        n912) );
  OAI221XL U423 ( .A0(n690), .A1(n1328), .B0(n588), .B1(n1326), .C0(n918), .Y(
        n913) );
  OAI221XL U424 ( .A0(n622), .A1(n1336), .B0(n656), .B1(n1334), .C0(n917), .Y(
        n914) );
  OR4X2 U425 ( .A(n904), .B(n905), .C(n906), .D(n907), .Y(N150) );
  OAI221XL U426 ( .A0(n757), .A1(n1319), .B0(n723), .B1(n1317), .C0(n911), .Y(
        n904) );
  OAI221XL U427 ( .A0(n689), .A1(n1328), .B0(n587), .B1(n888), .C0(n910), .Y(
        n905) );
  OAI221XL U428 ( .A0(n621), .A1(n1336), .B0(n655), .B1(n1334), .C0(n909), .Y(
        n906) );
  OR4X2 U429 ( .A(n896), .B(n897), .C(n898), .D(n899), .Y(N151) );
  OAI221XL U430 ( .A0(n756), .A1(n1319), .B0(n722), .B1(n1318), .C0(n903), .Y(
        n896) );
  OAI221XL U431 ( .A0(n688), .A1(n1328), .B0(n586), .B1(n888), .C0(n902), .Y(
        n897) );
  OAI221XL U432 ( .A0(n620), .A1(n882), .B0(n654), .B1(n1334), .C0(n901), .Y(
        n898) );
  OR4X2 U433 ( .A(n1080), .B(n1081), .C(n1082), .D(n1083), .Y(N128) );
  OAI221XL U434 ( .A0(n779), .A1(n1320), .B0(n745), .B1(n1318), .C0(n1087), 
        .Y(n1080) );
  OAI221XL U435 ( .A0(n711), .A1(n1329), .B0(n609), .B1(n1326), .C0(n1086), 
        .Y(n1081) );
  OAI221XL U436 ( .A0(n643), .A1(n882), .B0(n677), .B1(n1335), .C0(n1085), .Y(
        n1082) );
  OR4X2 U437 ( .A(n1056), .B(n1057), .C(n1058), .D(n1059), .Y(N131) );
  OAI221XL U438 ( .A0(n776), .A1(n1320), .B0(n742), .B1(n1317), .C0(n1063), 
        .Y(n1056) );
  OAI221XL U439 ( .A0(n708), .A1(n1329), .B0(n606), .B1(n1325), .C0(n1062), 
        .Y(n1057) );
  OAI221XL U440 ( .A0(n640), .A1(n882), .B0(n674), .B1(n1335), .C0(n1061), .Y(
        n1058) );
  OR4X2 U441 ( .A(n1152), .B(n1153), .C(n1154), .D(n1155), .Y(N119) );
  OAI221XL U442 ( .A0(n788), .A1(n1319), .B0(n754), .B1(n1318), .C0(n1164), 
        .Y(n1152) );
  OAI221XL U443 ( .A0(n720), .A1(n1329), .B0(n618), .B1(n1326), .C0(n1161), 
        .Y(n1153) );
  OAI221XL U444 ( .A0(n652), .A1(n1336), .B0(n686), .B1(n1335), .C0(n1160), 
        .Y(n1154) );
  OR4X2 U445 ( .A(n1144), .B(n1145), .C(n1146), .D(n1147), .Y(N120) );
  OAI221XL U446 ( .A0(n787), .A1(n1320), .B0(n753), .B1(n1318), .C0(n1151), 
        .Y(n1144) );
  OAI221XL U447 ( .A0(n719), .A1(n1328), .B0(n617), .B1(n1326), .C0(n1150), 
        .Y(n1145) );
  OAI221XL U448 ( .A0(n651), .A1(n1336), .B0(n685), .B1(n1334), .C0(n1149), 
        .Y(n1146) );
  OR4X2 U449 ( .A(n1136), .B(n1137), .C(n1138), .D(n1139), .Y(N121) );
  OAI221XL U450 ( .A0(n786), .A1(n1319), .B0(n752), .B1(n1318), .C0(n1143), 
        .Y(n1136) );
  OAI221XL U451 ( .A0(n718), .A1(n1329), .B0(n616), .B1(n1326), .C0(n1142), 
        .Y(n1137) );
  OAI221XL U452 ( .A0(n650), .A1(n1336), .B0(n684), .B1(n1335), .C0(n1141), 
        .Y(n1138) );
  OR4X2 U453 ( .A(n1128), .B(n1129), .C(n1130), .D(n1131), .Y(N122) );
  OAI221XL U454 ( .A0(n785), .A1(n1320), .B0(n751), .B1(n1318), .C0(n1135), 
        .Y(n1128) );
  OAI221XL U455 ( .A0(n717), .A1(n1328), .B0(n615), .B1(n1326), .C0(n1134), 
        .Y(n1129) );
  OAI221XL U456 ( .A0(n649), .A1(n1336), .B0(n683), .B1(n1334), .C0(n1133), 
        .Y(n1130) );
  OR4X2 U457 ( .A(n1120), .B(n1121), .C(n1122), .D(n1123), .Y(N123) );
  OAI221XL U458 ( .A0(n784), .A1(n1319), .B0(n750), .B1(n1318), .C0(n1127), 
        .Y(n1120) );
  OAI221XL U459 ( .A0(n716), .A1(n1329), .B0(n614), .B1(n1326), .C0(n1126), 
        .Y(n1121) );
  OAI221XL U460 ( .A0(n648), .A1(n1336), .B0(n682), .B1(n1335), .C0(n1125), 
        .Y(n1122) );
  OR4X2 U461 ( .A(n1112), .B(n1113), .C(n1114), .D(n1115), .Y(N124) );
  OAI221XL U462 ( .A0(n783), .A1(n1320), .B0(n749), .B1(n1318), .C0(n1119), 
        .Y(n1112) );
  OAI221XL U463 ( .A0(n715), .A1(n1328), .B0(n613), .B1(n1326), .C0(n1118), 
        .Y(n1113) );
  OAI221XL U464 ( .A0(n647), .A1(n1336), .B0(n681), .B1(n1334), .C0(n1117), 
        .Y(n1114) );
  OR4X2 U465 ( .A(n1104), .B(n1105), .C(n1106), .D(n1107), .Y(N125) );
  OAI221XL U466 ( .A0(n782), .A1(n1319), .B0(n748), .B1(n1318), .C0(n1111), 
        .Y(n1104) );
  OAI221XL U467 ( .A0(n714), .A1(n1329), .B0(n612), .B1(n1326), .C0(n1110), 
        .Y(n1105) );
  OAI221XL U468 ( .A0(n646), .A1(n1336), .B0(n680), .B1(n1335), .C0(n1109), 
        .Y(n1106) );
  OR4X2 U469 ( .A(n1096), .B(n1097), .C(n1098), .D(n1099), .Y(N126) );
  OAI221XL U470 ( .A0(n781), .A1(n1320), .B0(n747), .B1(n1318), .C0(n1103), 
        .Y(n1096) );
  OAI221XL U471 ( .A0(n713), .A1(n1328), .B0(n611), .B1(n1326), .C0(n1102), 
        .Y(n1097) );
  OAI221XL U472 ( .A0(n645), .A1(n1336), .B0(n679), .B1(n1334), .C0(n1101), 
        .Y(n1098) );
  OR4X2 U473 ( .A(n1088), .B(n1089), .C(n1090), .D(n1091), .Y(N127) );
  OAI221XL U474 ( .A0(n780), .A1(n1320), .B0(n746), .B1(n1318), .C0(n1095), 
        .Y(n1088) );
  OAI221XL U475 ( .A0(n712), .A1(n1329), .B0(n610), .B1(n1326), .C0(n1094), 
        .Y(n1089) );
  OAI221XL U476 ( .A0(n644), .A1(n882), .B0(n678), .B1(n1334), .C0(n1093), .Y(
        n1090) );
  OR4X2 U477 ( .A(n1016), .B(n1017), .C(n1018), .D(n1019), .Y(N136) );
  OAI221XL U478 ( .A0(n771), .A1(n1320), .B0(n737), .B1(n1317), .C0(n1023), 
        .Y(n1016) );
  OAI221XL U479 ( .A0(n703), .A1(n1329), .B0(n601), .B1(n1325), .C0(n1022), 
        .Y(n1017) );
  OAI221XL U480 ( .A0(n635), .A1(n882), .B0(n669), .B1(n1335), .C0(n1021), .Y(
        n1018) );
  OR4X2 U481 ( .A(n1008), .B(n1009), .C(n1010), .D(n1011), .Y(N137) );
  OAI221XL U482 ( .A0(n770), .A1(n1320), .B0(n736), .B1(n1317), .C0(n1015), 
        .Y(n1008) );
  OAI221XL U483 ( .A0(n702), .A1(n1329), .B0(n600), .B1(n1325), .C0(n1014), 
        .Y(n1009) );
  OAI221XL U484 ( .A0(n634), .A1(n1336), .B0(n668), .B1(n1335), .C0(n1013), 
        .Y(n1010) );
  OR4X2 U485 ( .A(n1000), .B(n1001), .C(n1002), .D(n1003), .Y(N138) );
  OAI221XL U486 ( .A0(n769), .A1(n1320), .B0(n735), .B1(n1317), .C0(n1007), 
        .Y(n1000) );
  OAI221XL U487 ( .A0(n701), .A1(n1329), .B0(n599), .B1(n1325), .C0(n1006), 
        .Y(n1001) );
  OAI221XL U488 ( .A0(n633), .A1(n1336), .B0(n667), .B1(n1335), .C0(n1005), 
        .Y(n1002) );
  OR4X2 U489 ( .A(n992), .B(n993), .C(n994), .D(n995), .Y(N139) );
  OAI221XL U490 ( .A0(n768), .A1(n1320), .B0(n734), .B1(n1317), .C0(n999), .Y(
        n992) );
  OAI221XL U491 ( .A0(n700), .A1(n1329), .B0(n598), .B1(n1325), .C0(n998), .Y(
        n993) );
  OAI221XL U492 ( .A0(n632), .A1(n1336), .B0(n666), .B1(n1335), .C0(n997), .Y(
        n994) );
  OR4X2 U493 ( .A(n984), .B(n985), .C(n986), .D(n987), .Y(N140) );
  OAI221XL U494 ( .A0(n767), .A1(n1319), .B0(n733), .B1(n1317), .C0(n991), .Y(
        n984) );
  OAI221XL U495 ( .A0(n699), .A1(n1328), .B0(n597), .B1(n1325), .C0(n990), .Y(
        n985) );
  OAI221XL U496 ( .A0(n631), .A1(n1336), .B0(n665), .B1(n1335), .C0(n989), .Y(
        n986) );
  OR4X2 U497 ( .A(n976), .B(n977), .C(n978), .D(n979), .Y(N141) );
  OAI221XL U498 ( .A0(n766), .A1(n1319), .B0(n732), .B1(n1317), .C0(n983), .Y(
        n976) );
  OAI221XL U499 ( .A0(n698), .A1(n1328), .B0(n596), .B1(n888), .C0(n982), .Y(
        n977) );
  OAI221XL U500 ( .A0(n630), .A1(n882), .B0(n664), .B1(n1334), .C0(n981), .Y(
        n978) );
  OR4X2 U501 ( .A(n968), .B(n969), .C(n970), .D(n971), .Y(N142) );
  OAI221XL U502 ( .A0(n765), .A1(n1319), .B0(n731), .B1(n1318), .C0(n975), .Y(
        n968) );
  OAI221XL U503 ( .A0(n697), .A1(n1328), .B0(n595), .B1(n888), .C0(n974), .Y(
        n969) );
  OAI221XL U504 ( .A0(n629), .A1(n882), .B0(n663), .B1(n1334), .C0(n973), .Y(
        n970) );
  OR4X2 U505 ( .A(n960), .B(n961), .C(n962), .D(n963), .Y(N143) );
  OAI221XL U506 ( .A0(n764), .A1(n1319), .B0(n730), .B1(n1317), .C0(n967), .Y(
        n960) );
  OAI221XL U507 ( .A0(n696), .A1(n1328), .B0(n594), .B1(n888), .C0(n966), .Y(
        n961) );
  OAI221XL U508 ( .A0(n628), .A1(n882), .B0(n662), .B1(n1334), .C0(n965), .Y(
        n962) );
  OR4X2 U509 ( .A(n952), .B(n953), .C(n954), .D(n955), .Y(N144) );
  OAI221XL U510 ( .A0(n763), .A1(n1319), .B0(n729), .B1(n1318), .C0(n959), .Y(
        n952) );
  OAI221XL U511 ( .A0(n695), .A1(n1328), .B0(n593), .B1(n888), .C0(n958), .Y(
        n953) );
  OAI221XL U512 ( .A0(n627), .A1(n882), .B0(n661), .B1(n1334), .C0(n957), .Y(
        n954) );
  OR4X2 U513 ( .A(n944), .B(n945), .C(n946), .D(n947), .Y(N145) );
  OAI221XL U514 ( .A0(n762), .A1(n1319), .B0(n728), .B1(n1317), .C0(n951), .Y(
        n944) );
  OAI221XL U515 ( .A0(n694), .A1(n1328), .B0(n592), .B1(n888), .C0(n950), .Y(
        n945) );
  OAI221XL U516 ( .A0(n626), .A1(n882), .B0(n660), .B1(n1334), .C0(n949), .Y(
        n946) );
  NOR2X1 U517 ( .A(n1405), .B(counter_2[1]), .Y(n872) );
  NOR2X1 U518 ( .A(counter_2[2]), .B(counter_2[1]), .Y(n1159) );
  OR3XL U519 ( .A(n584), .B(p_s_flag_in), .C(n1401), .Y(n225) );
  OR3XL U520 ( .A(counter_1[0]), .B(p_s_flag_in), .C(n1401), .Y(n226) );
  OR3XL U521 ( .A(counter_1[1]), .B(p_s_flag_in), .C(n584), .Y(n227) );
  INVX1 U522 ( .A(counter_1[1]), .Y(n1401) );
  INVX1 U523 ( .A(n870), .Y(n1403) );
  AOI221X1 U524 ( .A0(counter_2[0]), .A1(n871), .B0(n861), .B1(counter_2[2]), 
        .C0(n872), .Y(n870) );
  NAND2X1 U525 ( .A(n867), .B(n868), .Y(N52) );
  OAI2BB1X1 U526 ( .A0N(n869), .A1N(counter_2[0]), .B0(counter_2[3]), .Y(n868)
         );
  XNOR2X1 U527 ( .A(n1404), .B(counter_2[0]), .Y(N50) );
  XNOR2X1 U528 ( .A(n1401), .B(counter_1[0]), .Y(N26) );
  AOI22X1 U529 ( .A0(n1323), .A1(n145), .B0(n1322), .B1(R15[10]), .Y(n1078) );
  OAI221XL U530 ( .A0(n619), .A1(n882), .B0(n653), .B1(n1334), .C0(n884), .Y(
        n875) );
  OAI221XL U531 ( .A0(n687), .A1(n1328), .B0(n585), .B1(n888), .C0(n889), .Y(
        n874) );
  OAI221XL U532 ( .A0(n755), .A1(n1319), .B0(n721), .B1(n1318), .C0(n894), .Y(
        n873) );
  OAI221XL U533 ( .A0(n823), .A1(n1344), .B0(n789), .B1(n1343), .C0(n879), .Y(
        n876) );
  AOI22X1 U534 ( .A0(n1333), .A1(n147), .B0(n886), .B1(n91), .Y(n884) );
  AOI22X1 U535 ( .A0(n1323), .A1(n149), .B0(n1322), .B1(n93), .Y(n889) );
  AOI22X1 U536 ( .A0(n1402), .A1(n150), .B0(n1316), .B1(n89), .Y(n894) );
  AOI22X1 U537 ( .A0(n1341), .A1(n151), .B0(n1338), .B1(n90), .Y(n879) );
endmodule


module fft ( clk, rst_n, data_in, data_out );
  input [33:0] data_in;
  output [33:0] data_out;
  input clk, rst_n;
  wire   s_p_flag, mux_flag, demux_flag, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36;
  wire   [2:0] rotation;
  wire   [135:0] data_1;
  wire   [135:0] data_2;
  wire   [135:0] data_4;
  wire   [135:0] data_3;

  ctrl ctrl0 ( .clk(clk), .rst_n(rst_n), .s_p_flag_in(s_p_flag), .mux_flag(
        mux_flag), .rotation(rotation), .demux_flag(demux_flag) );
  s_p s_p0 ( .clk(clk), .rst_n(rst_n), .data_in_1(data_in), .data_out_1(data_1), .s_p_flag_out(s_p_flag) );
  mux mux0 ( .mux_flag(mux_flag), .clk(clk), .rst_n(rst_n), .data_in_1(data_2), 
        .data_in_2(data_1), .data_out(data_3), .data_in_3_33_(n9), 
        .data_in_3_32_(n26), .data_in_3_31_(n19), .data_in_3_30_(n20), 
        .data_in_3_29_(n25), .data_in_3_28_(n14), .data_in_3_27_(n32), 
        .data_in_3_26_(data_4[26]), .data_in_3_25_(data_4[25]), 
        .data_in_3_24_(data_4[24]), .data_in_3_23_(data_4[23]), 
        .data_in_3_22_(n7), .data_in_3_21_(data_4[21]), .data_in_3_20_(
        data_4[20]), .data_in_3_19_(data_4[19]), .data_in_3_18_(data_4[18]), 
        .data_in_3_17_(data_4[17]), .data_in_3_16_(n8), .data_in_3_15_(n29), 
        .data_in_3_14_(n2), .data_in_3_13_(n21), .data_in_3_12_(data_4[12]), 
        .data_in_3_11_(data_4[11]), .data_in_3_10_(n24), .data_in_3_9_(n1), 
        .data_in_3_8_(data_4[8]), .data_in_3_7_(data_4[7]), .data_in_3_6_(
        data_4[6]), .data_in_3_5_(data_4[5]), .data_in_3_4_(data_4[4]), 
        .data_in_3_3_(data_4[3]), .data_in_3_2_(data_4[2]), .data_in_3_1_(
        data_4[1]), .data_in_3_0_(data_4[0]) );
  butterfly butterfly0 ( .calc_in(data_3), .rotation(rotation), .calc_out(
        data_4) );
  reg1 reg10 ( .clk(clk), .rst_n(rst_n), .data_in_2({n30, data_4[134:133], n17, 
        data_4[131], n22, data_4[129:108], n11, data_4[106:101], n33, n15, n23, 
        n34, n18, data_4[95:85], n31, n12, n10, data_4[81:80], n35, 
        data_4[78:68], n27, n28, n13, data_4[64:50], n36, data_4[48:0]}), 
        .reg_datain_flag(demux_flag), .data_out_2(data_2) );
  p_s p_s0 ( .clk(clk), .rst_n(rst_n), .data_in_3({n30, data_4[134:131], n22, 
        n4, data_4[128:108], n11, data_4[106:101], n33, n15, n23, n34, n18, 
        data_4[95:85], n31, n12, n10, data_4[81:80], n35, n6, data_4[77:68], 
        n27, n28, n13, data_4[64:50], n36, data_4[48:0]}), .p_s_flag_in(
        demux_flag), .data_out_3(data_out) );
  BUFX3 U1 ( .A(data_4[15]), .Y(n29) );
  BUFX20 U2 ( .A(data_4[79]), .Y(n35) );
  BUFX20 U3 ( .A(data_4[66]), .Y(n28) );
  BUFX20 U4 ( .A(data_4[98]), .Y(n23) );
  BUFX20 U5 ( .A(data_4[96]), .Y(n18) );
  BUFX16 U6 ( .A(data_4[97]), .Y(n34) );
  BUFX16 U7 ( .A(data_4[83]), .Y(n12) );
  BUFX4 U8 ( .A(data_4[107]), .Y(n11) );
  BUFX3 U9 ( .A(data_4[22]), .Y(n7) );
  DLY1X1 U10 ( .A(data_4[9]), .Y(n1) );
  BUFX20 U11 ( .A(data_4[99]), .Y(n15) );
  BUFX16 U12 ( .A(data_4[82]), .Y(n10) );
  CLKINVX3 U13 ( .A(data_4[129]), .Y(n3) );
  BUFX16 U14 ( .A(data_4[135]), .Y(n30) );
  DLY1X1 U15 ( .A(data_4[14]), .Y(n2) );
  INVX4 U16 ( .A(n3), .Y(n4) );
  CLKINVX8 U17 ( .A(data_4[78]), .Y(n5) );
  INVX8 U18 ( .A(n5), .Y(n6) );
  BUFX20 U19 ( .A(data_4[65]), .Y(n13) );
  DLY1X1 U20 ( .A(data_4[16]), .Y(n8) );
  BUFX20 U21 ( .A(data_4[130]), .Y(n22) );
  DLY1X1 U22 ( .A(data_4[33]), .Y(n9) );
  BUFX20 U23 ( .A(data_4[67]), .Y(n27) );
  BUFX20 U24 ( .A(data_4[84]), .Y(n31) );
  BUFX20 U25 ( .A(data_4[100]), .Y(n33) );
  BUFX20 U26 ( .A(data_4[49]), .Y(n36) );
  DLY1X1 U27 ( .A(data_4[28]), .Y(n14) );
  CLKINVX8 U28 ( .A(data_4[132]), .Y(n16) );
  INVX8 U29 ( .A(n16), .Y(n17) );
  DLY1X1 U30 ( .A(data_4[31]), .Y(n19) );
  DLY1X1 U31 ( .A(data_4[30]), .Y(n20) );
  DLY1X1 U32 ( .A(data_4[13]), .Y(n21) );
  DLY1X1 U33 ( .A(data_4[10]), .Y(n24) );
  DLY1X1 U34 ( .A(data_4[29]), .Y(n25) );
  DLY1X1 U35 ( .A(data_4[32]), .Y(n26) );
  DLY1X1 U36 ( .A(data_4[27]), .Y(n32) );
endmodule


module fft_chip ( clk, rst_n, data_in, data_out );
  input [33:0] data_in;
  output [33:0] data_out;
  input clk, rst_n;
  wire   net_clk, net_rst_n;
  wire   [33:0] net_data_in;
  wire   [33:0] net_data_out;

  PIW PIW_clk ( .PAD(clk), .C(net_clk) );
  PIW PIW_rst_n ( .PAD(rst_n), .C(net_rst_n) );
  PIW PIW_data_in0 ( .PAD(data_in[0]), .C(net_data_in[0]) );
  PIW PIW_data_in1 ( .PAD(data_in[1]), .C(net_data_in[1]) );
  PIW PIW_data_in2 ( .PAD(data_in[2]), .C(net_data_in[2]) );
  PIW PIW_data_in3 ( .PAD(data_in[3]), .C(net_data_in[3]) );
  PIW PIW_data_in4 ( .PAD(data_in[4]), .C(net_data_in[4]) );
  PIW PIW_data_in5 ( .PAD(data_in[5]), .C(net_data_in[5]) );
  PIW PIW_data_in6 ( .PAD(data_in[6]), .C(net_data_in[6]) );
  PIW PIW_data_in7 ( .PAD(data_in[7]), .C(net_data_in[7]) );
  PIW PIW_data_in8 ( .PAD(data_in[8]), .C(net_data_in[8]) );
  PIW PIW_data_in9 ( .PAD(data_in[9]), .C(net_data_in[9]) );
  PIW PIW_data_in10 ( .PAD(data_in[10]), .C(net_data_in[10]) );
  PIW PIW_data_in11 ( .PAD(data_in[11]), .C(net_data_in[11]) );
  PIW PIW_data_in12 ( .PAD(data_in[12]), .C(net_data_in[12]) );
  PIW PIW_data_in13 ( .PAD(data_in[13]), .C(net_data_in[13]) );
  PIW PIW_data_in14 ( .PAD(data_in[14]), .C(net_data_in[14]) );
  PIW PIW_data_in15 ( .PAD(data_in[15]), .C(net_data_in[15]) );
  PIW PIW_data_in16 ( .PAD(data_in[16]), .C(net_data_in[16]) );
  PIW PIW_data_in17 ( .PAD(data_in[17]), .C(net_data_in[17]) );
  PIW PIW_data_in18 ( .PAD(data_in[18]), .C(net_data_in[18]) );
  PIW PIW_data_in19 ( .PAD(data_in[19]), .C(net_data_in[19]) );
  PIW PIW_data_in20 ( .PAD(data_in[20]), .C(net_data_in[20]) );
  PIW PIW_data_in21 ( .PAD(data_in[21]), .C(net_data_in[21]) );
  PIW PIW_data_in22 ( .PAD(data_in[22]), .C(net_data_in[22]) );
  PIW PIW_data_in23 ( .PAD(data_in[23]), .C(net_data_in[23]) );
  PIW PIW_data_in24 ( .PAD(data_in[24]), .C(net_data_in[24]) );
  PIW PIW_data_in25 ( .PAD(data_in[25]), .C(net_data_in[25]) );
  PIW PIW_data_in26 ( .PAD(data_in[26]), .C(net_data_in[26]) );
  PIW PIW_data_in27 ( .PAD(data_in[27]), .C(net_data_in[27]) );
  PIW PIW_data_in28 ( .PAD(data_in[28]), .C(net_data_in[28]) );
  PIW PIW_data_in29 ( .PAD(data_in[29]), .C(net_data_in[29]) );
  PIW PIW_data_in30 ( .PAD(data_in[30]), .C(net_data_in[30]) );
  PIW PIW_data_in31 ( .PAD(data_in[31]), .C(net_data_in[31]) );
  PIW PIW_data_in32 ( .PAD(data_in[32]), .C(net_data_in[32]) );
  PIW PIW_data_in33 ( .PAD(data_in[33]), .C(net_data_in[33]) );
  PO8W PO8W_data_out0 ( .I(net_data_out[0]), .PAD(data_out[0]) );
  PO8W PO8W_data_out1 ( .I(net_data_out[1]), .PAD(data_out[1]) );
  PO8W PO8W_data_out2 ( .I(net_data_out[2]), .PAD(data_out[2]) );
  PO8W PO8W_data_out3 ( .I(net_data_out[3]), .PAD(data_out[3]) );
  PO8W PO8W_data_out4 ( .I(net_data_out[4]), .PAD(data_out[4]) );
  PO8W PO8W_data_out5 ( .I(net_data_out[5]), .PAD(data_out[5]) );
  PO8W PO8W_data_out6 ( .I(net_data_out[6]), .PAD(data_out[6]) );
  PO8W PO8W_data_out7 ( .I(net_data_out[7]), .PAD(data_out[7]) );
  PO8W PO8W_data_out8 ( .I(net_data_out[8]), .PAD(data_out[8]) );
  PO8W PO8W_data_out9 ( .I(net_data_out[9]), .PAD(data_out[9]) );
  PO8W PO8W_data_out10 ( .I(net_data_out[10]), .PAD(data_out[10]) );
  PO8W PO8W_data_out11 ( .I(net_data_out[11]), .PAD(data_out[11]) );
  PO8W PO8W_data_out12 ( .I(net_data_out[12]), .PAD(data_out[12]) );
  PO8W PO8W_data_out13 ( .I(net_data_out[13]), .PAD(data_out[13]) );
  PO8W PO8W_data_out14 ( .I(net_data_out[14]), .PAD(data_out[14]) );
  PO8W PO8W_data_out15 ( .I(net_data_out[15]), .PAD(data_out[15]) );
  PO8W PO8W_data_out16 ( .I(net_data_out[16]), .PAD(data_out[16]) );
  PO8W PO8W_data_out17 ( .I(net_data_out[17]), .PAD(data_out[17]) );
  PO8W PO8W_data_out18 ( .I(net_data_out[18]), .PAD(data_out[18]) );
  PO8W PO8W_data_out19 ( .I(net_data_out[19]), .PAD(data_out[19]) );
  PO8W PO8W_data_out20 ( .I(net_data_out[20]), .PAD(data_out[20]) );
  PO8W PO8W_data_out21 ( .I(net_data_out[21]), .PAD(data_out[21]) );
  PO8W PO8W_data_out22 ( .I(net_data_out[22]), .PAD(data_out[22]) );
  PO8W PO8W_data_out23 ( .I(net_data_out[23]), .PAD(data_out[23]) );
  PO8W PO8W_data_out24 ( .I(net_data_out[24]), .PAD(data_out[24]) );
  PO8W PO8W_data_out25 ( .I(net_data_out[25]), .PAD(data_out[25]) );
  PO8W PO8W_data_out26 ( .I(net_data_out[26]), .PAD(data_out[26]) );
  PO8W PO8W_data_out27 ( .I(net_data_out[27]), .PAD(data_out[27]) );
  PO8W PO8W_data_out28 ( .I(net_data_out[28]), .PAD(data_out[28]) );
  PO8W PO8W_data_out29 ( .I(net_data_out[29]), .PAD(data_out[29]) );
  PO8W PO8W_data_out30 ( .I(net_data_out[30]), .PAD(data_out[30]) );
  PO8W PO8W_data_out31 ( .I(net_data_out[31]), .PAD(data_out[31]) );
  PO8W PO8W_data_out32 ( .I(net_data_out[32]), .PAD(data_out[32]) );
  PO8W PO8W_data_out33 ( .I(net_data_out[33]), .PAD(data_out[33]) );
  fft inst_fft ( .clk(net_clk), .rst_n(net_rst_n), .data_in(net_data_in), 
        .data_out(net_data_out) );
endmodule

