//
// Author: @xxx, copyright 2020
// e-mail: 
// School: Shanghai Jiao Tong University
//
// File Name:
//
// Type: 
//
// Purpose:
// xxx
//
// Details:
// - 
//
// Release History:
// - Version 1.0 20/03/19: Create;
//
// Notes:
// - xxx.
//

module template(xxx, yyy)

  input xxx; // xxx

  output yyy;

  parameter IDLE;

  wire xxx;

  reg yyy;

// aaa_bbb_ccc // xxx

always @ (*) begin
	if (xxx)
		yyy <= 1'b0;
	else
		yyy <= 1'b1;
end