
module ctrl ( clk, rst_n, s_p_flag_in, mux_flag, rotation, demux_flag );
  output [2:0] rotation;
  input clk, rst_n, s_p_flag_in;
  output mux_flag, demux_flag;
  wire   N17, N18, N19, n3, n1, n2;
  wire   [2:0] core_tick;

  DFFRHQX4 mux_flag_reg ( .D(core_tick[2]), .CK(clk), .RN(rst_n), .Q(mux_flag)
         );
  DFFRHQX1 core_tick_reg_2_ ( .D(N19), .CK(clk), .RN(rst_n), .Q(core_tick[2])
         );
  DFFRHQX1 core_tick_reg_1_ ( .D(N18), .CK(clk), .RN(rst_n), .Q(core_tick[1])
         );
  DFFRHQX1 core_tick_reg_0_ ( .D(N17), .CK(clk), .RN(rst_n), .Q(core_tick[0])
         );
  DFFRHQX1 demux_flag_reg ( .D(n2), .CK(clk), .RN(rst_n), .Q(demux_flag) );
  DFFRHQX4 rotation_reg_1_ ( .D(core_tick[1]), .CK(clk), .RN(rst_n), .Q(
        rotation[1]) );
  DFFRHQX4 rotation_reg_0_ ( .D(core_tick[0]), .CK(clk), .RN(rst_n), .Q(
        rotation[0]) );
  DFFRHQX4 rotation_reg_2_ ( .D(core_tick[2]), .CK(clk), .RN(rst_n), .Q(
        rotation[2]) );
  INVX1 U3 ( .A(core_tick[2]), .Y(n2) );
  AOI2BB1X1 U4 ( .A0N(n1), .A1N(core_tick[1]), .B0(core_tick[0]), .Y(N17) );
  OR2X2 U5 ( .A(s_p_flag_in), .B(core_tick[2]), .Y(n1) );
  XOR2X1 U6 ( .A(core_tick[1]), .B(core_tick[0]), .Y(N18) );
  XOR2X1 U7 ( .A(n2), .B(n3), .Y(N19) );
  NAND2X1 U8 ( .A(core_tick[1]), .B(core_tick[0]), .Y(n3) );
endmodule


module s_p ( clk, rst_n, data_in_1, data_out_1, s_p_flag_out );
  input [33:0] data_in_1;
  output [135:0] data_out_1;
  input clk, rst_n;
  output s_p_flag_out;
  wire   N13, N14, N15, N171, N230, n550, n551, n552, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n970, n971, n972, n973, n974, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
         n1037, n1038, n1039, n1040, n1041, n1042, n1043;
  wire   [3:0] counter;
  wire   [33:0] R15;
  wire   [33:0] R11;
  wire   [33:0] R7;
  wire   [33:0] R3;
  wire   [33:0] R12;
  wire   [33:0] R8;
  wire   [33:0] R4;
  wire   [33:0] R0;
  wire   [33:0] R13;
  wire   [33:0] R9;
  wire   [33:0] R5;
  wire   [33:0] R1;
  wire   [33:0] R14;
  wire   [33:0] R10;
  wire   [33:0] R6;
  wire   [33:0] R2;

  EDFFX1 R13_reg_33_ ( .D(data_in_1[33]), .E(n1010), .CK(clk), .Q(R13[33]) );
  EDFFX1 R13_reg_32_ ( .D(data_in_1[32]), .E(n1009), .CK(clk), .Q(R13[32]) );
  EDFFX1 R13_reg_31_ ( .D(data_in_1[31]), .E(n1011), .CK(clk), .Q(R13[31]) );
  EDFFX1 R13_reg_30_ ( .D(data_in_1[30]), .E(n1010), .CK(clk), .Q(R13[30]) );
  EDFFX1 R13_reg_29_ ( .D(data_in_1[29]), .E(n1009), .CK(clk), .Q(R13[29]) );
  EDFFX1 R13_reg_28_ ( .D(data_in_1[28]), .E(n1011), .CK(clk), .Q(R13[28]) );
  EDFFX1 R13_reg_27_ ( .D(data_in_1[27]), .E(n1010), .CK(clk), .Q(R13[27]) );
  EDFFX1 R13_reg_26_ ( .D(data_in_1[26]), .E(n1009), .CK(clk), .Q(R13[26]) );
  EDFFX1 R13_reg_25_ ( .D(data_in_1[25]), .E(n1011), .CK(clk), .Q(R13[25]) );
  EDFFX1 R13_reg_24_ ( .D(data_in_1[24]), .E(n1010), .CK(clk), .Q(R13[24]) );
  EDFFX1 R13_reg_23_ ( .D(data_in_1[23]), .E(n1009), .CK(clk), .Q(R13[23]) );
  EDFFX1 R13_reg_22_ ( .D(data_in_1[22]), .E(n1008), .CK(clk), .Q(R13[22]) );
  EDFFX1 R13_reg_21_ ( .D(data_in_1[21]), .E(n1010), .CK(clk), .Q(R13[21]) );
  EDFFX1 R13_reg_20_ ( .D(data_in_1[20]), .E(n1009), .CK(clk), .Q(R13[20]) );
  EDFFX1 R13_reg_19_ ( .D(data_in_1[19]), .E(n1011), .CK(clk), .Q(R13[19]) );
  EDFFX1 R13_reg_18_ ( .D(data_in_1[18]), .E(n1010), .CK(clk), .Q(R13[18]) );
  EDFFX1 R13_reg_17_ ( .D(data_in_1[17]), .E(n1010), .CK(clk), .Q(R13[17]) );
  EDFFX1 R13_reg_16_ ( .D(data_in_1[16]), .E(n1008), .CK(clk), .Q(R13[16]) );
  EDFFX1 R13_reg_15_ ( .D(data_in_1[15]), .E(n1011), .CK(clk), .Q(R13[15]) );
  EDFFX1 R13_reg_14_ ( .D(data_in_1[14]), .E(n1009), .CK(clk), .Q(R13[14]) );
  EDFFX1 R13_reg_13_ ( .D(data_in_1[13]), .E(n1011), .CK(clk), .Q(R13[13]) );
  EDFFX1 R13_reg_12_ ( .D(data_in_1[12]), .E(n1010), .CK(clk), .Q(R13[12]) );
  EDFFX1 R13_reg_11_ ( .D(data_in_1[11]), .E(n1009), .CK(clk), .Q(R13[11]) );
  EDFFX1 R13_reg_10_ ( .D(data_in_1[10]), .E(n1008), .CK(clk), .Q(R13[10]) );
  EDFFX1 R13_reg_9_ ( .D(data_in_1[9]), .E(n1009), .CK(clk), .Q(R13[9]) );
  EDFFX1 R13_reg_8_ ( .D(data_in_1[8]), .E(n1008), .CK(clk), .Q(R13[8]) );
  EDFFX1 R13_reg_7_ ( .D(data_in_1[7]), .E(n1008), .CK(clk), .Q(R13[7]) );
  EDFFX1 R13_reg_6_ ( .D(data_in_1[6]), .E(n1008), .CK(clk), .Q(R13[6]) );
  EDFFX1 R13_reg_5_ ( .D(data_in_1[5]), .E(n1010), .CK(clk), .Q(R13[5]) );
  EDFFX1 R13_reg_4_ ( .D(data_in_1[4]), .E(n1008), .CK(clk), .Q(R13[4]) );
  EDFFX1 R13_reg_3_ ( .D(data_in_1[3]), .E(n1008), .CK(clk), .Q(R13[3]) );
  EDFFX1 R13_reg_2_ ( .D(data_in_1[2]), .E(n1010), .CK(clk), .Q(R13[2]) );
  EDFFX1 R13_reg_1_ ( .D(data_in_1[1]), .E(n1011), .CK(clk), .Q(R13[1]) );
  EDFFX1 R13_reg_0_ ( .D(data_in_1[0]), .E(n1008), .CK(clk), .Q(R13[0]) );
  EDFFX1 R1_reg_33_ ( .D(data_in_1[33]), .E(n978), .CK(clk), .Q(R1[33]) );
  EDFFX1 R1_reg_32_ ( .D(data_in_1[32]), .E(n978), .CK(clk), .Q(R1[32]) );
  EDFFX1 R1_reg_31_ ( .D(data_in_1[31]), .E(n978), .CK(clk), .Q(R1[31]) );
  EDFFX1 R1_reg_30_ ( .D(data_in_1[30]), .E(n978), .CK(clk), .Q(R1[30]) );
  EDFFX1 R1_reg_29_ ( .D(data_in_1[29]), .E(n978), .CK(clk), .Q(R1[29]) );
  EDFFX1 R1_reg_28_ ( .D(data_in_1[28]), .E(n978), .CK(clk), .Q(R1[28]) );
  EDFFX1 R1_reg_27_ ( .D(data_in_1[27]), .E(n978), .CK(clk), .Q(R1[27]) );
  EDFFX1 R1_reg_26_ ( .D(data_in_1[26]), .E(n978), .CK(clk), .Q(R1[26]) );
  EDFFX1 R1_reg_25_ ( .D(data_in_1[25]), .E(n978), .CK(clk), .Q(R1[25]) );
  EDFFX1 R1_reg_24_ ( .D(data_in_1[24]), .E(n978), .CK(clk), .Q(R1[24]) );
  EDFFX1 R1_reg_23_ ( .D(data_in_1[23]), .E(n978), .CK(clk), .Q(R1[23]) );
  EDFFX1 R1_reg_22_ ( .D(data_in_1[22]), .E(n978), .CK(clk), .Q(R1[22]) );
  EDFFX1 R1_reg_21_ ( .D(data_in_1[21]), .E(n979), .CK(clk), .Q(R1[21]) );
  EDFFX1 R1_reg_20_ ( .D(data_in_1[20]), .E(n979), .CK(clk), .Q(R1[20]) );
  EDFFX1 R1_reg_19_ ( .D(data_in_1[19]), .E(n979), .CK(clk), .Q(R1[19]) );
  EDFFX1 R1_reg_18_ ( .D(data_in_1[18]), .E(n979), .CK(clk), .Q(R1[18]) );
  EDFFX1 R1_reg_17_ ( .D(data_in_1[17]), .E(n979), .CK(clk), .Q(R1[17]) );
  EDFFX1 R1_reg_16_ ( .D(data_in_1[16]), .E(n979), .CK(clk), .Q(R1[16]) );
  EDFFX1 R1_reg_15_ ( .D(data_in_1[15]), .E(n979), .CK(clk), .Q(R1[15]) );
  EDFFX1 R1_reg_14_ ( .D(data_in_1[14]), .E(n979), .CK(clk), .Q(R1[14]) );
  EDFFX1 R1_reg_13_ ( .D(data_in_1[13]), .E(n979), .CK(clk), .Q(R1[13]) );
  EDFFX1 R1_reg_12_ ( .D(data_in_1[12]), .E(n979), .CK(clk), .Q(R1[12]) );
  EDFFX1 R1_reg_11_ ( .D(data_in_1[11]), .E(n979), .CK(clk), .Q(R1[11]) );
  EDFFX1 R1_reg_10_ ( .D(data_in_1[10]), .E(n979), .CK(clk), .Q(R1[10]) );
  EDFFX1 R1_reg_9_ ( .D(data_in_1[9]), .E(n978), .CK(clk), .Q(R1[9]) );
  EDFFX1 R1_reg_8_ ( .D(data_in_1[8]), .E(n979), .CK(clk), .Q(R1[8]) );
  EDFFX1 R1_reg_7_ ( .D(data_in_1[7]), .E(n978), .CK(clk), .Q(R1[7]) );
  EDFFX1 R1_reg_6_ ( .D(data_in_1[6]), .E(n979), .CK(clk), .Q(R1[6]) );
  EDFFX1 R1_reg_5_ ( .D(data_in_1[5]), .E(n978), .CK(clk), .Q(R1[5]) );
  EDFFX1 R1_reg_4_ ( .D(data_in_1[4]), .E(n979), .CK(clk), .Q(R1[4]) );
  EDFFX1 R1_reg_3_ ( .D(data_in_1[3]), .E(n978), .CK(clk), .Q(R1[3]) );
  EDFFX1 R1_reg_2_ ( .D(data_in_1[2]), .E(n979), .CK(clk), .Q(R1[2]) );
  EDFFX1 R1_reg_1_ ( .D(data_in_1[1]), .E(n978), .CK(clk), .Q(R1[1]) );
  EDFFX1 R1_reg_0_ ( .D(data_in_1[0]), .E(n979), .CK(clk), .Q(R1[0]) );
  EDFFX1 R5_reg_33_ ( .D(data_in_1[33]), .E(n986), .CK(clk), .Q(R5[33]) );
  EDFFX1 R5_reg_32_ ( .D(data_in_1[32]), .E(n986), .CK(clk), .Q(R5[32]) );
  EDFFX1 R5_reg_31_ ( .D(data_in_1[31]), .E(n986), .CK(clk), .Q(R5[31]) );
  EDFFX1 R5_reg_30_ ( .D(data_in_1[30]), .E(n986), .CK(clk), .Q(R5[30]) );
  EDFFX1 R5_reg_29_ ( .D(data_in_1[29]), .E(n986), .CK(clk), .Q(R5[29]) );
  EDFFX1 R5_reg_28_ ( .D(data_in_1[28]), .E(n986), .CK(clk), .Q(R5[28]) );
  EDFFX1 R5_reg_27_ ( .D(data_in_1[27]), .E(n986), .CK(clk), .Q(R5[27]) );
  EDFFX1 R5_reg_26_ ( .D(data_in_1[26]), .E(n986), .CK(clk), .Q(R5[26]) );
  EDFFX1 R5_reg_25_ ( .D(data_in_1[25]), .E(n986), .CK(clk), .Q(R5[25]) );
  EDFFX1 R5_reg_24_ ( .D(data_in_1[24]), .E(n986), .CK(clk), .Q(R5[24]) );
  EDFFX1 R5_reg_23_ ( .D(data_in_1[23]), .E(n986), .CK(clk), .Q(R5[23]) );
  EDFFX1 R5_reg_22_ ( .D(data_in_1[22]), .E(n986), .CK(clk), .Q(R5[22]) );
  EDFFX1 R5_reg_21_ ( .D(data_in_1[21]), .E(n987), .CK(clk), .Q(R5[21]) );
  EDFFX1 R5_reg_20_ ( .D(data_in_1[20]), .E(n987), .CK(clk), .Q(R5[20]) );
  EDFFX1 R5_reg_19_ ( .D(data_in_1[19]), .E(n987), .CK(clk), .Q(R5[19]) );
  EDFFX1 R5_reg_18_ ( .D(data_in_1[18]), .E(n987), .CK(clk), .Q(R5[18]) );
  EDFFX1 R5_reg_17_ ( .D(data_in_1[17]), .E(n987), .CK(clk), .Q(R5[17]) );
  EDFFX1 R5_reg_16_ ( .D(data_in_1[16]), .E(n987), .CK(clk), .Q(R5[16]) );
  EDFFX1 R5_reg_15_ ( .D(data_in_1[15]), .E(n987), .CK(clk), .Q(R5[15]) );
  EDFFX1 R5_reg_14_ ( .D(data_in_1[14]), .E(n987), .CK(clk), .Q(R5[14]) );
  EDFFX1 R5_reg_13_ ( .D(data_in_1[13]), .E(n987), .CK(clk), .Q(R5[13]) );
  EDFFX1 R5_reg_12_ ( .D(data_in_1[12]), .E(n987), .CK(clk), .Q(R5[12]) );
  EDFFX1 R5_reg_11_ ( .D(data_in_1[11]), .E(n987), .CK(clk), .Q(R5[11]) );
  EDFFX1 R5_reg_10_ ( .D(data_in_1[10]), .E(n987), .CK(clk), .Q(R5[10]) );
  EDFFX1 R5_reg_9_ ( .D(data_in_1[9]), .E(n986), .CK(clk), .Q(R5[9]) );
  EDFFX1 R5_reg_8_ ( .D(data_in_1[8]), .E(n987), .CK(clk), .Q(R5[8]) );
  EDFFX1 R5_reg_7_ ( .D(data_in_1[7]), .E(n986), .CK(clk), .Q(R5[7]) );
  EDFFX1 R5_reg_6_ ( .D(data_in_1[6]), .E(n987), .CK(clk), .Q(R5[6]) );
  EDFFX1 R5_reg_5_ ( .D(data_in_1[5]), .E(n986), .CK(clk), .Q(R5[5]) );
  EDFFX1 R5_reg_4_ ( .D(data_in_1[4]), .E(n987), .CK(clk), .Q(R5[4]) );
  EDFFX1 R5_reg_3_ ( .D(data_in_1[3]), .E(n986), .CK(clk), .Q(R5[3]) );
  EDFFX1 R5_reg_2_ ( .D(data_in_1[2]), .E(n987), .CK(clk), .Q(R5[2]) );
  EDFFX1 R5_reg_1_ ( .D(data_in_1[1]), .E(n986), .CK(clk), .Q(R5[1]) );
  EDFFX1 R5_reg_0_ ( .D(data_in_1[0]), .E(n987), .CK(clk), .Q(R5[0]) );
  EDFFX1 R9_reg_33_ ( .D(data_in_1[33]), .E(n973), .CK(clk), .Q(R9[33]) );
  EDFFX1 R9_reg_32_ ( .D(data_in_1[32]), .E(n973), .CK(clk), .Q(R9[32]) );
  EDFFX1 R9_reg_31_ ( .D(data_in_1[31]), .E(n973), .CK(clk), .Q(R9[31]) );
  EDFFX1 R9_reg_30_ ( .D(data_in_1[30]), .E(n973), .CK(clk), .Q(R9[30]) );
  EDFFX1 R9_reg_29_ ( .D(data_in_1[29]), .E(n973), .CK(clk), .Q(R9[29]) );
  EDFFX1 R9_reg_28_ ( .D(data_in_1[28]), .E(n973), .CK(clk), .Q(R9[28]) );
  EDFFX1 R9_reg_27_ ( .D(data_in_1[27]), .E(n973), .CK(clk), .Q(R9[27]) );
  EDFFX1 R9_reg_26_ ( .D(data_in_1[26]), .E(n973), .CK(clk), .Q(R9[26]) );
  EDFFX1 R9_reg_25_ ( .D(data_in_1[25]), .E(n996), .CK(clk), .Q(R9[25]) );
  EDFFX1 R9_reg_24_ ( .D(data_in_1[24]), .E(n995), .CK(clk), .Q(R9[24]) );
  EDFFX1 R9_reg_23_ ( .D(data_in_1[23]), .E(n996), .CK(clk), .Q(R9[23]) );
  EDFFX1 R9_reg_22_ ( .D(data_in_1[22]), .E(n996), .CK(clk), .Q(R9[22]) );
  EDFFX1 R9_reg_21_ ( .D(data_in_1[21]), .E(n995), .CK(clk), .Q(R9[21]) );
  EDFFX1 R9_reg_20_ ( .D(data_in_1[20]), .E(n995), .CK(clk), .Q(R9[20]) );
  EDFFX1 R9_reg_19_ ( .D(data_in_1[19]), .E(n995), .CK(clk), .Q(R9[19]) );
  EDFFX1 R9_reg_18_ ( .D(data_in_1[18]), .E(n995), .CK(clk), .Q(R9[18]) );
  EDFFX1 R9_reg_17_ ( .D(data_in_1[17]), .E(n995), .CK(clk), .Q(R9[17]) );
  EDFFX1 R9_reg_16_ ( .D(data_in_1[16]), .E(n995), .CK(clk), .Q(R9[16]) );
  EDFFX1 R9_reg_15_ ( .D(data_in_1[15]), .E(n995), .CK(clk), .Q(R9[15]) );
  EDFFX1 R9_reg_14_ ( .D(data_in_1[14]), .E(n995), .CK(clk), .Q(R9[14]) );
  EDFFX1 R9_reg_13_ ( .D(data_in_1[13]), .E(n995), .CK(clk), .Q(R9[13]) );
  EDFFX1 R9_reg_12_ ( .D(data_in_1[12]), .E(n995), .CK(clk), .Q(R9[12]) );
  EDFFX1 R9_reg_11_ ( .D(data_in_1[11]), .E(n995), .CK(clk), .Q(R9[11]) );
  EDFFX1 R9_reg_10_ ( .D(data_in_1[10]), .E(n995), .CK(clk), .Q(R9[10]) );
  EDFFX1 R9_reg_9_ ( .D(data_in_1[9]), .E(n996), .CK(clk), .Q(R9[9]) );
  EDFFX1 R9_reg_8_ ( .D(data_in_1[8]), .E(n996), .CK(clk), .Q(R9[8]) );
  EDFFX1 R9_reg_7_ ( .D(data_in_1[7]), .E(n996), .CK(clk), .Q(R9[7]) );
  EDFFX1 R9_reg_6_ ( .D(data_in_1[6]), .E(n996), .CK(clk), .Q(R9[6]) );
  EDFFX1 R9_reg_5_ ( .D(data_in_1[5]), .E(n996), .CK(clk), .Q(R9[5]) );
  EDFFX1 R9_reg_4_ ( .D(data_in_1[4]), .E(n996), .CK(clk), .Q(R9[4]) );
  EDFFX1 R9_reg_3_ ( .D(data_in_1[3]), .E(n996), .CK(clk), .Q(R9[3]) );
  EDFFX1 R9_reg_2_ ( .D(data_in_1[2]), .E(n996), .CK(clk), .Q(R9[2]) );
  EDFFX1 R9_reg_1_ ( .D(data_in_1[1]), .E(n996), .CK(clk), .Q(R9[1]) );
  EDFFX1 R9_reg_0_ ( .D(data_in_1[0]), .E(n996), .CK(clk), .Q(R9[0]) );
  EDFFX1 R14_reg_33_ ( .D(data_in_1[33]), .E(n1015), .CK(clk), .Q(R14[33]) );
  EDFFX1 R14_reg_32_ ( .D(data_in_1[32]), .E(n1015), .CK(clk), .Q(R14[32]) );
  EDFFX1 R14_reg_31_ ( .D(data_in_1[31]), .E(n1015), .CK(clk), .Q(R14[31]) );
  EDFFX1 R14_reg_30_ ( .D(data_in_1[30]), .E(n1015), .CK(clk), .Q(R14[30]) );
  EDFFX1 R14_reg_29_ ( .D(data_in_1[29]), .E(n1015), .CK(clk), .Q(R14[29]) );
  EDFFX1 R14_reg_28_ ( .D(data_in_1[28]), .E(n1015), .CK(clk), .Q(R14[28]) );
  EDFFX1 R14_reg_27_ ( .D(data_in_1[27]), .E(n1015), .CK(clk), .Q(R14[27]) );
  EDFFX1 R14_reg_26_ ( .D(data_in_1[26]), .E(n1015), .CK(clk), .Q(R14[26]) );
  EDFFX1 R14_reg_25_ ( .D(data_in_1[25]), .E(n968), .CK(clk), .Q(R14[25]) );
  EDFFX1 R14_reg_24_ ( .D(data_in_1[24]), .E(n1014), .CK(clk), .Q(R14[24]) );
  EDFFX1 R14_reg_23_ ( .D(data_in_1[23]), .E(n1015), .CK(clk), .Q(R14[23]) );
  EDFFX1 R14_reg_22_ ( .D(data_in_1[22]), .E(n1015), .CK(clk), .Q(R14[22]) );
  EDFFX1 R14_reg_21_ ( .D(data_in_1[21]), .E(n968), .CK(clk), .Q(R14[21]) );
  EDFFX1 R14_reg_20_ ( .D(data_in_1[20]), .E(n1014), .CK(clk), .Q(R14[20]) );
  EDFFX1 R14_reg_19_ ( .D(data_in_1[19]), .E(n1015), .CK(clk), .Q(R14[19]) );
  EDFFX1 R14_reg_18_ ( .D(data_in_1[18]), .E(n1012), .CK(clk), .Q(R14[18]) );
  EDFFX1 R14_reg_17_ ( .D(data_in_1[17]), .E(n968), .CK(clk), .Q(R14[17]) );
  EDFFX1 R14_reg_16_ ( .D(data_in_1[16]), .E(n1014), .CK(clk), .Q(R14[16]) );
  EDFFX1 R14_reg_15_ ( .D(data_in_1[15]), .E(n1015), .CK(clk), .Q(R14[15]) );
  EDFFX1 R14_reg_14_ ( .D(data_in_1[14]), .E(n1014), .CK(clk), .Q(R14[14]) );
  EDFFX1 R14_reg_13_ ( .D(data_in_1[13]), .E(n968), .CK(clk), .Q(R14[13]) );
  EDFFX1 R14_reg_12_ ( .D(data_in_1[12]), .E(n1014), .CK(clk), .Q(R14[12]) );
  EDFFX1 R14_reg_11_ ( .D(data_in_1[11]), .E(n1015), .CK(clk), .Q(R14[11]) );
  EDFFX1 R14_reg_10_ ( .D(data_in_1[10]), .E(n1015), .CK(clk), .Q(R14[10]) );
  EDFFX1 R14_reg_9_ ( .D(data_in_1[9]), .E(n968), .CK(clk), .Q(R14[9]) );
  EDFFX1 R14_reg_8_ ( .D(data_in_1[8]), .E(n1014), .CK(clk), .Q(R14[8]) );
  EDFFX1 R14_reg_7_ ( .D(data_in_1[7]), .E(n1015), .CK(clk), .Q(R14[7]) );
  EDFFX1 R14_reg_6_ ( .D(data_in_1[6]), .E(n1012), .CK(clk), .Q(R14[6]) );
  EDFFX1 R14_reg_5_ ( .D(data_in_1[5]), .E(n968), .CK(clk), .Q(R14[5]) );
  EDFFX1 R14_reg_4_ ( .D(data_in_1[4]), .E(n1014), .CK(clk), .Q(R14[4]) );
  EDFFX1 R14_reg_3_ ( .D(data_in_1[3]), .E(n1013), .CK(clk), .Q(R14[3]) );
  EDFFX1 R14_reg_2_ ( .D(data_in_1[2]), .E(n1015), .CK(clk), .Q(R14[2]) );
  EDFFX1 R14_reg_1_ ( .D(data_in_1[1]), .E(n1013), .CK(clk), .Q(R14[1]) );
  EDFFX1 R14_reg_0_ ( .D(data_in_1[0]), .E(n1013), .CK(clk), .Q(R14[0]) );
  EDFFX1 R2_reg_33_ ( .D(data_in_1[33]), .E(n980), .CK(clk), .Q(R2[33]) );
  EDFFX1 R2_reg_32_ ( .D(data_in_1[32]), .E(n980), .CK(clk), .Q(R2[32]) );
  EDFFX1 R2_reg_31_ ( .D(data_in_1[31]), .E(n980), .CK(clk), .Q(R2[31]) );
  EDFFX1 R2_reg_30_ ( .D(data_in_1[30]), .E(n980), .CK(clk), .Q(R2[30]) );
  EDFFX1 R2_reg_29_ ( .D(data_in_1[29]), .E(n980), .CK(clk), .Q(R2[29]) );
  EDFFX1 R2_reg_28_ ( .D(data_in_1[28]), .E(n980), .CK(clk), .Q(R2[28]) );
  EDFFX1 R2_reg_27_ ( .D(data_in_1[27]), .E(n980), .CK(clk), .Q(R2[27]) );
  EDFFX1 R2_reg_26_ ( .D(data_in_1[26]), .E(n980), .CK(clk), .Q(R2[26]) );
  EDFFX1 R2_reg_25_ ( .D(data_in_1[25]), .E(n980), .CK(clk), .Q(R2[25]) );
  EDFFX1 R2_reg_24_ ( .D(data_in_1[24]), .E(n980), .CK(clk), .Q(R2[24]) );
  EDFFX1 R2_reg_23_ ( .D(data_in_1[23]), .E(n980), .CK(clk), .Q(R2[23]) );
  EDFFX1 R2_reg_22_ ( .D(data_in_1[22]), .E(n980), .CK(clk), .Q(R2[22]) );
  EDFFX1 R2_reg_21_ ( .D(data_in_1[21]), .E(n981), .CK(clk), .Q(R2[21]) );
  EDFFX1 R2_reg_20_ ( .D(data_in_1[20]), .E(n981), .CK(clk), .Q(R2[20]) );
  EDFFX1 R2_reg_19_ ( .D(data_in_1[19]), .E(n981), .CK(clk), .Q(R2[19]) );
  EDFFX1 R2_reg_18_ ( .D(data_in_1[18]), .E(n981), .CK(clk), .Q(R2[18]) );
  EDFFX1 R2_reg_17_ ( .D(data_in_1[17]), .E(n981), .CK(clk), .Q(R2[17]) );
  EDFFX1 R2_reg_16_ ( .D(data_in_1[16]), .E(n981), .CK(clk), .Q(R2[16]) );
  EDFFX1 R2_reg_15_ ( .D(data_in_1[15]), .E(n981), .CK(clk), .Q(R2[15]) );
  EDFFX1 R2_reg_14_ ( .D(data_in_1[14]), .E(n981), .CK(clk), .Q(R2[14]) );
  EDFFX1 R2_reg_13_ ( .D(data_in_1[13]), .E(n981), .CK(clk), .Q(R2[13]) );
  EDFFX1 R2_reg_12_ ( .D(data_in_1[12]), .E(n981), .CK(clk), .Q(R2[12]) );
  EDFFX1 R2_reg_11_ ( .D(data_in_1[11]), .E(n981), .CK(clk), .Q(R2[11]) );
  EDFFX1 R2_reg_10_ ( .D(data_in_1[10]), .E(n981), .CK(clk), .Q(R2[10]) );
  EDFFX1 R2_reg_9_ ( .D(data_in_1[9]), .E(n980), .CK(clk), .Q(R2[9]) );
  EDFFX1 R2_reg_8_ ( .D(data_in_1[8]), .E(n981), .CK(clk), .Q(R2[8]) );
  EDFFX1 R2_reg_7_ ( .D(data_in_1[7]), .E(n980), .CK(clk), .Q(R2[7]) );
  EDFFX1 R2_reg_6_ ( .D(data_in_1[6]), .E(n981), .CK(clk), .Q(R2[6]) );
  EDFFX1 R2_reg_5_ ( .D(data_in_1[5]), .E(n980), .CK(clk), .Q(R2[5]) );
  EDFFX1 R2_reg_4_ ( .D(data_in_1[4]), .E(n981), .CK(clk), .Q(R2[4]) );
  EDFFX1 R2_reg_3_ ( .D(data_in_1[3]), .E(n980), .CK(clk), .Q(R2[3]) );
  EDFFX1 R2_reg_2_ ( .D(data_in_1[2]), .E(n981), .CK(clk), .Q(R2[2]) );
  EDFFX1 R2_reg_1_ ( .D(data_in_1[1]), .E(n980), .CK(clk), .Q(R2[1]) );
  EDFFX1 R2_reg_0_ ( .D(data_in_1[0]), .E(n981), .CK(clk), .Q(R2[0]) );
  EDFFX1 R6_reg_33_ ( .D(data_in_1[33]), .E(n988), .CK(clk), .Q(R6[33]) );
  EDFFX1 R6_reg_32_ ( .D(data_in_1[32]), .E(n988), .CK(clk), .Q(R6[32]) );
  EDFFX1 R6_reg_31_ ( .D(data_in_1[31]), .E(n988), .CK(clk), .Q(R6[31]) );
  EDFFX1 R6_reg_30_ ( .D(data_in_1[30]), .E(n988), .CK(clk), .Q(R6[30]) );
  EDFFX1 R6_reg_29_ ( .D(data_in_1[29]), .E(n988), .CK(clk), .Q(R6[29]) );
  EDFFX1 R6_reg_28_ ( .D(data_in_1[28]), .E(n988), .CK(clk), .Q(R6[28]) );
  EDFFX1 R6_reg_27_ ( .D(data_in_1[27]), .E(n988), .CK(clk), .Q(R6[27]) );
  EDFFX1 R6_reg_26_ ( .D(data_in_1[26]), .E(n988), .CK(clk), .Q(R6[26]) );
  EDFFX1 R6_reg_25_ ( .D(data_in_1[25]), .E(n988), .CK(clk), .Q(R6[25]) );
  EDFFX1 R6_reg_24_ ( .D(data_in_1[24]), .E(n988), .CK(clk), .Q(R6[24]) );
  EDFFX1 R6_reg_23_ ( .D(data_in_1[23]), .E(n988), .CK(clk), .Q(R6[23]) );
  EDFFX1 R6_reg_22_ ( .D(data_in_1[22]), .E(n988), .CK(clk), .Q(R6[22]) );
  EDFFX1 R6_reg_21_ ( .D(data_in_1[21]), .E(n989), .CK(clk), .Q(R6[21]) );
  EDFFX1 R6_reg_20_ ( .D(data_in_1[20]), .E(n989), .CK(clk), .Q(R6[20]) );
  EDFFX1 R6_reg_19_ ( .D(data_in_1[19]), .E(n989), .CK(clk), .Q(R6[19]) );
  EDFFX1 R6_reg_18_ ( .D(data_in_1[18]), .E(n989), .CK(clk), .Q(R6[18]) );
  EDFFX1 R6_reg_17_ ( .D(data_in_1[17]), .E(n989), .CK(clk), .Q(R6[17]) );
  EDFFX1 R6_reg_16_ ( .D(data_in_1[16]), .E(n989), .CK(clk), .Q(R6[16]) );
  EDFFX1 R6_reg_15_ ( .D(data_in_1[15]), .E(n989), .CK(clk), .Q(R6[15]) );
  EDFFX1 R6_reg_14_ ( .D(data_in_1[14]), .E(n989), .CK(clk), .Q(R6[14]) );
  EDFFX1 R6_reg_13_ ( .D(data_in_1[13]), .E(n989), .CK(clk), .Q(R6[13]) );
  EDFFX1 R6_reg_12_ ( .D(data_in_1[12]), .E(n989), .CK(clk), .Q(R6[12]) );
  EDFFX1 R6_reg_11_ ( .D(data_in_1[11]), .E(n989), .CK(clk), .Q(R6[11]) );
  EDFFX1 R6_reg_10_ ( .D(data_in_1[10]), .E(n989), .CK(clk), .Q(R6[10]) );
  EDFFX1 R6_reg_9_ ( .D(data_in_1[9]), .E(n988), .CK(clk), .Q(R6[9]) );
  EDFFX1 R6_reg_8_ ( .D(data_in_1[8]), .E(n989), .CK(clk), .Q(R6[8]) );
  EDFFX1 R6_reg_7_ ( .D(data_in_1[7]), .E(n988), .CK(clk), .Q(R6[7]) );
  EDFFX1 R6_reg_6_ ( .D(data_in_1[6]), .E(n989), .CK(clk), .Q(R6[6]) );
  EDFFX1 R6_reg_5_ ( .D(data_in_1[5]), .E(n988), .CK(clk), .Q(R6[5]) );
  EDFFX1 R6_reg_4_ ( .D(data_in_1[4]), .E(n989), .CK(clk), .Q(R6[4]) );
  EDFFX1 R6_reg_3_ ( .D(data_in_1[3]), .E(n988), .CK(clk), .Q(R6[3]) );
  EDFFX1 R6_reg_2_ ( .D(data_in_1[2]), .E(n989), .CK(clk), .Q(R6[2]) );
  EDFFX1 R6_reg_1_ ( .D(data_in_1[1]), .E(n988), .CK(clk), .Q(R6[1]) );
  EDFFX1 R6_reg_0_ ( .D(data_in_1[0]), .E(n989), .CK(clk), .Q(R6[0]) );
  EDFFX1 R10_reg_33_ ( .D(data_in_1[33]), .E(n972), .CK(clk), .Q(R10[33]) );
  EDFFX1 R10_reg_32_ ( .D(data_in_1[32]), .E(n972), .CK(clk), .Q(R10[32]) );
  EDFFX1 R10_reg_31_ ( .D(data_in_1[31]), .E(n972), .CK(clk), .Q(R10[31]) );
  EDFFX1 R10_reg_30_ ( .D(data_in_1[30]), .E(n972), .CK(clk), .Q(R10[30]) );
  EDFFX1 R10_reg_29_ ( .D(data_in_1[29]), .E(n972), .CK(clk), .Q(R10[29]) );
  EDFFX1 R10_reg_28_ ( .D(data_in_1[28]), .E(n972), .CK(clk), .Q(R10[28]) );
  EDFFX1 R10_reg_27_ ( .D(data_in_1[27]), .E(n972), .CK(clk), .Q(R10[27]) );
  EDFFX1 R10_reg_26_ ( .D(data_in_1[26]), .E(n972), .CK(clk), .Q(R10[26]) );
  EDFFX1 R10_reg_25_ ( .D(data_in_1[25]), .E(n999), .CK(clk), .Q(R10[25]) );
  EDFFX1 R10_reg_24_ ( .D(data_in_1[24]), .E(n998), .CK(clk), .Q(R10[24]) );
  EDFFX1 R10_reg_23_ ( .D(data_in_1[23]), .E(n999), .CK(clk), .Q(R10[23]) );
  EDFFX1 R10_reg_22_ ( .D(data_in_1[22]), .E(n999), .CK(clk), .Q(R10[22]) );
  EDFFX1 R10_reg_21_ ( .D(data_in_1[21]), .E(n998), .CK(clk), .Q(R10[21]) );
  EDFFX1 R10_reg_20_ ( .D(data_in_1[20]), .E(n998), .CK(clk), .Q(R10[20]) );
  EDFFX1 R10_reg_19_ ( .D(data_in_1[19]), .E(n998), .CK(clk), .Q(R10[19]) );
  EDFFX1 R10_reg_18_ ( .D(data_in_1[18]), .E(n998), .CK(clk), .Q(R10[18]) );
  EDFFX1 R10_reg_17_ ( .D(data_in_1[17]), .E(n998), .CK(clk), .Q(R10[17]) );
  EDFFX1 R10_reg_16_ ( .D(data_in_1[16]), .E(n998), .CK(clk), .Q(R10[16]) );
  EDFFX1 R10_reg_15_ ( .D(data_in_1[15]), .E(n998), .CK(clk), .Q(R10[15]) );
  EDFFX1 R10_reg_14_ ( .D(data_in_1[14]), .E(n998), .CK(clk), .Q(R10[14]) );
  EDFFX1 R10_reg_13_ ( .D(data_in_1[13]), .E(n998), .CK(clk), .Q(R10[13]) );
  EDFFX1 R10_reg_12_ ( .D(data_in_1[12]), .E(n998), .CK(clk), .Q(R10[12]) );
  EDFFX1 R10_reg_11_ ( .D(data_in_1[11]), .E(n998), .CK(clk), .Q(R10[11]) );
  EDFFX1 R10_reg_10_ ( .D(data_in_1[10]), .E(n998), .CK(clk), .Q(R10[10]) );
  EDFFX1 R10_reg_9_ ( .D(data_in_1[9]), .E(n999), .CK(clk), .Q(R10[9]) );
  EDFFX1 R10_reg_8_ ( .D(data_in_1[8]), .E(n999), .CK(clk), .Q(R10[8]) );
  EDFFX1 R10_reg_7_ ( .D(data_in_1[7]), .E(n999), .CK(clk), .Q(R10[7]) );
  EDFFX1 R10_reg_6_ ( .D(data_in_1[6]), .E(n999), .CK(clk), .Q(R10[6]) );
  EDFFX1 R10_reg_5_ ( .D(data_in_1[5]), .E(n999), .CK(clk), .Q(R10[5]) );
  EDFFX1 R10_reg_4_ ( .D(data_in_1[4]), .E(n999), .CK(clk), .Q(R10[4]) );
  EDFFX1 R10_reg_3_ ( .D(data_in_1[3]), .E(n999), .CK(clk), .Q(R10[3]) );
  EDFFX1 R10_reg_2_ ( .D(data_in_1[2]), .E(n999), .CK(clk), .Q(R10[2]) );
  EDFFX1 R10_reg_1_ ( .D(data_in_1[1]), .E(n999), .CK(clk), .Q(R10[1]) );
  EDFFX1 R10_reg_0_ ( .D(data_in_1[0]), .E(n999), .CK(clk), .Q(R10[0]) );
  EDFFX1 R0_reg_33_ ( .D(data_in_1[33]), .E(n1039), .CK(clk), .Q(R0[33]) );
  EDFFX1 R0_reg_32_ ( .D(data_in_1[32]), .E(n1039), .CK(clk), .Q(R0[32]) );
  EDFFX1 R0_reg_31_ ( .D(data_in_1[31]), .E(n1039), .CK(clk), .Q(R0[31]) );
  EDFFX1 R0_reg_30_ ( .D(data_in_1[30]), .E(n1039), .CK(clk), .Q(R0[30]) );
  EDFFX1 R0_reg_29_ ( .D(data_in_1[29]), .E(n1039), .CK(clk), .Q(R0[29]) );
  EDFFX1 R0_reg_28_ ( .D(data_in_1[28]), .E(n1039), .CK(clk), .Q(R0[28]) );
  EDFFX1 R0_reg_27_ ( .D(data_in_1[27]), .E(n1039), .CK(clk), .Q(R0[27]) );
  EDFFX1 R0_reg_26_ ( .D(data_in_1[26]), .E(n1039), .CK(clk), .Q(R0[26]) );
  EDFFX1 R0_reg_25_ ( .D(data_in_1[25]), .E(n1039), .CK(clk), .Q(R0[25]) );
  EDFFX1 R0_reg_24_ ( .D(data_in_1[24]), .E(n1039), .CK(clk), .Q(R0[24]) );
  EDFFX1 R0_reg_23_ ( .D(data_in_1[23]), .E(n1031), .CK(clk), .Q(R0[23]) );
  EDFFX1 R0_reg_22_ ( .D(data_in_1[22]), .E(n1038), .CK(clk), .Q(R0[22]) );
  EDFFX1 R0_reg_21_ ( .D(data_in_1[21]), .E(n1033), .CK(clk), .Q(R0[21]) );
  EDFFX1 R0_reg_20_ ( .D(data_in_1[20]), .E(n1036), .CK(clk), .Q(R0[20]) );
  EDFFX1 R0_reg_19_ ( .D(data_in_1[19]), .E(n1030), .CK(clk), .Q(R0[19]) );
  EDFFX1 R0_reg_18_ ( .D(data_in_1[18]), .E(n1037), .CK(clk), .Q(R0[18]) );
  EDFFX1 R0_reg_17_ ( .D(data_in_1[17]), .E(n1035), .CK(clk), .Q(R0[17]) );
  EDFFX1 R0_reg_16_ ( .D(data_in_1[16]), .E(n1032), .CK(clk), .Q(R0[16]) );
  EDFFX1 R0_reg_15_ ( .D(data_in_1[15]), .E(n1034), .CK(clk), .Q(R0[15]) );
  EDFFX1 R0_reg_14_ ( .D(data_in_1[14]), .E(n1031), .CK(clk), .Q(R0[14]) );
  EDFFX1 R0_reg_13_ ( .D(data_in_1[13]), .E(n1038), .CK(clk), .Q(R0[13]) );
  EDFFX1 R0_reg_12_ ( .D(data_in_1[12]), .E(n1033), .CK(clk), .Q(R0[12]) );
  EDFFX1 R0_reg_11_ ( .D(data_in_1[11]), .E(n1036), .CK(clk), .Q(R0[11]) );
  EDFFX1 R0_reg_10_ ( .D(data_in_1[10]), .E(n1030), .CK(clk), .Q(R0[10]) );
  EDFFX1 R0_reg_9_ ( .D(data_in_1[9]), .E(n1037), .CK(clk), .Q(R0[9]) );
  EDFFX1 R0_reg_8_ ( .D(data_in_1[8]), .E(n1035), .CK(clk), .Q(R0[8]) );
  EDFFX1 R0_reg_7_ ( .D(data_in_1[7]), .E(n1032), .CK(clk), .Q(R0[7]) );
  EDFFX1 R0_reg_6_ ( .D(data_in_1[6]), .E(n1034), .CK(clk), .Q(R0[6]) );
  EDFFX1 R0_reg_5_ ( .D(data_in_1[5]), .E(n1031), .CK(clk), .Q(R0[5]) );
  EDFFX1 R0_reg_4_ ( .D(data_in_1[4]), .E(n1038), .CK(clk), .Q(R0[4]) );
  EDFFX1 R0_reg_3_ ( .D(data_in_1[3]), .E(n1033), .CK(clk), .Q(R0[3]) );
  EDFFX1 R0_reg_2_ ( .D(data_in_1[2]), .E(n1036), .CK(clk), .Q(R0[2]) );
  EDFFX1 R0_reg_1_ ( .D(data_in_1[1]), .E(n1033), .CK(clk), .Q(R0[1]) );
  EDFFX1 R0_reg_0_ ( .D(data_in_1[0]), .E(n1036), .CK(clk), .Q(R0[0]) );
  EDFFX1 R4_reg_33_ ( .D(data_in_1[33]), .E(n984), .CK(clk), .Q(R4[33]) );
  EDFFX1 R4_reg_32_ ( .D(data_in_1[32]), .E(n984), .CK(clk), .Q(R4[32]) );
  EDFFX1 R4_reg_31_ ( .D(data_in_1[31]), .E(n984), .CK(clk), .Q(R4[31]) );
  EDFFX1 R4_reg_30_ ( .D(data_in_1[30]), .E(n984), .CK(clk), .Q(R4[30]) );
  EDFFX1 R4_reg_29_ ( .D(data_in_1[29]), .E(n984), .CK(clk), .Q(R4[29]) );
  EDFFX1 R4_reg_28_ ( .D(data_in_1[28]), .E(n984), .CK(clk), .Q(R4[28]) );
  EDFFX1 R4_reg_27_ ( .D(data_in_1[27]), .E(n984), .CK(clk), .Q(R4[27]) );
  EDFFX1 R4_reg_26_ ( .D(data_in_1[26]), .E(n984), .CK(clk), .Q(R4[26]) );
  EDFFX1 R4_reg_25_ ( .D(data_in_1[25]), .E(n984), .CK(clk), .Q(R4[25]) );
  EDFFX1 R4_reg_24_ ( .D(data_in_1[24]), .E(n984), .CK(clk), .Q(R4[24]) );
  EDFFX1 R4_reg_23_ ( .D(data_in_1[23]), .E(n984), .CK(clk), .Q(R4[23]) );
  EDFFX1 R4_reg_22_ ( .D(data_in_1[22]), .E(n984), .CK(clk), .Q(R4[22]) );
  EDFFX1 R4_reg_21_ ( .D(data_in_1[21]), .E(n985), .CK(clk), .Q(R4[21]) );
  EDFFX1 R4_reg_20_ ( .D(data_in_1[20]), .E(n985), .CK(clk), .Q(R4[20]) );
  EDFFX1 R4_reg_19_ ( .D(data_in_1[19]), .E(n985), .CK(clk), .Q(R4[19]) );
  EDFFX1 R4_reg_18_ ( .D(data_in_1[18]), .E(n985), .CK(clk), .Q(R4[18]) );
  EDFFX1 R4_reg_17_ ( .D(data_in_1[17]), .E(n985), .CK(clk), .Q(R4[17]) );
  EDFFX1 R4_reg_16_ ( .D(data_in_1[16]), .E(n985), .CK(clk), .Q(R4[16]) );
  EDFFX1 R4_reg_15_ ( .D(data_in_1[15]), .E(n985), .CK(clk), .Q(R4[15]) );
  EDFFX1 R4_reg_14_ ( .D(data_in_1[14]), .E(n985), .CK(clk), .Q(R4[14]) );
  EDFFX1 R4_reg_13_ ( .D(data_in_1[13]), .E(n985), .CK(clk), .Q(R4[13]) );
  EDFFX1 R4_reg_12_ ( .D(data_in_1[12]), .E(n985), .CK(clk), .Q(R4[12]) );
  EDFFX1 R4_reg_11_ ( .D(data_in_1[11]), .E(n985), .CK(clk), .Q(R4[11]) );
  EDFFX1 R4_reg_10_ ( .D(data_in_1[10]), .E(n985), .CK(clk), .Q(R4[10]) );
  EDFFX1 R4_reg_9_ ( .D(data_in_1[9]), .E(n984), .CK(clk), .Q(R4[9]) );
  EDFFX1 R4_reg_8_ ( .D(data_in_1[8]), .E(n985), .CK(clk), .Q(R4[8]) );
  EDFFX1 R4_reg_7_ ( .D(data_in_1[7]), .E(n984), .CK(clk), .Q(R4[7]) );
  EDFFX1 R4_reg_6_ ( .D(data_in_1[6]), .E(n985), .CK(clk), .Q(R4[6]) );
  EDFFX1 R4_reg_5_ ( .D(data_in_1[5]), .E(n984), .CK(clk), .Q(R4[5]) );
  EDFFX1 R4_reg_4_ ( .D(data_in_1[4]), .E(n985), .CK(clk), .Q(R4[4]) );
  EDFFX1 R4_reg_3_ ( .D(data_in_1[3]), .E(n984), .CK(clk), .Q(R4[3]) );
  EDFFX1 R4_reg_2_ ( .D(data_in_1[2]), .E(n985), .CK(clk), .Q(R4[2]) );
  EDFFX1 R4_reg_1_ ( .D(data_in_1[1]), .E(n984), .CK(clk), .Q(R4[1]) );
  EDFFX1 R4_reg_0_ ( .D(data_in_1[0]), .E(n985), .CK(clk), .Q(R4[0]) );
  EDFFX1 R8_reg_33_ ( .D(data_in_1[33]), .E(n974), .CK(clk), .Q(R8[33]) );
  EDFFX1 R8_reg_32_ ( .D(data_in_1[32]), .E(n974), .CK(clk), .Q(R8[32]) );
  EDFFX1 R8_reg_31_ ( .D(data_in_1[31]), .E(n974), .CK(clk), .Q(R8[31]) );
  EDFFX1 R8_reg_30_ ( .D(data_in_1[30]), .E(n974), .CK(clk), .Q(R8[30]) );
  EDFFX1 R8_reg_29_ ( .D(data_in_1[29]), .E(n974), .CK(clk), .Q(R8[29]) );
  EDFFX1 R8_reg_28_ ( .D(data_in_1[28]), .E(n974), .CK(clk), .Q(R8[28]) );
  EDFFX1 R8_reg_27_ ( .D(data_in_1[27]), .E(n974), .CK(clk), .Q(R8[27]) );
  EDFFX1 R8_reg_26_ ( .D(data_in_1[26]), .E(n974), .CK(clk), .Q(R8[26]) );
  EDFFX1 R8_reg_25_ ( .D(data_in_1[25]), .E(n993), .CK(clk), .Q(R8[25]) );
  EDFFX1 R8_reg_24_ ( .D(data_in_1[24]), .E(n992), .CK(clk), .Q(R8[24]) );
  EDFFX1 R8_reg_23_ ( .D(data_in_1[23]), .E(n993), .CK(clk), .Q(R8[23]) );
  EDFFX1 R8_reg_22_ ( .D(data_in_1[22]), .E(n993), .CK(clk), .Q(R8[22]) );
  EDFFX1 R8_reg_21_ ( .D(data_in_1[21]), .E(n992), .CK(clk), .Q(R8[21]) );
  EDFFX1 R8_reg_20_ ( .D(data_in_1[20]), .E(n992), .CK(clk), .Q(R8[20]) );
  EDFFX1 R8_reg_19_ ( .D(data_in_1[19]), .E(n992), .CK(clk), .Q(R8[19]) );
  EDFFX1 R8_reg_18_ ( .D(data_in_1[18]), .E(n992), .CK(clk), .Q(R8[18]) );
  EDFFX1 R8_reg_17_ ( .D(data_in_1[17]), .E(n992), .CK(clk), .Q(R8[17]) );
  EDFFX1 R8_reg_16_ ( .D(data_in_1[16]), .E(n992), .CK(clk), .Q(R8[16]) );
  EDFFX1 R8_reg_15_ ( .D(data_in_1[15]), .E(n992), .CK(clk), .Q(R8[15]) );
  EDFFX1 R8_reg_14_ ( .D(data_in_1[14]), .E(n992), .CK(clk), .Q(R8[14]) );
  EDFFX1 R8_reg_13_ ( .D(data_in_1[13]), .E(n992), .CK(clk), .Q(R8[13]) );
  EDFFX1 R8_reg_12_ ( .D(data_in_1[12]), .E(n992), .CK(clk), .Q(R8[12]) );
  EDFFX1 R8_reg_11_ ( .D(data_in_1[11]), .E(n992), .CK(clk), .Q(R8[11]) );
  EDFFX1 R8_reg_10_ ( .D(data_in_1[10]), .E(n992), .CK(clk), .Q(R8[10]) );
  EDFFX1 R8_reg_9_ ( .D(data_in_1[9]), .E(n993), .CK(clk), .Q(R8[9]) );
  EDFFX1 R8_reg_8_ ( .D(data_in_1[8]), .E(n993), .CK(clk), .Q(R8[8]) );
  EDFFX1 R8_reg_7_ ( .D(data_in_1[7]), .E(n993), .CK(clk), .Q(R8[7]) );
  EDFFX1 R8_reg_6_ ( .D(data_in_1[6]), .E(n993), .CK(clk), .Q(R8[6]) );
  EDFFX1 R8_reg_5_ ( .D(data_in_1[5]), .E(n993), .CK(clk), .Q(R8[5]) );
  EDFFX1 R8_reg_4_ ( .D(data_in_1[4]), .E(n993), .CK(clk), .Q(R8[4]) );
  EDFFX1 R8_reg_3_ ( .D(data_in_1[3]), .E(n993), .CK(clk), .Q(R8[3]) );
  EDFFX1 R8_reg_2_ ( .D(data_in_1[2]), .E(n993), .CK(clk), .Q(R8[2]) );
  EDFFX1 R8_reg_1_ ( .D(data_in_1[1]), .E(n993), .CK(clk), .Q(R8[1]) );
  EDFFX1 R8_reg_0_ ( .D(data_in_1[0]), .E(n993), .CK(clk), .Q(R8[0]) );
  EDFFX1 R12_reg_33_ ( .D(data_in_1[33]), .E(n1005), .CK(clk), .Q(R12[33]) );
  EDFFX1 R12_reg_32_ ( .D(data_in_1[32]), .E(n1005), .CK(clk), .Q(R12[32]) );
  EDFFX1 R12_reg_31_ ( .D(data_in_1[31]), .E(n1005), .CK(clk), .Q(R12[31]) );
  EDFFX1 R12_reg_30_ ( .D(data_in_1[30]), .E(n1005), .CK(clk), .Q(R12[30]) );
  EDFFX1 R12_reg_29_ ( .D(data_in_1[29]), .E(n1005), .CK(clk), .Q(R12[29]) );
  EDFFX1 R12_reg_28_ ( .D(data_in_1[28]), .E(n1005), .CK(clk), .Q(R12[28]) );
  EDFFX1 R12_reg_27_ ( .D(data_in_1[27]), .E(n1005), .CK(clk), .Q(R12[27]) );
  EDFFX1 R12_reg_26_ ( .D(data_in_1[26]), .E(n1005), .CK(clk), .Q(R12[26]) );
  EDFFX1 R12_reg_25_ ( .D(data_in_1[25]), .E(n1005), .CK(clk), .Q(R12[25]) );
  EDFFX1 R12_reg_24_ ( .D(data_in_1[24]), .E(n1005), .CK(clk), .Q(R12[24]) );
  EDFFX1 R12_reg_23_ ( .D(data_in_1[23]), .E(n1004), .CK(clk), .Q(R12[23]) );
  EDFFX1 R12_reg_22_ ( .D(data_in_1[22]), .E(n1004), .CK(clk), .Q(R12[22]) );
  EDFFX1 R12_reg_21_ ( .D(data_in_1[21]), .E(n1004), .CK(clk), .Q(R12[21]) );
  EDFFX1 R12_reg_20_ ( .D(data_in_1[20]), .E(n1004), .CK(clk), .Q(R12[20]) );
  EDFFX1 R12_reg_19_ ( .D(data_in_1[19]), .E(n1004), .CK(clk), .Q(R12[19]) );
  EDFFX1 R12_reg_18_ ( .D(data_in_1[18]), .E(n1004), .CK(clk), .Q(R12[18]) );
  EDFFX1 R12_reg_17_ ( .D(data_in_1[17]), .E(n1004), .CK(clk), .Q(R12[17]) );
  EDFFX1 R12_reg_16_ ( .D(data_in_1[16]), .E(n1004), .CK(clk), .Q(R12[16]) );
  EDFFX1 R12_reg_15_ ( .D(data_in_1[15]), .E(n1004), .CK(clk), .Q(R12[15]) );
  EDFFX1 R12_reg_14_ ( .D(data_in_1[14]), .E(n1004), .CK(clk), .Q(R12[14]) );
  EDFFX1 R12_reg_13_ ( .D(data_in_1[13]), .E(n1004), .CK(clk), .Q(R12[13]) );
  EDFFX1 R12_reg_12_ ( .D(data_in_1[12]), .E(n1004), .CK(clk), .Q(R12[12]) );
  EDFFX1 R12_reg_11_ ( .D(data_in_1[11]), .E(n970), .CK(clk), .Q(R12[11]) );
  EDFFX1 R12_reg_10_ ( .D(data_in_1[10]), .E(n970), .CK(clk), .Q(R12[10]) );
  EDFFX1 R12_reg_9_ ( .D(data_in_1[9]), .E(n970), .CK(clk), .Q(R12[9]) );
  EDFFX1 R12_reg_8_ ( .D(data_in_1[8]), .E(n970), .CK(clk), .Q(R12[8]) );
  EDFFX1 R12_reg_7_ ( .D(data_in_1[7]), .E(n970), .CK(clk), .Q(R12[7]) );
  EDFFX1 R12_reg_6_ ( .D(data_in_1[6]), .E(n970), .CK(clk), .Q(R12[6]) );
  EDFFX1 R12_reg_5_ ( .D(data_in_1[5]), .E(n970), .CK(clk), .Q(R12[5]) );
  EDFFX1 R12_reg_4_ ( .D(data_in_1[4]), .E(n1004), .CK(clk), .Q(R12[4]) );
  EDFFX1 R12_reg_3_ ( .D(data_in_1[3]), .E(n1005), .CK(clk), .Q(R12[3]) );
  EDFFX1 R12_reg_2_ ( .D(data_in_1[2]), .E(n1004), .CK(clk), .Q(R12[2]) );
  EDFFX1 R12_reg_1_ ( .D(data_in_1[1]), .E(n1005), .CK(clk), .Q(R12[1]) );
  EDFFX1 R12_reg_0_ ( .D(data_in_1[0]), .E(n1005), .CK(clk), .Q(R12[0]) );
  EDFFX1 R15_reg_33_ ( .D(data_in_1[33]), .E(n1028), .CK(clk), .Q(R15[33]) );
  EDFFX1 R15_reg_32_ ( .D(data_in_1[32]), .E(n1028), .CK(clk), .Q(R15[32]) );
  EDFFX1 R15_reg_31_ ( .D(data_in_1[31]), .E(n1028), .CK(clk), .Q(R15[31]) );
  EDFFX1 R15_reg_30_ ( .D(data_in_1[30]), .E(n1028), .CK(clk), .Q(R15[30]) );
  EDFFX1 R15_reg_29_ ( .D(data_in_1[29]), .E(n1028), .CK(clk), .Q(R15[29]) );
  EDFFX1 R15_reg_28_ ( .D(data_in_1[28]), .E(n1028), .CK(clk), .Q(R15[28]) );
  EDFFX1 R15_reg_27_ ( .D(data_in_1[27]), .E(n1028), .CK(clk), .Q(R15[27]) );
  EDFFX1 R15_reg_26_ ( .D(data_in_1[26]), .E(n1028), .CK(clk), .Q(R15[26]) );
  EDFFX1 R15_reg_25_ ( .D(data_in_1[25]), .E(n1028), .CK(clk), .Q(R15[25]) );
  EDFFX1 R15_reg_24_ ( .D(data_in_1[24]), .E(n1028), .CK(clk), .Q(R15[24]) );
  EDFFX1 R15_reg_23_ ( .D(data_in_1[23]), .E(n1028), .CK(clk), .Q(R15[23]) );
  EDFFX1 R15_reg_22_ ( .D(data_in_1[22]), .E(n1028), .CK(clk), .Q(R15[22]) );
  EDFFX1 R15_reg_21_ ( .D(data_in_1[21]), .E(n1028), .CK(clk), .Q(R15[21]) );
  EDFFX1 R15_reg_20_ ( .D(data_in_1[20]), .E(n1028), .CK(clk), .Q(R15[20]) );
  EDFFX1 R15_reg_19_ ( .D(data_in_1[19]), .E(n1028), .CK(clk), .Q(R15[19]) );
  EDFFX1 R15_reg_18_ ( .D(data_in_1[18]), .E(n1028), .CK(clk), .Q(R15[18]) );
  EDFFX1 R15_reg_17_ ( .D(data_in_1[17]), .E(n1028), .CK(clk), .Q(R15[17]) );
  EDFFX1 R15_reg_16_ ( .D(data_in_1[16]), .E(n1028), .CK(clk), .Q(R15[16]) );
  EDFFX1 R15_reg_15_ ( .D(data_in_1[15]), .E(n1028), .CK(clk), .Q(R15[15]) );
  EDFFX1 R15_reg_14_ ( .D(data_in_1[14]), .E(n1028), .CK(clk), .Q(R15[14]) );
  EDFFX1 R15_reg_13_ ( .D(data_in_1[13]), .E(n1028), .CK(clk), .Q(R15[13]) );
  EDFFX1 R15_reg_12_ ( .D(data_in_1[12]), .E(n1028), .CK(clk), .Q(R15[12]) );
  EDFFX1 R15_reg_11_ ( .D(data_in_1[11]), .E(n1028), .CK(clk), .Q(R15[11]) );
  EDFFX1 R15_reg_10_ ( .D(data_in_1[10]), .E(n1028), .CK(clk), .Q(R15[10]) );
  EDFFX1 R15_reg_9_ ( .D(data_in_1[9]), .E(n1028), .CK(clk), .Q(R15[9]) );
  EDFFX1 R15_reg_8_ ( .D(data_in_1[8]), .E(n1028), .CK(clk), .Q(R15[8]) );
  EDFFX1 R15_reg_7_ ( .D(data_in_1[7]), .E(n1028), .CK(clk), .Q(R15[7]) );
  EDFFX1 R15_reg_6_ ( .D(data_in_1[6]), .E(n1028), .CK(clk), .Q(R15[6]) );
  EDFFX1 R15_reg_5_ ( .D(data_in_1[5]), .E(n1028), .CK(clk), .Q(R15[5]) );
  EDFFX1 R15_reg_4_ ( .D(data_in_1[4]), .E(n1028), .CK(clk), .Q(R15[4]) );
  EDFFX1 R15_reg_3_ ( .D(data_in_1[3]), .E(n1028), .CK(clk), .Q(R15[3]) );
  EDFFX1 R15_reg_2_ ( .D(data_in_1[2]), .E(n1028), .CK(clk), .Q(R15[2]) );
  EDFFX1 R15_reg_1_ ( .D(data_in_1[1]), .E(n1028), .CK(clk), .Q(R15[1]) );
  EDFFX1 R15_reg_0_ ( .D(data_in_1[0]), .E(n1028), .CK(clk), .Q(R15[0]) );
  EDFFX1 R3_reg_33_ ( .D(data_in_1[33]), .E(n982), .CK(clk), .Q(R3[33]) );
  EDFFX1 R3_reg_32_ ( .D(data_in_1[32]), .E(n982), .CK(clk), .Q(R3[32]) );
  EDFFX1 R3_reg_31_ ( .D(data_in_1[31]), .E(n982), .CK(clk), .Q(R3[31]) );
  EDFFX1 R3_reg_30_ ( .D(data_in_1[30]), .E(n982), .CK(clk), .Q(R3[30]) );
  EDFFX1 R3_reg_29_ ( .D(data_in_1[29]), .E(n982), .CK(clk), .Q(R3[29]) );
  EDFFX1 R3_reg_28_ ( .D(data_in_1[28]), .E(n982), .CK(clk), .Q(R3[28]) );
  EDFFX1 R3_reg_27_ ( .D(data_in_1[27]), .E(n982), .CK(clk), .Q(R3[27]) );
  EDFFX1 R3_reg_26_ ( .D(data_in_1[26]), .E(n982), .CK(clk), .Q(R3[26]) );
  EDFFX1 R3_reg_25_ ( .D(data_in_1[25]), .E(n982), .CK(clk), .Q(R3[25]) );
  EDFFX1 R3_reg_24_ ( .D(data_in_1[24]), .E(n982), .CK(clk), .Q(R3[24]) );
  EDFFX1 R3_reg_23_ ( .D(data_in_1[23]), .E(n982), .CK(clk), .Q(R3[23]) );
  EDFFX1 R3_reg_22_ ( .D(data_in_1[22]), .E(n982), .CK(clk), .Q(R3[22]) );
  EDFFX1 R3_reg_21_ ( .D(data_in_1[21]), .E(n983), .CK(clk), .Q(R3[21]) );
  EDFFX1 R3_reg_20_ ( .D(data_in_1[20]), .E(n983), .CK(clk), .Q(R3[20]) );
  EDFFX1 R3_reg_19_ ( .D(data_in_1[19]), .E(n983), .CK(clk), .Q(R3[19]) );
  EDFFX1 R3_reg_18_ ( .D(data_in_1[18]), .E(n983), .CK(clk), .Q(R3[18]) );
  EDFFX1 R3_reg_17_ ( .D(data_in_1[17]), .E(n983), .CK(clk), .Q(R3[17]) );
  EDFFX1 R3_reg_16_ ( .D(data_in_1[16]), .E(n983), .CK(clk), .Q(R3[16]) );
  EDFFX1 R3_reg_15_ ( .D(data_in_1[15]), .E(n983), .CK(clk), .Q(R3[15]) );
  EDFFX1 R3_reg_14_ ( .D(data_in_1[14]), .E(n983), .CK(clk), .Q(R3[14]) );
  EDFFX1 R3_reg_13_ ( .D(data_in_1[13]), .E(n983), .CK(clk), .Q(R3[13]) );
  EDFFX1 R3_reg_12_ ( .D(data_in_1[12]), .E(n983), .CK(clk), .Q(R3[12]) );
  EDFFX1 R3_reg_11_ ( .D(data_in_1[11]), .E(n983), .CK(clk), .Q(R3[11]) );
  EDFFX1 R3_reg_10_ ( .D(data_in_1[10]), .E(n983), .CK(clk), .Q(R3[10]) );
  EDFFX1 R3_reg_9_ ( .D(data_in_1[9]), .E(n982), .CK(clk), .Q(R3[9]) );
  EDFFX1 R3_reg_8_ ( .D(data_in_1[8]), .E(n983), .CK(clk), .Q(R3[8]) );
  EDFFX1 R3_reg_7_ ( .D(data_in_1[7]), .E(n982), .CK(clk), .Q(R3[7]) );
  EDFFX1 R3_reg_6_ ( .D(data_in_1[6]), .E(n983), .CK(clk), .Q(R3[6]) );
  EDFFX1 R3_reg_5_ ( .D(data_in_1[5]), .E(n982), .CK(clk), .Q(R3[5]) );
  EDFFX1 R3_reg_4_ ( .D(data_in_1[4]), .E(n983), .CK(clk), .Q(R3[4]) );
  EDFFX1 R3_reg_3_ ( .D(data_in_1[3]), .E(n982), .CK(clk), .Q(R3[3]) );
  EDFFX1 R3_reg_2_ ( .D(data_in_1[2]), .E(n983), .CK(clk), .Q(R3[2]) );
  EDFFX1 R3_reg_1_ ( .D(data_in_1[1]), .E(n982), .CK(clk), .Q(R3[1]) );
  EDFFX1 R3_reg_0_ ( .D(data_in_1[0]), .E(n983), .CK(clk), .Q(R3[0]) );
  EDFFX1 R7_reg_33_ ( .D(data_in_1[33]), .E(n990), .CK(clk), .Q(R7[33]) );
  EDFFX1 R7_reg_32_ ( .D(data_in_1[32]), .E(n991), .CK(clk), .Q(R7[32]) );
  EDFFX1 R7_reg_31_ ( .D(data_in_1[31]), .E(n990), .CK(clk), .Q(R7[31]) );
  EDFFX1 R7_reg_30_ ( .D(data_in_1[30]), .E(n991), .CK(clk), .Q(R7[30]) );
  EDFFX1 R7_reg_29_ ( .D(data_in_1[29]), .E(n990), .CK(clk), .Q(R7[29]) );
  EDFFX1 R7_reg_28_ ( .D(data_in_1[28]), .E(n991), .CK(clk), .Q(R7[28]) );
  EDFFX1 R7_reg_27_ ( .D(data_in_1[27]), .E(n990), .CK(clk), .Q(R7[27]) );
  EDFFX1 R7_reg_26_ ( .D(data_in_1[26]), .E(n991), .CK(clk), .Q(R7[26]) );
  EDFFX1 R7_reg_25_ ( .D(data_in_1[25]), .E(n990), .CK(clk), .Q(R7[25]) );
  EDFFX1 R7_reg_24_ ( .D(data_in_1[24]), .E(n991), .CK(clk), .Q(R7[24]) );
  EDFFX1 R7_reg_23_ ( .D(data_in_1[23]), .E(n991), .CK(clk), .Q(R7[23]) );
  EDFFX1 R7_reg_22_ ( .D(data_in_1[22]), .E(n991), .CK(clk), .Q(R7[22]) );
  EDFFX1 R7_reg_21_ ( .D(data_in_1[21]), .E(n991), .CK(clk), .Q(R7[21]) );
  EDFFX1 R7_reg_20_ ( .D(data_in_1[20]), .E(n991), .CK(clk), .Q(R7[20]) );
  EDFFX1 R7_reg_19_ ( .D(data_in_1[19]), .E(n991), .CK(clk), .Q(R7[19]) );
  EDFFX1 R7_reg_18_ ( .D(data_in_1[18]), .E(n991), .CK(clk), .Q(R7[18]) );
  EDFFX1 R7_reg_17_ ( .D(data_in_1[17]), .E(n991), .CK(clk), .Q(R7[17]) );
  EDFFX1 R7_reg_16_ ( .D(data_in_1[16]), .E(n991), .CK(clk), .Q(R7[16]) );
  EDFFX1 R7_reg_15_ ( .D(data_in_1[15]), .E(n991), .CK(clk), .Q(R7[15]) );
  EDFFX1 R7_reg_14_ ( .D(data_in_1[14]), .E(n991), .CK(clk), .Q(R7[14]) );
  EDFFX1 R7_reg_13_ ( .D(data_in_1[13]), .E(n991), .CK(clk), .Q(R7[13]) );
  EDFFX1 R7_reg_12_ ( .D(data_in_1[12]), .E(n991), .CK(clk), .Q(R7[12]) );
  EDFFX1 R7_reg_11_ ( .D(data_in_1[11]), .E(n990), .CK(clk), .Q(R7[11]) );
  EDFFX1 R7_reg_10_ ( .D(data_in_1[10]), .E(n990), .CK(clk), .Q(R7[10]) );
  EDFFX1 R7_reg_9_ ( .D(data_in_1[9]), .E(n990), .CK(clk), .Q(R7[9]) );
  EDFFX1 R7_reg_8_ ( .D(data_in_1[8]), .E(n990), .CK(clk), .Q(R7[8]) );
  EDFFX1 R7_reg_7_ ( .D(data_in_1[7]), .E(n990), .CK(clk), .Q(R7[7]) );
  EDFFX1 R7_reg_6_ ( .D(data_in_1[6]), .E(n990), .CK(clk), .Q(R7[6]) );
  EDFFX1 R7_reg_5_ ( .D(data_in_1[5]), .E(n990), .CK(clk), .Q(R7[5]) );
  EDFFX1 R7_reg_4_ ( .D(data_in_1[4]), .E(n990), .CK(clk), .Q(R7[4]) );
  EDFFX1 R7_reg_3_ ( .D(data_in_1[3]), .E(n990), .CK(clk), .Q(R7[3]) );
  EDFFX1 R7_reg_2_ ( .D(data_in_1[2]), .E(n990), .CK(clk), .Q(R7[2]) );
  EDFFX1 R7_reg_1_ ( .D(data_in_1[1]), .E(n990), .CK(clk), .Q(R7[1]) );
  EDFFX1 R7_reg_0_ ( .D(data_in_1[0]), .E(n990), .CK(clk), .Q(R7[0]) );
  EDFFX1 R11_reg_33_ ( .D(data_in_1[33]), .E(n971), .CK(clk), .Q(R11[33]) );
  EDFFX1 R11_reg_32_ ( .D(data_in_1[32]), .E(n971), .CK(clk), .Q(R11[32]) );
  EDFFX1 R11_reg_31_ ( .D(data_in_1[31]), .E(n971), .CK(clk), .Q(R11[31]) );
  EDFFX1 R11_reg_30_ ( .D(data_in_1[30]), .E(n971), .CK(clk), .Q(R11[30]) );
  EDFFX1 R11_reg_29_ ( .D(data_in_1[29]), .E(n971), .CK(clk), .Q(R11[29]) );
  EDFFX1 R11_reg_28_ ( .D(data_in_1[28]), .E(n971), .CK(clk), .Q(R11[28]) );
  EDFFX1 R11_reg_27_ ( .D(data_in_1[27]), .E(n971), .CK(clk), .Q(R11[27]) );
  EDFFX1 R11_reg_26_ ( .D(data_in_1[26]), .E(n971), .CK(clk), .Q(R11[26]) );
  EDFFX1 R11_reg_25_ ( .D(data_in_1[25]), .E(n1002), .CK(clk), .Q(R11[25]) );
  EDFFX1 R11_reg_24_ ( .D(data_in_1[24]), .E(n1001), .CK(clk), .Q(R11[24]) );
  EDFFX1 R11_reg_23_ ( .D(data_in_1[23]), .E(n1002), .CK(clk), .Q(R11[23]) );
  EDFFX1 R11_reg_22_ ( .D(data_in_1[22]), .E(n1002), .CK(clk), .Q(R11[22]) );
  EDFFX1 R11_reg_21_ ( .D(data_in_1[21]), .E(n1001), .CK(clk), .Q(R11[21]) );
  EDFFX1 R11_reg_20_ ( .D(data_in_1[20]), .E(n1001), .CK(clk), .Q(R11[20]) );
  EDFFX1 R11_reg_19_ ( .D(data_in_1[19]), .E(n1001), .CK(clk), .Q(R11[19]) );
  EDFFX1 R11_reg_18_ ( .D(data_in_1[18]), .E(n1001), .CK(clk), .Q(R11[18]) );
  EDFFX1 R11_reg_17_ ( .D(data_in_1[17]), .E(n1001), .CK(clk), .Q(R11[17]) );
  EDFFX1 R11_reg_16_ ( .D(data_in_1[16]), .E(n1001), .CK(clk), .Q(R11[16]) );
  EDFFX1 R11_reg_15_ ( .D(data_in_1[15]), .E(n1001), .CK(clk), .Q(R11[15]) );
  EDFFX1 R11_reg_14_ ( .D(data_in_1[14]), .E(n1001), .CK(clk), .Q(R11[14]) );
  EDFFX1 R11_reg_13_ ( .D(data_in_1[13]), .E(n1001), .CK(clk), .Q(R11[13]) );
  EDFFX1 R11_reg_12_ ( .D(data_in_1[12]), .E(n1001), .CK(clk), .Q(R11[12]) );
  EDFFX1 R11_reg_11_ ( .D(data_in_1[11]), .E(n1001), .CK(clk), .Q(R11[11]) );
  EDFFX1 R11_reg_10_ ( .D(data_in_1[10]), .E(n1001), .CK(clk), .Q(R11[10]) );
  EDFFX1 R11_reg_9_ ( .D(data_in_1[9]), .E(n1002), .CK(clk), .Q(R11[9]) );
  EDFFX1 R11_reg_8_ ( .D(data_in_1[8]), .E(n1002), .CK(clk), .Q(R11[8]) );
  EDFFX1 R11_reg_7_ ( .D(data_in_1[7]), .E(n1002), .CK(clk), .Q(R11[7]) );
  EDFFX1 R11_reg_6_ ( .D(data_in_1[6]), .E(n1002), .CK(clk), .Q(R11[6]) );
  EDFFX1 R11_reg_5_ ( .D(data_in_1[5]), .E(n1002), .CK(clk), .Q(R11[5]) );
  EDFFX1 R11_reg_4_ ( .D(data_in_1[4]), .E(n1002), .CK(clk), .Q(R11[4]) );
  EDFFX1 R11_reg_3_ ( .D(data_in_1[3]), .E(n1002), .CK(clk), .Q(R11[3]) );
  EDFFX1 R11_reg_2_ ( .D(data_in_1[2]), .E(n1002), .CK(clk), .Q(R11[2]) );
  EDFFX1 R11_reg_1_ ( .D(data_in_1[1]), .E(n1002), .CK(clk), .Q(R11[1]) );
  EDFFX1 R11_reg_0_ ( .D(data_in_1[0]), .E(n1002), .CK(clk), .Q(R11[0]) );
  DFFHQX1 data_out_1_reg_51_ ( .D(n916), .CK(clk), .Q(data_out_1[51]) );
  DFFHQX1 data_out_1_reg_34_ ( .D(n933), .CK(clk), .Q(data_out_1[34]) );
  DFFHQX1 data_out_1_reg_85_ ( .D(n882), .CK(clk), .Q(data_out_1[85]) );
  DFFHQX1 data_out_1_reg_68_ ( .D(n899), .CK(clk), .Q(data_out_1[68]) );
  DFFHQX1 data_out_1_reg_119_ ( .D(n848), .CK(clk), .Q(data_out_1[119]) );
  DFFHQX1 data_out_1_reg_102_ ( .D(n865), .CK(clk), .Q(data_out_1[102]) );
  DFFHQX1 data_out_1_reg_66_ ( .D(n901), .CK(clk), .Q(data_out_1[66]) );
  DFFHQX1 data_out_1_reg_65_ ( .D(n902), .CK(clk), .Q(data_out_1[65]) );
  DFFHQX1 data_out_1_reg_64_ ( .D(n903), .CK(clk), .Q(data_out_1[64]) );
  DFFHQX1 data_out_1_reg_63_ ( .D(n904), .CK(clk), .Q(data_out_1[63]) );
  DFFHQX1 data_out_1_reg_62_ ( .D(n905), .CK(clk), .Q(data_out_1[62]) );
  DFFHQX1 data_out_1_reg_61_ ( .D(n906), .CK(clk), .Q(data_out_1[61]) );
  DFFHQX1 data_out_1_reg_60_ ( .D(n907), .CK(clk), .Q(data_out_1[60]) );
  DFFHQX1 data_out_1_reg_59_ ( .D(n908), .CK(clk), .Q(data_out_1[59]) );
  DFFHQX1 data_out_1_reg_58_ ( .D(n909), .CK(clk), .Q(data_out_1[58]) );
  DFFHQX1 data_out_1_reg_57_ ( .D(n910), .CK(clk), .Q(data_out_1[57]) );
  DFFHQX1 data_out_1_reg_56_ ( .D(n911), .CK(clk), .Q(data_out_1[56]) );
  DFFHQX1 data_out_1_reg_55_ ( .D(n912), .CK(clk), .Q(data_out_1[55]) );
  DFFHQX1 data_out_1_reg_54_ ( .D(n913), .CK(clk), .Q(data_out_1[54]) );
  DFFHQX1 data_out_1_reg_53_ ( .D(n914), .CK(clk), .Q(data_out_1[53]) );
  DFFHQX1 data_out_1_reg_52_ ( .D(n915), .CK(clk), .Q(data_out_1[52]) );
  DFFHQX1 data_out_1_reg_49_ ( .D(n918), .CK(clk), .Q(data_out_1[49]) );
  DFFHQX1 data_out_1_reg_48_ ( .D(n919), .CK(clk), .Q(data_out_1[48]) );
  DFFHQX1 data_out_1_reg_47_ ( .D(n920), .CK(clk), .Q(data_out_1[47]) );
  DFFHQX1 data_out_1_reg_46_ ( .D(n921), .CK(clk), .Q(data_out_1[46]) );
  DFFHQX1 data_out_1_reg_45_ ( .D(n922), .CK(clk), .Q(data_out_1[45]) );
  DFFHQX1 data_out_1_reg_44_ ( .D(n923), .CK(clk), .Q(data_out_1[44]) );
  DFFHQX1 data_out_1_reg_43_ ( .D(n924), .CK(clk), .Q(data_out_1[43]) );
  DFFHQX1 data_out_1_reg_42_ ( .D(n925), .CK(clk), .Q(data_out_1[42]) );
  DFFHQX1 data_out_1_reg_41_ ( .D(n926), .CK(clk), .Q(data_out_1[41]) );
  DFFHQX1 data_out_1_reg_40_ ( .D(n927), .CK(clk), .Q(data_out_1[40]) );
  DFFHQX1 data_out_1_reg_39_ ( .D(n928), .CK(clk), .Q(data_out_1[39]) );
  DFFHQX1 data_out_1_reg_38_ ( .D(n929), .CK(clk), .Q(data_out_1[38]) );
  DFFHQX1 data_out_1_reg_37_ ( .D(n930), .CK(clk), .Q(data_out_1[37]) );
  DFFHQX1 data_out_1_reg_36_ ( .D(n931), .CK(clk), .Q(data_out_1[36]) );
  DFFHQX1 data_out_1_reg_35_ ( .D(n932), .CK(clk), .Q(data_out_1[35]) );
  DFFHQX1 data_out_1_reg_100_ ( .D(n867), .CK(clk), .Q(data_out_1[100]) );
  DFFHQX1 data_out_1_reg_99_ ( .D(n868), .CK(clk), .Q(data_out_1[99]) );
  DFFHQX1 data_out_1_reg_98_ ( .D(n869), .CK(clk), .Q(data_out_1[98]) );
  DFFHQX1 data_out_1_reg_97_ ( .D(n870), .CK(clk), .Q(data_out_1[97]) );
  DFFHQX1 data_out_1_reg_96_ ( .D(n871), .CK(clk), .Q(data_out_1[96]) );
  DFFHQX1 data_out_1_reg_95_ ( .D(n872), .CK(clk), .Q(data_out_1[95]) );
  DFFHQX1 data_out_1_reg_94_ ( .D(n873), .CK(clk), .Q(data_out_1[94]) );
  DFFHQX1 data_out_1_reg_93_ ( .D(n874), .CK(clk), .Q(data_out_1[93]) );
  DFFHQX1 data_out_1_reg_92_ ( .D(n875), .CK(clk), .Q(data_out_1[92]) );
  DFFHQX1 data_out_1_reg_91_ ( .D(n876), .CK(clk), .Q(data_out_1[91]) );
  DFFHQX1 data_out_1_reg_90_ ( .D(n877), .CK(clk), .Q(data_out_1[90]) );
  DFFHQX1 data_out_1_reg_89_ ( .D(n878), .CK(clk), .Q(data_out_1[89]) );
  DFFHQX1 data_out_1_reg_88_ ( .D(n879), .CK(clk), .Q(data_out_1[88]) );
  DFFHQX1 data_out_1_reg_87_ ( .D(n880), .CK(clk), .Q(data_out_1[87]) );
  DFFHQX1 data_out_1_reg_86_ ( .D(n881), .CK(clk), .Q(data_out_1[86]) );
  DFFHQX1 data_out_1_reg_83_ ( .D(n884), .CK(clk), .Q(data_out_1[83]) );
  DFFHQX1 data_out_1_reg_82_ ( .D(n885), .CK(clk), .Q(data_out_1[82]) );
  DFFHQX1 data_out_1_reg_81_ ( .D(n886), .CK(clk), .Q(data_out_1[81]) );
  DFFHQX1 data_out_1_reg_80_ ( .D(n887), .CK(clk), .Q(data_out_1[80]) );
  DFFHQX1 data_out_1_reg_79_ ( .D(n888), .CK(clk), .Q(data_out_1[79]) );
  DFFHQX1 data_out_1_reg_78_ ( .D(n889), .CK(clk), .Q(data_out_1[78]) );
  DFFHQX1 data_out_1_reg_77_ ( .D(n890), .CK(clk), .Q(data_out_1[77]) );
  DFFHQX1 data_out_1_reg_76_ ( .D(n891), .CK(clk), .Q(data_out_1[76]) );
  DFFHQX1 data_out_1_reg_75_ ( .D(n892), .CK(clk), .Q(data_out_1[75]) );
  DFFHQX1 data_out_1_reg_74_ ( .D(n893), .CK(clk), .Q(data_out_1[74]) );
  DFFHQX1 data_out_1_reg_73_ ( .D(n894), .CK(clk), .Q(data_out_1[73]) );
  DFFHQX1 data_out_1_reg_72_ ( .D(n895), .CK(clk), .Q(data_out_1[72]) );
  DFFHQX1 data_out_1_reg_71_ ( .D(n896), .CK(clk), .Q(data_out_1[71]) );
  DFFHQX1 data_out_1_reg_70_ ( .D(n897), .CK(clk), .Q(data_out_1[70]) );
  DFFHQX1 data_out_1_reg_69_ ( .D(n898), .CK(clk), .Q(data_out_1[69]) );
  DFFHQX1 data_out_1_reg_134_ ( .D(n833), .CK(clk), .Q(data_out_1[134]) );
  DFFHQX1 data_out_1_reg_133_ ( .D(n834), .CK(clk), .Q(data_out_1[133]) );
  DFFHQX1 data_out_1_reg_132_ ( .D(n835), .CK(clk), .Q(data_out_1[132]) );
  DFFHQX1 data_out_1_reg_131_ ( .D(n836), .CK(clk), .Q(data_out_1[131]) );
  DFFHQX1 data_out_1_reg_130_ ( .D(n837), .CK(clk), .Q(data_out_1[130]) );
  DFFHQX1 data_out_1_reg_129_ ( .D(n838), .CK(clk), .Q(data_out_1[129]) );
  DFFHQX1 data_out_1_reg_128_ ( .D(n839), .CK(clk), .Q(data_out_1[128]) );
  DFFHQX1 data_out_1_reg_127_ ( .D(n840), .CK(clk), .Q(data_out_1[127]) );
  DFFHQX1 data_out_1_reg_126_ ( .D(n841), .CK(clk), .Q(data_out_1[126]) );
  DFFHQX1 data_out_1_reg_125_ ( .D(n842), .CK(clk), .Q(data_out_1[125]) );
  DFFHQX1 data_out_1_reg_124_ ( .D(n843), .CK(clk), .Q(data_out_1[124]) );
  DFFHQX1 data_out_1_reg_123_ ( .D(n844), .CK(clk), .Q(data_out_1[123]) );
  DFFHQX1 data_out_1_reg_122_ ( .D(n845), .CK(clk), .Q(data_out_1[122]) );
  DFFHQX1 data_out_1_reg_121_ ( .D(n846), .CK(clk), .Q(data_out_1[121]) );
  DFFHQX1 data_out_1_reg_120_ ( .D(n847), .CK(clk), .Q(data_out_1[120]) );
  DFFHQX1 data_out_1_reg_117_ ( .D(n850), .CK(clk), .Q(data_out_1[117]) );
  DFFHQX1 data_out_1_reg_116_ ( .D(n851), .CK(clk), .Q(data_out_1[116]) );
  DFFHQX1 data_out_1_reg_115_ ( .D(n852), .CK(clk), .Q(data_out_1[115]) );
  DFFHQX1 data_out_1_reg_114_ ( .D(n853), .CK(clk), .Q(data_out_1[114]) );
  DFFHQX1 data_out_1_reg_113_ ( .D(n854), .CK(clk), .Q(data_out_1[113]) );
  DFFHQX1 data_out_1_reg_112_ ( .D(n855), .CK(clk), .Q(data_out_1[112]) );
  DFFHQX1 data_out_1_reg_111_ ( .D(n856), .CK(clk), .Q(data_out_1[111]) );
  DFFHQX1 data_out_1_reg_110_ ( .D(n857), .CK(clk), .Q(data_out_1[110]) );
  DFFHQX1 data_out_1_reg_109_ ( .D(n858), .CK(clk), .Q(data_out_1[109]) );
  DFFHQX1 data_out_1_reg_108_ ( .D(n859), .CK(clk), .Q(data_out_1[108]) );
  DFFHQX1 data_out_1_reg_107_ ( .D(n860), .CK(clk), .Q(data_out_1[107]) );
  DFFHQX1 data_out_1_reg_106_ ( .D(n861), .CK(clk), .Q(data_out_1[106]) );
  DFFHQX1 data_out_1_reg_105_ ( .D(n862), .CK(clk), .Q(data_out_1[105]) );
  DFFHQX1 data_out_1_reg_104_ ( .D(n863), .CK(clk), .Q(data_out_1[104]) );
  DFFHQX1 data_out_1_reg_103_ ( .D(n864), .CK(clk), .Q(data_out_1[103]) );
  DFFRHQX1 s_p_flag_out_reg ( .D(n1005), .CK(clk), .RN(rst_n), .Q(s_p_flag_out) );
  DFFHQX1 data_out_1_reg_33_ ( .D(n934), .CK(clk), .Q(data_out_1[33]) );
  DFFHQX1 data_out_1_reg_16_ ( .D(n951), .CK(clk), .Q(data_out_1[16]) );
  JKFFRXL counter_reg_0_ ( .J(1'b1), .K(1'b1), .CK(clk), .RN(rst_n), .Q(
        counter[0]), .QN(n550) );
  DFFHQX1 data_out_1_reg_32_ ( .D(n935), .CK(clk), .Q(data_out_1[32]) );
  DFFHQX1 data_out_1_reg_31_ ( .D(n936), .CK(clk), .Q(data_out_1[31]) );
  DFFHQX1 data_out_1_reg_15_ ( .D(n952), .CK(clk), .Q(data_out_1[15]) );
  DFFHQX1 data_out_1_reg_14_ ( .D(n953), .CK(clk), .Q(data_out_1[14]) );
  DFFHQX1 data_out_1_reg_13_ ( .D(n954), .CK(clk), .Q(data_out_1[13]) );
  DFFRHQX1 counter_reg_3_ ( .D(N15), .CK(clk), .RN(rst_n), .Q(counter[3]) );
  DFFRHQX1 counter_reg_1_ ( .D(N13), .CK(clk), .RN(rst_n), .Q(counter[1]) );
  DFFRHQX1 counter_reg_2_ ( .D(N14), .CK(clk), .RN(rst_n), .Q(counter[2]) );
  DFFHQX1 data_out_1_reg_30_ ( .D(n937), .CK(clk), .Q(data_out_1[30]) );
  DFFHQX1 data_out_1_reg_29_ ( .D(n938), .CK(clk), .Q(data_out_1[29]) );
  DFFHQX1 data_out_1_reg_28_ ( .D(n939), .CK(clk), .Q(data_out_1[28]) );
  DFFHQX1 data_out_1_reg_27_ ( .D(n940), .CK(clk), .Q(data_out_1[27]) );
  DFFHQX1 data_out_1_reg_26_ ( .D(n941), .CK(clk), .Q(data_out_1[26]) );
  DFFHQX1 data_out_1_reg_25_ ( .D(n942), .CK(clk), .Q(data_out_1[25]) );
  DFFHQX1 data_out_1_reg_23_ ( .D(n944), .CK(clk), .Q(data_out_1[23]) );
  DFFHQX1 data_out_1_reg_21_ ( .D(n946), .CK(clk), .Q(data_out_1[21]) );
  DFFHQX1 data_out_1_reg_20_ ( .D(n947), .CK(clk), .Q(data_out_1[20]) );
  DFFHQX1 data_out_1_reg_17_ ( .D(n950), .CK(clk), .Q(data_out_1[17]) );
  DFFHQX1 data_out_1_reg_12_ ( .D(n955), .CK(clk), .Q(data_out_1[12]) );
  DFFHQX1 data_out_1_reg_11_ ( .D(n956), .CK(clk), .Q(data_out_1[11]) );
  DFFHQX1 data_out_1_reg_10_ ( .D(n957), .CK(clk), .Q(data_out_1[10]) );
  DFFHQX1 data_out_1_reg_9_ ( .D(n958), .CK(clk), .Q(data_out_1[9]) );
  DFFHQX1 data_out_1_reg_8_ ( .D(n959), .CK(clk), .Q(data_out_1[8]) );
  DFFHQX1 data_out_1_reg_6_ ( .D(n961), .CK(clk), .Q(data_out_1[6]) );
  DFFHQX1 data_out_1_reg_5_ ( .D(n962), .CK(clk), .Q(data_out_1[5]) );
  DFFHQX1 data_out_1_reg_4_ ( .D(n963), .CK(clk), .Q(data_out_1[4]) );
  DFFHQX1 data_out_1_reg_24_ ( .D(n943), .CK(clk), .Q(data_out_1[24]) );
  DFFHQX1 data_out_1_reg_22_ ( .D(n945), .CK(clk), .Q(data_out_1[22]) );
  DFFHQX1 data_out_1_reg_7_ ( .D(n960), .CK(clk), .Q(data_out_1[7]) );
  DFFHQX1 data_out_1_reg_18_ ( .D(n949), .CK(clk), .Q(data_out_1[18]) );
  DFFHQX1 data_out_1_reg_3_ ( .D(n964), .CK(clk), .Q(data_out_1[3]) );
  DFFHQX1 data_out_1_reg_2_ ( .D(n965), .CK(clk), .Q(data_out_1[2]) );
  DFFHQX1 data_out_1_reg_1_ ( .D(n966), .CK(clk), .Q(data_out_1[1]) );
  DFFHQX1 data_out_1_reg_0_ ( .D(n967), .CK(clk), .Q(data_out_1[0]) );
  DFFHQX1 data_out_1_reg_19_ ( .D(n948), .CK(clk), .Q(data_out_1[19]) );
  DFFHQX1 data_out_1_reg_118_ ( .D(n849), .CK(clk), .Q(data_out_1[118]) );
  DFFHQX1 data_out_1_reg_135_ ( .D(n832), .CK(clk), .Q(data_out_1[135]) );
  DFFHQX1 data_out_1_reg_50_ ( .D(n917), .CK(clk), .Q(data_out_1[50]) );
  DFFHQX1 data_out_1_reg_67_ ( .D(n900), .CK(clk), .Q(data_out_1[67]) );
  DFFHQX2 data_out_1_reg_101_ ( .D(n866), .CK(clk), .Q(data_out_1[101]) );
  DFFHQX2 data_out_1_reg_84_ ( .D(n883), .CK(clk), .Q(data_out_1[84]) );
  OR3XL U4 ( .A(n1043), .B(n1042), .C(n825), .Y(n1) );
  OR2X2 U5 ( .A(n829), .B(n826), .Y(n2) );
  OR2X2 U6 ( .A(n826), .B(n830), .Y(n3) );
  OR2X2 U7 ( .A(n824), .B(n829), .Y(n4) );
  OR2X2 U8 ( .A(n824), .B(n830), .Y(n5) );
  OR2X2 U9 ( .A(n825), .B(n829), .Y(n6) );
  OR2X2 U10 ( .A(n825), .B(n830), .Y(n7) );
  OR2X2 U11 ( .A(n828), .B(n829), .Y(n8) );
  AOI22XL U12 ( .A0(R3[0]), .A1(n1039), .B0(data_out_1[0]), .B1(n1017), .Y(
        n822) );
  AOI22XL U13 ( .A0(R3[1]), .A1(n1039), .B0(data_out_1[1]), .B1(n1018), .Y(
        n820) );
  AOI22XL U14 ( .A0(R3[2]), .A1(n1039), .B0(data_out_1[2]), .B1(n1017), .Y(
        n818) );
  AOI22XL U15 ( .A0(R3[3]), .A1(n1039), .B0(data_out_1[3]), .B1(n1018), .Y(
        n816) );
  AOI22XL U16 ( .A0(R3[7]), .A1(n1038), .B0(data_out_1[7]), .B1(n1017), .Y(
        n808) );
  AOI22XL U17 ( .A0(R3[17]), .A1(n1038), .B0(data_out_1[17]), .B1(n1017), .Y(
        n788) );
  AOI22XL U18 ( .A0(R3[18]), .A1(n1038), .B0(data_out_1[18]), .B1(n1017), .Y(
        n786) );
  AOI22XL U19 ( .A0(R3[19]), .A1(n1038), .B0(data_out_1[19]), .B1(n1017), .Y(
        n784) );
  AOI22XL U20 ( .A0(R3[20]), .A1(n1037), .B0(data_out_1[20]), .B1(n1017), .Y(
        n782) );
  AOI22XL U21 ( .A0(R3[24]), .A1(n1037), .B0(data_out_1[24]), .B1(n1019), .Y(
        n774) );
  INVX1 U22 ( .A(n9), .Y(n1023) );
  INVX1 U23 ( .A(n9), .Y(n1024) );
  INVX1 U24 ( .A(n9), .Y(n1021) );
  INVX1 U25 ( .A(n9), .Y(n1022) );
  INVX1 U26 ( .A(n9), .Y(n1018) );
  INVX1 U27 ( .A(n9), .Y(n1019) );
  INVX1 U28 ( .A(n9), .Y(n1020) );
  INVX1 U29 ( .A(n9), .Y(n1017) );
  CLKINVX3 U30 ( .A(n1029), .Y(n1025) );
  CLKINVX3 U31 ( .A(n1016), .Y(n1012) );
  CLKINVX3 U32 ( .A(n1), .Y(n1007) );
  OR4X2 U33 ( .A(n1012), .B(n1007), .C(n1025), .D(N171), .Y(n9) );
  CLKINVX3 U34 ( .A(n1), .Y(n1009) );
  CLKINVX3 U35 ( .A(n1), .Y(n1008) );
  CLKINVX3 U36 ( .A(n1), .Y(n1011) );
  CLKINVX3 U37 ( .A(n1), .Y(n1010) );
  CLKINVX3 U38 ( .A(n1029), .Y(n1028) );
  INVX1 U39 ( .A(n1040), .Y(n1030) );
  INVX1 U40 ( .A(n1040), .Y(n1033) );
  INVX1 U41 ( .A(n1040), .Y(n1032) );
  INVX1 U42 ( .A(n1040), .Y(n1031) );
  INVX1 U43 ( .A(n1040), .Y(n1035) );
  INVX1 U44 ( .A(n1040), .Y(n1034) );
  INVX1 U45 ( .A(n1040), .Y(n1038) );
  INVX1 U46 ( .A(n1040), .Y(n1037) );
  INVX1 U47 ( .A(n1040), .Y(n1036) );
  CLKINVX3 U48 ( .A(n1029), .Y(n1026) );
  CLKINVX3 U49 ( .A(n1029), .Y(n1027) );
  INVX1 U50 ( .A(n1040), .Y(n1039) );
  CLKINVX3 U51 ( .A(n1016), .Y(n1013) );
  CLKINVX3 U52 ( .A(n1016), .Y(n1014) );
  CLKINVX3 U53 ( .A(n1016), .Y(n1015) );
  INVX1 U54 ( .A(n1006), .Y(n1004) );
  INVX1 U55 ( .A(n1003), .Y(n1001) );
  INVX1 U56 ( .A(n1000), .Y(n998) );
  INVX1 U57 ( .A(n997), .Y(n995) );
  INVX1 U58 ( .A(n994), .Y(n992) );
  INVX1 U59 ( .A(n2), .Y(n990) );
  INVX1 U60 ( .A(n2), .Y(n991) );
  INVX1 U61 ( .A(n4), .Y(n989) );
  INVX1 U62 ( .A(n6), .Y(n987) );
  INVX1 U63 ( .A(n8), .Y(n985) );
  INVX1 U64 ( .A(n3), .Y(n983) );
  INVX1 U65 ( .A(n5), .Y(n981) );
  INVX1 U66 ( .A(n7), .Y(n979) );
  INVX1 U67 ( .A(n1006), .Y(n1005) );
  INVX1 U68 ( .A(n1003), .Y(n1002) );
  INVX1 U69 ( .A(n1000), .Y(n999) );
  INVX1 U70 ( .A(n997), .Y(n996) );
  INVX1 U71 ( .A(n994), .Y(n993) );
  INVX1 U72 ( .A(N230), .Y(n1029) );
  INVX1 U73 ( .A(n968), .Y(n1016) );
  INVX1 U74 ( .A(N171), .Y(n1040) );
  INVX1 U75 ( .A(n4), .Y(n988) );
  INVX1 U76 ( .A(n6), .Y(n986) );
  INVX1 U77 ( .A(n8), .Y(n984) );
  INVX1 U78 ( .A(n3), .Y(n982) );
  INVX1 U79 ( .A(n5), .Y(n980) );
  INVX1 U80 ( .A(n7), .Y(n978) );
  INVX1 U81 ( .A(n970), .Y(n1006) );
  INVX1 U82 ( .A(n971), .Y(n1003) );
  INVX1 U83 ( .A(n972), .Y(n1000) );
  INVX1 U84 ( .A(n973), .Y(n997) );
  INVX1 U85 ( .A(n974), .Y(n994) );
  NOR3X1 U86 ( .A(n1043), .B(n1042), .C(n824), .Y(n968) );
  NOR3X1 U87 ( .A(n1042), .B(n826), .C(n1043), .Y(N230) );
  NOR2X1 U88 ( .A(n830), .B(n828), .Y(N171) );
  NAND2X1 U89 ( .A(n1042), .B(n1043), .Y(n830) );
  NOR3X1 U90 ( .A(n1043), .B(n1042), .C(n828), .Y(n970) );
  OAI211X1 U91 ( .A0(n831), .A1(n1043), .B0(n827), .C0(n2), .Y(N15) );
  NOR2X1 U92 ( .A(n826), .B(n827), .Y(n971) );
  NOR2X1 U93 ( .A(n824), .B(n827), .Y(n972) );
  NOR2X1 U94 ( .A(n825), .B(n827), .Y(n973) );
  NOR2X1 U95 ( .A(n828), .B(n827), .Y(n974) );
  NAND2X1 U96 ( .A(n824), .B(n825), .Y(N13) );
  INVX1 U97 ( .A(counter[2]), .Y(n1042) );
  INVX1 U98 ( .A(counter[3]), .Y(n1043) );
  NAND2X1 U99 ( .A(counter[0]), .B(n1041), .Y(n825) );
  NAND2X1 U100 ( .A(counter[1]), .B(counter[0]), .Y(n826) );
  NAND2X1 U101 ( .A(counter[1]), .B(n550), .Y(n824) );
  NAND2X1 U102 ( .A(n550), .B(n1041), .Y(n828) );
  INVX1 U103 ( .A(counter[1]), .Y(n1041) );
  NAND2X1 U104 ( .A(n618), .B(n619), .Y(n865) );
  AOI222X1 U105 ( .A0(R12[0]), .A1(n1011), .B0(R14[0]), .B1(n1028), .C0(R13[0]), .C1(n1013), .Y(n619) );
  AOI22X1 U106 ( .A0(R15[0]), .A1(n1031), .B0(data_out_1[102]), .B1(n1022), 
        .Y(n618) );
  NAND2X1 U107 ( .A(n616), .B(n617), .Y(n864) );
  AOI222X1 U108 ( .A0(R12[1]), .A1(n1008), .B0(R14[1]), .B1(n1026), .C0(R13[1]), .C1(n1013), .Y(n617) );
  AOI22X1 U109 ( .A0(R15[1]), .A1(n1031), .B0(data_out_1[103]), .B1(n1022), 
        .Y(n616) );
  NAND2X1 U110 ( .A(n614), .B(n615), .Y(n863) );
  AOI222X1 U111 ( .A0(R12[2]), .A1(n1008), .B0(R14[2]), .B1(n1027), .C0(R13[2]), .C1(n1013), .Y(n615) );
  AOI22X1 U112 ( .A0(R15[2]), .A1(n1031), .B0(data_out_1[104]), .B1(n1022), 
        .Y(n614) );
  NAND2X1 U113 ( .A(n612), .B(n613), .Y(n862) );
  AOI222X1 U114 ( .A0(R12[3]), .A1(n1008), .B0(R14[3]), .B1(n1027), .C0(R13[3]), .C1(n1013), .Y(n613) );
  AOI22X1 U115 ( .A0(R15[3]), .A1(n1031), .B0(data_out_1[105]), .B1(n1022), 
        .Y(n612) );
  NAND2X1 U116 ( .A(n610), .B(n611), .Y(n861) );
  AOI222X1 U117 ( .A0(R12[4]), .A1(n1009), .B0(R14[4]), .B1(n1026), .C0(R13[4]), .C1(n1013), .Y(n611) );
  AOI22X1 U118 ( .A0(R15[4]), .A1(n1031), .B0(data_out_1[106]), .B1(n1022), 
        .Y(n610) );
  NAND2X1 U119 ( .A(n608), .B(n609), .Y(n860) );
  AOI222X1 U120 ( .A0(R12[5]), .A1(n1008), .B0(R14[5]), .B1(n1026), .C0(R13[5]), .C1(n1013), .Y(n609) );
  AOI22X1 U121 ( .A0(R15[5]), .A1(n1031), .B0(data_out_1[107]), .B1(n1022), 
        .Y(n608) );
  NAND2X1 U122 ( .A(n606), .B(n607), .Y(n859) );
  AOI222X1 U123 ( .A0(R12[6]), .A1(n1010), .B0(R14[6]), .B1(n1027), .C0(R13[6]), .C1(n1013), .Y(n607) );
  AOI22X1 U124 ( .A0(R15[6]), .A1(n1031), .B0(data_out_1[108]), .B1(n1023), 
        .Y(n606) );
  NAND2X1 U125 ( .A(n604), .B(n605), .Y(n858) );
  AOI222X1 U126 ( .A0(R12[7]), .A1(n1008), .B0(R14[7]), .B1(n1027), .C0(R13[7]), .C1(n1013), .Y(n605) );
  AOI22X1 U127 ( .A0(R15[7]), .A1(n1031), .B0(data_out_1[109]), .B1(n1023), 
        .Y(n604) );
  NAND2X1 U128 ( .A(n602), .B(n603), .Y(n857) );
  AOI222X1 U129 ( .A0(R12[8]), .A1(n1011), .B0(R14[8]), .B1(n1027), .C0(R13[8]), .C1(n1013), .Y(n603) );
  AOI22X1 U130 ( .A0(R15[8]), .A1(n1030), .B0(data_out_1[110]), .B1(n1023), 
        .Y(n602) );
  NAND2X1 U131 ( .A(n600), .B(n601), .Y(n856) );
  AOI222X1 U132 ( .A0(R12[9]), .A1(n1009), .B0(R14[9]), .B1(n1026), .C0(R13[9]), .C1(n1013), .Y(n601) );
  AOI22X1 U133 ( .A0(R15[9]), .A1(n1030), .B0(data_out_1[111]), .B1(n1023), 
        .Y(n600) );
  NAND2X1 U134 ( .A(n598), .B(n599), .Y(n855) );
  AOI222X1 U135 ( .A0(R12[10]), .A1(n1010), .B0(R14[10]), .B1(n1027), .C0(
        R13[10]), .C1(n1013), .Y(n599) );
  AOI22X1 U136 ( .A0(R15[10]), .A1(n1030), .B0(data_out_1[112]), .B1(n1023), 
        .Y(n598) );
  NAND2X1 U137 ( .A(n596), .B(n597), .Y(n854) );
  AOI222X1 U138 ( .A0(R12[11]), .A1(n1011), .B0(R14[11]), .B1(n1028), .C0(
        R13[11]), .C1(n1013), .Y(n597) );
  AOI22X1 U139 ( .A0(R15[11]), .A1(n1030), .B0(data_out_1[113]), .B1(n1023), 
        .Y(n596) );
  NAND2X1 U140 ( .A(n594), .B(n595), .Y(n853) );
  AOI222X1 U141 ( .A0(R12[12]), .A1(n1008), .B0(R14[12]), .B1(n1026), .C0(
        R13[12]), .C1(n1013), .Y(n595) );
  AOI22X1 U142 ( .A0(R15[12]), .A1(n1030), .B0(data_out_1[114]), .B1(n1023), 
        .Y(n594) );
  NAND2X1 U143 ( .A(n592), .B(n593), .Y(n852) );
  AOI222X1 U144 ( .A0(R12[13]), .A1(n1011), .B0(R14[13]), .B1(n1027), .C0(
        R13[13]), .C1(n1013), .Y(n593) );
  AOI22X1 U145 ( .A0(R15[13]), .A1(n1030), .B0(data_out_1[115]), .B1(n1023), 
        .Y(n592) );
  NAND2X1 U146 ( .A(n590), .B(n591), .Y(n851) );
  AOI222X1 U147 ( .A0(R12[14]), .A1(n1011), .B0(R14[14]), .B1(n1027), .C0(
        R13[14]), .C1(n1013), .Y(n591) );
  AOI22X1 U148 ( .A0(R15[14]), .A1(n1030), .B0(data_out_1[116]), .B1(n1023), 
        .Y(n590) );
  NAND2X1 U149 ( .A(n588), .B(n589), .Y(n850) );
  AOI222X1 U150 ( .A0(R12[15]), .A1(n1009), .B0(R14[15]), .B1(N230), .C0(
        R13[15]), .C1(n1013), .Y(n589) );
  AOI22X1 U151 ( .A0(R15[15]), .A1(n1030), .B0(data_out_1[117]), .B1(n1023), 
        .Y(n588) );
  NAND2X1 U152 ( .A(n586), .B(n587), .Y(n849) );
  AOI222X1 U153 ( .A0(R12[16]), .A1(n1008), .B0(R14[16]), .B1(n1025), .C0(
        R13[16]), .C1(n1012), .Y(n587) );
  AOI22XL U154 ( .A0(R15[16]), .A1(n1030), .B0(data_out_1[118]), .B1(n1023), 
        .Y(n586) );
  NAND2X1 U155 ( .A(n584), .B(n585), .Y(n848) );
  AOI222X1 U156 ( .A0(R12[17]), .A1(n1007), .B0(R14[17]), .B1(n1025), .C0(
        R13[17]), .C1(n1012), .Y(n585) );
  AOI22X1 U157 ( .A0(R15[17]), .A1(n1030), .B0(data_out_1[119]), .B1(n1023), 
        .Y(n584) );
  NAND2X1 U158 ( .A(n582), .B(n583), .Y(n847) );
  AOI222X1 U159 ( .A0(R12[18]), .A1(n1007), .B0(R14[18]), .B1(n1025), .C0(
        R13[18]), .C1(n1012), .Y(n583) );
  AOI22X1 U160 ( .A0(R15[18]), .A1(n1030), .B0(data_out_1[120]), .B1(n1024), 
        .Y(n582) );
  NAND2X1 U161 ( .A(n580), .B(n581), .Y(n846) );
  AOI222X1 U162 ( .A0(R12[19]), .A1(n1007), .B0(R14[19]), .B1(n1025), .C0(
        R13[19]), .C1(n1012), .Y(n581) );
  AOI22X1 U163 ( .A0(R15[19]), .A1(n1030), .B0(data_out_1[121]), .B1(n1024), 
        .Y(n580) );
  NAND2X1 U164 ( .A(n578), .B(n579), .Y(n845) );
  AOI222X1 U165 ( .A0(R12[20]), .A1(n1007), .B0(R14[20]), .B1(n1025), .C0(
        R13[20]), .C1(n1012), .Y(n579) );
  AOI22X1 U166 ( .A0(R15[20]), .A1(n1030), .B0(data_out_1[122]), .B1(n1024), 
        .Y(n578) );
  NAND2X1 U167 ( .A(n576), .B(n577), .Y(n844) );
  AOI222X1 U168 ( .A0(R12[21]), .A1(n1007), .B0(R14[21]), .B1(n1025), .C0(
        R13[21]), .C1(n1012), .Y(n577) );
  AOI22X1 U169 ( .A0(R15[21]), .A1(n1032), .B0(data_out_1[123]), .B1(n1024), 
        .Y(n576) );
  NAND2X1 U170 ( .A(n574), .B(n575), .Y(n843) );
  AOI222X1 U171 ( .A0(R12[22]), .A1(n1007), .B0(R14[22]), .B1(n1025), .C0(
        R13[22]), .C1(n1012), .Y(n575) );
  AOI22X1 U172 ( .A0(R15[22]), .A1(n1034), .B0(data_out_1[124]), .B1(n1024), 
        .Y(n574) );
  NAND2X1 U173 ( .A(n572), .B(n573), .Y(n842) );
  AOI222X1 U174 ( .A0(R12[23]), .A1(n1007), .B0(R14[23]), .B1(n1025), .C0(
        R13[23]), .C1(n1012), .Y(n573) );
  AOI22X1 U175 ( .A0(R15[23]), .A1(n1037), .B0(data_out_1[125]), .B1(n1024), 
        .Y(n572) );
  NAND2X1 U176 ( .A(n570), .B(n571), .Y(n841) );
  AOI222X1 U177 ( .A0(R12[24]), .A1(n1007), .B0(R14[24]), .B1(n1025), .C0(
        R13[24]), .C1(n1012), .Y(n571) );
  AOI22X1 U178 ( .A0(R15[24]), .A1(n1035), .B0(data_out_1[126]), .B1(n1024), 
        .Y(n570) );
  NAND2X1 U179 ( .A(n568), .B(n569), .Y(n840) );
  AOI222X1 U180 ( .A0(R12[25]), .A1(n1007), .B0(R14[25]), .B1(n1025), .C0(
        R13[25]), .C1(n1012), .Y(n569) );
  AOI22X1 U181 ( .A0(R15[25]), .A1(n1030), .B0(data_out_1[127]), .B1(n1024), 
        .Y(n568) );
  NAND2X1 U182 ( .A(n566), .B(n567), .Y(n839) );
  AOI222X1 U183 ( .A0(R12[26]), .A1(n1007), .B0(R14[26]), .B1(n1025), .C0(
        R13[26]), .C1(n1012), .Y(n567) );
  AOI22X1 U184 ( .A0(R15[26]), .A1(n1032), .B0(data_out_1[128]), .B1(n1024), 
        .Y(n566) );
  NAND2X1 U185 ( .A(n564), .B(n565), .Y(n838) );
  AOI222X1 U186 ( .A0(R12[27]), .A1(n1007), .B0(R14[27]), .B1(n1025), .C0(
        R13[27]), .C1(n1012), .Y(n565) );
  AOI22X1 U187 ( .A0(R15[27]), .A1(n1034), .B0(data_out_1[129]), .B1(n1024), 
        .Y(n564) );
  NAND2X1 U188 ( .A(n562), .B(n563), .Y(n837) );
  AOI222X1 U189 ( .A0(R12[28]), .A1(n1007), .B0(R14[28]), .B1(n1025), .C0(
        R13[28]), .C1(n1012), .Y(n563) );
  AOI22X1 U190 ( .A0(R15[28]), .A1(n1037), .B0(data_out_1[130]), .B1(n1024), 
        .Y(n562) );
  NAND2X1 U191 ( .A(n560), .B(n561), .Y(n836) );
  AOI222X1 U192 ( .A0(R12[29]), .A1(n1007), .B0(R14[29]), .B1(n1025), .C0(
        R13[29]), .C1(n1012), .Y(n561) );
  AOI22X1 U193 ( .A0(R15[29]), .A1(n1035), .B0(data_out_1[131]), .B1(n1024), 
        .Y(n560) );
  NAND2X1 U194 ( .A(n686), .B(n687), .Y(n899) );
  AOI222X1 U195 ( .A0(R8[0]), .A1(n1008), .B0(R10[0]), .B1(n1026), .C0(R9[0]), 
        .C1(n1014), .Y(n687) );
  AOI22X1 U196 ( .A0(R11[0]), .A1(n1034), .B0(data_out_1[68]), .B1(n1020), .Y(
        n686) );
  NAND2X1 U197 ( .A(n684), .B(n685), .Y(n898) );
  AOI222X1 U198 ( .A0(R8[1]), .A1(n1008), .B0(R10[1]), .B1(n1026), .C0(R9[1]), 
        .C1(n1015), .Y(n685) );
  AOI22X1 U199 ( .A0(R11[1]), .A1(n1034), .B0(data_out_1[69]), .B1(n1020), .Y(
        n684) );
  NAND2X1 U200 ( .A(n682), .B(n683), .Y(n897) );
  AOI222X1 U201 ( .A0(R8[2]), .A1(n1008), .B0(R10[2]), .B1(n1026), .C0(R9[2]), 
        .C1(n1014), .Y(n683) );
  AOI22X1 U202 ( .A0(R11[2]), .A1(n1034), .B0(data_out_1[70]), .B1(n1020), .Y(
        n682) );
  NAND2X1 U203 ( .A(n680), .B(n681), .Y(n896) );
  AOI222X1 U204 ( .A0(R8[3]), .A1(n1008), .B0(R10[3]), .B1(n1026), .C0(R9[3]), 
        .C1(n1013), .Y(n681) );
  AOI22X1 U205 ( .A0(R11[3]), .A1(n1033), .B0(data_out_1[71]), .B1(n1020), .Y(
        n680) );
  NAND2X1 U206 ( .A(n678), .B(n679), .Y(n895) );
  AOI222X1 U207 ( .A0(R8[4]), .A1(n1008), .B0(R10[4]), .B1(n1026), .C0(R9[4]), 
        .C1(n1015), .Y(n679) );
  AOI22X1 U208 ( .A0(R11[4]), .A1(n1033), .B0(data_out_1[72]), .B1(n1021), .Y(
        n678) );
  NAND2X1 U209 ( .A(n676), .B(n677), .Y(n894) );
  AOI222X1 U210 ( .A0(R8[5]), .A1(n1008), .B0(R10[5]), .B1(n1026), .C0(R9[5]), 
        .C1(n1014), .Y(n677) );
  AOI22X1 U211 ( .A0(R11[5]), .A1(n1033), .B0(data_out_1[73]), .B1(n1021), .Y(
        n676) );
  NAND2X1 U212 ( .A(n674), .B(n675), .Y(n893) );
  AOI222X1 U213 ( .A0(R8[6]), .A1(n1008), .B0(R10[6]), .B1(n1026), .C0(R9[6]), 
        .C1(n1014), .Y(n675) );
  AOI22X1 U214 ( .A0(R11[6]), .A1(n1033), .B0(data_out_1[74]), .B1(n1021), .Y(
        n674) );
  NAND2X1 U215 ( .A(n672), .B(n673), .Y(n892) );
  AOI222X1 U216 ( .A0(R8[7]), .A1(n1008), .B0(R10[7]), .B1(n1026), .C0(R9[7]), 
        .C1(n1015), .Y(n673) );
  AOI22X1 U217 ( .A0(R11[7]), .A1(n1033), .B0(data_out_1[75]), .B1(n1021), .Y(
        n672) );
  NAND2X1 U218 ( .A(n670), .B(n671), .Y(n891) );
  AOI222X1 U219 ( .A0(R8[8]), .A1(n1008), .B0(R10[8]), .B1(n1026), .C0(R9[8]), 
        .C1(n1014), .Y(n671) );
  AOI22X1 U220 ( .A0(R11[8]), .A1(n1033), .B0(data_out_1[76]), .B1(n1021), .Y(
        n670) );
  NAND2X1 U221 ( .A(n668), .B(n669), .Y(n890) );
  AOI222X1 U222 ( .A0(R8[9]), .A1(n1008), .B0(R10[9]), .B1(n1026), .C0(R9[9]), 
        .C1(n1015), .Y(n669) );
  AOI22X1 U223 ( .A0(R11[9]), .A1(n1033), .B0(data_out_1[77]), .B1(n1021), .Y(
        n668) );
  NAND2X1 U224 ( .A(n666), .B(n667), .Y(n889) );
  AOI222X1 U225 ( .A0(R8[10]), .A1(n1008), .B0(R10[10]), .B1(n1026), .C0(
        R9[10]), .C1(n1015), .Y(n667) );
  AOI22X1 U226 ( .A0(R11[10]), .A1(n1033), .B0(data_out_1[78]), .B1(n1021), 
        .Y(n666) );
  NAND2X1 U227 ( .A(n664), .B(n665), .Y(n888) );
  AOI222X1 U228 ( .A0(R8[11]), .A1(n1008), .B0(R10[11]), .B1(n1026), .C0(
        R9[11]), .C1(n1014), .Y(n665) );
  AOI22X1 U229 ( .A0(R11[11]), .A1(n1033), .B0(data_out_1[79]), .B1(n1021), 
        .Y(n664) );
  NAND2X1 U230 ( .A(n662), .B(n663), .Y(n887) );
  AOI222X1 U231 ( .A0(R8[12]), .A1(n1008), .B0(R10[12]), .B1(n1026), .C0(
        R9[12]), .C1(n1013), .Y(n663) );
  AOI22X1 U232 ( .A0(R11[12]), .A1(n1033), .B0(data_out_1[80]), .B1(n1021), 
        .Y(n662) );
  NAND2X1 U233 ( .A(n660), .B(n661), .Y(n886) );
  AOI222X1 U234 ( .A0(R8[13]), .A1(n1008), .B0(R10[13]), .B1(n1026), .C0(
        R9[13]), .C1(n1015), .Y(n661) );
  AOI22X1 U235 ( .A0(R11[13]), .A1(n1033), .B0(data_out_1[81]), .B1(n1021), 
        .Y(n660) );
  NAND2X1 U236 ( .A(n658), .B(n659), .Y(n885) );
  AOI222X1 U237 ( .A0(R8[14]), .A1(n1008), .B0(R10[14]), .B1(n1026), .C0(
        R9[14]), .C1(n1015), .Y(n659) );
  AOI22X1 U238 ( .A0(R11[14]), .A1(n1033), .B0(data_out_1[82]), .B1(n1021), 
        .Y(n658) );
  NAND2X1 U239 ( .A(n656), .B(n657), .Y(n884) );
  AOI222X1 U240 ( .A0(R8[15]), .A1(n1009), .B0(R10[15]), .B1(n1025), .C0(
        R9[15]), .C1(n1013), .Y(n657) );
  AOI22X1 U241 ( .A0(R11[15]), .A1(n1033), .B0(data_out_1[83]), .B1(n1021), 
        .Y(n656) );
  NAND2X1 U242 ( .A(n654), .B(n655), .Y(n883) );
  AOI222X1 U243 ( .A0(R8[16]), .A1(n1009), .B0(R10[16]), .B1(n1028), .C0(
        R9[16]), .C1(n1015), .Y(n655) );
  AOI22XL U244 ( .A0(R11[16]), .A1(n1032), .B0(data_out_1[84]), .B1(n1021), 
        .Y(n654) );
  NAND2X1 U245 ( .A(n652), .B(n653), .Y(n882) );
  AOI222X1 U246 ( .A0(R8[17]), .A1(n1010), .B0(R10[17]), .B1(n1027), .C0(
        R9[17]), .C1(n1014), .Y(n653) );
  AOI22X1 U247 ( .A0(R11[17]), .A1(n1032), .B0(data_out_1[85]), .B1(n1024), 
        .Y(n652) );
  NAND2X1 U248 ( .A(n650), .B(n651), .Y(n881) );
  AOI222X1 U249 ( .A0(R8[18]), .A1(n1011), .B0(R10[18]), .B1(n1028), .C0(
        R9[18]), .C1(n1015), .Y(n651) );
  AOI22X1 U250 ( .A0(R11[18]), .A1(n1032), .B0(data_out_1[86]), .B1(n1021), 
        .Y(n650) );
  NAND2X1 U251 ( .A(n648), .B(n649), .Y(n880) );
  AOI222X1 U252 ( .A0(R8[19]), .A1(n1008), .B0(R10[19]), .B1(n1026), .C0(
        R9[19]), .C1(n1013), .Y(n649) );
  AOI22X1 U253 ( .A0(R11[19]), .A1(n1032), .B0(data_out_1[87]), .B1(n1024), 
        .Y(n648) );
  NAND2X1 U254 ( .A(n646), .B(n647), .Y(n879) );
  AOI222X1 U255 ( .A0(R8[20]), .A1(n1009), .B0(R10[20]), .B1(n1025), .C0(
        R9[20]), .C1(n1014), .Y(n647) );
  AOI22X1 U256 ( .A0(R11[20]), .A1(n1032), .B0(data_out_1[88]), .B1(n1023), 
        .Y(n646) );
  NAND2X1 U257 ( .A(n644), .B(n645), .Y(n878) );
  AOI222X1 U258 ( .A0(R8[21]), .A1(n1010), .B0(R10[21]), .B1(n1027), .C0(
        R9[21]), .C1(n1015), .Y(n645) );
  AOI22X1 U259 ( .A0(R11[21]), .A1(n1032), .B0(data_out_1[89]), .B1(n1024), 
        .Y(n644) );
  NAND2X1 U260 ( .A(n642), .B(n643), .Y(n877) );
  AOI222X1 U261 ( .A0(R8[22]), .A1(n1011), .B0(R10[22]), .B1(n1027), .C0(
        R9[22]), .C1(n1013), .Y(n643) );
  AOI22X1 U262 ( .A0(R11[22]), .A1(n1032), .B0(data_out_1[90]), .B1(n1021), 
        .Y(n642) );
  NAND2X1 U263 ( .A(n640), .B(n641), .Y(n876) );
  AOI222X1 U264 ( .A0(R8[23]), .A1(n1008), .B0(R10[23]), .B1(n1026), .C0(
        R9[23]), .C1(n1014), .Y(n641) );
  AOI22X1 U265 ( .A0(R11[23]), .A1(n1032), .B0(data_out_1[91]), .B1(n1024), 
        .Y(n640) );
  NAND2X1 U266 ( .A(n638), .B(n639), .Y(n875) );
  AOI222X1 U267 ( .A0(R8[24]), .A1(n1009), .B0(R10[24]), .B1(N230), .C0(R9[24]), .C1(n1015), .Y(n639) );
  AOI22X1 U268 ( .A0(R11[24]), .A1(n1032), .B0(data_out_1[92]), .B1(n1022), 
        .Y(n638) );
  NAND2X1 U269 ( .A(n636), .B(n637), .Y(n874) );
  AOI222X1 U270 ( .A0(R8[25]), .A1(n1010), .B0(R10[25]), .B1(n1027), .C0(
        R9[25]), .C1(n1013), .Y(n637) );
  AOI22X1 U271 ( .A0(R11[25]), .A1(n1032), .B0(data_out_1[93]), .B1(n1021), 
        .Y(n636) );
  NAND2X1 U272 ( .A(n634), .B(n635), .Y(n873) );
  AOI222X1 U273 ( .A0(R8[26]), .A1(n1011), .B0(R10[26]), .B1(n1026), .C0(
        R9[26]), .C1(n1014), .Y(n635) );
  AOI22X1 U274 ( .A0(R11[26]), .A1(n1032), .B0(data_out_1[94]), .B1(n1024), 
        .Y(n634) );
  NAND2X1 U275 ( .A(n632), .B(n633), .Y(n872) );
  AOI222X1 U276 ( .A0(R8[27]), .A1(n1008), .B0(R10[27]), .B1(n1026), .C0(
        R9[27]), .C1(n1015), .Y(n633) );
  AOI22X1 U277 ( .A0(R11[27]), .A1(n1032), .B0(data_out_1[95]), .B1(n1021), 
        .Y(n632) );
  NAND2X1 U278 ( .A(n630), .B(n631), .Y(n871) );
  AOI222X1 U279 ( .A0(R8[28]), .A1(n1009), .B0(R10[28]), .B1(N230), .C0(R9[28]), .C1(n1013), .Y(n631) );
  AOI22X1 U280 ( .A0(R11[28]), .A1(n1032), .B0(data_out_1[96]), .B1(n1022), 
        .Y(n630) );
  NAND2X1 U281 ( .A(n628), .B(n629), .Y(n870) );
  AOI222X1 U282 ( .A0(R8[29]), .A1(n1010), .B0(R10[29]), .B1(n1027), .C0(
        R9[29]), .C1(n1014), .Y(n629) );
  AOI22X1 U283 ( .A0(R11[29]), .A1(n1031), .B0(data_out_1[97]), .B1(n1022), 
        .Y(n628) );
  NAND2X1 U284 ( .A(n626), .B(n627), .Y(n869) );
  AOI222X1 U285 ( .A0(R8[30]), .A1(n1011), .B0(R10[30]), .B1(n1026), .C0(
        R9[30]), .C1(n1015), .Y(n627) );
  AOI22X1 U286 ( .A0(R11[30]), .A1(n1031), .B0(data_out_1[98]), .B1(n1022), 
        .Y(n626) );
  NAND2X1 U287 ( .A(n624), .B(n625), .Y(n868) );
  AOI222X1 U288 ( .A0(R8[31]), .A1(n1008), .B0(R10[31]), .B1(n1026), .C0(
        R9[31]), .C1(n1013), .Y(n625) );
  AOI22X1 U289 ( .A0(R11[31]), .A1(n1031), .B0(data_out_1[99]), .B1(n1022), 
        .Y(n624) );
  NAND2X1 U290 ( .A(n622), .B(n623), .Y(n867) );
  AOI222X1 U291 ( .A0(R8[32]), .A1(n1008), .B0(R10[32]), .B1(n1028), .C0(
        R9[32]), .C1(n1013), .Y(n623) );
  AOI22X1 U292 ( .A0(R11[32]), .A1(n1031), .B0(data_out_1[100]), .B1(n1022), 
        .Y(n622) );
  NAND2X1 U293 ( .A(n620), .B(n621), .Y(n866) );
  AOI222X1 U294 ( .A0(R8[33]), .A1(n1010), .B0(R10[33]), .B1(n1027), .C0(
        R9[33]), .C1(n1013), .Y(n621) );
  AOI22XL U295 ( .A0(R11[33]), .A1(n1031), .B0(data_out_1[101]), .B1(n1022), 
        .Y(n620) );
  NAND2X1 U296 ( .A(n754), .B(n755), .Y(n933) );
  AOI222X1 U297 ( .A0(R4[0]), .A1(n1010), .B0(R6[0]), .B1(n1028), .C0(R5[0]), 
        .C1(n1014), .Y(n755) );
  AOI22X1 U298 ( .A0(R7[0]), .A1(n1036), .B0(data_out_1[34]), .B1(n1020), .Y(
        n754) );
  NAND2X1 U299 ( .A(n752), .B(n753), .Y(n932) );
  AOI222X1 U300 ( .A0(R4[1]), .A1(n1010), .B0(R6[1]), .B1(n1027), .C0(R5[1]), 
        .C1(n1014), .Y(n753) );
  AOI22X1 U301 ( .A0(R7[1]), .A1(n1036), .B0(data_out_1[35]), .B1(n1020), .Y(
        n752) );
  NAND2X1 U302 ( .A(n750), .B(n751), .Y(n931) );
  AOI222X1 U303 ( .A0(R4[2]), .A1(n1010), .B0(R6[2]), .B1(n1026), .C0(R5[2]), 
        .C1(n1014), .Y(n751) );
  AOI22X1 U304 ( .A0(R7[2]), .A1(n1036), .B0(data_out_1[36]), .B1(n1018), .Y(
        n750) );
  NAND2X1 U305 ( .A(n748), .B(n749), .Y(n930) );
  AOI222X1 U306 ( .A0(R4[3]), .A1(n1010), .B0(R6[3]), .B1(n1028), .C0(R5[3]), 
        .C1(n1014), .Y(n749) );
  AOI22X1 U307 ( .A0(R7[3]), .A1(n1036), .B0(data_out_1[37]), .B1(n1018), .Y(
        n748) );
  NAND2X1 U308 ( .A(n746), .B(n747), .Y(n929) );
  AOI222X1 U309 ( .A0(R4[4]), .A1(n1010), .B0(R6[4]), .B1(n1027), .C0(R5[4]), 
        .C1(n1014), .Y(n747) );
  AOI22X1 U310 ( .A0(R7[4]), .A1(n1036), .B0(data_out_1[38]), .B1(n1018), .Y(
        n746) );
  NAND2X1 U311 ( .A(n744), .B(n745), .Y(n928) );
  AOI222X1 U312 ( .A0(R4[5]), .A1(n1010), .B0(R6[5]), .B1(n1026), .C0(R5[5]), 
        .C1(n1014), .Y(n745) );
  AOI22X1 U313 ( .A0(R7[5]), .A1(n1036), .B0(data_out_1[39]), .B1(n1018), .Y(
        n744) );
  NAND2X1 U314 ( .A(n742), .B(n743), .Y(n927) );
  AOI222X1 U315 ( .A0(R4[6]), .A1(n1010), .B0(R6[6]), .B1(n1028), .C0(R5[6]), 
        .C1(n1014), .Y(n743) );
  AOI22X1 U316 ( .A0(R7[6]), .A1(n1036), .B0(data_out_1[40]), .B1(n1018), .Y(
        n742) );
  NAND2X1 U317 ( .A(n740), .B(n741), .Y(n926) );
  AOI222X1 U318 ( .A0(R4[7]), .A1(n1010), .B0(R6[7]), .B1(n1027), .C0(R5[7]), 
        .C1(n1014), .Y(n741) );
  AOI22X1 U319 ( .A0(R7[7]), .A1(n1036), .B0(data_out_1[41]), .B1(n1018), .Y(
        n740) );
  NAND2X1 U320 ( .A(n738), .B(n739), .Y(n925) );
  AOI222X1 U321 ( .A0(R4[8]), .A1(n1010), .B0(R6[8]), .B1(n1026), .C0(R5[8]), 
        .C1(n1014), .Y(n739) );
  AOI22X1 U322 ( .A0(R7[8]), .A1(n1036), .B0(data_out_1[42]), .B1(n1018), .Y(
        n738) );
  NAND2X1 U323 ( .A(n736), .B(n737), .Y(n924) );
  AOI222X1 U324 ( .A0(R4[9]), .A1(n1010), .B0(R6[9]), .B1(n1028), .C0(R5[9]), 
        .C1(n1014), .Y(n737) );
  AOI22X1 U325 ( .A0(R7[9]), .A1(n1036), .B0(data_out_1[43]), .B1(n1018), .Y(
        n736) );
  NAND2X1 U326 ( .A(n734), .B(n735), .Y(n923) );
  AOI222X1 U327 ( .A0(R4[10]), .A1(n1010), .B0(R6[10]), .B1(n1027), .C0(R5[10]), .C1(n1014), .Y(n735) );
  AOI22X1 U328 ( .A0(R7[10]), .A1(n1036), .B0(data_out_1[44]), .B1(n1018), .Y(
        n734) );
  NAND2X1 U329 ( .A(n732), .B(n733), .Y(n922) );
  AOI222X1 U330 ( .A0(R4[11]), .A1(n1010), .B0(R6[11]), .B1(n1026), .C0(R5[11]), .C1(n1014), .Y(n733) );
  AOI22X1 U331 ( .A0(R7[11]), .A1(n1036), .B0(data_out_1[45]), .B1(n1018), .Y(
        n732) );
  NAND2X1 U332 ( .A(n730), .B(n731), .Y(n921) );
  AOI222X1 U333 ( .A0(R4[12]), .A1(n1010), .B0(R6[12]), .B1(n1028), .C0(R5[12]), .C1(n1014), .Y(n731) );
  AOI22X1 U334 ( .A0(R7[12]), .A1(n1035), .B0(data_out_1[46]), .B1(n1018), .Y(
        n730) );
  NAND2X1 U335 ( .A(n728), .B(n729), .Y(n920) );
  AOI222X1 U336 ( .A0(R4[13]), .A1(n1010), .B0(R6[13]), .B1(n1026), .C0(R5[13]), .C1(n1013), .Y(n729) );
  AOI22X1 U337 ( .A0(R7[13]), .A1(n1035), .B0(data_out_1[47]), .B1(n1018), .Y(
        n728) );
  NAND2X1 U338 ( .A(n726), .B(n727), .Y(n919) );
  AOI222X1 U339 ( .A0(R4[14]), .A1(n1009), .B0(R6[14]), .B1(n1026), .C0(R5[14]), .C1(n1013), .Y(n727) );
  AOI22X1 U340 ( .A0(R7[14]), .A1(n1035), .B0(data_out_1[48]), .B1(n1019), .Y(
        n726) );
  NAND2X1 U341 ( .A(n724), .B(n725), .Y(n918) );
  AOI222X1 U342 ( .A0(R4[15]), .A1(n1009), .B0(R6[15]), .B1(n1027), .C0(R5[15]), .C1(n1013), .Y(n725) );
  AOI22X1 U343 ( .A0(R7[15]), .A1(n1035), .B0(data_out_1[49]), .B1(n1019), .Y(
        n724) );
  NAND2X1 U344 ( .A(n722), .B(n723), .Y(n917) );
  AOI222X1 U345 ( .A0(R4[16]), .A1(n1009), .B0(R6[16]), .B1(n1026), .C0(R5[16]), .C1(n1013), .Y(n723) );
  AOI22XL U346 ( .A0(R7[16]), .A1(n1035), .B0(data_out_1[50]), .B1(n1019), .Y(
        n722) );
  NAND2X1 U347 ( .A(n720), .B(n721), .Y(n916) );
  AOI222X1 U348 ( .A0(R4[17]), .A1(n1009), .B0(R6[17]), .B1(n1028), .C0(R5[17]), .C1(n1013), .Y(n721) );
  AOI22X1 U349 ( .A0(R7[17]), .A1(n1035), .B0(data_out_1[51]), .B1(n1019), .Y(
        n720) );
  NAND2X1 U350 ( .A(n718), .B(n719), .Y(n915) );
  AOI222X1 U351 ( .A0(R4[18]), .A1(n1009), .B0(R6[18]), .B1(n1026), .C0(R5[18]), .C1(n1013), .Y(n719) );
  AOI22X1 U352 ( .A0(R7[18]), .A1(n1035), .B0(data_out_1[52]), .B1(n1019), .Y(
        n718) );
  NAND2X1 U353 ( .A(n716), .B(n717), .Y(n914) );
  AOI222X1 U354 ( .A0(R4[19]), .A1(n1009), .B0(R6[19]), .B1(n1028), .C0(R5[19]), .C1(n1013), .Y(n717) );
  AOI22X1 U355 ( .A0(R7[19]), .A1(n1035), .B0(data_out_1[53]), .B1(n1019), .Y(
        n716) );
  NAND2X1 U356 ( .A(n714), .B(n715), .Y(n913) );
  AOI222X1 U357 ( .A0(R4[20]), .A1(n1009), .B0(R6[20]), .B1(n1027), .C0(R5[20]), .C1(n1013), .Y(n715) );
  AOI22X1 U358 ( .A0(R7[20]), .A1(n1035), .B0(data_out_1[54]), .B1(n1019), .Y(
        n714) );
  NAND2X1 U359 ( .A(n712), .B(n713), .Y(n912) );
  AOI222X1 U360 ( .A0(R4[21]), .A1(n1009), .B0(R6[21]), .B1(n1027), .C0(R5[21]), .C1(n1013), .Y(n713) );
  AOI22X1 U361 ( .A0(R7[21]), .A1(n1035), .B0(data_out_1[55]), .B1(n1019), .Y(
        n712) );
  NAND2X1 U362 ( .A(n710), .B(n711), .Y(n911) );
  AOI222X1 U363 ( .A0(R4[22]), .A1(n1009), .B0(R6[22]), .B1(n1026), .C0(R5[22]), .C1(n1013), .Y(n711) );
  AOI22X1 U364 ( .A0(R7[22]), .A1(n1035), .B0(data_out_1[56]), .B1(n1019), .Y(
        n710) );
  NAND2X1 U365 ( .A(n708), .B(n709), .Y(n910) );
  AOI222X1 U366 ( .A0(R4[23]), .A1(n1009), .B0(R6[23]), .B1(n1028), .C0(R5[23]), .C1(n1013), .Y(n709) );
  AOI22X1 U367 ( .A0(R7[23]), .A1(n1035), .B0(data_out_1[57]), .B1(n1019), .Y(
        n708) );
  NAND2X1 U368 ( .A(n706), .B(n707), .Y(n909) );
  AOI222X1 U369 ( .A0(R4[24]), .A1(n1009), .B0(R6[24]), .B1(n1027), .C0(R5[24]), .C1(n1013), .Y(n707) );
  AOI22X1 U370 ( .A0(R7[24]), .A1(n1034), .B0(data_out_1[58]), .B1(n1019), .Y(
        n706) );
  NAND2X1 U371 ( .A(n704), .B(n705), .Y(n908) );
  AOI222X1 U372 ( .A0(R4[25]), .A1(n1009), .B0(R6[25]), .B1(n1026), .C0(R5[25]), .C1(n1013), .Y(n705) );
  AOI22X1 U373 ( .A0(R7[25]), .A1(n1034), .B0(data_out_1[59]), .B1(n1019), .Y(
        n704) );
  NAND2X1 U374 ( .A(n702), .B(n703), .Y(n907) );
  AOI222X1 U375 ( .A0(R4[26]), .A1(n1009), .B0(R6[26]), .B1(n1026), .C0(R5[26]), .C1(n1013), .Y(n703) );
  AOI22X1 U376 ( .A0(R7[26]), .A1(n1034), .B0(data_out_1[60]), .B1(n1020), .Y(
        n702) );
  NAND2X1 U377 ( .A(n700), .B(n701), .Y(n906) );
  AOI222X1 U378 ( .A0(R4[27]), .A1(n1009), .B0(R6[27]), .B1(n1028), .C0(R5[27]), .C1(n1013), .Y(n701) );
  AOI22X1 U379 ( .A0(R7[27]), .A1(n1034), .B0(data_out_1[61]), .B1(n1020), .Y(
        n700) );
  NAND2X1 U380 ( .A(n698), .B(n699), .Y(n905) );
  AOI222X1 U381 ( .A0(R4[28]), .A1(n1009), .B0(R6[28]), .B1(n1027), .C0(R5[28]), .C1(n1013), .Y(n699) );
  AOI22X1 U382 ( .A0(R7[28]), .A1(n1034), .B0(data_out_1[62]), .B1(n1020), .Y(
        n698) );
  NAND2X1 U383 ( .A(n696), .B(n697), .Y(n904) );
  AOI222X1 U384 ( .A0(R4[29]), .A1(n1009), .B0(R6[29]), .B1(n1026), .C0(R5[29]), .C1(n1014), .Y(n697) );
  AOI22X1 U385 ( .A0(R7[29]), .A1(n1034), .B0(data_out_1[63]), .B1(n1020), .Y(
        n696) );
  NAND2X1 U386 ( .A(n694), .B(n695), .Y(n903) );
  AOI222X1 U387 ( .A0(R4[30]), .A1(n1009), .B0(R6[30]), .B1(n1026), .C0(R5[30]), .C1(n1014), .Y(n695) );
  AOI22X1 U388 ( .A0(R7[30]), .A1(n1034), .B0(data_out_1[64]), .B1(n1020), .Y(
        n694) );
  NAND2X1 U389 ( .A(n692), .B(n693), .Y(n902) );
  AOI222X1 U390 ( .A0(R4[31]), .A1(n1008), .B0(R6[31]), .B1(n1026), .C0(R5[31]), .C1(n1014), .Y(n693) );
  AOI22X1 U391 ( .A0(R7[31]), .A1(n1034), .B0(data_out_1[65]), .B1(n1020), .Y(
        n692) );
  NAND2X1 U392 ( .A(n690), .B(n691), .Y(n901) );
  AOI222X1 U393 ( .A0(R4[32]), .A1(n1008), .B0(R6[32]), .B1(n1026), .C0(R5[32]), .C1(n1015), .Y(n691) );
  AOI22X1 U394 ( .A0(R7[32]), .A1(n1034), .B0(data_out_1[66]), .B1(n1020), .Y(
        n690) );
  NAND2X1 U395 ( .A(n688), .B(n689), .Y(n900) );
  AOI222X1 U396 ( .A0(R4[33]), .A1(n1008), .B0(R6[33]), .B1(n1026), .C0(R5[33]), .C1(n1014), .Y(n689) );
  AOI22XL U397 ( .A0(R7[33]), .A1(n1034), .B0(data_out_1[67]), .B1(n1020), .Y(
        n688) );
  NAND2X1 U398 ( .A(n822), .B(n823), .Y(n967) );
  AOI222X1 U399 ( .A0(R0[0]), .A1(n1009), .B0(R2[0]), .B1(n1027), .C0(R1[0]), 
        .C1(n1015), .Y(n823) );
  NAND2X1 U400 ( .A(n820), .B(n821), .Y(n966) );
  AOI222X1 U401 ( .A0(R0[1]), .A1(n1010), .B0(R2[1]), .B1(n1026), .C0(R1[1]), 
        .C1(n1015), .Y(n821) );
  NAND2X1 U402 ( .A(n818), .B(n819), .Y(n965) );
  AOI222X1 U403 ( .A0(R0[2]), .A1(n1011), .B0(R2[2]), .B1(n1027), .C0(R1[2]), 
        .C1(n1015), .Y(n819) );
  NAND2X1 U404 ( .A(n816), .B(n817), .Y(n964) );
  AOI222X1 U405 ( .A0(R0[3]), .A1(n1009), .B0(R2[3]), .B1(n1026), .C0(R1[3]), 
        .C1(n1015), .Y(n817) );
  NAND2X1 U406 ( .A(n814), .B(n815), .Y(n963) );
  AOI222X1 U407 ( .A0(R0[4]), .A1(n1011), .B0(R2[4]), .B1(n1026), .C0(R1[4]), 
        .C1(n1015), .Y(n815) );
  AOI22X1 U408 ( .A0(R3[4]), .A1(n1039), .B0(data_out_1[4]), .B1(n1022), .Y(
        n814) );
  NAND2X1 U409 ( .A(n812), .B(n813), .Y(n962) );
  AOI222X1 U410 ( .A0(R0[5]), .A1(n1011), .B0(R2[5]), .B1(n1027), .C0(R1[5]), 
        .C1(n1015), .Y(n813) );
  AOI22X1 U411 ( .A0(R3[5]), .A1(n1039), .B0(data_out_1[5]), .B1(n1018), .Y(
        n812) );
  NAND2X1 U412 ( .A(n810), .B(n811), .Y(n961) );
  AOI222X1 U413 ( .A0(R0[6]), .A1(n1009), .B0(R2[6]), .B1(n1027), .C0(R1[6]), 
        .C1(n1015), .Y(n811) );
  AOI22X1 U414 ( .A0(R3[6]), .A1(n1039), .B0(data_out_1[6]), .B1(n1017), .Y(
        n810) );
  NAND2X1 U415 ( .A(n808), .B(n809), .Y(n960) );
  AOI222X1 U416 ( .A0(R0[7]), .A1(n1010), .B0(R2[7]), .B1(n1026), .C0(R1[7]), 
        .C1(n1015), .Y(n809) );
  NAND2X1 U417 ( .A(n806), .B(n807), .Y(n959) );
  AOI222X1 U418 ( .A0(R0[8]), .A1(n1010), .B0(R2[8]), .B1(n1027), .C0(R1[8]), 
        .C1(n1015), .Y(n807) );
  AOI22X1 U419 ( .A0(R3[8]), .A1(n1038), .B0(data_out_1[8]), .B1(n1023), .Y(
        n806) );
  NAND2X1 U420 ( .A(n804), .B(n805), .Y(n958) );
  AOI222X1 U421 ( .A0(R0[9]), .A1(n1011), .B0(R2[9]), .B1(n1026), .C0(R1[9]), 
        .C1(n1015), .Y(n805) );
  AOI22X1 U422 ( .A0(R3[9]), .A1(n1038), .B0(data_out_1[9]), .B1(n1018), .Y(
        n804) );
  NAND2X1 U423 ( .A(n802), .B(n803), .Y(n957) );
  AOI222X1 U424 ( .A0(R0[10]), .A1(n1009), .B0(R2[10]), .B1(N230), .C0(R1[10]), 
        .C1(n1015), .Y(n803) );
  AOI22X1 U425 ( .A0(R3[10]), .A1(n1038), .B0(data_out_1[10]), .B1(n1017), .Y(
        n802) );
  NAND2X1 U426 ( .A(n800), .B(n801), .Y(n956) );
  AOI222X1 U427 ( .A0(R0[11]), .A1(n1010), .B0(R2[11]), .B1(n1027), .C0(R1[11]), .C1(n1014), .Y(n801) );
  AOI22X1 U428 ( .A0(R3[11]), .A1(n1038), .B0(data_out_1[11]), .B1(n1022), .Y(
        n800) );
  NAND2X1 U429 ( .A(n798), .B(n799), .Y(n955) );
  AOI222X1 U430 ( .A0(R0[12]), .A1(n1011), .B0(R2[12]), .B1(n1027), .C0(R1[12]), .C1(n1014), .Y(n799) );
  AOI22X1 U431 ( .A0(R3[12]), .A1(n1038), .B0(data_out_1[12]), .B1(n1017), .Y(
        n798) );
  NAND2X1 U432 ( .A(n796), .B(n797), .Y(n954) );
  AOI222X1 U433 ( .A0(R0[13]), .A1(n1011), .B0(R2[13]), .B1(n1027), .C0(R1[13]), .C1(n1015), .Y(n797) );
  AOI22X1 U434 ( .A0(R3[13]), .A1(n1038), .B0(data_out_1[13]), .B1(n1017), .Y(
        n796) );
  NAND2X1 U435 ( .A(n794), .B(n795), .Y(n953) );
  AOI222X1 U436 ( .A0(R0[14]), .A1(n1011), .B0(R2[14]), .B1(n1027), .C0(R1[14]), .C1(n1014), .Y(n795) );
  AOI22X1 U437 ( .A0(R3[14]), .A1(n1038), .B0(data_out_1[14]), .B1(n1017), .Y(
        n794) );
  NAND2X1 U438 ( .A(n792), .B(n793), .Y(n952) );
  AOI222X1 U439 ( .A0(R0[15]), .A1(n1011), .B0(R2[15]), .B1(n1027), .C0(R1[15]), .C1(n1015), .Y(n793) );
  AOI22X1 U440 ( .A0(R3[15]), .A1(n1038), .B0(data_out_1[15]), .B1(n1017), .Y(
        n792) );
  NAND2X1 U441 ( .A(n790), .B(n791), .Y(n951) );
  AOI222X1 U442 ( .A0(R0[16]), .A1(n1011), .B0(R2[16]), .B1(n1027), .C0(R1[16]), .C1(n1014), .Y(n791) );
  AOI22X1 U443 ( .A0(R3[16]), .A1(n1038), .B0(data_out_1[16]), .B1(n1017), .Y(
        n790) );
  NAND2X1 U444 ( .A(n788), .B(n789), .Y(n950) );
  AOI222X1 U445 ( .A0(R0[17]), .A1(n1011), .B0(R2[17]), .B1(n1027), .C0(R1[17]), .C1(n1015), .Y(n789) );
  NAND2X1 U446 ( .A(n786), .B(n787), .Y(n949) );
  AOI222X1 U447 ( .A0(R0[18]), .A1(n1011), .B0(R2[18]), .B1(n1027), .C0(R1[18]), .C1(n1015), .Y(n787) );
  NAND2X1 U448 ( .A(n784), .B(n785), .Y(n948) );
  AOI222X1 U449 ( .A0(R0[19]), .A1(n1011), .B0(R2[19]), .B1(n1027), .C0(R1[19]), .C1(n1013), .Y(n785) );
  NAND2X1 U450 ( .A(n782), .B(n783), .Y(n947) );
  AOI222X1 U451 ( .A0(R0[20]), .A1(n1011), .B0(R2[20]), .B1(n1027), .C0(R1[20]), .C1(n1014), .Y(n783) );
  NAND2X1 U452 ( .A(n780), .B(n781), .Y(n946) );
  AOI222X1 U453 ( .A0(R0[21]), .A1(n1011), .B0(R2[21]), .B1(n1027), .C0(R1[21]), .C1(n1013), .Y(n781) );
  AOI22X1 U454 ( .A0(R3[21]), .A1(n1037), .B0(data_out_1[21]), .B1(n1017), .Y(
        n780) );
  NAND2X1 U455 ( .A(n778), .B(n779), .Y(n945) );
  AOI222X1 U456 ( .A0(R0[22]), .A1(n1011), .B0(R2[22]), .B1(n1027), .C0(R1[22]), .C1(n1014), .Y(n779) );
  AOI22X1 U457 ( .A0(R3[22]), .A1(n1037), .B0(data_out_1[22]), .B1(n1017), .Y(
        n778) );
  NAND2X1 U458 ( .A(n776), .B(n777), .Y(n944) );
  AOI222X1 U459 ( .A0(R0[23]), .A1(n1011), .B0(R2[23]), .B1(n1027), .C0(R1[23]), .C1(n1015), .Y(n777) );
  AOI22X1 U460 ( .A0(R3[23]), .A1(n1037), .B0(data_out_1[23]), .B1(n1017), .Y(
        n776) );
  NAND2X1 U461 ( .A(n774), .B(n775), .Y(n943) );
  AOI222X1 U462 ( .A0(R0[24]), .A1(n1011), .B0(R2[24]), .B1(n1027), .C0(R1[24]), .C1(n1015), .Y(n775) );
  NAND2X1 U463 ( .A(n772), .B(n773), .Y(n942) );
  AOI222X1 U464 ( .A0(R0[25]), .A1(n1011), .B0(R2[25]), .B1(n1027), .C0(R1[25]), .C1(n1014), .Y(n773) );
  AOI22X1 U465 ( .A0(R3[25]), .A1(n1037), .B0(data_out_1[25]), .B1(n1020), .Y(
        n772) );
  NAND2X1 U466 ( .A(n770), .B(n771), .Y(n941) );
  AOI222X1 U467 ( .A0(R0[26]), .A1(n1011), .B0(R2[26]), .B1(n1027), .C0(R1[26]), .C1(n1014), .Y(n771) );
  AOI22X1 U468 ( .A0(R3[26]), .A1(n1037), .B0(data_out_1[26]), .B1(n1019), .Y(
        n770) );
  NAND2X1 U469 ( .A(n768), .B(n769), .Y(n940) );
  AOI222X1 U470 ( .A0(R0[27]), .A1(n1011), .B0(R2[27]), .B1(n1027), .C0(R1[27]), .C1(n1015), .Y(n769) );
  AOI22X1 U471 ( .A0(R3[27]), .A1(n1037), .B0(data_out_1[27]), .B1(n1020), .Y(
        n768) );
  NAND2X1 U472 ( .A(n766), .B(n767), .Y(n939) );
  AOI222X1 U473 ( .A0(R0[28]), .A1(n1011), .B0(R2[28]), .B1(n1027), .C0(R1[28]), .C1(n1015), .Y(n767) );
  AOI22X1 U474 ( .A0(R3[28]), .A1(n1037), .B0(data_out_1[28]), .B1(n1019), .Y(
        n766) );
  NAND2X1 U475 ( .A(n764), .B(n765), .Y(n938) );
  AOI222X1 U476 ( .A0(R0[29]), .A1(n1011), .B0(R2[29]), .B1(n1027), .C0(R1[29]), .C1(n1014), .Y(n765) );
  AOI22X1 U477 ( .A0(R3[29]), .A1(n1037), .B0(data_out_1[29]), .B1(n1020), .Y(
        n764) );
  NAND2X1 U478 ( .A(n762), .B(n763), .Y(n937) );
  AOI222X1 U479 ( .A0(R0[30]), .A1(n1010), .B0(R2[30]), .B1(n1027), .C0(R1[30]), .C1(n1014), .Y(n763) );
  AOI22X1 U480 ( .A0(R3[30]), .A1(n1037), .B0(data_out_1[30]), .B1(n1019), .Y(
        n762) );
  NAND2X1 U481 ( .A(n760), .B(n761), .Y(n936) );
  AOI222X1 U482 ( .A0(R0[31]), .A1(n1010), .B0(R2[31]), .B1(n1026), .C0(R1[31]), .C1(n1014), .Y(n761) );
  AOI22X1 U483 ( .A0(R3[31]), .A1(n1037), .B0(data_out_1[31]), .B1(n1023), .Y(
        n760) );
  NAND2X1 U484 ( .A(n758), .B(n759), .Y(n935) );
  AOI222X1 U485 ( .A0(R0[32]), .A1(n1010), .B0(R2[32]), .B1(n1028), .C0(R1[32]), .C1(n1014), .Y(n759) );
  AOI22X1 U486 ( .A0(R3[32]), .A1(n1037), .B0(data_out_1[32]), .B1(n1018), .Y(
        n758) );
  NAND2X1 U487 ( .A(n756), .B(n757), .Y(n934) );
  AOI222X1 U488 ( .A0(R0[33]), .A1(n1010), .B0(R2[33]), .B1(n1027), .C0(R1[33]), .C1(n1014), .Y(n757) );
  AOI22X1 U489 ( .A0(R3[33]), .A1(n1036), .B0(data_out_1[33]), .B1(n1019), .Y(
        n756) );
  NAND2X1 U490 ( .A(n558), .B(n559), .Y(n835) );
  AOI222X1 U491 ( .A0(R12[30]), .A1(n1007), .B0(R14[30]), .B1(n1025), .C0(
        R13[30]), .C1(n1012), .Y(n559) );
  AOI22X1 U492 ( .A0(R15[30]), .A1(n1038), .B0(data_out_1[132]), .B1(n1022), 
        .Y(n558) );
  NAND2X1 U493 ( .A(n556), .B(n557), .Y(n834) );
  AOI222X1 U494 ( .A0(R12[31]), .A1(n1007), .B0(R14[31]), .B1(n1025), .C0(
        R13[31]), .C1(n1012), .Y(n557) );
  AOI22X1 U495 ( .A0(R15[31]), .A1(n1031), .B0(data_out_1[133]), .B1(n1023), 
        .Y(n556) );
  NAND2X1 U496 ( .A(n554), .B(n555), .Y(n833) );
  AOI222X1 U497 ( .A0(R12[32]), .A1(n1007), .B0(R14[32]), .B1(n1025), .C0(
        R13[32]), .C1(n1012), .Y(n555) );
  AOI22X1 U498 ( .A0(R15[32]), .A1(n1030), .B0(data_out_1[134]), .B1(n1022), 
        .Y(n554) );
  NAND2X1 U499 ( .A(n551), .B(n552), .Y(n832) );
  AOI222X1 U500 ( .A0(R12[33]), .A1(n1009), .B0(R14[33]), .B1(n1026), .C0(
        R13[33]), .C1(n1013), .Y(n552) );
  AOI22XL U501 ( .A0(R15[33]), .A1(n1035), .B0(data_out_1[135]), .B1(n1023), 
        .Y(n551) );
  NAND2X1 U502 ( .A(counter[3]), .B(n1042), .Y(n827) );
  NAND2X1 U503 ( .A(counter[2]), .B(n1043), .Y(n829) );
  NOR2X1 U504 ( .A(n550), .B(n1041), .Y(n831) );
  OAI22X1 U505 ( .A0(n831), .A1(n1042), .B0(counter[2]), .B1(n826), .Y(N14) );
endmodule


module mux ( mux_flag, clk, rst_n, data_in_1, data_in_2, data_out, 
        data_in_3_33_, data_in_3_32_, data_in_3_31_, data_in_3_30_, 
        data_in_3_29_, data_in_3_28_, data_in_3_27_, data_in_3_26_, 
        data_in_3_25_, data_in_3_24_, data_in_3_23_, data_in_3_22_, 
        data_in_3_21_, data_in_3_20_, data_in_3_19_, data_in_3_18_, 
        data_in_3_17_, data_in_3_16_, data_in_3_15_, data_in_3_14_, 
        data_in_3_13_, data_in_3_12_, data_in_3_11_, data_in_3_10_, 
        data_in_3_9_, data_in_3_8_, data_in_3_7_, data_in_3_6_, data_in_3_5_, 
        data_in_3_4_, data_in_3_3_, data_in_3_2_, data_in_3_1_, data_in_3_0_
 );
  input [135:0] data_in_1;
  input [135:0] data_in_2;
  output [135:0] data_out;
  input mux_flag, clk, rst_n, data_in_3_33_, data_in_3_32_, data_in_3_31_,
         data_in_3_30_, data_in_3_29_, data_in_3_28_, data_in_3_27_,
         data_in_3_26_, data_in_3_25_, data_in_3_24_, data_in_3_23_,
         data_in_3_22_, data_in_3_21_, data_in_3_20_, data_in_3_19_,
         data_in_3_18_, data_in_3_17_, data_in_3_16_, data_in_3_15_,
         data_in_3_14_, data_in_3_13_, data_in_3_12_, data_in_3_11_,
         data_in_3_10_, data_in_3_9_, data_in_3_8_, data_in_3_7_, data_in_3_6_,
         data_in_3_5_, data_in_3_4_, data_in_3_3_, data_in_3_2_, data_in_3_1_,
         data_in_3_0_;
  wire   N6, N7, N8, n140, n141, n281, n282, n285, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n51, n52, n53,
         n54, n55, n56, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n283, n284, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n557, n558;
  wire   [3:1] counter;
  wire   [33:0] R4;
  wire   [32:0] R3;
  wire   [32:0] R2;
  wire   [33:0] R1;

  JKFFRX4 counter_reg_0_ ( .J(1'b1), .K(1'b1), .CK(clk), .RN(rst_n), .Q(n3), 
        .QN(n140) );
  DFFRHQX4 counter_reg_1_ ( .D(N6), .CK(clk), .RN(rst_n), .Q(counter[1]) );
  DFFRHQX4 counter_reg_2_ ( .D(N7), .CK(clk), .RN(rst_n), .Q(counter[2]) );
  DFFRHQX4 counter_reg_3_ ( .D(N8), .CK(clk), .RN(rst_n), .Q(counter[3]) );
  TLATXL R4_reg_16_ ( .G(n191), .D(data_in_3_16_), .QN(n7) );
  TLATXL R3_reg_16_ ( .G(n189), .D(data_in_3_16_), .QN(n54) );
  TLATXL R2_reg_16_ ( .G(n193), .D(data_in_3_16_), .Q(R2[16]) );
  TLATXL R1_reg_16_ ( .G(n186), .D(data_in_3_16_), .Q(R1[16]) );
  TLATXL R4_reg_13_ ( .G(n191), .D(data_in_3_13_), .Q(R4[13]) );
  TLATXL R3_reg_13_ ( .G(n189), .D(data_in_3_13_), .Q(R3[13]) );
  TLATXL R2_reg_13_ ( .G(n193), .D(data_in_3_13_), .Q(R2[13]) );
  TLATXL R1_reg_13_ ( .G(n186), .D(data_in_3_13_), .Q(R1[13]) );
  TLATXL R4_reg_14_ ( .G(n191), .D(data_in_3_14_), .Q(R4[14]) );
  TLATXL R3_reg_14_ ( .G(n189), .D(data_in_3_14_), .Q(R3[14]) );
  TLATXL R2_reg_14_ ( .G(n193), .D(data_in_3_14_), .Q(R2[14]) );
  TLATXL R1_reg_14_ ( .G(n186), .D(data_in_3_14_), .Q(R1[14]) );
  TLATXL R4_reg_33_ ( .G(n190), .D(data_in_3_33_), .Q(R4[33]) );
  TLATXL R2_reg_33_ ( .G(n192), .D(data_in_3_33_), .QN(n51) );
  TLATXL R1_reg_24_ ( .G(n186), .D(data_in_3_24_), .Q(R1[24]) );
  TLATXL R2_reg_32_ ( .G(n193), .D(data_in_3_32_), .Q(R2[32]) );
  TLATXL R2_reg_31_ ( .G(n192), .D(data_in_3_31_), .Q(R2[31]) );
  TLATXL R2_reg_30_ ( .G(n193), .D(data_in_3_30_), .Q(R2[30]) );
  TLATXL R2_reg_29_ ( .G(n192), .D(data_in_3_29_), .Q(R2[29]) );
  TLATXL R2_reg_28_ ( .G(n193), .D(data_in_3_28_), .Q(R2[28]) );
  TLATXL R2_reg_27_ ( .G(n192), .D(data_in_3_27_), .Q(R2[27]) );
  TLATXL R2_reg_26_ ( .G(n193), .D(data_in_3_26_), .Q(R2[26]) );
  TLATXL R2_reg_25_ ( .G(n192), .D(data_in_3_25_), .Q(R2[25]) );
  TLATXL R2_reg_24_ ( .G(n193), .D(data_in_3_24_), .Q(R2[24]) );
  TLATXL R3_reg_9_ ( .G(n188), .D(data_in_3_9_), .Q(R3[9]) );
  TLATXL R3_reg_8_ ( .G(n189), .D(data_in_3_8_), .Q(R3[8]) );
  TLATXL R3_reg_7_ ( .G(n188), .D(data_in_3_7_), .Q(R3[7]) );
  TLATXL R3_reg_6_ ( .G(n189), .D(data_in_3_6_), .Q(R3[6]) );
  TLATXL R3_reg_5_ ( .G(n188), .D(data_in_3_5_), .Q(R3[5]) );
  TLATXL R3_reg_4_ ( .G(n189), .D(data_in_3_4_), .Q(R3[4]) );
  TLATXL R4_reg_9_ ( .G(n190), .D(data_in_3_9_), .Q(R4[9]) );
  TLATXL R4_reg_8_ ( .G(n191), .D(data_in_3_8_), .Q(R4[8]) );
  TLATXL R4_reg_7_ ( .G(n190), .D(data_in_3_7_), .Q(R4[7]) );
  TLATXL R4_reg_6_ ( .G(n191), .D(data_in_3_6_), .Q(R4[6]) );
  TLATXL R4_reg_5_ ( .G(n190), .D(data_in_3_5_), .Q(R4[5]) );
  TLATXL R4_reg_4_ ( .G(n191), .D(data_in_3_4_), .Q(R4[4]) );
  TLATXL R1_reg_22_ ( .G(n186), .D(data_in_3_22_), .Q(R1[22]) );
  TLATXL R2_reg_23_ ( .G(n193), .D(data_in_3_23_), .Q(R2[23]) );
  TLATXL R2_reg_22_ ( .G(n193), .D(data_in_3_22_), .Q(R2[22]) );
  TLATXL R2_reg_21_ ( .G(n193), .D(data_in_3_21_), .Q(R2[21]) );
  TLATXL R2_reg_15_ ( .G(n193), .D(data_in_3_15_), .Q(R2[15]) );
  TLATXL R2_reg_12_ ( .G(n193), .D(data_in_3_12_), .Q(R2[12]) );
  TLATXL R3_reg_21_ ( .G(n189), .D(data_in_3_21_), .Q(R3[21]) );
  TLATXL R3_reg_15_ ( .G(n189), .D(data_in_3_15_), .Q(R3[15]) );
  TLATXL R3_reg_12_ ( .G(n189), .D(data_in_3_12_), .Q(R3[12]) );
  TLATXL R3_reg_11_ ( .G(n189), .D(data_in_3_11_), .Q(R3[11]) );
  TLATXL R3_reg_10_ ( .G(n189), .D(data_in_3_10_), .Q(R3[10]) );
  TLATXL R4_reg_21_ ( .G(n191), .D(data_in_3_21_), .Q(R4[21]) );
  TLATXL R4_reg_15_ ( .G(n191), .D(data_in_3_15_), .Q(R4[15]) );
  TLATXL R4_reg_12_ ( .G(n191), .D(data_in_3_12_), .Q(R4[12]) );
  TLATXL R4_reg_11_ ( .G(n191), .D(data_in_3_11_), .Q(R4[11]) );
  TLATXL R4_reg_10_ ( .G(n191), .D(data_in_3_10_), .Q(R4[10]) );
  TLATXL R1_reg_7_ ( .G(n185), .D(data_in_3_7_), .Q(R1[7]) );
  TLATXL R2_reg_11_ ( .G(n192), .D(data_in_3_11_), .Q(R2[11]) );
  TLATXL R2_reg_10_ ( .G(n192), .D(data_in_3_10_), .Q(R2[10]) );
  TLATXL R2_reg_9_ ( .G(n192), .D(data_in_3_9_), .Q(R2[9]) );
  TLATXL R2_reg_8_ ( .G(n192), .D(data_in_3_8_), .Q(R2[8]) );
  TLATXL R2_reg_7_ ( .G(n192), .D(data_in_3_7_), .Q(R2[7]) );
  TLATXL R2_reg_6_ ( .G(n192), .D(data_in_3_6_), .Q(R2[6]) );
  TLATXL R2_reg_5_ ( .G(n192), .D(data_in_3_5_), .Q(R2[5]) );
  TLATXL R2_reg_4_ ( .G(n192), .D(data_in_3_4_), .Q(R2[4]) );
  TLATXL R3_reg_33_ ( .G(n188), .D(data_in_3_33_), .Q(n52) );
  TLATXL R3_reg_32_ ( .G(n188), .D(data_in_3_32_), .Q(R3[32]) );
  TLATXL R3_reg_31_ ( .G(n188), .D(data_in_3_31_), .Q(R3[31]) );
  TLATXL R3_reg_30_ ( .G(n188), .D(data_in_3_30_), .Q(R3[30]) );
  TLATXL R3_reg_29_ ( .G(n188), .D(data_in_3_29_), .Q(R3[29]) );
  TLATXL R3_reg_28_ ( .G(n188), .D(data_in_3_28_), .Q(R3[28]) );
  TLATXL R3_reg_27_ ( .G(n188), .D(data_in_3_27_), .Q(R3[27]) );
  TLATXL R3_reg_26_ ( .G(n188), .D(data_in_3_26_), .Q(R3[26]) );
  TLATXL R3_reg_25_ ( .G(n188), .D(data_in_3_25_), .Q(R3[25]) );
  TLATXL R3_reg_24_ ( .G(n188), .D(data_in_3_24_), .Q(R3[24]) );
  TLATXL R3_reg_23_ ( .G(n188), .D(data_in_3_23_), .Q(R3[23]) );
  TLATXL R3_reg_22_ ( .G(n188), .D(data_in_3_22_), .Q(R3[22]) );
  TLATXL R4_reg_32_ ( .G(n190), .D(data_in_3_32_), .Q(R4[32]) );
  TLATXL R4_reg_31_ ( .G(n190), .D(data_in_3_31_), .Q(R4[31]) );
  TLATXL R4_reg_30_ ( .G(n190), .D(data_in_3_30_), .Q(R4[30]) );
  TLATXL R4_reg_29_ ( .G(n190), .D(data_in_3_29_), .Q(R4[29]) );
  TLATXL R4_reg_28_ ( .G(n190), .D(data_in_3_28_), .Q(R4[28]) );
  TLATXL R4_reg_27_ ( .G(n190), .D(data_in_3_27_), .Q(R4[27]) );
  TLATXL R4_reg_26_ ( .G(n190), .D(data_in_3_26_), .Q(R4[26]) );
  TLATXL R4_reg_25_ ( .G(n190), .D(data_in_3_25_), .Q(R4[25]) );
  TLATXL R4_reg_24_ ( .G(n190), .D(data_in_3_24_), .Q(R4[24]) );
  TLATXL R4_reg_23_ ( .G(n190), .D(data_in_3_23_), .Q(R4[23]) );
  TLATXL R4_reg_22_ ( .G(n190), .D(data_in_3_22_), .Q(R4[22]) );
  TLATXL R1_reg_33_ ( .G(n185), .D(data_in_3_33_), .Q(R1[33]) );
  TLATXL R1_reg_32_ ( .G(n186), .D(data_in_3_32_), .Q(R1[32]) );
  TLATXL R1_reg_31_ ( .G(n185), .D(data_in_3_31_), .Q(R1[31]) );
  TLATXL R1_reg_30_ ( .G(n186), .D(data_in_3_30_), .Q(R1[30]) );
  TLATXL R1_reg_29_ ( .G(n285), .D(data_in_3_29_), .Q(R1[29]) );
  TLATXL R1_reg_28_ ( .G(n285), .D(data_in_3_28_), .Q(R1[28]) );
  TLATXL R1_reg_27_ ( .G(n285), .D(data_in_3_27_), .Q(R1[27]) );
  TLATXL R1_reg_26_ ( .G(n285), .D(data_in_3_26_), .Q(R1[26]) );
  TLATXL R1_reg_25_ ( .G(n285), .D(data_in_3_25_), .Q(R1[25]) );
  TLATXL R1_reg_23_ ( .G(n186), .D(data_in_3_23_), .Q(R1[23]) );
  TLATXL R1_reg_21_ ( .G(n186), .D(data_in_3_21_), .Q(R1[21]) );
  TLATXL R1_reg_15_ ( .G(n186), .D(data_in_3_15_), .Q(R1[15]) );
  TLATXL R1_reg_12_ ( .G(n186), .D(data_in_3_12_), .Q(R1[12]) );
  TLATXL R1_reg_11_ ( .G(n185), .D(data_in_3_11_), .Q(R1[11]) );
  TLATXL R1_reg_10_ ( .G(n185), .D(data_in_3_10_), .Q(R1[10]) );
  TLATXL R1_reg_9_ ( .G(n185), .D(data_in_3_9_), .Q(R1[9]) );
  TLATXL R1_reg_8_ ( .G(n185), .D(data_in_3_8_), .Q(R1[8]) );
  TLATXL R1_reg_6_ ( .G(n185), .D(data_in_3_6_), .Q(R1[6]) );
  TLATXL R1_reg_5_ ( .G(n185), .D(data_in_3_5_), .Q(R1[5]) );
  TLATXL R1_reg_4_ ( .G(n185), .D(data_in_3_4_), .Q(R1[4]) );
  TLATXL R2_reg_1_ ( .G(n192), .D(data_in_3_1_), .Q(R2[1]) );
  TLATXL R2_reg_2_ ( .G(n192), .D(data_in_3_2_), .Q(R2[2]) );
  TLATXL R2_reg_3_ ( .G(n192), .D(data_in_3_3_), .Q(R2[3]) );
  TLATXL R4_reg_20_ ( .G(n191), .D(data_in_3_20_), .Q(R4[20]) );
  TLATXL R1_reg_20_ ( .G(n186), .D(data_in_3_20_), .Q(R1[20]) );
  TLATXL R1_reg_2_ ( .G(n185), .D(data_in_3_2_), .Q(R1[2]) );
  TLATXL R4_reg_1_ ( .G(n190), .D(data_in_3_1_), .Q(R4[1]) );
  TLATXL R2_reg_18_ ( .G(n193), .D(data_in_3_18_), .Q(R2[18]) );
  TLATXL R4_reg_18_ ( .G(n191), .D(data_in_3_18_), .Q(R4[18]) );
  TLATXL R4_reg_2_ ( .G(n191), .D(data_in_3_2_), .Q(R4[2]) );
  TLATXL R2_reg_19_ ( .G(n193), .D(data_in_3_19_), .Q(R2[19]) );
  TLATXL R4_reg_19_ ( .G(n191), .D(data_in_3_19_), .Q(R4[19]) );
  TLATXL R3_reg_1_ ( .G(n188), .D(data_in_3_1_), .Q(R3[1]) );
  TLATXL R3_reg_18_ ( .G(n189), .D(data_in_3_18_), .Q(R3[18]) );
  TLATXL R3_reg_2_ ( .G(n189), .D(data_in_3_2_), .Q(R3[2]) );
  TLATXL R3_reg_19_ ( .G(n189), .D(data_in_3_19_), .Q(R3[19]) );
  TLATXL R2_reg_20_ ( .G(n193), .D(data_in_3_20_), .Q(R2[20]) );
  TLATXL R3_reg_20_ ( .G(n189), .D(data_in_3_20_), .Q(R3[20]) );
  TLATXL R3_reg_3_ ( .G(n188), .D(data_in_3_3_), .Q(R3[3]) );
  TLATXL R4_reg_3_ ( .G(n190), .D(data_in_3_3_), .Q(R4[3]) );
  TLATXL R1_reg_3_ ( .G(n185), .D(data_in_3_3_), .Q(R1[3]) );
  TLATXL R1_reg_18_ ( .G(n186), .D(data_in_3_18_), .Q(R1[18]) );
  TLATXL R1_reg_0_ ( .G(n185), .D(data_in_3_0_), .Q(R1[0]) );
  TLATXL R1_reg_1_ ( .G(n185), .D(data_in_3_1_), .Q(R1[1]) );
  TLATXL R2_reg_17_ ( .G(n193), .D(data_in_3_17_), .Q(R2[17]) );
  TLATXL R2_reg_0_ ( .G(n192), .D(data_in_3_0_), .Q(R2[0]) );
  TLATXL R3_reg_17_ ( .G(n189), .D(data_in_3_17_), .Q(R3[17]) );
  TLATXL R3_reg_0_ ( .G(n189), .D(data_in_3_0_), .Q(R3[0]) );
  TLATXL R4_reg_17_ ( .G(n191), .D(data_in_3_17_), .Q(R4[17]) );
  TLATXL R4_reg_0_ ( .G(n191), .D(data_in_3_0_), .Q(R4[0]) );
  TLATXL R1_reg_19_ ( .G(n186), .D(data_in_3_19_), .Q(R1[19]) );
  TLATXL R1_reg_17_ ( .G(n186), .D(data_in_3_17_), .Q(R1[17]) );
  AND2X4 U4 ( .A(n16), .B(n11), .Y(n55) );
  NAND2X4 U5 ( .A(data_in_1[84]), .B(n160), .Y(n399) );
  BUFX3 U6 ( .A(n195), .Y(n1) );
  OAI21X2 U7 ( .A0(n160), .A1(n450), .B0(n449), .Y(n452) );
  NAND2X2 U8 ( .A(data_in_1[101]), .B(n160), .Y(n449) );
  OAI2BB1X2 U9 ( .A0N(data_in_2[6]), .A1N(n238), .B0(n203), .Y(data_out[6]) );
  OAI2BB1X2 U10 ( .A0N(data_in_2[9]), .A1N(n238), .B0(n209), .Y(data_out[9])
         );
  OAI2BB1X2 U11 ( .A0N(data_in_2[27]), .A1N(n167), .B0(n240), .Y(data_out[27])
         );
  OAI2BB1X2 U12 ( .A0N(data_in_2[29]), .A1N(n226), .B0(n244), .Y(data_out[29])
         );
  INVX1 U13 ( .A(data_in_1[50]), .Y(n13) );
  INVX1 U14 ( .A(data_in_2[101]), .Y(n450) );
  NAND2X1 U15 ( .A(n451), .B(R4[33]), .Y(n551) );
  INVX1 U16 ( .A(n160), .Y(n8) );
  CLKINVX3 U17 ( .A(n545), .Y(n177) );
  INVX4 U18 ( .A(n183), .Y(n178) );
  INVX4 U19 ( .A(n183), .Y(n182) );
  CLKINVX3 U20 ( .A(n177), .Y(n170) );
  OR3XL U21 ( .A(n14), .B(n2), .C(n10), .Y(n141) );
  BUFX8 U22 ( .A(counter[2]), .Y(n2) );
  NOR3BX4 U23 ( .AN(counter[1]), .B(n2), .C(n10), .Y(n298) );
  INVX8 U24 ( .A(n184), .Y(n181) );
  INVX2 U25 ( .A(n53), .Y(n241) );
  CLKINVX3 U26 ( .A(n233), .Y(n545) );
  INVX4 U27 ( .A(n184), .Y(n180) );
  OR2XL U28 ( .A(n140), .B(n141), .Y(n4) );
  INVX1 U29 ( .A(n176), .Y(n171) );
  OR3XL U30 ( .A(n282), .B(n557), .C(n558), .Y(n5) );
  OR2XL U31 ( .A(n3), .B(n141), .Y(n6) );
  INVXL U32 ( .A(n238), .Y(n168) );
  INVX1 U33 ( .A(n546), .Y(n183) );
  BUFX12 U34 ( .A(mux_flag), .Y(n160) );
  INVX1 U35 ( .A(n160), .Y(n194) );
  OAI2BB1X2 U36 ( .A0N(data_in_2[5]), .A1N(n202), .B0(n201), .Y(data_out[5])
         );
  OAI2BB1X2 U37 ( .A0N(data_in_2[30]), .A1N(n167), .B0(n245), .Y(data_out[30])
         );
  NAND3X2 U38 ( .A(n8), .B(data_in_2[118]), .C(n18), .Y(n500) );
  INVX2 U39 ( .A(n18), .Y(n17) );
  AOI22X1 U40 ( .A0(data_in_1[30]), .A1(n170), .B0(R1[30]), .B1(n181), .Y(n245) );
  NAND2X4 U41 ( .A(n140), .B(n298), .Y(n553) );
  NAND2X4 U42 ( .A(n9), .B(n352), .Y(data_out[67]) );
  AND2X4 U43 ( .A(n350), .B(n351), .Y(n9) );
  INVX8 U44 ( .A(n451), .Y(n18) );
  BUFX12 U45 ( .A(counter[3]), .Y(n10) );
  NAND2X4 U46 ( .A(n140), .B(n349), .Y(n550) );
  OAI2BB1X4 U47 ( .A0N(R2[16]), .A1N(n299), .B0(n300), .Y(n301) );
  NAND3X1 U48 ( .A(n194), .B(data_in_2[135]), .C(n553), .Y(n552) );
  AND3X2 U49 ( .A(n553), .B(n160), .C(data_in_1[135]), .Y(n56) );
  AND2X2 U50 ( .A(n1), .B(n194), .Y(n53) );
  AND2X1 U51 ( .A(data_in_1[118]), .B(n160), .Y(n11) );
  NAND2BX2 U52 ( .AN(n54), .B(n299), .Y(n401) );
  NAND2X1 U53 ( .A(n52), .B(n451), .Y(n12) );
  NAND3BX4 U54 ( .AN(n13), .B(n16), .C(n160), .Y(n300) );
  OAI2BB1X2 U55 ( .A0N(data_in_2[8]), .A1N(n226), .B0(n208), .Y(data_out[8])
         );
  INVX12 U56 ( .A(n1), .Y(n546) );
  OR2X4 U57 ( .A(n18), .B(n7), .Y(n499) );
  NOR3BX2 U58 ( .AN(data_in_2[50]), .B(n299), .C(n160), .Y(n302) );
  NAND2X4 U59 ( .A(n500), .B(n499), .Y(n501) );
  NAND2X2 U60 ( .A(n160), .B(n1), .Y(n233) );
  XOR2XL U61 ( .A(n14), .B(n3), .Y(N6) );
  NAND2BX4 U62 ( .AN(n51), .B(n17), .Y(n352) );
  INVX8 U63 ( .A(n553), .Y(n299) );
  NAND2BXL U64 ( .AN(n3), .B(n298), .Y(n195) );
  DLY1X1 U65 ( .A(counter[1]), .Y(n14) );
  AOI22X2 U66 ( .A0(data_in_1[31]), .A1(n170), .B0(R1[31]), .B1(n15), .Y(n246)
         );
  OAI2BB1X4 U67 ( .A0N(n452), .A1N(n18), .B0(n12), .Y(data_out[101]) );
  NAND3X1 U68 ( .A(data_in_1[67]), .B(n160), .C(n550), .Y(n351) );
  INVX8 U69 ( .A(n177), .Y(n169) );
  NAND3BX1 U70 ( .AN(n160), .B(data_in_2[67]), .C(n550), .Y(n350) );
  OAI2BB1X4 U71 ( .A0N(n402), .A1N(n16), .B0(n401), .Y(data_out[84]) );
  AOI22X1 U72 ( .A0(data_in_1[27]), .A1(n169), .B0(R1[27]), .B1(n181), .Y(n240) );
  CLKINVX8 U73 ( .A(n550), .Y(n451) );
  INVX12 U74 ( .A(n183), .Y(n15) );
  INVX12 U75 ( .A(n184), .Y(n179) );
  CLKINVX4 U76 ( .A(n546), .Y(n184) );
  INVX8 U77 ( .A(n299), .Y(n16) );
  INVX4 U78 ( .A(n241), .Y(n167) );
  AOI22X1 U79 ( .A0(data_in_1[0]), .A1(n545), .B0(R1[0]), .B1(n180), .Y(n196)
         );
  INVX4 U80 ( .A(data_in_2[84]), .Y(n400) );
  OAI21XL U81 ( .A0(n160), .A1(n400), .B0(n399), .Y(n402) );
  AOI22X2 U82 ( .A0(data_in_1[18]), .A1(n169), .B0(R1[18]), .B1(n180), .Y(n219) );
  AOI22X2 U83 ( .A0(data_in_1[17]), .A1(n169), .B0(R1[17]), .B1(n181), .Y(n218) );
  AOI22XL U84 ( .A0(data_in_1[2]), .A1(n169), .B0(R1[2]), .B1(n180), .Y(n198)
         );
  AOI22XL U85 ( .A0(data_in_1[29]), .A1(n169), .B0(R1[29]), .B1(n181), .Y(n244) );
  AOI22XL U86 ( .A0(data_in_1[32]), .A1(n170), .B0(R1[32]), .B1(n178), .Y(n247) );
  OAI2BB1X1 U87 ( .A0N(data_in_2[12]), .A1N(n167), .B0(n213), .Y(data_out[12])
         );
  AOI22XL U88 ( .A0(data_in_1[33]), .A1(n170), .B0(R1[33]), .B1(n181), .Y(n248) );
  AOI22XL U89 ( .A0(data_in_1[68]), .A1(n170), .B0(R3[0]), .B1(n179), .Y(n353)
         );
  AOI22XL U90 ( .A0(data_in_1[51]), .A1(n170), .B0(R2[17]), .B1(n15), .Y(n303)
         );
  AOI22XL U91 ( .A0(data_in_1[34]), .A1(n170), .B0(R2[0]), .B1(n182), .Y(n249)
         );
  AOI22XL U92 ( .A0(data_in_1[85]), .A1(n170), .B0(R3[17]), .B1(n181), .Y(n403) );
  AOI22XL U93 ( .A0(data_in_1[119]), .A1(n170), .B0(R4[17]), .B1(n181), .Y(
        n502) );
  AOI22XL U94 ( .A0(data_in_1[102]), .A1(n170), .B0(R4[0]), .B1(n181), .Y(n453) );
  NAND2XL U95 ( .A(R4[21]), .B(n181), .Y(n512) );
  NAND2XL U96 ( .A(R4[22]), .B(n181), .Y(n515) );
  NAND2XL U97 ( .A(R4[23]), .B(n546), .Y(n518) );
  NAND2XL U98 ( .A(R4[24]), .B(n15), .Y(n521) );
  NAND2XL U99 ( .A(R4[25]), .B(n15), .Y(n524) );
  NAND2XL U100 ( .A(R4[26]), .B(n180), .Y(n527) );
  NAND2XL U101 ( .A(R4[27]), .B(n178), .Y(n530) );
  NAND2XL U102 ( .A(R4[28]), .B(n181), .Y(n533) );
  NAND2XL U103 ( .A(R4[29]), .B(n179), .Y(n536) );
  NAND2XL U104 ( .A(data_in_1[132]), .B(n170), .Y(n540) );
  NAND2XL U105 ( .A(R4[30]), .B(n15), .Y(n539) );
  NAND2XL U106 ( .A(data_in_1[133]), .B(n170), .Y(n543) );
  NAND2XL U107 ( .A(R4[31]), .B(n182), .Y(n542) );
  NAND2XL U108 ( .A(R4[20]), .B(n181), .Y(n509) );
  NAND2XL U109 ( .A(R4[14]), .B(n181), .Y(n493) );
  NAND2XL U110 ( .A(data_in_1[35]), .B(n170), .Y(n251) );
  INVX1 U111 ( .A(n176), .Y(n174) );
  INVX1 U112 ( .A(n176), .Y(n172) );
  INVX1 U113 ( .A(n176), .Y(n173) );
  INVX1 U114 ( .A(n176), .Y(n175) );
  INVX1 U115 ( .A(n168), .Y(n165) );
  INVX1 U116 ( .A(n168), .Y(n164) );
  INVX1 U117 ( .A(n168), .Y(n163) );
  INVX1 U118 ( .A(n168), .Y(n162) );
  INVX1 U119 ( .A(n168), .Y(n166) );
  INVX1 U120 ( .A(n168), .Y(n161) );
  INVX1 U121 ( .A(n5), .Y(n193) );
  INVXL U122 ( .A(n545), .Y(n176) );
  INVX1 U123 ( .A(n5), .Y(n192) );
  INVX1 U124 ( .A(n4), .Y(n191) );
  INVX1 U125 ( .A(n6), .Y(n189) );
  INVX1 U126 ( .A(n187), .Y(n186) );
  XOR2X1 U127 ( .A(n557), .B(n282), .Y(N7) );
  INVX1 U128 ( .A(n4), .Y(n190) );
  INVX1 U129 ( .A(n6), .Y(n188) );
  INVX1 U130 ( .A(n187), .Y(n185) );
  INVX1 U131 ( .A(n285), .Y(n187) );
  OR2X4 U132 ( .A(n501), .B(n55), .Y(data_out[118]) );
  OR2X4 U133 ( .A(n554), .B(n56), .Y(data_out[135]) );
  NAND2BX2 U134 ( .AN(n236), .B(n235), .Y(data_out[24]) );
  OAI22XL U135 ( .A0(n241), .A1(n234), .B0(n233), .B1(n232), .Y(n236) );
  NAND2X1 U136 ( .A(R1[24]), .B(n180), .Y(n235) );
  INVX1 U137 ( .A(data_in_2[24]), .Y(n234) );
  NAND2BX2 U138 ( .AN(n207), .B(n206), .Y(data_out[7]) );
  OAI22XL U139 ( .A0(n241), .A1(n205), .B0(n233), .B1(n204), .Y(n207) );
  NAND2X1 U140 ( .A(R1[7]), .B(n179), .Y(n206) );
  INVX1 U141 ( .A(data_in_2[7]), .Y(n205) );
  OAI22XL U142 ( .A0(n241), .A1(n228), .B0(n233), .B1(n227), .Y(n230) );
  NAND2X1 U143 ( .A(R1[22]), .B(n15), .Y(n229) );
  INVX1 U144 ( .A(data_in_2[22]), .Y(n228) );
  OAI22XL U145 ( .A0(n241), .A1(n221), .B0(n233), .B1(n220), .Y(n223) );
  NAND2X2 U146 ( .A(R1[19]), .B(n15), .Y(n222) );
  INVX1 U147 ( .A(data_in_2[19]), .Y(n221) );
  INVXL U148 ( .A(n241), .Y(n202) );
  AOI22XL U149 ( .A0(data_in_1[5]), .A1(n545), .B0(R1[5]), .B1(n179), .Y(n201)
         );
  AOI22X2 U150 ( .A0(data_in_1[3]), .A1(n169), .B0(R1[3]), .B1(n181), .Y(n199)
         );
  OAI2BB1X2 U151 ( .A0N(data_in_2[28]), .A1N(n243), .B0(n242), .Y(data_out[28]) );
  INVXL U152 ( .A(n241), .Y(n243) );
  AOI22XL U153 ( .A0(data_in_1[28]), .A1(n169), .B0(R1[28]), .B1(n179), .Y(
        n242) );
  INVXL U154 ( .A(n241), .Y(n238) );
  AOI22XL U155 ( .A0(data_in_1[25]), .A1(n169), .B0(R1[25]), .B1(n181), .Y(
        n237) );
  INVXL U156 ( .A(n241), .Y(n226) );
  AOI22XL U157 ( .A0(data_in_1[21]), .A1(n169), .B0(R1[21]), .B1(n15), .Y(n225) );
  OAI2BB1X2 U158 ( .A0N(data_in_2[11]), .A1N(n212), .B0(n211), .Y(data_out[11]) );
  INVXL U159 ( .A(n241), .Y(n212) );
  AOI22XL U160 ( .A0(data_in_1[11]), .A1(n169), .B0(R1[11]), .B1(n181), .Y(
        n211) );
  AOI22XL U161 ( .A0(data_in_1[26]), .A1(n169), .B0(R1[26]), .B1(n181), .Y(
        n239) );
  OAI2BB1X2 U162 ( .A0N(data_in_2[10]), .A1N(n212), .B0(n210), .Y(data_out[10]) );
  AOI22XL U163 ( .A0(data_in_1[10]), .A1(n169), .B0(R1[10]), .B1(n178), .Y(
        n210) );
  AOI22XL U164 ( .A0(data_in_1[9]), .A1(n169), .B0(R1[9]), .B1(n546), .Y(n209)
         );
  AOI22XL U165 ( .A0(data_in_1[4]), .A1(n169), .B0(R1[4]), .B1(n15), .Y(n200)
         );
  AOI22XL U166 ( .A0(data_in_1[6]), .A1(n169), .B0(R1[6]), .B1(n182), .Y(n203)
         );
  OAI2BB1X1 U167 ( .A0N(data_in_2[13]), .A1N(n167), .B0(n214), .Y(data_out[13]) );
  OAI2BB1X1 U168 ( .A0N(data_in_2[14]), .A1N(n167), .B0(n215), .Y(data_out[14]) );
  AOI22XL U169 ( .A0(data_in_1[14]), .A1(n169), .B0(R1[14]), .B1(n15), .Y(n215) );
  AOI22XL U170 ( .A0(data_in_1[20]), .A1(n169), .B0(R1[20]), .B1(n178), .Y(
        n224) );
  OAI2BB1X1 U171 ( .A0N(data_in_2[31]), .A1N(n167), .B0(n246), .Y(data_out[31]) );
  AOI22XL U172 ( .A0(data_in_1[12]), .A1(n169), .B0(R1[12]), .B1(n546), .Y(
        n213) );
  AOI22XL U173 ( .A0(data_in_1[23]), .A1(n169), .B0(R1[23]), .B1(n546), .Y(
        n231) );
  AOI22XL U174 ( .A0(data_in_1[8]), .A1(n169), .B0(R1[8]), .B1(n181), .Y(n208)
         );
  OAI2BB1X1 U175 ( .A0N(data_in_2[15]), .A1N(n212), .B0(n216), .Y(data_out[15]) );
  AOI22XL U176 ( .A0(data_in_1[15]), .A1(n169), .B0(R1[15]), .B1(n181), .Y(
        n216) );
  OAI2BB1X1 U177 ( .A0N(data_in_2[32]), .A1N(n212), .B0(n247), .Y(data_out[32]) );
  INVX1 U178 ( .A(data_in_1[19]), .Y(n220) );
  OAI2BB1X1 U179 ( .A0N(data_in_2[16]), .A1N(n243), .B0(n217), .Y(data_out[16]) );
  OAI2BB1X1 U180 ( .A0N(data_in_2[33]), .A1N(n212), .B0(n248), .Y(data_out[33]) );
  INVX1 U181 ( .A(data_in_1[24]), .Y(n232) );
  INVX1 U182 ( .A(data_in_1[7]), .Y(n204) );
  INVX1 U183 ( .A(data_in_1[22]), .Y(n227) );
  INVXL U184 ( .A(n2), .Y(n557) );
  XOR2X1 U185 ( .A(n10), .B(n281), .Y(N8) );
  NOR2X1 U186 ( .A(n557), .B(n282), .Y(n281) );
  OAI2BB1X1 U187 ( .A0N(data_in_2[102]), .A1N(n165), .B0(n453), .Y(
        data_out[102]) );
  NAND3X1 U188 ( .A(n291), .B(n290), .C(n289), .Y(data_out[47]) );
  NAND2X1 U189 ( .A(data_in_1[47]), .B(n175), .Y(n290) );
  NAND2X1 U190 ( .A(data_in_2[47]), .B(n166), .Y(n291) );
  NAND3X1 U191 ( .A(n392), .B(n391), .C(n390), .Y(data_out[81]) );
  NAND2X1 U192 ( .A(data_in_1[81]), .B(n173), .Y(n391) );
  NAND2X1 U193 ( .A(data_in_2[81]), .B(n164), .Y(n392) );
  NAND3X1 U194 ( .A(n492), .B(n491), .C(n490), .Y(data_out[115]) );
  NAND2X1 U195 ( .A(data_in_1[115]), .B(n171), .Y(n491) );
  NAND2X1 U196 ( .A(data_in_2[115]), .B(n162), .Y(n492) );
  NAND3X1 U197 ( .A(n456), .B(n455), .C(n454), .Y(data_out[103]) );
  NAND2X1 U198 ( .A(data_in_1[103]), .B(n172), .Y(n455) );
  NAND2X1 U199 ( .A(R4[1]), .B(n546), .Y(n454) );
  NAND2X1 U200 ( .A(data_in_2[103]), .B(n163), .Y(n456) );
  NAND3X1 U201 ( .A(n255), .B(n254), .C(n253), .Y(data_out[36]) );
  NAND2X1 U202 ( .A(data_in_1[36]), .B(n171), .Y(n254) );
  NAND2XL U203 ( .A(R2[2]), .B(n181), .Y(n253) );
  NAND2X1 U204 ( .A(data_in_2[36]), .B(n165), .Y(n255) );
  NAND3X1 U205 ( .A(n459), .B(n458), .C(n457), .Y(data_out[104]) );
  NAND2X1 U206 ( .A(data_in_1[104]), .B(n172), .Y(n458) );
  NAND2X1 U207 ( .A(R4[2]), .B(n15), .Y(n457) );
  NAND2X1 U208 ( .A(data_in_2[104]), .B(n163), .Y(n459) );
  NAND3X1 U209 ( .A(n312), .B(n311), .C(n310), .Y(data_out[54]) );
  NAND2X1 U210 ( .A(data_in_1[54]), .B(n175), .Y(n311) );
  NAND2X1 U211 ( .A(R2[20]), .B(n182), .Y(n310) );
  NAND2X1 U212 ( .A(data_in_2[54]), .B(n166), .Y(n312) );
  NAND3X1 U213 ( .A(n362), .B(n361), .C(n360), .Y(data_out[71]) );
  NAND2X1 U214 ( .A(data_in_1[71]), .B(n173), .Y(n361) );
  NAND2X1 U215 ( .A(data_in_2[71]), .B(n165), .Y(n362) );
  NAND2X1 U216 ( .A(R3[3]), .B(n179), .Y(n360) );
  NAND3X1 U217 ( .A(n462), .B(n461), .C(n460), .Y(data_out[105]) );
  NAND2X1 U218 ( .A(data_in_1[105]), .B(n172), .Y(n461) );
  NAND2X1 U219 ( .A(R4[3]), .B(n181), .Y(n460) );
  NAND2X1 U220 ( .A(data_in_2[105]), .B(n163), .Y(n462) );
  NAND3X1 U221 ( .A(n315), .B(n314), .C(n313), .Y(data_out[55]) );
  NAND2X1 U222 ( .A(data_in_1[55]), .B(n174), .Y(n314) );
  NAND2X1 U223 ( .A(R2[21]), .B(n181), .Y(n313) );
  NAND2X1 U224 ( .A(data_in_2[55]), .B(n166), .Y(n315) );
  NAND3X1 U225 ( .A(n261), .B(n260), .C(n259), .Y(data_out[38]) );
  NAND2X1 U226 ( .A(data_in_1[38]), .B(n175), .Y(n260) );
  NAND2XL U227 ( .A(R2[4]), .B(n546), .Y(n259) );
  NAND2X1 U228 ( .A(data_in_2[38]), .B(n164), .Y(n261) );
  NAND3X1 U229 ( .A(n365), .B(n364), .C(n363), .Y(data_out[72]) );
  NAND2X1 U230 ( .A(data_in_1[72]), .B(n173), .Y(n364) );
  NAND2X1 U231 ( .A(data_in_2[72]), .B(n165), .Y(n365) );
  NAND2X1 U232 ( .A(R3[4]), .B(n15), .Y(n363) );
  NAND3X1 U233 ( .A(n514), .B(n513), .C(n512), .Y(data_out[123]) );
  NAND2X1 U234 ( .A(data_in_1[123]), .B(n171), .Y(n513) );
  NAND2X1 U235 ( .A(data_in_2[123]), .B(n161), .Y(n514) );
  NAND3X1 U236 ( .A(n465), .B(n464), .C(n463), .Y(data_out[106]) );
  NAND2X1 U237 ( .A(data_in_1[106]), .B(n172), .Y(n464) );
  NAND2X1 U238 ( .A(data_in_2[106]), .B(n162), .Y(n465) );
  NAND2X1 U239 ( .A(R4[4]), .B(n15), .Y(n463) );
  NAND3X1 U240 ( .A(n318), .B(n317), .C(n316), .Y(data_out[56]) );
  NAND2X1 U241 ( .A(data_in_1[56]), .B(n174), .Y(n317) );
  NAND2X1 U242 ( .A(R2[22]), .B(n181), .Y(n316) );
  NAND2X1 U243 ( .A(data_in_2[56]), .B(n166), .Y(n318) );
  NAND3X1 U244 ( .A(n264), .B(n263), .C(n262), .Y(data_out[39]) );
  NAND2XL U245 ( .A(R2[5]), .B(n15), .Y(n262) );
  NAND2X1 U246 ( .A(data_in_1[39]), .B(n175), .Y(n263) );
  NAND2X1 U247 ( .A(data_in_2[39]), .B(n163), .Y(n264) );
  NAND3X1 U248 ( .A(n368), .B(n367), .C(n366), .Y(data_out[73]) );
  NAND2X1 U249 ( .A(data_in_1[73]), .B(n173), .Y(n367) );
  NAND2X1 U250 ( .A(data_in_2[73]), .B(n165), .Y(n368) );
  NAND2X1 U251 ( .A(R3[5]), .B(n182), .Y(n366) );
  NAND3X1 U252 ( .A(n517), .B(n516), .C(n515), .Y(data_out[124]) );
  NAND2X1 U253 ( .A(data_in_1[124]), .B(n171), .Y(n516) );
  NAND2X1 U254 ( .A(data_in_2[124]), .B(n161), .Y(n517) );
  NAND3X1 U255 ( .A(n468), .B(n467), .C(n466), .Y(data_out[107]) );
  NAND2X1 U256 ( .A(data_in_1[107]), .B(n172), .Y(n467) );
  NAND2X1 U257 ( .A(R4[5]), .B(n180), .Y(n466) );
  NAND2X1 U258 ( .A(data_in_2[107]), .B(n162), .Y(n468) );
  NAND3X1 U259 ( .A(n321), .B(n320), .C(n319), .Y(data_out[57]) );
  NAND2X1 U260 ( .A(data_in_1[57]), .B(n174), .Y(n320) );
  NAND2X1 U261 ( .A(R2[23]), .B(n181), .Y(n319) );
  NAND2X1 U262 ( .A(data_in_2[57]), .B(n165), .Y(n321) );
  NAND3X1 U263 ( .A(n267), .B(n266), .C(n265), .Y(data_out[40]) );
  NAND2XL U264 ( .A(R2[6]), .B(n15), .Y(n265) );
  NAND2X1 U265 ( .A(data_in_1[40]), .B(n175), .Y(n266) );
  NAND2X1 U266 ( .A(data_in_2[40]), .B(n162), .Y(n267) );
  NAND3X1 U267 ( .A(n371), .B(n370), .C(n369), .Y(data_out[74]) );
  NAND2X1 U268 ( .A(data_in_1[74]), .B(n173), .Y(n370) );
  NAND2X1 U269 ( .A(R3[6]), .B(n178), .Y(n369) );
  NAND2X1 U270 ( .A(data_in_2[74]), .B(n165), .Y(n371) );
  NAND3X1 U271 ( .A(n520), .B(n519), .C(n518), .Y(data_out[125]) );
  NAND2X1 U272 ( .A(data_in_1[125]), .B(n171), .Y(n519) );
  NAND2X1 U273 ( .A(data_in_2[125]), .B(n161), .Y(n520) );
  NAND3X1 U274 ( .A(n471), .B(n470), .C(n469), .Y(data_out[108]) );
  NAND2X1 U275 ( .A(data_in_1[108]), .B(n172), .Y(n470) );
  NAND2X1 U276 ( .A(R4[6]), .B(n178), .Y(n469) );
  NAND2X1 U277 ( .A(data_in_2[108]), .B(n162), .Y(n471) );
  NAND3X1 U278 ( .A(n324), .B(n323), .C(n322), .Y(data_out[58]) );
  NAND2X1 U279 ( .A(data_in_1[58]), .B(n174), .Y(n323) );
  NAND2X1 U280 ( .A(data_in_2[58]), .B(n166), .Y(n324) );
  NAND2X1 U281 ( .A(R2[24]), .B(n181), .Y(n322) );
  NAND3X1 U282 ( .A(n270), .B(n269), .C(n268), .Y(data_out[41]) );
  NAND2XL U283 ( .A(R2[7]), .B(n180), .Y(n268) );
  NAND2X1 U284 ( .A(data_in_1[41]), .B(n175), .Y(n269) );
  NAND2X1 U285 ( .A(data_in_2[41]), .B(n161), .Y(n270) );
  NAND3X1 U286 ( .A(n374), .B(n373), .C(n372), .Y(data_out[75]) );
  NAND2X1 U287 ( .A(data_in_1[75]), .B(n173), .Y(n373) );
  NAND2X1 U288 ( .A(R3[7]), .B(n181), .Y(n372) );
  NAND2X1 U289 ( .A(data_in_2[75]), .B(n165), .Y(n374) );
  NAND3X1 U290 ( .A(n523), .B(n522), .C(n521), .Y(data_out[126]) );
  NAND2X1 U291 ( .A(data_in_1[126]), .B(n171), .Y(n522) );
  NAND2X1 U292 ( .A(data_in_2[126]), .B(n161), .Y(n523) );
  NAND3X1 U293 ( .A(n474), .B(n473), .C(n472), .Y(data_out[109]) );
  NAND2X1 U294 ( .A(data_in_1[109]), .B(n172), .Y(n473) );
  NAND2X1 U295 ( .A(R4[7]), .B(n181), .Y(n472) );
  NAND2X1 U296 ( .A(data_in_2[109]), .B(n162), .Y(n474) );
  NAND3X1 U297 ( .A(n327), .B(n326), .C(n325), .Y(data_out[59]) );
  NAND2X1 U298 ( .A(data_in_1[59]), .B(n174), .Y(n326) );
  NAND2X1 U299 ( .A(data_in_2[59]), .B(n166), .Y(n327) );
  NAND2X1 U300 ( .A(R2[25]), .B(n181), .Y(n325) );
  NAND3X1 U301 ( .A(n273), .B(n272), .C(n271), .Y(data_out[42]) );
  NAND2X1 U302 ( .A(data_in_1[42]), .B(n175), .Y(n272) );
  NAND2X1 U303 ( .A(data_in_2[42]), .B(n166), .Y(n273) );
  NAND2X1 U304 ( .A(R2[8]), .B(n546), .Y(n271) );
  NAND3X1 U305 ( .A(n427), .B(n426), .C(n425), .Y(data_out[93]) );
  NAND2X1 U306 ( .A(data_in_1[93]), .B(n172), .Y(n426) );
  NAND2X1 U307 ( .A(data_in_2[93]), .B(n163), .Y(n427) );
  NAND2X1 U308 ( .A(R3[25]), .B(n180), .Y(n425) );
  NAND3X1 U309 ( .A(n377), .B(n376), .C(n375), .Y(data_out[76]) );
  NAND2X1 U310 ( .A(data_in_1[76]), .B(n173), .Y(n376) );
  NAND2X1 U311 ( .A(R3[8]), .B(n179), .Y(n375) );
  NAND2X1 U312 ( .A(data_in_2[76]), .B(n164), .Y(n377) );
  NAND3X1 U313 ( .A(n526), .B(n525), .C(n524), .Y(data_out[127]) );
  NAND2X1 U314 ( .A(data_in_1[127]), .B(n171), .Y(n525) );
  NAND2X1 U315 ( .A(data_in_2[127]), .B(n161), .Y(n526) );
  NAND3X1 U316 ( .A(n477), .B(n476), .C(n475), .Y(data_out[110]) );
  NAND2X1 U317 ( .A(data_in_1[110]), .B(n172), .Y(n476) );
  NAND2X1 U318 ( .A(R4[8]), .B(n179), .Y(n475) );
  NAND2X1 U319 ( .A(data_in_2[110]), .B(n162), .Y(n477) );
  NAND3X1 U320 ( .A(n330), .B(n329), .C(n328), .Y(data_out[60]) );
  NAND2X1 U321 ( .A(data_in_1[60]), .B(n174), .Y(n329) );
  NAND2X1 U322 ( .A(data_in_2[60]), .B(n166), .Y(n330) );
  NAND2X1 U323 ( .A(R2[26]), .B(n181), .Y(n328) );
  NAND3X1 U324 ( .A(n276), .B(n275), .C(n274), .Y(data_out[43]) );
  NAND2X1 U325 ( .A(data_in_1[43]), .B(n175), .Y(n275) );
  NAND2X1 U326 ( .A(data_in_2[43]), .B(n165), .Y(n276) );
  NAND2X1 U327 ( .A(R2[9]), .B(n15), .Y(n274) );
  NAND3X1 U328 ( .A(n430), .B(n429), .C(n428), .Y(data_out[94]) );
  NAND2X1 U329 ( .A(data_in_1[94]), .B(n173), .Y(n429) );
  NAND2X1 U330 ( .A(data_in_2[94]), .B(n163), .Y(n430) );
  NAND2X1 U331 ( .A(R3[26]), .B(n178), .Y(n428) );
  NAND3X1 U332 ( .A(n380), .B(n379), .C(n378), .Y(data_out[77]) );
  NAND2X1 U333 ( .A(data_in_1[77]), .B(n173), .Y(n379) );
  NAND2X1 U334 ( .A(R3[9]), .B(n15), .Y(n378) );
  NAND2X1 U335 ( .A(data_in_2[77]), .B(n164), .Y(n380) );
  NAND3X1 U336 ( .A(n529), .B(n528), .C(n527), .Y(data_out[128]) );
  NAND2X1 U337 ( .A(data_in_1[128]), .B(n171), .Y(n528) );
  NAND2X1 U338 ( .A(data_in_2[128]), .B(n161), .Y(n529) );
  NAND3X1 U339 ( .A(n480), .B(n479), .C(n478), .Y(data_out[111]) );
  NAND2X1 U340 ( .A(data_in_1[111]), .B(n172), .Y(n479) );
  NAND2X1 U341 ( .A(R4[9]), .B(n15), .Y(n478) );
  NAND2X1 U342 ( .A(data_in_2[111]), .B(n162), .Y(n480) );
  NAND3X1 U343 ( .A(n333), .B(n332), .C(n331), .Y(data_out[61]) );
  NAND2X1 U344 ( .A(data_in_1[61]), .B(n174), .Y(n332) );
  NAND2X1 U345 ( .A(data_in_2[61]), .B(n166), .Y(n333) );
  NAND2X1 U346 ( .A(R2[27]), .B(n546), .Y(n331) );
  NAND3X1 U347 ( .A(n279), .B(n278), .C(n277), .Y(data_out[44]) );
  NAND2X1 U348 ( .A(data_in_1[44]), .B(n175), .Y(n278) );
  NAND2X1 U349 ( .A(data_in_2[44]), .B(n164), .Y(n279) );
  NAND2X1 U350 ( .A(R2[10]), .B(n15), .Y(n277) );
  NAND3X1 U351 ( .A(n433), .B(n432), .C(n431), .Y(data_out[95]) );
  NAND2X1 U352 ( .A(data_in_1[95]), .B(n171), .Y(n432) );
  NAND2X1 U353 ( .A(data_in_2[95]), .B(n163), .Y(n433) );
  NAND2X1 U354 ( .A(R3[27]), .B(n181), .Y(n431) );
  NAND3X1 U355 ( .A(n383), .B(n382), .C(n381), .Y(data_out[78]) );
  NAND2X1 U356 ( .A(data_in_1[78]), .B(n173), .Y(n382) );
  NAND2X1 U357 ( .A(R3[10]), .B(n182), .Y(n381) );
  NAND2X1 U358 ( .A(data_in_2[78]), .B(n164), .Y(n383) );
  NAND3X1 U359 ( .A(n532), .B(n531), .C(n530), .Y(data_out[129]) );
  NAND2X1 U360 ( .A(data_in_1[129]), .B(n171), .Y(n531) );
  NAND2X1 U361 ( .A(data_in_2[129]), .B(n161), .Y(n532) );
  NAND3X1 U362 ( .A(n483), .B(n482), .C(n481), .Y(data_out[112]) );
  NAND2X1 U363 ( .A(data_in_1[112]), .B(n172), .Y(n482) );
  NAND2X1 U364 ( .A(R4[10]), .B(n182), .Y(n481) );
  NAND2X1 U365 ( .A(data_in_2[112]), .B(n162), .Y(n483) );
  NAND3X1 U366 ( .A(n336), .B(n335), .C(n334), .Y(data_out[62]) );
  NAND2X1 U367 ( .A(data_in_1[62]), .B(n174), .Y(n335) );
  NAND2X1 U368 ( .A(data_in_2[62]), .B(n166), .Y(n336) );
  NAND2X1 U369 ( .A(R2[28]), .B(n15), .Y(n334) );
  NAND3X1 U370 ( .A(n284), .B(n283), .C(n280), .Y(data_out[45]) );
  NAND2X1 U371 ( .A(data_in_1[45]), .B(n175), .Y(n283) );
  NAND2X1 U372 ( .A(R2[11]), .B(n180), .Y(n280) );
  NAND2X1 U373 ( .A(data_in_2[45]), .B(n166), .Y(n284) );
  NAND3X1 U374 ( .A(n436), .B(n435), .C(n434), .Y(data_out[96]) );
  NAND2X1 U375 ( .A(data_in_1[96]), .B(n172), .Y(n435) );
  NAND2X1 U376 ( .A(data_in_2[96]), .B(n163), .Y(n436) );
  NAND2X1 U377 ( .A(R3[28]), .B(n179), .Y(n434) );
  NAND3X1 U378 ( .A(n386), .B(n385), .C(n384), .Y(data_out[79]) );
  NAND2X1 U379 ( .A(data_in_1[79]), .B(n173), .Y(n385) );
  NAND2X1 U380 ( .A(R3[11]), .B(n181), .Y(n384) );
  NAND2X1 U381 ( .A(data_in_2[79]), .B(n164), .Y(n386) );
  NAND3X1 U382 ( .A(n535), .B(n534), .C(n533), .Y(data_out[130]) );
  NAND2X1 U383 ( .A(data_in_1[130]), .B(n171), .Y(n534) );
  NAND2X1 U384 ( .A(data_in_2[130]), .B(n161), .Y(n535) );
  NAND3X1 U385 ( .A(n486), .B(n485), .C(n484), .Y(data_out[113]) );
  NAND2X1 U386 ( .A(data_in_1[113]), .B(n172), .Y(n485) );
  NAND2X1 U387 ( .A(R4[11]), .B(n181), .Y(n484) );
  NAND2X1 U388 ( .A(data_in_2[113]), .B(n162), .Y(n486) );
  NAND3X1 U389 ( .A(n339), .B(n338), .C(n337), .Y(data_out[63]) );
  NAND2X1 U390 ( .A(data_in_1[63]), .B(n174), .Y(n338) );
  NAND2X1 U391 ( .A(data_in_2[63]), .B(n165), .Y(n339) );
  NAND2X1 U392 ( .A(R2[29]), .B(n15), .Y(n337) );
  NAND3X1 U393 ( .A(n288), .B(n287), .C(n286), .Y(data_out[46]) );
  NAND2X1 U394 ( .A(data_in_1[46]), .B(n175), .Y(n287) );
  NAND2X1 U395 ( .A(data_in_2[46]), .B(n163), .Y(n288) );
  NAND2X1 U396 ( .A(R2[12]), .B(n178), .Y(n286) );
  NAND3X1 U397 ( .A(n439), .B(n438), .C(n437), .Y(data_out[97]) );
  NAND2X1 U398 ( .A(data_in_1[97]), .B(n175), .Y(n438) );
  NAND2X1 U399 ( .A(data_in_2[97]), .B(n163), .Y(n439) );
  NAND2X1 U400 ( .A(R3[29]), .B(n15), .Y(n437) );
  NAND3X1 U401 ( .A(n389), .B(n388), .C(n387), .Y(data_out[80]) );
  NAND2X1 U402 ( .A(data_in_1[80]), .B(n173), .Y(n388) );
  NAND2X1 U403 ( .A(R3[12]), .B(n181), .Y(n387) );
  NAND2X1 U404 ( .A(data_in_2[80]), .B(n164), .Y(n389) );
  NAND3X1 U405 ( .A(n538), .B(n537), .C(n536), .Y(data_out[131]) );
  NAND2X1 U406 ( .A(data_in_1[131]), .B(n171), .Y(n537) );
  NAND2X1 U407 ( .A(data_in_2[131]), .B(n161), .Y(n538) );
  NAND3X1 U408 ( .A(n489), .B(n488), .C(n487), .Y(data_out[114]) );
  NAND2X1 U409 ( .A(data_in_1[114]), .B(n172), .Y(n488) );
  NAND2X1 U410 ( .A(R4[12]), .B(n181), .Y(n487) );
  NAND2X1 U411 ( .A(data_in_2[114]), .B(n162), .Y(n489) );
  NAND3X1 U412 ( .A(n342), .B(n341), .C(n340), .Y(data_out[64]) );
  NAND2X1 U413 ( .A(data_in_1[64]), .B(n174), .Y(n341) );
  NAND2X1 U414 ( .A(data_in_2[64]), .B(n165), .Y(n342) );
  NAND2X1 U415 ( .A(R2[30]), .B(n180), .Y(n340) );
  NAND3X1 U416 ( .A(n442), .B(n441), .C(n440), .Y(data_out[98]) );
  NAND2X1 U417 ( .A(data_in_1[98]), .B(n174), .Y(n441) );
  NAND2X1 U418 ( .A(data_in_2[98]), .B(n163), .Y(n442) );
  NAND2X1 U419 ( .A(R3[30]), .B(n182), .Y(n440) );
  NAND3X1 U420 ( .A(n541), .B(n540), .C(n539), .Y(data_out[132]) );
  NAND2X1 U421 ( .A(data_in_2[132]), .B(n161), .Y(n541) );
  NAND3X1 U422 ( .A(n345), .B(n344), .C(n343), .Y(data_out[65]) );
  NAND2X1 U423 ( .A(data_in_1[65]), .B(n174), .Y(n344) );
  NAND2X1 U424 ( .A(data_in_2[65]), .B(n165), .Y(n345) );
  NAND2X1 U425 ( .A(R2[31]), .B(n178), .Y(n343) );
  NAND3X1 U426 ( .A(n294), .B(n293), .C(n292), .Y(data_out[48]) );
  NAND2X1 U427 ( .A(data_in_1[48]), .B(n175), .Y(n293) );
  NAND2X1 U428 ( .A(data_in_2[48]), .B(n166), .Y(n294) );
  NAND2X1 U429 ( .A(R2[14]), .B(n181), .Y(n292) );
  NAND3X1 U430 ( .A(n445), .B(n444), .C(n443), .Y(data_out[99]) );
  NAND2X1 U431 ( .A(data_in_1[99]), .B(n173), .Y(n444) );
  NAND2X1 U432 ( .A(data_in_2[99]), .B(n163), .Y(n445) );
  NAND2X1 U433 ( .A(R3[31]), .B(n181), .Y(n443) );
  NAND3X1 U434 ( .A(n395), .B(n394), .C(n393), .Y(data_out[82]) );
  NAND2X1 U435 ( .A(data_in_1[82]), .B(n173), .Y(n394) );
  NAND2X1 U436 ( .A(data_in_2[82]), .B(n164), .Y(n395) );
  NAND2X1 U437 ( .A(R3[14]), .B(n181), .Y(n393) );
  NAND3X1 U438 ( .A(n544), .B(n543), .C(n542), .Y(data_out[133]) );
  NAND2X1 U439 ( .A(data_in_2[133]), .B(n161), .Y(n544) );
  NAND3X1 U440 ( .A(n495), .B(n494), .C(n493), .Y(data_out[116]) );
  NAND2X1 U441 ( .A(data_in_1[116]), .B(n172), .Y(n494) );
  NAND2X1 U442 ( .A(data_in_2[116]), .B(n162), .Y(n495) );
  NAND3X1 U443 ( .A(n348), .B(n347), .C(n346), .Y(data_out[66]) );
  NAND2X1 U444 ( .A(data_in_1[66]), .B(n174), .Y(n347) );
  NAND2X1 U445 ( .A(data_in_2[66]), .B(n165), .Y(n348) );
  NAND2X1 U446 ( .A(R2[32]), .B(n181), .Y(n346) );
  NAND3X1 U447 ( .A(n297), .B(n296), .C(n295), .Y(data_out[49]) );
  NAND2X1 U448 ( .A(data_in_1[49]), .B(n175), .Y(n296) );
  NAND2X1 U449 ( .A(R2[15]), .B(n179), .Y(n295) );
  NAND2X1 U450 ( .A(data_in_2[49]), .B(n166), .Y(n297) );
  NAND3X1 U451 ( .A(n448), .B(n447), .C(n446), .Y(data_out[100]) );
  NAND2X1 U452 ( .A(data_in_1[100]), .B(n172), .Y(n447) );
  NAND2X1 U453 ( .A(data_in_2[100]), .B(n163), .Y(n448) );
  NAND2X1 U454 ( .A(R3[32]), .B(n181), .Y(n446) );
  NAND3X1 U455 ( .A(n398), .B(n397), .C(n396), .Y(data_out[83]) );
  NAND2X1 U456 ( .A(data_in_1[83]), .B(n173), .Y(n397) );
  NAND2X1 U457 ( .A(R3[15]), .B(n546), .Y(n396) );
  NAND2X1 U458 ( .A(data_in_2[83]), .B(n164), .Y(n398) );
  NAND3X1 U459 ( .A(n549), .B(n548), .C(n547), .Y(data_out[134]) );
  NAND2X1 U460 ( .A(data_in_1[134]), .B(n171), .Y(n548) );
  NAND2X1 U461 ( .A(R4[32]), .B(n15), .Y(n547) );
  NAND2X1 U462 ( .A(data_in_2[134]), .B(n165), .Y(n549) );
  NAND3X1 U463 ( .A(n498), .B(n497), .C(n496), .Y(data_out[117]) );
  NAND2X1 U464 ( .A(data_in_1[117]), .B(n171), .Y(n497) );
  NAND2X1 U465 ( .A(R4[15]), .B(n181), .Y(n496) );
  NAND2X1 U466 ( .A(data_in_2[117]), .B(n162), .Y(n498) );
  NAND3X1 U467 ( .A(n252), .B(n251), .C(n250), .Y(data_out[35]) );
  NAND2XL U468 ( .A(R2[1]), .B(n178), .Y(n250) );
  NAND2X1 U469 ( .A(data_in_2[35]), .B(n162), .Y(n252) );
  NAND3X1 U470 ( .A(n356), .B(n355), .C(n354), .Y(data_out[69]) );
  NAND2X1 U471 ( .A(data_in_1[69]), .B(n174), .Y(n355) );
  NAND2X1 U472 ( .A(data_in_2[69]), .B(n165), .Y(n356) );
  NAND2X1 U473 ( .A(R3[1]), .B(n179), .Y(n354) );
  NAND3X1 U474 ( .A(n359), .B(n358), .C(n357), .Y(data_out[70]) );
  NAND2X1 U475 ( .A(data_in_1[70]), .B(n174), .Y(n358) );
  NAND2X1 U476 ( .A(data_in_2[70]), .B(n165), .Y(n359) );
  NAND2X1 U477 ( .A(R3[2]), .B(n15), .Y(n357) );
  NAND3X1 U478 ( .A(n258), .B(n257), .C(n256), .Y(data_out[37]) );
  NAND2X1 U479 ( .A(data_in_1[37]), .B(n174), .Y(n257) );
  NAND2XL U480 ( .A(R2[3]), .B(n181), .Y(n256) );
  NAND2X1 U481 ( .A(data_in_2[37]), .B(n161), .Y(n258) );
  NAND3X1 U482 ( .A(n511), .B(n510), .C(n509), .Y(data_out[122]) );
  NAND2X1 U483 ( .A(data_in_1[122]), .B(n171), .Y(n510) );
  NAND2X1 U484 ( .A(data_in_2[122]), .B(n161), .Y(n511) );
  NAND3X1 U485 ( .A(n406), .B(n405), .C(n404), .Y(data_out[86]) );
  NAND2X1 U486 ( .A(data_in_1[86]), .B(n173), .Y(n405) );
  NAND2X1 U487 ( .A(R3[18]), .B(n15), .Y(n404) );
  NAND2X1 U488 ( .A(data_in_2[86]), .B(n164), .Y(n406) );
  NAND3X1 U489 ( .A(n409), .B(n408), .C(n407), .Y(data_out[87]) );
  NAND2X1 U490 ( .A(data_in_1[87]), .B(n172), .Y(n408) );
  NAND2X1 U491 ( .A(R3[19]), .B(n180), .Y(n407) );
  NAND2X1 U492 ( .A(data_in_2[87]), .B(n164), .Y(n409) );
  NAND3X1 U493 ( .A(n412), .B(n411), .C(n410), .Y(data_out[88]) );
  NAND2X1 U494 ( .A(data_in_1[88]), .B(n175), .Y(n411) );
  NAND2X1 U495 ( .A(data_in_2[88]), .B(n164), .Y(n412) );
  NAND2X1 U496 ( .A(R3[20]), .B(n181), .Y(n410) );
  NAND3X1 U497 ( .A(n415), .B(n414), .C(n413), .Y(data_out[89]) );
  NAND2X1 U498 ( .A(data_in_1[89]), .B(n174), .Y(n414) );
  NAND2X1 U499 ( .A(data_in_2[89]), .B(n164), .Y(n415) );
  NAND2X1 U500 ( .A(R3[21]), .B(n546), .Y(n413) );
  NAND3X1 U501 ( .A(n418), .B(n417), .C(n416), .Y(data_out[90]) );
  NAND2X1 U502 ( .A(data_in_1[90]), .B(n173), .Y(n417) );
  NAND2X1 U503 ( .A(data_in_2[90]), .B(n164), .Y(n418) );
  NAND2X1 U504 ( .A(R3[22]), .B(n15), .Y(n416) );
  NAND3X1 U505 ( .A(n421), .B(n420), .C(n419), .Y(data_out[91]) );
  NAND2X1 U506 ( .A(data_in_1[91]), .B(n171), .Y(n420) );
  NAND2X1 U507 ( .A(data_in_2[91]), .B(n163), .Y(n421) );
  NAND2X1 U508 ( .A(R3[23]), .B(n15), .Y(n419) );
  NAND3X1 U509 ( .A(n424), .B(n423), .C(n422), .Y(data_out[92]) );
  NAND2X1 U510 ( .A(data_in_1[92]), .B(n172), .Y(n423) );
  NAND2X1 U511 ( .A(data_in_2[92]), .B(n163), .Y(n424) );
  NAND2X1 U512 ( .A(R3[24]), .B(n180), .Y(n422) );
  NAND3X1 U513 ( .A(n508), .B(n507), .C(n506), .Y(data_out[121]) );
  NAND2X1 U514 ( .A(data_in_1[121]), .B(n171), .Y(n507) );
  NAND2X1 U515 ( .A(R4[19]), .B(n178), .Y(n506) );
  NAND2X1 U516 ( .A(data_in_2[121]), .B(n161), .Y(n508) );
  NAND3X1 U517 ( .A(n306), .B(n305), .C(n304), .Y(data_out[52]) );
  NAND2X1 U518 ( .A(data_in_1[52]), .B(n175), .Y(n305) );
  NAND2X1 U519 ( .A(R2[18]), .B(n15), .Y(n304) );
  NAND2X1 U520 ( .A(data_in_2[52]), .B(n166), .Y(n306) );
  NAND3X1 U521 ( .A(n309), .B(n308), .C(n307), .Y(data_out[53]) );
  NAND2X1 U522 ( .A(data_in_1[53]), .B(n175), .Y(n308) );
  NAND2X1 U523 ( .A(R2[19]), .B(n182), .Y(n307) );
  NAND2X1 U524 ( .A(data_in_2[53]), .B(n166), .Y(n309) );
  OAI2BB1X1 U525 ( .A0N(data_in_2[51]), .A1N(n164), .B0(n303), .Y(data_out[51]) );
  OAI2BB1X1 U526 ( .A0N(data_in_2[34]), .A1N(n163), .B0(n249), .Y(data_out[34]) );
  OAI2BB1X1 U527 ( .A0N(data_in_2[85]), .A1N(n166), .B0(n403), .Y(data_out[85]) );
  OAI2BB1X1 U528 ( .A0N(data_in_2[68]), .A1N(n162), .B0(n353), .Y(data_out[68]) );
  NAND3X1 U529 ( .A(n505), .B(n504), .C(n503), .Y(data_out[120]) );
  NAND2X1 U530 ( .A(data_in_1[120]), .B(n171), .Y(n504) );
  NAND2X1 U531 ( .A(R4[18]), .B(n546), .Y(n503) );
  NAND2X1 U532 ( .A(data_in_2[120]), .B(n162), .Y(n505) );
  OAI2BB1X1 U533 ( .A0N(data_in_2[119]), .A1N(n161), .B0(n502), .Y(
        data_out[119]) );
  INVXL U534 ( .A(n10), .Y(n558) );
  AOI22XL U535 ( .A0(data_in_1[13]), .A1(n169), .B0(R1[13]), .B1(n182), .Y(
        n214) );
  NAND2X1 U536 ( .A(R2[13]), .B(n181), .Y(n289) );
  NAND2X1 U537 ( .A(R3[13]), .B(n181), .Y(n390) );
  NAND2X1 U538 ( .A(R4[13]), .B(n15), .Y(n490) );
  AOI22XL U539 ( .A0(data_in_1[16]), .A1(n169), .B0(R1[16]), .B1(n182), .Y(
        n217) );
  NAND2X2 U540 ( .A(n551), .B(n552), .Y(n554) );
  NOR4BXL U541 ( .AN(n14), .B(n557), .C(n558), .D(n3), .Y(n285) );
  NAND2XL U542 ( .A(n14), .B(n3), .Y(n282) );
  NOR3BX4 U543 ( .AN(counter[1]), .B(n2), .C(n10), .Y(n349) );
  OAI2BB1X4 U544 ( .A0N(data_in_2[0]), .A1N(n167), .B0(n196), .Y(data_out[0])
         );
  AOI22X4 U545 ( .A0(data_in_1[1]), .A1(n169), .B0(R1[1]), .B1(n15), .Y(n197)
         );
  OAI2BB1X4 U546 ( .A0N(data_in_2[1]), .A1N(n167), .B0(n197), .Y(data_out[1])
         );
  OAI2BB1X4 U547 ( .A0N(data_in_2[2]), .A1N(n243), .B0(n198), .Y(data_out[2])
         );
  OAI2BB1X4 U548 ( .A0N(data_in_2[3]), .A1N(n167), .B0(n199), .Y(data_out[3])
         );
  OAI2BB1X4 U549 ( .A0N(data_in_2[4]), .A1N(n167), .B0(n200), .Y(data_out[4])
         );
  OAI2BB1X4 U550 ( .A0N(data_in_2[17]), .A1N(n167), .B0(n218), .Y(data_out[17]) );
  OAI2BB1X4 U551 ( .A0N(data_in_2[18]), .A1N(n167), .B0(n219), .Y(data_out[18]) );
  NAND2BX4 U552 ( .AN(n223), .B(n222), .Y(data_out[19]) );
  OAI2BB1X4 U553 ( .A0N(data_in_2[20]), .A1N(n243), .B0(n224), .Y(data_out[20]) );
  OAI2BB1X4 U554 ( .A0N(data_in_2[21]), .A1N(n226), .B0(n225), .Y(data_out[21]) );
  NAND2BX4 U555 ( .AN(n230), .B(n229), .Y(data_out[22]) );
  OAI2BB1X4 U556 ( .A0N(data_in_2[23]), .A1N(n226), .B0(n231), .Y(data_out[23]) );
  OAI2BB1X4 U557 ( .A0N(data_in_2[25]), .A1N(n238), .B0(n237), .Y(data_out[25]) );
  OAI2BB1X4 U558 ( .A0N(data_in_2[26]), .A1N(n238), .B0(n239), .Y(data_out[26]) );
  OR2X4 U559 ( .A(n301), .B(n302), .Y(data_out[50]) );
endmodule


module multi16_0_DW01_add_5 ( A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, 
        A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, 
        A_4_, B_23_, B_22_, B_21_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, 
        B_14_, B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, 
        SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, 
        SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, 
        SUM_7_ );
  input A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_,
         A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, B_23_, B_22_,
         B_21_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_,
         B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_;
  output SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_,
         SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_,
         SUM_8_, SUM_7_;
  wire   n1, n2, n3, n4;
  wire   [23:7] carry;

  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry[7]), .CO(carry[8]), .S(SUM_7_)
         );
  ADDFX2 U1_21 ( .A(A_21_), .B(B_21_), .CI(carry[21]), .CO(carry[22]), .S(
        SUM_21_) );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry[20]), .CO(carry[21]), .S(
        SUM_20_) );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry[19]), .CO(carry[20]), .S(
        SUM_19_) );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry[18]), .CO(carry[19]), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry[17]), .CO(carry[18]), .S(
        SUM_17_) );
  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry[16]), .CO(carry[17]), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry[15]), .CO(carry[16]), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry[14]), .CO(carry[15]), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry[13]), .CO(carry[14]), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry[12]), .CO(carry[13]), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry[11]), .CO(carry[12]), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry[10]), .CO(carry[11]), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry[9]), .CO(carry[10]), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry[8]), .CO(carry[9]), .S(SUM_8_)
         );
  ADDFX2 U1_22 ( .A(A_22_), .B(B_22_), .CI(carry[22]), .CO(carry[23]), .S(
        SUM_22_) );
  AND2X2 U1 ( .A(A_4_), .B(B_4_), .Y(n1) );
  XOR2X1 U2 ( .A(B_23_), .B(carry[23]), .Y(SUM_23_) );
  OAI2BB1X1 U3 ( .A0N(n2), .A1N(A_6_), .B0(n3), .Y(carry[7]) );
  OAI21XL U4 ( .A0(A_6_), .A1(n2), .B0(B_6_), .Y(n3) );
  OAI2BB1X1 U5 ( .A0N(n1), .A1N(A_5_), .B0(n4), .Y(n2) );
  OAI21XL U6 ( .A0(A_5_), .A1(n1), .B0(B_5_), .Y(n4) );
endmodule


module multi16_0_DW01_add_3 ( A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, 
        A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, 
        B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, 
        B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, SUM_22_, SUM_21_, SUM_20_, 
        SUM_19_, SUM_18_, SUM_17_, SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, 
        SUM_11_, SUM_10_, SUM_9_, SUM_8_, SUM_7_ );
  input A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_,
         A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, B_20_, B_19_,
         B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, B_10_, B_9_,
         B_8_, B_7_, B_6_, B_5_;
  output SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_,
         SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_,
         SUM_7_;
  wire   carry_21_, carry_20_, carry_19_, carry_18_, carry_17_, carry_16_,
         carry_15_, carry_14_, carry_13_, carry_12_, carry_11_, carry_10_,
         carry_9_, carry_8_, carry_7_, n1;

  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry_16_), .CO(carry_17_), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry_15_), .CO(carry_16_), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry_14_), .CO(carry_15_), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry_13_), .CO(carry_14_), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry_12_), .CO(carry_13_), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry_11_), .CO(carry_12_), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry_10_), .CO(carry_11_), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry_9_), .CO(carry_10_), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry_8_), .CO(carry_9_), .S(SUM_8_)
         );
  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry_7_), .CO(carry_8_), .S(SUM_7_)
         );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry_20_), .CO(carry_21_), .S(
        SUM_20_) );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry_19_), .CO(carry_20_), .S(
        SUM_19_) );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry_18_), .CO(carry_19_), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry_17_), .CO(carry_18_), .S(
        SUM_17_) );
  ADDFX2 U1_21 ( .A(A_21_), .B(B_21_), .CI(carry_21_), .CO(SUM_22_), .S(
        SUM_21_) );
  OAI2BB1X1 U1 ( .A0N(A_6_), .A1N(B_6_), .B0(n1), .Y(carry_7_) );
  OAI211X1 U2 ( .A0(B_6_), .A1(A_6_), .B0(A_5_), .C0(B_5_), .Y(n1) );
endmodule


module multi16_0_DW01_add_0 ( A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, 
        A_16_, A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, 
        A_6_, A_5_, A_4_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, 
        B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, 
        SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, 
        SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, 
        SUM_7_ );
  input A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_,
         A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, B_20_,
         B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, B_10_,
         B_9_, B_8_, B_7_, B_6_, B_5_, B_4_;
  output SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_,
         SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_,
         SUM_8_, SUM_7_;
  wire   n1, n2, n3, n4, n5, n6;
  wire   [21:7] carry;

  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry[7]), .CO(carry[8]), .S(SUM_7_)
         );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry[18]), .CO(carry[19]), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry[17]), .CO(carry[18]), .S(
        SUM_17_) );
  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry[16]), .CO(carry[17]), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry[15]), .CO(carry[16]), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry[14]), .CO(carry[15]), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry[13]), .CO(carry[14]), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry[12]), .CO(carry[13]), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry[11]), .CO(carry[12]), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry[10]), .CO(carry[11]), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry[9]), .CO(carry[10]), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry[8]), .CO(carry[9]), .S(SUM_8_)
         );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry[19]), .CO(carry[20]), .S(
        SUM_19_) );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry[20]), .CO(carry[21]), .S(
        SUM_20_) );
  AND2X2 U1 ( .A(A_22_), .B(n2), .Y(n1) );
  AND2X2 U2 ( .A(A_21_), .B(carry[21]), .Y(n2) );
  AND2X2 U3 ( .A(A_4_), .B(B_4_), .Y(n3) );
  XOR2X1 U4 ( .A(A_23_), .B(n1), .Y(SUM_23_) );
  XOR2X1 U5 ( .A(A_21_), .B(carry[21]), .Y(SUM_21_) );
  XOR2X1 U6 ( .A(A_22_), .B(n2), .Y(SUM_22_) );
  OAI2BB1X1 U7 ( .A0N(n4), .A1N(A_6_), .B0(n5), .Y(carry[7]) );
  OAI21XL U8 ( .A0(A_6_), .A1(n4), .B0(B_6_), .Y(n5) );
  OAI2BB1X1 U9 ( .A0N(n3), .A1N(A_5_), .B0(n6), .Y(n4) );
  OAI21XL U10 ( .A0(A_5_), .A1(n3), .B0(B_5_), .Y(n6) );
endmodule


module multi16_0 ( in_17bit, in_8bit, out );
  input [16:0] in_17bit;
  input [7:0] in_8bit;
  output [16:0] out;
  wire   n197, n198, n199, n200, N14, N15, N16, N17, N18, N19, N20, N21, N22,
         N23, N24, N25, N26, N27, N28, N29, N108, N109, N110, N111, N112, N113,
         N114, N115, N116, N117, N118, N119, N120, N121, N122, N123, N205,
         N206, N207, N208, N209, N210, N211, N212, N213, N214, N215, N216,
         N217, N218, N219, N220, N221, N347, N348, N349, N350, N351, N352,
         N353, N354, N355, N356, N357, N358, N359, N360, N361, N362, N363,
         N446, N447, N448, N449, N450, N451, N452, N453, N454, N455, N456,
         N457, N458, N459, N460, N461, N462, N463, N477, N478, N479, N480,
         N481, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, add_2_root_r115_carry_10_,
         add_2_root_r115_carry_11_, add_2_root_r115_carry_12_,
         add_2_root_r115_carry_13_, add_2_root_r115_carry_14_,
         add_2_root_r115_carry_15_, add_2_root_r115_carry_16_,
         add_2_root_r115_carry_17_, add_2_root_r115_carry_18_,
         add_2_root_r115_carry_19_, add_2_root_r115_carry_4_,
         add_2_root_r115_carry_5_, add_2_root_r115_carry_6_,
         add_2_root_r115_carry_7_, add_2_root_r115_carry_8_,
         add_2_root_r115_carry_9_, add_2_root_r115_SUM_3_,
         add_2_root_r115_SUM_4_, add_2_root_r115_SUM_5_,
         add_2_root_r115_SUM_6_, add_2_root_r115_SUM_7_,
         add_2_root_r115_SUM_8_, add_2_root_r115_SUM_9_,
         add_2_root_r115_SUM_10_, add_2_root_r115_SUM_11_,
         add_2_root_r115_SUM_12_, add_2_root_r115_SUM_13_,
         add_2_root_r115_SUM_14_, add_2_root_r115_SUM_15_,
         add_2_root_r115_SUM_16_, add_2_root_r115_SUM_17_,
         add_2_root_r115_SUM_18_, add_2_root_r115_SUM_19_,
         add_2_root_r115_SUM_20_, add_1_root_r115_carry_10_,
         add_1_root_r115_carry_11_, add_1_root_r115_carry_12_,
         add_1_root_r115_carry_13_, add_1_root_r115_carry_14_,
         add_1_root_r115_carry_15_, add_1_root_r115_carry_16_,
         add_1_root_r115_carry_17_, add_1_root_r115_carry_18_,
         add_1_root_r115_carry_19_, add_1_root_r115_carry_20_,
         add_1_root_r115_carry_21_, add_1_root_r115_carry_22_,
         add_1_root_r115_carry_7_, add_1_root_r115_carry_8_,
         add_1_root_r115_carry_9_, add_1_root_r115_SUM_6_,
         add_1_root_r115_SUM_7_, add_1_root_r115_SUM_8_,
         add_1_root_r115_SUM_9_, add_1_root_r115_SUM_10_,
         add_1_root_r115_SUM_11_, add_1_root_r115_SUM_12_,
         add_1_root_r115_SUM_13_, add_1_root_r115_SUM_14_,
         add_1_root_r115_SUM_15_, add_1_root_r115_SUM_16_,
         add_1_root_r115_SUM_17_, add_1_root_r115_SUM_18_,
         add_1_root_r115_SUM_19_, add_1_root_r115_SUM_20_,
         add_1_root_r115_SUM_21_, add_1_root_r115_SUM_22_,
         add_1_root_r115_SUM_23_, add_1_root_r112_carry_10_,
         add_1_root_r112_carry_11_, add_1_root_r112_carry_12_,
         add_1_root_r112_carry_13_, add_1_root_r112_carry_14_,
         add_1_root_r112_carry_15_, add_1_root_r112_carry_16_,
         add_1_root_r112_carry_17_, add_1_root_r112_carry_18_,
         add_1_root_r112_carry_19_, add_1_root_r112_carry_20_,
         add_1_root_r112_carry_5_, add_1_root_r112_carry_6_,
         add_1_root_r112_carry_7_, add_1_root_r112_carry_8_,
         add_1_root_r112_carry_9_, add_1_root_r112_SUM_1_,
         add_1_root_r112_SUM_2_, add_1_root_r112_SUM_3_,
         add_1_root_r112_SUM_4_, add_1_root_r112_SUM_5_,
         add_1_root_r112_SUM_6_, add_1_root_r112_SUM_7_,
         add_1_root_r112_SUM_8_, add_1_root_r112_SUM_9_,
         add_1_root_r112_SUM_10_, add_1_root_r112_SUM_11_,
         add_1_root_r112_SUM_12_, add_1_root_r112_SUM_13_,
         add_1_root_r112_SUM_14_, add_1_root_r112_SUM_15_,
         add_1_root_r112_SUM_16_, add_1_root_r112_SUM_17_,
         add_1_root_r112_SUM_18_, add_1_root_r112_SUM_19_,
         add_1_root_r112_SUM_20_, add_1_root_r112_SUM_21_,
         add_2_root_r119_carry_10_, add_2_root_r119_carry_11_,
         add_2_root_r119_carry_12_, add_2_root_r119_carry_13_,
         add_2_root_r119_carry_14_, add_2_root_r119_carry_15_,
         add_2_root_r119_carry_16_, add_2_root_r119_carry_17_,
         add_2_root_r119_carry_18_, add_2_root_r119_carry_19_,
         add_2_root_r119_carry_20_, add_2_root_r119_carry_21_,
         add_2_root_r119_carry_6_, add_2_root_r119_carry_7_,
         add_2_root_r119_carry_8_, add_2_root_r119_carry_9_,
         add_2_root_r119_SUM_5_, add_2_root_r119_SUM_6_,
         add_2_root_r119_SUM_7_, add_2_root_r119_SUM_8_,
         add_2_root_r119_SUM_9_, add_2_root_r119_SUM_10_,
         add_2_root_r119_SUM_11_, add_2_root_r119_SUM_12_,
         add_2_root_r119_SUM_13_, add_2_root_r119_SUM_14_,
         add_2_root_r119_SUM_15_, add_2_root_r119_SUM_16_,
         add_2_root_r119_SUM_17_, add_2_root_r119_SUM_18_,
         add_2_root_r119_SUM_19_, add_2_root_r119_SUM_20_,
         add_2_root_r119_SUM_21_, add_2_root_r119_SUM_22_,
         add_1_root_r119_SUM_6_, add_1_root_r119_SUM_7_,
         add_1_root_r119_SUM_8_, add_1_root_r119_SUM_9_,
         add_1_root_r119_SUM_10_, add_1_root_r119_SUM_11_,
         add_1_root_r119_SUM_12_, add_1_root_r119_SUM_13_,
         add_1_root_r119_SUM_14_, add_1_root_r119_SUM_15_,
         add_1_root_r119_SUM_16_, add_1_root_r119_SUM_17_,
         add_1_root_r119_SUM_18_, add_1_root_r119_SUM_19_,
         add_1_root_r119_SUM_20_, add_1_root_r119_SUM_21_,
         add_1_root_r119_SUM_22_, add_1_root_r119_SUM_23_,
         add_1_root_r119_A_2_, add_1_root_r119_A_3_, add_1_root_r119_A_4_,
         add_1_root_r119_A_5_, add_1_root_r119_A_6_, add_1_root_r119_A_7_,
         add_1_root_r119_A_8_, add_1_root_r119_A_9_, add_1_root_r119_A_10_,
         add_1_root_r119_A_11_, add_1_root_r119_A_12_, add_1_root_r119_A_13_,
         add_1_root_r119_A_14_, add_1_root_r119_A_15_, add_1_root_r119_A_16_,
         add_1_root_r119_A_17_, add_1_root_r119_A_18_, add_1_root_r119_A_19_,
         add_3_root_r119_carry_10_, add_3_root_r119_carry_11_,
         add_3_root_r119_carry_12_, add_3_root_r119_carry_13_,
         add_3_root_r119_carry_14_, add_3_root_r119_carry_15_,
         add_3_root_r119_carry_16_, add_3_root_r119_carry_17_,
         add_3_root_r119_carry_18_, add_3_root_r119_carry_3_,
         add_3_root_r119_carry_4_, add_3_root_r119_carry_5_,
         add_3_root_r119_carry_6_, add_3_root_r119_carry_7_,
         add_3_root_r119_carry_8_, add_3_root_r119_carry_9_, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n170, n171, n172, n173, n174, n175, n176,
         n177;
  wire   [16:0] in_17bit_b;
  wire   [23:8] neg_mul;
  wire   [16:11] sub_add_75_b0_carry;
  wire   [16:2] sub_add_54_b0_carry;
  wire   [22:7] add_1_root_r119_carry;

  multi16_0_DW01_add_5 add_0_root_r119 ( .A_22_(add_2_root_r119_SUM_22_), 
        .A_21_(add_2_root_r119_SUM_21_), .A_20_(add_2_root_r119_SUM_20_), 
        .A_19_(add_2_root_r119_SUM_19_), .A_18_(add_2_root_r119_SUM_18_), 
        .A_17_(add_2_root_r119_SUM_17_), .A_16_(add_2_root_r119_SUM_16_), 
        .A_15_(add_2_root_r119_SUM_15_), .A_14_(add_2_root_r119_SUM_14_), 
        .A_13_(add_2_root_r119_SUM_13_), .A_12_(add_2_root_r119_SUM_12_), 
        .A_11_(add_2_root_r119_SUM_11_), .A_10_(add_2_root_r119_SUM_10_), 
        .A_9_(add_2_root_r119_SUM_9_), .A_8_(add_2_root_r119_SUM_8_), .A_7_(
        add_2_root_r119_SUM_7_), .A_6_(add_2_root_r119_SUM_6_), .A_5_(
        add_2_root_r119_SUM_5_), .A_4_(in_17bit_b[0]), .B_23_(
        add_1_root_r119_SUM_23_), .B_22_(add_1_root_r119_SUM_22_), .B_21_(
        add_1_root_r119_SUM_21_), .B_20_(add_1_root_r119_SUM_20_), .B_19_(
        add_1_root_r119_SUM_19_), .B_18_(add_1_root_r119_SUM_18_), .B_17_(
        add_1_root_r119_SUM_17_), .B_16_(add_1_root_r119_SUM_16_), .B_15_(
        add_1_root_r119_SUM_15_), .B_14_(add_1_root_r119_SUM_14_), .B_13_(
        add_1_root_r119_SUM_13_), .B_12_(add_1_root_r119_SUM_12_), .B_11_(
        add_1_root_r119_SUM_11_), .B_10_(add_1_root_r119_SUM_10_), .B_9_(
        add_1_root_r119_SUM_9_), .B_8_(add_1_root_r119_SUM_8_), .B_7_(
        add_1_root_r119_SUM_7_), .B_6_(add_1_root_r119_SUM_6_), .B_5_(
        add_1_root_r119_A_5_), .B_4_(add_1_root_r119_A_4_), .SUM_23_(N363), 
        .SUM_22_(N362), .SUM_21_(N361), .SUM_20_(N360), .SUM_19_(N359), 
        .SUM_18_(N358), .SUM_17_(N357), .SUM_16_(N356), .SUM_15_(N355), 
        .SUM_14_(N354), .SUM_13_(N353), .SUM_12_(N352), .SUM_11_(N351), 
        .SUM_10_(N350), .SUM_9_(N349), .SUM_8_(N348), .SUM_7_(N347) );
  multi16_0_DW01_add_3 add_0_root_r112 ( .A_21_(n42), .A_20_(in_17bit_b[15]), 
        .A_19_(in_17bit_b[14]), .A_18_(in_17bit_b[13]), .A_17_(in_17bit_b[12]), 
        .A_16_(in_17bit_b[11]), .A_15_(in_17bit_b[10]), .A_14_(in_17bit_b[9]), 
        .A_13_(in_17bit_b[8]), .A_12_(in_17bit_b[7]), .A_11_(in_17bit_b[6]), 
        .A_10_(in_17bit_b[5]), .A_9_(in_17bit_b[4]), .A_8_(in_17bit_b[3]), 
        .A_7_(in_17bit_b[2]), .A_6_(in_17bit_b[1]), .A_5_(in_17bit_b[0]), 
        .B_21_(add_1_root_r112_SUM_21_), .B_20_(add_1_root_r112_SUM_20_), 
        .B_19_(add_1_root_r112_SUM_19_), .B_18_(add_1_root_r112_SUM_18_), 
        .B_17_(add_1_root_r112_SUM_17_), .B_16_(add_1_root_r112_SUM_16_), 
        .B_15_(add_1_root_r112_SUM_15_), .B_14_(add_1_root_r112_SUM_14_), 
        .B_13_(add_1_root_r112_SUM_13_), .B_12_(add_1_root_r112_SUM_12_), 
        .B_11_(add_1_root_r112_SUM_11_), .B_10_(add_1_root_r112_SUM_10_), 
        .B_9_(add_1_root_r112_SUM_9_), .B_8_(add_1_root_r112_SUM_8_), .B_7_(
        add_1_root_r112_SUM_7_), .B_6_(add_1_root_r112_SUM_6_), .B_5_(
        add_1_root_r112_SUM_5_), .SUM_22_(N123), .SUM_21_(N122), .SUM_20_(N121), .SUM_19_(N120), .SUM_18_(N119), .SUM_17_(N118), .SUM_16_(N117), .SUM_15_(
        N116), .SUM_14_(N115), .SUM_13_(N114), .SUM_12_(N113), .SUM_11_(N112), 
        .SUM_10_(N111), .SUM_9_(N110), .SUM_8_(N109), .SUM_7_(N108) );
  multi16_0_DW01_add_0 add_0_root_r115 ( .A_23_(add_1_root_r115_SUM_23_), 
        .A_22_(add_1_root_r115_SUM_22_), .A_21_(add_1_root_r115_SUM_21_), 
        .A_20_(add_1_root_r115_SUM_20_), .A_19_(add_1_root_r115_SUM_19_), 
        .A_18_(add_1_root_r115_SUM_18_), .A_17_(add_1_root_r115_SUM_17_), 
        .A_16_(add_1_root_r115_SUM_16_), .A_15_(add_1_root_r115_SUM_15_), 
        .A_14_(add_1_root_r115_SUM_14_), .A_13_(add_1_root_r115_SUM_13_), 
        .A_12_(add_1_root_r115_SUM_12_), .A_11_(add_1_root_r115_SUM_11_), 
        .A_10_(add_1_root_r115_SUM_10_), .A_9_(add_1_root_r115_SUM_9_), .A_8_(
        add_1_root_r115_SUM_8_), .A_7_(add_1_root_r115_SUM_7_), .A_6_(
        add_1_root_r115_SUM_6_), .A_5_(in_17bit_b[1]), .A_4_(in_17bit_b[0]), 
        .B_20_(add_2_root_r115_SUM_20_), .B_19_(add_2_root_r115_SUM_19_), 
        .B_18_(add_2_root_r115_SUM_18_), .B_17_(add_2_root_r115_SUM_17_), 
        .B_16_(add_2_root_r115_SUM_16_), .B_15_(add_2_root_r115_SUM_15_), 
        .B_14_(add_2_root_r115_SUM_14_), .B_13_(add_2_root_r115_SUM_13_), 
        .B_12_(add_2_root_r115_SUM_12_), .B_11_(add_2_root_r115_SUM_11_), 
        .B_10_(add_2_root_r115_SUM_10_), .B_9_(add_2_root_r115_SUM_9_), .B_8_(
        add_2_root_r115_SUM_8_), .B_7_(add_2_root_r115_SUM_7_), .B_6_(
        add_2_root_r115_SUM_6_), .B_5_(add_2_root_r115_SUM_5_), .B_4_(
        add_2_root_r115_SUM_4_), .SUM_23_(N221), .SUM_22_(N220), .SUM_21_(N219), .SUM_20_(N218), .SUM_19_(N217), .SUM_18_(N216), .SUM_17_(N215), .SUM_16_(
        N214), .SUM_15_(N213), .SUM_14_(N212), .SUM_13_(N211), .SUM_12_(N210), 
        .SUM_11_(N209), .SUM_10_(N208), .SUM_9_(N207), .SUM_8_(N206), .SUM_7_(
        N205) );
  TLATX1 neg_mul_reg_17_ ( .G(N446), .D(N457), .QN(n7) );
  TLATX1 neg_mul_reg_16_ ( .G(N446), .D(N456), .QN(n5) );
  TLATX1 neg_mul_reg_15_ ( .G(N446), .D(N455), .QN(n3) );
  TLATX1 neg_mul_reg_14_ ( .G(N446), .D(N454), .QN(n4) );
  TLATX1 neg_mul_reg_13_ ( .G(N446), .D(N453), .Q(neg_mul[13]), .QN(n16) );
  TLATX1 neg_mul_reg_12_ ( .G(N446), .D(N452), .QN(n6) );
  TLATX1 neg_mul_reg_11_ ( .G(N446), .D(N451), .Q(neg_mul[11]), .QN(n15) );
  TLATX1 neg_mul_reg_23_ ( .G(N446), .D(N463), .Q(neg_mul[23]), .QN(n13) );
  TLATX1 neg_mul_reg_22_ ( .G(N446), .D(N462), .Q(neg_mul[22]), .QN(n10) );
  TLATX1 neg_mul_reg_21_ ( .G(N446), .D(N461), .Q(neg_mul[21]), .QN(n8) );
  TLATX1 neg_mul_reg_20_ ( .G(N446), .D(N460), .Q(neg_mul[20]), .QN(n9) );
  TLATX1 neg_mul_reg_19_ ( .G(N446), .D(N459), .Q(neg_mul[19]), .QN(n11) );
  TLATX1 neg_mul_reg_18_ ( .G(N446), .D(N458), .QN(n12) );
  TLATX1 neg_mul_reg_8_ ( .G(N446), .D(N448), .Q(neg_mul[8]) );
  TLATX1 neg_mul_reg_9_ ( .G(N446), .D(N449), .Q(neg_mul[9]), .QN(n14) );
  TLATX1 neg_mul_reg_10_ ( .G(N446), .D(N450), .Q(neg_mul[10]) );
  TLATX1 neg_mul_reg_7_ ( .G(N446), .D(N447), .Q(out[0]) );
  BUFX12 U2 ( .A(n30), .Y(n2) );
  BUFX8 U3 ( .A(n199), .Y(out[2]) );
  BUFX4 U4 ( .A(n197), .Y(out[12]) );
  INVX1 U5 ( .A(n67), .Y(n18) );
  MX2X1 U6 ( .A(neg_mul[21]), .B(N479), .S0(n2), .Y(out[14]) );
  MX2X1 U7 ( .A(neg_mul[20]), .B(N478), .S0(n2), .Y(out[13]) );
  BUFX4 U8 ( .A(n198), .Y(out[3]) );
  CLKINVX3 U9 ( .A(n39), .Y(n49) );
  INVX4 U10 ( .A(n53), .Y(n39) );
  XOR2X4 U11 ( .A(n49), .B(in_8bit[7]), .Y(n30) );
  INVXL U12 ( .A(n49), .Y(n54) );
  XNOR2X2 U13 ( .A(n53), .B(in_8bit[7]), .Y(n88) );
  XOR2X4 U14 ( .A(n84), .B(neg_mul[13]), .Y(out[6]) );
  BUFX12 U15 ( .A(n200), .Y(out[1]) );
  INVX2 U16 ( .A(in_17bit[16]), .Y(n17) );
  XOR2X4 U17 ( .A(n80), .B(neg_mul[11]), .Y(out[4]) );
  INVX8 U18 ( .A(n50), .Y(n38) );
  INVX8 U19 ( .A(n50), .Y(n53) );
  NOR2X4 U20 ( .A(n28), .B(n86), .Y(n87) );
  NOR2X1 U21 ( .A(n76), .B(in_17bit[16]), .Y(n77) );
  AND2X4 U22 ( .A(n17), .B(n18), .Y(n69) );
  CLKINVX2 U23 ( .A(n50), .Y(n52) );
  XNOR2X4 U24 ( .A(n53), .B(in_8bit[7]), .Y(n81) );
  AOI211X2 U25 ( .A0(n53), .A1(n62), .B0(n61), .C0(n32), .Y(n200) );
  NOR2X4 U26 ( .A(n23), .B(n81), .Y(n82) );
  AOI211X2 U27 ( .A0(n38), .A1(n70), .B0(n69), .C0(n68), .Y(n199) );
  OR2X4 U28 ( .A(n26), .B(n85), .Y(n20) );
  XNOR2X4 U29 ( .A(n53), .B(in_8bit[7]), .Y(n85) );
  INVX8 U30 ( .A(in_17bit[16]), .Y(n50) );
  INVXL U31 ( .A(n48), .Y(n55) );
  INVXL U32 ( .A(in_8bit[0]), .Y(n47) );
  INVX1 U33 ( .A(n152), .Y(in_17bit_b[1]) );
  INVX1 U34 ( .A(n113), .Y(in_17bit_b[14]) );
  INVX1 U35 ( .A(n116), .Y(in_17bit_b[13]) );
  INVX1 U36 ( .A(n149), .Y(in_17bit_b[2]) );
  INVX1 U37 ( .A(n140), .Y(in_17bit_b[5]) );
  INVX1 U38 ( .A(n137), .Y(in_17bit_b[6]) );
  INVX1 U39 ( .A(n134), .Y(in_17bit_b[7]) );
  INVX1 U40 ( .A(n131), .Y(in_17bit_b[8]) );
  INVX1 U41 ( .A(n128), .Y(in_17bit_b[9]) );
  INVX1 U42 ( .A(n125), .Y(in_17bit_b[10]) );
  INVX1 U43 ( .A(n122), .Y(in_17bit_b[11]) );
  INVX1 U44 ( .A(n119), .Y(in_17bit_b[12]) );
  INVX1 U45 ( .A(n143), .Y(in_17bit_b[4]) );
  INVX1 U46 ( .A(n146), .Y(in_17bit_b[3]) );
  XOR2X4 U47 ( .A(n20), .B(n5), .Y(out[9]) );
  XOR2X4 U48 ( .A(n21), .B(n3), .Y(out[8]) );
  OR2X4 U49 ( .A(n88), .B(n27), .Y(n21) );
  XOR2X4 U50 ( .A(n22), .B(n4), .Y(out[7]) );
  OR2X4 U51 ( .A(n25), .B(n85), .Y(n22) );
  INVX1 U52 ( .A(n54), .Y(n48) );
  INVX1 U53 ( .A(n47), .Y(n46) );
  ADDFX2 U54 ( .A(n42), .B(in_17bit_b[12]), .CI(add_1_root_r112_carry_16_), 
        .CO(add_1_root_r112_carry_17_), .S(add_1_root_r112_SUM_16_) );
  ADDFX2 U55 ( .A(add_1_root_r119_A_19_), .B(in_17bit_b[13]), .CI(
        add_1_root_r119_carry[19]), .CO(add_1_root_r119_carry[20]), .S(
        add_1_root_r119_SUM_19_) );
  ADDFX2 U56 ( .A(n42), .B(in_17bit_b[15]), .CI(add_3_root_r119_carry_17_), 
        .CO(add_3_root_r119_carry_18_), .S(add_1_root_r119_A_17_) );
  ADDFX2 U57 ( .A(n42), .B(in_17bit_b[14]), .CI(add_2_root_r115_carry_17_), 
        .CO(add_2_root_r115_carry_18_), .S(add_2_root_r115_SUM_17_) );
  ADDFX2 U58 ( .A(n42), .B(in_17bit_b[14]), .CI(add_1_root_r115_carry_20_), 
        .CO(add_1_root_r115_carry_21_), .S(add_1_root_r115_SUM_20_) );
  ADDFX2 U59 ( .A(n42), .B(in_17bit_b[15]), .CI(add_2_root_r119_carry_20_), 
        .CO(add_2_root_r119_carry_21_), .S(add_2_root_r119_SUM_20_) );
  INVX1 U60 ( .A(n55), .Y(n51) );
  ADDFX2 U61 ( .A(in_17bit_b[3]), .B(in_17bit_b[1]), .CI(
        add_2_root_r115_carry_4_), .CO(add_2_root_r115_carry_5_), .S(
        add_2_root_r115_SUM_4_) );
  ADDFX2 U62 ( .A(in_17bit_b[4]), .B(in_17bit_b[2]), .CI(
        add_2_root_r115_carry_5_), .CO(add_2_root_r115_carry_6_), .S(
        add_2_root_r115_SUM_5_) );
  ADDFX2 U63 ( .A(in_17bit_b[5]), .B(in_17bit_b[1]), .CI(
        add_1_root_r112_carry_5_), .CO(add_1_root_r112_carry_6_), .S(
        add_1_root_r112_SUM_5_) );
  ADDFX2 U64 ( .A(in_17bit_b[6]), .B(in_17bit_b[5]), .CI(
        add_3_root_r119_carry_7_), .CO(add_3_root_r119_carry_8_), .S(
        add_1_root_r119_A_7_) );
  ADDFX2 U65 ( .A(in_17bit_b[6]), .B(in_17bit_b[2]), .CI(
        add_1_root_r112_carry_6_), .CO(add_1_root_r112_carry_7_), .S(
        add_1_root_r112_SUM_6_) );
  ADDFX2 U66 ( .A(in_17bit_b[3]), .B(in_17bit_b[1]), .CI(
        add_1_root_r115_carry_7_), .CO(add_1_root_r115_carry_8_), .S(
        add_1_root_r115_SUM_7_) );
  ADDFX2 U67 ( .A(in_17bit_b[7]), .B(in_17bit_b[6]), .CI(
        add_3_root_r119_carry_8_), .CO(add_3_root_r119_carry_9_), .S(
        add_1_root_r119_A_8_) );
  ADDFX2 U68 ( .A(add_1_root_r119_A_7_), .B(in_17bit_b[1]), .CI(
        add_1_root_r119_carry[7]), .CO(add_1_root_r119_carry[8]), .S(
        add_1_root_r119_SUM_7_) );
  ADDFX2 U69 ( .A(in_17bit_b[2]), .B(in_17bit_b[1]), .CI(
        add_2_root_r119_carry_6_), .CO(add_2_root_r119_carry_7_), .S(
        add_2_root_r119_SUM_6_) );
  ADDFX2 U70 ( .A(in_17bit_b[4]), .B(in_17bit_b[2]), .CI(
        add_1_root_r115_carry_8_), .CO(add_1_root_r115_carry_9_), .S(
        add_1_root_r115_SUM_8_) );
  ADDFX2 U71 ( .A(in_17bit_b[8]), .B(in_17bit_b[7]), .CI(
        add_3_root_r119_carry_9_), .CO(add_3_root_r119_carry_10_), .S(
        add_1_root_r119_A_9_) );
  ADDFX2 U72 ( .A(in_17bit_b[3]), .B(in_17bit_b[2]), .CI(
        add_2_root_r119_carry_7_), .CO(add_2_root_r119_carry_8_), .S(
        add_2_root_r119_SUM_7_) );
  ADDFX2 U73 ( .A(in_17bit_b[6]), .B(in_17bit_b[4]), .CI(
        add_2_root_r115_carry_7_), .CO(add_2_root_r115_carry_8_), .S(
        add_2_root_r115_SUM_7_) );
  ADDFX2 U74 ( .A(in_17bit_b[8]), .B(in_17bit_b[4]), .CI(
        add_1_root_r112_carry_8_), .CO(add_1_root_r112_carry_9_), .S(
        add_1_root_r112_SUM_8_) );
  ADDFX2 U75 ( .A(in_17bit_b[9]), .B(in_17bit_b[8]), .CI(
        add_3_root_r119_carry_10_), .CO(add_3_root_r119_carry_11_), .S(
        add_1_root_r119_A_10_) );
  ADDFX2 U76 ( .A(in_17bit_b[7]), .B(in_17bit_b[5]), .CI(
        add_2_root_r115_carry_8_), .CO(add_2_root_r115_carry_9_), .S(
        add_2_root_r115_SUM_8_) );
  ADDFX2 U77 ( .A(in_17bit_b[9]), .B(in_17bit_b[5]), .CI(
        add_1_root_r112_carry_9_), .CO(add_1_root_r112_carry_10_), .S(
        add_1_root_r112_SUM_9_) );
  ADDFX2 U78 ( .A(in_17bit_b[6]), .B(in_17bit_b[4]), .CI(
        add_1_root_r115_carry_10_), .CO(add_1_root_r115_carry_11_), .S(
        add_1_root_r115_SUM_10_) );
  ADDFX2 U79 ( .A(in_17bit_b[10]), .B(in_17bit_b[9]), .CI(
        add_3_root_r119_carry_11_), .CO(add_3_root_r119_carry_12_), .S(
        add_1_root_r119_A_11_) );
  ADDFX2 U80 ( .A(add_1_root_r119_A_10_), .B(in_17bit_b[4]), .CI(
        add_1_root_r119_carry[10]), .CO(add_1_root_r119_carry[11]), .S(
        add_1_root_r119_SUM_10_) );
  ADDFX2 U81 ( .A(in_17bit_b[8]), .B(in_17bit_b[6]), .CI(
        add_2_root_r115_carry_9_), .CO(add_2_root_r115_carry_10_), .S(
        add_2_root_r115_SUM_9_) );
  ADDFX2 U82 ( .A(in_17bit_b[10]), .B(in_17bit_b[6]), .CI(
        add_1_root_r112_carry_10_), .CO(add_1_root_r112_carry_11_), .S(
        add_1_root_r112_SUM_10_) );
  ADDFX2 U83 ( .A(in_17bit_b[7]), .B(in_17bit_b[5]), .CI(
        add_1_root_r115_carry_11_), .CO(add_1_root_r115_carry_12_), .S(
        add_1_root_r115_SUM_11_) );
  ADDFX2 U84 ( .A(in_17bit_b[6]), .B(in_17bit_b[5]), .CI(
        add_2_root_r119_carry_10_), .CO(add_2_root_r119_carry_11_), .S(
        add_2_root_r119_SUM_10_) );
  ADDFX2 U85 ( .A(in_17bit_b[11]), .B(in_17bit_b[7]), .CI(
        add_1_root_r112_carry_11_), .CO(add_1_root_r112_carry_12_), .S(
        add_1_root_r112_SUM_11_) );
  ADDFX2 U86 ( .A(in_17bit_b[8]), .B(in_17bit_b[6]), .CI(
        add_1_root_r115_carry_12_), .CO(add_1_root_r115_carry_13_), .S(
        add_1_root_r115_SUM_12_) );
  ADDFX2 U87 ( .A(in_17bit_b[12]), .B(in_17bit_b[11]), .CI(
        add_3_root_r119_carry_13_), .CO(add_3_root_r119_carry_14_), .S(
        add_1_root_r119_A_13_) );
  ADDFX2 U88 ( .A(in_17bit_b[7]), .B(in_17bit_b[6]), .CI(
        add_2_root_r119_carry_11_), .CO(add_2_root_r119_carry_12_), .S(
        add_2_root_r119_SUM_11_) );
  ADDFX2 U89 ( .A(in_17bit_b[10]), .B(in_17bit_b[8]), .CI(
        add_2_root_r115_carry_11_), .CO(add_2_root_r115_carry_12_), .S(
        add_2_root_r115_SUM_11_) );
  ADDFX2 U90 ( .A(in_17bit_b[12]), .B(in_17bit_b[8]), .CI(
        add_1_root_r112_carry_12_), .CO(add_1_root_r112_carry_13_), .S(
        add_1_root_r112_SUM_12_) );
  ADDFX2 U91 ( .A(in_17bit_b[9]), .B(in_17bit_b[7]), .CI(
        add_1_root_r115_carry_13_), .CO(add_1_root_r115_carry_14_), .S(
        add_1_root_r115_SUM_13_) );
  ADDFX2 U92 ( .A(in_17bit_b[13]), .B(in_17bit_b[12]), .CI(
        add_3_root_r119_carry_14_), .CO(add_3_root_r119_carry_15_), .S(
        add_1_root_r119_A_14_) );
  ADDFX2 U93 ( .A(add_1_root_r119_A_13_), .B(in_17bit_b[7]), .CI(
        add_1_root_r119_carry[13]), .CO(add_1_root_r119_carry[14]), .S(
        add_1_root_r119_SUM_13_) );
  ADDFX2 U94 ( .A(in_17bit_b[8]), .B(in_17bit_b[7]), .CI(
        add_2_root_r119_carry_12_), .CO(add_2_root_r119_carry_13_), .S(
        add_2_root_r119_SUM_12_) );
  ADDFX2 U95 ( .A(in_17bit_b[11]), .B(in_17bit_b[9]), .CI(
        add_2_root_r115_carry_12_), .CO(add_2_root_r115_carry_13_), .S(
        add_2_root_r115_SUM_12_) );
  ADDFX2 U96 ( .A(in_17bit_b[13]), .B(in_17bit_b[9]), .CI(
        add_1_root_r112_carry_13_), .CO(add_1_root_r112_carry_14_), .S(
        add_1_root_r112_SUM_13_) );
  ADDFX2 U97 ( .A(in_17bit_b[10]), .B(in_17bit_b[8]), .CI(
        add_1_root_r115_carry_14_), .CO(add_1_root_r115_carry_15_), .S(
        add_1_root_r115_SUM_14_) );
  ADDFX2 U98 ( .A(in_17bit_b[14]), .B(in_17bit_b[13]), .CI(
        add_3_root_r119_carry_15_), .CO(add_3_root_r119_carry_16_), .S(
        add_1_root_r119_A_15_) );
  ADDFX2 U99 ( .A(add_1_root_r119_A_14_), .B(in_17bit_b[8]), .CI(
        add_1_root_r119_carry[14]), .CO(add_1_root_r119_carry[15]), .S(
        add_1_root_r119_SUM_14_) );
  ADDFX2 U100 ( .A(in_17bit_b[9]), .B(in_17bit_b[8]), .CI(
        add_2_root_r119_carry_13_), .CO(add_2_root_r119_carry_14_), .S(
        add_2_root_r119_SUM_13_) );
  ADDFX2 U101 ( .A(in_17bit_b[12]), .B(in_17bit_b[10]), .CI(
        add_2_root_r115_carry_13_), .CO(add_2_root_r115_carry_14_), .S(
        add_2_root_r115_SUM_13_) );
  ADDFX2 U102 ( .A(in_17bit_b[14]), .B(in_17bit_b[10]), .CI(
        add_1_root_r112_carry_14_), .CO(add_1_root_r112_carry_15_), .S(
        add_1_root_r112_SUM_14_) );
  ADDFX2 U103 ( .A(in_17bit_b[11]), .B(in_17bit_b[9]), .CI(
        add_1_root_r115_carry_15_), .CO(add_1_root_r115_carry_16_), .S(
        add_1_root_r115_SUM_15_) );
  ADDFX2 U104 ( .A(add_1_root_r119_A_15_), .B(in_17bit_b[9]), .CI(
        add_1_root_r119_carry[15]), .CO(add_1_root_r119_carry[16]), .S(
        add_1_root_r119_SUM_15_) );
  ADDFX2 U105 ( .A(in_17bit_b[3]), .B(in_17bit_b[2]), .CI(
        add_3_root_r119_carry_4_), .CO(add_3_root_r119_carry_5_), .S(
        add_1_root_r119_A_4_) );
  ADDFX2 U106 ( .A(in_17bit_b[2]), .B(in_17bit_b[1]), .CI(
        add_3_root_r119_carry_3_), .CO(add_3_root_r119_carry_4_), .S(
        add_1_root_r119_A_3_) );
  ADDFX2 U107 ( .A(in_17bit_b[10]), .B(in_17bit_b[9]), .CI(
        add_2_root_r119_carry_14_), .CO(add_2_root_r119_carry_15_), .S(
        add_2_root_r119_SUM_14_) );
  ADDFX2 U108 ( .A(in_17bit_b[13]), .B(in_17bit_b[11]), .CI(
        add_2_root_r115_carry_14_), .CO(add_2_root_r115_carry_15_), .S(
        add_2_root_r115_SUM_14_) );
  ADDFX2 U109 ( .A(in_17bit_b[15]), .B(in_17bit_b[11]), .CI(
        add_1_root_r112_carry_15_), .CO(add_1_root_r112_carry_16_), .S(
        add_1_root_r112_SUM_15_) );
  ADDFX2 U110 ( .A(in_17bit_b[12]), .B(in_17bit_b[10]), .CI(
        add_1_root_r115_carry_16_), .CO(add_1_root_r115_carry_17_), .S(
        add_1_root_r115_SUM_16_) );
  ADDFX2 U111 ( .A(add_1_root_r119_A_16_), .B(in_17bit_b[10]), .CI(
        add_1_root_r119_carry[16]), .CO(add_1_root_r119_carry[17]), .S(
        add_1_root_r119_SUM_16_) );
  ADDFX2 U112 ( .A(in_17bit_b[11]), .B(in_17bit_b[10]), .CI(
        add_2_root_r119_carry_15_), .CO(add_2_root_r119_carry_16_), .S(
        add_2_root_r119_SUM_15_) );
  ADDFX2 U113 ( .A(in_17bit_b[14]), .B(in_17bit_b[12]), .CI(
        add_2_root_r115_carry_15_), .CO(add_2_root_r115_carry_16_), .S(
        add_2_root_r115_SUM_15_) );
  ADDFX2 U114 ( .A(in_17bit_b[13]), .B(in_17bit_b[11]), .CI(
        add_1_root_r115_carry_17_), .CO(add_1_root_r115_carry_18_), .S(
        add_1_root_r115_SUM_17_) );
  ADDFX2 U115 ( .A(add_1_root_r119_A_17_), .B(in_17bit_b[11]), .CI(
        add_1_root_r119_carry[17]), .CO(add_1_root_r119_carry[18]), .S(
        add_1_root_r119_SUM_17_) );
  ADDFX2 U116 ( .A(in_17bit_b[12]), .B(in_17bit_b[11]), .CI(
        add_2_root_r119_carry_16_), .CO(add_2_root_r119_carry_17_), .S(
        add_2_root_r119_SUM_16_) );
  ADDFX2 U117 ( .A(in_17bit_b[14]), .B(in_17bit_b[12]), .CI(
        add_1_root_r115_carry_18_), .CO(add_1_root_r115_carry_19_), .S(
        add_1_root_r115_SUM_18_) );
  ADDFX2 U118 ( .A(add_1_root_r119_A_18_), .B(in_17bit_b[12]), .CI(
        add_1_root_r119_carry[18]), .CO(add_1_root_r119_carry[19]), .S(
        add_1_root_r119_SUM_18_) );
  ADDFX2 U119 ( .A(in_17bit_b[13]), .B(in_17bit_b[12]), .CI(
        add_2_root_r119_carry_17_), .CO(add_2_root_r119_carry_18_), .S(
        add_2_root_r119_SUM_17_) );
  ADDFX2 U120 ( .A(add_1_root_r119_A_8_), .B(in_17bit_b[2]), .CI(
        add_1_root_r119_carry[8]), .CO(add_1_root_r119_carry[9]), .S(
        add_1_root_r119_SUM_8_) );
  ADDFX2 U121 ( .A(in_17bit_b[11]), .B(in_17bit_b[10]), .CI(
        add_3_root_r119_carry_12_), .CO(add_3_root_r119_carry_13_), .S(
        add_1_root_r119_A_12_) );
  ADDFX2 U122 ( .A(in_17bit_b[15]), .B(in_17bit_b[13]), .CI(
        add_2_root_r115_carry_16_), .CO(add_2_root_r115_carry_17_), .S(
        add_2_root_r115_SUM_16_) );
  ADDFX2 U123 ( .A(in_17bit_b[15]), .B(in_17bit_b[13]), .CI(
        add_1_root_r115_carry_19_), .CO(add_1_root_r115_carry_20_), .S(
        add_1_root_r115_SUM_19_) );
  ADDFX2 U124 ( .A(in_17bit_b[5]), .B(in_17bit_b[3]), .CI(
        add_2_root_r115_carry_6_), .CO(add_2_root_r115_carry_7_), .S(
        add_2_root_r115_SUM_6_) );
  ADDFX2 U125 ( .A(in_17bit_b[7]), .B(in_17bit_b[3]), .CI(
        add_1_root_r112_carry_7_), .CO(add_1_root_r112_carry_8_), .S(
        add_1_root_r112_SUM_7_) );
  ADDFX2 U126 ( .A(in_17bit_b[5]), .B(in_17bit_b[3]), .CI(
        add_1_root_r115_carry_9_), .CO(add_1_root_r115_carry_10_), .S(
        add_1_root_r115_SUM_9_) );
  ADDFX2 U127 ( .A(in_17bit_b[4]), .B(in_17bit_b[3]), .CI(
        add_2_root_r119_carry_8_), .CO(add_2_root_r119_carry_9_), .S(
        add_2_root_r119_SUM_8_) );
  ADDFX2 U128 ( .A(in_17bit_b[9]), .B(in_17bit_b[7]), .CI(
        add_2_root_r115_carry_10_), .CO(add_2_root_r115_carry_11_), .S(
        add_2_root_r115_SUM_10_) );
  ADDFX2 U129 ( .A(add_1_root_r119_A_12_), .B(in_17bit_b[6]), .CI(
        add_1_root_r119_carry[12]), .CO(add_1_root_r119_carry[13]), .S(
        add_1_root_r119_SUM_12_) );
  ADDFX2 U130 ( .A(in_17bit_b[15]), .B(in_17bit_b[14]), .CI(
        add_3_root_r119_carry_16_), .CO(add_3_root_r119_carry_17_), .S(
        add_1_root_r119_A_16_) );
  ADDFX2 U131 ( .A(in_17bit_b[14]), .B(in_17bit_b[13]), .CI(
        add_2_root_r119_carry_18_), .CO(add_2_root_r119_carry_19_), .S(
        add_2_root_r119_SUM_18_) );
  ADDFX2 U132 ( .A(in_17bit_b[5]), .B(in_17bit_b[4]), .CI(
        add_2_root_r119_carry_9_), .CO(add_2_root_r119_carry_10_), .S(
        add_2_root_r119_SUM_9_) );
  ADDFX2 U133 ( .A(add_1_root_r119_A_11_), .B(in_17bit_b[5]), .CI(
        add_1_root_r119_carry[11]), .CO(add_1_root_r119_carry[12]), .S(
        add_1_root_r119_SUM_11_) );
  ADDFX2 U134 ( .A(add_1_root_r119_A_9_), .B(in_17bit_b[3]), .CI(
        add_1_root_r119_carry[9]), .CO(add_1_root_r119_carry[10]), .S(
        add_1_root_r119_SUM_9_) );
  ADDFX2 U135 ( .A(in_17bit_b[4]), .B(in_17bit_b[3]), .CI(
        add_3_root_r119_carry_5_), .CO(add_3_root_r119_carry_6_), .S(
        add_1_root_r119_A_5_) );
  ADDFX2 U136 ( .A(in_17bit_b[5]), .B(in_17bit_b[4]), .CI(
        add_3_root_r119_carry_6_), .CO(add_3_root_r119_carry_7_), .S(
        add_1_root_r119_A_6_) );
  ADDFX2 U137 ( .A(in_17bit_b[15]), .B(in_17bit_b[14]), .CI(
        add_2_root_r119_carry_19_), .CO(add_2_root_r119_carry_20_), .S(
        add_2_root_r119_SUM_19_) );
  BUFX3 U138 ( .A(in_17bit_b[16]), .Y(n42) );
  INVX1 U139 ( .A(n102), .Y(in_17bit_b[16]) );
  BUFX3 U140 ( .A(in_8bit[6]), .Y(n45) );
  BUFX3 U141 ( .A(in_8bit[1]), .Y(n44) );
  INVX1 U142 ( .A(in_8bit[2]), .Y(n43) );
  NOR3X1 U143 ( .A(n43), .B(n177), .C(n47), .Y(n157) );
  CLKINVX3 U144 ( .A(n155), .Y(in_17bit_b[0]) );
  INVX1 U145 ( .A(n103), .Y(n174) );
  OAI21XL U146 ( .A0(n103), .A1(n102), .B0(n104), .Y(N463) );
  AOI22X1 U147 ( .A0(N221), .A1(n41), .B0(N363), .B1(n40), .Y(n104) );
  NAND2XL U148 ( .A(N29), .B(n53), .Y(n102) );
  CLKINVX3 U149 ( .A(n110), .Y(in_17bit_b[15]) );
  AOI32X1 U150 ( .A0(n157), .A1(n175), .A2(in_8bit[5]), .B0(n158), .B1(n159), 
        .Y(n103) );
  INVX1 U151 ( .A(n160), .Y(n175) );
  INVXL U152 ( .A(in_8bit[3]), .Y(n177) );
  NAND3BXL U153 ( .AN(in_8bit[5]), .B(n43), .C(in_8bit[3]), .Y(n166) );
  NOR4BX1 U154 ( .AN(n165), .B(n47), .C(n44), .D(in_8bit[2]), .Y(n159) );
  NOR2XL U155 ( .A(n45), .B(in_8bit[3]), .Y(n165) );
  AOI22XL U156 ( .A0(in_17bit[0]), .A1(n48), .B0(in_17bit[0]), .B1(n55), .Y(
        n155) );
  AOI22X1 U157 ( .A0(N28), .A1(n51), .B0(in_17bit[15]), .B1(n54), .Y(n110) );
  AOI22X1 U158 ( .A0(N17), .A1(n51), .B0(in_17bit[4]), .B1(n54), .Y(n143) );
  AOI22X1 U159 ( .A0(N27), .A1(n51), .B0(in_17bit[14]), .B1(n55), .Y(n113) );
  AOI22X1 U160 ( .A0(N26), .A1(n51), .B0(in_17bit[13]), .B1(n54), .Y(n116) );
  AOI22XL U161 ( .A0(N14), .A1(n48), .B0(in_17bit[1]), .B1(n55), .Y(n152) );
  AOI22XL U162 ( .A0(N15), .A1(n48), .B0(in_17bit[2]), .B1(n55), .Y(n149) );
  AOI22X1 U163 ( .A0(N16), .A1(n51), .B0(in_17bit[3]), .B1(n55), .Y(n146) );
  AOI22X1 U164 ( .A0(N18), .A1(n51), .B0(in_17bit[5]), .B1(n54), .Y(n140) );
  AOI22X1 U165 ( .A0(N19), .A1(n51), .B0(in_17bit[6]), .B1(n54), .Y(n137) );
  AOI22X1 U166 ( .A0(N20), .A1(n51), .B0(in_17bit[7]), .B1(n54), .Y(n134) );
  AOI22X1 U167 ( .A0(N21), .A1(n51), .B0(in_17bit[8]), .B1(n55), .Y(n131) );
  AOI22X1 U168 ( .A0(N22), .A1(n51), .B0(in_17bit[9]), .B1(n54), .Y(n128) );
  AOI22X1 U169 ( .A0(N23), .A1(n51), .B0(in_17bit[10]), .B1(n55), .Y(n125) );
  AOI22X1 U170 ( .A0(N24), .A1(n51), .B0(in_17bit[11]), .B1(n55), .Y(n122) );
  AOI22X1 U171 ( .A0(N25), .A1(n51), .B0(in_17bit[12]), .B1(n54), .Y(n119) );
  NAND3X1 U172 ( .A(in_8bit[2]), .B(n177), .C(in_8bit[5]), .Y(n167) );
  AND2X2 U173 ( .A(n31), .B(n15), .Y(n23) );
  AND2X2 U174 ( .A(n23), .B(n6), .Y(n24) );
  AND2X2 U175 ( .A(n24), .B(n16), .Y(n25) );
  AND2X2 U176 ( .A(n27), .B(n3), .Y(n26) );
  AND2X2 U177 ( .A(n25), .B(n4), .Y(n27) );
  BUFX3 U178 ( .A(n106), .Y(n40) );
  OAI32X1 U179 ( .A0(n167), .A1(n46), .A2(n160), .B0(n166), .B1(n168), .Y(n106) );
  BUFX3 U180 ( .A(n105), .Y(n41) );
  OAI32X1 U181 ( .A0(n160), .A1(n46), .A2(n166), .B0(n167), .B1(n168), .Y(n105) );
  AND2X2 U182 ( .A(n26), .B(n5), .Y(n28) );
  INVX1 U183 ( .A(in_17bit[3]), .Y(n92) );
  INVX1 U184 ( .A(in_17bit[4]), .Y(n93) );
  INVX1 U185 ( .A(in_17bit[5]), .Y(n94) );
  INVX1 U186 ( .A(in_17bit[6]), .Y(n95) );
  INVX1 U187 ( .A(in_17bit[7]), .Y(n96) );
  INVX1 U188 ( .A(in_17bit[8]), .Y(n97) );
  INVX1 U189 ( .A(in_17bit[9]), .Y(n98) );
  INVX1 U190 ( .A(in_17bit[10]), .Y(n99) );
  INVX1 U191 ( .A(in_17bit[11]), .Y(n100) );
  INVX1 U192 ( .A(in_17bit[12]), .Y(n101) );
  INVX1 U193 ( .A(in_17bit[13]), .Y(n170) );
  INVX1 U194 ( .A(in_17bit[14]), .Y(n171) );
  INVX1 U195 ( .A(in_17bit[15]), .Y(n172) );
  INVX1 U196 ( .A(in_17bit[1]), .Y(n90) );
  INVX1 U197 ( .A(in_17bit[2]), .Y(n91) );
  INVX1 U198 ( .A(in_17bit[0]), .Y(n89) );
  NAND2X1 U199 ( .A(n153), .B(n154), .Y(N447) );
  AOI22X1 U200 ( .A0(N108), .A1(n109), .B0(N205), .B1(n41), .Y(n154) );
  AOI22X1 U201 ( .A0(N347), .A1(n40), .B0(n174), .B1(in_17bit_b[0]), .Y(n153)
         );
  NAND2X1 U202 ( .A(n150), .B(n151), .Y(N448) );
  AOI22X1 U203 ( .A0(N109), .A1(n109), .B0(N206), .B1(n41), .Y(n151) );
  AOI22X1 U204 ( .A0(N348), .A1(n40), .B0(n174), .B1(n173), .Y(n150) );
  INVX1 U205 ( .A(n152), .Y(n173) );
  NAND2X1 U206 ( .A(n147), .B(n148), .Y(N449) );
  AOI22X1 U207 ( .A0(N110), .A1(n109), .B0(N207), .B1(n41), .Y(n148) );
  AOI22X1 U208 ( .A0(N349), .A1(n40), .B0(n174), .B1(in_17bit_b[2]), .Y(n147)
         );
  NAND2X1 U209 ( .A(n144), .B(n145), .Y(N450) );
  AOI22X1 U210 ( .A0(N111), .A1(n109), .B0(N208), .B1(n41), .Y(n145) );
  AOI22X1 U211 ( .A0(N350), .A1(n40), .B0(n174), .B1(in_17bit_b[3]), .Y(n144)
         );
  NAND2X1 U212 ( .A(n141), .B(n142), .Y(N451) );
  AOI22X1 U213 ( .A0(N112), .A1(n109), .B0(N209), .B1(n41), .Y(n142) );
  AOI22X1 U214 ( .A0(N351), .A1(n40), .B0(n174), .B1(in_17bit_b[4]), .Y(n141)
         );
  NAND2X1 U215 ( .A(n138), .B(n139), .Y(N452) );
  AOI22X1 U216 ( .A0(N113), .A1(n109), .B0(N210), .B1(n41), .Y(n139) );
  AOI22X1 U217 ( .A0(N352), .A1(n40), .B0(n174), .B1(in_17bit_b[5]), .Y(n138)
         );
  NAND2X1 U218 ( .A(n135), .B(n136), .Y(N453) );
  AOI22X1 U219 ( .A0(N114), .A1(n109), .B0(N211), .B1(n41), .Y(n136) );
  AOI22X1 U220 ( .A0(N353), .A1(n40), .B0(n174), .B1(in_17bit_b[6]), .Y(n135)
         );
  NAND2X1 U221 ( .A(n132), .B(n133), .Y(N454) );
  AOI22X1 U222 ( .A0(N115), .A1(n109), .B0(N212), .B1(n41), .Y(n133) );
  AOI22X1 U223 ( .A0(N354), .A1(n40), .B0(n174), .B1(in_17bit_b[7]), .Y(n132)
         );
  NAND2X1 U224 ( .A(n129), .B(n130), .Y(N455) );
  AOI22X1 U225 ( .A0(N116), .A1(n109), .B0(N213), .B1(n41), .Y(n130) );
  AOI22X1 U226 ( .A0(N355), .A1(n40), .B0(n174), .B1(in_17bit_b[8]), .Y(n129)
         );
  NAND2X1 U227 ( .A(n126), .B(n127), .Y(N456) );
  AOI22X1 U228 ( .A0(N117), .A1(n109), .B0(N214), .B1(n41), .Y(n127) );
  AOI22X1 U229 ( .A0(N356), .A1(n40), .B0(n174), .B1(in_17bit_b[9]), .Y(n126)
         );
  NAND2X1 U230 ( .A(n123), .B(n124), .Y(N457) );
  AOI22X1 U231 ( .A0(N118), .A1(n109), .B0(N215), .B1(n41), .Y(n124) );
  AOI22X1 U232 ( .A0(N357), .A1(n40), .B0(n174), .B1(in_17bit_b[10]), .Y(n123)
         );
  NAND2X1 U233 ( .A(n120), .B(n121), .Y(N458) );
  AOI22X1 U234 ( .A0(N119), .A1(n109), .B0(N216), .B1(n41), .Y(n121) );
  AOI22X1 U235 ( .A0(N358), .A1(n40), .B0(n174), .B1(in_17bit_b[11]), .Y(n120)
         );
  NAND2X1 U236 ( .A(n117), .B(n118), .Y(N459) );
  AOI22X1 U237 ( .A0(N120), .A1(n109), .B0(N217), .B1(n41), .Y(n118) );
  AOI22X1 U238 ( .A0(N359), .A1(n40), .B0(n174), .B1(in_17bit_b[12]), .Y(n117)
         );
  NAND2X1 U239 ( .A(n114), .B(n115), .Y(N460) );
  AOI22X1 U240 ( .A0(N121), .A1(n109), .B0(N218), .B1(n41), .Y(n115) );
  AOI22X1 U241 ( .A0(N360), .A1(n40), .B0(n174), .B1(in_17bit_b[13]), .Y(n114)
         );
  NAND2X1 U242 ( .A(n111), .B(n112), .Y(N461) );
  AOI22X1 U243 ( .A0(N122), .A1(n109), .B0(N219), .B1(n41), .Y(n112) );
  AOI22X1 U244 ( .A0(N361), .A1(n40), .B0(n174), .B1(in_17bit_b[14]), .Y(n111)
         );
  NAND2X1 U245 ( .A(n107), .B(n108), .Y(N462) );
  AOI22X1 U246 ( .A0(N123), .A1(n109), .B0(N220), .B1(n41), .Y(n108) );
  AOI22X1 U247 ( .A0(N362), .A1(n40), .B0(n174), .B1(in_17bit_b[15]), .Y(n107)
         );
  INVX1 U248 ( .A(n71), .Y(n68) );
  OAI21XL U249 ( .A0(in_8bit[7]), .A1(n64), .B0(n63), .Y(n70) );
  XNOR2X1 U250 ( .A(n12), .B(sub_add_75_b0_carry[11]), .Y(n29) );
  AOI21X1 U251 ( .A0(n66), .A1(in_8bit[7]), .B0(n65), .Y(n67) );
  INVX1 U252 ( .A(n64), .Y(n66) );
  NOR2X1 U253 ( .A(in_8bit[7]), .B(neg_mul[9]), .Y(n65) );
  OAI21XL U254 ( .A0(in_8bit[7]), .A1(n73), .B0(n72), .Y(n78) );
  MX2X1 U255 ( .A(neg_mul[22]), .B(N480), .S0(n2), .Y(out[15]) );
  MX2X1 U256 ( .A(neg_mul[19]), .B(N477), .S0(n2), .Y(n197) );
  XNOR2X1 U257 ( .A(n38), .B(in_8bit[7]), .Y(n86) );
  MX2X1 U258 ( .A(neg_mul[23]), .B(N481), .S0(n2), .Y(out[16]) );
  NAND4BBX1 U259 ( .AN(n40), .BN(n41), .C(n156), .D(n103), .Y(N446) );
  AOI2BB1X1 U260 ( .A0N(n161), .A1N(n162), .B0(n109), .Y(n156) );
  OR4X2 U261 ( .A(in_8bit[4]), .B(in_8bit[5]), .C(n45), .D(in_8bit[7]), .Y(
        n161) );
  OR4XL U262 ( .A(n44), .B(n46), .C(in_8bit[2]), .D(in_8bit[3]), .Y(n162) );
  NOR3X1 U263 ( .A(in_8bit[4]), .B(in_8bit[5]), .C(n176), .Y(n158) );
  NAND4X1 U264 ( .A(n45), .B(in_8bit[4]), .C(n44), .D(n176), .Y(n160) );
  NOR2X1 U265 ( .A(n71), .B(neg_mul[10]), .Y(n31) );
  NAND4X1 U266 ( .A(n44), .B(in_8bit[7]), .C(n169), .D(n47), .Y(n168) );
  NOR2X1 U267 ( .A(n45), .B(in_8bit[4]), .Y(n169) );
  NOR2X1 U268 ( .A(out[0]), .B(neg_mul[8]), .Y(n32) );
  NAND2X1 U269 ( .A(n32), .B(n14), .Y(n71) );
  NAND2X1 U270 ( .A(out[0]), .B(neg_mul[8]), .Y(n57) );
  NAND2X1 U271 ( .A(neg_mul[10]), .B(n71), .Y(n73) );
  NAND2BX1 U272 ( .AN(n32), .B(neg_mul[9]), .Y(n64) );
  NAND2X1 U273 ( .A(n163), .B(n164), .Y(n109) );
  NAND4X1 U274 ( .A(n158), .B(n157), .C(n45), .D(n44), .Y(n164) );
  NAND4X1 U275 ( .A(n159), .B(in_8bit[5]), .C(in_8bit[4]), .D(n176), .Y(n163)
         );
  NOR2X1 U276 ( .A(n59), .B(n58), .Y(n60) );
  NOR2X1 U277 ( .A(in_8bit[7]), .B(neg_mul[8]), .Y(n58) );
  NOR2X1 U278 ( .A(n176), .B(n57), .Y(n59) );
  NOR2X1 U279 ( .A(n75), .B(n74), .Y(n76) );
  NOR2X1 U280 ( .A(in_8bit[7]), .B(neg_mul[10]), .Y(n74) );
  NOR2X1 U281 ( .A(n176), .B(n73), .Y(n75) );
  NAND2BX1 U282 ( .AN(neg_mul[10]), .B(in_8bit[7]), .Y(n72) );
  NAND2BX1 U283 ( .AN(neg_mul[9]), .B(in_8bit[7]), .Y(n63) );
  NAND2BX1 U284 ( .AN(neg_mul[8]), .B(in_8bit[7]), .Y(n56) );
  INVX1 U285 ( .A(in_8bit[7]), .Y(n176) );
  AOI211X2 U286 ( .A0(n38), .A1(n78), .B0(n77), .C0(n31), .Y(n198) );
  OAI21X4 U287 ( .A0(in_8bit[7]), .A1(n57), .B0(n56), .Y(n62) );
  NOR2X4 U288 ( .A(n38), .B(n60), .Y(n61) );
  XNOR2X4 U289 ( .A(n52), .B(in_8bit[7]), .Y(n79) );
  NOR2X4 U290 ( .A(n31), .B(n79), .Y(n80) );
  XNOR2X4 U291 ( .A(n82), .B(n6), .Y(out[5]) );
  XNOR2X4 U292 ( .A(n38), .B(in_8bit[7]), .Y(n83) );
  NOR2X4 U293 ( .A(n24), .B(n83), .Y(n84) );
  XNOR2X4 U294 ( .A(n87), .B(n7), .Y(out[10]) );
  MXI2X4 U295 ( .A(n12), .B(n29), .S0(n2), .Y(out[11]) );
  AND2X1 U296 ( .A(add_1_root_r112_carry_20_), .B(n42), .Y(
        add_1_root_r112_SUM_21_) );
  XOR2X1 U297 ( .A(n42), .B(add_1_root_r112_carry_20_), .Y(
        add_1_root_r112_SUM_20_) );
  AND2X1 U298 ( .A(add_1_root_r112_carry_19_), .B(in_17bit_b[15]), .Y(
        add_1_root_r112_carry_20_) );
  XOR2X1 U299 ( .A(in_17bit_b[15]), .B(add_1_root_r112_carry_19_), .Y(
        add_1_root_r112_SUM_19_) );
  AND2X1 U300 ( .A(add_1_root_r112_carry_18_), .B(in_17bit_b[14]), .Y(
        add_1_root_r112_carry_19_) );
  XOR2X1 U301 ( .A(in_17bit_b[14]), .B(add_1_root_r112_carry_18_), .Y(
        add_1_root_r112_SUM_18_) );
  AND2X1 U302 ( .A(add_1_root_r112_carry_17_), .B(in_17bit_b[13]), .Y(
        add_1_root_r112_carry_18_) );
  XOR2X1 U303 ( .A(in_17bit_b[13]), .B(add_1_root_r112_carry_17_), .Y(
        add_1_root_r112_SUM_17_) );
  AND2X1 U304 ( .A(add_2_root_r119_carry_21_), .B(n42), .Y(
        add_2_root_r119_SUM_22_) );
  XOR2X1 U305 ( .A(n42), .B(add_2_root_r119_carry_21_), .Y(
        add_2_root_r119_SUM_21_) );
  AND2X1 U306 ( .A(in_17bit_b[1]), .B(in_17bit_b[0]), .Y(
        add_2_root_r119_carry_6_) );
  XOR2X1 U307 ( .A(in_17bit_b[0]), .B(in_17bit_b[1]), .Y(
        add_2_root_r119_SUM_5_) );
  AND2X1 U308 ( .A(add_1_root_r119_carry[22]), .B(n42), .Y(
        add_1_root_r119_SUM_23_) );
  XOR2X1 U309 ( .A(n42), .B(add_1_root_r119_carry[22]), .Y(
        add_1_root_r119_SUM_22_) );
  AND2X1 U310 ( .A(add_1_root_r119_carry[21]), .B(in_17bit_b[15]), .Y(
        add_1_root_r119_carry[22]) );
  XOR2X1 U311 ( .A(in_17bit_b[15]), .B(add_1_root_r119_carry[21]), .Y(
        add_1_root_r119_SUM_21_) );
  AND2X1 U312 ( .A(add_1_root_r119_carry[20]), .B(in_17bit_b[14]), .Y(
        add_1_root_r119_carry[21]) );
  XOR2X1 U313 ( .A(in_17bit_b[14]), .B(add_1_root_r119_carry[20]), .Y(
        add_1_root_r119_SUM_20_) );
  AND2X1 U314 ( .A(add_1_root_r119_A_6_), .B(in_17bit_b[0]), .Y(
        add_1_root_r119_carry[7]) );
  XOR2X1 U315 ( .A(in_17bit_b[0]), .B(add_1_root_r119_A_6_), .Y(
        add_1_root_r119_SUM_6_) );
  AND2X1 U316 ( .A(add_3_root_r119_carry_18_), .B(n42), .Y(
        add_1_root_r119_A_19_) );
  XOR2X1 U317 ( .A(n42), .B(add_3_root_r119_carry_18_), .Y(
        add_1_root_r119_A_18_) );
  AND2X1 U318 ( .A(in_17bit_b[1]), .B(in_17bit_b[0]), .Y(
        add_3_root_r119_carry_3_) );
  XOR2X1 U319 ( .A(in_17bit_b[0]), .B(in_17bit_b[1]), .Y(add_1_root_r119_A_2_)
         );
  AND2X1 U320 ( .A(add_2_root_r115_carry_19_), .B(n42), .Y(
        add_2_root_r115_SUM_20_) );
  XOR2X1 U321 ( .A(n42), .B(add_2_root_r115_carry_19_), .Y(
        add_2_root_r115_SUM_19_) );
  AND2X1 U322 ( .A(add_2_root_r115_carry_18_), .B(in_17bit_b[15]), .Y(
        add_2_root_r115_carry_19_) );
  XOR2X1 U323 ( .A(in_17bit_b[15]), .B(add_2_root_r115_carry_18_), .Y(
        add_2_root_r115_SUM_18_) );
  AND2X1 U324 ( .A(in_17bit_b[2]), .B(in_17bit_b[0]), .Y(
        add_2_root_r115_carry_4_) );
  XOR2X1 U325 ( .A(in_17bit_b[0]), .B(in_17bit_b[2]), .Y(
        add_2_root_r115_SUM_3_) );
  AND2X1 U326 ( .A(add_1_root_r115_carry_22_), .B(n42), .Y(
        add_1_root_r115_SUM_23_) );
  XOR2X1 U327 ( .A(n42), .B(add_1_root_r115_carry_22_), .Y(
        add_1_root_r115_SUM_22_) );
  AND2X1 U328 ( .A(add_1_root_r115_carry_21_), .B(in_17bit_b[15]), .Y(
        add_1_root_r115_carry_22_) );
  XOR2X1 U329 ( .A(in_17bit_b[15]), .B(add_1_root_r115_carry_21_), .Y(
        add_1_root_r115_SUM_21_) );
  AND2X1 U330 ( .A(in_17bit_b[2]), .B(in_17bit_b[0]), .Y(
        add_1_root_r115_carry_7_) );
  XOR2X1 U331 ( .A(in_17bit_b[0]), .B(in_17bit_b[2]), .Y(
        add_1_root_r115_SUM_6_) );
  XOR2X1 U332 ( .A(n55), .B(sub_add_54_b0_carry[16]), .Y(N29) );
  AND2X1 U333 ( .A(sub_add_54_b0_carry[15]), .B(n172), .Y(
        sub_add_54_b0_carry[16]) );
  XOR2X1 U334 ( .A(n172), .B(sub_add_54_b0_carry[15]), .Y(N28) );
  AND2X1 U335 ( .A(sub_add_54_b0_carry[14]), .B(n171), .Y(
        sub_add_54_b0_carry[15]) );
  XOR2X1 U336 ( .A(n171), .B(sub_add_54_b0_carry[14]), .Y(N27) );
  AND2X1 U337 ( .A(sub_add_54_b0_carry[13]), .B(n170), .Y(
        sub_add_54_b0_carry[14]) );
  XOR2X1 U338 ( .A(n170), .B(sub_add_54_b0_carry[13]), .Y(N26) );
  AND2X1 U339 ( .A(sub_add_54_b0_carry[12]), .B(n101), .Y(
        sub_add_54_b0_carry[13]) );
  XOR2X1 U340 ( .A(n101), .B(sub_add_54_b0_carry[12]), .Y(N25) );
  AND2X1 U341 ( .A(sub_add_54_b0_carry[11]), .B(n100), .Y(
        sub_add_54_b0_carry[12]) );
  XOR2X1 U342 ( .A(n100), .B(sub_add_54_b0_carry[11]), .Y(N24) );
  AND2X1 U343 ( .A(sub_add_54_b0_carry[10]), .B(n99), .Y(
        sub_add_54_b0_carry[11]) );
  XOR2X1 U344 ( .A(n99), .B(sub_add_54_b0_carry[10]), .Y(N23) );
  AND2X1 U345 ( .A(sub_add_54_b0_carry[9]), .B(n98), .Y(
        sub_add_54_b0_carry[10]) );
  XOR2X1 U346 ( .A(n98), .B(sub_add_54_b0_carry[9]), .Y(N22) );
  AND2X1 U347 ( .A(sub_add_54_b0_carry[8]), .B(n97), .Y(sub_add_54_b0_carry[9]) );
  XOR2X1 U348 ( .A(n97), .B(sub_add_54_b0_carry[8]), .Y(N21) );
  AND2X1 U349 ( .A(sub_add_54_b0_carry[7]), .B(n96), .Y(sub_add_54_b0_carry[8]) );
  XOR2X1 U350 ( .A(n96), .B(sub_add_54_b0_carry[7]), .Y(N20) );
  AND2X1 U351 ( .A(sub_add_54_b0_carry[6]), .B(n95), .Y(sub_add_54_b0_carry[7]) );
  XOR2X1 U352 ( .A(n95), .B(sub_add_54_b0_carry[6]), .Y(N19) );
  AND2X1 U353 ( .A(sub_add_54_b0_carry[5]), .B(n94), .Y(sub_add_54_b0_carry[6]) );
  XOR2X1 U354 ( .A(n94), .B(sub_add_54_b0_carry[5]), .Y(N18) );
  AND2X1 U355 ( .A(sub_add_54_b0_carry[4]), .B(n93), .Y(sub_add_54_b0_carry[5]) );
  XOR2X1 U356 ( .A(n93), .B(sub_add_54_b0_carry[4]), .Y(N17) );
  AND2X1 U357 ( .A(sub_add_54_b0_carry[3]), .B(n92), .Y(sub_add_54_b0_carry[4]) );
  XOR2X1 U358 ( .A(n92), .B(sub_add_54_b0_carry[3]), .Y(N16) );
  AND2X1 U359 ( .A(sub_add_54_b0_carry[2]), .B(n91), .Y(sub_add_54_b0_carry[3]) );
  XOR2X1 U360 ( .A(n91), .B(sub_add_54_b0_carry[2]), .Y(N15) );
  AND2X1 U361 ( .A(n89), .B(n90), .Y(sub_add_54_b0_carry[2]) );
  XOR2X1 U362 ( .A(n90), .B(n89), .Y(N14) );
  XOR2X1 U363 ( .A(n13), .B(sub_add_75_b0_carry[16]), .Y(N481) );
  AND2X1 U364 ( .A(sub_add_75_b0_carry[15]), .B(n10), .Y(
        sub_add_75_b0_carry[16]) );
  XOR2X1 U365 ( .A(n10), .B(sub_add_75_b0_carry[15]), .Y(N480) );
  AND2X1 U366 ( .A(sub_add_75_b0_carry[14]), .B(n8), .Y(
        sub_add_75_b0_carry[15]) );
  XOR2X1 U367 ( .A(n8), .B(sub_add_75_b0_carry[14]), .Y(N479) );
  AND2X1 U368 ( .A(sub_add_75_b0_carry[13]), .B(n9), .Y(
        sub_add_75_b0_carry[14]) );
  XOR2X1 U369 ( .A(n9), .B(sub_add_75_b0_carry[13]), .Y(N478) );
  AND2X1 U370 ( .A(sub_add_75_b0_carry[12]), .B(n11), .Y(
        sub_add_75_b0_carry[13]) );
  XOR2X1 U371 ( .A(n11), .B(sub_add_75_b0_carry[12]), .Y(N477) );
  AND2X1 U372 ( .A(sub_add_75_b0_carry[11]), .B(n12), .Y(
        sub_add_75_b0_carry[12]) );
  AND2X1 U373 ( .A(n28), .B(n7), .Y(sub_add_75_b0_carry[11]) );
  AND2X1 U374 ( .A(in_17bit_b[0]), .B(in_17bit_b[4]), .Y(
        add_1_root_r112_carry_5_) );
endmodule


module multi16_11_DW01_add_0 ( A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, 
        A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, 
        A_4_, B_23_, B_22_, B_21_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, 
        B_14_, B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, 
        SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, 
        SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, 
        SUM_7_ );
  input A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_,
         A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, B_23_, B_22_,
         B_21_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_,
         B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_;
  output SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_,
         SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_,
         SUM_8_, SUM_7_;
  wire   n1, n2, n3, n4;
  wire   [23:7] carry;

  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry[7]), .CO(carry[8]), .S(SUM_7_)
         );
  ADDFX2 U1_21 ( .A(A_21_), .B(B_21_), .CI(carry[21]), .CO(carry[22]), .S(
        SUM_21_) );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry[20]), .CO(carry[21]), .S(
        SUM_20_) );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry[19]), .CO(carry[20]), .S(
        SUM_19_) );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry[18]), .CO(carry[19]), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry[17]), .CO(carry[18]), .S(
        SUM_17_) );
  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry[16]), .CO(carry[17]), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry[15]), .CO(carry[16]), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry[14]), .CO(carry[15]), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry[13]), .CO(carry[14]), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry[12]), .CO(carry[13]), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry[11]), .CO(carry[12]), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry[10]), .CO(carry[11]), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry[9]), .CO(carry[10]), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry[8]), .CO(carry[9]), .S(SUM_8_)
         );
  ADDFX2 U1_22 ( .A(A_22_), .B(B_22_), .CI(carry[22]), .CO(carry[23]), .S(
        SUM_22_) );
  AND2X2 U1 ( .A(A_4_), .B(B_4_), .Y(n1) );
  XOR2X1 U2 ( .A(B_23_), .B(carry[23]), .Y(SUM_23_) );
  OAI2BB1X1 U3 ( .A0N(n2), .A1N(A_6_), .B0(n3), .Y(carry[7]) );
  OAI21XL U4 ( .A0(A_6_), .A1(n2), .B0(B_6_), .Y(n3) );
  OAI2BB1X1 U5 ( .A0N(n1), .A1N(A_5_), .B0(n4), .Y(n2) );
  OAI21XL U6 ( .A0(A_5_), .A1(n1), .B0(B_5_), .Y(n4) );
endmodule


module multi16_11_DW01_add_4 ( A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, 
        A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, 
        B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, 
        B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, SUM_22_, SUM_21_, SUM_20_, 
        SUM_19_, SUM_18_, SUM_17_, SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, 
        SUM_11_, SUM_10_, SUM_9_, SUM_8_, SUM_7_ );
  input A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_,
         A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, B_20_, B_19_,
         B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, B_10_, B_9_,
         B_8_, B_7_, B_6_, B_5_;
  output SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_,
         SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_,
         SUM_7_;
  wire   carry_21_, carry_20_, carry_19_, carry_18_, carry_17_, carry_16_,
         carry_15_, carry_14_, carry_13_, carry_12_, carry_11_, carry_10_,
         carry_9_, carry_8_, carry_7_, n1;

  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry_16_), .CO(carry_17_), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry_15_), .CO(carry_16_), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry_14_), .CO(carry_15_), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry_13_), .CO(carry_14_), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry_12_), .CO(carry_13_), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry_11_), .CO(carry_12_), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry_10_), .CO(carry_11_), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry_9_), .CO(carry_10_), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry_8_), .CO(carry_9_), .S(SUM_8_)
         );
  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry_7_), .CO(carry_8_), .S(SUM_7_)
         );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry_20_), .CO(carry_21_), .S(
        SUM_20_) );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry_19_), .CO(carry_20_), .S(
        SUM_19_) );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry_18_), .CO(carry_19_), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry_17_), .CO(carry_18_), .S(
        SUM_17_) );
  ADDFX2 U1_21 ( .A(A_21_), .B(B_21_), .CI(carry_21_), .CO(SUM_22_), .S(
        SUM_21_) );
  OAI2BB1X1 U1 ( .A0N(A_6_), .A1N(B_6_), .B0(n1), .Y(carry_7_) );
  OAI211X1 U2 ( .A0(B_6_), .A1(A_6_), .B0(A_5_), .C0(B_5_), .Y(n1) );
endmodule


module multi16_11_DW01_add_6 ( A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, 
        A_16_, A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, 
        A_6_, A_5_, A_4_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, 
        B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, 
        SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, 
        SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, 
        SUM_7_ );
  input A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_,
         A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, B_20_,
         B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, B_10_,
         B_9_, B_8_, B_7_, B_6_, B_5_, B_4_;
  output SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_,
         SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_,
         SUM_8_, SUM_7_;
  wire   n1, n2, n3, n4, n5, n6;
  wire   [21:7] carry;

  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry[7]), .CO(carry[8]), .S(SUM_7_)
         );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry[18]), .CO(carry[19]), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry[17]), .CO(carry[18]), .S(
        SUM_17_) );
  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry[16]), .CO(carry[17]), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry[15]), .CO(carry[16]), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry[14]), .CO(carry[15]), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry[13]), .CO(carry[14]), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry[12]), .CO(carry[13]), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry[11]), .CO(carry[12]), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry[10]), .CO(carry[11]), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry[9]), .CO(carry[10]), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry[8]), .CO(carry[9]), .S(SUM_8_)
         );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry[19]), .CO(carry[20]), .S(
        SUM_19_) );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry[20]), .CO(carry[21]), .S(
        SUM_20_) );
  AND2X2 U1 ( .A(A_22_), .B(n2), .Y(n1) );
  AND2X2 U2 ( .A(A_21_), .B(carry[21]), .Y(n2) );
  AND2X2 U3 ( .A(A_4_), .B(B_4_), .Y(n3) );
  XOR2X1 U4 ( .A(A_23_), .B(n1), .Y(SUM_23_) );
  XOR2X1 U5 ( .A(A_21_), .B(carry[21]), .Y(SUM_21_) );
  XOR2X1 U6 ( .A(A_22_), .B(n2), .Y(SUM_22_) );
  OAI2BB1X1 U7 ( .A0N(n4), .A1N(A_6_), .B0(n5), .Y(carry[7]) );
  OAI21XL U8 ( .A0(A_6_), .A1(n4), .B0(B_6_), .Y(n5) );
  OAI2BB1X1 U9 ( .A0N(n3), .A1N(A_5_), .B0(n6), .Y(n4) );
  OAI21XL U10 ( .A0(A_5_), .A1(n3), .B0(B_5_), .Y(n6) );
endmodule


module multi16_11 ( in_17bit, in_8bit, out );
  input [16:0] in_17bit;
  input [7:0] in_8bit;
  output [16:0] out;
  wire   n252, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26,
         N27, N28, N29, N108, N109, N110, N111, N112, N113, N114, N115, N116,
         N117, N118, N119, N120, N121, N122, N123, N205, N206, N207, N208,
         N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, N219,
         N220, N221, N347, N348, N349, N350, N351, N352, N353, N354, N355,
         N356, N357, N358, N359, N360, N361, N362, N363, N446, N447, N448,
         N449, N450, N451, N452, N453, N454, N455, N456, N457, N458, N459,
         N460, N461, N462, N463, N476, N477, N478, N479, N480,
         add_2_root_r119_carry_10_, add_2_root_r119_carry_11_,
         add_2_root_r119_carry_12_, add_2_root_r119_carry_13_,
         add_2_root_r119_carry_14_, add_2_root_r119_carry_15_,
         add_2_root_r119_carry_16_, add_2_root_r119_carry_17_,
         add_2_root_r119_carry_18_, add_2_root_r119_carry_19_,
         add_2_root_r119_carry_20_, add_2_root_r119_carry_21_,
         add_2_root_r119_carry_6_, add_2_root_r119_carry_7_,
         add_2_root_r119_carry_8_, add_2_root_r119_carry_9_,
         add_2_root_r119_SUM_5_, add_2_root_r119_SUM_6_,
         add_2_root_r119_SUM_7_, add_2_root_r119_SUM_8_,
         add_2_root_r119_SUM_9_, add_2_root_r119_SUM_10_,
         add_2_root_r119_SUM_11_, add_2_root_r119_SUM_12_,
         add_2_root_r119_SUM_13_, add_2_root_r119_SUM_14_,
         add_2_root_r119_SUM_15_, add_2_root_r119_SUM_16_,
         add_2_root_r119_SUM_17_, add_2_root_r119_SUM_18_,
         add_2_root_r119_SUM_19_, add_2_root_r119_SUM_20_,
         add_2_root_r119_SUM_21_, add_2_root_r119_SUM_22_,
         add_1_root_r119_SUM_6_, add_1_root_r119_SUM_7_,
         add_1_root_r119_SUM_8_, add_1_root_r119_SUM_9_,
         add_1_root_r119_SUM_10_, add_1_root_r119_SUM_11_,
         add_1_root_r119_SUM_12_, add_1_root_r119_SUM_13_,
         add_1_root_r119_SUM_14_, add_1_root_r119_SUM_15_,
         add_1_root_r119_SUM_16_, add_1_root_r119_SUM_17_,
         add_1_root_r119_SUM_18_, add_1_root_r119_SUM_19_,
         add_1_root_r119_SUM_20_, add_1_root_r119_SUM_21_,
         add_1_root_r119_SUM_22_, add_1_root_r119_SUM_23_,
         add_1_root_r119_A_2_, add_1_root_r119_A_3_, add_1_root_r119_A_4_,
         add_1_root_r119_A_5_, add_1_root_r119_A_6_, add_1_root_r119_A_7_,
         add_1_root_r119_A_8_, add_1_root_r119_A_9_, add_1_root_r119_A_10_,
         add_1_root_r119_A_11_, add_1_root_r119_A_12_, add_1_root_r119_A_13_,
         add_1_root_r119_A_14_, add_1_root_r119_A_15_, add_1_root_r119_A_16_,
         add_1_root_r119_A_17_, add_1_root_r119_A_18_, add_1_root_r119_A_19_,
         add_3_root_r119_carry_10_, add_3_root_r119_carry_11_,
         add_3_root_r119_carry_12_, add_3_root_r119_carry_13_,
         add_3_root_r119_carry_14_, add_3_root_r119_carry_15_,
         add_3_root_r119_carry_16_, add_3_root_r119_carry_17_,
         add_3_root_r119_carry_18_, add_3_root_r119_carry_3_,
         add_3_root_r119_carry_4_, add_3_root_r119_carry_5_,
         add_3_root_r119_carry_6_, add_3_root_r119_carry_7_,
         add_3_root_r119_carry_8_, add_3_root_r119_carry_9_,
         add_1_root_r112_carry_10_, add_1_root_r112_carry_11_,
         add_1_root_r112_carry_12_, add_1_root_r112_carry_13_,
         add_1_root_r112_carry_14_, add_1_root_r112_carry_15_,
         add_1_root_r112_carry_16_, add_1_root_r112_carry_17_,
         add_1_root_r112_carry_18_, add_1_root_r112_carry_19_,
         add_1_root_r112_carry_20_, add_1_root_r112_carry_5_,
         add_1_root_r112_carry_6_, add_1_root_r112_carry_7_,
         add_1_root_r112_carry_8_, add_1_root_r112_carry_9_,
         add_1_root_r112_SUM_1_, add_1_root_r112_SUM_2_,
         add_1_root_r112_SUM_3_, add_1_root_r112_SUM_4_,
         add_1_root_r112_SUM_5_, add_1_root_r112_SUM_6_,
         add_1_root_r112_SUM_7_, add_1_root_r112_SUM_8_,
         add_1_root_r112_SUM_9_, add_1_root_r112_SUM_10_,
         add_1_root_r112_SUM_11_, add_1_root_r112_SUM_12_,
         add_1_root_r112_SUM_13_, add_1_root_r112_SUM_14_,
         add_1_root_r112_SUM_15_, add_1_root_r112_SUM_16_,
         add_1_root_r112_SUM_17_, add_1_root_r112_SUM_18_,
         add_1_root_r112_SUM_19_, add_1_root_r112_SUM_20_,
         add_1_root_r112_SUM_21_, add_2_root_r115_carry_10_,
         add_2_root_r115_carry_11_, add_2_root_r115_carry_12_,
         add_2_root_r115_carry_13_, add_2_root_r115_carry_14_,
         add_2_root_r115_carry_15_, add_2_root_r115_carry_16_,
         add_2_root_r115_carry_17_, add_2_root_r115_carry_18_,
         add_2_root_r115_carry_19_, add_2_root_r115_carry_4_,
         add_2_root_r115_carry_5_, add_2_root_r115_carry_6_,
         add_2_root_r115_carry_7_, add_2_root_r115_carry_8_,
         add_2_root_r115_carry_9_, add_2_root_r115_SUM_3_,
         add_2_root_r115_SUM_4_, add_2_root_r115_SUM_5_,
         add_2_root_r115_SUM_6_, add_2_root_r115_SUM_7_,
         add_2_root_r115_SUM_8_, add_2_root_r115_SUM_9_,
         add_2_root_r115_SUM_10_, add_2_root_r115_SUM_11_,
         add_2_root_r115_SUM_12_, add_2_root_r115_SUM_13_,
         add_2_root_r115_SUM_14_, add_2_root_r115_SUM_15_,
         add_2_root_r115_SUM_16_, add_2_root_r115_SUM_17_,
         add_2_root_r115_SUM_18_, add_2_root_r115_SUM_19_,
         add_2_root_r115_SUM_20_, add_1_root_r115_carry_10_,
         add_1_root_r115_carry_11_, add_1_root_r115_carry_12_,
         add_1_root_r115_carry_13_, add_1_root_r115_carry_14_,
         add_1_root_r115_carry_15_, add_1_root_r115_carry_16_,
         add_1_root_r115_carry_17_, add_1_root_r115_carry_18_,
         add_1_root_r115_carry_19_, add_1_root_r115_carry_20_,
         add_1_root_r115_carry_21_, add_1_root_r115_carry_22_,
         add_1_root_r115_carry_7_, add_1_root_r115_carry_8_,
         add_1_root_r115_carry_9_, add_1_root_r115_SUM_6_,
         add_1_root_r115_SUM_7_, add_1_root_r115_SUM_8_,
         add_1_root_r115_SUM_9_, add_1_root_r115_SUM_10_,
         add_1_root_r115_SUM_11_, add_1_root_r115_SUM_12_,
         add_1_root_r115_SUM_13_, add_1_root_r115_SUM_14_,
         add_1_root_r115_SUM_15_, add_1_root_r115_SUM_16_,
         add_1_root_r115_SUM_17_, add_1_root_r115_SUM_18_,
         add_1_root_r115_SUM_19_, add_1_root_r115_SUM_20_,
         add_1_root_r115_SUM_21_, add_1_root_r115_SUM_22_,
         add_1_root_r115_SUM_23_, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n158, n160, n161, n162, n163, n164, n168, n170,
         n171, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251;
  wire   [16:0] in_17bit_b;
  wire   [23:8] neg_mul;
  wire   [15:10] sub_add_75_b0_carry;
  wire   [16:2] sub_add_54_b0_carry;
  wire   [22:7] add_1_root_r119_carry;

  multi16_11_DW01_add_0 add_0_root_r119 ( .A_22_(add_2_root_r119_SUM_22_), 
        .A_21_(add_2_root_r119_SUM_21_), .A_20_(add_2_root_r119_SUM_20_), 
        .A_19_(add_2_root_r119_SUM_19_), .A_18_(add_2_root_r119_SUM_18_), 
        .A_17_(add_2_root_r119_SUM_17_), .A_16_(add_2_root_r119_SUM_16_), 
        .A_15_(add_2_root_r119_SUM_15_), .A_14_(add_2_root_r119_SUM_14_), 
        .A_13_(add_2_root_r119_SUM_13_), .A_12_(add_2_root_r119_SUM_12_), 
        .A_11_(add_2_root_r119_SUM_11_), .A_10_(add_2_root_r119_SUM_10_), 
        .A_9_(add_2_root_r119_SUM_9_), .A_8_(add_2_root_r119_SUM_8_), .A_7_(
        add_2_root_r119_SUM_7_), .A_6_(add_2_root_r119_SUM_6_), .A_5_(
        add_2_root_r119_SUM_5_), .A_4_(in_17bit_b[0]), .B_23_(
        add_1_root_r119_SUM_23_), .B_22_(add_1_root_r119_SUM_22_), .B_21_(
        add_1_root_r119_SUM_21_), .B_20_(add_1_root_r119_SUM_20_), .B_19_(
        add_1_root_r119_SUM_19_), .B_18_(add_1_root_r119_SUM_18_), .B_17_(
        add_1_root_r119_SUM_17_), .B_16_(add_1_root_r119_SUM_16_), .B_15_(
        add_1_root_r119_SUM_15_), .B_14_(add_1_root_r119_SUM_14_), .B_13_(
        add_1_root_r119_SUM_13_), .B_12_(add_1_root_r119_SUM_12_), .B_11_(
        add_1_root_r119_SUM_11_), .B_10_(add_1_root_r119_SUM_10_), .B_9_(
        add_1_root_r119_SUM_9_), .B_8_(add_1_root_r119_SUM_8_), .B_7_(
        add_1_root_r119_SUM_7_), .B_6_(add_1_root_r119_SUM_6_), .B_5_(
        add_1_root_r119_A_5_), .B_4_(add_1_root_r119_A_4_), .SUM_23_(N363), 
        .SUM_22_(N362), .SUM_21_(N361), .SUM_20_(N360), .SUM_19_(N359), 
        .SUM_18_(N358), .SUM_17_(N357), .SUM_16_(N356), .SUM_15_(N355), 
        .SUM_14_(N354), .SUM_13_(N353), .SUM_12_(N352), .SUM_11_(N351), 
        .SUM_10_(N350), .SUM_9_(N349), .SUM_8_(N348), .SUM_7_(N347) );
  multi16_11_DW01_add_4 add_0_root_r112 ( .A_21_(n40), .A_20_(in_17bit_b[15]), 
        .A_19_(in_17bit_b[14]), .A_18_(in_17bit_b[13]), .A_17_(in_17bit_b[12]), 
        .A_16_(in_17bit_b[11]), .A_15_(in_17bit_b[10]), .A_14_(in_17bit_b[9]), 
        .A_13_(in_17bit_b[8]), .A_12_(in_17bit_b[7]), .A_11_(in_17bit_b[6]), 
        .A_10_(in_17bit_b[5]), .A_9_(in_17bit_b[4]), .A_8_(in_17bit_b[3]), 
        .A_7_(in_17bit_b[2]), .A_6_(in_17bit_b[1]), .A_5_(in_17bit_b[0]), 
        .B_21_(add_1_root_r112_SUM_21_), .B_20_(add_1_root_r112_SUM_20_), 
        .B_19_(add_1_root_r112_SUM_19_), .B_18_(add_1_root_r112_SUM_18_), 
        .B_17_(add_1_root_r112_SUM_17_), .B_16_(add_1_root_r112_SUM_16_), 
        .B_15_(add_1_root_r112_SUM_15_), .B_14_(add_1_root_r112_SUM_14_), 
        .B_13_(add_1_root_r112_SUM_13_), .B_12_(add_1_root_r112_SUM_12_), 
        .B_11_(add_1_root_r112_SUM_11_), .B_10_(add_1_root_r112_SUM_10_), 
        .B_9_(add_1_root_r112_SUM_9_), .B_8_(add_1_root_r112_SUM_8_), .B_7_(
        add_1_root_r112_SUM_7_), .B_6_(add_1_root_r112_SUM_6_), .B_5_(
        add_1_root_r112_SUM_5_), .SUM_22_(N123), .SUM_21_(N122), .SUM_20_(N121), .SUM_19_(N120), .SUM_18_(N119), .SUM_17_(N118), .SUM_16_(N117), .SUM_15_(
        N116), .SUM_14_(N115), .SUM_13_(N114), .SUM_12_(N113), .SUM_11_(N112), 
        .SUM_10_(N111), .SUM_9_(N110), .SUM_8_(N109), .SUM_7_(N108) );
  multi16_11_DW01_add_6 add_0_root_r115 ( .A_23_(add_1_root_r115_SUM_23_), 
        .A_22_(add_1_root_r115_SUM_22_), .A_21_(add_1_root_r115_SUM_21_), 
        .A_20_(add_1_root_r115_SUM_20_), .A_19_(add_1_root_r115_SUM_19_), 
        .A_18_(add_1_root_r115_SUM_18_), .A_17_(add_1_root_r115_SUM_17_), 
        .A_16_(add_1_root_r115_SUM_16_), .A_15_(add_1_root_r115_SUM_15_), 
        .A_14_(add_1_root_r115_SUM_14_), .A_13_(add_1_root_r115_SUM_13_), 
        .A_12_(add_1_root_r115_SUM_12_), .A_11_(add_1_root_r115_SUM_11_), 
        .A_10_(add_1_root_r115_SUM_10_), .A_9_(add_1_root_r115_SUM_9_), .A_8_(
        add_1_root_r115_SUM_8_), .A_7_(add_1_root_r115_SUM_7_), .A_6_(
        add_1_root_r115_SUM_6_), .A_5_(in_17bit_b[1]), .A_4_(in_17bit_b[0]), 
        .B_20_(add_2_root_r115_SUM_20_), .B_19_(add_2_root_r115_SUM_19_), 
        .B_18_(add_2_root_r115_SUM_18_), .B_17_(add_2_root_r115_SUM_17_), 
        .B_16_(add_2_root_r115_SUM_16_), .B_15_(add_2_root_r115_SUM_15_), 
        .B_14_(add_2_root_r115_SUM_14_), .B_13_(add_2_root_r115_SUM_13_), 
        .B_12_(add_2_root_r115_SUM_12_), .B_11_(add_2_root_r115_SUM_11_), 
        .B_10_(add_2_root_r115_SUM_10_), .B_9_(add_2_root_r115_SUM_9_), .B_8_(
        add_2_root_r115_SUM_8_), .B_7_(add_2_root_r115_SUM_7_), .B_6_(
        add_2_root_r115_SUM_6_), .B_5_(add_2_root_r115_SUM_5_), .B_4_(
        add_2_root_r115_SUM_4_), .SUM_23_(N221), .SUM_22_(N220), .SUM_21_(N219), .SUM_20_(N218), .SUM_19_(N217), .SUM_18_(N216), .SUM_17_(N215), .SUM_16_(
        N214), .SUM_15_(N213), .SUM_14_(N212), .SUM_13_(N211), .SUM_12_(N210), 
        .SUM_11_(N209), .SUM_10_(N208), .SUM_9_(N207), .SUM_8_(N206), .SUM_7_(
        N205) );
  TLATX1 neg_mul_reg_16_ ( .G(N446), .D(N456), .QN(n7) );
  TLATX1 neg_mul_reg_15_ ( .G(N446), .D(N455), .QN(n3) );
  TLATX1 neg_mul_reg_14_ ( .G(N446), .D(N454), .QN(n6) );
  TLATX1 neg_mul_reg_13_ ( .G(N446), .D(N453), .Q(neg_mul[13]), .QN(n1) );
  TLATX1 neg_mul_reg_12_ ( .G(N446), .D(N452), .QN(n5) );
  TLATX1 neg_mul_reg_11_ ( .G(N446), .D(N451), .QN(n4) );
  TLATX1 neg_mul_reg_23_ ( .G(N446), .D(N463), .Q(neg_mul[23]), .QN(n2) );
  TLATX1 neg_mul_reg_22_ ( .G(N446), .D(N462), .Q(neg_mul[22]), .QN(n9) );
  TLATX1 neg_mul_reg_21_ ( .G(N446), .D(N461), .Q(neg_mul[21]), .QN(n10) );
  TLATX1 neg_mul_reg_20_ ( .G(N446), .D(N460), .Q(neg_mul[20]), .QN(n11) );
  TLATX1 neg_mul_reg_19_ ( .G(N446), .D(N459), .Q(neg_mul[19]), .QN(n12) );
  TLATX1 neg_mul_reg_18_ ( .G(N446), .D(N458), .Q(neg_mul[18]), .QN(n13) );
  TLATX1 neg_mul_reg_17_ ( .G(N446), .D(N457), .QN(n14) );
  TLATX1 neg_mul_reg_9_ ( .G(N446), .D(N449), .Q(neg_mul[9]), .QN(n15) );
  TLATX1 neg_mul_reg_10_ ( .G(N446), .D(N450), .Q(neg_mul[10]), .QN(n8) );
  TLATX1 neg_mul_reg_8_ ( .G(N446), .D(N448), .Q(neg_mul[8]), .QN(n16) );
  TLATX1 neg_mul_reg_7_ ( .G(N446), .D(N447), .Q(out[0]) );
  NAND2X1 U2 ( .A(n36), .B(n16), .Y(n54) );
  AOI211X2 U3 ( .A0(n37), .A1(n59), .B0(n58), .C0(n33), .Y(out[1]) );
  NOR2X2 U4 ( .A(n57), .B(n48), .Y(n58) );
  BUFX8 U5 ( .A(n252), .Y(out[3]) );
  OAI21X1 U6 ( .A0(n36), .A1(n68), .B0(n67), .Y(n72) );
  NAND2X1 U7 ( .A(n36), .B(n8), .Y(n67) );
  MX2X1 U8 ( .A(neg_mul[20]), .B(N478), .S0(n81), .Y(out[13]) );
  MX2X1 U9 ( .A(neg_mul[22]), .B(N480), .S0(n81), .Y(out[15]) );
  NAND2X1 U10 ( .A(n36), .B(n15), .Y(n60) );
  MX2X1 U11 ( .A(neg_mul[21]), .B(N479), .S0(n81), .Y(out[14]) );
  INVX1 U12 ( .A(n90), .Y(n86) );
  BUFX8 U13 ( .A(in_8bit[7]), .Y(n36) );
  CLKINVX8 U14 ( .A(in_17bit[16]), .Y(n49) );
  INVX1 U15 ( .A(n19), .Y(n50) );
  INVX1 U16 ( .A(in_8bit[7]), .Y(n42) );
  XNOR2X1 U17 ( .A(neg_mul[23]), .B(n34), .Y(n17) );
  NOR2BX4 U18 ( .AN(n53), .B(n73), .Y(n75) );
  NOR2X2 U19 ( .A(n70), .B(n48), .Y(n71) );
  INVXL U20 ( .A(n37), .Y(n19) );
  XOR2X4 U21 ( .A(n77), .B(neg_mul[13]), .Y(out[6]) );
  NOR2X2 U22 ( .A(n48), .B(n62), .Y(n64) );
  INVXL U23 ( .A(n19), .Y(n20) );
  AOI211X2 U24 ( .A0(n37), .A1(n72), .B0(n71), .C0(n74), .Y(n252) );
  INVX8 U25 ( .A(n80), .Y(n81) );
  XNOR2X4 U26 ( .A(n37), .B(n36), .Y(n78) );
  INVX8 U27 ( .A(n49), .Y(n48) );
  XNOR2X4 U28 ( .A(n37), .B(n36), .Y(n73) );
  INVX8 U29 ( .A(n49), .Y(n37) );
  XNOR2X4 U30 ( .A(n22), .B(n7), .Y(out[9]) );
  NOR2X4 U31 ( .A(n80), .B(n31), .Y(n22) );
  XNOR2X4 U32 ( .A(n21), .B(n3), .Y(out[8]) );
  NOR2X4 U33 ( .A(n80), .B(n29), .Y(n21) );
  NOR2X4 U34 ( .A(n27), .B(n73), .Y(n77) );
  AOI2BB2X1 U35 ( .B0(n42), .B1(n15), .A0N(n61), .A1N(n42), .Y(n62) );
  MX2X4 U36 ( .A(neg_mul[19]), .B(N477), .S0(n81), .Y(out[12]) );
  AOI2BB2X1 U37 ( .B0(n56), .B1(n36), .A0N(in_8bit[7]), .A1N(neg_mul[8]), .Y(
        n57) );
  XNOR2X4 U38 ( .A(n37), .B(n36), .Y(n80) );
  INVX1 U39 ( .A(n201), .Y(in_17bit_b[1]) );
  INVX1 U40 ( .A(n240), .Y(in_17bit_b[14]) );
  INVX1 U41 ( .A(n237), .Y(in_17bit_b[13]) );
  INVX1 U42 ( .A(n204), .Y(in_17bit_b[2]) );
  INVX1 U43 ( .A(n213), .Y(in_17bit_b[5]) );
  INVX1 U44 ( .A(n222), .Y(in_17bit_b[8]) );
  INVX1 U45 ( .A(n216), .Y(in_17bit_b[6]) );
  INVX1 U46 ( .A(n219), .Y(in_17bit_b[7]) );
  INVX1 U47 ( .A(n225), .Y(in_17bit_b[9]) );
  INVX1 U48 ( .A(n231), .Y(in_17bit_b[11]) );
  INVX1 U49 ( .A(n228), .Y(in_17bit_b[10]) );
  INVX1 U50 ( .A(n234), .Y(in_17bit_b[12]) );
  INVX1 U51 ( .A(n210), .Y(in_17bit_b[4]) );
  INVX1 U52 ( .A(n207), .Y(in_17bit_b[3]) );
  AOI21X1 U53 ( .A0(n23), .A1(n24), .B0(n244), .Y(n197) );
  NOR4XL U54 ( .A(in_8bit[4]), .B(in_8bit[5]), .C(in_8bit[6]), .D(n36), .Y(n23) );
  NOR4X1 U55 ( .A(n41), .B(in_8bit[0]), .C(n46), .D(in_8bit[3]), .Y(n24) );
  AND4X1 U56 ( .A(n41), .B(n36), .C(n191), .D(n43), .Y(n25) );
  BUFX3 U57 ( .A(in_8bit[1]), .Y(n41) );
  INVX1 U58 ( .A(n47), .Y(n46) );
  INVX1 U59 ( .A(in_8bit[2]), .Y(n47) );
  INVX1 U60 ( .A(in_8bit[6]), .Y(n44) );
  NOR3X1 U61 ( .A(n47), .B(n45), .C(n43), .Y(n196) );
  NOR4BX1 U62 ( .AN(n194), .B(n43), .C(n41), .D(n46), .Y(n195) );
  NOR2X1 U63 ( .A(in_8bit[6]), .B(in_8bit[3]), .Y(n194) );
  NAND3X1 U64 ( .A(n46), .B(n45), .C(in_8bit[5]), .Y(n192) );
  ADDFX2 U65 ( .A(n40), .B(in_17bit_b[12]), .CI(add_1_root_r112_carry_16_), 
        .CO(add_1_root_r112_carry_17_), .S(add_1_root_r112_SUM_16_) );
  ADDFX2 U66 ( .A(add_1_root_r119_A_19_), .B(in_17bit_b[13]), .CI(
        add_1_root_r119_carry[19]), .CO(add_1_root_r119_carry[20]), .S(
        add_1_root_r119_SUM_19_) );
  ADDFX2 U67 ( .A(n40), .B(in_17bit_b[15]), .CI(add_3_root_r119_carry_17_), 
        .CO(add_3_root_r119_carry_18_), .S(add_1_root_r119_A_17_) );
  ADDFX2 U68 ( .A(n40), .B(in_17bit_b[14]), .CI(add_2_root_r115_carry_17_), 
        .CO(add_2_root_r115_carry_18_), .S(add_2_root_r115_SUM_17_) );
  ADDFX2 U69 ( .A(n40), .B(in_17bit_b[14]), .CI(add_1_root_r115_carry_20_), 
        .CO(add_1_root_r115_carry_21_), .S(add_1_root_r115_SUM_20_) );
  ADDFX2 U70 ( .A(n40), .B(in_17bit_b[15]), .CI(add_2_root_r119_carry_20_), 
        .CO(add_2_root_r119_carry_21_), .S(add_2_root_r119_SUM_20_) );
  ADDFX2 U71 ( .A(in_17bit_b[3]), .B(in_17bit_b[1]), .CI(
        add_2_root_r115_carry_4_), .CO(add_2_root_r115_carry_5_), .S(
        add_2_root_r115_SUM_4_) );
  ADDFX2 U72 ( .A(in_17bit_b[4]), .B(in_17bit_b[2]), .CI(
        add_2_root_r115_carry_5_), .CO(add_2_root_r115_carry_6_), .S(
        add_2_root_r115_SUM_5_) );
  ADDFX2 U73 ( .A(in_17bit_b[5]), .B(in_17bit_b[1]), .CI(
        add_1_root_r112_carry_5_), .CO(add_1_root_r112_carry_6_), .S(
        add_1_root_r112_SUM_5_) );
  ADDFX2 U74 ( .A(in_17bit_b[6]), .B(in_17bit_b[5]), .CI(
        add_3_root_r119_carry_7_), .CO(add_3_root_r119_carry_8_), .S(
        add_1_root_r119_A_7_) );
  ADDFX2 U75 ( .A(in_17bit_b[6]), .B(in_17bit_b[2]), .CI(
        add_1_root_r112_carry_6_), .CO(add_1_root_r112_carry_7_), .S(
        add_1_root_r112_SUM_6_) );
  ADDFX2 U76 ( .A(in_17bit_b[3]), .B(in_17bit_b[1]), .CI(
        add_1_root_r115_carry_7_), .CO(add_1_root_r115_carry_8_), .S(
        add_1_root_r115_SUM_7_) );
  ADDFX2 U77 ( .A(in_17bit_b[7]), .B(in_17bit_b[6]), .CI(
        add_3_root_r119_carry_8_), .CO(add_3_root_r119_carry_9_), .S(
        add_1_root_r119_A_8_) );
  ADDFX2 U78 ( .A(add_1_root_r119_A_7_), .B(in_17bit_b[1]), .CI(
        add_1_root_r119_carry[7]), .CO(add_1_root_r119_carry[8]), .S(
        add_1_root_r119_SUM_7_) );
  ADDFX2 U79 ( .A(in_17bit_b[2]), .B(in_17bit_b[1]), .CI(
        add_2_root_r119_carry_6_), .CO(add_2_root_r119_carry_7_), .S(
        add_2_root_r119_SUM_6_) );
  ADDFX2 U80 ( .A(in_17bit_b[4]), .B(in_17bit_b[2]), .CI(
        add_1_root_r115_carry_8_), .CO(add_1_root_r115_carry_9_), .S(
        add_1_root_r115_SUM_8_) );
  ADDFX2 U81 ( .A(in_17bit_b[8]), .B(in_17bit_b[7]), .CI(
        add_3_root_r119_carry_9_), .CO(add_3_root_r119_carry_10_), .S(
        add_1_root_r119_A_9_) );
  ADDFX2 U82 ( .A(add_1_root_r119_A_8_), .B(in_17bit_b[2]), .CI(
        add_1_root_r119_carry[8]), .CO(add_1_root_r119_carry[9]), .S(
        add_1_root_r119_SUM_8_) );
  ADDFX2 U83 ( .A(in_17bit_b[3]), .B(in_17bit_b[2]), .CI(
        add_2_root_r119_carry_7_), .CO(add_2_root_r119_carry_8_), .S(
        add_2_root_r119_SUM_7_) );
  ADDFX2 U84 ( .A(in_17bit_b[6]), .B(in_17bit_b[4]), .CI(
        add_2_root_r115_carry_7_), .CO(add_2_root_r115_carry_8_), .S(
        add_2_root_r115_SUM_7_) );
  ADDFX2 U85 ( .A(in_17bit_b[8]), .B(in_17bit_b[4]), .CI(
        add_1_root_r112_carry_8_), .CO(add_1_root_r112_carry_9_), .S(
        add_1_root_r112_SUM_8_) );
  ADDFX2 U86 ( .A(in_17bit_b[9]), .B(in_17bit_b[8]), .CI(
        add_3_root_r119_carry_10_), .CO(add_3_root_r119_carry_11_), .S(
        add_1_root_r119_A_10_) );
  ADDFX2 U87 ( .A(in_17bit_b[6]), .B(in_17bit_b[4]), .CI(
        add_1_root_r115_carry_10_), .CO(add_1_root_r115_carry_11_), .S(
        add_1_root_r115_SUM_10_) );
  ADDFX2 U88 ( .A(in_17bit_b[7]), .B(in_17bit_b[5]), .CI(
        add_2_root_r115_carry_8_), .CO(add_2_root_r115_carry_9_), .S(
        add_2_root_r115_SUM_8_) );
  ADDFX2 U89 ( .A(in_17bit_b[9]), .B(in_17bit_b[5]), .CI(
        add_1_root_r112_carry_9_), .CO(add_1_root_r112_carry_10_), .S(
        add_1_root_r112_SUM_9_) );
  ADDFX2 U90 ( .A(in_17bit_b[10]), .B(in_17bit_b[9]), .CI(
        add_3_root_r119_carry_11_), .CO(add_3_root_r119_carry_12_), .S(
        add_1_root_r119_A_11_) );
  ADDFX2 U91 ( .A(add_1_root_r119_A_10_), .B(in_17bit_b[4]), .CI(
        add_1_root_r119_carry[10]), .CO(add_1_root_r119_carry[11]), .S(
        add_1_root_r119_SUM_10_) );
  ADDFX2 U92 ( .A(in_17bit_b[5]), .B(in_17bit_b[4]), .CI(
        add_2_root_r119_carry_9_), .CO(add_2_root_r119_carry_10_), .S(
        add_2_root_r119_SUM_9_) );
  ADDFX2 U93 ( .A(in_17bit_b[8]), .B(in_17bit_b[6]), .CI(
        add_2_root_r115_carry_9_), .CO(add_2_root_r115_carry_10_), .S(
        add_2_root_r115_SUM_9_) );
  ADDFX2 U94 ( .A(in_17bit_b[10]), .B(in_17bit_b[6]), .CI(
        add_1_root_r112_carry_10_), .CO(add_1_root_r112_carry_11_), .S(
        add_1_root_r112_SUM_10_) );
  ADDFX2 U95 ( .A(in_17bit_b[7]), .B(in_17bit_b[5]), .CI(
        add_1_root_r115_carry_11_), .CO(add_1_root_r115_carry_12_), .S(
        add_1_root_r115_SUM_11_) );
  ADDFX2 U96 ( .A(in_17bit_b[11]), .B(in_17bit_b[10]), .CI(
        add_3_root_r119_carry_12_), .CO(add_3_root_r119_carry_13_), .S(
        add_1_root_r119_A_12_) );
  ADDFX2 U97 ( .A(add_1_root_r119_A_11_), .B(in_17bit_b[5]), .CI(
        add_1_root_r119_carry[11]), .CO(add_1_root_r119_carry[12]), .S(
        add_1_root_r119_SUM_11_) );
  ADDFX2 U98 ( .A(in_17bit_b[6]), .B(in_17bit_b[5]), .CI(
        add_2_root_r119_carry_10_), .CO(add_2_root_r119_carry_11_), .S(
        add_2_root_r119_SUM_10_) );
  ADDFX2 U99 ( .A(in_17bit_b[9]), .B(in_17bit_b[7]), .CI(
        add_2_root_r115_carry_10_), .CO(add_2_root_r115_carry_11_), .S(
        add_2_root_r115_SUM_10_) );
  ADDFX2 U100 ( .A(in_17bit_b[11]), .B(in_17bit_b[7]), .CI(
        add_1_root_r112_carry_11_), .CO(add_1_root_r112_carry_12_), .S(
        add_1_root_r112_SUM_11_) );
  ADDFX2 U101 ( .A(in_17bit_b[8]), .B(in_17bit_b[6]), .CI(
        add_1_root_r115_carry_12_), .CO(add_1_root_r115_carry_13_), .S(
        add_1_root_r115_SUM_12_) );
  ADDFX2 U102 ( .A(in_17bit_b[12]), .B(in_17bit_b[11]), .CI(
        add_3_root_r119_carry_13_), .CO(add_3_root_r119_carry_14_), .S(
        add_1_root_r119_A_13_) );
  ADDFX2 U103 ( .A(add_1_root_r119_A_12_), .B(in_17bit_b[6]), .CI(
        add_1_root_r119_carry[12]), .CO(add_1_root_r119_carry[13]), .S(
        add_1_root_r119_SUM_12_) );
  ADDFX2 U104 ( .A(in_17bit_b[7]), .B(in_17bit_b[6]), .CI(
        add_2_root_r119_carry_11_), .CO(add_2_root_r119_carry_12_), .S(
        add_2_root_r119_SUM_11_) );
  ADDFX2 U105 ( .A(in_17bit_b[12]), .B(in_17bit_b[8]), .CI(
        add_1_root_r112_carry_12_), .CO(add_1_root_r112_carry_13_), .S(
        add_1_root_r112_SUM_12_) );
  ADDFX2 U106 ( .A(in_17bit_b[9]), .B(in_17bit_b[7]), .CI(
        add_1_root_r115_carry_13_), .CO(add_1_root_r115_carry_14_), .S(
        add_1_root_r115_SUM_13_) );
  ADDFX2 U107 ( .A(in_17bit_b[13]), .B(in_17bit_b[12]), .CI(
        add_3_root_r119_carry_14_), .CO(add_3_root_r119_carry_15_), .S(
        add_1_root_r119_A_14_) );
  ADDFX2 U108 ( .A(add_1_root_r119_A_13_), .B(in_17bit_b[7]), .CI(
        add_1_root_r119_carry[13]), .CO(add_1_root_r119_carry[14]), .S(
        add_1_root_r119_SUM_13_) );
  ADDFX2 U109 ( .A(in_17bit_b[8]), .B(in_17bit_b[7]), .CI(
        add_2_root_r119_carry_12_), .CO(add_2_root_r119_carry_13_), .S(
        add_2_root_r119_SUM_12_) );
  ADDFX2 U110 ( .A(in_17bit_b[11]), .B(in_17bit_b[9]), .CI(
        add_2_root_r115_carry_12_), .CO(add_2_root_r115_carry_13_), .S(
        add_2_root_r115_SUM_12_) );
  ADDFX2 U111 ( .A(in_17bit_b[13]), .B(in_17bit_b[9]), .CI(
        add_1_root_r112_carry_13_), .CO(add_1_root_r112_carry_14_), .S(
        add_1_root_r112_SUM_13_) );
  ADDFX2 U112 ( .A(in_17bit_b[10]), .B(in_17bit_b[8]), .CI(
        add_1_root_r115_carry_14_), .CO(add_1_root_r115_carry_15_), .S(
        add_1_root_r115_SUM_14_) );
  ADDFX2 U113 ( .A(in_17bit_b[14]), .B(in_17bit_b[13]), .CI(
        add_3_root_r119_carry_15_), .CO(add_3_root_r119_carry_16_), .S(
        add_1_root_r119_A_15_) );
  ADDFX2 U114 ( .A(add_1_root_r119_A_14_), .B(in_17bit_b[8]), .CI(
        add_1_root_r119_carry[14]), .CO(add_1_root_r119_carry[15]), .S(
        add_1_root_r119_SUM_14_) );
  ADDFX2 U115 ( .A(in_17bit_b[9]), .B(in_17bit_b[8]), .CI(
        add_2_root_r119_carry_13_), .CO(add_2_root_r119_carry_14_), .S(
        add_2_root_r119_SUM_13_) );
  ADDFX2 U116 ( .A(in_17bit_b[12]), .B(in_17bit_b[10]), .CI(
        add_2_root_r115_carry_13_), .CO(add_2_root_r115_carry_14_), .S(
        add_2_root_r115_SUM_13_) );
  ADDFX2 U117 ( .A(in_17bit_b[14]), .B(in_17bit_b[10]), .CI(
        add_1_root_r112_carry_14_), .CO(add_1_root_r112_carry_15_), .S(
        add_1_root_r112_SUM_14_) );
  ADDFX2 U118 ( .A(in_17bit_b[11]), .B(in_17bit_b[9]), .CI(
        add_1_root_r115_carry_15_), .CO(add_1_root_r115_carry_16_), .S(
        add_1_root_r115_SUM_15_) );
  ADDFX2 U119 ( .A(add_1_root_r119_A_15_), .B(in_17bit_b[9]), .CI(
        add_1_root_r119_carry[15]), .CO(add_1_root_r119_carry[16]), .S(
        add_1_root_r119_SUM_15_) );
  ADDFX2 U120 ( .A(in_17bit_b[3]), .B(in_17bit_b[2]), .CI(
        add_3_root_r119_carry_4_), .CO(add_3_root_r119_carry_5_), .S(
        add_1_root_r119_A_4_) );
  ADDFX2 U121 ( .A(in_17bit_b[2]), .B(in_17bit_b[1]), .CI(
        add_3_root_r119_carry_3_), .CO(add_3_root_r119_carry_4_), .S(
        add_1_root_r119_A_3_) );
  ADDFX2 U122 ( .A(in_17bit_b[10]), .B(in_17bit_b[9]), .CI(
        add_2_root_r119_carry_14_), .CO(add_2_root_r119_carry_15_), .S(
        add_2_root_r119_SUM_14_) );
  ADDFX2 U123 ( .A(in_17bit_b[13]), .B(in_17bit_b[11]), .CI(
        add_2_root_r115_carry_14_), .CO(add_2_root_r115_carry_15_), .S(
        add_2_root_r115_SUM_14_) );
  ADDFX2 U124 ( .A(in_17bit_b[15]), .B(in_17bit_b[11]), .CI(
        add_1_root_r112_carry_15_), .CO(add_1_root_r112_carry_16_), .S(
        add_1_root_r112_SUM_15_) );
  ADDFX2 U125 ( .A(in_17bit_b[12]), .B(in_17bit_b[10]), .CI(
        add_1_root_r115_carry_16_), .CO(add_1_root_r115_carry_17_), .S(
        add_1_root_r115_SUM_16_) );
  ADDFX2 U126 ( .A(add_1_root_r119_A_16_), .B(in_17bit_b[10]), .CI(
        add_1_root_r119_carry[16]), .CO(add_1_root_r119_carry[17]), .S(
        add_1_root_r119_SUM_16_) );
  ADDFX2 U127 ( .A(in_17bit_b[11]), .B(in_17bit_b[10]), .CI(
        add_2_root_r119_carry_15_), .CO(add_2_root_r119_carry_16_), .S(
        add_2_root_r119_SUM_15_) );
  ADDFX2 U128 ( .A(in_17bit_b[14]), .B(in_17bit_b[12]), .CI(
        add_2_root_r115_carry_15_), .CO(add_2_root_r115_carry_16_), .S(
        add_2_root_r115_SUM_15_) );
  ADDFX2 U129 ( .A(in_17bit_b[13]), .B(in_17bit_b[11]), .CI(
        add_1_root_r115_carry_17_), .CO(add_1_root_r115_carry_18_), .S(
        add_1_root_r115_SUM_17_) );
  ADDFX2 U130 ( .A(add_1_root_r119_A_17_), .B(in_17bit_b[11]), .CI(
        add_1_root_r119_carry[17]), .CO(add_1_root_r119_carry[18]), .S(
        add_1_root_r119_SUM_17_) );
  ADDFX2 U131 ( .A(in_17bit_b[12]), .B(in_17bit_b[11]), .CI(
        add_2_root_r119_carry_16_), .CO(add_2_root_r119_carry_17_), .S(
        add_2_root_r119_SUM_16_) );
  ADDFX2 U132 ( .A(in_17bit_b[15]), .B(in_17bit_b[13]), .CI(
        add_2_root_r115_carry_16_), .CO(add_2_root_r115_carry_17_), .S(
        add_2_root_r115_SUM_16_) );
  ADDFX2 U133 ( .A(in_17bit_b[14]), .B(in_17bit_b[12]), .CI(
        add_1_root_r115_carry_18_), .CO(add_1_root_r115_carry_19_), .S(
        add_1_root_r115_SUM_18_) );
  ADDFX2 U134 ( .A(add_1_root_r119_A_18_), .B(in_17bit_b[12]), .CI(
        add_1_root_r119_carry[18]), .CO(add_1_root_r119_carry[19]), .S(
        add_1_root_r119_SUM_18_) );
  ADDFX2 U135 ( .A(in_17bit_b[13]), .B(in_17bit_b[12]), .CI(
        add_2_root_r119_carry_17_), .CO(add_2_root_r119_carry_18_), .S(
        add_2_root_r119_SUM_17_) );
  ADDFX2 U136 ( .A(in_17bit_b[5]), .B(in_17bit_b[3]), .CI(
        add_2_root_r115_carry_6_), .CO(add_2_root_r115_carry_7_), .S(
        add_2_root_r115_SUM_6_) );
  ADDFX2 U137 ( .A(in_17bit_b[7]), .B(in_17bit_b[3]), .CI(
        add_1_root_r112_carry_7_), .CO(add_1_root_r112_carry_8_), .S(
        add_1_root_r112_SUM_7_) );
  ADDFX2 U138 ( .A(in_17bit_b[5]), .B(in_17bit_b[3]), .CI(
        add_1_root_r115_carry_9_), .CO(add_1_root_r115_carry_10_), .S(
        add_1_root_r115_SUM_9_) );
  ADDFX2 U139 ( .A(in_17bit_b[15]), .B(in_17bit_b[13]), .CI(
        add_1_root_r115_carry_19_), .CO(add_1_root_r115_carry_20_), .S(
        add_1_root_r115_SUM_19_) );
  ADDFX2 U140 ( .A(add_1_root_r119_A_9_), .B(in_17bit_b[3]), .CI(
        add_1_root_r119_carry[9]), .CO(add_1_root_r119_carry[10]), .S(
        add_1_root_r119_SUM_9_) );
  ADDFX2 U141 ( .A(in_17bit_b[4]), .B(in_17bit_b[3]), .CI(
        add_2_root_r119_carry_8_), .CO(add_2_root_r119_carry_9_), .S(
        add_2_root_r119_SUM_8_) );
  ADDFX2 U142 ( .A(in_17bit_b[10]), .B(in_17bit_b[8]), .CI(
        add_2_root_r115_carry_11_), .CO(add_2_root_r115_carry_12_), .S(
        add_2_root_r115_SUM_11_) );
  ADDFX2 U143 ( .A(in_17bit_b[15]), .B(in_17bit_b[14]), .CI(
        add_3_root_r119_carry_16_), .CO(add_3_root_r119_carry_17_), .S(
        add_1_root_r119_A_16_) );
  ADDFX2 U144 ( .A(in_17bit_b[14]), .B(in_17bit_b[13]), .CI(
        add_2_root_r119_carry_18_), .CO(add_2_root_r119_carry_19_), .S(
        add_2_root_r119_SUM_18_) );
  ADDFX2 U145 ( .A(in_17bit_b[4]), .B(in_17bit_b[3]), .CI(
        add_3_root_r119_carry_5_), .CO(add_3_root_r119_carry_6_), .S(
        add_1_root_r119_A_5_) );
  ADDFX2 U146 ( .A(in_17bit_b[5]), .B(in_17bit_b[4]), .CI(
        add_3_root_r119_carry_6_), .CO(add_3_root_r119_carry_7_), .S(
        add_1_root_r119_A_6_) );
  ADDFX2 U147 ( .A(in_17bit_b[15]), .B(in_17bit_b[14]), .CI(
        add_2_root_r119_carry_19_), .CO(add_2_root_r119_carry_20_), .S(
        add_2_root_r119_SUM_19_) );
  BUFX3 U148 ( .A(in_17bit_b[16]), .Y(n40) );
  INVX1 U149 ( .A(n251), .Y(in_17bit_b[16]) );
  INVX1 U150 ( .A(n193), .Y(n89) );
  NAND3BX1 U151 ( .AN(in_8bit[5]), .B(n47), .C(in_8bit[3]), .Y(n193) );
  INVX1 U152 ( .A(in_8bit[0]), .Y(n43) );
  INVXL U153 ( .A(n20), .Y(n52) );
  INVXL U154 ( .A(n50), .Y(n51) );
  CLKINVX3 U155 ( .A(n198), .Y(in_17bit_b[0]) );
  INVX1 U156 ( .A(n171), .Y(n250) );
  NAND2XL U157 ( .A(N29), .B(n50), .Y(n251) );
  OAI21XL U158 ( .A0(n250), .A1(n251), .B0(n249), .Y(N463) );
  AOI22X1 U159 ( .A0(N221), .A1(n39), .B0(N363), .B1(n38), .Y(n249) );
  CLKINVX3 U160 ( .A(n243), .Y(in_17bit_b[15]) );
  NAND2X1 U161 ( .A(n200), .B(n199), .Y(N447) );
  AOI22X1 U162 ( .A0(N108), .A1(n244), .B0(N205), .B1(n39), .Y(n199) );
  AOI22X1 U163 ( .A0(N347), .A1(n38), .B0(n171), .B1(in_17bit_b[0]), .Y(n200)
         );
  NAND2X1 U164 ( .A(n203), .B(n202), .Y(N448) );
  AOI22X1 U165 ( .A0(N109), .A1(n244), .B0(N206), .B1(n39), .Y(n202) );
  AOI22X1 U166 ( .A0(N348), .A1(n38), .B0(n171), .B1(n170), .Y(n203) );
  INVX1 U167 ( .A(n201), .Y(n170) );
  NAND2X1 U168 ( .A(n206), .B(n205), .Y(N449) );
  AOI22X1 U169 ( .A0(N110), .A1(n244), .B0(N207), .B1(n39), .Y(n205) );
  AOI22X1 U170 ( .A0(N349), .A1(n38), .B0(n171), .B1(in_17bit_b[2]), .Y(n206)
         );
  NAND2X1 U171 ( .A(n209), .B(n208), .Y(N450) );
  AOI22X1 U172 ( .A0(N111), .A1(n244), .B0(N208), .B1(n39), .Y(n208) );
  AOI22X1 U173 ( .A0(N350), .A1(n38), .B0(n171), .B1(in_17bit_b[3]), .Y(n209)
         );
  NAND2X1 U174 ( .A(n212), .B(n211), .Y(N451) );
  AOI22X1 U175 ( .A0(N112), .A1(n244), .B0(N209), .B1(n39), .Y(n211) );
  AOI22X1 U176 ( .A0(N351), .A1(n38), .B0(n171), .B1(in_17bit_b[4]), .Y(n212)
         );
  NAND2X1 U177 ( .A(n215), .B(n214), .Y(N452) );
  AOI22X1 U178 ( .A0(N113), .A1(n244), .B0(N210), .B1(n39), .Y(n214) );
  AOI22X1 U179 ( .A0(N352), .A1(n38), .B0(n171), .B1(in_17bit_b[5]), .Y(n215)
         );
  NAND2X1 U180 ( .A(n218), .B(n217), .Y(N453) );
  AOI22X1 U181 ( .A0(N114), .A1(n244), .B0(N211), .B1(n39), .Y(n217) );
  AOI22X1 U182 ( .A0(N353), .A1(n38), .B0(n171), .B1(in_17bit_b[6]), .Y(n218)
         );
  NAND2X1 U183 ( .A(n221), .B(n220), .Y(N454) );
  AOI22X1 U184 ( .A0(N115), .A1(n244), .B0(N212), .B1(n39), .Y(n220) );
  AOI22X1 U185 ( .A0(N354), .A1(n38), .B0(n171), .B1(in_17bit_b[7]), .Y(n221)
         );
  NAND2X1 U186 ( .A(n224), .B(n223), .Y(N455) );
  AOI22X1 U187 ( .A0(N116), .A1(n244), .B0(N213), .B1(n39), .Y(n223) );
  AOI22X1 U188 ( .A0(N355), .A1(n38), .B0(n171), .B1(in_17bit_b[8]), .Y(n224)
         );
  NAND2X1 U189 ( .A(n227), .B(n226), .Y(N456) );
  AOI22X1 U190 ( .A0(N117), .A1(n244), .B0(N214), .B1(n39), .Y(n226) );
  AOI22X1 U191 ( .A0(N356), .A1(n38), .B0(n171), .B1(in_17bit_b[9]), .Y(n227)
         );
  NAND2X1 U192 ( .A(n230), .B(n229), .Y(N457) );
  AOI22X1 U193 ( .A0(N118), .A1(n244), .B0(N215), .B1(n39), .Y(n229) );
  AOI22X1 U194 ( .A0(N357), .A1(n38), .B0(n171), .B1(in_17bit_b[10]), .Y(n230)
         );
  NAND2X1 U195 ( .A(n233), .B(n232), .Y(N458) );
  AOI22X1 U196 ( .A0(N119), .A1(n244), .B0(N216), .B1(n39), .Y(n232) );
  AOI22X1 U197 ( .A0(N358), .A1(n38), .B0(n171), .B1(in_17bit_b[11]), .Y(n233)
         );
  NAND2X1 U198 ( .A(n236), .B(n235), .Y(N459) );
  AOI22X1 U199 ( .A0(N120), .A1(n244), .B0(N217), .B1(n39), .Y(n235) );
  AOI22X1 U200 ( .A0(N359), .A1(n38), .B0(n171), .B1(in_17bit_b[12]), .Y(n236)
         );
  NAND2X1 U201 ( .A(n239), .B(n238), .Y(N460) );
  AOI22X1 U202 ( .A0(N121), .A1(n244), .B0(N218), .B1(n39), .Y(n238) );
  AOI22X1 U203 ( .A0(N360), .A1(n38), .B0(n171), .B1(in_17bit_b[13]), .Y(n239)
         );
  NAND2X1 U204 ( .A(n242), .B(n241), .Y(N461) );
  AOI22X1 U205 ( .A0(N122), .A1(n244), .B0(N219), .B1(n39), .Y(n241) );
  AOI22X1 U206 ( .A0(N361), .A1(n38), .B0(n171), .B1(in_17bit_b[14]), .Y(n242)
         );
  NAND2X1 U207 ( .A(n246), .B(n245), .Y(N462) );
  AOI22X1 U208 ( .A0(N123), .A1(n244), .B0(N220), .B1(n39), .Y(n245) );
  AOI22X1 U209 ( .A0(N362), .A1(n38), .B0(n171), .B1(in_17bit_b[15]), .Y(n246)
         );
  INVX1 U210 ( .A(in_8bit[3]), .Y(n45) );
  OAI21XL U211 ( .A0(n36), .A1(n55), .B0(n54), .Y(n59) );
  INVX1 U212 ( .A(n66), .Y(n63) );
  OAI21XL U213 ( .A0(n36), .A1(n61), .B0(n60), .Y(n65) );
  MXI2XL U214 ( .A(n2), .B(n17), .S0(n81), .Y(out[16]) );
  AOI22XL U215 ( .A0(in_17bit[0]), .A1(n20), .B0(in_17bit[0]), .B1(n52), .Y(
        n198) );
  AOI22X1 U216 ( .A0(N27), .A1(n50), .B0(in_17bit[14]), .B1(n19), .Y(n240) );
  AOI22X1 U217 ( .A0(N28), .A1(n50), .B0(in_17bit[15]), .B1(n52), .Y(n243) );
  AOI22XL U218 ( .A0(N14), .A1(n50), .B0(in_17bit[1]), .B1(n52), .Y(n201) );
  AOI22XL U219 ( .A0(N15), .A1(n20), .B0(in_17bit[2]), .B1(n51), .Y(n204) );
  AOI22X1 U220 ( .A0(N16), .A1(n50), .B0(in_17bit[3]), .B1(n51), .Y(n207) );
  AOI22X1 U221 ( .A0(N17), .A1(n50), .B0(in_17bit[4]), .B1(n19), .Y(n210) );
  AOI22X1 U222 ( .A0(N18), .A1(n50), .B0(in_17bit[5]), .B1(n52), .Y(n213) );
  AOI22X1 U223 ( .A0(N19), .A1(n50), .B0(in_17bit[6]), .B1(n19), .Y(n216) );
  AOI22X1 U224 ( .A0(N20), .A1(n50), .B0(in_17bit[7]), .B1(n51), .Y(n219) );
  AOI22X1 U225 ( .A0(N21), .A1(n50), .B0(in_17bit[8]), .B1(n51), .Y(n222) );
  AOI22X1 U226 ( .A0(N22), .A1(n50), .B0(in_17bit[9]), .B1(n51), .Y(n225) );
  AOI22X1 U227 ( .A0(N23), .A1(n50), .B0(in_17bit[10]), .B1(n19), .Y(n228) );
  AOI22X1 U228 ( .A0(N24), .A1(n50), .B0(in_17bit[11]), .B1(n19), .Y(n231) );
  AOI22X1 U229 ( .A0(N25), .A1(n50), .B0(in_17bit[12]), .B1(n51), .Y(n234) );
  AOI22X1 U230 ( .A0(N26), .A1(n50), .B0(in_17bit[13]), .B1(n52), .Y(n237) );
  INVX1 U231 ( .A(n53), .Y(n74) );
  NAND2BX1 U232 ( .AN(n66), .B(n8), .Y(n53) );
  NAND2X1 U233 ( .A(n33), .B(n15), .Y(n66) );
  AND2X2 U234 ( .A(n74), .B(n4), .Y(n26) );
  AND2X2 U235 ( .A(n26), .B(n5), .Y(n27) );
  AND2X2 U236 ( .A(n27), .B(n1), .Y(n28) );
  AND2X2 U237 ( .A(n28), .B(n6), .Y(n29) );
  BUFX3 U238 ( .A(n247), .Y(n38) );
  OAI2BB1X1 U239 ( .A0N(n89), .A1N(n25), .B0(n87), .Y(n247) );
  NAND2BX1 U240 ( .AN(n192), .B(n30), .Y(n87) );
  BUFX3 U241 ( .A(n248), .Y(n39) );
  OAI2BB1X1 U242 ( .A0N(n30), .A1N(n89), .B0(n88), .Y(n248) );
  NAND2BX1 U243 ( .AN(n192), .B(n25), .Y(n88) );
  NAND2X1 U244 ( .A(n85), .B(n84), .Y(n244) );
  NAND3X1 U245 ( .A(n195), .B(in_8bit[5]), .C(n83), .Y(n84) );
  NAND4BXL U246 ( .AN(n44), .B(n196), .C(n92), .D(n41), .Y(n85) );
  OAI2BB1X1 U247 ( .A0N(n195), .A1N(n92), .B0(n91), .Y(n171) );
  NAND3BX1 U248 ( .AN(n90), .B(n196), .C(in_8bit[5]), .Y(n91) );
  AND2X2 U249 ( .A(n86), .B(n43), .Y(n30) );
  AND2X2 U250 ( .A(n29), .B(n3), .Y(n31) );
  INVX1 U251 ( .A(in_17bit[13]), .Y(n163) );
  INVX1 U252 ( .A(in_17bit[2]), .Y(n95) );
  INVX1 U253 ( .A(in_17bit[4]), .Y(n97) );
  INVX1 U254 ( .A(in_17bit[5]), .Y(n98) );
  INVX1 U255 ( .A(in_17bit[6]), .Y(n99) );
  INVX1 U256 ( .A(in_17bit[7]), .Y(n100) );
  INVX1 U257 ( .A(in_17bit[8]), .Y(n101) );
  INVX1 U258 ( .A(in_17bit[9]), .Y(n158) );
  INVX1 U259 ( .A(in_17bit[10]), .Y(n160) );
  INVX1 U260 ( .A(in_17bit[11]), .Y(n161) );
  INVX1 U261 ( .A(in_17bit[12]), .Y(n162) );
  INVX1 U262 ( .A(in_17bit[14]), .Y(n164) );
  INVX1 U263 ( .A(in_17bit[15]), .Y(n168) );
  INVX1 U264 ( .A(in_17bit[1]), .Y(n94) );
  INVX1 U265 ( .A(in_17bit[3]), .Y(n96) );
  INVX1 U266 ( .A(in_17bit[0]), .Y(n93) );
  XNOR2X1 U267 ( .A(n14), .B(sub_add_75_b0_carry[10]), .Y(n32) );
  MX2X4 U268 ( .A(neg_mul[18]), .B(N476), .S0(n81), .Y(out[11]) );
  INVX1 U269 ( .A(n55), .Y(n56) );
  AOI2BB2X2 U270 ( .B0(n69), .B1(n36), .A0N(in_8bit[7]), .A1N(neg_mul[10]), 
        .Y(n70) );
  INVX1 U271 ( .A(n68), .Y(n69) );
  NAND4BBX1 U272 ( .AN(n38), .BN(n39), .C(n197), .D(n250), .Y(N446) );
  NOR3BXL U273 ( .AN(in_8bit[7]), .B(in_8bit[5]), .C(in_8bit[4]), .Y(n92) );
  NAND4BXL U274 ( .AN(in_8bit[7]), .B(in_8bit[4]), .C(n41), .D(in_8bit[6]), 
        .Y(n90) );
  NOR2X1 U275 ( .A(out[0]), .B(neg_mul[8]), .Y(n33) );
  NAND2X1 U276 ( .A(out[0]), .B(neg_mul[8]), .Y(n55) );
  NAND2X1 U277 ( .A(neg_mul[10]), .B(n66), .Y(n68) );
  NOR2X1 U278 ( .A(in_8bit[6]), .B(in_8bit[4]), .Y(n191) );
  NOR2XL U279 ( .A(n36), .B(n82), .Y(n83) );
  INVX1 U280 ( .A(in_8bit[4]), .Y(n82) );
  NAND2X1 U281 ( .A(sub_add_75_b0_carry[15]), .B(n9), .Y(n34) );
  NAND2BX1 U282 ( .AN(n33), .B(neg_mul[9]), .Y(n61) );
  AOI211X4 U283 ( .A0(n48), .A1(n65), .B0(n64), .C0(n63), .Y(out[2]) );
  XNOR2X4 U284 ( .A(n75), .B(n4), .Y(out[4]) );
  NOR2X4 U285 ( .A(n26), .B(n78), .Y(n76) );
  XNOR2X4 U286 ( .A(n76), .B(n5), .Y(out[5]) );
  NOR2X4 U287 ( .A(n28), .B(n78), .Y(n79) );
  XNOR2X4 U288 ( .A(n79), .B(n6), .Y(out[7]) );
  MXI2X4 U289 ( .A(n14), .B(n32), .S0(n81), .Y(out[10]) );
  AND2X1 U290 ( .A(add_1_root_r112_carry_20_), .B(n40), .Y(
        add_1_root_r112_SUM_21_) );
  XOR2X1 U291 ( .A(n40), .B(add_1_root_r112_carry_20_), .Y(
        add_1_root_r112_SUM_20_) );
  AND2X1 U292 ( .A(add_1_root_r112_carry_19_), .B(in_17bit_b[15]), .Y(
        add_1_root_r112_carry_20_) );
  XOR2X1 U293 ( .A(in_17bit_b[15]), .B(add_1_root_r112_carry_19_), .Y(
        add_1_root_r112_SUM_19_) );
  AND2X1 U294 ( .A(add_1_root_r112_carry_18_), .B(in_17bit_b[14]), .Y(
        add_1_root_r112_carry_19_) );
  XOR2X1 U295 ( .A(in_17bit_b[14]), .B(add_1_root_r112_carry_18_), .Y(
        add_1_root_r112_SUM_18_) );
  AND2X1 U296 ( .A(add_1_root_r112_carry_17_), .B(in_17bit_b[13]), .Y(
        add_1_root_r112_carry_18_) );
  XOR2X1 U297 ( .A(in_17bit_b[13]), .B(add_1_root_r112_carry_17_), .Y(
        add_1_root_r112_SUM_17_) );
  AND2X1 U298 ( .A(add_2_root_r119_carry_21_), .B(n40), .Y(
        add_2_root_r119_SUM_22_) );
  XOR2X1 U299 ( .A(n40), .B(add_2_root_r119_carry_21_), .Y(
        add_2_root_r119_SUM_21_) );
  AND2X1 U300 ( .A(in_17bit_b[1]), .B(in_17bit_b[0]), .Y(
        add_2_root_r119_carry_6_) );
  XOR2X1 U301 ( .A(in_17bit_b[0]), .B(in_17bit_b[1]), .Y(
        add_2_root_r119_SUM_5_) );
  AND2X1 U302 ( .A(add_1_root_r119_carry[22]), .B(n40), .Y(
        add_1_root_r119_SUM_23_) );
  XOR2X1 U303 ( .A(n40), .B(add_1_root_r119_carry[22]), .Y(
        add_1_root_r119_SUM_22_) );
  AND2X1 U304 ( .A(add_1_root_r119_carry[21]), .B(in_17bit_b[15]), .Y(
        add_1_root_r119_carry[22]) );
  XOR2X1 U305 ( .A(in_17bit_b[15]), .B(add_1_root_r119_carry[21]), .Y(
        add_1_root_r119_SUM_21_) );
  AND2X1 U306 ( .A(add_1_root_r119_carry[20]), .B(in_17bit_b[14]), .Y(
        add_1_root_r119_carry[21]) );
  XOR2X1 U307 ( .A(in_17bit_b[14]), .B(add_1_root_r119_carry[20]), .Y(
        add_1_root_r119_SUM_20_) );
  AND2X1 U308 ( .A(add_1_root_r119_A_6_), .B(in_17bit_b[0]), .Y(
        add_1_root_r119_carry[7]) );
  XOR2X1 U309 ( .A(in_17bit_b[0]), .B(add_1_root_r119_A_6_), .Y(
        add_1_root_r119_SUM_6_) );
  AND2X1 U310 ( .A(add_3_root_r119_carry_18_), .B(n40), .Y(
        add_1_root_r119_A_19_) );
  XOR2X1 U311 ( .A(n40), .B(add_3_root_r119_carry_18_), .Y(
        add_1_root_r119_A_18_) );
  AND2X1 U312 ( .A(in_17bit_b[1]), .B(in_17bit_b[0]), .Y(
        add_3_root_r119_carry_3_) );
  XOR2X1 U313 ( .A(in_17bit_b[0]), .B(in_17bit_b[1]), .Y(add_1_root_r119_A_2_)
         );
  AND2X1 U314 ( .A(add_2_root_r115_carry_19_), .B(n40), .Y(
        add_2_root_r115_SUM_20_) );
  XOR2X1 U315 ( .A(n40), .B(add_2_root_r115_carry_19_), .Y(
        add_2_root_r115_SUM_19_) );
  AND2X1 U316 ( .A(add_2_root_r115_carry_18_), .B(in_17bit_b[15]), .Y(
        add_2_root_r115_carry_19_) );
  XOR2X1 U317 ( .A(in_17bit_b[15]), .B(add_2_root_r115_carry_18_), .Y(
        add_2_root_r115_SUM_18_) );
  AND2X1 U318 ( .A(in_17bit_b[2]), .B(in_17bit_b[0]), .Y(
        add_2_root_r115_carry_4_) );
  XOR2X1 U319 ( .A(in_17bit_b[0]), .B(in_17bit_b[2]), .Y(
        add_2_root_r115_SUM_3_) );
  AND2X1 U320 ( .A(add_1_root_r115_carry_22_), .B(n40), .Y(
        add_1_root_r115_SUM_23_) );
  XOR2X1 U321 ( .A(n40), .B(add_1_root_r115_carry_22_), .Y(
        add_1_root_r115_SUM_22_) );
  AND2X1 U322 ( .A(add_1_root_r115_carry_21_), .B(in_17bit_b[15]), .Y(
        add_1_root_r115_carry_22_) );
  XOR2X1 U323 ( .A(in_17bit_b[15]), .B(add_1_root_r115_carry_21_), .Y(
        add_1_root_r115_SUM_21_) );
  AND2X1 U324 ( .A(in_17bit_b[2]), .B(in_17bit_b[0]), .Y(
        add_1_root_r115_carry_7_) );
  XOR2X1 U325 ( .A(in_17bit_b[0]), .B(in_17bit_b[2]), .Y(
        add_1_root_r115_SUM_6_) );
  XOR2X1 U326 ( .A(n52), .B(sub_add_54_b0_carry[16]), .Y(N29) );
  AND2X1 U327 ( .A(sub_add_54_b0_carry[15]), .B(n168), .Y(
        sub_add_54_b0_carry[16]) );
  XOR2X1 U328 ( .A(n168), .B(sub_add_54_b0_carry[15]), .Y(N28) );
  AND2X1 U329 ( .A(sub_add_54_b0_carry[14]), .B(n164), .Y(
        sub_add_54_b0_carry[15]) );
  XOR2X1 U330 ( .A(n164), .B(sub_add_54_b0_carry[14]), .Y(N27) );
  AND2X1 U331 ( .A(sub_add_54_b0_carry[13]), .B(n163), .Y(
        sub_add_54_b0_carry[14]) );
  XOR2X1 U332 ( .A(n163), .B(sub_add_54_b0_carry[13]), .Y(N26) );
  AND2X1 U333 ( .A(sub_add_54_b0_carry[12]), .B(n162), .Y(
        sub_add_54_b0_carry[13]) );
  XOR2X1 U334 ( .A(n162), .B(sub_add_54_b0_carry[12]), .Y(N25) );
  AND2X1 U335 ( .A(sub_add_54_b0_carry[11]), .B(n161), .Y(
        sub_add_54_b0_carry[12]) );
  XOR2X1 U336 ( .A(n161), .B(sub_add_54_b0_carry[11]), .Y(N24) );
  AND2X1 U337 ( .A(sub_add_54_b0_carry[10]), .B(n160), .Y(
        sub_add_54_b0_carry[11]) );
  XOR2X1 U338 ( .A(n160), .B(sub_add_54_b0_carry[10]), .Y(N23) );
  AND2X1 U339 ( .A(sub_add_54_b0_carry[9]), .B(n158), .Y(
        sub_add_54_b0_carry[10]) );
  XOR2X1 U340 ( .A(n158), .B(sub_add_54_b0_carry[9]), .Y(N22) );
  AND2X1 U341 ( .A(sub_add_54_b0_carry[8]), .B(n101), .Y(
        sub_add_54_b0_carry[9]) );
  XOR2X1 U342 ( .A(n101), .B(sub_add_54_b0_carry[8]), .Y(N21) );
  AND2X1 U343 ( .A(sub_add_54_b0_carry[7]), .B(n100), .Y(
        sub_add_54_b0_carry[8]) );
  XOR2X1 U344 ( .A(n100), .B(sub_add_54_b0_carry[7]), .Y(N20) );
  AND2X1 U345 ( .A(sub_add_54_b0_carry[6]), .B(n99), .Y(sub_add_54_b0_carry[7]) );
  XOR2X1 U346 ( .A(n99), .B(sub_add_54_b0_carry[6]), .Y(N19) );
  AND2X1 U347 ( .A(sub_add_54_b0_carry[5]), .B(n98), .Y(sub_add_54_b0_carry[6]) );
  XOR2X1 U348 ( .A(n98), .B(sub_add_54_b0_carry[5]), .Y(N18) );
  AND2X1 U349 ( .A(sub_add_54_b0_carry[4]), .B(n97), .Y(sub_add_54_b0_carry[5]) );
  XOR2X1 U350 ( .A(n97), .B(sub_add_54_b0_carry[4]), .Y(N17) );
  AND2X1 U351 ( .A(sub_add_54_b0_carry[3]), .B(n96), .Y(sub_add_54_b0_carry[4]) );
  XOR2X1 U352 ( .A(n96), .B(sub_add_54_b0_carry[3]), .Y(N16) );
  AND2X1 U353 ( .A(sub_add_54_b0_carry[2]), .B(n95), .Y(sub_add_54_b0_carry[3]) );
  XOR2X1 U354 ( .A(n95), .B(sub_add_54_b0_carry[2]), .Y(N15) );
  AND2X1 U355 ( .A(n93), .B(n94), .Y(sub_add_54_b0_carry[2]) );
  XOR2X1 U356 ( .A(n94), .B(n93), .Y(N14) );
  XOR2X1 U357 ( .A(n9), .B(sub_add_75_b0_carry[15]), .Y(N480) );
  AND2X1 U358 ( .A(sub_add_75_b0_carry[14]), .B(n10), .Y(
        sub_add_75_b0_carry[15]) );
  XOR2X1 U359 ( .A(n10), .B(sub_add_75_b0_carry[14]), .Y(N479) );
  AND2X1 U360 ( .A(sub_add_75_b0_carry[13]), .B(n11), .Y(
        sub_add_75_b0_carry[14]) );
  XOR2X1 U361 ( .A(n11), .B(sub_add_75_b0_carry[13]), .Y(N478) );
  AND2X1 U362 ( .A(sub_add_75_b0_carry[12]), .B(n12), .Y(
        sub_add_75_b0_carry[13]) );
  XOR2X1 U363 ( .A(n12), .B(sub_add_75_b0_carry[12]), .Y(N477) );
  AND2X1 U364 ( .A(sub_add_75_b0_carry[11]), .B(n13), .Y(
        sub_add_75_b0_carry[12]) );
  XOR2X1 U365 ( .A(n13), .B(sub_add_75_b0_carry[11]), .Y(N476) );
  AND2X1 U366 ( .A(sub_add_75_b0_carry[10]), .B(n14), .Y(
        sub_add_75_b0_carry[11]) );
  AND2X1 U367 ( .A(n31), .B(n7), .Y(sub_add_75_b0_carry[10]) );
  AND2X1 U368 ( .A(in_17bit_b[0]), .B(in_17bit_b[4]), .Y(
        add_1_root_r112_carry_5_) );
endmodule


module multi16_10_DW01_add_0 ( A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, 
        A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, 
        A_4_, B_23_, B_22_, B_21_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, 
        B_14_, B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, 
        SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, 
        SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, 
        SUM_7_ );
  input A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_,
         A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, B_23_, B_22_,
         B_21_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_,
         B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_;
  output SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_,
         SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_,
         SUM_8_, SUM_7_;
  wire   n1, n2, n3, n4;
  wire   [23:7] carry;

  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry[7]), .CO(carry[8]), .S(SUM_7_)
         );
  ADDFX2 U1_21 ( .A(A_21_), .B(B_21_), .CI(carry[21]), .CO(carry[22]), .S(
        SUM_21_) );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry[20]), .CO(carry[21]), .S(
        SUM_20_) );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry[19]), .CO(carry[20]), .S(
        SUM_19_) );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry[18]), .CO(carry[19]), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry[17]), .CO(carry[18]), .S(
        SUM_17_) );
  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry[16]), .CO(carry[17]), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry[15]), .CO(carry[16]), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry[14]), .CO(carry[15]), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry[13]), .CO(carry[14]), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry[12]), .CO(carry[13]), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry[11]), .CO(carry[12]), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry[10]), .CO(carry[11]), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry[9]), .CO(carry[10]), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry[8]), .CO(carry[9]), .S(SUM_8_)
         );
  ADDFX2 U1_22 ( .A(A_22_), .B(B_22_), .CI(carry[22]), .CO(carry[23]), .S(
        SUM_22_) );
  AND2X2 U1 ( .A(A_4_), .B(B_4_), .Y(n1) );
  XOR2X1 U2 ( .A(B_23_), .B(carry[23]), .Y(SUM_23_) );
  OAI2BB1X1 U3 ( .A0N(n2), .A1N(A_6_), .B0(n3), .Y(carry[7]) );
  OAI21XL U4 ( .A0(A_6_), .A1(n2), .B0(B_6_), .Y(n3) );
  OAI2BB1X1 U5 ( .A0N(n1), .A1N(A_5_), .B0(n4), .Y(n2) );
  OAI21XL U6 ( .A0(A_5_), .A1(n1), .B0(B_5_), .Y(n4) );
endmodule


module multi16_10_DW01_add_4 ( A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, 
        A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, 
        B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, 
        B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, SUM_22_, SUM_21_, SUM_20_, 
        SUM_19_, SUM_18_, SUM_17_, SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, 
        SUM_11_, SUM_10_, SUM_9_, SUM_8_, SUM_7_ );
  input A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_,
         A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, B_20_, B_19_,
         B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, B_10_, B_9_,
         B_8_, B_7_, B_6_, B_5_;
  output SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_,
         SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_,
         SUM_7_;
  wire   carry_21_, carry_20_, carry_19_, carry_18_, carry_17_, carry_16_,
         carry_15_, carry_14_, carry_13_, carry_12_, carry_11_, carry_10_,
         carry_9_, carry_8_, carry_7_, n1;

  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry_16_), .CO(carry_17_), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry_15_), .CO(carry_16_), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry_14_), .CO(carry_15_), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry_13_), .CO(carry_14_), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry_12_), .CO(carry_13_), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry_11_), .CO(carry_12_), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry_10_), .CO(carry_11_), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry_9_), .CO(carry_10_), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry_8_), .CO(carry_9_), .S(SUM_8_)
         );
  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry_7_), .CO(carry_8_), .S(SUM_7_)
         );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry_20_), .CO(carry_21_), .S(
        SUM_20_) );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry_19_), .CO(carry_20_), .S(
        SUM_19_) );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry_18_), .CO(carry_19_), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry_17_), .CO(carry_18_), .S(
        SUM_17_) );
  ADDFX2 U1_21 ( .A(A_21_), .B(B_21_), .CI(carry_21_), .CO(SUM_22_), .S(
        SUM_21_) );
  OAI2BB1X1 U1 ( .A0N(A_6_), .A1N(B_6_), .B0(n1), .Y(carry_7_) );
  OAI211X1 U2 ( .A0(B_6_), .A1(A_6_), .B0(A_5_), .C0(B_5_), .Y(n1) );
endmodule


module multi16_10_DW01_add_6 ( A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, 
        A_16_, A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, 
        A_6_, A_5_, A_4_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, 
        B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, 
        SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, 
        SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, 
        SUM_7_ );
  input A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_,
         A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, B_20_,
         B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, B_10_,
         B_9_, B_8_, B_7_, B_6_, B_5_, B_4_;
  output SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_,
         SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_,
         SUM_8_, SUM_7_;
  wire   n1, n2, n3, n4, n5, n6;
  wire   [21:7] carry;

  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry[7]), .CO(carry[8]), .S(SUM_7_)
         );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry[18]), .CO(carry[19]), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry[17]), .CO(carry[18]), .S(
        SUM_17_) );
  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry[16]), .CO(carry[17]), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry[15]), .CO(carry[16]), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry[14]), .CO(carry[15]), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry[13]), .CO(carry[14]), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry[12]), .CO(carry[13]), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry[11]), .CO(carry[12]), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry[10]), .CO(carry[11]), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry[9]), .CO(carry[10]), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry[8]), .CO(carry[9]), .S(SUM_8_)
         );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry[19]), .CO(carry[20]), .S(
        SUM_19_) );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry[20]), .CO(carry[21]), .S(
        SUM_20_) );
  AND2X2 U1 ( .A(A_22_), .B(n2), .Y(n1) );
  AND2X2 U2 ( .A(A_21_), .B(carry[21]), .Y(n2) );
  AND2X2 U3 ( .A(A_4_), .B(B_4_), .Y(n3) );
  XOR2X1 U4 ( .A(A_23_), .B(n1), .Y(SUM_23_) );
  XOR2X1 U5 ( .A(A_21_), .B(carry[21]), .Y(SUM_21_) );
  XOR2X1 U6 ( .A(A_22_), .B(n2), .Y(SUM_22_) );
  OAI2BB1X1 U7 ( .A0N(n4), .A1N(A_6_), .B0(n5), .Y(carry[7]) );
  OAI21XL U8 ( .A0(A_6_), .A1(n4), .B0(B_6_), .Y(n5) );
  OAI2BB1X1 U9 ( .A0N(n3), .A1N(A_5_), .B0(n6), .Y(n4) );
  OAI21XL U10 ( .A0(A_5_), .A1(n3), .B0(B_5_), .Y(n6) );
endmodule


module multi16_10 ( in_17bit, in_8bit, out );
  input [16:0] in_17bit;
  input [7:0] in_8bit;
  output [16:0] out;
  wire   n263, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26,
         N27, N28, N29, N108, N109, N110, N111, N112, N113, N114, N115, N116,
         N117, N118, N119, N120, N121, N122, N123, N205, N206, N207, N208,
         N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, N219,
         N220, N221, N347, N348, N349, N350, N351, N352, N353, N354, N355,
         N356, N357, N358, N359, N360, N361, N362, N363, N446, N447, N448,
         N449, N450, N451, N452, N453, N454, N455, N456, N457, N458, N459,
         N460, N461, N462, N463, N478, N479, N480, add_2_root_r119_carry_10_,
         add_2_root_r119_carry_11_, add_2_root_r119_carry_12_,
         add_2_root_r119_carry_13_, add_2_root_r119_carry_14_,
         add_2_root_r119_carry_15_, add_2_root_r119_carry_16_,
         add_2_root_r119_carry_17_, add_2_root_r119_carry_18_,
         add_2_root_r119_carry_19_, add_2_root_r119_carry_20_,
         add_2_root_r119_carry_21_, add_2_root_r119_carry_6_,
         add_2_root_r119_carry_7_, add_2_root_r119_carry_8_,
         add_2_root_r119_carry_9_, add_2_root_r119_SUM_5_,
         add_2_root_r119_SUM_6_, add_2_root_r119_SUM_7_,
         add_2_root_r119_SUM_8_, add_2_root_r119_SUM_9_,
         add_2_root_r119_SUM_10_, add_2_root_r119_SUM_11_,
         add_2_root_r119_SUM_12_, add_2_root_r119_SUM_13_,
         add_2_root_r119_SUM_14_, add_2_root_r119_SUM_15_,
         add_2_root_r119_SUM_16_, add_2_root_r119_SUM_17_,
         add_2_root_r119_SUM_18_, add_2_root_r119_SUM_19_,
         add_2_root_r119_SUM_20_, add_2_root_r119_SUM_21_,
         add_2_root_r119_SUM_22_, add_1_root_r119_SUM_6_,
         add_1_root_r119_SUM_7_, add_1_root_r119_SUM_8_,
         add_1_root_r119_SUM_9_, add_1_root_r119_SUM_10_,
         add_1_root_r119_SUM_11_, add_1_root_r119_SUM_12_,
         add_1_root_r119_SUM_13_, add_1_root_r119_SUM_14_,
         add_1_root_r119_SUM_15_, add_1_root_r119_SUM_16_,
         add_1_root_r119_SUM_17_, add_1_root_r119_SUM_18_,
         add_1_root_r119_SUM_19_, add_1_root_r119_SUM_20_,
         add_1_root_r119_SUM_21_, add_1_root_r119_SUM_22_,
         add_1_root_r119_SUM_23_, add_1_root_r119_A_2_, add_1_root_r119_A_3_,
         add_1_root_r119_A_4_, add_1_root_r119_A_5_, add_1_root_r119_A_6_,
         add_1_root_r119_A_7_, add_1_root_r119_A_8_, add_1_root_r119_A_9_,
         add_1_root_r119_A_10_, add_1_root_r119_A_11_, add_1_root_r119_A_12_,
         add_1_root_r119_A_13_, add_1_root_r119_A_14_, add_1_root_r119_A_15_,
         add_1_root_r119_A_16_, add_1_root_r119_A_17_, add_1_root_r119_A_18_,
         add_1_root_r119_A_19_, add_3_root_r119_carry_10_,
         add_3_root_r119_carry_11_, add_3_root_r119_carry_12_,
         add_3_root_r119_carry_13_, add_3_root_r119_carry_14_,
         add_3_root_r119_carry_15_, add_3_root_r119_carry_16_,
         add_3_root_r119_carry_17_, add_3_root_r119_carry_18_,
         add_3_root_r119_carry_3_, add_3_root_r119_carry_4_,
         add_3_root_r119_carry_5_, add_3_root_r119_carry_6_,
         add_3_root_r119_carry_7_, add_3_root_r119_carry_8_,
         add_3_root_r119_carry_9_, add_1_root_r112_carry_10_,
         add_1_root_r112_carry_11_, add_1_root_r112_carry_12_,
         add_1_root_r112_carry_13_, add_1_root_r112_carry_14_,
         add_1_root_r112_carry_15_, add_1_root_r112_carry_16_,
         add_1_root_r112_carry_17_, add_1_root_r112_carry_18_,
         add_1_root_r112_carry_19_, add_1_root_r112_carry_20_,
         add_1_root_r112_carry_5_, add_1_root_r112_carry_6_,
         add_1_root_r112_carry_7_, add_1_root_r112_carry_8_,
         add_1_root_r112_carry_9_, add_1_root_r112_SUM_1_,
         add_1_root_r112_SUM_2_, add_1_root_r112_SUM_3_,
         add_1_root_r112_SUM_4_, add_1_root_r112_SUM_5_,
         add_1_root_r112_SUM_6_, add_1_root_r112_SUM_7_,
         add_1_root_r112_SUM_8_, add_1_root_r112_SUM_9_,
         add_1_root_r112_SUM_10_, add_1_root_r112_SUM_11_,
         add_1_root_r112_SUM_12_, add_1_root_r112_SUM_13_,
         add_1_root_r112_SUM_14_, add_1_root_r112_SUM_15_,
         add_1_root_r112_SUM_16_, add_1_root_r112_SUM_17_,
         add_1_root_r112_SUM_18_, add_1_root_r112_SUM_19_,
         add_1_root_r112_SUM_20_, add_1_root_r112_SUM_21_,
         add_2_root_r115_carry_10_, add_2_root_r115_carry_11_,
         add_2_root_r115_carry_12_, add_2_root_r115_carry_13_,
         add_2_root_r115_carry_14_, add_2_root_r115_carry_15_,
         add_2_root_r115_carry_16_, add_2_root_r115_carry_17_,
         add_2_root_r115_carry_18_, add_2_root_r115_carry_19_,
         add_2_root_r115_carry_4_, add_2_root_r115_carry_5_,
         add_2_root_r115_carry_6_, add_2_root_r115_carry_7_,
         add_2_root_r115_carry_8_, add_2_root_r115_carry_9_,
         add_2_root_r115_SUM_3_, add_2_root_r115_SUM_4_,
         add_2_root_r115_SUM_5_, add_2_root_r115_SUM_6_,
         add_2_root_r115_SUM_7_, add_2_root_r115_SUM_8_,
         add_2_root_r115_SUM_9_, add_2_root_r115_SUM_10_,
         add_2_root_r115_SUM_11_, add_2_root_r115_SUM_12_,
         add_2_root_r115_SUM_13_, add_2_root_r115_SUM_14_,
         add_2_root_r115_SUM_15_, add_2_root_r115_SUM_16_,
         add_2_root_r115_SUM_17_, add_2_root_r115_SUM_18_,
         add_2_root_r115_SUM_19_, add_2_root_r115_SUM_20_,
         add_1_root_r115_carry_10_, add_1_root_r115_carry_11_,
         add_1_root_r115_carry_12_, add_1_root_r115_carry_13_,
         add_1_root_r115_carry_14_, add_1_root_r115_carry_15_,
         add_1_root_r115_carry_16_, add_1_root_r115_carry_17_,
         add_1_root_r115_carry_18_, add_1_root_r115_carry_19_,
         add_1_root_r115_carry_20_, add_1_root_r115_carry_21_,
         add_1_root_r115_carry_22_, add_1_root_r115_carry_7_,
         add_1_root_r115_carry_8_, add_1_root_r115_carry_9_,
         add_1_root_r115_SUM_6_, add_1_root_r115_SUM_7_,
         add_1_root_r115_SUM_8_, add_1_root_r115_SUM_9_,
         add_1_root_r115_SUM_10_, add_1_root_r115_SUM_11_,
         add_1_root_r115_SUM_12_, add_1_root_r115_SUM_13_,
         add_1_root_r115_SUM_14_, add_1_root_r115_SUM_15_,
         add_1_root_r115_SUM_16_, add_1_root_r115_SUM_17_,
         add_1_root_r115_SUM_18_, add_1_root_r115_SUM_19_,
         add_1_root_r115_SUM_20_, add_1_root_r115_SUM_21_,
         add_1_root_r115_SUM_22_, add_1_root_r115_SUM_23_, n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n158, n160, n161, n162,
         n163, n164, n168, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262;
  wire   [16:0] in_17bit_b;
  wire   [23:8] neg_mul;
  wire   [15:11] sub_add_75_b0_carry;
  wire   [15:2] sub_add_54_b0_carry;
  wire   [22:7] add_1_root_r119_carry;

  multi16_10_DW01_add_0 add_0_root_r119 ( .A_22_(add_2_root_r119_SUM_22_), 
        .A_21_(add_2_root_r119_SUM_21_), .A_20_(add_2_root_r119_SUM_20_), 
        .A_19_(add_2_root_r119_SUM_19_), .A_18_(add_2_root_r119_SUM_18_), 
        .A_17_(add_2_root_r119_SUM_17_), .A_16_(add_2_root_r119_SUM_16_), 
        .A_15_(add_2_root_r119_SUM_15_), .A_14_(add_2_root_r119_SUM_14_), 
        .A_13_(add_2_root_r119_SUM_13_), .A_12_(add_2_root_r119_SUM_12_), 
        .A_11_(add_2_root_r119_SUM_11_), .A_10_(add_2_root_r119_SUM_10_), 
        .A_9_(add_2_root_r119_SUM_9_), .A_8_(add_2_root_r119_SUM_8_), .A_7_(
        add_2_root_r119_SUM_7_), .A_6_(add_2_root_r119_SUM_6_), .A_5_(
        add_2_root_r119_SUM_5_), .A_4_(in_17bit_b[0]), .B_23_(
        add_1_root_r119_SUM_23_), .B_22_(add_1_root_r119_SUM_22_), .B_21_(
        add_1_root_r119_SUM_21_), .B_20_(add_1_root_r119_SUM_20_), .B_19_(
        add_1_root_r119_SUM_19_), .B_18_(add_1_root_r119_SUM_18_), .B_17_(
        add_1_root_r119_SUM_17_), .B_16_(add_1_root_r119_SUM_16_), .B_15_(
        add_1_root_r119_SUM_15_), .B_14_(add_1_root_r119_SUM_14_), .B_13_(
        add_1_root_r119_SUM_13_), .B_12_(add_1_root_r119_SUM_12_), .B_11_(
        add_1_root_r119_SUM_11_), .B_10_(add_1_root_r119_SUM_10_), .B_9_(
        add_1_root_r119_SUM_9_), .B_8_(add_1_root_r119_SUM_8_), .B_7_(
        add_1_root_r119_SUM_7_), .B_6_(add_1_root_r119_SUM_6_), .B_5_(
        add_1_root_r119_A_5_), .B_4_(add_1_root_r119_A_4_), .SUM_23_(N363), 
        .SUM_22_(N362), .SUM_21_(N361), .SUM_20_(N360), .SUM_19_(N359), 
        .SUM_18_(N358), .SUM_17_(N357), .SUM_16_(N356), .SUM_15_(N355), 
        .SUM_14_(N354), .SUM_13_(N353), .SUM_12_(N352), .SUM_11_(N351), 
        .SUM_10_(N350), .SUM_9_(N349), .SUM_8_(N348), .SUM_7_(N347) );
  multi16_10_DW01_add_4 add_0_root_r112 ( .A_21_(n42), .A_20_(in_17bit_b[15]), 
        .A_19_(in_17bit_b[14]), .A_18_(in_17bit_b[13]), .A_17_(in_17bit_b[12]), 
        .A_16_(in_17bit_b[11]), .A_15_(in_17bit_b[10]), .A_14_(in_17bit_b[9]), 
        .A_13_(in_17bit_b[8]), .A_12_(in_17bit_b[7]), .A_11_(in_17bit_b[6]), 
        .A_10_(in_17bit_b[5]), .A_9_(in_17bit_b[4]), .A_8_(in_17bit_b[3]), 
        .A_7_(in_17bit_b[2]), .A_6_(in_17bit_b[1]), .A_5_(in_17bit_b[0]), 
        .B_21_(add_1_root_r112_SUM_21_), .B_20_(add_1_root_r112_SUM_20_), 
        .B_19_(add_1_root_r112_SUM_19_), .B_18_(add_1_root_r112_SUM_18_), 
        .B_17_(add_1_root_r112_SUM_17_), .B_16_(add_1_root_r112_SUM_16_), 
        .B_15_(add_1_root_r112_SUM_15_), .B_14_(add_1_root_r112_SUM_14_), 
        .B_13_(add_1_root_r112_SUM_13_), .B_12_(add_1_root_r112_SUM_12_), 
        .B_11_(add_1_root_r112_SUM_11_), .B_10_(add_1_root_r112_SUM_10_), 
        .B_9_(add_1_root_r112_SUM_9_), .B_8_(add_1_root_r112_SUM_8_), .B_7_(
        add_1_root_r112_SUM_7_), .B_6_(add_1_root_r112_SUM_6_), .B_5_(
        add_1_root_r112_SUM_5_), .SUM_22_(N123), .SUM_21_(N122), .SUM_20_(N121), .SUM_19_(N120), .SUM_18_(N119), .SUM_17_(N118), .SUM_16_(N117), .SUM_15_(
        N116), .SUM_14_(N115), .SUM_13_(N114), .SUM_12_(N113), .SUM_11_(N112), 
        .SUM_10_(N111), .SUM_9_(N110), .SUM_8_(N109), .SUM_7_(N108) );
  multi16_10_DW01_add_6 add_0_root_r115 ( .A_23_(add_1_root_r115_SUM_23_), 
        .A_22_(add_1_root_r115_SUM_22_), .A_21_(add_1_root_r115_SUM_21_), 
        .A_20_(add_1_root_r115_SUM_20_), .A_19_(add_1_root_r115_SUM_19_), 
        .A_18_(add_1_root_r115_SUM_18_), .A_17_(add_1_root_r115_SUM_17_), 
        .A_16_(add_1_root_r115_SUM_16_), .A_15_(add_1_root_r115_SUM_15_), 
        .A_14_(add_1_root_r115_SUM_14_), .A_13_(add_1_root_r115_SUM_13_), 
        .A_12_(add_1_root_r115_SUM_12_), .A_11_(add_1_root_r115_SUM_11_), 
        .A_10_(add_1_root_r115_SUM_10_), .A_9_(add_1_root_r115_SUM_9_), .A_8_(
        add_1_root_r115_SUM_8_), .A_7_(add_1_root_r115_SUM_7_), .A_6_(
        add_1_root_r115_SUM_6_), .A_5_(in_17bit_b[1]), .A_4_(in_17bit_b[0]), 
        .B_20_(add_2_root_r115_SUM_20_), .B_19_(add_2_root_r115_SUM_19_), 
        .B_18_(add_2_root_r115_SUM_18_), .B_17_(add_2_root_r115_SUM_17_), 
        .B_16_(add_2_root_r115_SUM_16_), .B_15_(add_2_root_r115_SUM_15_), 
        .B_14_(add_2_root_r115_SUM_14_), .B_13_(add_2_root_r115_SUM_13_), 
        .B_12_(add_2_root_r115_SUM_12_), .B_11_(add_2_root_r115_SUM_11_), 
        .B_10_(add_2_root_r115_SUM_10_), .B_9_(add_2_root_r115_SUM_9_), .B_8_(
        add_2_root_r115_SUM_8_), .B_7_(add_2_root_r115_SUM_7_), .B_6_(
        add_2_root_r115_SUM_6_), .B_5_(add_2_root_r115_SUM_5_), .B_4_(
        add_2_root_r115_SUM_4_), .SUM_23_(N221), .SUM_22_(N220), .SUM_21_(N219), .SUM_20_(N218), .SUM_19_(N217), .SUM_18_(N216), .SUM_17_(N215), .SUM_16_(
        N214), .SUM_15_(N213), .SUM_14_(N212), .SUM_13_(N211), .SUM_12_(N210), 
        .SUM_11_(N209), .SUM_10_(N208), .SUM_9_(N207), .SUM_8_(N206), .SUM_7_(
        N205) );
  TLATX1 neg_mul_reg_17_ ( .G(N446), .D(N457), .QN(n8) );
  TLATX1 neg_mul_reg_16_ ( .G(N446), .D(N456), .QN(n7) );
  TLATX1 neg_mul_reg_15_ ( .G(N446), .D(N455), .QN(n6) );
  TLATX1 neg_mul_reg_14_ ( .G(N446), .D(N454), .QN(n5) );
  TLATX1 neg_mul_reg_13_ ( .G(N446), .D(N453), .QN(n4) );
  TLATX1 neg_mul_reg_12_ ( .G(N446), .D(N452), .QN(n3) );
  TLATX1 neg_mul_reg_11_ ( .G(N446), .D(N451), .Q(n1), .QN(n16) );
  TLATX1 neg_mul_reg_23_ ( .G(N446), .D(N463), .Q(neg_mul[23]), .QN(n2) );
  TLATX1 neg_mul_reg_22_ ( .G(N446), .D(N462), .Q(neg_mul[22]), .QN(n10) );
  TLATX1 neg_mul_reg_21_ ( .G(N446), .D(N461), .Q(neg_mul[21]), .QN(n13) );
  TLATX1 neg_mul_reg_20_ ( .G(N446), .D(N460), .Q(neg_mul[20]), .QN(n11) );
  TLATX1 neg_mul_reg_19_ ( .G(N446), .D(N459), .QN(n17) );
  TLATX1 neg_mul_reg_18_ ( .G(N446), .D(N458), .QN(n12) );
  TLATX1 neg_mul_reg_9_ ( .G(N446), .D(N449), .Q(neg_mul[9]), .QN(n9) );
  TLATX1 neg_mul_reg_10_ ( .G(N446), .D(N450), .Q(neg_mul[10]), .QN(n14) );
  TLATX1 neg_mul_reg_8_ ( .G(N446), .D(N448), .Q(neg_mul[8]), .QN(n15) );
  TLATX1 neg_mul_reg_7_ ( .G(N446), .D(N447), .Q(out[0]) );
  NOR2X2 U2 ( .A(n57), .B(n70), .Y(n72) );
  XNOR2X4 U3 ( .A(n57), .B(n43), .Y(n81) );
  XNOR2X2 U4 ( .A(n57), .B(n43), .Y(n83) );
  XNOR2X2 U5 ( .A(n57), .B(n43), .Y(n86) );
  INVX2 U6 ( .A(in_17bit[16]), .Y(n55) );
  NOR2BX2 U7 ( .AN(n59), .B(n78), .Y(n79) );
  INVX4 U8 ( .A(n53), .Y(n59) );
  AOI2BB2X1 U9 ( .B0(n63), .B1(n43), .A0N(n44), .A1N(neg_mul[8]), .Y(n64) );
  INVX12 U10 ( .A(n45), .Y(n44) );
  CLKINVX20 U11 ( .A(n45), .Y(n43) );
  XNOR2X2 U12 ( .A(n57), .B(n43), .Y(n88) );
  AOI2BB2X1 U13 ( .B0(n77), .B1(n43), .A0N(n44), .A1N(neg_mul[10]), .Y(n78) );
  OAI21XL U14 ( .A0(n43), .A1(n62), .B0(n61), .Y(n66) );
  NAND2X2 U15 ( .A(n43), .B(n15), .Y(n61) );
  AOI2BB2X1 U16 ( .B0(n69), .B1(n43), .A0N(n44), .A1N(neg_mul[9]), .Y(n70) );
  NAND2X1 U17 ( .A(n44), .B(n9), .Y(n67) );
  MXI2X2 U18 ( .A(n12), .B(n18), .S0(n27), .Y(out[11]) );
  NOR2X2 U19 ( .A(n92), .B(n35), .Y(n91) );
  MXI2X1 U20 ( .A(n17), .B(n36), .S0(n27), .Y(out[12]) );
  MX2X1 U21 ( .A(neg_mul[20]), .B(N478), .S0(n27), .Y(out[13]) );
  CLKINVX3 U22 ( .A(n54), .Y(n53) );
  INVX4 U23 ( .A(in_8bit[7]), .Y(n45) );
  INVX1 U24 ( .A(n101), .Y(n97) );
  INVX4 U25 ( .A(in_17bit[16]), .Y(n22) );
  INVX1 U26 ( .A(n55), .Y(n51) );
  INVX1 U27 ( .A(in_17bit[16]), .Y(n54) );
  INVX1 U28 ( .A(n55), .Y(n52) );
  XNOR2X2 U29 ( .A(n57), .B(n43), .Y(n92) );
  XNOR2X1 U30 ( .A(n12), .B(sub_add_75_b0_carry[11]), .Y(n18) );
  XNOR2X1 U31 ( .A(neg_mul[23]), .B(n38), .Y(n19) );
  CLKINVX8 U32 ( .A(n20), .Y(out[1]) );
  INVX8 U33 ( .A(n22), .Y(n57) );
  INVX4 U34 ( .A(n263), .Y(n20) );
  AOI211X2 U35 ( .A0(n51), .A1(n66), .B0(n65), .C0(n37), .Y(n263) );
  XOR2X4 U36 ( .A(n57), .B(n43), .Y(n27) );
  NOR2X2 U37 ( .A(n57), .B(n64), .Y(n65) );
  NOR2X2 U38 ( .A(n92), .B(n33), .Y(n90) );
  OAI21XL U39 ( .A0(n43), .A1(n68), .B0(n67), .Y(n73) );
  NOR2X4 U40 ( .A(n82), .B(n81), .Y(n23) );
  INVX1 U41 ( .A(n212), .Y(in_17bit_b[1]) );
  INVX1 U42 ( .A(n251), .Y(in_17bit_b[14]) );
  INVX1 U43 ( .A(n248), .Y(in_17bit_b[13]) );
  INVX1 U44 ( .A(n215), .Y(in_17bit_b[2]) );
  INVX1 U45 ( .A(n224), .Y(in_17bit_b[5]) );
  INVX1 U46 ( .A(n227), .Y(in_17bit_b[6]) );
  INVX1 U47 ( .A(n230), .Y(in_17bit_b[7]) );
  INVX1 U48 ( .A(n233), .Y(in_17bit_b[8]) );
  INVX1 U49 ( .A(n236), .Y(in_17bit_b[9]) );
  INVX1 U50 ( .A(n239), .Y(in_17bit_b[10]) );
  INVX1 U51 ( .A(n242), .Y(in_17bit_b[11]) );
  INVX1 U52 ( .A(n245), .Y(in_17bit_b[12]) );
  INVX1 U53 ( .A(n221), .Y(in_17bit_b[4]) );
  INVX1 U54 ( .A(n218), .Y(in_17bit_b[3]) );
  XOR2X4 U55 ( .A(n23), .B(n1), .Y(out[4]) );
  NAND2XL U56 ( .A(n44), .B(n14), .Y(n75) );
  AOI21X1 U57 ( .A0(n24), .A1(n25), .B0(n255), .Y(n208) );
  NOR4XL U58 ( .A(in_8bit[4]), .B(in_8bit[5]), .C(in_8bit[6]), .D(n43), .Y(n24) );
  NOR4X1 U59 ( .A(in_8bit[1]), .B(in_8bit[0]), .C(n49), .D(in_8bit[3]), .Y(n25) );
  AND4X1 U60 ( .A(in_8bit[1]), .B(in_8bit[7]), .C(n202), .D(n46), .Y(n26) );
  INVX1 U61 ( .A(n50), .Y(n49) );
  INVX1 U62 ( .A(in_8bit[2]), .Y(n50) );
  INVX1 U63 ( .A(in_8bit[6]), .Y(n47) );
  NOR3X1 U64 ( .A(n50), .B(n48), .C(n46), .Y(n207) );
  NOR4BX1 U65 ( .AN(n205), .B(n46), .C(in_8bit[1]), .D(n49), .Y(n206) );
  NOR2X1 U66 ( .A(in_8bit[6]), .B(in_8bit[3]), .Y(n205) );
  NAND3X1 U67 ( .A(n49), .B(n48), .C(in_8bit[5]), .Y(n203) );
  ADDFX2 U68 ( .A(n42), .B(in_17bit_b[12]), .CI(add_1_root_r112_carry_16_), 
        .CO(add_1_root_r112_carry_17_), .S(add_1_root_r112_SUM_16_) );
  ADDFX2 U69 ( .A(add_1_root_r119_A_19_), .B(in_17bit_b[13]), .CI(
        add_1_root_r119_carry[19]), .CO(add_1_root_r119_carry[20]), .S(
        add_1_root_r119_SUM_19_) );
  ADDFX2 U70 ( .A(n42), .B(in_17bit_b[15]), .CI(add_3_root_r119_carry_17_), 
        .CO(add_3_root_r119_carry_18_), .S(add_1_root_r119_A_17_) );
  ADDFX2 U71 ( .A(n42), .B(in_17bit_b[14]), .CI(add_2_root_r115_carry_17_), 
        .CO(add_2_root_r115_carry_18_), .S(add_2_root_r115_SUM_17_) );
  ADDFX2 U72 ( .A(n42), .B(in_17bit_b[14]), .CI(add_1_root_r115_carry_20_), 
        .CO(add_1_root_r115_carry_21_), .S(add_1_root_r115_SUM_20_) );
  ADDFX2 U73 ( .A(n42), .B(in_17bit_b[15]), .CI(add_2_root_r119_carry_20_), 
        .CO(add_2_root_r119_carry_21_), .S(add_2_root_r119_SUM_20_) );
  INVX1 U74 ( .A(n59), .Y(n56) );
  ADDFX2 U75 ( .A(in_17bit_b[3]), .B(in_17bit_b[1]), .CI(
        add_2_root_r115_carry_4_), .CO(add_2_root_r115_carry_5_), .S(
        add_2_root_r115_SUM_4_) );
  ADDFX2 U76 ( .A(in_17bit_b[4]), .B(in_17bit_b[2]), .CI(
        add_2_root_r115_carry_5_), .CO(add_2_root_r115_carry_6_), .S(
        add_2_root_r115_SUM_5_) );
  ADDFX2 U77 ( .A(in_17bit_b[5]), .B(in_17bit_b[1]), .CI(
        add_1_root_r112_carry_5_), .CO(add_1_root_r112_carry_6_), .S(
        add_1_root_r112_SUM_5_) );
  ADDFX2 U78 ( .A(in_17bit_b[6]), .B(in_17bit_b[5]), .CI(
        add_3_root_r119_carry_7_), .CO(add_3_root_r119_carry_8_), .S(
        add_1_root_r119_A_7_) );
  ADDFX2 U79 ( .A(in_17bit_b[6]), .B(in_17bit_b[2]), .CI(
        add_1_root_r112_carry_6_), .CO(add_1_root_r112_carry_7_), .S(
        add_1_root_r112_SUM_6_) );
  ADDFX2 U80 ( .A(in_17bit_b[3]), .B(in_17bit_b[1]), .CI(
        add_1_root_r115_carry_7_), .CO(add_1_root_r115_carry_8_), .S(
        add_1_root_r115_SUM_7_) );
  ADDFX2 U81 ( .A(in_17bit_b[7]), .B(in_17bit_b[6]), .CI(
        add_3_root_r119_carry_8_), .CO(add_3_root_r119_carry_9_), .S(
        add_1_root_r119_A_8_) );
  ADDFX2 U82 ( .A(add_1_root_r119_A_7_), .B(in_17bit_b[1]), .CI(
        add_1_root_r119_carry[7]), .CO(add_1_root_r119_carry[8]), .S(
        add_1_root_r119_SUM_7_) );
  ADDFX2 U83 ( .A(in_17bit_b[2]), .B(in_17bit_b[1]), .CI(
        add_2_root_r119_carry_6_), .CO(add_2_root_r119_carry_7_), .S(
        add_2_root_r119_SUM_6_) );
  ADDFX2 U84 ( .A(in_17bit_b[4]), .B(in_17bit_b[2]), .CI(
        add_1_root_r115_carry_8_), .CO(add_1_root_r115_carry_9_), .S(
        add_1_root_r115_SUM_8_) );
  ADDFX2 U85 ( .A(in_17bit_b[8]), .B(in_17bit_b[7]), .CI(
        add_3_root_r119_carry_9_), .CO(add_3_root_r119_carry_10_), .S(
        add_1_root_r119_A_9_) );
  ADDFX2 U86 ( .A(add_1_root_r119_A_8_), .B(in_17bit_b[2]), .CI(
        add_1_root_r119_carry[8]), .CO(add_1_root_r119_carry[9]), .S(
        add_1_root_r119_SUM_8_) );
  ADDFX2 U87 ( .A(in_17bit_b[3]), .B(in_17bit_b[2]), .CI(
        add_2_root_r119_carry_7_), .CO(add_2_root_r119_carry_8_), .S(
        add_2_root_r119_SUM_7_) );
  ADDFX2 U88 ( .A(in_17bit_b[6]), .B(in_17bit_b[4]), .CI(
        add_2_root_r115_carry_7_), .CO(add_2_root_r115_carry_8_), .S(
        add_2_root_r115_SUM_7_) );
  ADDFX2 U89 ( .A(in_17bit_b[8]), .B(in_17bit_b[4]), .CI(
        add_1_root_r112_carry_8_), .CO(add_1_root_r112_carry_9_), .S(
        add_1_root_r112_SUM_8_) );
  ADDFX2 U90 ( .A(in_17bit_b[9]), .B(in_17bit_b[8]), .CI(
        add_3_root_r119_carry_10_), .CO(add_3_root_r119_carry_11_), .S(
        add_1_root_r119_A_10_) );
  ADDFX2 U91 ( .A(in_17bit_b[7]), .B(in_17bit_b[5]), .CI(
        add_2_root_r115_carry_8_), .CO(add_2_root_r115_carry_9_), .S(
        add_2_root_r115_SUM_8_) );
  ADDFX2 U92 ( .A(in_17bit_b[9]), .B(in_17bit_b[5]), .CI(
        add_1_root_r112_carry_9_), .CO(add_1_root_r112_carry_10_), .S(
        add_1_root_r112_SUM_9_) );
  ADDFX2 U93 ( .A(in_17bit_b[6]), .B(in_17bit_b[4]), .CI(
        add_1_root_r115_carry_10_), .CO(add_1_root_r115_carry_11_), .S(
        add_1_root_r115_SUM_10_) );
  ADDFX2 U94 ( .A(in_17bit_b[10]), .B(in_17bit_b[9]), .CI(
        add_3_root_r119_carry_11_), .CO(add_3_root_r119_carry_12_), .S(
        add_1_root_r119_A_11_) );
  ADDFX2 U95 ( .A(add_1_root_r119_A_9_), .B(in_17bit_b[3]), .CI(
        add_1_root_r119_carry[9]), .CO(add_1_root_r119_carry[10]), .S(
        add_1_root_r119_SUM_9_) );
  ADDFX2 U96 ( .A(in_17bit_b[5]), .B(in_17bit_b[4]), .CI(
        add_2_root_r119_carry_9_), .CO(add_2_root_r119_carry_10_), .S(
        add_2_root_r119_SUM_9_) );
  ADDFX2 U97 ( .A(in_17bit_b[8]), .B(in_17bit_b[6]), .CI(
        add_2_root_r115_carry_9_), .CO(add_2_root_r115_carry_10_), .S(
        add_2_root_r115_SUM_9_) );
  ADDFX2 U98 ( .A(in_17bit_b[10]), .B(in_17bit_b[6]), .CI(
        add_1_root_r112_carry_10_), .CO(add_1_root_r112_carry_11_), .S(
        add_1_root_r112_SUM_10_) );
  ADDFX2 U99 ( .A(in_17bit_b[7]), .B(in_17bit_b[5]), .CI(
        add_1_root_r115_carry_11_), .CO(add_1_root_r115_carry_12_), .S(
        add_1_root_r115_SUM_11_) );
  ADDFX2 U100 ( .A(in_17bit_b[11]), .B(in_17bit_b[10]), .CI(
        add_3_root_r119_carry_12_), .CO(add_3_root_r119_carry_13_), .S(
        add_1_root_r119_A_12_) );
  ADDFX2 U101 ( .A(add_1_root_r119_A_11_), .B(in_17bit_b[5]), .CI(
        add_1_root_r119_carry[11]), .CO(add_1_root_r119_carry[12]), .S(
        add_1_root_r119_SUM_11_) );
  ADDFX2 U102 ( .A(in_17bit_b[6]), .B(in_17bit_b[5]), .CI(
        add_2_root_r119_carry_10_), .CO(add_2_root_r119_carry_11_), .S(
        add_2_root_r119_SUM_10_) );
  ADDFX2 U103 ( .A(in_17bit_b[9]), .B(in_17bit_b[7]), .CI(
        add_2_root_r115_carry_10_), .CO(add_2_root_r115_carry_11_), .S(
        add_2_root_r115_SUM_10_) );
  ADDFX2 U104 ( .A(in_17bit_b[8]), .B(in_17bit_b[6]), .CI(
        add_1_root_r115_carry_12_), .CO(add_1_root_r115_carry_13_), .S(
        add_1_root_r115_SUM_12_) );
  ADDFX2 U105 ( .A(in_17bit_b[12]), .B(in_17bit_b[11]), .CI(
        add_3_root_r119_carry_13_), .CO(add_3_root_r119_carry_14_), .S(
        add_1_root_r119_A_13_) );
  ADDFX2 U106 ( .A(add_1_root_r119_A_12_), .B(in_17bit_b[6]), .CI(
        add_1_root_r119_carry[12]), .CO(add_1_root_r119_carry[13]), .S(
        add_1_root_r119_SUM_12_) );
  ADDFX2 U107 ( .A(in_17bit_b[7]), .B(in_17bit_b[6]), .CI(
        add_2_root_r119_carry_11_), .CO(add_2_root_r119_carry_12_), .S(
        add_2_root_r119_SUM_11_) );
  ADDFX2 U108 ( .A(in_17bit_b[10]), .B(in_17bit_b[8]), .CI(
        add_2_root_r115_carry_11_), .CO(add_2_root_r115_carry_12_), .S(
        add_2_root_r115_SUM_11_) );
  ADDFX2 U109 ( .A(in_17bit_b[12]), .B(in_17bit_b[8]), .CI(
        add_1_root_r112_carry_12_), .CO(add_1_root_r112_carry_13_), .S(
        add_1_root_r112_SUM_12_) );
  ADDFX2 U110 ( .A(in_17bit_b[9]), .B(in_17bit_b[7]), .CI(
        add_1_root_r115_carry_13_), .CO(add_1_root_r115_carry_14_), .S(
        add_1_root_r115_SUM_13_) );
  ADDFX2 U111 ( .A(in_17bit_b[13]), .B(in_17bit_b[12]), .CI(
        add_3_root_r119_carry_14_), .CO(add_3_root_r119_carry_15_), .S(
        add_1_root_r119_A_14_) );
  ADDFX2 U112 ( .A(add_1_root_r119_A_13_), .B(in_17bit_b[7]), .CI(
        add_1_root_r119_carry[13]), .CO(add_1_root_r119_carry[14]), .S(
        add_1_root_r119_SUM_13_) );
  ADDFX2 U113 ( .A(in_17bit_b[8]), .B(in_17bit_b[7]), .CI(
        add_2_root_r119_carry_12_), .CO(add_2_root_r119_carry_13_), .S(
        add_2_root_r119_SUM_12_) );
  ADDFX2 U114 ( .A(in_17bit_b[11]), .B(in_17bit_b[9]), .CI(
        add_2_root_r115_carry_12_), .CO(add_2_root_r115_carry_13_), .S(
        add_2_root_r115_SUM_12_) );
  ADDFX2 U115 ( .A(in_17bit_b[13]), .B(in_17bit_b[9]), .CI(
        add_1_root_r112_carry_13_), .CO(add_1_root_r112_carry_14_), .S(
        add_1_root_r112_SUM_13_) );
  ADDFX2 U116 ( .A(in_17bit_b[10]), .B(in_17bit_b[8]), .CI(
        add_1_root_r115_carry_14_), .CO(add_1_root_r115_carry_15_), .S(
        add_1_root_r115_SUM_14_) );
  ADDFX2 U117 ( .A(in_17bit_b[14]), .B(in_17bit_b[13]), .CI(
        add_3_root_r119_carry_15_), .CO(add_3_root_r119_carry_16_), .S(
        add_1_root_r119_A_15_) );
  ADDFX2 U118 ( .A(add_1_root_r119_A_14_), .B(in_17bit_b[8]), .CI(
        add_1_root_r119_carry[14]), .CO(add_1_root_r119_carry[15]), .S(
        add_1_root_r119_SUM_14_) );
  ADDFX2 U119 ( .A(in_17bit_b[3]), .B(in_17bit_b[2]), .CI(
        add_3_root_r119_carry_4_), .CO(add_3_root_r119_carry_5_), .S(
        add_1_root_r119_A_4_) );
  ADDFX2 U120 ( .A(in_17bit_b[2]), .B(in_17bit_b[1]), .CI(
        add_3_root_r119_carry_3_), .CO(add_3_root_r119_carry_4_), .S(
        add_1_root_r119_A_3_) );
  ADDFX2 U121 ( .A(in_17bit_b[9]), .B(in_17bit_b[8]), .CI(
        add_2_root_r119_carry_13_), .CO(add_2_root_r119_carry_14_), .S(
        add_2_root_r119_SUM_13_) );
  ADDFX2 U122 ( .A(in_17bit_b[12]), .B(in_17bit_b[10]), .CI(
        add_2_root_r115_carry_13_), .CO(add_2_root_r115_carry_14_), .S(
        add_2_root_r115_SUM_13_) );
  ADDFX2 U123 ( .A(in_17bit_b[14]), .B(in_17bit_b[10]), .CI(
        add_1_root_r112_carry_14_), .CO(add_1_root_r112_carry_15_), .S(
        add_1_root_r112_SUM_14_) );
  ADDFX2 U124 ( .A(in_17bit_b[11]), .B(in_17bit_b[9]), .CI(
        add_1_root_r115_carry_15_), .CO(add_1_root_r115_carry_16_), .S(
        add_1_root_r115_SUM_15_) );
  ADDFX2 U125 ( .A(add_1_root_r119_A_15_), .B(in_17bit_b[9]), .CI(
        add_1_root_r119_carry[15]), .CO(add_1_root_r119_carry[16]), .S(
        add_1_root_r119_SUM_15_) );
  ADDFX2 U126 ( .A(in_17bit_b[10]), .B(in_17bit_b[9]), .CI(
        add_2_root_r119_carry_14_), .CO(add_2_root_r119_carry_15_), .S(
        add_2_root_r119_SUM_14_) );
  ADDFX2 U127 ( .A(in_17bit_b[13]), .B(in_17bit_b[11]), .CI(
        add_2_root_r115_carry_14_), .CO(add_2_root_r115_carry_15_), .S(
        add_2_root_r115_SUM_14_) );
  ADDFX2 U128 ( .A(in_17bit_b[15]), .B(in_17bit_b[11]), .CI(
        add_1_root_r112_carry_15_), .CO(add_1_root_r112_carry_16_), .S(
        add_1_root_r112_SUM_15_) );
  ADDFX2 U129 ( .A(in_17bit_b[12]), .B(in_17bit_b[10]), .CI(
        add_1_root_r115_carry_16_), .CO(add_1_root_r115_carry_17_), .S(
        add_1_root_r115_SUM_16_) );
  ADDFX2 U130 ( .A(add_1_root_r119_A_16_), .B(in_17bit_b[10]), .CI(
        add_1_root_r119_carry[16]), .CO(add_1_root_r119_carry[17]), .S(
        add_1_root_r119_SUM_16_) );
  ADDFX2 U131 ( .A(in_17bit_b[11]), .B(in_17bit_b[10]), .CI(
        add_2_root_r119_carry_15_), .CO(add_2_root_r119_carry_16_), .S(
        add_2_root_r119_SUM_15_) );
  ADDFX2 U132 ( .A(in_17bit_b[14]), .B(in_17bit_b[12]), .CI(
        add_2_root_r115_carry_15_), .CO(add_2_root_r115_carry_16_), .S(
        add_2_root_r115_SUM_15_) );
  ADDFX2 U133 ( .A(in_17bit_b[13]), .B(in_17bit_b[11]), .CI(
        add_1_root_r115_carry_17_), .CO(add_1_root_r115_carry_18_), .S(
        add_1_root_r115_SUM_17_) );
  ADDFX2 U134 ( .A(add_1_root_r119_A_17_), .B(in_17bit_b[11]), .CI(
        add_1_root_r119_carry[17]), .CO(add_1_root_r119_carry[18]), .S(
        add_1_root_r119_SUM_17_) );
  ADDFX2 U135 ( .A(in_17bit_b[5]), .B(in_17bit_b[4]), .CI(
        add_3_root_r119_carry_6_), .CO(add_3_root_r119_carry_7_), .S(
        add_1_root_r119_A_6_) );
  ADDFX2 U136 ( .A(in_17bit_b[12]), .B(in_17bit_b[11]), .CI(
        add_2_root_r119_carry_16_), .CO(add_2_root_r119_carry_17_), .S(
        add_2_root_r119_SUM_16_) );
  ADDFX2 U137 ( .A(in_17bit_b[15]), .B(in_17bit_b[13]), .CI(
        add_2_root_r115_carry_16_), .CO(add_2_root_r115_carry_17_), .S(
        add_2_root_r115_SUM_16_) );
  ADDFX2 U138 ( .A(in_17bit_b[14]), .B(in_17bit_b[12]), .CI(
        add_1_root_r115_carry_18_), .CO(add_1_root_r115_carry_19_), .S(
        add_1_root_r115_SUM_18_) );
  ADDFX2 U139 ( .A(add_1_root_r119_A_18_), .B(in_17bit_b[12]), .CI(
        add_1_root_r119_carry[18]), .CO(add_1_root_r119_carry[19]), .S(
        add_1_root_r119_SUM_18_) );
  ADDFX2 U140 ( .A(in_17bit_b[13]), .B(in_17bit_b[12]), .CI(
        add_2_root_r119_carry_17_), .CO(add_2_root_r119_carry_18_), .S(
        add_2_root_r119_SUM_17_) );
  ADDFX2 U141 ( .A(in_17bit_b[5]), .B(in_17bit_b[3]), .CI(
        add_2_root_r115_carry_6_), .CO(add_2_root_r115_carry_7_), .S(
        add_2_root_r115_SUM_6_) );
  ADDFX2 U142 ( .A(in_17bit_b[5]), .B(in_17bit_b[3]), .CI(
        add_1_root_r115_carry_9_), .CO(add_1_root_r115_carry_10_), .S(
        add_1_root_r115_SUM_9_) );
  ADDFX2 U143 ( .A(add_1_root_r119_A_10_), .B(in_17bit_b[4]), .CI(
        add_1_root_r119_carry[10]), .CO(add_1_root_r119_carry[11]), .S(
        add_1_root_r119_SUM_10_) );
  ADDFX2 U144 ( .A(in_17bit_b[11]), .B(in_17bit_b[7]), .CI(
        add_1_root_r112_carry_11_), .CO(add_1_root_r112_carry_12_), .S(
        add_1_root_r112_SUM_11_) );
  ADDFX2 U145 ( .A(in_17bit_b[15]), .B(in_17bit_b[14]), .CI(
        add_3_root_r119_carry_16_), .CO(add_3_root_r119_carry_17_), .S(
        add_1_root_r119_A_16_) );
  ADDFX2 U146 ( .A(in_17bit_b[15]), .B(in_17bit_b[13]), .CI(
        add_1_root_r115_carry_19_), .CO(add_1_root_r115_carry_20_), .S(
        add_1_root_r115_SUM_19_) );
  ADDFX2 U147 ( .A(in_17bit_b[7]), .B(in_17bit_b[3]), .CI(
        add_1_root_r112_carry_7_), .CO(add_1_root_r112_carry_8_), .S(
        add_1_root_r112_SUM_7_) );
  ADDFX2 U148 ( .A(in_17bit_b[4]), .B(in_17bit_b[3]), .CI(
        add_2_root_r119_carry_8_), .CO(add_2_root_r119_carry_9_), .S(
        add_2_root_r119_SUM_8_) );
  ADDFX2 U149 ( .A(in_17bit_b[4]), .B(in_17bit_b[3]), .CI(
        add_3_root_r119_carry_5_), .CO(add_3_root_r119_carry_6_), .S(
        add_1_root_r119_A_5_) );
  ADDFX2 U150 ( .A(in_17bit_b[14]), .B(in_17bit_b[13]), .CI(
        add_2_root_r119_carry_18_), .CO(add_2_root_r119_carry_19_), .S(
        add_2_root_r119_SUM_18_) );
  ADDFX2 U151 ( .A(in_17bit_b[15]), .B(in_17bit_b[14]), .CI(
        add_2_root_r119_carry_19_), .CO(add_2_root_r119_carry_20_), .S(
        add_2_root_r119_SUM_19_) );
  BUFX3 U152 ( .A(in_17bit_b[16]), .Y(n42) );
  INVX1 U153 ( .A(n262), .Y(in_17bit_b[16]) );
  INVX1 U154 ( .A(n204), .Y(n100) );
  NAND3BX1 U155 ( .AN(in_8bit[5]), .B(n50), .C(in_8bit[3]), .Y(n204) );
  INVX1 U156 ( .A(in_8bit[0]), .Y(n46) );
  INVX1 U157 ( .A(n56), .Y(n58) );
  XNOR2X1 U158 ( .A(n58), .B(n28), .Y(N29) );
  NAND2X1 U159 ( .A(sub_add_54_b0_carry[15]), .B(n180), .Y(n28) );
  CLKINVX3 U160 ( .A(n209), .Y(in_17bit_b[0]) );
  OAI21XL U161 ( .A0(n261), .A1(n262), .B0(n260), .Y(N463) );
  AOI22X1 U162 ( .A0(N221), .A1(n41), .B0(N363), .B1(n40), .Y(n260) );
  INVX1 U163 ( .A(n182), .Y(n261) );
  CLKINVX3 U164 ( .A(n254), .Y(in_17bit_b[15]) );
  NAND2X1 U165 ( .A(n211), .B(n210), .Y(N447) );
  AOI22X1 U166 ( .A0(N108), .A1(n255), .B0(N205), .B1(n41), .Y(n210) );
  AOI22X1 U167 ( .A0(N347), .A1(n40), .B0(n182), .B1(in_17bit_b[0]), .Y(n211)
         );
  NAND2X1 U168 ( .A(n214), .B(n213), .Y(N448) );
  AOI22X1 U169 ( .A0(N109), .A1(n255), .B0(N206), .B1(n41), .Y(n213) );
  AOI22X1 U170 ( .A0(N348), .A1(n40), .B0(n182), .B1(n181), .Y(n214) );
  INVX1 U171 ( .A(n212), .Y(n181) );
  NAND2X1 U172 ( .A(n217), .B(n216), .Y(N449) );
  AOI22X1 U173 ( .A0(N110), .A1(n255), .B0(N207), .B1(n41), .Y(n216) );
  AOI22X1 U174 ( .A0(N349), .A1(n40), .B0(n182), .B1(in_17bit_b[2]), .Y(n217)
         );
  NAND2X1 U175 ( .A(n220), .B(n219), .Y(N450) );
  AOI22X1 U176 ( .A0(N111), .A1(n255), .B0(N208), .B1(n41), .Y(n219) );
  AOI22X1 U177 ( .A0(N350), .A1(n40), .B0(n182), .B1(in_17bit_b[3]), .Y(n220)
         );
  NAND2X1 U178 ( .A(n223), .B(n222), .Y(N451) );
  AOI22X1 U179 ( .A0(N112), .A1(n255), .B0(N209), .B1(n41), .Y(n222) );
  AOI22X1 U180 ( .A0(N351), .A1(n40), .B0(n182), .B1(in_17bit_b[4]), .Y(n223)
         );
  NAND2X1 U181 ( .A(n226), .B(n225), .Y(N452) );
  AOI22X1 U182 ( .A0(N113), .A1(n255), .B0(N210), .B1(n41), .Y(n225) );
  AOI22X1 U183 ( .A0(N352), .A1(n40), .B0(n182), .B1(in_17bit_b[5]), .Y(n226)
         );
  NAND2X1 U184 ( .A(n229), .B(n228), .Y(N453) );
  AOI22X1 U185 ( .A0(N114), .A1(n255), .B0(N211), .B1(n41), .Y(n228) );
  AOI22X1 U186 ( .A0(N353), .A1(n40), .B0(n182), .B1(in_17bit_b[6]), .Y(n229)
         );
  NAND2X1 U187 ( .A(n232), .B(n231), .Y(N454) );
  AOI22X1 U188 ( .A0(N115), .A1(n255), .B0(N212), .B1(n41), .Y(n231) );
  AOI22X1 U189 ( .A0(N354), .A1(n40), .B0(n182), .B1(in_17bit_b[7]), .Y(n232)
         );
  NAND2X1 U190 ( .A(n235), .B(n234), .Y(N455) );
  AOI22X1 U191 ( .A0(N116), .A1(n255), .B0(N213), .B1(n41), .Y(n234) );
  AOI22X1 U192 ( .A0(N355), .A1(n40), .B0(n182), .B1(in_17bit_b[8]), .Y(n235)
         );
  NAND2X1 U193 ( .A(n238), .B(n237), .Y(N456) );
  AOI22X1 U194 ( .A0(N117), .A1(n255), .B0(N214), .B1(n41), .Y(n237) );
  AOI22X1 U195 ( .A0(N356), .A1(n40), .B0(n182), .B1(in_17bit_b[9]), .Y(n238)
         );
  NAND2X1 U196 ( .A(n241), .B(n240), .Y(N457) );
  AOI22X1 U197 ( .A0(N118), .A1(n255), .B0(N215), .B1(n41), .Y(n240) );
  AOI22X1 U198 ( .A0(N357), .A1(n40), .B0(n182), .B1(in_17bit_b[10]), .Y(n241)
         );
  NAND2X1 U199 ( .A(n244), .B(n243), .Y(N458) );
  AOI22X1 U200 ( .A0(N119), .A1(n255), .B0(N216), .B1(n41), .Y(n243) );
  AOI22X1 U201 ( .A0(N358), .A1(n40), .B0(n182), .B1(in_17bit_b[11]), .Y(n244)
         );
  NAND2X1 U202 ( .A(n247), .B(n246), .Y(N459) );
  AOI22X1 U203 ( .A0(N120), .A1(n255), .B0(N217), .B1(n41), .Y(n246) );
  AOI22X1 U204 ( .A0(N359), .A1(n40), .B0(n182), .B1(in_17bit_b[12]), .Y(n247)
         );
  NAND2X1 U205 ( .A(n250), .B(n249), .Y(N460) );
  AOI22X1 U206 ( .A0(N121), .A1(n255), .B0(N218), .B1(n41), .Y(n249) );
  AOI22X1 U207 ( .A0(N360), .A1(n40), .B0(n182), .B1(in_17bit_b[13]), .Y(n250)
         );
  NAND2X1 U208 ( .A(n253), .B(n252), .Y(N461) );
  AOI22X1 U209 ( .A0(N122), .A1(n255), .B0(N219), .B1(n41), .Y(n252) );
  AOI22X1 U210 ( .A0(N361), .A1(n40), .B0(n182), .B1(in_17bit_b[14]), .Y(n253)
         );
  NAND2X1 U211 ( .A(n257), .B(n256), .Y(N462) );
  AOI22X1 U212 ( .A0(N123), .A1(n255), .B0(N220), .B1(n41), .Y(n256) );
  AOI22X1 U213 ( .A0(N362), .A1(n40), .B0(n182), .B1(in_17bit_b[15]), .Y(n257)
         );
  INVX1 U214 ( .A(in_8bit[3]), .Y(n48) );
  INVX1 U215 ( .A(n74), .Y(n71) );
  OAI21XL U216 ( .A0(n43), .A1(n76), .B0(n75), .Y(n80) );
  MXI2XL U217 ( .A(n2), .B(n19), .S0(n27), .Y(out[16]) );
  AOI22X1 U218 ( .A0(N27), .A1(n56), .B0(in_17bit[14]), .B1(n58), .Y(n251) );
  AOI22X1 U219 ( .A0(N28), .A1(n56), .B0(in_17bit[15]), .B1(n58), .Y(n254) );
  AOI22X1 U220 ( .A0(N17), .A1(n56), .B0(in_17bit[4]), .B1(n58), .Y(n221) );
  AOI22X1 U221 ( .A0(N18), .A1(n56), .B0(in_17bit[5]), .B1(n58), .Y(n224) );
  AOI22X1 U222 ( .A0(N19), .A1(n56), .B0(in_17bit[6]), .B1(n58), .Y(n227) );
  AOI22X1 U223 ( .A0(N26), .A1(n56), .B0(in_17bit[13]), .B1(n58), .Y(n248) );
  AOI22X1 U224 ( .A0(N20), .A1(n56), .B0(in_17bit[7]), .B1(n58), .Y(n230) );
  AOI22X1 U225 ( .A0(N21), .A1(n56), .B0(in_17bit[8]), .B1(n58), .Y(n233) );
  AOI22X1 U226 ( .A0(N22), .A1(n56), .B0(in_17bit[9]), .B1(n58), .Y(n236) );
  AOI22X1 U227 ( .A0(N23), .A1(n56), .B0(in_17bit[10]), .B1(n58), .Y(n239) );
  AOI22X1 U228 ( .A0(N24), .A1(n56), .B0(in_17bit[11]), .B1(n58), .Y(n242) );
  AOI22X1 U229 ( .A0(N25), .A1(n56), .B0(in_17bit[12]), .B1(n58), .Y(n245) );
  AOI22X1 U230 ( .A0(N16), .A1(n56), .B0(in_17bit[3]), .B1(n58), .Y(n218) );
  INVX1 U231 ( .A(n60), .Y(n82) );
  NAND2BX1 U232 ( .AN(n74), .B(n14), .Y(n60) );
  NAND2X1 U233 ( .A(n37), .B(n9), .Y(n74) );
  AND2X2 U234 ( .A(n82), .B(n16), .Y(n29) );
  AND2X2 U235 ( .A(n29), .B(n3), .Y(n30) );
  AND2X2 U236 ( .A(n30), .B(n4), .Y(n31) );
  AND2X2 U237 ( .A(n31), .B(n5), .Y(n32) );
  AND2X2 U238 ( .A(n32), .B(n6), .Y(n33) );
  BUFX3 U239 ( .A(n258), .Y(n40) );
  OAI2BB1X1 U240 ( .A0N(n100), .A1N(n26), .B0(n98), .Y(n258) );
  NAND2BX1 U241 ( .AN(n203), .B(n34), .Y(n98) );
  BUFX3 U242 ( .A(n259), .Y(n41) );
  OAI2BB1X1 U243 ( .A0N(n34), .A1N(n100), .B0(n99), .Y(n259) );
  NAND2BX1 U244 ( .AN(n203), .B(n26), .Y(n99) );
  NAND2X1 U245 ( .A(n96), .B(n95), .Y(n255) );
  NAND3X1 U246 ( .A(n206), .B(in_8bit[5]), .C(n94), .Y(n95) );
  NAND4BXL U247 ( .AN(n47), .B(n207), .C(n160), .D(in_8bit[1]), .Y(n96) );
  OAI2BB1X1 U248 ( .A0N(n206), .A1N(n160), .B0(n158), .Y(n182) );
  NAND3BX1 U249 ( .AN(n101), .B(n207), .C(in_8bit[5]), .Y(n158) );
  AND2X2 U250 ( .A(n97), .B(n46), .Y(n34) );
  AND2X2 U251 ( .A(n33), .B(n7), .Y(n35) );
  INVX1 U252 ( .A(in_17bit[3]), .Y(n164) );
  INVX1 U253 ( .A(in_17bit[4]), .Y(n168) );
  INVX1 U254 ( .A(in_17bit[5]), .Y(n170) );
  INVX1 U255 ( .A(in_17bit[6]), .Y(n171) );
  INVX1 U256 ( .A(in_17bit[7]), .Y(n172) );
  INVX1 U257 ( .A(in_17bit[8]), .Y(n173) );
  INVX1 U258 ( .A(in_17bit[9]), .Y(n174) );
  INVX1 U259 ( .A(in_17bit[10]), .Y(n175) );
  INVX1 U260 ( .A(in_17bit[11]), .Y(n176) );
  INVX1 U261 ( .A(in_17bit[12]), .Y(n177) );
  INVX1 U262 ( .A(in_17bit[13]), .Y(n178) );
  INVX1 U263 ( .A(in_17bit[14]), .Y(n179) );
  INVX1 U264 ( .A(in_17bit[15]), .Y(n180) );
  INVX1 U265 ( .A(in_17bit[1]), .Y(n162) );
  INVX1 U266 ( .A(in_17bit[2]), .Y(n163) );
  INVX1 U267 ( .A(in_17bit[0]), .Y(n161) );
  XNOR2X1 U268 ( .A(n17), .B(sub_add_75_b0_carry[12]), .Y(n36) );
  INVX1 U269 ( .A(n62), .Y(n63) );
  MX2X1 U270 ( .A(neg_mul[21]), .B(N479), .S0(n27), .Y(out[14]) );
  MX2X1 U271 ( .A(neg_mul[22]), .B(N480), .S0(n27), .Y(out[15]) );
  INVX1 U272 ( .A(n76), .Y(n77) );
  INVX1 U273 ( .A(n68), .Y(n69) );
  NAND4BBX1 U274 ( .AN(n40), .BN(n41), .C(n208), .D(n261), .Y(N446) );
  NOR3BXL U275 ( .AN(in_8bit[7]), .B(in_8bit[5]), .C(in_8bit[4]), .Y(n160) );
  NOR2X1 U276 ( .A(out[0]), .B(neg_mul[8]), .Y(n37) );
  NAND4BXL U277 ( .AN(in_8bit[7]), .B(in_8bit[4]), .C(in_8bit[1]), .D(
        in_8bit[6]), .Y(n101) );
  NAND2BX1 U278 ( .AN(n37), .B(neg_mul[9]), .Y(n68) );
  NAND2X1 U279 ( .A(out[0]), .B(neg_mul[8]), .Y(n62) );
  NAND2X1 U280 ( .A(neg_mul[10]), .B(n74), .Y(n76) );
  NOR2X1 U281 ( .A(in_8bit[6]), .B(in_8bit[4]), .Y(n202) );
  NOR2XL U282 ( .A(n43), .B(n93), .Y(n94) );
  INVX1 U283 ( .A(in_8bit[4]), .Y(n93) );
  NAND2X1 U284 ( .A(sub_add_75_b0_carry[15]), .B(n10), .Y(n38) );
  NAND2XL U285 ( .A(N29), .B(n57), .Y(n262) );
  AOI22XL U286 ( .A0(N15), .A1(n57), .B0(in_17bit[2]), .B1(n58), .Y(n215) );
  AOI22XL U287 ( .A0(in_17bit[0]), .A1(n57), .B0(in_17bit[0]), .B1(n58), .Y(
        n209) );
  AOI22XL U288 ( .A0(N14), .A1(n57), .B0(in_17bit[1]), .B1(n58), .Y(n212) );
  AOI211X4 U289 ( .A0(n52), .A1(n80), .B0(n79), .C0(n82), .Y(out[3]) );
  AOI211X4 U290 ( .A0(n52), .A1(n73), .B0(n72), .C0(n71), .Y(out[2]) );
  NOR2X4 U291 ( .A(n29), .B(n83), .Y(n84) );
  XNOR2X4 U292 ( .A(n84), .B(n3), .Y(out[5]) );
  NOR2X4 U293 ( .A(n30), .B(n88), .Y(n85) );
  XNOR2X4 U294 ( .A(n85), .B(n4), .Y(out[6]) );
  NOR2X4 U295 ( .A(n31), .B(n86), .Y(n87) );
  XNOR2X4 U296 ( .A(n87), .B(n5), .Y(out[7]) );
  NOR2X4 U297 ( .A(n32), .B(n88), .Y(n89) );
  XNOR2X4 U298 ( .A(n89), .B(n6), .Y(out[8]) );
  XNOR2X4 U299 ( .A(n90), .B(n7), .Y(out[9]) );
  XNOR2X4 U300 ( .A(n91), .B(n8), .Y(out[10]) );
  AND2X1 U301 ( .A(add_1_root_r112_carry_20_), .B(n42), .Y(
        add_1_root_r112_SUM_21_) );
  XOR2X1 U302 ( .A(n42), .B(add_1_root_r112_carry_20_), .Y(
        add_1_root_r112_SUM_20_) );
  AND2X1 U303 ( .A(add_1_root_r112_carry_19_), .B(in_17bit_b[15]), .Y(
        add_1_root_r112_carry_20_) );
  XOR2X1 U304 ( .A(in_17bit_b[15]), .B(add_1_root_r112_carry_19_), .Y(
        add_1_root_r112_SUM_19_) );
  AND2X1 U305 ( .A(add_1_root_r112_carry_18_), .B(in_17bit_b[14]), .Y(
        add_1_root_r112_carry_19_) );
  XOR2X1 U306 ( .A(in_17bit_b[14]), .B(add_1_root_r112_carry_18_), .Y(
        add_1_root_r112_SUM_18_) );
  AND2X1 U307 ( .A(add_1_root_r112_carry_17_), .B(in_17bit_b[13]), .Y(
        add_1_root_r112_carry_18_) );
  XOR2X1 U308 ( .A(in_17bit_b[13]), .B(add_1_root_r112_carry_17_), .Y(
        add_1_root_r112_SUM_17_) );
  AND2X1 U309 ( .A(add_2_root_r119_carry_21_), .B(n42), .Y(
        add_2_root_r119_SUM_22_) );
  XOR2X1 U310 ( .A(n42), .B(add_2_root_r119_carry_21_), .Y(
        add_2_root_r119_SUM_21_) );
  AND2X1 U311 ( .A(in_17bit_b[1]), .B(in_17bit_b[0]), .Y(
        add_2_root_r119_carry_6_) );
  XOR2X1 U312 ( .A(in_17bit_b[0]), .B(in_17bit_b[1]), .Y(
        add_2_root_r119_SUM_5_) );
  AND2X1 U313 ( .A(add_1_root_r119_carry[22]), .B(n42), .Y(
        add_1_root_r119_SUM_23_) );
  XOR2X1 U314 ( .A(n42), .B(add_1_root_r119_carry[22]), .Y(
        add_1_root_r119_SUM_22_) );
  AND2X1 U315 ( .A(add_1_root_r119_carry[21]), .B(in_17bit_b[15]), .Y(
        add_1_root_r119_carry[22]) );
  XOR2X1 U316 ( .A(in_17bit_b[15]), .B(add_1_root_r119_carry[21]), .Y(
        add_1_root_r119_SUM_21_) );
  AND2X1 U317 ( .A(add_1_root_r119_carry[20]), .B(in_17bit_b[14]), .Y(
        add_1_root_r119_carry[21]) );
  XOR2X1 U318 ( .A(in_17bit_b[14]), .B(add_1_root_r119_carry[20]), .Y(
        add_1_root_r119_SUM_20_) );
  AND2X1 U319 ( .A(add_1_root_r119_A_6_), .B(in_17bit_b[0]), .Y(
        add_1_root_r119_carry[7]) );
  XOR2X1 U320 ( .A(in_17bit_b[0]), .B(add_1_root_r119_A_6_), .Y(
        add_1_root_r119_SUM_6_) );
  AND2X1 U321 ( .A(add_3_root_r119_carry_18_), .B(n42), .Y(
        add_1_root_r119_A_19_) );
  XOR2X1 U322 ( .A(n42), .B(add_3_root_r119_carry_18_), .Y(
        add_1_root_r119_A_18_) );
  AND2X1 U323 ( .A(in_17bit_b[1]), .B(in_17bit_b[0]), .Y(
        add_3_root_r119_carry_3_) );
  XOR2X1 U324 ( .A(in_17bit_b[0]), .B(in_17bit_b[1]), .Y(add_1_root_r119_A_2_)
         );
  AND2X1 U325 ( .A(add_2_root_r115_carry_19_), .B(n42), .Y(
        add_2_root_r115_SUM_20_) );
  XOR2X1 U326 ( .A(n42), .B(add_2_root_r115_carry_19_), .Y(
        add_2_root_r115_SUM_19_) );
  AND2X1 U327 ( .A(add_2_root_r115_carry_18_), .B(in_17bit_b[15]), .Y(
        add_2_root_r115_carry_19_) );
  XOR2X1 U328 ( .A(in_17bit_b[15]), .B(add_2_root_r115_carry_18_), .Y(
        add_2_root_r115_SUM_18_) );
  AND2X1 U329 ( .A(in_17bit_b[2]), .B(in_17bit_b[0]), .Y(
        add_2_root_r115_carry_4_) );
  XOR2X1 U330 ( .A(in_17bit_b[0]), .B(in_17bit_b[2]), .Y(
        add_2_root_r115_SUM_3_) );
  AND2X1 U331 ( .A(add_1_root_r115_carry_22_), .B(n42), .Y(
        add_1_root_r115_SUM_23_) );
  XOR2X1 U332 ( .A(n42), .B(add_1_root_r115_carry_22_), .Y(
        add_1_root_r115_SUM_22_) );
  AND2X1 U333 ( .A(add_1_root_r115_carry_21_), .B(in_17bit_b[15]), .Y(
        add_1_root_r115_carry_22_) );
  XOR2X1 U334 ( .A(in_17bit_b[15]), .B(add_1_root_r115_carry_21_), .Y(
        add_1_root_r115_SUM_21_) );
  AND2X1 U335 ( .A(in_17bit_b[2]), .B(in_17bit_b[0]), .Y(
        add_1_root_r115_carry_7_) );
  XOR2X1 U336 ( .A(in_17bit_b[0]), .B(in_17bit_b[2]), .Y(
        add_1_root_r115_SUM_6_) );
  XOR2X1 U337 ( .A(n180), .B(sub_add_54_b0_carry[15]), .Y(N28) );
  AND2X1 U338 ( .A(sub_add_54_b0_carry[14]), .B(n179), .Y(
        sub_add_54_b0_carry[15]) );
  XOR2X1 U339 ( .A(n179), .B(sub_add_54_b0_carry[14]), .Y(N27) );
  AND2X1 U340 ( .A(sub_add_54_b0_carry[13]), .B(n178), .Y(
        sub_add_54_b0_carry[14]) );
  XOR2X1 U341 ( .A(n178), .B(sub_add_54_b0_carry[13]), .Y(N26) );
  AND2X1 U342 ( .A(sub_add_54_b0_carry[12]), .B(n177), .Y(
        sub_add_54_b0_carry[13]) );
  XOR2X1 U343 ( .A(n177), .B(sub_add_54_b0_carry[12]), .Y(N25) );
  AND2X1 U344 ( .A(sub_add_54_b0_carry[11]), .B(n176), .Y(
        sub_add_54_b0_carry[12]) );
  XOR2X1 U345 ( .A(n176), .B(sub_add_54_b0_carry[11]), .Y(N24) );
  AND2X1 U346 ( .A(sub_add_54_b0_carry[10]), .B(n175), .Y(
        sub_add_54_b0_carry[11]) );
  XOR2X1 U347 ( .A(n175), .B(sub_add_54_b0_carry[10]), .Y(N23) );
  AND2X1 U348 ( .A(sub_add_54_b0_carry[9]), .B(n174), .Y(
        sub_add_54_b0_carry[10]) );
  XOR2X1 U349 ( .A(n174), .B(sub_add_54_b0_carry[9]), .Y(N22) );
  AND2X1 U350 ( .A(sub_add_54_b0_carry[8]), .B(n173), .Y(
        sub_add_54_b0_carry[9]) );
  XOR2X1 U351 ( .A(n173), .B(sub_add_54_b0_carry[8]), .Y(N21) );
  AND2X1 U352 ( .A(sub_add_54_b0_carry[7]), .B(n172), .Y(
        sub_add_54_b0_carry[8]) );
  XOR2X1 U353 ( .A(n172), .B(sub_add_54_b0_carry[7]), .Y(N20) );
  AND2X1 U354 ( .A(sub_add_54_b0_carry[6]), .B(n171), .Y(
        sub_add_54_b0_carry[7]) );
  XOR2X1 U355 ( .A(n171), .B(sub_add_54_b0_carry[6]), .Y(N19) );
  AND2X1 U356 ( .A(sub_add_54_b0_carry[5]), .B(n170), .Y(
        sub_add_54_b0_carry[6]) );
  XOR2X1 U357 ( .A(n170), .B(sub_add_54_b0_carry[5]), .Y(N18) );
  AND2X1 U358 ( .A(sub_add_54_b0_carry[4]), .B(n168), .Y(
        sub_add_54_b0_carry[5]) );
  XOR2X1 U359 ( .A(n168), .B(sub_add_54_b0_carry[4]), .Y(N17) );
  AND2X1 U360 ( .A(sub_add_54_b0_carry[3]), .B(n164), .Y(
        sub_add_54_b0_carry[4]) );
  XOR2X1 U361 ( .A(n164), .B(sub_add_54_b0_carry[3]), .Y(N16) );
  AND2X1 U362 ( .A(sub_add_54_b0_carry[2]), .B(n163), .Y(
        sub_add_54_b0_carry[3]) );
  XOR2X1 U363 ( .A(n163), .B(sub_add_54_b0_carry[2]), .Y(N15) );
  AND2X1 U364 ( .A(n161), .B(n162), .Y(sub_add_54_b0_carry[2]) );
  XOR2X1 U365 ( .A(n162), .B(n161), .Y(N14) );
  XOR2X1 U366 ( .A(n10), .B(sub_add_75_b0_carry[15]), .Y(N480) );
  AND2X1 U367 ( .A(sub_add_75_b0_carry[14]), .B(n13), .Y(
        sub_add_75_b0_carry[15]) );
  XOR2X1 U368 ( .A(n13), .B(sub_add_75_b0_carry[14]), .Y(N479) );
  AND2X1 U369 ( .A(sub_add_75_b0_carry[13]), .B(n11), .Y(
        sub_add_75_b0_carry[14]) );
  XOR2X1 U370 ( .A(n11), .B(sub_add_75_b0_carry[13]), .Y(N478) );
  AND2X1 U371 ( .A(sub_add_75_b0_carry[12]), .B(n17), .Y(
        sub_add_75_b0_carry[13]) );
  AND2X1 U372 ( .A(sub_add_75_b0_carry[11]), .B(n12), .Y(
        sub_add_75_b0_carry[12]) );
  AND2X1 U373 ( .A(n35), .B(n8), .Y(sub_add_75_b0_carry[11]) );
  AND2X1 U374 ( .A(in_17bit_b[0]), .B(in_17bit_b[4]), .Y(
        add_1_root_r112_carry_5_) );
endmodule


module multi16_9_DW01_add_0 ( A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, 
        A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, 
        A_4_, B_23_, B_22_, B_21_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, 
        B_14_, B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, 
        SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, 
        SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, 
        SUM_7_ );
  input A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_,
         A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, B_23_, B_22_,
         B_21_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_,
         B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_;
  output SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_,
         SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_,
         SUM_8_, SUM_7_;
  wire   n1, n2, n3, n4;
  wire   [23:7] carry;

  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry[7]), .CO(carry[8]), .S(SUM_7_)
         );
  ADDFX2 U1_21 ( .A(A_21_), .B(B_21_), .CI(carry[21]), .CO(carry[22]), .S(
        SUM_21_) );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry[20]), .CO(carry[21]), .S(
        SUM_20_) );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry[19]), .CO(carry[20]), .S(
        SUM_19_) );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry[18]), .CO(carry[19]), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry[17]), .CO(carry[18]), .S(
        SUM_17_) );
  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry[16]), .CO(carry[17]), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry[15]), .CO(carry[16]), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry[14]), .CO(carry[15]), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry[13]), .CO(carry[14]), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry[12]), .CO(carry[13]), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry[11]), .CO(carry[12]), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry[10]), .CO(carry[11]), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry[9]), .CO(carry[10]), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry[8]), .CO(carry[9]), .S(SUM_8_)
         );
  ADDFX2 U1_22 ( .A(A_22_), .B(B_22_), .CI(carry[22]), .CO(carry[23]), .S(
        SUM_22_) );
  AND2X2 U1 ( .A(A_4_), .B(B_4_), .Y(n1) );
  XOR2X1 U2 ( .A(B_23_), .B(carry[23]), .Y(SUM_23_) );
  OAI2BB1X1 U3 ( .A0N(n2), .A1N(A_6_), .B0(n3), .Y(carry[7]) );
  OAI21XL U4 ( .A0(A_6_), .A1(n2), .B0(B_6_), .Y(n3) );
  OAI2BB1X1 U5 ( .A0N(n1), .A1N(A_5_), .B0(n4), .Y(n2) );
  OAI21XL U6 ( .A0(A_5_), .A1(n1), .B0(B_5_), .Y(n4) );
endmodule


module multi16_9_DW01_add_4 ( A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, 
        A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, 
        B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, 
        B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, SUM_22_, SUM_21_, SUM_20_, 
        SUM_19_, SUM_18_, SUM_17_, SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, 
        SUM_11_, SUM_10_, SUM_9_, SUM_8_, SUM_7_ );
  input A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_,
         A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, B_20_, B_19_,
         B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, B_10_, B_9_,
         B_8_, B_7_, B_6_, B_5_;
  output SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_,
         SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_,
         SUM_7_;
  wire   carry_21_, carry_20_, carry_19_, carry_18_, carry_17_, carry_16_,
         carry_15_, carry_14_, carry_13_, carry_12_, carry_11_, carry_10_,
         carry_9_, carry_8_, carry_7_, n1;

  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry_16_), .CO(carry_17_), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry_15_), .CO(carry_16_), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry_14_), .CO(carry_15_), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry_13_), .CO(carry_14_), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry_12_), .CO(carry_13_), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry_11_), .CO(carry_12_), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry_10_), .CO(carry_11_), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry_9_), .CO(carry_10_), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry_8_), .CO(carry_9_), .S(SUM_8_)
         );
  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry_7_), .CO(carry_8_), .S(SUM_7_)
         );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry_20_), .CO(carry_21_), .S(
        SUM_20_) );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry_19_), .CO(carry_20_), .S(
        SUM_19_) );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry_18_), .CO(carry_19_), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry_17_), .CO(carry_18_), .S(
        SUM_17_) );
  ADDFX2 U1_21 ( .A(A_21_), .B(B_21_), .CI(carry_21_), .CO(SUM_22_), .S(
        SUM_21_) );
  OAI2BB1X1 U1 ( .A0N(A_6_), .A1N(B_6_), .B0(n1), .Y(carry_7_) );
  OAI211X1 U2 ( .A0(B_6_), .A1(A_6_), .B0(A_5_), .C0(B_5_), .Y(n1) );
endmodule


module multi16_9_DW01_add_6 ( A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, 
        A_16_, A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, 
        A_6_, A_5_, A_4_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, 
        B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, 
        SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, 
        SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, 
        SUM_7_ );
  input A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_,
         A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, B_20_,
         B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, B_10_,
         B_9_, B_8_, B_7_, B_6_, B_5_, B_4_;
  output SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_,
         SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_,
         SUM_8_, SUM_7_;
  wire   n1, n2, n3, n4, n5, n6;
  wire   [21:7] carry;

  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry[7]), .CO(carry[8]), .S(SUM_7_)
         );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry[18]), .CO(carry[19]), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry[17]), .CO(carry[18]), .S(
        SUM_17_) );
  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry[16]), .CO(carry[17]), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry[15]), .CO(carry[16]), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry[14]), .CO(carry[15]), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry[13]), .CO(carry[14]), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry[12]), .CO(carry[13]), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry[11]), .CO(carry[12]), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry[10]), .CO(carry[11]), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry[9]), .CO(carry[10]), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry[8]), .CO(carry[9]), .S(SUM_8_)
         );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry[19]), .CO(carry[20]), .S(
        SUM_19_) );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry[20]), .CO(carry[21]), .S(
        SUM_20_) );
  AND2X2 U1 ( .A(A_22_), .B(n2), .Y(n1) );
  AND2X2 U2 ( .A(A_21_), .B(carry[21]), .Y(n2) );
  AND2X2 U3 ( .A(A_4_), .B(B_4_), .Y(n3) );
  XOR2X1 U4 ( .A(A_23_), .B(n1), .Y(SUM_23_) );
  XOR2X1 U5 ( .A(A_21_), .B(carry[21]), .Y(SUM_21_) );
  XOR2X1 U6 ( .A(A_22_), .B(n2), .Y(SUM_22_) );
  OAI2BB1X1 U7 ( .A0N(n4), .A1N(A_6_), .B0(n5), .Y(carry[7]) );
  OAI21XL U8 ( .A0(A_6_), .A1(n4), .B0(B_6_), .Y(n5) );
  OAI2BB1X1 U9 ( .A0N(n3), .A1N(A_5_), .B0(n6), .Y(n4) );
  OAI21XL U10 ( .A0(A_5_), .A1(n3), .B0(B_5_), .Y(n6) );
endmodule


module multi16_9 ( in_17bit, in_8bit, out );
  input [16:0] in_17bit;
  input [7:0] in_8bit;
  output [16:0] out;
  wire   n250, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26,
         N27, N28, N29, N108, N109, N110, N111, N112, N113, N114, N115, N116,
         N117, N118, N119, N120, N121, N122, N123, N205, N206, N207, N208,
         N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, N219,
         N220, N221, N347, N348, N349, N350, N351, N352, N353, N354, N355,
         N356, N357, N358, N359, N360, N361, N362, N363, N446, N447, N448,
         N449, N450, N451, N452, N453, N454, N455, N456, N457, N458, N459,
         N460, N461, N462, N463, N476, N477, N478, N479, N480, N481,
         add_2_root_r119_carry_10_, add_2_root_r119_carry_11_,
         add_2_root_r119_carry_12_, add_2_root_r119_carry_13_,
         add_2_root_r119_carry_14_, add_2_root_r119_carry_15_,
         add_2_root_r119_carry_16_, add_2_root_r119_carry_17_,
         add_2_root_r119_carry_18_, add_2_root_r119_carry_19_,
         add_2_root_r119_carry_20_, add_2_root_r119_carry_21_,
         add_2_root_r119_carry_6_, add_2_root_r119_carry_7_,
         add_2_root_r119_carry_8_, add_2_root_r119_carry_9_,
         add_2_root_r119_SUM_5_, add_2_root_r119_SUM_6_,
         add_2_root_r119_SUM_7_, add_2_root_r119_SUM_8_,
         add_2_root_r119_SUM_9_, add_2_root_r119_SUM_10_,
         add_2_root_r119_SUM_11_, add_2_root_r119_SUM_12_,
         add_2_root_r119_SUM_13_, add_2_root_r119_SUM_14_,
         add_2_root_r119_SUM_15_, add_2_root_r119_SUM_16_,
         add_2_root_r119_SUM_17_, add_2_root_r119_SUM_18_,
         add_2_root_r119_SUM_19_, add_2_root_r119_SUM_20_,
         add_2_root_r119_SUM_21_, add_2_root_r119_SUM_22_,
         add_1_root_r119_SUM_6_, add_1_root_r119_SUM_7_,
         add_1_root_r119_SUM_8_, add_1_root_r119_SUM_9_,
         add_1_root_r119_SUM_10_, add_1_root_r119_SUM_11_,
         add_1_root_r119_SUM_12_, add_1_root_r119_SUM_13_,
         add_1_root_r119_SUM_14_, add_1_root_r119_SUM_15_,
         add_1_root_r119_SUM_16_, add_1_root_r119_SUM_17_,
         add_1_root_r119_SUM_18_, add_1_root_r119_SUM_19_,
         add_1_root_r119_SUM_20_, add_1_root_r119_SUM_21_,
         add_1_root_r119_SUM_22_, add_1_root_r119_SUM_23_,
         add_1_root_r119_A_2_, add_1_root_r119_A_3_, add_1_root_r119_A_4_,
         add_1_root_r119_A_5_, add_1_root_r119_A_6_, add_1_root_r119_A_7_,
         add_1_root_r119_A_8_, add_1_root_r119_A_9_, add_1_root_r119_A_10_,
         add_1_root_r119_A_11_, add_1_root_r119_A_12_, add_1_root_r119_A_13_,
         add_1_root_r119_A_14_, add_1_root_r119_A_15_, add_1_root_r119_A_16_,
         add_1_root_r119_A_17_, add_1_root_r119_A_18_, add_1_root_r119_A_19_,
         add_3_root_r119_carry_10_, add_3_root_r119_carry_11_,
         add_3_root_r119_carry_12_, add_3_root_r119_carry_13_,
         add_3_root_r119_carry_14_, add_3_root_r119_carry_15_,
         add_3_root_r119_carry_16_, add_3_root_r119_carry_17_,
         add_3_root_r119_carry_18_, add_3_root_r119_carry_3_,
         add_3_root_r119_carry_4_, add_3_root_r119_carry_5_,
         add_3_root_r119_carry_6_, add_3_root_r119_carry_7_,
         add_3_root_r119_carry_8_, add_3_root_r119_carry_9_,
         add_1_root_r112_carry_10_, add_1_root_r112_carry_11_,
         add_1_root_r112_carry_12_, add_1_root_r112_carry_13_,
         add_1_root_r112_carry_14_, add_1_root_r112_carry_15_,
         add_1_root_r112_carry_16_, add_1_root_r112_carry_17_,
         add_1_root_r112_carry_18_, add_1_root_r112_carry_19_,
         add_1_root_r112_carry_20_, add_1_root_r112_carry_5_,
         add_1_root_r112_carry_6_, add_1_root_r112_carry_7_,
         add_1_root_r112_carry_8_, add_1_root_r112_carry_9_,
         add_1_root_r112_SUM_1_, add_1_root_r112_SUM_2_,
         add_1_root_r112_SUM_3_, add_1_root_r112_SUM_4_,
         add_1_root_r112_SUM_5_, add_1_root_r112_SUM_6_,
         add_1_root_r112_SUM_7_, add_1_root_r112_SUM_8_,
         add_1_root_r112_SUM_9_, add_1_root_r112_SUM_10_,
         add_1_root_r112_SUM_11_, add_1_root_r112_SUM_12_,
         add_1_root_r112_SUM_13_, add_1_root_r112_SUM_14_,
         add_1_root_r112_SUM_15_, add_1_root_r112_SUM_16_,
         add_1_root_r112_SUM_17_, add_1_root_r112_SUM_18_,
         add_1_root_r112_SUM_19_, add_1_root_r112_SUM_20_,
         add_1_root_r112_SUM_21_, add_2_root_r115_carry_10_,
         add_2_root_r115_carry_11_, add_2_root_r115_carry_12_,
         add_2_root_r115_carry_13_, add_2_root_r115_carry_14_,
         add_2_root_r115_carry_15_, add_2_root_r115_carry_16_,
         add_2_root_r115_carry_17_, add_2_root_r115_carry_18_,
         add_2_root_r115_carry_19_, add_2_root_r115_carry_4_,
         add_2_root_r115_carry_5_, add_2_root_r115_carry_6_,
         add_2_root_r115_carry_7_, add_2_root_r115_carry_8_,
         add_2_root_r115_carry_9_, add_2_root_r115_SUM_3_,
         add_2_root_r115_SUM_4_, add_2_root_r115_SUM_5_,
         add_2_root_r115_SUM_6_, add_2_root_r115_SUM_7_,
         add_2_root_r115_SUM_8_, add_2_root_r115_SUM_9_,
         add_2_root_r115_SUM_10_, add_2_root_r115_SUM_11_,
         add_2_root_r115_SUM_12_, add_2_root_r115_SUM_13_,
         add_2_root_r115_SUM_14_, add_2_root_r115_SUM_15_,
         add_2_root_r115_SUM_16_, add_2_root_r115_SUM_17_,
         add_2_root_r115_SUM_18_, add_2_root_r115_SUM_19_,
         add_2_root_r115_SUM_20_, add_1_root_r115_carry_10_,
         add_1_root_r115_carry_11_, add_1_root_r115_carry_12_,
         add_1_root_r115_carry_13_, add_1_root_r115_carry_14_,
         add_1_root_r115_carry_15_, add_1_root_r115_carry_16_,
         add_1_root_r115_carry_17_, add_1_root_r115_carry_18_,
         add_1_root_r115_carry_19_, add_1_root_r115_carry_20_,
         add_1_root_r115_carry_21_, add_1_root_r115_carry_22_,
         add_1_root_r115_carry_7_, add_1_root_r115_carry_8_,
         add_1_root_r115_carry_9_, add_1_root_r115_SUM_6_,
         add_1_root_r115_SUM_7_, add_1_root_r115_SUM_8_,
         add_1_root_r115_SUM_9_, add_1_root_r115_SUM_10_,
         add_1_root_r115_SUM_11_, add_1_root_r115_SUM_12_,
         add_1_root_r115_SUM_13_, add_1_root_r115_SUM_14_,
         add_1_root_r115_SUM_15_, add_1_root_r115_SUM_16_,
         add_1_root_r115_SUM_17_, add_1_root_r115_SUM_18_,
         add_1_root_r115_SUM_19_, add_1_root_r115_SUM_20_,
         add_1_root_r115_SUM_21_, add_1_root_r115_SUM_22_,
         add_1_root_r115_SUM_23_, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249;
  wire   [16:0] in_17bit_b;
  wire   [23:8] neg_mul;
  wire   [16:10] sub_add_75_b0_carry;
  wire   [15:2] sub_add_54_b0_carry;
  wire   [22:7] add_1_root_r119_carry;

  multi16_9_DW01_add_0 add_0_root_r119 ( .A_22_(add_2_root_r119_SUM_22_), 
        .A_21_(add_2_root_r119_SUM_21_), .A_20_(add_2_root_r119_SUM_20_), 
        .A_19_(add_2_root_r119_SUM_19_), .A_18_(add_2_root_r119_SUM_18_), 
        .A_17_(add_2_root_r119_SUM_17_), .A_16_(add_2_root_r119_SUM_16_), 
        .A_15_(add_2_root_r119_SUM_15_), .A_14_(add_2_root_r119_SUM_14_), 
        .A_13_(add_2_root_r119_SUM_13_), .A_12_(add_2_root_r119_SUM_12_), 
        .A_11_(add_2_root_r119_SUM_11_), .A_10_(add_2_root_r119_SUM_10_), 
        .A_9_(add_2_root_r119_SUM_9_), .A_8_(add_2_root_r119_SUM_8_), .A_7_(
        add_2_root_r119_SUM_7_), .A_6_(add_2_root_r119_SUM_6_), .A_5_(
        add_2_root_r119_SUM_5_), .A_4_(in_17bit_b[0]), .B_23_(
        add_1_root_r119_SUM_23_), .B_22_(add_1_root_r119_SUM_22_), .B_21_(
        add_1_root_r119_SUM_21_), .B_20_(add_1_root_r119_SUM_20_), .B_19_(
        add_1_root_r119_SUM_19_), .B_18_(add_1_root_r119_SUM_18_), .B_17_(
        add_1_root_r119_SUM_17_), .B_16_(add_1_root_r119_SUM_16_), .B_15_(
        add_1_root_r119_SUM_15_), .B_14_(add_1_root_r119_SUM_14_), .B_13_(
        add_1_root_r119_SUM_13_), .B_12_(add_1_root_r119_SUM_12_), .B_11_(
        add_1_root_r119_SUM_11_), .B_10_(add_1_root_r119_SUM_10_), .B_9_(
        add_1_root_r119_SUM_9_), .B_8_(add_1_root_r119_SUM_8_), .B_7_(
        add_1_root_r119_SUM_7_), .B_6_(add_1_root_r119_SUM_6_), .B_5_(
        add_1_root_r119_A_5_), .B_4_(add_1_root_r119_A_4_), .SUM_23_(N363), 
        .SUM_22_(N362), .SUM_21_(N361), .SUM_20_(N360), .SUM_19_(N359), 
        .SUM_18_(N358), .SUM_17_(N357), .SUM_16_(N356), .SUM_15_(N355), 
        .SUM_14_(N354), .SUM_13_(N353), .SUM_12_(N352), .SUM_11_(N351), 
        .SUM_10_(N350), .SUM_9_(N349), .SUM_8_(N348), .SUM_7_(N347) );
  multi16_9_DW01_add_4 add_0_root_r112 ( .A_21_(n36), .A_20_(in_17bit_b[15]), 
        .A_19_(in_17bit_b[14]), .A_18_(in_17bit_b[13]), .A_17_(in_17bit_b[12]), 
        .A_16_(in_17bit_b[11]), .A_15_(in_17bit_b[10]), .A_14_(in_17bit_b[9]), 
        .A_13_(in_17bit_b[8]), .A_12_(in_17bit_b[7]), .A_11_(in_17bit_b[6]), 
        .A_10_(in_17bit_b[5]), .A_9_(in_17bit_b[4]), .A_8_(in_17bit_b[3]), 
        .A_7_(in_17bit_b[2]), .A_6_(in_17bit_b[1]), .A_5_(in_17bit_b[0]), 
        .B_21_(add_1_root_r112_SUM_21_), .B_20_(add_1_root_r112_SUM_20_), 
        .B_19_(add_1_root_r112_SUM_19_), .B_18_(add_1_root_r112_SUM_18_), 
        .B_17_(add_1_root_r112_SUM_17_), .B_16_(add_1_root_r112_SUM_16_), 
        .B_15_(add_1_root_r112_SUM_15_), .B_14_(add_1_root_r112_SUM_14_), 
        .B_13_(add_1_root_r112_SUM_13_), .B_12_(add_1_root_r112_SUM_12_), 
        .B_11_(add_1_root_r112_SUM_11_), .B_10_(add_1_root_r112_SUM_10_), 
        .B_9_(add_1_root_r112_SUM_9_), .B_8_(add_1_root_r112_SUM_8_), .B_7_(
        add_1_root_r112_SUM_7_), .B_6_(add_1_root_r112_SUM_6_), .B_5_(
        add_1_root_r112_SUM_5_), .SUM_22_(N123), .SUM_21_(N122), .SUM_20_(N121), .SUM_19_(N120), .SUM_18_(N119), .SUM_17_(N118), .SUM_16_(N117), .SUM_15_(
        N116), .SUM_14_(N115), .SUM_13_(N114), .SUM_12_(N113), .SUM_11_(N112), 
        .SUM_10_(N111), .SUM_9_(N110), .SUM_8_(N109), .SUM_7_(N108) );
  multi16_9_DW01_add_6 add_0_root_r115 ( .A_23_(add_1_root_r115_SUM_23_), 
        .A_22_(add_1_root_r115_SUM_22_), .A_21_(add_1_root_r115_SUM_21_), 
        .A_20_(add_1_root_r115_SUM_20_), .A_19_(add_1_root_r115_SUM_19_), 
        .A_18_(add_1_root_r115_SUM_18_), .A_17_(add_1_root_r115_SUM_17_), 
        .A_16_(add_1_root_r115_SUM_16_), .A_15_(add_1_root_r115_SUM_15_), 
        .A_14_(add_1_root_r115_SUM_14_), .A_13_(add_1_root_r115_SUM_13_), 
        .A_12_(add_1_root_r115_SUM_12_), .A_11_(add_1_root_r115_SUM_11_), 
        .A_10_(add_1_root_r115_SUM_10_), .A_9_(add_1_root_r115_SUM_9_), .A_8_(
        add_1_root_r115_SUM_8_), .A_7_(add_1_root_r115_SUM_7_), .A_6_(
        add_1_root_r115_SUM_6_), .A_5_(in_17bit_b[1]), .A_4_(in_17bit_b[0]), 
        .B_20_(add_2_root_r115_SUM_20_), .B_19_(add_2_root_r115_SUM_19_), 
        .B_18_(add_2_root_r115_SUM_18_), .B_17_(add_2_root_r115_SUM_17_), 
        .B_16_(add_2_root_r115_SUM_16_), .B_15_(add_2_root_r115_SUM_15_), 
        .B_14_(add_2_root_r115_SUM_14_), .B_13_(add_2_root_r115_SUM_13_), 
        .B_12_(add_2_root_r115_SUM_12_), .B_11_(add_2_root_r115_SUM_11_), 
        .B_10_(add_2_root_r115_SUM_10_), .B_9_(add_2_root_r115_SUM_9_), .B_8_(
        add_2_root_r115_SUM_8_), .B_7_(add_2_root_r115_SUM_7_), .B_6_(
        add_2_root_r115_SUM_6_), .B_5_(add_2_root_r115_SUM_5_), .B_4_(
        add_2_root_r115_SUM_4_), .SUM_23_(N221), .SUM_22_(N220), .SUM_21_(N219), .SUM_20_(N218), .SUM_19_(N217), .SUM_18_(N216), .SUM_17_(N215), .SUM_16_(
        N214), .SUM_15_(N213), .SUM_14_(N212), .SUM_13_(N211), .SUM_12_(N210), 
        .SUM_11_(N209), .SUM_10_(N208), .SUM_9_(N207), .SUM_8_(N206), .SUM_7_(
        N205) );
  TLATX1 neg_mul_reg_16_ ( .G(N446), .D(N456), .QN(n7) );
  TLATX1 neg_mul_reg_15_ ( .G(N446), .D(N455), .QN(n6) );
  TLATX1 neg_mul_reg_14_ ( .G(N446), .D(N454), .QN(n5) );
  TLATX1 neg_mul_reg_13_ ( .G(N446), .D(N453), .Q(neg_mul[13]), .QN(n3) );
  TLATX1 neg_mul_reg_12_ ( .G(N446), .D(N452), .Q(neg_mul[12]), .QN(n4) );
  TLATX1 neg_mul_reg_11_ ( .G(N446), .D(N451), .Q(neg_mul[11]), .QN(n2) );
  TLATX1 neg_mul_reg_23_ ( .G(N446), .D(N463), .Q(neg_mul[23]), .QN(n14) );
  TLATX1 neg_mul_reg_22_ ( .G(N446), .D(N462), .Q(neg_mul[22]), .QN(n8) );
  TLATX1 neg_mul_reg_21_ ( .G(N446), .D(N461), .Q(neg_mul[21]), .QN(n9) );
  TLATX1 neg_mul_reg_20_ ( .G(N446), .D(N460), .Q(neg_mul[20]), .QN(n10) );
  TLATX1 neg_mul_reg_19_ ( .G(N446), .D(N459), .Q(neg_mul[19]), .QN(n11) );
  TLATX1 neg_mul_reg_18_ ( .G(N446), .D(N458), .Q(neg_mul[18]), .QN(n12) );
  TLATX1 neg_mul_reg_17_ ( .G(N446), .D(N457), .QN(n13) );
  TLATX1 neg_mul_reg_8_ ( .G(N446), .D(N448), .Q(neg_mul[8]) );
  TLATX1 neg_mul_reg_9_ ( .G(N446), .D(N449), .Q(neg_mul[9]), .QN(n15) );
  TLATX1 neg_mul_reg_10_ ( .G(N446), .D(N450), .Q(neg_mul[10]) );
  TLATX1 neg_mul_reg_7_ ( .G(N446), .D(N447), .Q(out[0]) );
  NOR2X2 U2 ( .A(n72), .B(n25), .Y(n20) );
  MXI2X4 U3 ( .A(n13), .B(n28), .S0(n73), .Y(out[10]) );
  CLKBUFX8 U4 ( .A(n250), .Y(out[11]) );
  MX2X2 U5 ( .A(neg_mul[18]), .B(N476), .S0(n73), .Y(n250) );
  MX2X2 U6 ( .A(neg_mul[19]), .B(N477), .S0(n73), .Y(out[12]) );
  INVX8 U7 ( .A(n72), .Y(n73) );
  MX2X1 U8 ( .A(neg_mul[20]), .B(N478), .S0(n73), .Y(out[13]) );
  MX2X1 U9 ( .A(neg_mul[21]), .B(N479), .S0(n73), .Y(out[14]) );
  MX2X1 U10 ( .A(neg_mul[22]), .B(N480), .S0(n73), .Y(out[15]) );
  OAI21XL U11 ( .A0(in_8bit[7]), .A1(n64), .B0(n63), .Y(n69) );
  NAND2BX1 U12 ( .AN(neg_mul[10]), .B(in_8bit[7]), .Y(n63) );
  CLKINVX4 U13 ( .A(in_17bit[16]), .Y(n42) );
  INVXL U14 ( .A(n44), .Y(n16) );
  XOR2X4 U15 ( .A(n70), .B(neg_mul[12]), .Y(out[5]) );
  OR2X4 U16 ( .A(n72), .B(n27), .Y(n17) );
  NOR2X4 U17 ( .A(n29), .B(n71), .Y(n19) );
  NOR2X2 U18 ( .A(n44), .B(n51), .Y(n52) );
  NOR2X1 U19 ( .A(n44), .B(n58), .Y(n60) );
  XNOR2X4 U20 ( .A(n21), .B(n6), .Y(out[8]) );
  NOR2XL U21 ( .A(n67), .B(n44), .Y(n68) );
  XNOR2X4 U22 ( .A(n44), .B(in_8bit[7]), .Y(n72) );
  INVX8 U23 ( .A(n42), .Y(n44) );
  INVXL U24 ( .A(n16), .Y(n41) );
  NOR2X2 U25 ( .A(n72), .B(n26), .Y(n21) );
  INVX1 U26 ( .A(n199), .Y(in_17bit_b[1]) );
  INVX1 U27 ( .A(n238), .Y(in_17bit_b[14]) );
  INVX1 U28 ( .A(n235), .Y(in_17bit_b[13]) );
  INVX1 U29 ( .A(n202), .Y(in_17bit_b[2]) );
  INVX1 U30 ( .A(n211), .Y(in_17bit_b[5]) );
  INVX1 U31 ( .A(n214), .Y(in_17bit_b[6]) );
  INVX1 U32 ( .A(n217), .Y(in_17bit_b[7]) );
  INVX1 U33 ( .A(n220), .Y(in_17bit_b[8]) );
  INVX1 U34 ( .A(n223), .Y(in_17bit_b[9]) );
  INVX1 U35 ( .A(n226), .Y(in_17bit_b[10]) );
  INVX1 U36 ( .A(n229), .Y(in_17bit_b[11]) );
  INVX1 U37 ( .A(n232), .Y(in_17bit_b[12]) );
  INVX1 U38 ( .A(n208), .Y(in_17bit_b[4]) );
  INVX1 U39 ( .A(n205), .Y(in_17bit_b[3]) );
  XNOR2X4 U40 ( .A(n18), .B(n5), .Y(out[7]) );
  NOR2X4 U41 ( .A(n24), .B(n71), .Y(n18) );
  XOR2X4 U42 ( .A(n19), .B(neg_mul[11]), .Y(out[4]) );
  XOR2X4 U43 ( .A(n20), .B(neg_mul[13]), .Y(out[6]) );
  INVX1 U44 ( .A(n46), .Y(n43) );
  ADDFX2 U45 ( .A(n36), .B(in_17bit_b[12]), .CI(add_1_root_r112_carry_16_), 
        .CO(add_1_root_r112_carry_17_), .S(add_1_root_r112_SUM_16_) );
  ADDFX2 U46 ( .A(add_1_root_r119_A_19_), .B(in_17bit_b[13]), .CI(
        add_1_root_r119_carry[19]), .CO(add_1_root_r119_carry[20]), .S(
        add_1_root_r119_SUM_19_) );
  ADDFX2 U47 ( .A(n36), .B(in_17bit_b[15]), .CI(add_3_root_r119_carry_17_), 
        .CO(add_3_root_r119_carry_18_), .S(add_1_root_r119_A_17_) );
  ADDFX2 U48 ( .A(n36), .B(in_17bit_b[14]), .CI(add_2_root_r115_carry_17_), 
        .CO(add_2_root_r115_carry_18_), .S(add_2_root_r115_SUM_17_) );
  ADDFX2 U49 ( .A(n36), .B(in_17bit_b[14]), .CI(add_1_root_r115_carry_20_), 
        .CO(add_1_root_r115_carry_21_), .S(add_1_root_r115_SUM_20_) );
  ADDFX2 U50 ( .A(n36), .B(in_17bit_b[15]), .CI(add_2_root_r119_carry_20_), 
        .CO(add_2_root_r119_carry_21_), .S(add_2_root_r119_SUM_20_) );
  ADDFX2 U51 ( .A(in_17bit_b[3]), .B(in_17bit_b[1]), .CI(
        add_2_root_r115_carry_4_), .CO(add_2_root_r115_carry_5_), .S(
        add_2_root_r115_SUM_4_) );
  ADDFX2 U52 ( .A(in_17bit_b[4]), .B(in_17bit_b[2]), .CI(
        add_2_root_r115_carry_5_), .CO(add_2_root_r115_carry_6_), .S(
        add_2_root_r115_SUM_5_) );
  ADDFX2 U53 ( .A(in_17bit_b[5]), .B(in_17bit_b[1]), .CI(
        add_1_root_r112_carry_5_), .CO(add_1_root_r112_carry_6_), .S(
        add_1_root_r112_SUM_5_) );
  ADDFX2 U54 ( .A(in_17bit_b[6]), .B(in_17bit_b[5]), .CI(
        add_3_root_r119_carry_7_), .CO(add_3_root_r119_carry_8_), .S(
        add_1_root_r119_A_7_) );
  ADDFX2 U55 ( .A(in_17bit_b[6]), .B(in_17bit_b[2]), .CI(
        add_1_root_r112_carry_6_), .CO(add_1_root_r112_carry_7_), .S(
        add_1_root_r112_SUM_6_) );
  ADDFX2 U56 ( .A(in_17bit_b[3]), .B(in_17bit_b[1]), .CI(
        add_1_root_r115_carry_7_), .CO(add_1_root_r115_carry_8_), .S(
        add_1_root_r115_SUM_7_) );
  ADDFX2 U57 ( .A(in_17bit_b[7]), .B(in_17bit_b[6]), .CI(
        add_3_root_r119_carry_8_), .CO(add_3_root_r119_carry_9_), .S(
        add_1_root_r119_A_8_) );
  ADDFX2 U58 ( .A(add_1_root_r119_A_7_), .B(in_17bit_b[1]), .CI(
        add_1_root_r119_carry[7]), .CO(add_1_root_r119_carry[8]), .S(
        add_1_root_r119_SUM_7_) );
  ADDFX2 U59 ( .A(in_17bit_b[2]), .B(in_17bit_b[1]), .CI(
        add_2_root_r119_carry_6_), .CO(add_2_root_r119_carry_7_), .S(
        add_2_root_r119_SUM_6_) );
  ADDFX2 U60 ( .A(in_17bit_b[4]), .B(in_17bit_b[2]), .CI(
        add_1_root_r115_carry_8_), .CO(add_1_root_r115_carry_9_), .S(
        add_1_root_r115_SUM_8_) );
  ADDFX2 U61 ( .A(in_17bit_b[8]), .B(in_17bit_b[7]), .CI(
        add_3_root_r119_carry_9_), .CO(add_3_root_r119_carry_10_), .S(
        add_1_root_r119_A_9_) );
  ADDFX2 U62 ( .A(add_1_root_r119_A_8_), .B(in_17bit_b[2]), .CI(
        add_1_root_r119_carry[8]), .CO(add_1_root_r119_carry[9]), .S(
        add_1_root_r119_SUM_8_) );
  ADDFX2 U63 ( .A(in_17bit_b[3]), .B(in_17bit_b[2]), .CI(
        add_2_root_r119_carry_7_), .CO(add_2_root_r119_carry_8_), .S(
        add_2_root_r119_SUM_7_) );
  ADDFX2 U64 ( .A(in_17bit_b[6]), .B(in_17bit_b[4]), .CI(
        add_2_root_r115_carry_7_), .CO(add_2_root_r115_carry_8_), .S(
        add_2_root_r115_SUM_7_) );
  ADDFX2 U65 ( .A(in_17bit_b[8]), .B(in_17bit_b[4]), .CI(
        add_1_root_r112_carry_8_), .CO(add_1_root_r112_carry_9_), .S(
        add_1_root_r112_SUM_8_) );
  ADDFX2 U66 ( .A(in_17bit_b[9]), .B(in_17bit_b[8]), .CI(
        add_3_root_r119_carry_10_), .CO(add_3_root_r119_carry_11_), .S(
        add_1_root_r119_A_10_) );
  ADDFX2 U67 ( .A(in_17bit_b[7]), .B(in_17bit_b[5]), .CI(
        add_2_root_r115_carry_8_), .CO(add_2_root_r115_carry_9_), .S(
        add_2_root_r115_SUM_8_) );
  ADDFX2 U68 ( .A(in_17bit_b[9]), .B(in_17bit_b[5]), .CI(
        add_1_root_r112_carry_9_), .CO(add_1_root_r112_carry_10_), .S(
        add_1_root_r112_SUM_9_) );
  ADDFX2 U69 ( .A(in_17bit_b[10]), .B(in_17bit_b[9]), .CI(
        add_3_root_r119_carry_11_), .CO(add_3_root_r119_carry_12_), .S(
        add_1_root_r119_A_11_) );
  ADDFX2 U70 ( .A(in_17bit_b[6]), .B(in_17bit_b[4]), .CI(
        add_1_root_r115_carry_10_), .CO(add_1_root_r115_carry_11_), .S(
        add_1_root_r115_SUM_10_) );
  ADDFX2 U71 ( .A(add_1_root_r119_A_10_), .B(in_17bit_b[4]), .CI(
        add_1_root_r119_carry[10]), .CO(add_1_root_r119_carry[11]), .S(
        add_1_root_r119_SUM_10_) );
  ADDFX2 U72 ( .A(in_17bit_b[5]), .B(in_17bit_b[4]), .CI(
        add_2_root_r119_carry_9_), .CO(add_2_root_r119_carry_10_), .S(
        add_2_root_r119_SUM_9_) );
  ADDFX2 U73 ( .A(in_17bit_b[8]), .B(in_17bit_b[6]), .CI(
        add_2_root_r115_carry_9_), .CO(add_2_root_r115_carry_10_), .S(
        add_2_root_r115_SUM_9_) );
  ADDFX2 U74 ( .A(in_17bit_b[10]), .B(in_17bit_b[6]), .CI(
        add_1_root_r112_carry_10_), .CO(add_1_root_r112_carry_11_), .S(
        add_1_root_r112_SUM_10_) );
  ADDFX2 U75 ( .A(in_17bit_b[7]), .B(in_17bit_b[5]), .CI(
        add_1_root_r115_carry_11_), .CO(add_1_root_r115_carry_12_), .S(
        add_1_root_r115_SUM_11_) );
  ADDFX2 U76 ( .A(in_17bit_b[11]), .B(in_17bit_b[10]), .CI(
        add_3_root_r119_carry_12_), .CO(add_3_root_r119_carry_13_), .S(
        add_1_root_r119_A_12_) );
  ADDFX2 U77 ( .A(in_17bit_b[6]), .B(in_17bit_b[5]), .CI(
        add_2_root_r119_carry_10_), .CO(add_2_root_r119_carry_11_), .S(
        add_2_root_r119_SUM_10_) );
  ADDFX2 U78 ( .A(in_17bit_b[9]), .B(in_17bit_b[7]), .CI(
        add_2_root_r115_carry_10_), .CO(add_2_root_r115_carry_11_), .S(
        add_2_root_r115_SUM_10_) );
  ADDFX2 U79 ( .A(in_17bit_b[11]), .B(in_17bit_b[7]), .CI(
        add_1_root_r112_carry_11_), .CO(add_1_root_r112_carry_12_), .S(
        add_1_root_r112_SUM_11_) );
  ADDFX2 U80 ( .A(in_17bit_b[8]), .B(in_17bit_b[6]), .CI(
        add_1_root_r115_carry_12_), .CO(add_1_root_r115_carry_13_), .S(
        add_1_root_r115_SUM_12_) );
  ADDFX2 U81 ( .A(in_17bit_b[12]), .B(in_17bit_b[11]), .CI(
        add_3_root_r119_carry_13_), .CO(add_3_root_r119_carry_14_), .S(
        add_1_root_r119_A_13_) );
  ADDFX2 U82 ( .A(add_1_root_r119_A_12_), .B(in_17bit_b[6]), .CI(
        add_1_root_r119_carry[12]), .CO(add_1_root_r119_carry[13]), .S(
        add_1_root_r119_SUM_12_) );
  ADDFX2 U83 ( .A(in_17bit_b[7]), .B(in_17bit_b[6]), .CI(
        add_2_root_r119_carry_11_), .CO(add_2_root_r119_carry_12_), .S(
        add_2_root_r119_SUM_11_) );
  ADDFX2 U84 ( .A(in_17bit_b[10]), .B(in_17bit_b[8]), .CI(
        add_2_root_r115_carry_11_), .CO(add_2_root_r115_carry_12_), .S(
        add_2_root_r115_SUM_11_) );
  ADDFX2 U85 ( .A(in_17bit_b[12]), .B(in_17bit_b[8]), .CI(
        add_1_root_r112_carry_12_), .CO(add_1_root_r112_carry_13_), .S(
        add_1_root_r112_SUM_12_) );
  ADDFX2 U86 ( .A(in_17bit_b[9]), .B(in_17bit_b[7]), .CI(
        add_1_root_r115_carry_13_), .CO(add_1_root_r115_carry_14_), .S(
        add_1_root_r115_SUM_13_) );
  ADDFX2 U87 ( .A(add_1_root_r119_A_13_), .B(in_17bit_b[7]), .CI(
        add_1_root_r119_carry[13]), .CO(add_1_root_r119_carry[14]), .S(
        add_1_root_r119_SUM_13_) );
  ADDFX2 U88 ( .A(in_17bit_b[8]), .B(in_17bit_b[7]), .CI(
        add_2_root_r119_carry_12_), .CO(add_2_root_r119_carry_13_), .S(
        add_2_root_r119_SUM_12_) );
  ADDFX2 U89 ( .A(in_17bit_b[11]), .B(in_17bit_b[9]), .CI(
        add_2_root_r115_carry_12_), .CO(add_2_root_r115_carry_13_), .S(
        add_2_root_r115_SUM_12_) );
  ADDFX2 U90 ( .A(in_17bit_b[13]), .B(in_17bit_b[9]), .CI(
        add_1_root_r112_carry_13_), .CO(add_1_root_r112_carry_14_), .S(
        add_1_root_r112_SUM_13_) );
  ADDFX2 U91 ( .A(in_17bit_b[10]), .B(in_17bit_b[8]), .CI(
        add_1_root_r115_carry_14_), .CO(add_1_root_r115_carry_15_), .S(
        add_1_root_r115_SUM_14_) );
  ADDFX2 U92 ( .A(in_17bit_b[14]), .B(in_17bit_b[13]), .CI(
        add_3_root_r119_carry_15_), .CO(add_3_root_r119_carry_16_), .S(
        add_1_root_r119_A_15_) );
  ADDFX2 U93 ( .A(add_1_root_r119_A_14_), .B(in_17bit_b[8]), .CI(
        add_1_root_r119_carry[14]), .CO(add_1_root_r119_carry[15]), .S(
        add_1_root_r119_SUM_14_) );
  ADDFX2 U94 ( .A(in_17bit_b[3]), .B(in_17bit_b[2]), .CI(
        add_3_root_r119_carry_4_), .CO(add_3_root_r119_carry_5_), .S(
        add_1_root_r119_A_4_) );
  ADDFX2 U95 ( .A(in_17bit_b[2]), .B(in_17bit_b[1]), .CI(
        add_3_root_r119_carry_3_), .CO(add_3_root_r119_carry_4_), .S(
        add_1_root_r119_A_3_) );
  ADDFX2 U96 ( .A(in_17bit_b[9]), .B(in_17bit_b[8]), .CI(
        add_2_root_r119_carry_13_), .CO(add_2_root_r119_carry_14_), .S(
        add_2_root_r119_SUM_13_) );
  ADDFX2 U97 ( .A(in_17bit_b[12]), .B(in_17bit_b[10]), .CI(
        add_2_root_r115_carry_13_), .CO(add_2_root_r115_carry_14_), .S(
        add_2_root_r115_SUM_13_) );
  ADDFX2 U98 ( .A(in_17bit_b[14]), .B(in_17bit_b[10]), .CI(
        add_1_root_r112_carry_14_), .CO(add_1_root_r112_carry_15_), .S(
        add_1_root_r112_SUM_14_) );
  ADDFX2 U99 ( .A(in_17bit_b[11]), .B(in_17bit_b[9]), .CI(
        add_1_root_r115_carry_15_), .CO(add_1_root_r115_carry_16_), .S(
        add_1_root_r115_SUM_15_) );
  ADDFX2 U100 ( .A(add_1_root_r119_A_15_), .B(in_17bit_b[9]), .CI(
        add_1_root_r119_carry[15]), .CO(add_1_root_r119_carry[16]), .S(
        add_1_root_r119_SUM_15_) );
  ADDFX2 U101 ( .A(in_17bit_b[10]), .B(in_17bit_b[9]), .CI(
        add_2_root_r119_carry_14_), .CO(add_2_root_r119_carry_15_), .S(
        add_2_root_r119_SUM_14_) );
  ADDFX2 U102 ( .A(in_17bit_b[13]), .B(in_17bit_b[11]), .CI(
        add_2_root_r115_carry_14_), .CO(add_2_root_r115_carry_15_), .S(
        add_2_root_r115_SUM_14_) );
  ADDFX2 U103 ( .A(in_17bit_b[15]), .B(in_17bit_b[11]), .CI(
        add_1_root_r112_carry_15_), .CO(add_1_root_r112_carry_16_), .S(
        add_1_root_r112_SUM_15_) );
  ADDFX2 U104 ( .A(in_17bit_b[12]), .B(in_17bit_b[10]), .CI(
        add_1_root_r115_carry_16_), .CO(add_1_root_r115_carry_17_), .S(
        add_1_root_r115_SUM_16_) );
  ADDFX2 U105 ( .A(add_1_root_r119_A_16_), .B(in_17bit_b[10]), .CI(
        add_1_root_r119_carry[16]), .CO(add_1_root_r119_carry[17]), .S(
        add_1_root_r119_SUM_16_) );
  ADDFX2 U106 ( .A(in_17bit_b[11]), .B(in_17bit_b[10]), .CI(
        add_2_root_r119_carry_15_), .CO(add_2_root_r119_carry_16_), .S(
        add_2_root_r119_SUM_15_) );
  ADDFX2 U107 ( .A(in_17bit_b[14]), .B(in_17bit_b[12]), .CI(
        add_2_root_r115_carry_15_), .CO(add_2_root_r115_carry_16_), .S(
        add_2_root_r115_SUM_15_) );
  ADDFX2 U108 ( .A(in_17bit_b[13]), .B(in_17bit_b[11]), .CI(
        add_1_root_r115_carry_17_), .CO(add_1_root_r115_carry_18_), .S(
        add_1_root_r115_SUM_17_) );
  ADDFX2 U109 ( .A(add_1_root_r119_A_17_), .B(in_17bit_b[11]), .CI(
        add_1_root_r119_carry[17]), .CO(add_1_root_r119_carry[18]), .S(
        add_1_root_r119_SUM_17_) );
  ADDFX2 U110 ( .A(in_17bit_b[12]), .B(in_17bit_b[11]), .CI(
        add_2_root_r119_carry_16_), .CO(add_2_root_r119_carry_17_), .S(
        add_2_root_r119_SUM_16_) );
  ADDFX2 U111 ( .A(in_17bit_b[14]), .B(in_17bit_b[12]), .CI(
        add_1_root_r115_carry_18_), .CO(add_1_root_r115_carry_19_), .S(
        add_1_root_r115_SUM_18_) );
  ADDFX2 U112 ( .A(add_1_root_r119_A_18_), .B(in_17bit_b[12]), .CI(
        add_1_root_r119_carry[18]), .CO(add_1_root_r119_carry[19]), .S(
        add_1_root_r119_SUM_18_) );
  ADDFX2 U113 ( .A(in_17bit_b[13]), .B(in_17bit_b[12]), .CI(
        add_2_root_r119_carry_17_), .CO(add_2_root_r119_carry_18_), .S(
        add_2_root_r119_SUM_17_) );
  ADDFX2 U114 ( .A(in_17bit_b[5]), .B(in_17bit_b[3]), .CI(
        add_2_root_r115_carry_6_), .CO(add_2_root_r115_carry_7_), .S(
        add_2_root_r115_SUM_6_) );
  ADDFX2 U115 ( .A(in_17bit_b[7]), .B(in_17bit_b[3]), .CI(
        add_1_root_r112_carry_7_), .CO(add_1_root_r112_carry_8_), .S(
        add_1_root_r112_SUM_7_) );
  ADDFX2 U116 ( .A(in_17bit_b[5]), .B(in_17bit_b[3]), .CI(
        add_1_root_r115_carry_9_), .CO(add_1_root_r115_carry_10_), .S(
        add_1_root_r115_SUM_9_) );
  ADDFX2 U117 ( .A(in_17bit_b[14]), .B(in_17bit_b[13]), .CI(
        add_2_root_r119_carry_18_), .CO(add_2_root_r119_carry_19_), .S(
        add_2_root_r119_SUM_18_) );
  ADDFX2 U118 ( .A(add_1_root_r119_A_9_), .B(in_17bit_b[3]), .CI(
        add_1_root_r119_carry[9]), .CO(add_1_root_r119_carry[10]), .S(
        add_1_root_r119_SUM_9_) );
  ADDFX2 U119 ( .A(in_17bit_b[4]), .B(in_17bit_b[3]), .CI(
        add_2_root_r119_carry_8_), .CO(add_2_root_r119_carry_9_), .S(
        add_2_root_r119_SUM_8_) );
  ADDFX2 U120 ( .A(add_1_root_r119_A_11_), .B(in_17bit_b[5]), .CI(
        add_1_root_r119_carry[11]), .CO(add_1_root_r119_carry[12]), .S(
        add_1_root_r119_SUM_11_) );
  ADDFX2 U121 ( .A(in_17bit_b[15]), .B(in_17bit_b[13]), .CI(
        add_2_root_r115_carry_16_), .CO(add_2_root_r115_carry_17_), .S(
        add_2_root_r115_SUM_16_) );
  ADDFX2 U122 ( .A(in_17bit_b[15]), .B(in_17bit_b[13]), .CI(
        add_1_root_r115_carry_19_), .CO(add_1_root_r115_carry_20_), .S(
        add_1_root_r115_SUM_19_) );
  ADDFX2 U123 ( .A(in_17bit_b[13]), .B(in_17bit_b[12]), .CI(
        add_3_root_r119_carry_14_), .CO(add_3_root_r119_carry_15_), .S(
        add_1_root_r119_A_14_) );
  ADDFX2 U124 ( .A(in_17bit_b[15]), .B(in_17bit_b[14]), .CI(
        add_3_root_r119_carry_16_), .CO(add_3_root_r119_carry_17_), .S(
        add_1_root_r119_A_16_) );
  ADDFX2 U125 ( .A(in_17bit_b[4]), .B(in_17bit_b[3]), .CI(
        add_3_root_r119_carry_5_), .CO(add_3_root_r119_carry_6_), .S(
        add_1_root_r119_A_5_) );
  ADDFX2 U126 ( .A(in_17bit_b[5]), .B(in_17bit_b[4]), .CI(
        add_3_root_r119_carry_6_), .CO(add_3_root_r119_carry_7_), .S(
        add_1_root_r119_A_6_) );
  ADDFX2 U127 ( .A(in_17bit_b[15]), .B(in_17bit_b[14]), .CI(
        add_2_root_r119_carry_19_), .CO(add_2_root_r119_carry_20_), .S(
        add_2_root_r119_SUM_19_) );
  BUFX3 U128 ( .A(in_17bit_b[16]), .Y(n36) );
  INVX1 U129 ( .A(n249), .Y(in_17bit_b[16]) );
  BUFX3 U130 ( .A(in_8bit[6]), .Y(n39) );
  BUFX3 U131 ( .A(in_8bit[1]), .Y(n38) );
  INVX1 U132 ( .A(n41), .Y(n45) );
  INVX1 U133 ( .A(in_8bit[2]), .Y(n37) );
  INVX1 U134 ( .A(in_8bit[0]), .Y(n40) );
  XNOR2X1 U135 ( .A(n46), .B(n22), .Y(N29) );
  NAND2X1 U136 ( .A(sub_add_54_b0_carry[15]), .B(n89), .Y(n22) );
  CLKINVX3 U137 ( .A(n196), .Y(in_17bit_b[0]) );
  NOR3X1 U138 ( .A(n37), .B(n94), .C(n40), .Y(n194) );
  INVX1 U139 ( .A(n248), .Y(n91) );
  OAI21XL U140 ( .A0(n248), .A1(n249), .B0(n247), .Y(N463) );
  AOI22X1 U141 ( .A0(N221), .A1(n35), .B0(N363), .B1(n34), .Y(n247) );
  CLKINVX3 U142 ( .A(n241), .Y(in_17bit_b[15]) );
  XOR2X4 U143 ( .A(n17), .B(n7), .Y(out[9]) );
  AOI32X1 U144 ( .A0(n194), .A1(n92), .A2(in_8bit[5]), .B0(n193), .B1(n192), 
        .Y(n248) );
  INVX1 U145 ( .A(n191), .Y(n92) );
  INVXL U146 ( .A(in_8bit[3]), .Y(n94) );
  NAND3BXL U147 ( .AN(in_8bit[5]), .B(n37), .C(in_8bit[3]), .Y(n185) );
  NOR4BX1 U148 ( .AN(n186), .B(n40), .C(n38), .D(in_8bit[2]), .Y(n192) );
  NOR2XL U149 ( .A(n39), .B(in_8bit[3]), .Y(n186) );
  AOI22X1 U150 ( .A0(N27), .A1(n43), .B0(in_17bit[14]), .B1(n45), .Y(n238) );
  AOI22X1 U151 ( .A0(N28), .A1(n43), .B0(in_17bit[15]), .B1(n45), .Y(n241) );
  AOI22X1 U152 ( .A0(N17), .A1(n43), .B0(in_17bit[4]), .B1(n45), .Y(n208) );
  AOI22X1 U153 ( .A0(N18), .A1(n43), .B0(in_17bit[5]), .B1(n45), .Y(n211) );
  AOI22X1 U154 ( .A0(N19), .A1(n43), .B0(in_17bit[6]), .B1(n16), .Y(n214) );
  AOI22X1 U155 ( .A0(N20), .A1(n43), .B0(in_17bit[7]), .B1(n46), .Y(n217) );
  AOI22X1 U156 ( .A0(N21), .A1(n43), .B0(in_17bit[8]), .B1(n16), .Y(n220) );
  AOI22X1 U157 ( .A0(N22), .A1(n43), .B0(in_17bit[9]), .B1(n45), .Y(n223) );
  AOI22X1 U158 ( .A0(N23), .A1(n43), .B0(in_17bit[10]), .B1(n16), .Y(n226) );
  AOI22X1 U159 ( .A0(N24), .A1(n43), .B0(in_17bit[11]), .B1(n46), .Y(n229) );
  AOI22X1 U160 ( .A0(N25), .A1(n43), .B0(in_17bit[12]), .B1(n45), .Y(n232) );
  AOI22X1 U161 ( .A0(N26), .A1(n43), .B0(in_17bit[13]), .B1(n16), .Y(n235) );
  AOI22X1 U162 ( .A0(N15), .A1(n43), .B0(in_17bit[2]), .B1(n16), .Y(n202) );
  NAND3X1 U163 ( .A(in_8bit[2]), .B(n94), .C(in_8bit[5]), .Y(n184) );
  AND2X2 U164 ( .A(n29), .B(n2), .Y(n23) );
  AND2X2 U165 ( .A(n25), .B(n3), .Y(n24) );
  BUFX3 U166 ( .A(n245), .Y(n34) );
  OAI32X1 U167 ( .A0(n184), .A1(in_8bit[0]), .A2(n191), .B0(n185), .B1(n183), 
        .Y(n245) );
  AND2X2 U168 ( .A(n23), .B(n4), .Y(n25) );
  BUFX3 U169 ( .A(n246), .Y(n35) );
  OAI32X1 U170 ( .A0(n191), .A1(in_8bit[0]), .A2(n185), .B0(n184), .B1(n183), 
        .Y(n246) );
  AND2X2 U171 ( .A(n24), .B(n5), .Y(n26) );
  INVX1 U172 ( .A(in_17bit[13]), .Y(n87) );
  INVX1 U173 ( .A(in_17bit[2]), .Y(n76) );
  INVX1 U174 ( .A(in_17bit[4]), .Y(n78) );
  INVX1 U175 ( .A(in_17bit[5]), .Y(n79) );
  INVX1 U176 ( .A(in_17bit[6]), .Y(n80) );
  INVX1 U177 ( .A(in_17bit[7]), .Y(n81) );
  INVX1 U178 ( .A(in_17bit[8]), .Y(n82) );
  INVX1 U179 ( .A(in_17bit[9]), .Y(n83) );
  INVX1 U180 ( .A(in_17bit[10]), .Y(n84) );
  INVX1 U181 ( .A(in_17bit[11]), .Y(n85) );
  INVX1 U182 ( .A(in_17bit[12]), .Y(n86) );
  INVX1 U183 ( .A(in_17bit[14]), .Y(n88) );
  INVX1 U184 ( .A(in_17bit[15]), .Y(n89) );
  INVX1 U185 ( .A(in_17bit[1]), .Y(n75) );
  INVX1 U186 ( .A(in_17bit[3]), .Y(n77) );
  INVX1 U187 ( .A(in_17bit[0]), .Y(n74) );
  NAND2X1 U188 ( .A(n198), .B(n197), .Y(N447) );
  AOI22X1 U189 ( .A0(N108), .A1(n242), .B0(N205), .B1(n35), .Y(n197) );
  AOI22X1 U190 ( .A0(N347), .A1(n34), .B0(n91), .B1(in_17bit_b[0]), .Y(n198)
         );
  NAND2X1 U191 ( .A(n201), .B(n200), .Y(N448) );
  AOI22X1 U192 ( .A0(N109), .A1(n242), .B0(N206), .B1(n35), .Y(n200) );
  AOI22X1 U193 ( .A0(N348), .A1(n34), .B0(n91), .B1(n90), .Y(n201) );
  INVX1 U194 ( .A(n199), .Y(n90) );
  NAND2X1 U195 ( .A(n204), .B(n203), .Y(N449) );
  AOI22X1 U196 ( .A0(N110), .A1(n242), .B0(N207), .B1(n35), .Y(n203) );
  AOI22X1 U197 ( .A0(N349), .A1(n34), .B0(n91), .B1(in_17bit_b[2]), .Y(n204)
         );
  NAND2X1 U198 ( .A(n207), .B(n206), .Y(N450) );
  AOI22X1 U199 ( .A0(N111), .A1(n242), .B0(N208), .B1(n35), .Y(n206) );
  AOI22X1 U200 ( .A0(N350), .A1(n34), .B0(n91), .B1(in_17bit_b[3]), .Y(n207)
         );
  NAND2X1 U201 ( .A(n210), .B(n209), .Y(N451) );
  AOI22X1 U202 ( .A0(N112), .A1(n242), .B0(N209), .B1(n35), .Y(n209) );
  AOI22X1 U203 ( .A0(N351), .A1(n34), .B0(n91), .B1(in_17bit_b[4]), .Y(n210)
         );
  NAND2X1 U204 ( .A(n213), .B(n212), .Y(N452) );
  AOI22X1 U205 ( .A0(N113), .A1(n242), .B0(N210), .B1(n35), .Y(n212) );
  AOI22X1 U206 ( .A0(N352), .A1(n34), .B0(n91), .B1(in_17bit_b[5]), .Y(n213)
         );
  NAND2X1 U207 ( .A(n216), .B(n215), .Y(N453) );
  AOI22X1 U208 ( .A0(N114), .A1(n242), .B0(N211), .B1(n35), .Y(n215) );
  AOI22X1 U209 ( .A0(N353), .A1(n34), .B0(n91), .B1(in_17bit_b[6]), .Y(n216)
         );
  NAND2X1 U210 ( .A(n219), .B(n218), .Y(N454) );
  AOI22X1 U211 ( .A0(N115), .A1(n242), .B0(N212), .B1(n35), .Y(n218) );
  AOI22X1 U212 ( .A0(N354), .A1(n34), .B0(n91), .B1(in_17bit_b[7]), .Y(n219)
         );
  NAND2X1 U213 ( .A(n222), .B(n221), .Y(N455) );
  AOI22X1 U214 ( .A0(N116), .A1(n242), .B0(N213), .B1(n35), .Y(n221) );
  AOI22X1 U215 ( .A0(N355), .A1(n34), .B0(n91), .B1(in_17bit_b[8]), .Y(n222)
         );
  NAND2X1 U216 ( .A(n225), .B(n224), .Y(N456) );
  AOI22X1 U217 ( .A0(N117), .A1(n242), .B0(N214), .B1(n35), .Y(n224) );
  AOI22X1 U218 ( .A0(N356), .A1(n34), .B0(n91), .B1(in_17bit_b[9]), .Y(n225)
         );
  NAND2X1 U219 ( .A(n228), .B(n227), .Y(N457) );
  AOI22X1 U220 ( .A0(N118), .A1(n242), .B0(N215), .B1(n35), .Y(n227) );
  AOI22X1 U221 ( .A0(N357), .A1(n34), .B0(n91), .B1(in_17bit_b[10]), .Y(n228)
         );
  NAND2X1 U222 ( .A(n231), .B(n230), .Y(N458) );
  AOI22X1 U223 ( .A0(N119), .A1(n242), .B0(N216), .B1(n35), .Y(n230) );
  AOI22X1 U224 ( .A0(N358), .A1(n34), .B0(n91), .B1(in_17bit_b[11]), .Y(n231)
         );
  NAND2X1 U225 ( .A(n234), .B(n233), .Y(N459) );
  AOI22X1 U226 ( .A0(N120), .A1(n242), .B0(N217), .B1(n35), .Y(n233) );
  AOI22X1 U227 ( .A0(N359), .A1(n34), .B0(n91), .B1(in_17bit_b[12]), .Y(n234)
         );
  NAND2X1 U228 ( .A(n237), .B(n236), .Y(N460) );
  AOI22X1 U229 ( .A0(N121), .A1(n242), .B0(N218), .B1(n35), .Y(n236) );
  AOI22X1 U230 ( .A0(N360), .A1(n34), .B0(n91), .B1(in_17bit_b[13]), .Y(n237)
         );
  NAND2X1 U231 ( .A(n240), .B(n239), .Y(N461) );
  AOI22X1 U232 ( .A0(N122), .A1(n242), .B0(N219), .B1(n35), .Y(n239) );
  AOI22X1 U233 ( .A0(N361), .A1(n34), .B0(n91), .B1(in_17bit_b[14]), .Y(n240)
         );
  NAND2X1 U234 ( .A(n244), .B(n243), .Y(N462) );
  AOI22X1 U235 ( .A0(N123), .A1(n242), .B0(N220), .B1(n35), .Y(n243) );
  AOI22X1 U236 ( .A0(N362), .A1(n34), .B0(n91), .B1(in_17bit_b[15]), .Y(n244)
         );
  AND2X2 U237 ( .A(n26), .B(n6), .Y(n27) );
  XNOR2X1 U238 ( .A(n13), .B(sub_add_75_b0_carry[10]), .Y(n28) );
  OAI21XL U239 ( .A0(in_8bit[7]), .A1(n48), .B0(n47), .Y(n53) );
  NAND2BX1 U240 ( .AN(neg_mul[8]), .B(in_8bit[7]), .Y(n47) );
  INVX1 U241 ( .A(n62), .Y(n59) );
  OAI21XL U242 ( .A0(in_8bit[7]), .A1(n55), .B0(n54), .Y(n61) );
  MX2X1 U243 ( .A(neg_mul[23]), .B(N481), .S0(n73), .Y(out[16]) );
  NAND4BBX1 U244 ( .AN(n34), .BN(n35), .C(n195), .D(n248), .Y(N446) );
  AOI2BB1X1 U245 ( .A0N(n190), .A1N(n189), .B0(n242), .Y(n195) );
  OR4X2 U246 ( .A(in_8bit[4]), .B(in_8bit[5]), .C(n39), .D(in_8bit[7]), .Y(
        n190) );
  OR4XL U247 ( .A(n38), .B(in_8bit[0]), .C(in_8bit[2]), .D(in_8bit[3]), .Y(
        n189) );
  NOR3X1 U248 ( .A(in_8bit[4]), .B(in_8bit[5]), .C(n93), .Y(n193) );
  NAND4X1 U249 ( .A(n39), .B(in_8bit[4]), .C(n38), .D(n93), .Y(n191) );
  NOR2X1 U250 ( .A(n62), .B(neg_mul[10]), .Y(n29) );
  NAND4X1 U251 ( .A(n38), .B(in_8bit[7]), .C(n182), .D(n40), .Y(n183) );
  NOR2X1 U252 ( .A(n39), .B(in_8bit[4]), .Y(n182) );
  NOR2X1 U253 ( .A(out[0]), .B(neg_mul[8]), .Y(n30) );
  NAND2X1 U254 ( .A(n30), .B(n15), .Y(n62) );
  NAND2X1 U255 ( .A(out[0]), .B(neg_mul[8]), .Y(n48) );
  NAND2X1 U256 ( .A(neg_mul[10]), .B(n62), .Y(n64) );
  NAND2BX1 U257 ( .AN(n30), .B(neg_mul[9]), .Y(n55) );
  NAND2X1 U258 ( .A(n188), .B(n187), .Y(n242) );
  NAND4X1 U259 ( .A(n193), .B(n194), .C(n39), .D(n38), .Y(n187) );
  NAND4X1 U260 ( .A(n192), .B(in_8bit[5]), .C(in_8bit[4]), .D(n93), .Y(n188)
         );
  NOR2X1 U261 ( .A(n50), .B(n49), .Y(n51) );
  NOR2X1 U262 ( .A(in_8bit[7]), .B(neg_mul[8]), .Y(n49) );
  NOR2X1 U263 ( .A(n93), .B(n48), .Y(n50) );
  AOI21X1 U264 ( .A0(n57), .A1(in_8bit[7]), .B0(n56), .Y(n58) );
  INVX1 U265 ( .A(n55), .Y(n57) );
  NOR2X1 U266 ( .A(in_8bit[7]), .B(neg_mul[9]), .Y(n56) );
  NAND2BX1 U267 ( .AN(neg_mul[9]), .B(in_8bit[7]), .Y(n54) );
  NOR2X1 U268 ( .A(n66), .B(n65), .Y(n67) );
  NOR2X1 U269 ( .A(in_8bit[7]), .B(neg_mul[10]), .Y(n65) );
  NOR2X1 U270 ( .A(n93), .B(n64), .Y(n66) );
  INVX1 U271 ( .A(in_8bit[7]), .Y(n93) );
  INVX1 U272 ( .A(n41), .Y(n46) );
  AOI211X4 U273 ( .A0(n44), .A1(n53), .B0(n52), .C0(n30), .Y(out[1]) );
  XNOR2X4 U274 ( .A(n44), .B(in_8bit[7]), .Y(n71) );
  NAND2XL U275 ( .A(N29), .B(n41), .Y(n249) );
  AOI22XL U276 ( .A0(N16), .A1(n41), .B0(in_17bit[3]), .B1(n16), .Y(n205) );
  AOI22XL U277 ( .A0(in_17bit[0]), .A1(n41), .B0(in_17bit[0]), .B1(n46), .Y(
        n196) );
  AOI22XL U278 ( .A0(N14), .A1(n41), .B0(in_17bit[1]), .B1(n46), .Y(n199) );
  AOI211X4 U279 ( .A0(n44), .A1(n69), .B0(n68), .C0(n29), .Y(out[3]) );
  AOI211X4 U280 ( .A0(n44), .A1(n61), .B0(n60), .C0(n59), .Y(out[2]) );
  NOR2X4 U281 ( .A(n23), .B(n71), .Y(n70) );
  AND2X1 U282 ( .A(add_1_root_r112_carry_20_), .B(n36), .Y(
        add_1_root_r112_SUM_21_) );
  XOR2X1 U283 ( .A(n36), .B(add_1_root_r112_carry_20_), .Y(
        add_1_root_r112_SUM_20_) );
  AND2X1 U284 ( .A(add_1_root_r112_carry_19_), .B(in_17bit_b[15]), .Y(
        add_1_root_r112_carry_20_) );
  XOR2X1 U285 ( .A(in_17bit_b[15]), .B(add_1_root_r112_carry_19_), .Y(
        add_1_root_r112_SUM_19_) );
  AND2X1 U286 ( .A(add_1_root_r112_carry_18_), .B(in_17bit_b[14]), .Y(
        add_1_root_r112_carry_19_) );
  XOR2X1 U287 ( .A(in_17bit_b[14]), .B(add_1_root_r112_carry_18_), .Y(
        add_1_root_r112_SUM_18_) );
  AND2X1 U288 ( .A(add_1_root_r112_carry_17_), .B(in_17bit_b[13]), .Y(
        add_1_root_r112_carry_18_) );
  XOR2X1 U289 ( .A(in_17bit_b[13]), .B(add_1_root_r112_carry_17_), .Y(
        add_1_root_r112_SUM_17_) );
  AND2X1 U290 ( .A(add_2_root_r119_carry_21_), .B(n36), .Y(
        add_2_root_r119_SUM_22_) );
  XOR2X1 U291 ( .A(n36), .B(add_2_root_r119_carry_21_), .Y(
        add_2_root_r119_SUM_21_) );
  AND2X1 U292 ( .A(in_17bit_b[1]), .B(in_17bit_b[0]), .Y(
        add_2_root_r119_carry_6_) );
  XOR2X1 U293 ( .A(in_17bit_b[0]), .B(in_17bit_b[1]), .Y(
        add_2_root_r119_SUM_5_) );
  AND2X1 U294 ( .A(add_1_root_r119_carry[22]), .B(n36), .Y(
        add_1_root_r119_SUM_23_) );
  XOR2X1 U295 ( .A(n36), .B(add_1_root_r119_carry[22]), .Y(
        add_1_root_r119_SUM_22_) );
  AND2X1 U296 ( .A(add_1_root_r119_carry[21]), .B(in_17bit_b[15]), .Y(
        add_1_root_r119_carry[22]) );
  XOR2X1 U297 ( .A(in_17bit_b[15]), .B(add_1_root_r119_carry[21]), .Y(
        add_1_root_r119_SUM_21_) );
  AND2X1 U298 ( .A(add_1_root_r119_carry[20]), .B(in_17bit_b[14]), .Y(
        add_1_root_r119_carry[21]) );
  XOR2X1 U299 ( .A(in_17bit_b[14]), .B(add_1_root_r119_carry[20]), .Y(
        add_1_root_r119_SUM_20_) );
  AND2X1 U300 ( .A(add_1_root_r119_A_6_), .B(in_17bit_b[0]), .Y(
        add_1_root_r119_carry[7]) );
  XOR2X1 U301 ( .A(in_17bit_b[0]), .B(add_1_root_r119_A_6_), .Y(
        add_1_root_r119_SUM_6_) );
  AND2X1 U302 ( .A(add_3_root_r119_carry_18_), .B(n36), .Y(
        add_1_root_r119_A_19_) );
  XOR2X1 U303 ( .A(n36), .B(add_3_root_r119_carry_18_), .Y(
        add_1_root_r119_A_18_) );
  AND2X1 U304 ( .A(in_17bit_b[1]), .B(in_17bit_b[0]), .Y(
        add_3_root_r119_carry_3_) );
  XOR2X1 U305 ( .A(in_17bit_b[0]), .B(in_17bit_b[1]), .Y(add_1_root_r119_A_2_)
         );
  AND2X1 U306 ( .A(add_2_root_r115_carry_19_), .B(n36), .Y(
        add_2_root_r115_SUM_20_) );
  XOR2X1 U307 ( .A(n36), .B(add_2_root_r115_carry_19_), .Y(
        add_2_root_r115_SUM_19_) );
  AND2X1 U308 ( .A(add_2_root_r115_carry_18_), .B(in_17bit_b[15]), .Y(
        add_2_root_r115_carry_19_) );
  XOR2X1 U309 ( .A(in_17bit_b[15]), .B(add_2_root_r115_carry_18_), .Y(
        add_2_root_r115_SUM_18_) );
  AND2X1 U310 ( .A(in_17bit_b[2]), .B(in_17bit_b[0]), .Y(
        add_2_root_r115_carry_4_) );
  XOR2X1 U311 ( .A(in_17bit_b[0]), .B(in_17bit_b[2]), .Y(
        add_2_root_r115_SUM_3_) );
  AND2X1 U312 ( .A(add_1_root_r115_carry_22_), .B(n36), .Y(
        add_1_root_r115_SUM_23_) );
  XOR2X1 U313 ( .A(n36), .B(add_1_root_r115_carry_22_), .Y(
        add_1_root_r115_SUM_22_) );
  AND2X1 U314 ( .A(add_1_root_r115_carry_21_), .B(in_17bit_b[15]), .Y(
        add_1_root_r115_carry_22_) );
  XOR2X1 U315 ( .A(in_17bit_b[15]), .B(add_1_root_r115_carry_21_), .Y(
        add_1_root_r115_SUM_21_) );
  AND2X1 U316 ( .A(in_17bit_b[2]), .B(in_17bit_b[0]), .Y(
        add_1_root_r115_carry_7_) );
  XOR2X1 U317 ( .A(in_17bit_b[0]), .B(in_17bit_b[2]), .Y(
        add_1_root_r115_SUM_6_) );
  XOR2X1 U318 ( .A(n89), .B(sub_add_54_b0_carry[15]), .Y(N28) );
  AND2X1 U319 ( .A(sub_add_54_b0_carry[14]), .B(n88), .Y(
        sub_add_54_b0_carry[15]) );
  XOR2X1 U320 ( .A(n88), .B(sub_add_54_b0_carry[14]), .Y(N27) );
  AND2X1 U321 ( .A(sub_add_54_b0_carry[13]), .B(n87), .Y(
        sub_add_54_b0_carry[14]) );
  XOR2X1 U322 ( .A(n87), .B(sub_add_54_b0_carry[13]), .Y(N26) );
  AND2X1 U323 ( .A(sub_add_54_b0_carry[12]), .B(n86), .Y(
        sub_add_54_b0_carry[13]) );
  XOR2X1 U324 ( .A(n86), .B(sub_add_54_b0_carry[12]), .Y(N25) );
  AND2X1 U325 ( .A(sub_add_54_b0_carry[11]), .B(n85), .Y(
        sub_add_54_b0_carry[12]) );
  XOR2X1 U326 ( .A(n85), .B(sub_add_54_b0_carry[11]), .Y(N24) );
  AND2X1 U327 ( .A(sub_add_54_b0_carry[10]), .B(n84), .Y(
        sub_add_54_b0_carry[11]) );
  XOR2X1 U328 ( .A(n84), .B(sub_add_54_b0_carry[10]), .Y(N23) );
  AND2X1 U329 ( .A(sub_add_54_b0_carry[9]), .B(n83), .Y(
        sub_add_54_b0_carry[10]) );
  XOR2X1 U330 ( .A(n83), .B(sub_add_54_b0_carry[9]), .Y(N22) );
  AND2X1 U331 ( .A(sub_add_54_b0_carry[8]), .B(n82), .Y(sub_add_54_b0_carry[9]) );
  XOR2X1 U332 ( .A(n82), .B(sub_add_54_b0_carry[8]), .Y(N21) );
  AND2X1 U333 ( .A(sub_add_54_b0_carry[7]), .B(n81), .Y(sub_add_54_b0_carry[8]) );
  XOR2X1 U334 ( .A(n81), .B(sub_add_54_b0_carry[7]), .Y(N20) );
  AND2X1 U335 ( .A(sub_add_54_b0_carry[6]), .B(n80), .Y(sub_add_54_b0_carry[7]) );
  XOR2X1 U336 ( .A(n80), .B(sub_add_54_b0_carry[6]), .Y(N19) );
  AND2X1 U337 ( .A(sub_add_54_b0_carry[5]), .B(n79), .Y(sub_add_54_b0_carry[6]) );
  XOR2X1 U338 ( .A(n79), .B(sub_add_54_b0_carry[5]), .Y(N18) );
  AND2X1 U339 ( .A(sub_add_54_b0_carry[4]), .B(n78), .Y(sub_add_54_b0_carry[5]) );
  XOR2X1 U340 ( .A(n78), .B(sub_add_54_b0_carry[4]), .Y(N17) );
  AND2X1 U341 ( .A(sub_add_54_b0_carry[3]), .B(n77), .Y(sub_add_54_b0_carry[4]) );
  XOR2X1 U342 ( .A(n77), .B(sub_add_54_b0_carry[3]), .Y(N16) );
  AND2X1 U343 ( .A(sub_add_54_b0_carry[2]), .B(n76), .Y(sub_add_54_b0_carry[3]) );
  XOR2X1 U344 ( .A(n76), .B(sub_add_54_b0_carry[2]), .Y(N15) );
  AND2X1 U345 ( .A(n74), .B(n75), .Y(sub_add_54_b0_carry[2]) );
  XOR2X1 U346 ( .A(n75), .B(n74), .Y(N14) );
  XOR2X1 U347 ( .A(n14), .B(sub_add_75_b0_carry[16]), .Y(N481) );
  AND2X1 U348 ( .A(sub_add_75_b0_carry[15]), .B(n8), .Y(
        sub_add_75_b0_carry[16]) );
  XOR2X1 U349 ( .A(n8), .B(sub_add_75_b0_carry[15]), .Y(N480) );
  AND2X1 U350 ( .A(sub_add_75_b0_carry[14]), .B(n9), .Y(
        sub_add_75_b0_carry[15]) );
  XOR2X1 U351 ( .A(n9), .B(sub_add_75_b0_carry[14]), .Y(N479) );
  AND2X1 U352 ( .A(sub_add_75_b0_carry[13]), .B(n10), .Y(
        sub_add_75_b0_carry[14]) );
  XOR2X1 U353 ( .A(n10), .B(sub_add_75_b0_carry[13]), .Y(N478) );
  AND2X1 U354 ( .A(sub_add_75_b0_carry[12]), .B(n11), .Y(
        sub_add_75_b0_carry[13]) );
  XOR2X1 U355 ( .A(n11), .B(sub_add_75_b0_carry[12]), .Y(N477) );
  AND2X1 U356 ( .A(sub_add_75_b0_carry[11]), .B(n12), .Y(
        sub_add_75_b0_carry[12]) );
  XOR2X1 U357 ( .A(n12), .B(sub_add_75_b0_carry[11]), .Y(N476) );
  AND2X1 U358 ( .A(sub_add_75_b0_carry[10]), .B(n13), .Y(
        sub_add_75_b0_carry[11]) );
  AND2X1 U359 ( .A(n27), .B(n7), .Y(sub_add_75_b0_carry[10]) );
  AND2X1 U360 ( .A(in_17bit_b[0]), .B(in_17bit_b[4]), .Y(
        add_1_root_r112_carry_5_) );
endmodule


module multi16_8_DW01_add_0 ( A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, 
        A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, 
        A_4_, B_23_, B_22_, B_21_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, 
        B_14_, B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, 
        SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, 
        SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, 
        SUM_7_ );
  input A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_,
         A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, B_23_, B_22_,
         B_21_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_,
         B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_;
  output SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_,
         SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_,
         SUM_8_, SUM_7_;
  wire   n1, n2, n3, n4;
  wire   [23:7] carry;

  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry[7]), .CO(carry[8]), .S(SUM_7_)
         );
  ADDFX2 U1_21 ( .A(A_21_), .B(B_21_), .CI(carry[21]), .CO(carry[22]), .S(
        SUM_21_) );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry[20]), .CO(carry[21]), .S(
        SUM_20_) );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry[19]), .CO(carry[20]), .S(
        SUM_19_) );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry[18]), .CO(carry[19]), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry[17]), .CO(carry[18]), .S(
        SUM_17_) );
  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry[16]), .CO(carry[17]), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry[15]), .CO(carry[16]), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry[14]), .CO(carry[15]), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry[13]), .CO(carry[14]), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry[12]), .CO(carry[13]), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry[11]), .CO(carry[12]), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry[10]), .CO(carry[11]), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry[9]), .CO(carry[10]), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry[8]), .CO(carry[9]), .S(SUM_8_)
         );
  ADDFX2 U1_22 ( .A(A_22_), .B(B_22_), .CI(carry[22]), .CO(carry[23]), .S(
        SUM_22_) );
  AND2X2 U1 ( .A(A_4_), .B(B_4_), .Y(n1) );
  XOR2X1 U2 ( .A(B_23_), .B(carry[23]), .Y(SUM_23_) );
  OAI2BB1X1 U3 ( .A0N(n2), .A1N(A_6_), .B0(n3), .Y(carry[7]) );
  OAI21XL U4 ( .A0(A_6_), .A1(n2), .B0(B_6_), .Y(n3) );
  OAI2BB1X1 U5 ( .A0N(n1), .A1N(A_5_), .B0(n4), .Y(n2) );
  OAI21XL U6 ( .A0(A_5_), .A1(n1), .B0(B_5_), .Y(n4) );
endmodule


module multi16_8_DW01_add_4 ( A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, 
        A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, 
        B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, 
        B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, SUM_22_, SUM_21_, SUM_20_, 
        SUM_19_, SUM_18_, SUM_17_, SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, 
        SUM_11_, SUM_10_, SUM_9_, SUM_8_, SUM_7_ );
  input A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_,
         A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, B_20_, B_19_,
         B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, B_10_, B_9_,
         B_8_, B_7_, B_6_, B_5_;
  output SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_,
         SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_,
         SUM_7_;
  wire   carry_21_, carry_20_, carry_19_, carry_18_, carry_17_, carry_16_,
         carry_15_, carry_14_, carry_13_, carry_12_, carry_11_, carry_10_,
         carry_9_, carry_8_, carry_7_, n1;

  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry_16_), .CO(carry_17_), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry_15_), .CO(carry_16_), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry_14_), .CO(carry_15_), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry_13_), .CO(carry_14_), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry_12_), .CO(carry_13_), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry_11_), .CO(carry_12_), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry_10_), .CO(carry_11_), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry_9_), .CO(carry_10_), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry_8_), .CO(carry_9_), .S(SUM_8_)
         );
  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry_7_), .CO(carry_8_), .S(SUM_7_)
         );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry_20_), .CO(carry_21_), .S(
        SUM_20_) );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry_19_), .CO(carry_20_), .S(
        SUM_19_) );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry_18_), .CO(carry_19_), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry_17_), .CO(carry_18_), .S(
        SUM_17_) );
  ADDFX2 U1_21 ( .A(A_21_), .B(B_21_), .CI(carry_21_), .CO(SUM_22_), .S(
        SUM_21_) );
  OAI2BB1X1 U1 ( .A0N(A_6_), .A1N(B_6_), .B0(n1), .Y(carry_7_) );
  OAI211X1 U2 ( .A0(B_6_), .A1(A_6_), .B0(A_5_), .C0(B_5_), .Y(n1) );
endmodule


module multi16_8_DW01_add_6 ( A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, 
        A_16_, A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, 
        A_6_, A_5_, A_4_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, 
        B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, 
        SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, 
        SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, 
        SUM_7_ );
  input A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_,
         A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, B_20_,
         B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, B_10_,
         B_9_, B_8_, B_7_, B_6_, B_5_, B_4_;
  output SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_,
         SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_,
         SUM_8_, SUM_7_;
  wire   n1, n2, n3, n4, n5, n6;
  wire   [21:7] carry;

  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry[7]), .CO(carry[8]), .S(SUM_7_)
         );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry[18]), .CO(carry[19]), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry[17]), .CO(carry[18]), .S(
        SUM_17_) );
  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry[16]), .CO(carry[17]), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry[15]), .CO(carry[16]), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry[14]), .CO(carry[15]), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry[13]), .CO(carry[14]), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry[12]), .CO(carry[13]), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry[11]), .CO(carry[12]), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry[10]), .CO(carry[11]), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry[9]), .CO(carry[10]), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry[8]), .CO(carry[9]), .S(SUM_8_)
         );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry[19]), .CO(carry[20]), .S(
        SUM_19_) );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry[20]), .CO(carry[21]), .S(
        SUM_20_) );
  AND2X2 U1 ( .A(A_22_), .B(n2), .Y(n1) );
  AND2X2 U2 ( .A(A_21_), .B(carry[21]), .Y(n2) );
  XOR2X1 U3 ( .A(A_23_), .B(n1), .Y(SUM_23_) );
  AND2X2 U4 ( .A(A_4_), .B(B_4_), .Y(n3) );
  XOR2X1 U5 ( .A(A_21_), .B(carry[21]), .Y(SUM_21_) );
  XOR2X1 U6 ( .A(A_22_), .B(n2), .Y(SUM_22_) );
  OAI2BB1X1 U7 ( .A0N(n4), .A1N(A_6_), .B0(n5), .Y(carry[7]) );
  OAI21XL U8 ( .A0(A_6_), .A1(n4), .B0(B_6_), .Y(n5) );
  OAI2BB1X1 U9 ( .A0N(n3), .A1N(A_5_), .B0(n6), .Y(n4) );
  OAI21XL U10 ( .A0(A_5_), .A1(n3), .B0(B_5_), .Y(n6) );
endmodule


module multi16_8 ( in_17bit, in_8bit, out );
  input [16:0] in_17bit;
  input [7:0] in_8bit;
  output [16:0] out;
  wire   N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27,
         N28, N29, N108, N109, N110, N111, N112, N113, N114, N115, N116, N117,
         N118, N119, N120, N121, N122, N123, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220,
         N221, N347, N348, N349, N350, N351, N352, N353, N354, N355, N356,
         N357, N358, N359, N360, N361, N362, N363, N446, N447, N448, N449,
         N450, N451, N452, N453, N454, N455, N456, N457, N458, N459, N460,
         N461, N462, N463, N477, N478, N479, N480, add_2_root_r119_carry_10_,
         add_2_root_r119_carry_11_, add_2_root_r119_carry_12_,
         add_2_root_r119_carry_13_, add_2_root_r119_carry_14_,
         add_2_root_r119_carry_15_, add_2_root_r119_carry_16_,
         add_2_root_r119_carry_17_, add_2_root_r119_carry_18_,
         add_2_root_r119_carry_19_, add_2_root_r119_carry_20_,
         add_2_root_r119_carry_21_, add_2_root_r119_carry_6_,
         add_2_root_r119_carry_7_, add_2_root_r119_carry_8_,
         add_2_root_r119_carry_9_, add_2_root_r119_SUM_5_,
         add_2_root_r119_SUM_6_, add_2_root_r119_SUM_7_,
         add_2_root_r119_SUM_8_, add_2_root_r119_SUM_9_,
         add_2_root_r119_SUM_10_, add_2_root_r119_SUM_11_,
         add_2_root_r119_SUM_12_, add_2_root_r119_SUM_13_,
         add_2_root_r119_SUM_14_, add_2_root_r119_SUM_15_,
         add_2_root_r119_SUM_16_, add_2_root_r119_SUM_17_,
         add_2_root_r119_SUM_18_, add_2_root_r119_SUM_19_,
         add_2_root_r119_SUM_20_, add_2_root_r119_SUM_21_,
         add_2_root_r119_SUM_22_, add_1_root_r119_SUM_6_,
         add_1_root_r119_SUM_7_, add_1_root_r119_SUM_8_,
         add_1_root_r119_SUM_9_, add_1_root_r119_SUM_10_,
         add_1_root_r119_SUM_11_, add_1_root_r119_SUM_12_,
         add_1_root_r119_SUM_13_, add_1_root_r119_SUM_14_,
         add_1_root_r119_SUM_15_, add_1_root_r119_SUM_16_,
         add_1_root_r119_SUM_17_, add_1_root_r119_SUM_18_,
         add_1_root_r119_SUM_19_, add_1_root_r119_SUM_20_,
         add_1_root_r119_SUM_21_, add_1_root_r119_SUM_22_,
         add_1_root_r119_SUM_23_, add_1_root_r119_A_2_, add_1_root_r119_A_3_,
         add_1_root_r119_A_4_, add_1_root_r119_A_5_, add_1_root_r119_A_6_,
         add_1_root_r119_A_7_, add_1_root_r119_A_8_, add_1_root_r119_A_9_,
         add_1_root_r119_A_10_, add_1_root_r119_A_11_, add_1_root_r119_A_12_,
         add_1_root_r119_A_13_, add_1_root_r119_A_14_, add_1_root_r119_A_15_,
         add_1_root_r119_A_16_, add_1_root_r119_A_17_, add_1_root_r119_A_18_,
         add_1_root_r119_A_19_, add_3_root_r119_carry_10_,
         add_3_root_r119_carry_11_, add_3_root_r119_carry_12_,
         add_3_root_r119_carry_13_, add_3_root_r119_carry_14_,
         add_3_root_r119_carry_15_, add_3_root_r119_carry_16_,
         add_3_root_r119_carry_17_, add_3_root_r119_carry_18_,
         add_3_root_r119_carry_3_, add_3_root_r119_carry_4_,
         add_3_root_r119_carry_5_, add_3_root_r119_carry_6_,
         add_3_root_r119_carry_7_, add_3_root_r119_carry_8_,
         add_3_root_r119_carry_9_, add_1_root_r112_carry_10_,
         add_1_root_r112_carry_11_, add_1_root_r112_carry_12_,
         add_1_root_r112_carry_13_, add_1_root_r112_carry_14_,
         add_1_root_r112_carry_15_, add_1_root_r112_carry_16_,
         add_1_root_r112_carry_17_, add_1_root_r112_carry_18_,
         add_1_root_r112_carry_19_, add_1_root_r112_carry_20_,
         add_1_root_r112_carry_5_, add_1_root_r112_carry_6_,
         add_1_root_r112_carry_7_, add_1_root_r112_carry_8_,
         add_1_root_r112_carry_9_, add_1_root_r112_SUM_1_,
         add_1_root_r112_SUM_2_, add_1_root_r112_SUM_3_,
         add_1_root_r112_SUM_4_, add_1_root_r112_SUM_5_,
         add_1_root_r112_SUM_6_, add_1_root_r112_SUM_7_,
         add_1_root_r112_SUM_8_, add_1_root_r112_SUM_9_,
         add_1_root_r112_SUM_10_, add_1_root_r112_SUM_11_,
         add_1_root_r112_SUM_12_, add_1_root_r112_SUM_13_,
         add_1_root_r112_SUM_14_, add_1_root_r112_SUM_15_,
         add_1_root_r112_SUM_16_, add_1_root_r112_SUM_17_,
         add_1_root_r112_SUM_18_, add_1_root_r112_SUM_19_,
         add_1_root_r112_SUM_20_, add_1_root_r112_SUM_21_,
         add_2_root_r115_carry_10_, add_2_root_r115_carry_11_,
         add_2_root_r115_carry_12_, add_2_root_r115_carry_13_,
         add_2_root_r115_carry_14_, add_2_root_r115_carry_15_,
         add_2_root_r115_carry_16_, add_2_root_r115_carry_17_,
         add_2_root_r115_carry_18_, add_2_root_r115_carry_19_,
         add_2_root_r115_carry_4_, add_2_root_r115_carry_5_,
         add_2_root_r115_carry_6_, add_2_root_r115_carry_7_,
         add_2_root_r115_carry_8_, add_2_root_r115_carry_9_,
         add_2_root_r115_SUM_3_, add_2_root_r115_SUM_4_,
         add_2_root_r115_SUM_5_, add_2_root_r115_SUM_6_,
         add_2_root_r115_SUM_7_, add_2_root_r115_SUM_8_,
         add_2_root_r115_SUM_9_, add_2_root_r115_SUM_10_,
         add_2_root_r115_SUM_11_, add_2_root_r115_SUM_12_,
         add_2_root_r115_SUM_13_, add_2_root_r115_SUM_14_,
         add_2_root_r115_SUM_15_, add_2_root_r115_SUM_16_,
         add_2_root_r115_SUM_17_, add_2_root_r115_SUM_18_,
         add_2_root_r115_SUM_19_, add_2_root_r115_SUM_20_,
         add_1_root_r115_carry_10_, add_1_root_r115_carry_11_,
         add_1_root_r115_carry_12_, add_1_root_r115_carry_13_,
         add_1_root_r115_carry_14_, add_1_root_r115_carry_15_,
         add_1_root_r115_carry_16_, add_1_root_r115_carry_17_,
         add_1_root_r115_carry_18_, add_1_root_r115_carry_19_,
         add_1_root_r115_carry_20_, add_1_root_r115_carry_21_,
         add_1_root_r115_carry_22_, add_1_root_r115_carry_7_,
         add_1_root_r115_carry_8_, add_1_root_r115_carry_9_,
         add_1_root_r115_SUM_6_, add_1_root_r115_SUM_7_,
         add_1_root_r115_SUM_8_, add_1_root_r115_SUM_9_,
         add_1_root_r115_SUM_10_, add_1_root_r115_SUM_11_,
         add_1_root_r115_SUM_12_, add_1_root_r115_SUM_13_,
         add_1_root_r115_SUM_14_, add_1_root_r115_SUM_15_,
         add_1_root_r115_SUM_16_, add_1_root_r115_SUM_17_,
         add_1_root_r115_SUM_18_, add_1_root_r115_SUM_19_,
         add_1_root_r115_SUM_20_, add_1_root_r115_SUM_21_,
         add_1_root_r115_SUM_22_, add_1_root_r115_SUM_23_, n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245;
  wire   [16:0] in_17bit_b;
  wire   [23:8] neg_mul;
  wire   [15:10] sub_add_75_b0_carry;
  wire   [16:2] sub_add_54_b0_carry;
  wire   [22:7] add_1_root_r119_carry;

  multi16_8_DW01_add_0 add_0_root_r119 ( .A_22_(add_2_root_r119_SUM_22_), 
        .A_21_(add_2_root_r119_SUM_21_), .A_20_(add_2_root_r119_SUM_20_), 
        .A_19_(add_2_root_r119_SUM_19_), .A_18_(add_2_root_r119_SUM_18_), 
        .A_17_(add_2_root_r119_SUM_17_), .A_16_(add_2_root_r119_SUM_16_), 
        .A_15_(add_2_root_r119_SUM_15_), .A_14_(add_2_root_r119_SUM_14_), 
        .A_13_(add_2_root_r119_SUM_13_), .A_12_(add_2_root_r119_SUM_12_), 
        .A_11_(add_2_root_r119_SUM_11_), .A_10_(add_2_root_r119_SUM_10_), 
        .A_9_(add_2_root_r119_SUM_9_), .A_8_(add_2_root_r119_SUM_8_), .A_7_(
        add_2_root_r119_SUM_7_), .A_6_(add_2_root_r119_SUM_6_), .A_5_(
        add_2_root_r119_SUM_5_), .A_4_(in_17bit_b[0]), .B_23_(
        add_1_root_r119_SUM_23_), .B_22_(add_1_root_r119_SUM_22_), .B_21_(
        add_1_root_r119_SUM_21_), .B_20_(add_1_root_r119_SUM_20_), .B_19_(
        add_1_root_r119_SUM_19_), .B_18_(add_1_root_r119_SUM_18_), .B_17_(
        add_1_root_r119_SUM_17_), .B_16_(add_1_root_r119_SUM_16_), .B_15_(
        add_1_root_r119_SUM_15_), .B_14_(add_1_root_r119_SUM_14_), .B_13_(
        add_1_root_r119_SUM_13_), .B_12_(add_1_root_r119_SUM_12_), .B_11_(
        add_1_root_r119_SUM_11_), .B_10_(add_1_root_r119_SUM_10_), .B_9_(
        add_1_root_r119_SUM_9_), .B_8_(add_1_root_r119_SUM_8_), .B_7_(
        add_1_root_r119_SUM_7_), .B_6_(add_1_root_r119_SUM_6_), .B_5_(
        add_1_root_r119_A_5_), .B_4_(add_1_root_r119_A_4_), .SUM_23_(N363), 
        .SUM_22_(N362), .SUM_21_(N361), .SUM_20_(N360), .SUM_19_(N359), 
        .SUM_18_(N358), .SUM_17_(N357), .SUM_16_(N356), .SUM_15_(N355), 
        .SUM_14_(N354), .SUM_13_(N353), .SUM_12_(N352), .SUM_11_(N351), 
        .SUM_10_(N350), .SUM_9_(N349), .SUM_8_(N348), .SUM_7_(N347) );
  multi16_8_DW01_add_4 add_0_root_r112 ( .A_21_(n37), .A_20_(in_17bit_b[15]), 
        .A_19_(in_17bit_b[14]), .A_18_(in_17bit_b[13]), .A_17_(in_17bit_b[12]), 
        .A_16_(in_17bit_b[11]), .A_15_(in_17bit_b[10]), .A_14_(in_17bit_b[9]), 
        .A_13_(in_17bit_b[8]), .A_12_(in_17bit_b[7]), .A_11_(in_17bit_b[6]), 
        .A_10_(in_17bit_b[5]), .A_9_(in_17bit_b[4]), .A_8_(in_17bit_b[3]), 
        .A_7_(in_17bit_b[2]), .A_6_(in_17bit_b[1]), .A_5_(in_17bit_b[0]), 
        .B_21_(add_1_root_r112_SUM_21_), .B_20_(add_1_root_r112_SUM_20_), 
        .B_19_(add_1_root_r112_SUM_19_), .B_18_(add_1_root_r112_SUM_18_), 
        .B_17_(add_1_root_r112_SUM_17_), .B_16_(add_1_root_r112_SUM_16_), 
        .B_15_(add_1_root_r112_SUM_15_), .B_14_(add_1_root_r112_SUM_14_), 
        .B_13_(add_1_root_r112_SUM_13_), .B_12_(add_1_root_r112_SUM_12_), 
        .B_11_(add_1_root_r112_SUM_11_), .B_10_(add_1_root_r112_SUM_10_), 
        .B_9_(add_1_root_r112_SUM_9_), .B_8_(add_1_root_r112_SUM_8_), .B_7_(
        add_1_root_r112_SUM_7_), .B_6_(add_1_root_r112_SUM_6_), .B_5_(
        add_1_root_r112_SUM_5_), .SUM_22_(N123), .SUM_21_(N122), .SUM_20_(N121), .SUM_19_(N120), .SUM_18_(N119), .SUM_17_(N118), .SUM_16_(N117), .SUM_15_(
        N116), .SUM_14_(N115), .SUM_13_(N114), .SUM_12_(N113), .SUM_11_(N112), 
        .SUM_10_(N111), .SUM_9_(N110), .SUM_8_(N109), .SUM_7_(N108) );
  multi16_8_DW01_add_6 add_0_root_r115 ( .A_23_(add_1_root_r115_SUM_23_), 
        .A_22_(add_1_root_r115_SUM_22_), .A_21_(add_1_root_r115_SUM_21_), 
        .A_20_(add_1_root_r115_SUM_20_), .A_19_(add_1_root_r115_SUM_19_), 
        .A_18_(add_1_root_r115_SUM_18_), .A_17_(add_1_root_r115_SUM_17_), 
        .A_16_(add_1_root_r115_SUM_16_), .A_15_(add_1_root_r115_SUM_15_), 
        .A_14_(add_1_root_r115_SUM_14_), .A_13_(add_1_root_r115_SUM_13_), 
        .A_12_(add_1_root_r115_SUM_12_), .A_11_(add_1_root_r115_SUM_11_), 
        .A_10_(add_1_root_r115_SUM_10_), .A_9_(add_1_root_r115_SUM_9_), .A_8_(
        add_1_root_r115_SUM_8_), .A_7_(add_1_root_r115_SUM_7_), .A_6_(
        add_1_root_r115_SUM_6_), .A_5_(in_17bit_b[1]), .A_4_(in_17bit_b[0]), 
        .B_20_(add_2_root_r115_SUM_20_), .B_19_(add_2_root_r115_SUM_19_), 
        .B_18_(add_2_root_r115_SUM_18_), .B_17_(add_2_root_r115_SUM_17_), 
        .B_16_(add_2_root_r115_SUM_16_), .B_15_(add_2_root_r115_SUM_15_), 
        .B_14_(add_2_root_r115_SUM_14_), .B_13_(add_2_root_r115_SUM_13_), 
        .B_12_(add_2_root_r115_SUM_12_), .B_11_(add_2_root_r115_SUM_11_), 
        .B_10_(add_2_root_r115_SUM_10_), .B_9_(add_2_root_r115_SUM_9_), .B_8_(
        add_2_root_r115_SUM_8_), .B_7_(add_2_root_r115_SUM_7_), .B_6_(
        add_2_root_r115_SUM_6_), .B_5_(add_2_root_r115_SUM_5_), .B_4_(
        add_2_root_r115_SUM_4_), .SUM_23_(N221), .SUM_22_(N220), .SUM_21_(N219), .SUM_20_(N218), .SUM_19_(N217), .SUM_18_(N216), .SUM_17_(N215), .SUM_16_(
        N214), .SUM_15_(N213), .SUM_14_(N212), .SUM_13_(N211), .SUM_12_(N210), 
        .SUM_11_(N209), .SUM_10_(N208), .SUM_9_(N207), .SUM_8_(N206), .SUM_7_(
        N205) );
  TLATX1 neg_mul_reg_16_ ( .G(N446), .D(N456), .QN(n8) );
  TLATX1 neg_mul_reg_15_ ( .G(N446), .D(N455), .QN(n3) );
  TLATX1 neg_mul_reg_14_ ( .G(N446), .D(N454), .QN(n7) );
  TLATX1 neg_mul_reg_13_ ( .G(N446), .D(N453), .QN(n6) );
  TLATX1 neg_mul_reg_12_ ( .G(N446), .D(N452), .QN(n5) );
  TLATX1 neg_mul_reg_11_ ( .G(N446), .D(N451), .QN(n4) );
  TLATX1 neg_mul_reg_10_ ( .G(N446), .D(N450), .QN(n2) );
  TLATX1 neg_mul_reg_9_ ( .G(N446), .D(N449), .Q(neg_mul[9]), .QN(n15) );
  TLATX1 neg_mul_reg_23_ ( .G(N446), .D(N463), .Q(neg_mul[23]), .QN(n1) );
  TLATX1 neg_mul_reg_22_ ( .G(N446), .D(N462), .Q(neg_mul[22]), .QN(n9) );
  TLATX1 neg_mul_reg_21_ ( .G(N446), .D(N461), .Q(neg_mul[21]), .QN(n11) );
  TLATX1 neg_mul_reg_20_ ( .G(N446), .D(N460), .Q(neg_mul[20]), .QN(n12) );
  TLATX1 neg_mul_reg_19_ ( .G(N446), .D(N459), .Q(neg_mul[19]), .QN(n10) );
  TLATX1 neg_mul_reg_18_ ( .G(N446), .D(N458), .QN(n13) );
  TLATX1 neg_mul_reg_17_ ( .G(N446), .D(N457), .QN(n16) );
  TLATX1 neg_mul_reg_8_ ( .G(N446), .D(N448), .Q(neg_mul[8]) );
  TLATX1 neg_mul_reg_7_ ( .G(N446), .D(N447), .Q(out[0]), .QN(n14) );
  NOR2X4 U2 ( .A(n60), .B(n52), .Y(n61) );
  OR2X4 U3 ( .A(n52), .B(n29), .Y(n18) );
  INVX8 U4 ( .A(in_8bit[7]), .Y(n42) );
  NAND4XL U5 ( .A(in_8bit[1]), .B(in_8bit[7]), .C(n182), .D(n98), .Y(n183) );
  XNOR2X1 U6 ( .A(neg_mul[23]), .B(n34), .Y(n17) );
  INVX20 U7 ( .A(n52), .Y(n66) );
  XNOR2X4 U8 ( .A(in_8bit[7]), .B(n45), .Y(n65) );
  XOR2X4 U9 ( .A(n18), .B(n3), .Y(out[8]) );
  CLKINVX3 U10 ( .A(in_17bit[16]), .Y(n19) );
  INVX4 U11 ( .A(in_17bit[16]), .Y(n47) );
  XOR2X4 U12 ( .A(n20), .B(n8), .Y(out[9]) );
  OR2X4 U13 ( .A(n30), .B(n65), .Y(n20) );
  NOR2X4 U14 ( .A(n28), .B(n21), .Y(n64) );
  XOR2X4 U15 ( .A(n55), .B(neg_mul[9]), .Y(out[2]) );
  NOR2X2 U16 ( .A(n57), .B(n14), .Y(n53) );
  XOR2X4 U17 ( .A(n42), .B(n45), .Y(n21) );
  NOR2X4 U18 ( .A(n26), .B(n65), .Y(n62) );
  MX2X4 U19 ( .A(neg_mul[19]), .B(N477), .S0(n66), .Y(out[12]) );
  XOR2X4 U20 ( .A(n42), .B(n45), .Y(n52) );
  NAND2X4 U21 ( .A(n16), .B(n22), .Y(n23) );
  NAND2X2 U22 ( .A(n32), .B(n66), .Y(n24) );
  NAND2X4 U23 ( .A(n23), .B(n24), .Y(n25) );
  INVX2 U24 ( .A(n66), .Y(n22) );
  INVX8 U25 ( .A(n25), .Y(out[10]) );
  INVX8 U26 ( .A(n47), .Y(n45) );
  NAND3XL U27 ( .A(in_8bit[7]), .B(n40), .C(n44), .Y(n76) );
  INVXL U28 ( .A(n45), .Y(n36) );
  INVX1 U29 ( .A(n195), .Y(in_17bit_b[1]) );
  INVX1 U30 ( .A(n234), .Y(in_17bit_b[14]) );
  INVX1 U31 ( .A(n231), .Y(in_17bit_b[13]) );
  INVX1 U32 ( .A(n198), .Y(in_17bit_b[2]) );
  INVX1 U33 ( .A(n207), .Y(in_17bit_b[5]) );
  INVX1 U34 ( .A(n210), .Y(in_17bit_b[6]) );
  INVX1 U35 ( .A(n213), .Y(in_17bit_b[7]) );
  INVX1 U36 ( .A(n204), .Y(in_17bit_b[4]) );
  INVX1 U37 ( .A(n216), .Y(in_17bit_b[8]) );
  INVX1 U38 ( .A(n219), .Y(in_17bit_b[9]) );
  INVX1 U39 ( .A(n222), .Y(in_17bit_b[10]) );
  INVX1 U40 ( .A(n225), .Y(in_17bit_b[11]) );
  INVX1 U41 ( .A(n228), .Y(in_17bit_b[12]) );
  INVX1 U42 ( .A(n201), .Y(in_17bit_b[3]) );
  MX2X1 U43 ( .A(neg_mul[20]), .B(N478), .S0(n66), .Y(out[13]) );
  INVX1 U44 ( .A(n36), .Y(n48) );
  INVX1 U45 ( .A(n46), .Y(n50) );
  INVX1 U46 ( .A(n46), .Y(n49) );
  NAND3X1 U47 ( .A(in_8bit[2]), .B(n41), .C(in_8bit[5]), .Y(n184) );
  NAND3BX1 U48 ( .AN(in_8bit[5]), .B(n43), .C(in_8bit[3]), .Y(n185) );
  INVX1 U49 ( .A(n39), .Y(n38) );
  INVX1 U50 ( .A(n97), .Y(n244) );
  OAI21XL U51 ( .A0(n244), .A1(n245), .B0(n243), .Y(N463) );
  AOI22X1 U52 ( .A0(N221), .A1(n242), .B0(N363), .B1(n241), .Y(n243) );
  ADDFX2 U53 ( .A(n37), .B(in_17bit_b[12]), .CI(add_1_root_r112_carry_16_), 
        .CO(add_1_root_r112_carry_17_), .S(add_1_root_r112_SUM_16_) );
  ADDFX2 U54 ( .A(add_1_root_r119_A_19_), .B(in_17bit_b[13]), .CI(
        add_1_root_r119_carry[19]), .CO(add_1_root_r119_carry[20]), .S(
        add_1_root_r119_SUM_19_) );
  ADDFX2 U55 ( .A(n37), .B(in_17bit_b[15]), .CI(add_3_root_r119_carry_17_), 
        .CO(add_3_root_r119_carry_18_), .S(add_1_root_r119_A_17_) );
  ADDFX2 U56 ( .A(n37), .B(in_17bit_b[14]), .CI(add_2_root_r115_carry_17_), 
        .CO(add_2_root_r115_carry_18_), .S(add_2_root_r115_SUM_17_) );
  ADDFX2 U57 ( .A(n37), .B(in_17bit_b[14]), .CI(add_1_root_r115_carry_20_), 
        .CO(add_1_root_r115_carry_21_), .S(add_1_root_r115_SUM_20_) );
  ADDFX2 U58 ( .A(n37), .B(in_17bit_b[15]), .CI(add_2_root_r119_carry_20_), 
        .CO(add_2_root_r119_carry_21_), .S(add_2_root_r119_SUM_20_) );
  ADDFX2 U59 ( .A(in_17bit_b[3]), .B(in_17bit_b[1]), .CI(
        add_2_root_r115_carry_4_), .CO(add_2_root_r115_carry_5_), .S(
        add_2_root_r115_SUM_4_) );
  ADDFX2 U60 ( .A(in_17bit_b[4]), .B(in_17bit_b[2]), .CI(
        add_2_root_r115_carry_5_), .CO(add_2_root_r115_carry_6_), .S(
        add_2_root_r115_SUM_5_) );
  ADDFX2 U61 ( .A(in_17bit_b[5]), .B(in_17bit_b[1]), .CI(
        add_1_root_r112_carry_5_), .CO(add_1_root_r112_carry_6_), .S(
        add_1_root_r112_SUM_5_) );
  ADDFX2 U62 ( .A(in_17bit_b[6]), .B(in_17bit_b[5]), .CI(
        add_3_root_r119_carry_7_), .CO(add_3_root_r119_carry_8_), .S(
        add_1_root_r119_A_7_) );
  ADDFX2 U63 ( .A(in_17bit_b[6]), .B(in_17bit_b[2]), .CI(
        add_1_root_r112_carry_6_), .CO(add_1_root_r112_carry_7_), .S(
        add_1_root_r112_SUM_6_) );
  ADDFX2 U64 ( .A(in_17bit_b[3]), .B(in_17bit_b[1]), .CI(
        add_1_root_r115_carry_7_), .CO(add_1_root_r115_carry_8_), .S(
        add_1_root_r115_SUM_7_) );
  ADDFX2 U65 ( .A(in_17bit_b[7]), .B(in_17bit_b[6]), .CI(
        add_3_root_r119_carry_8_), .CO(add_3_root_r119_carry_9_), .S(
        add_1_root_r119_A_8_) );
  ADDFX2 U66 ( .A(add_1_root_r119_A_7_), .B(in_17bit_b[1]), .CI(
        add_1_root_r119_carry[7]), .CO(add_1_root_r119_carry[8]), .S(
        add_1_root_r119_SUM_7_) );
  ADDFX2 U67 ( .A(in_17bit_b[2]), .B(in_17bit_b[1]), .CI(
        add_2_root_r119_carry_6_), .CO(add_2_root_r119_carry_7_), .S(
        add_2_root_r119_SUM_6_) );
  ADDFX2 U68 ( .A(in_17bit_b[4]), .B(in_17bit_b[2]), .CI(
        add_1_root_r115_carry_8_), .CO(add_1_root_r115_carry_9_), .S(
        add_1_root_r115_SUM_8_) );
  ADDFX2 U69 ( .A(in_17bit_b[8]), .B(in_17bit_b[7]), .CI(
        add_3_root_r119_carry_9_), .CO(add_3_root_r119_carry_10_), .S(
        add_1_root_r119_A_9_) );
  ADDFX2 U70 ( .A(add_1_root_r119_A_8_), .B(in_17bit_b[2]), .CI(
        add_1_root_r119_carry[8]), .CO(add_1_root_r119_carry[9]), .S(
        add_1_root_r119_SUM_8_) );
  ADDFX2 U71 ( .A(in_17bit_b[3]), .B(in_17bit_b[2]), .CI(
        add_2_root_r119_carry_7_), .CO(add_2_root_r119_carry_8_), .S(
        add_2_root_r119_SUM_7_) );
  ADDFX2 U72 ( .A(in_17bit_b[6]), .B(in_17bit_b[4]), .CI(
        add_2_root_r115_carry_7_), .CO(add_2_root_r115_carry_8_), .S(
        add_2_root_r115_SUM_7_) );
  ADDFX2 U73 ( .A(in_17bit_b[8]), .B(in_17bit_b[4]), .CI(
        add_1_root_r112_carry_8_), .CO(add_1_root_r112_carry_9_), .S(
        add_1_root_r112_SUM_8_) );
  ADDFX2 U74 ( .A(in_17bit_b[9]), .B(in_17bit_b[8]), .CI(
        add_3_root_r119_carry_10_), .CO(add_3_root_r119_carry_11_), .S(
        add_1_root_r119_A_10_) );
  ADDFX2 U75 ( .A(in_17bit_b[7]), .B(in_17bit_b[5]), .CI(
        add_2_root_r115_carry_8_), .CO(add_2_root_r115_carry_9_), .S(
        add_2_root_r115_SUM_8_) );
  ADDFX2 U76 ( .A(in_17bit_b[9]), .B(in_17bit_b[5]), .CI(
        add_1_root_r112_carry_9_), .CO(add_1_root_r112_carry_10_), .S(
        add_1_root_r112_SUM_9_) );
  ADDFX2 U77 ( .A(in_17bit_b[6]), .B(in_17bit_b[4]), .CI(
        add_1_root_r115_carry_10_), .CO(add_1_root_r115_carry_11_), .S(
        add_1_root_r115_SUM_10_) );
  ADDFX2 U78 ( .A(in_17bit_b[10]), .B(in_17bit_b[9]), .CI(
        add_3_root_r119_carry_11_), .CO(add_3_root_r119_carry_12_), .S(
        add_1_root_r119_A_11_) );
  ADDFX2 U79 ( .A(in_17bit_b[5]), .B(in_17bit_b[4]), .CI(
        add_2_root_r119_carry_9_), .CO(add_2_root_r119_carry_10_), .S(
        add_2_root_r119_SUM_9_) );
  ADDFX2 U80 ( .A(in_17bit_b[8]), .B(in_17bit_b[6]), .CI(
        add_2_root_r115_carry_9_), .CO(add_2_root_r115_carry_10_), .S(
        add_2_root_r115_SUM_9_) );
  ADDFX2 U81 ( .A(in_17bit_b[10]), .B(in_17bit_b[6]), .CI(
        add_1_root_r112_carry_10_), .CO(add_1_root_r112_carry_11_), .S(
        add_1_root_r112_SUM_10_) );
  ADDFX2 U82 ( .A(in_17bit_b[7]), .B(in_17bit_b[5]), .CI(
        add_1_root_r115_carry_11_), .CO(add_1_root_r115_carry_12_), .S(
        add_1_root_r115_SUM_11_) );
  ADDFX2 U83 ( .A(in_17bit_b[11]), .B(in_17bit_b[10]), .CI(
        add_3_root_r119_carry_12_), .CO(add_3_root_r119_carry_13_), .S(
        add_1_root_r119_A_12_) );
  ADDFX2 U84 ( .A(in_17bit_b[6]), .B(in_17bit_b[5]), .CI(
        add_2_root_r119_carry_10_), .CO(add_2_root_r119_carry_11_), .S(
        add_2_root_r119_SUM_10_) );
  ADDFX2 U85 ( .A(in_17bit_b[9]), .B(in_17bit_b[7]), .CI(
        add_2_root_r115_carry_10_), .CO(add_2_root_r115_carry_11_), .S(
        add_2_root_r115_SUM_10_) );
  ADDFX2 U86 ( .A(in_17bit_b[11]), .B(in_17bit_b[7]), .CI(
        add_1_root_r112_carry_11_), .CO(add_1_root_r112_carry_12_), .S(
        add_1_root_r112_SUM_11_) );
  ADDFX2 U87 ( .A(in_17bit_b[8]), .B(in_17bit_b[6]), .CI(
        add_1_root_r115_carry_12_), .CO(add_1_root_r115_carry_13_), .S(
        add_1_root_r115_SUM_12_) );
  ADDFX2 U88 ( .A(in_17bit_b[12]), .B(in_17bit_b[11]), .CI(
        add_3_root_r119_carry_13_), .CO(add_3_root_r119_carry_14_), .S(
        add_1_root_r119_A_13_) );
  ADDFX2 U89 ( .A(add_1_root_r119_A_12_), .B(in_17bit_b[6]), .CI(
        add_1_root_r119_carry[12]), .CO(add_1_root_r119_carry[13]), .S(
        add_1_root_r119_SUM_12_) );
  ADDFX2 U90 ( .A(in_17bit_b[7]), .B(in_17bit_b[6]), .CI(
        add_2_root_r119_carry_11_), .CO(add_2_root_r119_carry_12_), .S(
        add_2_root_r119_SUM_11_) );
  ADDFX2 U91 ( .A(in_17bit_b[10]), .B(in_17bit_b[8]), .CI(
        add_2_root_r115_carry_11_), .CO(add_2_root_r115_carry_12_), .S(
        add_2_root_r115_SUM_11_) );
  ADDFX2 U92 ( .A(in_17bit_b[12]), .B(in_17bit_b[8]), .CI(
        add_1_root_r112_carry_12_), .CO(add_1_root_r112_carry_13_), .S(
        add_1_root_r112_SUM_12_) );
  ADDFX2 U93 ( .A(in_17bit_b[9]), .B(in_17bit_b[7]), .CI(
        add_1_root_r115_carry_13_), .CO(add_1_root_r115_carry_14_), .S(
        add_1_root_r115_SUM_13_) );
  ADDFX2 U94 ( .A(in_17bit_b[13]), .B(in_17bit_b[12]), .CI(
        add_3_root_r119_carry_14_), .CO(add_3_root_r119_carry_15_), .S(
        add_1_root_r119_A_14_) );
  ADDFX2 U95 ( .A(add_1_root_r119_A_13_), .B(in_17bit_b[7]), .CI(
        add_1_root_r119_carry[13]), .CO(add_1_root_r119_carry[14]), .S(
        add_1_root_r119_SUM_13_) );
  ADDFX2 U96 ( .A(in_17bit_b[11]), .B(in_17bit_b[9]), .CI(
        add_2_root_r115_carry_12_), .CO(add_2_root_r115_carry_13_), .S(
        add_2_root_r115_SUM_12_) );
  ADDFX2 U97 ( .A(in_17bit_b[13]), .B(in_17bit_b[9]), .CI(
        add_1_root_r112_carry_13_), .CO(add_1_root_r112_carry_14_), .S(
        add_1_root_r112_SUM_13_) );
  ADDFX2 U98 ( .A(in_17bit_b[10]), .B(in_17bit_b[8]), .CI(
        add_1_root_r115_carry_14_), .CO(add_1_root_r115_carry_15_), .S(
        add_1_root_r115_SUM_14_) );
  ADDFX2 U99 ( .A(in_17bit_b[14]), .B(in_17bit_b[13]), .CI(
        add_3_root_r119_carry_15_), .CO(add_3_root_r119_carry_16_), .S(
        add_1_root_r119_A_15_) );
  ADDFX2 U100 ( .A(add_1_root_r119_A_14_), .B(in_17bit_b[8]), .CI(
        add_1_root_r119_carry[14]), .CO(add_1_root_r119_carry[15]), .S(
        add_1_root_r119_SUM_14_) );
  ADDFX2 U101 ( .A(in_17bit_b[3]), .B(in_17bit_b[2]), .CI(
        add_3_root_r119_carry_4_), .CO(add_3_root_r119_carry_5_), .S(
        add_1_root_r119_A_4_) );
  ADDFX2 U102 ( .A(in_17bit_b[2]), .B(in_17bit_b[1]), .CI(
        add_3_root_r119_carry_3_), .CO(add_3_root_r119_carry_4_), .S(
        add_1_root_r119_A_3_) );
  ADDFX2 U103 ( .A(in_17bit_b[9]), .B(in_17bit_b[8]), .CI(
        add_2_root_r119_carry_13_), .CO(add_2_root_r119_carry_14_), .S(
        add_2_root_r119_SUM_13_) );
  ADDFX2 U104 ( .A(in_17bit_b[12]), .B(in_17bit_b[10]), .CI(
        add_2_root_r115_carry_13_), .CO(add_2_root_r115_carry_14_), .S(
        add_2_root_r115_SUM_13_) );
  ADDFX2 U105 ( .A(in_17bit_b[14]), .B(in_17bit_b[10]), .CI(
        add_1_root_r112_carry_14_), .CO(add_1_root_r112_carry_15_), .S(
        add_1_root_r112_SUM_14_) );
  ADDFX2 U106 ( .A(in_17bit_b[11]), .B(in_17bit_b[9]), .CI(
        add_1_root_r115_carry_15_), .CO(add_1_root_r115_carry_16_), .S(
        add_1_root_r115_SUM_15_) );
  ADDFX2 U107 ( .A(add_1_root_r119_A_15_), .B(in_17bit_b[9]), .CI(
        add_1_root_r119_carry[15]), .CO(add_1_root_r119_carry[16]), .S(
        add_1_root_r119_SUM_15_) );
  ADDFX2 U108 ( .A(in_17bit_b[10]), .B(in_17bit_b[9]), .CI(
        add_2_root_r119_carry_14_), .CO(add_2_root_r119_carry_15_), .S(
        add_2_root_r119_SUM_14_) );
  ADDFX2 U109 ( .A(in_17bit_b[13]), .B(in_17bit_b[11]), .CI(
        add_2_root_r115_carry_14_), .CO(add_2_root_r115_carry_15_), .S(
        add_2_root_r115_SUM_14_) );
  ADDFX2 U110 ( .A(in_17bit_b[15]), .B(in_17bit_b[11]), .CI(
        add_1_root_r112_carry_15_), .CO(add_1_root_r112_carry_16_), .S(
        add_1_root_r112_SUM_15_) );
  ADDFX2 U111 ( .A(in_17bit_b[12]), .B(in_17bit_b[10]), .CI(
        add_1_root_r115_carry_16_), .CO(add_1_root_r115_carry_17_), .S(
        add_1_root_r115_SUM_16_) );
  ADDFX2 U112 ( .A(add_1_root_r119_A_16_), .B(in_17bit_b[10]), .CI(
        add_1_root_r119_carry[16]), .CO(add_1_root_r119_carry[17]), .S(
        add_1_root_r119_SUM_16_) );
  ADDFX2 U113 ( .A(in_17bit_b[11]), .B(in_17bit_b[10]), .CI(
        add_2_root_r119_carry_15_), .CO(add_2_root_r119_carry_16_), .S(
        add_2_root_r119_SUM_15_) );
  ADDFX2 U114 ( .A(in_17bit_b[14]), .B(in_17bit_b[12]), .CI(
        add_2_root_r115_carry_15_), .CO(add_2_root_r115_carry_16_), .S(
        add_2_root_r115_SUM_15_) );
  ADDFX2 U115 ( .A(in_17bit_b[13]), .B(in_17bit_b[11]), .CI(
        add_1_root_r115_carry_17_), .CO(add_1_root_r115_carry_18_), .S(
        add_1_root_r115_SUM_17_) );
  ADDFX2 U116 ( .A(add_1_root_r119_A_17_), .B(in_17bit_b[11]), .CI(
        add_1_root_r119_carry[17]), .CO(add_1_root_r119_carry[18]), .S(
        add_1_root_r119_SUM_17_) );
  ADDFX2 U117 ( .A(in_17bit_b[12]), .B(in_17bit_b[11]), .CI(
        add_2_root_r119_carry_16_), .CO(add_2_root_r119_carry_17_), .S(
        add_2_root_r119_SUM_16_) );
  ADDFX2 U118 ( .A(in_17bit_b[14]), .B(in_17bit_b[12]), .CI(
        add_1_root_r115_carry_18_), .CO(add_1_root_r115_carry_19_), .S(
        add_1_root_r115_SUM_18_) );
  ADDFX2 U119 ( .A(add_1_root_r119_A_18_), .B(in_17bit_b[12]), .CI(
        add_1_root_r119_carry[18]), .CO(add_1_root_r119_carry[19]), .S(
        add_1_root_r119_SUM_18_) );
  ADDFX2 U120 ( .A(in_17bit_b[13]), .B(in_17bit_b[12]), .CI(
        add_2_root_r119_carry_17_), .CO(add_2_root_r119_carry_18_), .S(
        add_2_root_r119_SUM_17_) );
  ADDFX2 U121 ( .A(in_17bit_b[5]), .B(in_17bit_b[3]), .CI(
        add_2_root_r115_carry_6_), .CO(add_2_root_r115_carry_7_), .S(
        add_2_root_r115_SUM_6_) );
  ADDFX2 U122 ( .A(in_17bit_b[7]), .B(in_17bit_b[3]), .CI(
        add_1_root_r112_carry_7_), .CO(add_1_root_r112_carry_8_), .S(
        add_1_root_r112_SUM_7_) );
  ADDFX2 U123 ( .A(add_1_root_r119_A_11_), .B(in_17bit_b[5]), .CI(
        add_1_root_r119_carry[11]), .CO(add_1_root_r119_carry[12]), .S(
        add_1_root_r119_SUM_11_) );
  ADDFX2 U124 ( .A(in_17bit_b[5]), .B(in_17bit_b[3]), .CI(
        add_1_root_r115_carry_9_), .CO(add_1_root_r115_carry_10_), .S(
        add_1_root_r115_SUM_9_) );
  ADDFX2 U125 ( .A(add_1_root_r119_A_9_), .B(in_17bit_b[3]), .CI(
        add_1_root_r119_carry[9]), .CO(add_1_root_r119_carry[10]), .S(
        add_1_root_r119_SUM_9_) );
  ADDFX2 U126 ( .A(in_17bit_b[4]), .B(in_17bit_b[3]), .CI(
        add_3_root_r119_carry_5_), .CO(add_3_root_r119_carry_6_), .S(
        add_1_root_r119_A_5_) );
  ADDFX2 U127 ( .A(in_17bit_b[15]), .B(in_17bit_b[13]), .CI(
        add_1_root_r115_carry_19_), .CO(add_1_root_r115_carry_20_), .S(
        add_1_root_r115_SUM_19_) );
  ADDFX2 U128 ( .A(in_17bit_b[4]), .B(in_17bit_b[3]), .CI(
        add_2_root_r119_carry_8_), .CO(add_2_root_r119_carry_9_), .S(
        add_2_root_r119_SUM_8_) );
  ADDFX2 U129 ( .A(add_1_root_r119_A_10_), .B(in_17bit_b[4]), .CI(
        add_1_root_r119_carry[10]), .CO(add_1_root_r119_carry[11]), .S(
        add_1_root_r119_SUM_10_) );
  ADDFX2 U130 ( .A(in_17bit_b[8]), .B(in_17bit_b[7]), .CI(
        add_2_root_r119_carry_12_), .CO(add_2_root_r119_carry_13_), .S(
        add_2_root_r119_SUM_12_) );
  ADDFX2 U131 ( .A(in_17bit_b[15]), .B(in_17bit_b[14]), .CI(
        add_3_root_r119_carry_16_), .CO(add_3_root_r119_carry_17_), .S(
        add_1_root_r119_A_16_) );
  ADDFX2 U132 ( .A(in_17bit_b[15]), .B(in_17bit_b[13]), .CI(
        add_2_root_r115_carry_16_), .CO(add_2_root_r115_carry_17_), .S(
        add_2_root_r115_SUM_16_) );
  ADDFX2 U133 ( .A(in_17bit_b[5]), .B(in_17bit_b[4]), .CI(
        add_3_root_r119_carry_6_), .CO(add_3_root_r119_carry_7_), .S(
        add_1_root_r119_A_6_) );
  ADDFX2 U134 ( .A(in_17bit_b[14]), .B(in_17bit_b[13]), .CI(
        add_2_root_r119_carry_18_), .CO(add_2_root_r119_carry_19_), .S(
        add_2_root_r119_SUM_18_) );
  ADDFX2 U135 ( .A(in_17bit_b[15]), .B(in_17bit_b[14]), .CI(
        add_2_root_r119_carry_19_), .CO(add_2_root_r119_carry_20_), .S(
        add_2_root_r119_SUM_19_) );
  INVX1 U136 ( .A(n190), .Y(n67) );
  BUFX3 U137 ( .A(in_17bit_b[16]), .Y(n37) );
  INVX1 U138 ( .A(n245), .Y(in_17bit_b[16]) );
  INVX1 U139 ( .A(in_8bit[2]), .Y(n43) );
  INVX1 U140 ( .A(in_8bit[3]), .Y(n41) );
  INVX1 U141 ( .A(in_8bit[6]), .Y(n39) );
  INVX1 U142 ( .A(in_8bit[5]), .Y(n44) );
  INVX1 U143 ( .A(in_8bit[4]), .Y(n40) );
  CLKINVX3 U144 ( .A(n192), .Y(in_17bit_b[0]) );
  NOR3X1 U145 ( .A(n43), .B(n41), .C(n98), .Y(n190) );
  NAND2X1 U146 ( .A(N29), .B(n48), .Y(n245) );
  NAND4BXL U147 ( .AN(in_8bit[7]), .B(in_8bit[4]), .C(in_8bit[5]), .D(n189), 
        .Y(n68) );
  CLKINVX3 U148 ( .A(n237), .Y(in_17bit_b[15]) );
  OR2X2 U149 ( .A(n72), .B(n71), .Y(n241) );
  NOR2X1 U150 ( .A(n73), .B(n184), .Y(n71) );
  NOR2X1 U151 ( .A(n185), .B(n183), .Y(n72) );
  OR2X2 U152 ( .A(n75), .B(n74), .Y(n242) );
  NOR2X1 U153 ( .A(n73), .B(n185), .Y(n74) );
  NOR2X1 U154 ( .A(n184), .B(n183), .Y(n75) );
  OAI2BB1X1 U155 ( .A0N(n189), .A1N(n79), .B0(n78), .Y(n97) );
  INVX1 U156 ( .A(n76), .Y(n79) );
  NAND3BX1 U157 ( .AN(n77), .B(n190), .C(in_8bit[5]), .Y(n78) );
  NAND2X1 U158 ( .A(n194), .B(n193), .Y(N447) );
  AOI22X1 U159 ( .A0(N108), .A1(n238), .B0(N205), .B1(n242), .Y(n193) );
  AOI22X1 U160 ( .A0(N347), .A1(n241), .B0(n97), .B1(in_17bit_b[0]), .Y(n194)
         );
  NAND2X1 U161 ( .A(n197), .B(n196), .Y(N448) );
  AOI22X1 U162 ( .A0(N109), .A1(n238), .B0(N206), .B1(n242), .Y(n196) );
  AOI22X1 U163 ( .A0(N348), .A1(n241), .B0(n97), .B1(n96), .Y(n197) );
  INVX1 U164 ( .A(n195), .Y(n96) );
  NAND2X1 U165 ( .A(n200), .B(n199), .Y(N449) );
  AOI22X1 U166 ( .A0(N110), .A1(n238), .B0(N207), .B1(n242), .Y(n199) );
  AOI22X1 U167 ( .A0(N349), .A1(n241), .B0(n97), .B1(in_17bit_b[2]), .Y(n200)
         );
  NAND2X1 U168 ( .A(n203), .B(n202), .Y(N450) );
  AOI22X1 U169 ( .A0(N111), .A1(n238), .B0(N208), .B1(n242), .Y(n202) );
  AOI22X1 U170 ( .A0(N350), .A1(n241), .B0(n97), .B1(in_17bit_b[3]), .Y(n203)
         );
  NAND2X1 U171 ( .A(n206), .B(n205), .Y(N451) );
  AOI22X1 U172 ( .A0(N112), .A1(n238), .B0(N209), .B1(n242), .Y(n205) );
  AOI22X1 U173 ( .A0(N351), .A1(n241), .B0(n97), .B1(in_17bit_b[4]), .Y(n206)
         );
  NAND2X1 U174 ( .A(n209), .B(n208), .Y(N452) );
  AOI22X1 U175 ( .A0(N113), .A1(n238), .B0(N210), .B1(n242), .Y(n208) );
  AOI22X1 U176 ( .A0(N352), .A1(n241), .B0(n97), .B1(in_17bit_b[5]), .Y(n209)
         );
  NAND2X1 U177 ( .A(n212), .B(n211), .Y(N453) );
  AOI22X1 U178 ( .A0(N114), .A1(n238), .B0(N211), .B1(n242), .Y(n211) );
  AOI22X1 U179 ( .A0(N353), .A1(n241), .B0(n97), .B1(in_17bit_b[6]), .Y(n212)
         );
  NAND2X1 U180 ( .A(n215), .B(n214), .Y(N454) );
  AOI22X1 U181 ( .A0(N115), .A1(n238), .B0(N212), .B1(n242), .Y(n214) );
  AOI22X1 U182 ( .A0(N354), .A1(n241), .B0(n97), .B1(in_17bit_b[7]), .Y(n215)
         );
  NAND2X1 U183 ( .A(n218), .B(n217), .Y(N455) );
  AOI22X1 U184 ( .A0(N116), .A1(n238), .B0(N213), .B1(n242), .Y(n217) );
  AOI22X1 U185 ( .A0(N355), .A1(n241), .B0(n97), .B1(in_17bit_b[8]), .Y(n218)
         );
  NAND2X1 U186 ( .A(n221), .B(n220), .Y(N456) );
  AOI22X1 U187 ( .A0(N117), .A1(n238), .B0(N214), .B1(n242), .Y(n220) );
  AOI22X1 U188 ( .A0(N356), .A1(n241), .B0(n97), .B1(in_17bit_b[9]), .Y(n221)
         );
  NAND2X1 U189 ( .A(n224), .B(n223), .Y(N457) );
  AOI22X1 U190 ( .A0(N118), .A1(n238), .B0(N215), .B1(n242), .Y(n223) );
  AOI22X1 U191 ( .A0(N357), .A1(n241), .B0(n97), .B1(in_17bit_b[10]), .Y(n224)
         );
  NAND2X1 U192 ( .A(n227), .B(n226), .Y(N458) );
  AOI22X1 U193 ( .A0(N119), .A1(n238), .B0(N216), .B1(n242), .Y(n226) );
  AOI22X1 U194 ( .A0(N358), .A1(n241), .B0(n97), .B1(in_17bit_b[11]), .Y(n227)
         );
  NAND2X1 U195 ( .A(n230), .B(n229), .Y(N459) );
  AOI22X1 U196 ( .A0(N120), .A1(n238), .B0(N217), .B1(n242), .Y(n229) );
  AOI22X1 U197 ( .A0(N359), .A1(n241), .B0(n97), .B1(in_17bit_b[12]), .Y(n230)
         );
  NAND2X1 U198 ( .A(n233), .B(n232), .Y(N460) );
  AOI22X1 U199 ( .A0(N121), .A1(n238), .B0(N218), .B1(n242), .Y(n232) );
  AOI22X1 U200 ( .A0(N360), .A1(n241), .B0(n97), .B1(in_17bit_b[13]), .Y(n233)
         );
  NAND2X1 U201 ( .A(n236), .B(n235), .Y(N461) );
  AOI22X1 U202 ( .A0(N122), .A1(n238), .B0(N219), .B1(n242), .Y(n235) );
  AOI22X1 U203 ( .A0(N361), .A1(n241), .B0(n97), .B1(in_17bit_b[14]), .Y(n236)
         );
  NAND2X1 U204 ( .A(n240), .B(n239), .Y(N462) );
  AOI22X1 U205 ( .A0(N123), .A1(n238), .B0(N220), .B1(n242), .Y(n239) );
  AOI22X1 U206 ( .A0(N362), .A1(n241), .B0(n97), .B1(in_17bit_b[15]), .Y(n240)
         );
  INVX1 U207 ( .A(n56), .Y(n58) );
  MXI2XL U208 ( .A(n1), .B(n17), .S0(n66), .Y(out[16]) );
  NAND4BBX1 U209 ( .AN(n241), .BN(n242), .C(n191), .D(n244), .Y(N446) );
  AOI2BB1X1 U210 ( .A0N(n188), .A1N(n187), .B0(n238), .Y(n191) );
  OR4XL U211 ( .A(in_8bit[4]), .B(in_8bit[5]), .C(n38), .D(in_8bit[7]), .Y(
        n188) );
  NOR2X1 U212 ( .A(n38), .B(in_8bit[4]), .Y(n182) );
  NOR4BX1 U213 ( .AN(n186), .B(n98), .C(in_8bit[1]), .D(in_8bit[2]), .Y(n189)
         );
  NOR2X1 U214 ( .A(n38), .B(in_8bit[3]), .Y(n186) );
  INVXL U215 ( .A(in_8bit[0]), .Y(n98) );
  NAND4BXL U216 ( .AN(in_8bit[7]), .B(n38), .C(in_8bit[1]), .D(in_8bit[4]), 
        .Y(n77) );
  AOI22X1 U217 ( .A0(N22), .A1(n48), .B0(in_17bit[9]), .B1(n36), .Y(n219) );
  AOI22X1 U218 ( .A0(N23), .A1(n48), .B0(in_17bit[10]), .B1(n36), .Y(n222) );
  AOI22X1 U219 ( .A0(N27), .A1(n48), .B0(in_17bit[14]), .B1(n49), .Y(n234) );
  AOI22X1 U220 ( .A0(N28), .A1(n48), .B0(in_17bit[15]), .B1(n36), .Y(n237) );
  AOI22X1 U221 ( .A0(N24), .A1(n48), .B0(in_17bit[11]), .B1(n49), .Y(n225) );
  AOI22X1 U222 ( .A0(N25), .A1(n48), .B0(in_17bit[12]), .B1(n36), .Y(n228) );
  AOI22X1 U223 ( .A0(N26), .A1(n48), .B0(in_17bit[13]), .B1(n50), .Y(n231) );
  AOI22X1 U224 ( .A0(N21), .A1(n48), .B0(in_17bit[8]), .B1(n49), .Y(n216) );
  INVX1 U225 ( .A(n51), .Y(n60) );
  NAND2BX1 U226 ( .AN(n56), .B(n2), .Y(n51) );
  AND2X2 U227 ( .A(n60), .B(n4), .Y(n26) );
  AND2X2 U228 ( .A(n26), .B(n5), .Y(n27) );
  AND2X2 U229 ( .A(n27), .B(n6), .Y(n28) );
  OR2XL U230 ( .A(n77), .B(in_8bit[0]), .Y(n73) );
  AND2X2 U231 ( .A(n28), .B(n7), .Y(n29) );
  OAI2BB1X1 U232 ( .A0N(n70), .A1N(n69), .B0(n68), .Y(n238) );
  NOR2X1 U233 ( .A(n39), .B(n67), .Y(n70) );
  NOR2BX1 U234 ( .AN(in_8bit[1]), .B(n76), .Y(n69) );
  AND2X2 U235 ( .A(n29), .B(n3), .Y(n30) );
  NAND2X1 U236 ( .A(n33), .B(n15), .Y(n56) );
  INVX1 U237 ( .A(in_17bit[8]), .Y(n88) );
  INVX1 U238 ( .A(in_17bit[9]), .Y(n89) );
  INVX1 U239 ( .A(in_17bit[10]), .Y(n90) );
  INVX1 U240 ( .A(in_17bit[11]), .Y(n91) );
  INVX1 U241 ( .A(in_17bit[12]), .Y(n92) );
  INVX1 U242 ( .A(in_17bit[13]), .Y(n93) );
  INVX1 U243 ( .A(in_17bit[14]), .Y(n94) );
  INVX1 U244 ( .A(in_17bit[15]), .Y(n95) );
  INVX1 U245 ( .A(in_17bit[1]), .Y(n81) );
  INVX1 U246 ( .A(in_17bit[2]), .Y(n82) );
  INVX1 U247 ( .A(in_17bit[3]), .Y(n83) );
  INVX1 U248 ( .A(in_17bit[4]), .Y(n84) );
  INVX1 U249 ( .A(in_17bit[5]), .Y(n85) );
  INVX1 U250 ( .A(in_17bit[6]), .Y(n86) );
  INVX1 U251 ( .A(in_17bit[7]), .Y(n87) );
  INVX1 U252 ( .A(in_17bit[0]), .Y(n80) );
  XNOR2X1 U253 ( .A(n13), .B(sub_add_75_b0_carry[11]), .Y(n31) );
  XNOR2X1 U254 ( .A(n16), .B(sub_add_75_b0_carry[10]), .Y(n32) );
  MX2X1 U255 ( .A(neg_mul[21]), .B(N479), .S0(n66), .Y(out[14]) );
  MX2X1 U256 ( .A(neg_mul[22]), .B(N480), .S0(n66), .Y(out[15]) );
  NOR2X1 U257 ( .A(out[0]), .B(neg_mul[8]), .Y(n33) );
  NAND2X1 U258 ( .A(sub_add_75_b0_carry[15]), .B(n9), .Y(n34) );
  XNOR2X4 U259 ( .A(n19), .B(n42), .Y(n54) );
  INVX1 U260 ( .A(n36), .Y(n46) );
  AOI22XL U261 ( .A0(in_17bit[0]), .A1(n46), .B0(in_17bit[0]), .B1(n50), .Y(
        n192) );
  AOI22XL U262 ( .A0(N14), .A1(n46), .B0(in_17bit[1]), .B1(n50), .Y(n195) );
  AOI22XL U263 ( .A0(N15), .A1(n46), .B0(in_17bit[2]), .B1(n49), .Y(n198) );
  AOI22XL U264 ( .A0(N16), .A1(n46), .B0(in_17bit[3]), .B1(n49), .Y(n201) );
  AOI22XL U265 ( .A0(N17), .A1(n46), .B0(in_17bit[4]), .B1(n50), .Y(n204) );
  AOI22XL U266 ( .A0(N18), .A1(n46), .B0(in_17bit[5]), .B1(n36), .Y(n207) );
  AOI22XL U267 ( .A0(N19), .A1(n46), .B0(in_17bit[6]), .B1(n36), .Y(n210) );
  AOI22XL U268 ( .A0(N20), .A1(n46), .B0(in_17bit[7]), .B1(n36), .Y(n213) );
  OR4X1 U269 ( .A(in_8bit[1]), .B(in_8bit[0]), .C(in_8bit[2]), .D(in_8bit[3]), 
        .Y(n187) );
  XOR2X4 U270 ( .A(n53), .B(neg_mul[8]), .Y(out[1]) );
  NOR2X4 U271 ( .A(n54), .B(n33), .Y(n55) );
  XOR2X4 U272 ( .A(in_17bit[16]), .B(n42), .Y(n57) );
  NOR2X4 U273 ( .A(n58), .B(n57), .Y(n59) );
  XNOR2X4 U274 ( .A(n59), .B(n2), .Y(out[3]) );
  XNOR2X4 U275 ( .A(n61), .B(n4), .Y(out[4]) );
  XNOR2X4 U276 ( .A(n62), .B(n5), .Y(out[5]) );
  NOR2X4 U277 ( .A(n27), .B(n21), .Y(n63) );
  XNOR2X4 U278 ( .A(n63), .B(n6), .Y(out[6]) );
  XNOR2X4 U279 ( .A(n64), .B(n7), .Y(out[7]) );
  MXI2X4 U280 ( .A(n13), .B(n31), .S0(n66), .Y(out[11]) );
  AND2X1 U281 ( .A(add_1_root_r112_carry_20_), .B(n37), .Y(
        add_1_root_r112_SUM_21_) );
  XOR2X1 U282 ( .A(n37), .B(add_1_root_r112_carry_20_), .Y(
        add_1_root_r112_SUM_20_) );
  AND2X1 U283 ( .A(add_1_root_r112_carry_19_), .B(in_17bit_b[15]), .Y(
        add_1_root_r112_carry_20_) );
  XOR2X1 U284 ( .A(in_17bit_b[15]), .B(add_1_root_r112_carry_19_), .Y(
        add_1_root_r112_SUM_19_) );
  AND2X1 U285 ( .A(add_1_root_r112_carry_18_), .B(in_17bit_b[14]), .Y(
        add_1_root_r112_carry_19_) );
  XOR2X1 U286 ( .A(in_17bit_b[14]), .B(add_1_root_r112_carry_18_), .Y(
        add_1_root_r112_SUM_18_) );
  AND2X1 U287 ( .A(add_1_root_r112_carry_17_), .B(in_17bit_b[13]), .Y(
        add_1_root_r112_carry_18_) );
  XOR2X1 U288 ( .A(in_17bit_b[13]), .B(add_1_root_r112_carry_17_), .Y(
        add_1_root_r112_SUM_17_) );
  AND2X1 U289 ( .A(add_2_root_r119_carry_21_), .B(n37), .Y(
        add_2_root_r119_SUM_22_) );
  XOR2X1 U290 ( .A(n37), .B(add_2_root_r119_carry_21_), .Y(
        add_2_root_r119_SUM_21_) );
  AND2X1 U291 ( .A(in_17bit_b[1]), .B(in_17bit_b[0]), .Y(
        add_2_root_r119_carry_6_) );
  XOR2X1 U292 ( .A(in_17bit_b[0]), .B(in_17bit_b[1]), .Y(
        add_2_root_r119_SUM_5_) );
  AND2X1 U293 ( .A(add_1_root_r119_carry[22]), .B(n37), .Y(
        add_1_root_r119_SUM_23_) );
  XOR2X1 U294 ( .A(n37), .B(add_1_root_r119_carry[22]), .Y(
        add_1_root_r119_SUM_22_) );
  AND2X1 U295 ( .A(add_1_root_r119_carry[21]), .B(in_17bit_b[15]), .Y(
        add_1_root_r119_carry[22]) );
  XOR2X1 U296 ( .A(in_17bit_b[15]), .B(add_1_root_r119_carry[21]), .Y(
        add_1_root_r119_SUM_21_) );
  AND2X1 U297 ( .A(add_1_root_r119_carry[20]), .B(in_17bit_b[14]), .Y(
        add_1_root_r119_carry[21]) );
  XOR2X1 U298 ( .A(in_17bit_b[14]), .B(add_1_root_r119_carry[20]), .Y(
        add_1_root_r119_SUM_20_) );
  AND2X1 U299 ( .A(add_1_root_r119_A_6_), .B(in_17bit_b[0]), .Y(
        add_1_root_r119_carry[7]) );
  XOR2X1 U300 ( .A(in_17bit_b[0]), .B(add_1_root_r119_A_6_), .Y(
        add_1_root_r119_SUM_6_) );
  AND2X1 U301 ( .A(add_3_root_r119_carry_18_), .B(n37), .Y(
        add_1_root_r119_A_19_) );
  XOR2X1 U302 ( .A(n37), .B(add_3_root_r119_carry_18_), .Y(
        add_1_root_r119_A_18_) );
  AND2X1 U303 ( .A(in_17bit_b[1]), .B(in_17bit_b[0]), .Y(
        add_3_root_r119_carry_3_) );
  XOR2X1 U304 ( .A(in_17bit_b[0]), .B(in_17bit_b[1]), .Y(add_1_root_r119_A_2_)
         );
  AND2X1 U305 ( .A(add_2_root_r115_carry_19_), .B(n37), .Y(
        add_2_root_r115_SUM_20_) );
  XOR2X1 U306 ( .A(n37), .B(add_2_root_r115_carry_19_), .Y(
        add_2_root_r115_SUM_19_) );
  AND2X1 U307 ( .A(add_2_root_r115_carry_18_), .B(in_17bit_b[15]), .Y(
        add_2_root_r115_carry_19_) );
  XOR2X1 U308 ( .A(in_17bit_b[15]), .B(add_2_root_r115_carry_18_), .Y(
        add_2_root_r115_SUM_18_) );
  AND2X1 U309 ( .A(in_17bit_b[2]), .B(in_17bit_b[0]), .Y(
        add_2_root_r115_carry_4_) );
  XOR2X1 U310 ( .A(in_17bit_b[0]), .B(in_17bit_b[2]), .Y(
        add_2_root_r115_SUM_3_) );
  AND2X1 U311 ( .A(add_1_root_r115_carry_22_), .B(n37), .Y(
        add_1_root_r115_SUM_23_) );
  XOR2X1 U312 ( .A(n37), .B(add_1_root_r115_carry_22_), .Y(
        add_1_root_r115_SUM_22_) );
  AND2X1 U313 ( .A(add_1_root_r115_carry_21_), .B(in_17bit_b[15]), .Y(
        add_1_root_r115_carry_22_) );
  XOR2X1 U314 ( .A(in_17bit_b[15]), .B(add_1_root_r115_carry_21_), .Y(
        add_1_root_r115_SUM_21_) );
  AND2X1 U315 ( .A(in_17bit_b[2]), .B(in_17bit_b[0]), .Y(
        add_1_root_r115_carry_7_) );
  XOR2X1 U316 ( .A(in_17bit_b[0]), .B(in_17bit_b[2]), .Y(
        add_1_root_r115_SUM_6_) );
  XOR2X1 U317 ( .A(n50), .B(sub_add_54_b0_carry[16]), .Y(N29) );
  AND2X1 U318 ( .A(sub_add_54_b0_carry[15]), .B(n95), .Y(
        sub_add_54_b0_carry[16]) );
  XOR2X1 U319 ( .A(n95), .B(sub_add_54_b0_carry[15]), .Y(N28) );
  AND2X1 U320 ( .A(sub_add_54_b0_carry[14]), .B(n94), .Y(
        sub_add_54_b0_carry[15]) );
  XOR2X1 U321 ( .A(n94), .B(sub_add_54_b0_carry[14]), .Y(N27) );
  AND2X1 U322 ( .A(sub_add_54_b0_carry[13]), .B(n93), .Y(
        sub_add_54_b0_carry[14]) );
  XOR2X1 U323 ( .A(n93), .B(sub_add_54_b0_carry[13]), .Y(N26) );
  AND2X1 U324 ( .A(sub_add_54_b0_carry[12]), .B(n92), .Y(
        sub_add_54_b0_carry[13]) );
  XOR2X1 U325 ( .A(n92), .B(sub_add_54_b0_carry[12]), .Y(N25) );
  AND2X1 U326 ( .A(sub_add_54_b0_carry[11]), .B(n91), .Y(
        sub_add_54_b0_carry[12]) );
  XOR2X1 U327 ( .A(n91), .B(sub_add_54_b0_carry[11]), .Y(N24) );
  AND2X1 U328 ( .A(sub_add_54_b0_carry[10]), .B(n90), .Y(
        sub_add_54_b0_carry[11]) );
  XOR2X1 U329 ( .A(n90), .B(sub_add_54_b0_carry[10]), .Y(N23) );
  AND2X1 U330 ( .A(sub_add_54_b0_carry[9]), .B(n89), .Y(
        sub_add_54_b0_carry[10]) );
  XOR2X1 U331 ( .A(n89), .B(sub_add_54_b0_carry[9]), .Y(N22) );
  AND2X1 U332 ( .A(sub_add_54_b0_carry[8]), .B(n88), .Y(sub_add_54_b0_carry[9]) );
  XOR2X1 U333 ( .A(n88), .B(sub_add_54_b0_carry[8]), .Y(N21) );
  AND2X1 U334 ( .A(sub_add_54_b0_carry[7]), .B(n87), .Y(sub_add_54_b0_carry[8]) );
  XOR2X1 U335 ( .A(n87), .B(sub_add_54_b0_carry[7]), .Y(N20) );
  AND2X1 U336 ( .A(sub_add_54_b0_carry[6]), .B(n86), .Y(sub_add_54_b0_carry[7]) );
  XOR2X1 U337 ( .A(n86), .B(sub_add_54_b0_carry[6]), .Y(N19) );
  AND2X1 U338 ( .A(sub_add_54_b0_carry[5]), .B(n85), .Y(sub_add_54_b0_carry[6]) );
  XOR2X1 U339 ( .A(n85), .B(sub_add_54_b0_carry[5]), .Y(N18) );
  AND2X1 U340 ( .A(sub_add_54_b0_carry[4]), .B(n84), .Y(sub_add_54_b0_carry[5]) );
  XOR2X1 U341 ( .A(n84), .B(sub_add_54_b0_carry[4]), .Y(N17) );
  AND2X1 U342 ( .A(sub_add_54_b0_carry[3]), .B(n83), .Y(sub_add_54_b0_carry[4]) );
  XOR2X1 U343 ( .A(n83), .B(sub_add_54_b0_carry[3]), .Y(N16) );
  AND2X1 U344 ( .A(sub_add_54_b0_carry[2]), .B(n82), .Y(sub_add_54_b0_carry[3]) );
  XOR2X1 U345 ( .A(n82), .B(sub_add_54_b0_carry[2]), .Y(N15) );
  AND2X1 U346 ( .A(n80), .B(n81), .Y(sub_add_54_b0_carry[2]) );
  XOR2X1 U347 ( .A(n81), .B(n80), .Y(N14) );
  XOR2X1 U348 ( .A(n9), .B(sub_add_75_b0_carry[15]), .Y(N480) );
  AND2X1 U349 ( .A(sub_add_75_b0_carry[14]), .B(n11), .Y(
        sub_add_75_b0_carry[15]) );
  XOR2X1 U350 ( .A(n11), .B(sub_add_75_b0_carry[14]), .Y(N479) );
  AND2X1 U351 ( .A(sub_add_75_b0_carry[13]), .B(n12), .Y(
        sub_add_75_b0_carry[14]) );
  XOR2X1 U352 ( .A(n12), .B(sub_add_75_b0_carry[13]), .Y(N478) );
  AND2X1 U353 ( .A(sub_add_75_b0_carry[12]), .B(n10), .Y(
        sub_add_75_b0_carry[13]) );
  XOR2X1 U354 ( .A(n10), .B(sub_add_75_b0_carry[12]), .Y(N477) );
  AND2X1 U355 ( .A(sub_add_75_b0_carry[11]), .B(n13), .Y(
        sub_add_75_b0_carry[12]) );
  AND2X1 U356 ( .A(sub_add_75_b0_carry[10]), .B(n16), .Y(
        sub_add_75_b0_carry[11]) );
  AND2X1 U357 ( .A(n30), .B(n8), .Y(sub_add_75_b0_carry[10]) );
  AND2X1 U358 ( .A(in_17bit_b[0]), .B(in_17bit_b[4]), .Y(
        add_1_root_r112_carry_5_) );
endmodule


module multi16_7_DW01_add_0 ( A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, 
        A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, 
        A_4_, B_23_, B_22_, B_21_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, 
        B_14_, B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, 
        SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, 
        SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, 
        SUM_7_ );
  input A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_,
         A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, B_23_, B_22_,
         B_21_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_,
         B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_;
  output SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_,
         SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_,
         SUM_8_, SUM_7_;
  wire   n1, n2, n3, n4;
  wire   [23:7] carry;

  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry[7]), .CO(carry[8]), .S(SUM_7_)
         );
  ADDFX2 U1_21 ( .A(A_21_), .B(B_21_), .CI(carry[21]), .CO(carry[22]), .S(
        SUM_21_) );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry[20]), .CO(carry[21]), .S(
        SUM_20_) );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry[19]), .CO(carry[20]), .S(
        SUM_19_) );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry[18]), .CO(carry[19]), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry[17]), .CO(carry[18]), .S(
        SUM_17_) );
  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry[16]), .CO(carry[17]), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry[15]), .CO(carry[16]), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry[14]), .CO(carry[15]), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry[13]), .CO(carry[14]), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry[12]), .CO(carry[13]), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry[11]), .CO(carry[12]), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry[10]), .CO(carry[11]), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry[9]), .CO(carry[10]), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry[8]), .CO(carry[9]), .S(SUM_8_)
         );
  ADDFX2 U1_22 ( .A(A_22_), .B(B_22_), .CI(carry[22]), .CO(carry[23]), .S(
        SUM_22_) );
  AND2X2 U1 ( .A(A_4_), .B(B_4_), .Y(n1) );
  XOR2X1 U2 ( .A(B_23_), .B(carry[23]), .Y(SUM_23_) );
  OAI2BB1X1 U3 ( .A0N(n2), .A1N(A_6_), .B0(n3), .Y(carry[7]) );
  OAI21XL U4 ( .A0(A_6_), .A1(n2), .B0(B_6_), .Y(n3) );
  OAI2BB1X1 U5 ( .A0N(n1), .A1N(A_5_), .B0(n4), .Y(n2) );
  OAI21XL U6 ( .A0(A_5_), .A1(n1), .B0(B_5_), .Y(n4) );
endmodule


module multi16_7_DW01_add_4 ( A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, 
        A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, 
        B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, 
        B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, SUM_22_, SUM_21_, SUM_20_, 
        SUM_19_, SUM_18_, SUM_17_, SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, 
        SUM_11_, SUM_10_, SUM_9_, SUM_8_, SUM_7_ );
  input A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_,
         A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, B_20_, B_19_,
         B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, B_10_, B_9_,
         B_8_, B_7_, B_6_, B_5_;
  output SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_,
         SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_,
         SUM_7_;
  wire   carry_21_, carry_20_, carry_19_, carry_18_, carry_17_, carry_16_,
         carry_15_, carry_14_, carry_13_, carry_12_, carry_11_, carry_10_,
         carry_9_, carry_8_, carry_7_, n1;

  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry_16_), .CO(carry_17_), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry_15_), .CO(carry_16_), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry_14_), .CO(carry_15_), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry_13_), .CO(carry_14_), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry_12_), .CO(carry_13_), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry_11_), .CO(carry_12_), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry_10_), .CO(carry_11_), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry_9_), .CO(carry_10_), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry_8_), .CO(carry_9_), .S(SUM_8_)
         );
  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry_7_), .CO(carry_8_), .S(SUM_7_)
         );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry_20_), .CO(carry_21_), .S(
        SUM_20_) );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry_19_), .CO(carry_20_), .S(
        SUM_19_) );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry_18_), .CO(carry_19_), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry_17_), .CO(carry_18_), .S(
        SUM_17_) );
  ADDFX2 U1_21 ( .A(A_21_), .B(B_21_), .CI(carry_21_), .CO(SUM_22_), .S(
        SUM_21_) );
  OAI2BB1X1 U1 ( .A0N(A_6_), .A1N(B_6_), .B0(n1), .Y(carry_7_) );
  OAI211X1 U2 ( .A0(B_6_), .A1(A_6_), .B0(A_5_), .C0(B_5_), .Y(n1) );
endmodule


module multi16_7_DW01_add_6 ( A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, 
        A_16_, A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, 
        A_6_, A_5_, A_4_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, 
        B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, 
        SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, 
        SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, 
        SUM_7_ );
  input A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_,
         A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, B_20_,
         B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, B_10_,
         B_9_, B_8_, B_7_, B_6_, B_5_, B_4_;
  output SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_,
         SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_,
         SUM_8_, SUM_7_;
  wire   n1, n2, n3, n4, n5, n6;
  wire   [21:7] carry;

  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry[7]), .CO(carry[8]), .S(SUM_7_)
         );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry[18]), .CO(carry[19]), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry[17]), .CO(carry[18]), .S(
        SUM_17_) );
  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry[16]), .CO(carry[17]), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry[15]), .CO(carry[16]), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry[14]), .CO(carry[15]), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry[13]), .CO(carry[14]), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry[12]), .CO(carry[13]), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry[11]), .CO(carry[12]), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry[10]), .CO(carry[11]), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry[9]), .CO(carry[10]), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry[8]), .CO(carry[9]), .S(SUM_8_)
         );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry[19]), .CO(carry[20]), .S(
        SUM_19_) );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry[20]), .CO(carry[21]), .S(
        SUM_20_) );
  AND2X2 U1 ( .A(A_22_), .B(n2), .Y(n1) );
  AND2X2 U2 ( .A(A_21_), .B(carry[21]), .Y(n2) );
  AND2X2 U3 ( .A(A_4_), .B(B_4_), .Y(n3) );
  XOR2X1 U4 ( .A(A_23_), .B(n1), .Y(SUM_23_) );
  XOR2X1 U5 ( .A(A_21_), .B(carry[21]), .Y(SUM_21_) );
  XOR2X1 U6 ( .A(A_22_), .B(n2), .Y(SUM_22_) );
  OAI2BB1X1 U7 ( .A0N(n4), .A1N(A_6_), .B0(n5), .Y(carry[7]) );
  OAI21XL U8 ( .A0(A_6_), .A1(n4), .B0(B_6_), .Y(n5) );
  OAI2BB1X1 U9 ( .A0N(n3), .A1N(A_5_), .B0(n6), .Y(n4) );
  OAI21XL U10 ( .A0(A_5_), .A1(n3), .B0(B_5_), .Y(n6) );
endmodule


module multi16_7 ( in_17bit, in_8bit, out );
  input [16:0] in_17bit;
  input [7:0] in_8bit;
  output [16:0] out;
  wire   N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27,
         N28, N29, N108, N109, N110, N111, N112, N113, N114, N115, N116, N117,
         N118, N119, N120, N121, N122, N123, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220,
         N221, N347, N348, N349, N350, N351, N352, N353, N354, N355, N356,
         N357, N358, N359, N360, N361, N362, N363, N446, N447, N448, N449,
         N450, N451, N452, N453, N454, N455, N456, N457, N458, N459, N460,
         N461, N462, N463, N475, N477, N479, N480, N481,
         add_2_root_r119_carry_10_, add_2_root_r119_carry_11_,
         add_2_root_r119_carry_12_, add_2_root_r119_carry_13_,
         add_2_root_r119_carry_14_, add_2_root_r119_carry_15_,
         add_2_root_r119_carry_16_, add_2_root_r119_carry_17_,
         add_2_root_r119_carry_18_, add_2_root_r119_carry_19_,
         add_2_root_r119_carry_20_, add_2_root_r119_carry_21_,
         add_2_root_r119_carry_6_, add_2_root_r119_carry_7_,
         add_2_root_r119_carry_8_, add_2_root_r119_carry_9_,
         add_2_root_r119_SUM_5_, add_2_root_r119_SUM_6_,
         add_2_root_r119_SUM_7_, add_2_root_r119_SUM_8_,
         add_2_root_r119_SUM_9_, add_2_root_r119_SUM_10_,
         add_2_root_r119_SUM_11_, add_2_root_r119_SUM_12_,
         add_2_root_r119_SUM_13_, add_2_root_r119_SUM_14_,
         add_2_root_r119_SUM_15_, add_2_root_r119_SUM_16_,
         add_2_root_r119_SUM_17_, add_2_root_r119_SUM_18_,
         add_2_root_r119_SUM_19_, add_2_root_r119_SUM_20_,
         add_2_root_r119_SUM_21_, add_2_root_r119_SUM_22_,
         add_1_root_r119_SUM_6_, add_1_root_r119_SUM_7_,
         add_1_root_r119_SUM_8_, add_1_root_r119_SUM_9_,
         add_1_root_r119_SUM_10_, add_1_root_r119_SUM_11_,
         add_1_root_r119_SUM_12_, add_1_root_r119_SUM_13_,
         add_1_root_r119_SUM_14_, add_1_root_r119_SUM_15_,
         add_1_root_r119_SUM_16_, add_1_root_r119_SUM_17_,
         add_1_root_r119_SUM_18_, add_1_root_r119_SUM_19_,
         add_1_root_r119_SUM_20_, add_1_root_r119_SUM_21_,
         add_1_root_r119_SUM_22_, add_1_root_r119_SUM_23_,
         add_1_root_r119_A_2_, add_1_root_r119_A_3_, add_1_root_r119_A_4_,
         add_1_root_r119_A_5_, add_1_root_r119_A_6_, add_1_root_r119_A_7_,
         add_1_root_r119_A_8_, add_1_root_r119_A_9_, add_1_root_r119_A_10_,
         add_1_root_r119_A_11_, add_1_root_r119_A_12_, add_1_root_r119_A_13_,
         add_1_root_r119_A_14_, add_1_root_r119_A_15_, add_1_root_r119_A_16_,
         add_1_root_r119_A_17_, add_1_root_r119_A_18_, add_1_root_r119_A_19_,
         add_3_root_r119_carry_10_, add_3_root_r119_carry_11_,
         add_3_root_r119_carry_12_, add_3_root_r119_carry_13_,
         add_3_root_r119_carry_14_, add_3_root_r119_carry_15_,
         add_3_root_r119_carry_16_, add_3_root_r119_carry_17_,
         add_3_root_r119_carry_18_, add_3_root_r119_carry_3_,
         add_3_root_r119_carry_4_, add_3_root_r119_carry_5_,
         add_3_root_r119_carry_6_, add_3_root_r119_carry_7_,
         add_3_root_r119_carry_8_, add_3_root_r119_carry_9_,
         add_1_root_r112_carry_10_, add_1_root_r112_carry_11_,
         add_1_root_r112_carry_12_, add_1_root_r112_carry_13_,
         add_1_root_r112_carry_14_, add_1_root_r112_carry_15_,
         add_1_root_r112_carry_16_, add_1_root_r112_carry_17_,
         add_1_root_r112_carry_18_, add_1_root_r112_carry_19_,
         add_1_root_r112_carry_20_, add_1_root_r112_carry_5_,
         add_1_root_r112_carry_6_, add_1_root_r112_carry_7_,
         add_1_root_r112_carry_8_, add_1_root_r112_carry_9_,
         add_1_root_r112_SUM_1_, add_1_root_r112_SUM_2_,
         add_1_root_r112_SUM_3_, add_1_root_r112_SUM_4_,
         add_1_root_r112_SUM_5_, add_1_root_r112_SUM_6_,
         add_1_root_r112_SUM_7_, add_1_root_r112_SUM_8_,
         add_1_root_r112_SUM_9_, add_1_root_r112_SUM_10_,
         add_1_root_r112_SUM_11_, add_1_root_r112_SUM_12_,
         add_1_root_r112_SUM_13_, add_1_root_r112_SUM_14_,
         add_1_root_r112_SUM_15_, add_1_root_r112_SUM_16_,
         add_1_root_r112_SUM_17_, add_1_root_r112_SUM_18_,
         add_1_root_r112_SUM_19_, add_1_root_r112_SUM_20_,
         add_1_root_r112_SUM_21_, add_2_root_r115_carry_10_,
         add_2_root_r115_carry_11_, add_2_root_r115_carry_12_,
         add_2_root_r115_carry_13_, add_2_root_r115_carry_14_,
         add_2_root_r115_carry_15_, add_2_root_r115_carry_16_,
         add_2_root_r115_carry_17_, add_2_root_r115_carry_18_,
         add_2_root_r115_carry_19_, add_2_root_r115_carry_4_,
         add_2_root_r115_carry_5_, add_2_root_r115_carry_6_,
         add_2_root_r115_carry_7_, add_2_root_r115_carry_8_,
         add_2_root_r115_carry_9_, add_2_root_r115_SUM_3_,
         add_2_root_r115_SUM_4_, add_2_root_r115_SUM_5_,
         add_2_root_r115_SUM_6_, add_2_root_r115_SUM_7_,
         add_2_root_r115_SUM_8_, add_2_root_r115_SUM_9_,
         add_2_root_r115_SUM_10_, add_2_root_r115_SUM_11_,
         add_2_root_r115_SUM_12_, add_2_root_r115_SUM_13_,
         add_2_root_r115_SUM_14_, add_2_root_r115_SUM_15_,
         add_2_root_r115_SUM_16_, add_2_root_r115_SUM_17_,
         add_2_root_r115_SUM_18_, add_2_root_r115_SUM_19_,
         add_2_root_r115_SUM_20_, add_1_root_r115_carry_10_,
         add_1_root_r115_carry_11_, add_1_root_r115_carry_12_,
         add_1_root_r115_carry_13_, add_1_root_r115_carry_14_,
         add_1_root_r115_carry_15_, add_1_root_r115_carry_16_,
         add_1_root_r115_carry_17_, add_1_root_r115_carry_18_,
         add_1_root_r115_carry_19_, add_1_root_r115_carry_20_,
         add_1_root_r115_carry_21_, add_1_root_r115_carry_22_,
         add_1_root_r115_carry_7_, add_1_root_r115_carry_8_,
         add_1_root_r115_carry_9_, add_1_root_r115_SUM_6_,
         add_1_root_r115_SUM_7_, add_1_root_r115_SUM_8_,
         add_1_root_r115_SUM_9_, add_1_root_r115_SUM_10_,
         add_1_root_r115_SUM_11_, add_1_root_r115_SUM_12_,
         add_1_root_r115_SUM_13_, add_1_root_r115_SUM_14_,
         add_1_root_r115_SUM_15_, add_1_root_r115_SUM_16_,
         add_1_root_r115_SUM_17_, add_1_root_r115_SUM_18_,
         add_1_root_r115_SUM_19_, add_1_root_r115_SUM_20_,
         add_1_root_r115_SUM_21_, add_1_root_r115_SUM_22_,
         add_1_root_r115_SUM_23_, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234;
  wire   [16:0] in_17bit_b;
  wire   [23:8] neg_mul;
  wire   [16:10] sub_add_75_b0_carry;
  wire   [16:2] sub_add_54_b0_carry;
  wire   [22:7] add_1_root_r119_carry;

  multi16_7_DW01_add_0 add_0_root_r119 ( .A_22_(add_2_root_r119_SUM_22_), 
        .A_21_(add_2_root_r119_SUM_21_), .A_20_(add_2_root_r119_SUM_20_), 
        .A_19_(add_2_root_r119_SUM_19_), .A_18_(add_2_root_r119_SUM_18_), 
        .A_17_(add_2_root_r119_SUM_17_), .A_16_(add_2_root_r119_SUM_16_), 
        .A_15_(add_2_root_r119_SUM_15_), .A_14_(add_2_root_r119_SUM_14_), 
        .A_13_(add_2_root_r119_SUM_13_), .A_12_(add_2_root_r119_SUM_12_), 
        .A_11_(add_2_root_r119_SUM_11_), .A_10_(add_2_root_r119_SUM_10_), 
        .A_9_(add_2_root_r119_SUM_9_), .A_8_(add_2_root_r119_SUM_8_), .A_7_(
        add_2_root_r119_SUM_7_), .A_6_(add_2_root_r119_SUM_6_), .A_5_(
        add_2_root_r119_SUM_5_), .A_4_(in_17bit_b[0]), .B_23_(
        add_1_root_r119_SUM_23_), .B_22_(add_1_root_r119_SUM_22_), .B_21_(
        add_1_root_r119_SUM_21_), .B_20_(add_1_root_r119_SUM_20_), .B_19_(
        add_1_root_r119_SUM_19_), .B_18_(add_1_root_r119_SUM_18_), .B_17_(
        add_1_root_r119_SUM_17_), .B_16_(add_1_root_r119_SUM_16_), .B_15_(
        add_1_root_r119_SUM_15_), .B_14_(add_1_root_r119_SUM_14_), .B_13_(
        add_1_root_r119_SUM_13_), .B_12_(add_1_root_r119_SUM_12_), .B_11_(
        add_1_root_r119_SUM_11_), .B_10_(add_1_root_r119_SUM_10_), .B_9_(
        add_1_root_r119_SUM_9_), .B_8_(add_1_root_r119_SUM_8_), .B_7_(
        add_1_root_r119_SUM_7_), .B_6_(add_1_root_r119_SUM_6_), .B_5_(
        add_1_root_r119_A_5_), .B_4_(add_1_root_r119_A_4_), .SUM_23_(N363), 
        .SUM_22_(N362), .SUM_21_(N361), .SUM_20_(N360), .SUM_19_(N359), 
        .SUM_18_(N358), .SUM_17_(N357), .SUM_16_(N356), .SUM_15_(N355), 
        .SUM_14_(N354), .SUM_13_(N353), .SUM_12_(N352), .SUM_11_(N351), 
        .SUM_10_(N350), .SUM_9_(N349), .SUM_8_(N348), .SUM_7_(N347) );
  multi16_7_DW01_add_4 add_0_root_r112 ( .A_21_(n39), .A_20_(in_17bit_b[15]), 
        .A_19_(in_17bit_b[14]), .A_18_(in_17bit_b[13]), .A_17_(in_17bit_b[12]), 
        .A_16_(in_17bit_b[11]), .A_15_(in_17bit_b[10]), .A_14_(in_17bit_b[9]), 
        .A_13_(in_17bit_b[8]), .A_12_(in_17bit_b[7]), .A_11_(in_17bit_b[6]), 
        .A_10_(in_17bit_b[5]), .A_9_(in_17bit_b[4]), .A_8_(in_17bit_b[3]), 
        .A_7_(in_17bit_b[2]), .A_6_(in_17bit_b[1]), .A_5_(in_17bit_b[0]), 
        .B_21_(add_1_root_r112_SUM_21_), .B_20_(add_1_root_r112_SUM_20_), 
        .B_19_(add_1_root_r112_SUM_19_), .B_18_(add_1_root_r112_SUM_18_), 
        .B_17_(add_1_root_r112_SUM_17_), .B_16_(add_1_root_r112_SUM_16_), 
        .B_15_(add_1_root_r112_SUM_15_), .B_14_(add_1_root_r112_SUM_14_), 
        .B_13_(add_1_root_r112_SUM_13_), .B_12_(add_1_root_r112_SUM_12_), 
        .B_11_(add_1_root_r112_SUM_11_), .B_10_(add_1_root_r112_SUM_10_), 
        .B_9_(add_1_root_r112_SUM_9_), .B_8_(add_1_root_r112_SUM_8_), .B_7_(
        add_1_root_r112_SUM_7_), .B_6_(add_1_root_r112_SUM_6_), .B_5_(
        add_1_root_r112_SUM_5_), .SUM_22_(N123), .SUM_21_(N122), .SUM_20_(N121), .SUM_19_(N120), .SUM_18_(N119), .SUM_17_(N118), .SUM_16_(N117), .SUM_15_(
        N116), .SUM_14_(N115), .SUM_13_(N114), .SUM_12_(N113), .SUM_11_(N112), 
        .SUM_10_(N111), .SUM_9_(N110), .SUM_8_(N109), .SUM_7_(N108) );
  multi16_7_DW01_add_6 add_0_root_r115 ( .A_23_(add_1_root_r115_SUM_23_), 
        .A_22_(add_1_root_r115_SUM_22_), .A_21_(add_1_root_r115_SUM_21_), 
        .A_20_(add_1_root_r115_SUM_20_), .A_19_(add_1_root_r115_SUM_19_), 
        .A_18_(add_1_root_r115_SUM_18_), .A_17_(add_1_root_r115_SUM_17_), 
        .A_16_(add_1_root_r115_SUM_16_), .A_15_(add_1_root_r115_SUM_15_), 
        .A_14_(add_1_root_r115_SUM_14_), .A_13_(add_1_root_r115_SUM_13_), 
        .A_12_(add_1_root_r115_SUM_12_), .A_11_(add_1_root_r115_SUM_11_), 
        .A_10_(add_1_root_r115_SUM_10_), .A_9_(add_1_root_r115_SUM_9_), .A_8_(
        add_1_root_r115_SUM_8_), .A_7_(add_1_root_r115_SUM_7_), .A_6_(
        add_1_root_r115_SUM_6_), .A_5_(in_17bit_b[1]), .A_4_(in_17bit_b[0]), 
        .B_20_(add_2_root_r115_SUM_20_), .B_19_(add_2_root_r115_SUM_19_), 
        .B_18_(add_2_root_r115_SUM_18_), .B_17_(add_2_root_r115_SUM_17_), 
        .B_16_(add_2_root_r115_SUM_16_), .B_15_(add_2_root_r115_SUM_15_), 
        .B_14_(add_2_root_r115_SUM_14_), .B_13_(add_2_root_r115_SUM_13_), 
        .B_12_(add_2_root_r115_SUM_12_), .B_11_(add_2_root_r115_SUM_11_), 
        .B_10_(add_2_root_r115_SUM_10_), .B_9_(add_2_root_r115_SUM_9_), .B_8_(
        add_2_root_r115_SUM_8_), .B_7_(add_2_root_r115_SUM_7_), .B_6_(
        add_2_root_r115_SUM_6_), .B_5_(add_2_root_r115_SUM_5_), .B_4_(
        add_2_root_r115_SUM_4_), .SUM_23_(N221), .SUM_22_(N220), .SUM_21_(N219), .SUM_20_(N218), .SUM_19_(N217), .SUM_18_(N216), .SUM_17_(N215), .SUM_16_(
        N214), .SUM_15_(N213), .SUM_14_(N212), .SUM_13_(N211), .SUM_12_(N210), 
        .SUM_11_(N209), .SUM_10_(N208), .SUM_9_(N207), .SUM_8_(N206), .SUM_7_(
        N205) );
  TLATX1 neg_mul_reg_16_ ( .G(N446), .D(N456), .QN(n6) );
  TLATX1 neg_mul_reg_15_ ( .G(N446), .D(N455), .QN(n5) );
  TLATX1 neg_mul_reg_14_ ( .G(N446), .D(N454), .QN(n8) );
  TLATX1 neg_mul_reg_13_ ( .G(N446), .D(N453), .QN(n7) );
  TLATX1 neg_mul_reg_12_ ( .G(N446), .D(N452), .QN(n3) );
  TLATX1 neg_mul_reg_11_ ( .G(N446), .D(N451), .QN(n4) );
  TLATX1 neg_mul_reg_10_ ( .G(N446), .D(N450), .QN(n2) );
  TLATX1 neg_mul_reg_9_ ( .G(N446), .D(N449), .QN(n1) );
  TLATX1 neg_mul_reg_23_ ( .G(N446), .D(N463), .Q(neg_mul[23]), .QN(n16) );
  TLATX1 neg_mul_reg_22_ ( .G(N446), .D(N462), .Q(neg_mul[22]), .QN(n12) );
  TLATX1 neg_mul_reg_21_ ( .G(N446), .D(N461), .Q(neg_mul[21]), .QN(n13) );
  TLATX1 neg_mul_reg_20_ ( .G(N446), .D(N460), .QN(n14) );
  TLATX1 neg_mul_reg_19_ ( .G(N446), .D(N459), .Q(neg_mul[19]), .QN(n10) );
  TLATX1 neg_mul_reg_18_ ( .G(N446), .D(N458), .QN(n15) );
  TLATX1 neg_mul_reg_17_ ( .G(N446), .D(N457), .Q(neg_mul[17]), .QN(n11) );
  TLATX1 neg_mul_reg_8_ ( .G(N446), .D(N448), .Q(neg_mul[8]) );
  TLATX1 neg_mul_reg_7_ ( .G(N446), .D(N447), .Q(out[0]), .QN(n9) );
  NAND2X2 U2 ( .A(n24), .B(n63), .Y(n19) );
  NAND2X2 U3 ( .A(n24), .B(n61), .Y(n62) );
  INVX12 U4 ( .A(n67), .Y(n68) );
  INVX8 U5 ( .A(n42), .Y(n41) );
  INVX1 U6 ( .A(in_8bit[7]), .Y(n42) );
  INVX1 U7 ( .A(n63), .Y(n50) );
  INVX1 U8 ( .A(n18), .Y(n46) );
  INVX4 U9 ( .A(n41), .Y(n43) );
  AOI22X1 U10 ( .A0(N27), .A1(n46), .B0(in_17bit[14]), .B1(n18), .Y(n223) );
  XOR2X4 U11 ( .A(n17), .B(n5), .Y(out[8]) );
  OR2X4 U12 ( .A(n65), .B(n26), .Y(n17) );
  DLY1X1 U13 ( .A(n48), .Y(n18) );
  INVX8 U14 ( .A(n48), .Y(n37) );
  INVX2 U15 ( .A(n65), .Y(n66) );
  CLKBUFX8 U16 ( .A(in_17bit[16]), .Y(n38) );
  XNOR2X4 U17 ( .A(n38), .B(n43), .Y(n53) );
  XOR2X4 U18 ( .A(n37), .B(n41), .Y(n24) );
  MXI2X2 U19 ( .A(n15), .B(n34), .S0(n24), .Y(out[11]) );
  XNOR2X4 U20 ( .A(n43), .B(n48), .Y(n67) );
  NOR2X4 U21 ( .A(n65), .B(n58), .Y(n20) );
  NOR2X4 U22 ( .A(n67), .B(n9), .Y(n51) );
  NAND2X4 U23 ( .A(n56), .B(n55), .Y(n57) );
  XOR2X4 U24 ( .A(n41), .B(n38), .Y(n56) );
  XOR2X4 U25 ( .A(n37), .B(n43), .Y(n65) );
  INVX4 U26 ( .A(in_17bit[16]), .Y(n48) );
  XOR2X4 U27 ( .A(n8), .B(n19), .Y(out[7]) );
  NOR2X2 U28 ( .A(n65), .B(n32), .Y(n64) );
  AOI22XL U29 ( .A0(N355), .A1(n230), .B0(n94), .B1(in_17bit_b[8]), .Y(n207)
         );
  AOI22XL U30 ( .A0(N356), .A1(n230), .B0(n94), .B1(in_17bit_b[9]), .Y(n210)
         );
  AOI22XL U31 ( .A0(N357), .A1(n230), .B0(n94), .B1(in_17bit_b[10]), .Y(n213)
         );
  AOI22XL U32 ( .A0(N358), .A1(n230), .B0(n94), .B1(in_17bit_b[11]), .Y(n216)
         );
  AOI22XL U33 ( .A0(N120), .A1(n227), .B0(N217), .B1(n231), .Y(n218) );
  AOI22XL U34 ( .A0(N359), .A1(n230), .B0(n94), .B1(in_17bit_b[12]), .Y(n219)
         );
  AOI22XL U35 ( .A0(N121), .A1(n227), .B0(N218), .B1(n231), .Y(n221) );
  AOI22XL U36 ( .A0(N360), .A1(n230), .B0(n94), .B1(in_17bit_b[13]), .Y(n222)
         );
  AOI22XL U37 ( .A0(N122), .A1(n227), .B0(N219), .B1(n231), .Y(n224) );
  AOI22XL U38 ( .A0(N361), .A1(n230), .B0(n94), .B1(in_17bit_b[14]), .Y(n225)
         );
  AOI22XL U39 ( .A0(N123), .A1(n227), .B0(N220), .B1(n231), .Y(n228) );
  AOI22XL U40 ( .A0(N362), .A1(n230), .B0(n94), .B1(in_17bit_b[15]), .Y(n229)
         );
  INVX1 U41 ( .A(n223), .Y(in_17bit_b[14]) );
  INVX1 U42 ( .A(n184), .Y(in_17bit_b[1]) );
  INVX1 U43 ( .A(n220), .Y(in_17bit_b[13]) );
  INVX1 U44 ( .A(n196), .Y(in_17bit_b[5]) );
  INVX1 U45 ( .A(n199), .Y(in_17bit_b[6]) );
  INVX1 U46 ( .A(n202), .Y(in_17bit_b[7]) );
  INVX1 U47 ( .A(n205), .Y(in_17bit_b[8]) );
  INVX1 U48 ( .A(n208), .Y(in_17bit_b[9]) );
  INVX1 U49 ( .A(n211), .Y(in_17bit_b[10]) );
  INVX1 U50 ( .A(n214), .Y(in_17bit_b[11]) );
  INVX1 U51 ( .A(n217), .Y(in_17bit_b[12]) );
  INVX1 U52 ( .A(n187), .Y(in_17bit_b[2]) );
  INVX1 U53 ( .A(n193), .Y(in_17bit_b[4]) );
  INVX1 U54 ( .A(n190), .Y(in_17bit_b[3]) );
  XNOR2X4 U55 ( .A(n20), .B(n4), .Y(out[4]) );
  AOI21X1 U56 ( .A0(n21), .A1(n22), .B0(n227), .Y(n180) );
  NOR4XL U57 ( .A(in_8bit[4]), .B(in_8bit[5]), .C(in_8bit[6]), .D(n41), .Y(n21) );
  NOR4X1 U58 ( .A(in_8bit[1]), .B(in_8bit[0]), .C(in_8bit[2]), .D(in_8bit[3]), 
        .Y(n22) );
  AND4X1 U59 ( .A(in_8bit[1]), .B(n41), .C(n175), .D(n40), .Y(n23) );
  INVX1 U60 ( .A(n46), .Y(n47) );
  ADDFX2 U61 ( .A(n39), .B(in_17bit_b[12]), .CI(add_1_root_r112_carry_16_), 
        .CO(add_1_root_r112_carry_17_), .S(add_1_root_r112_SUM_16_) );
  ADDFX2 U62 ( .A(add_1_root_r119_A_19_), .B(in_17bit_b[13]), .CI(
        add_1_root_r119_carry[19]), .CO(add_1_root_r119_carry[20]), .S(
        add_1_root_r119_SUM_19_) );
  ADDFX2 U63 ( .A(n39), .B(in_17bit_b[15]), .CI(add_3_root_r119_carry_17_), 
        .CO(add_3_root_r119_carry_18_), .S(add_1_root_r119_A_17_) );
  ADDFX2 U64 ( .A(n39), .B(in_17bit_b[14]), .CI(add_2_root_r115_carry_17_), 
        .CO(add_2_root_r115_carry_18_), .S(add_2_root_r115_SUM_17_) );
  ADDFX2 U65 ( .A(n39), .B(in_17bit_b[14]), .CI(add_1_root_r115_carry_20_), 
        .CO(add_1_root_r115_carry_21_), .S(add_1_root_r115_SUM_20_) );
  ADDFX2 U66 ( .A(n39), .B(in_17bit_b[15]), .CI(add_2_root_r119_carry_20_), 
        .CO(add_2_root_r119_carry_21_), .S(add_2_root_r119_SUM_20_) );
  ADDFX2 U67 ( .A(in_17bit_b[3]), .B(in_17bit_b[1]), .CI(
        add_2_root_r115_carry_4_), .CO(add_2_root_r115_carry_5_), .S(
        add_2_root_r115_SUM_4_) );
  ADDFX2 U68 ( .A(in_17bit_b[4]), .B(in_17bit_b[2]), .CI(
        add_2_root_r115_carry_5_), .CO(add_2_root_r115_carry_6_), .S(
        add_2_root_r115_SUM_5_) );
  ADDFX2 U69 ( .A(in_17bit_b[5]), .B(in_17bit_b[1]), .CI(
        add_1_root_r112_carry_5_), .CO(add_1_root_r112_carry_6_), .S(
        add_1_root_r112_SUM_5_) );
  ADDFX2 U70 ( .A(in_17bit_b[6]), .B(in_17bit_b[5]), .CI(
        add_3_root_r119_carry_7_), .CO(add_3_root_r119_carry_8_), .S(
        add_1_root_r119_A_7_) );
  ADDFX2 U71 ( .A(in_17bit_b[6]), .B(in_17bit_b[2]), .CI(
        add_1_root_r112_carry_6_), .CO(add_1_root_r112_carry_7_), .S(
        add_1_root_r112_SUM_6_) );
  ADDFX2 U72 ( .A(in_17bit_b[3]), .B(in_17bit_b[1]), .CI(
        add_1_root_r115_carry_7_), .CO(add_1_root_r115_carry_8_), .S(
        add_1_root_r115_SUM_7_) );
  ADDFX2 U73 ( .A(in_17bit_b[7]), .B(in_17bit_b[6]), .CI(
        add_3_root_r119_carry_8_), .CO(add_3_root_r119_carry_9_), .S(
        add_1_root_r119_A_8_) );
  ADDFX2 U74 ( .A(add_1_root_r119_A_7_), .B(in_17bit_b[1]), .CI(
        add_1_root_r119_carry[7]), .CO(add_1_root_r119_carry[8]), .S(
        add_1_root_r119_SUM_7_) );
  ADDFX2 U75 ( .A(in_17bit_b[2]), .B(in_17bit_b[1]), .CI(
        add_2_root_r119_carry_6_), .CO(add_2_root_r119_carry_7_), .S(
        add_2_root_r119_SUM_6_) );
  ADDFX2 U76 ( .A(in_17bit_b[4]), .B(in_17bit_b[2]), .CI(
        add_1_root_r115_carry_8_), .CO(add_1_root_r115_carry_9_), .S(
        add_1_root_r115_SUM_8_) );
  ADDFX2 U77 ( .A(in_17bit_b[8]), .B(in_17bit_b[7]), .CI(
        add_3_root_r119_carry_9_), .CO(add_3_root_r119_carry_10_), .S(
        add_1_root_r119_A_9_) );
  ADDFX2 U78 ( .A(add_1_root_r119_A_8_), .B(in_17bit_b[2]), .CI(
        add_1_root_r119_carry[8]), .CO(add_1_root_r119_carry[9]), .S(
        add_1_root_r119_SUM_8_) );
  ADDFX2 U79 ( .A(in_17bit_b[3]), .B(in_17bit_b[2]), .CI(
        add_2_root_r119_carry_7_), .CO(add_2_root_r119_carry_8_), .S(
        add_2_root_r119_SUM_7_) );
  ADDFX2 U80 ( .A(in_17bit_b[6]), .B(in_17bit_b[4]), .CI(
        add_2_root_r115_carry_7_), .CO(add_2_root_r115_carry_8_), .S(
        add_2_root_r115_SUM_7_) );
  ADDFX2 U81 ( .A(in_17bit_b[9]), .B(in_17bit_b[8]), .CI(
        add_3_root_r119_carry_10_), .CO(add_3_root_r119_carry_11_), .S(
        add_1_root_r119_A_10_) );
  ADDFX2 U82 ( .A(in_17bit_b[7]), .B(in_17bit_b[5]), .CI(
        add_2_root_r115_carry_8_), .CO(add_2_root_r115_carry_9_), .S(
        add_2_root_r115_SUM_8_) );
  ADDFX2 U83 ( .A(in_17bit_b[9]), .B(in_17bit_b[5]), .CI(
        add_1_root_r112_carry_9_), .CO(add_1_root_r112_carry_10_), .S(
        add_1_root_r112_SUM_9_) );
  ADDFX2 U84 ( .A(in_17bit_b[10]), .B(in_17bit_b[9]), .CI(
        add_3_root_r119_carry_11_), .CO(add_3_root_r119_carry_12_), .S(
        add_1_root_r119_A_11_) );
  ADDFX2 U85 ( .A(in_17bit_b[6]), .B(in_17bit_b[4]), .CI(
        add_1_root_r115_carry_10_), .CO(add_1_root_r115_carry_11_), .S(
        add_1_root_r115_SUM_10_) );
  ADDFX2 U86 ( .A(add_1_root_r119_A_10_), .B(in_17bit_b[4]), .CI(
        add_1_root_r119_carry[10]), .CO(add_1_root_r119_carry[11]), .S(
        add_1_root_r119_SUM_10_) );
  ADDFX2 U87 ( .A(in_17bit_b[5]), .B(in_17bit_b[4]), .CI(
        add_2_root_r119_carry_9_), .CO(add_2_root_r119_carry_10_), .S(
        add_2_root_r119_SUM_9_) );
  ADDFX2 U88 ( .A(in_17bit_b[8]), .B(in_17bit_b[6]), .CI(
        add_2_root_r115_carry_9_), .CO(add_2_root_r115_carry_10_), .S(
        add_2_root_r115_SUM_9_) );
  ADDFX2 U89 ( .A(in_17bit_b[10]), .B(in_17bit_b[6]), .CI(
        add_1_root_r112_carry_10_), .CO(add_1_root_r112_carry_11_), .S(
        add_1_root_r112_SUM_10_) );
  ADDFX2 U90 ( .A(in_17bit_b[7]), .B(in_17bit_b[5]), .CI(
        add_1_root_r115_carry_11_), .CO(add_1_root_r115_carry_12_), .S(
        add_1_root_r115_SUM_11_) );
  ADDFX2 U91 ( .A(in_17bit_b[11]), .B(in_17bit_b[10]), .CI(
        add_3_root_r119_carry_12_), .CO(add_3_root_r119_carry_13_), .S(
        add_1_root_r119_A_12_) );
  ADDFX2 U92 ( .A(add_1_root_r119_A_11_), .B(in_17bit_b[5]), .CI(
        add_1_root_r119_carry[11]), .CO(add_1_root_r119_carry[12]), .S(
        add_1_root_r119_SUM_11_) );
  ADDFX2 U93 ( .A(in_17bit_b[6]), .B(in_17bit_b[5]), .CI(
        add_2_root_r119_carry_10_), .CO(add_2_root_r119_carry_11_), .S(
        add_2_root_r119_SUM_10_) );
  ADDFX2 U94 ( .A(in_17bit_b[9]), .B(in_17bit_b[7]), .CI(
        add_2_root_r115_carry_10_), .CO(add_2_root_r115_carry_11_), .S(
        add_2_root_r115_SUM_10_) );
  ADDFX2 U95 ( .A(in_17bit_b[11]), .B(in_17bit_b[7]), .CI(
        add_1_root_r112_carry_11_), .CO(add_1_root_r112_carry_12_), .S(
        add_1_root_r112_SUM_11_) );
  ADDFX2 U96 ( .A(in_17bit_b[8]), .B(in_17bit_b[6]), .CI(
        add_1_root_r115_carry_12_), .CO(add_1_root_r115_carry_13_), .S(
        add_1_root_r115_SUM_12_) );
  ADDFX2 U97 ( .A(in_17bit_b[12]), .B(in_17bit_b[11]), .CI(
        add_3_root_r119_carry_13_), .CO(add_3_root_r119_carry_14_), .S(
        add_1_root_r119_A_13_) );
  ADDFX2 U98 ( .A(add_1_root_r119_A_12_), .B(in_17bit_b[6]), .CI(
        add_1_root_r119_carry[12]), .CO(add_1_root_r119_carry[13]), .S(
        add_1_root_r119_SUM_12_) );
  ADDFX2 U99 ( .A(in_17bit_b[7]), .B(in_17bit_b[6]), .CI(
        add_2_root_r119_carry_11_), .CO(add_2_root_r119_carry_12_), .S(
        add_2_root_r119_SUM_11_) );
  ADDFX2 U100 ( .A(in_17bit_b[10]), .B(in_17bit_b[8]), .CI(
        add_2_root_r115_carry_11_), .CO(add_2_root_r115_carry_12_), .S(
        add_2_root_r115_SUM_11_) );
  ADDFX2 U101 ( .A(in_17bit_b[12]), .B(in_17bit_b[8]), .CI(
        add_1_root_r112_carry_12_), .CO(add_1_root_r112_carry_13_), .S(
        add_1_root_r112_SUM_12_) );
  ADDFX2 U102 ( .A(in_17bit_b[9]), .B(in_17bit_b[7]), .CI(
        add_1_root_r115_carry_13_), .CO(add_1_root_r115_carry_14_), .S(
        add_1_root_r115_SUM_13_) );
  ADDFX2 U103 ( .A(in_17bit_b[13]), .B(in_17bit_b[12]), .CI(
        add_3_root_r119_carry_14_), .CO(add_3_root_r119_carry_15_), .S(
        add_1_root_r119_A_14_) );
  ADDFX2 U104 ( .A(add_1_root_r119_A_13_), .B(in_17bit_b[7]), .CI(
        add_1_root_r119_carry[13]), .CO(add_1_root_r119_carry[14]), .S(
        add_1_root_r119_SUM_13_) );
  ADDFX2 U105 ( .A(in_17bit_b[8]), .B(in_17bit_b[7]), .CI(
        add_2_root_r119_carry_12_), .CO(add_2_root_r119_carry_13_), .S(
        add_2_root_r119_SUM_12_) );
  ADDFX2 U106 ( .A(in_17bit_b[11]), .B(in_17bit_b[9]), .CI(
        add_2_root_r115_carry_12_), .CO(add_2_root_r115_carry_13_), .S(
        add_2_root_r115_SUM_12_) );
  ADDFX2 U107 ( .A(in_17bit_b[13]), .B(in_17bit_b[9]), .CI(
        add_1_root_r112_carry_13_), .CO(add_1_root_r112_carry_14_), .S(
        add_1_root_r112_SUM_13_) );
  ADDFX2 U108 ( .A(in_17bit_b[10]), .B(in_17bit_b[8]), .CI(
        add_1_root_r115_carry_14_), .CO(add_1_root_r115_carry_15_), .S(
        add_1_root_r115_SUM_14_) );
  ADDFX2 U109 ( .A(in_17bit_b[14]), .B(in_17bit_b[13]), .CI(
        add_3_root_r119_carry_15_), .CO(add_3_root_r119_carry_16_), .S(
        add_1_root_r119_A_15_) );
  ADDFX2 U110 ( .A(add_1_root_r119_A_14_), .B(in_17bit_b[8]), .CI(
        add_1_root_r119_carry[14]), .CO(add_1_root_r119_carry[15]), .S(
        add_1_root_r119_SUM_14_) );
  ADDFX2 U111 ( .A(in_17bit_b[9]), .B(in_17bit_b[8]), .CI(
        add_2_root_r119_carry_13_), .CO(add_2_root_r119_carry_14_), .S(
        add_2_root_r119_SUM_13_) );
  ADDFX2 U112 ( .A(in_17bit_b[12]), .B(in_17bit_b[10]), .CI(
        add_2_root_r115_carry_13_), .CO(add_2_root_r115_carry_14_), .S(
        add_2_root_r115_SUM_13_) );
  ADDFX2 U113 ( .A(in_17bit_b[11]), .B(in_17bit_b[9]), .CI(
        add_1_root_r115_carry_15_), .CO(add_1_root_r115_carry_16_), .S(
        add_1_root_r115_SUM_15_) );
  ADDFX2 U114 ( .A(add_1_root_r119_A_15_), .B(in_17bit_b[9]), .CI(
        add_1_root_r119_carry[15]), .CO(add_1_root_r119_carry[16]), .S(
        add_1_root_r119_SUM_15_) );
  ADDFX2 U115 ( .A(in_17bit_b[3]), .B(in_17bit_b[2]), .CI(
        add_3_root_r119_carry_4_), .CO(add_3_root_r119_carry_5_), .S(
        add_1_root_r119_A_4_) );
  ADDFX2 U116 ( .A(in_17bit_b[2]), .B(in_17bit_b[1]), .CI(
        add_3_root_r119_carry_3_), .CO(add_3_root_r119_carry_4_), .S(
        add_1_root_r119_A_3_) );
  ADDFX2 U117 ( .A(in_17bit_b[13]), .B(in_17bit_b[11]), .CI(
        add_2_root_r115_carry_14_), .CO(add_2_root_r115_carry_15_), .S(
        add_2_root_r115_SUM_14_) );
  ADDFX2 U118 ( .A(in_17bit_b[15]), .B(in_17bit_b[11]), .CI(
        add_1_root_r112_carry_15_), .CO(add_1_root_r112_carry_16_), .S(
        add_1_root_r112_SUM_15_) );
  ADDFX2 U119 ( .A(in_17bit_b[12]), .B(in_17bit_b[10]), .CI(
        add_1_root_r115_carry_16_), .CO(add_1_root_r115_carry_17_), .S(
        add_1_root_r115_SUM_16_) );
  ADDFX2 U120 ( .A(add_1_root_r119_A_16_), .B(in_17bit_b[10]), .CI(
        add_1_root_r119_carry[16]), .CO(add_1_root_r119_carry[17]), .S(
        add_1_root_r119_SUM_16_) );
  ADDFX2 U121 ( .A(in_17bit_b[11]), .B(in_17bit_b[10]), .CI(
        add_2_root_r119_carry_15_), .CO(add_2_root_r119_carry_16_), .S(
        add_2_root_r119_SUM_15_) );
  ADDFX2 U122 ( .A(in_17bit_b[14]), .B(in_17bit_b[12]), .CI(
        add_2_root_r115_carry_15_), .CO(add_2_root_r115_carry_16_), .S(
        add_2_root_r115_SUM_15_) );
  ADDFX2 U123 ( .A(in_17bit_b[13]), .B(in_17bit_b[11]), .CI(
        add_1_root_r115_carry_17_), .CO(add_1_root_r115_carry_18_), .S(
        add_1_root_r115_SUM_17_) );
  ADDFX2 U124 ( .A(add_1_root_r119_A_17_), .B(in_17bit_b[11]), .CI(
        add_1_root_r119_carry[17]), .CO(add_1_root_r119_carry[18]), .S(
        add_1_root_r119_SUM_17_) );
  ADDFX2 U125 ( .A(in_17bit_b[12]), .B(in_17bit_b[11]), .CI(
        add_2_root_r119_carry_16_), .CO(add_2_root_r119_carry_17_), .S(
        add_2_root_r119_SUM_16_) );
  ADDFX2 U126 ( .A(in_17bit_b[15]), .B(in_17bit_b[13]), .CI(
        add_2_root_r115_carry_16_), .CO(add_2_root_r115_carry_17_), .S(
        add_2_root_r115_SUM_16_) );
  ADDFX2 U127 ( .A(in_17bit_b[14]), .B(in_17bit_b[12]), .CI(
        add_1_root_r115_carry_18_), .CO(add_1_root_r115_carry_19_), .S(
        add_1_root_r115_SUM_18_) );
  ADDFX2 U128 ( .A(in_17bit_b[15]), .B(in_17bit_b[13]), .CI(
        add_1_root_r115_carry_19_), .CO(add_1_root_r115_carry_20_), .S(
        add_1_root_r115_SUM_19_) );
  ADDFX2 U129 ( .A(in_17bit_b[13]), .B(in_17bit_b[12]), .CI(
        add_2_root_r119_carry_17_), .CO(add_2_root_r119_carry_18_), .S(
        add_2_root_r119_SUM_17_) );
  ADDFX2 U130 ( .A(in_17bit_b[14]), .B(in_17bit_b[13]), .CI(
        add_2_root_r119_carry_18_), .CO(add_2_root_r119_carry_19_), .S(
        add_2_root_r119_SUM_18_) );
  ADDFX2 U131 ( .A(in_17bit_b[5]), .B(in_17bit_b[3]), .CI(
        add_2_root_r115_carry_6_), .CO(add_2_root_r115_carry_7_), .S(
        add_2_root_r115_SUM_6_) );
  ADDFX2 U132 ( .A(in_17bit_b[7]), .B(in_17bit_b[3]), .CI(
        add_1_root_r112_carry_7_), .CO(add_1_root_r112_carry_8_), .S(
        add_1_root_r112_SUM_7_) );
  ADDFX2 U133 ( .A(in_17bit_b[14]), .B(in_17bit_b[10]), .CI(
        add_1_root_r112_carry_14_), .CO(add_1_root_r112_carry_15_), .S(
        add_1_root_r112_SUM_14_) );
  ADDFX2 U134 ( .A(in_17bit_b[8]), .B(in_17bit_b[4]), .CI(
        add_1_root_r112_carry_8_), .CO(add_1_root_r112_carry_9_), .S(
        add_1_root_r112_SUM_8_) );
  ADDFX2 U135 ( .A(in_17bit_b[5]), .B(in_17bit_b[3]), .CI(
        add_1_root_r115_carry_9_), .CO(add_1_root_r115_carry_10_), .S(
        add_1_root_r115_SUM_9_) );
  ADDFX2 U136 ( .A(add_1_root_r119_A_9_), .B(in_17bit_b[3]), .CI(
        add_1_root_r119_carry[9]), .CO(add_1_root_r119_carry[10]), .S(
        add_1_root_r119_SUM_9_) );
  ADDFX2 U137 ( .A(in_17bit_b[10]), .B(in_17bit_b[9]), .CI(
        add_2_root_r119_carry_14_), .CO(add_2_root_r119_carry_15_), .S(
        add_2_root_r119_SUM_14_) );
  ADDFX2 U138 ( .A(in_17bit_b[15]), .B(in_17bit_b[14]), .CI(
        add_3_root_r119_carry_16_), .CO(add_3_root_r119_carry_17_), .S(
        add_1_root_r119_A_16_) );
  ADDFX2 U139 ( .A(in_17bit_b[4]), .B(in_17bit_b[3]), .CI(
        add_2_root_r119_carry_8_), .CO(add_2_root_r119_carry_9_), .S(
        add_2_root_r119_SUM_8_) );
  ADDFX2 U140 ( .A(add_1_root_r119_A_18_), .B(in_17bit_b[12]), .CI(
        add_1_root_r119_carry[18]), .CO(add_1_root_r119_carry[19]), .S(
        add_1_root_r119_SUM_18_) );
  ADDFX2 U141 ( .A(in_17bit_b[4]), .B(in_17bit_b[3]), .CI(
        add_3_root_r119_carry_5_), .CO(add_3_root_r119_carry_6_), .S(
        add_1_root_r119_A_5_) );
  ADDFX2 U142 ( .A(in_17bit_b[5]), .B(in_17bit_b[4]), .CI(
        add_3_root_r119_carry_6_), .CO(add_3_root_r119_carry_7_), .S(
        add_1_root_r119_A_6_) );
  ADDFX2 U143 ( .A(in_17bit_b[15]), .B(in_17bit_b[14]), .CI(
        add_2_root_r119_carry_19_), .CO(add_2_root_r119_carry_20_), .S(
        add_2_root_r119_SUM_19_) );
  BUFX3 U144 ( .A(in_17bit_b[16]), .Y(n39) );
  INVX1 U145 ( .A(n234), .Y(in_17bit_b[16]) );
  NAND2XL U146 ( .A(N29), .B(n46), .Y(n234) );
  CLKINVX3 U147 ( .A(n181), .Y(in_17bit_b[0]) );
  INVX1 U148 ( .A(n94), .Y(n233) );
  OAI21XL U149 ( .A0(n233), .A1(n234), .B0(n232), .Y(N463) );
  AOI22XL U150 ( .A0(N221), .A1(n231), .B0(N363), .B1(n230), .Y(n232) );
  CLKINVX3 U151 ( .A(n226), .Y(in_17bit_b[15]) );
  NAND2X1 U152 ( .A(n31), .B(in_8bit[1]), .Y(n69) );
  INVX1 U153 ( .A(in_8bit[0]), .Y(n40) );
  INVX1 U154 ( .A(in_8bit[2]), .Y(n44) );
  INVX1 U155 ( .A(in_8bit[5]), .Y(n45) );
  AOI22XL U156 ( .A0(N28), .A1(n46), .B0(in_17bit[15]), .B1(n47), .Y(n226) );
  AOI22XL U157 ( .A0(N18), .A1(n46), .B0(in_17bit[5]), .B1(n47), .Y(n196) );
  AOI22XL U158 ( .A0(N19), .A1(n46), .B0(in_17bit[6]), .B1(n18), .Y(n199) );
  AOI22XL U159 ( .A0(N20), .A1(n46), .B0(in_17bit[7]), .B1(n18), .Y(n202) );
  AOI22XL U160 ( .A0(N21), .A1(n46), .B0(in_17bit[8]), .B1(n18), .Y(n205) );
  AOI22XL U161 ( .A0(N22), .A1(n46), .B0(in_17bit[9]), .B1(n47), .Y(n208) );
  AOI22XL U162 ( .A0(N23), .A1(n46), .B0(in_17bit[10]), .B1(n47), .Y(n211) );
  AOI22XL U163 ( .A0(N24), .A1(n46), .B0(in_17bit[11]), .B1(n47), .Y(n214) );
  AOI22XL U164 ( .A0(N25), .A1(n46), .B0(in_17bit[12]), .B1(n47), .Y(n217) );
  AOI22XL U165 ( .A0(N26), .A1(n46), .B0(in_17bit[13]), .B1(n47), .Y(n220) );
  NOR3X1 U166 ( .A(n44), .B(n95), .C(n40), .Y(n179) );
  AOI22X1 U167 ( .A0(in_17bit[0]), .A1(n46), .B0(in_17bit[0]), .B1(n47), .Y(
        n181) );
  AOI22X1 U168 ( .A0(N14), .A1(n46), .B0(in_17bit[1]), .B1(n18), .Y(n184) );
  AOI22X1 U169 ( .A0(N15), .A1(n46), .B0(in_17bit[2]), .B1(n47), .Y(n187) );
  AOI22X1 U170 ( .A0(N16), .A1(n46), .B0(in_17bit[3]), .B1(n47), .Y(n190) );
  AOI22X1 U171 ( .A0(N17), .A1(n46), .B0(in_17bit[4]), .B1(n18), .Y(n193) );
  NOR2X1 U172 ( .A(in_8bit[0]), .B(n75), .Y(n25) );
  INVX1 U173 ( .A(n49), .Y(n58) );
  NAND2BX1 U174 ( .AN(n55), .B(n2), .Y(n49) );
  AND2X2 U175 ( .A(n50), .B(n8), .Y(n26) );
  AOI21X1 U176 ( .A0(n74), .A1(n23), .B0(n28), .Y(n27) );
  INVX1 U177 ( .A(n27), .Y(n230) );
  AND2X2 U178 ( .A(n25), .B(n33), .Y(n28) );
  AOI21X1 U179 ( .A0(n33), .A1(n23), .B0(n30), .Y(n29) );
  INVX1 U180 ( .A(n29), .Y(n231) );
  AND2X2 U181 ( .A(n25), .B(n74), .Y(n30) );
  NAND2X1 U182 ( .A(n58), .B(n4), .Y(n59) );
  NAND2BX1 U183 ( .AN(n59), .B(n3), .Y(n61) );
  NAND2BX1 U184 ( .AN(n61), .B(n7), .Y(n63) );
  OAI2BB1X1 U185 ( .A0N(n178), .A1N(n31), .B0(n76), .Y(n94) );
  NAND3BX1 U186 ( .AN(n75), .B(n179), .C(in_8bit[5]), .Y(n76) );
  AND3X1 U187 ( .A(n41), .B(n70), .C(n45), .Y(n31) );
  NAND2BX1 U188 ( .AN(n52), .B(n1), .Y(n55) );
  AND2X2 U189 ( .A(n26), .B(n5), .Y(n32) );
  NOR2XL U190 ( .A(n41), .B(n70), .Y(n71) );
  INVX1 U191 ( .A(in_17bit[13]), .Y(n90) );
  INVX1 U192 ( .A(in_17bit[3]), .Y(n80) );
  INVX1 U193 ( .A(in_17bit[4]), .Y(n81) );
  INVX1 U194 ( .A(in_17bit[5]), .Y(n82) );
  INVX1 U195 ( .A(in_17bit[6]), .Y(n83) );
  INVX1 U196 ( .A(in_17bit[7]), .Y(n84) );
  INVX1 U197 ( .A(in_17bit[8]), .Y(n85) );
  INVX1 U198 ( .A(in_17bit[9]), .Y(n86) );
  INVX1 U199 ( .A(in_17bit[10]), .Y(n87) );
  INVX1 U200 ( .A(in_17bit[11]), .Y(n88) );
  INVX1 U201 ( .A(in_17bit[12]), .Y(n89) );
  INVX1 U202 ( .A(in_17bit[14]), .Y(n91) );
  INVX1 U203 ( .A(in_17bit[15]), .Y(n92) );
  INVX1 U204 ( .A(in_17bit[1]), .Y(n78) );
  INVX1 U205 ( .A(in_17bit[2]), .Y(n79) );
  INVX1 U206 ( .A(in_17bit[0]), .Y(n77) );
  AND3X2 U207 ( .A(in_8bit[2]), .B(n95), .C(in_8bit[5]), .Y(n33) );
  NAND2X1 U208 ( .A(n183), .B(n182), .Y(N447) );
  AOI22X1 U209 ( .A0(N108), .A1(n227), .B0(N205), .B1(n231), .Y(n182) );
  AOI22X1 U210 ( .A0(N347), .A1(n230), .B0(n94), .B1(in_17bit_b[0]), .Y(n183)
         );
  NAND2X1 U211 ( .A(n186), .B(n185), .Y(N448) );
  AOI22X1 U212 ( .A0(N109), .A1(n227), .B0(N206), .B1(n231), .Y(n185) );
  AOI22X1 U213 ( .A0(N348), .A1(n230), .B0(n94), .B1(n93), .Y(n186) );
  INVX1 U214 ( .A(n184), .Y(n93) );
  NAND2X1 U215 ( .A(n189), .B(n188), .Y(N449) );
  AOI22X1 U216 ( .A0(N110), .A1(n227), .B0(N207), .B1(n231), .Y(n188) );
  AOI22X1 U217 ( .A0(N349), .A1(n230), .B0(n94), .B1(in_17bit_b[2]), .Y(n189)
         );
  NAND2X1 U218 ( .A(n192), .B(n191), .Y(N450) );
  AOI22X1 U219 ( .A0(N111), .A1(n227), .B0(N208), .B1(n231), .Y(n191) );
  AOI22X1 U220 ( .A0(N350), .A1(n230), .B0(n94), .B1(in_17bit_b[3]), .Y(n192)
         );
  NAND2X1 U221 ( .A(n195), .B(n194), .Y(N451) );
  AOI22X1 U222 ( .A0(N112), .A1(n227), .B0(N209), .B1(n231), .Y(n194) );
  AOI22X1 U223 ( .A0(N351), .A1(n230), .B0(n94), .B1(in_17bit_b[4]), .Y(n195)
         );
  NAND2X1 U224 ( .A(n198), .B(n197), .Y(N452) );
  AOI22X1 U225 ( .A0(N113), .A1(n227), .B0(N210), .B1(n231), .Y(n197) );
  AOI22X1 U226 ( .A0(N352), .A1(n230), .B0(n94), .B1(in_17bit_b[5]), .Y(n198)
         );
  NAND2X1 U227 ( .A(n201), .B(n200), .Y(N453) );
  AOI22X1 U228 ( .A0(N114), .A1(n227), .B0(N211), .B1(n231), .Y(n200) );
  AOI22X1 U229 ( .A0(N353), .A1(n230), .B0(n94), .B1(in_17bit_b[6]), .Y(n201)
         );
  NAND2X1 U230 ( .A(n204), .B(n203), .Y(N454) );
  AOI22X1 U231 ( .A0(N115), .A1(n227), .B0(N212), .B1(n231), .Y(n203) );
  AOI22X1 U232 ( .A0(N354), .A1(n230), .B0(n94), .B1(in_17bit_b[7]), .Y(n204)
         );
  NAND2X1 U233 ( .A(n207), .B(n206), .Y(N455) );
  AOI22X1 U234 ( .A0(N116), .A1(n227), .B0(N213), .B1(n231), .Y(n206) );
  NAND2X1 U235 ( .A(n210), .B(n209), .Y(N456) );
  AOI22X1 U236 ( .A0(N117), .A1(n227), .B0(N214), .B1(n231), .Y(n209) );
  NAND2X1 U237 ( .A(n213), .B(n212), .Y(N457) );
  AOI22X1 U238 ( .A0(N118), .A1(n227), .B0(N215), .B1(n231), .Y(n212) );
  NAND2X1 U239 ( .A(n216), .B(n215), .Y(N458) );
  AOI22X1 U240 ( .A0(N119), .A1(n227), .B0(N216), .B1(n231), .Y(n215) );
  NAND2X1 U241 ( .A(n219), .B(n218), .Y(N459) );
  NAND2X1 U242 ( .A(n222), .B(n221), .Y(N460) );
  NAND2X1 U243 ( .A(n225), .B(n224), .Y(N461) );
  NAND2X1 U244 ( .A(n229), .B(n228), .Y(N462) );
  MX2X4 U245 ( .A(neg_mul[17]), .B(N475), .S0(n66), .Y(out[10]) );
  XNOR2X1 U246 ( .A(n15), .B(sub_add_75_b0_carry[11]), .Y(n34) );
  XNOR2X1 U247 ( .A(n14), .B(sub_add_75_b0_carry[13]), .Y(n35) );
  MX2X4 U248 ( .A(neg_mul[19]), .B(N477), .S0(n68), .Y(out[12]) );
  MX2X1 U249 ( .A(neg_mul[21]), .B(N479), .S0(n68), .Y(out[14]) );
  MX2X1 U250 ( .A(neg_mul[22]), .B(N480), .S0(n68), .Y(out[15]) );
  MX2X1 U251 ( .A(neg_mul[23]), .B(N481), .S0(n68), .Y(out[16]) );
  NAND4BBX1 U252 ( .AN(n230), .BN(n231), .C(n180), .D(n233), .Y(N446) );
  NOR4BX1 U253 ( .AN(n177), .B(n40), .C(in_8bit[1]), .D(in_8bit[2]), .Y(n178)
         );
  NOR2X1 U254 ( .A(in_8bit[6]), .B(in_8bit[3]), .Y(n177) );
  NAND4BXL U255 ( .AN(n41), .B(in_8bit[6]), .C(in_8bit[1]), .D(in_8bit[4]), 
        .Y(n75) );
  NAND2X1 U256 ( .A(n73), .B(n72), .Y(n227) );
  NAND3BX1 U257 ( .AN(n69), .B(n179), .C(in_8bit[6]), .Y(n73) );
  NAND3X1 U258 ( .A(n178), .B(in_8bit[5]), .C(n71), .Y(n72) );
  OR2X2 U259 ( .A(out[0]), .B(neg_mul[8]), .Y(n52) );
  INVX1 U260 ( .A(n176), .Y(n74) );
  NAND3BX1 U261 ( .AN(in_8bit[5]), .B(n44), .C(in_8bit[3]), .Y(n176) );
  NOR2X1 U262 ( .A(in_8bit[6]), .B(in_8bit[4]), .Y(n175) );
  INVX1 U263 ( .A(in_8bit[4]), .Y(n70) );
  INVX1 U264 ( .A(in_8bit[3]), .Y(n95) );
  XOR2X4 U265 ( .A(n51), .B(neg_mul[8]), .Y(out[1]) );
  NAND2X4 U266 ( .A(n53), .B(n52), .Y(n54) );
  XOR2X4 U267 ( .A(n54), .B(n1), .Y(out[2]) );
  XOR2X4 U268 ( .A(n57), .B(n2), .Y(out[3]) );
  NAND2X4 U269 ( .A(n24), .B(n59), .Y(n60) );
  XOR2X4 U270 ( .A(n60), .B(n3), .Y(out[5]) );
  XOR2X4 U271 ( .A(n7), .B(n62), .Y(out[6]) );
  XNOR2X4 U272 ( .A(n64), .B(n6), .Y(out[9]) );
  MXI2X4 U273 ( .A(n14), .B(n35), .S0(n68), .Y(out[13]) );
  AND2X1 U274 ( .A(add_1_root_r112_carry_20_), .B(n39), .Y(
        add_1_root_r112_SUM_21_) );
  XOR2X1 U275 ( .A(n39), .B(add_1_root_r112_carry_20_), .Y(
        add_1_root_r112_SUM_20_) );
  AND2X1 U276 ( .A(add_1_root_r112_carry_19_), .B(in_17bit_b[15]), .Y(
        add_1_root_r112_carry_20_) );
  XOR2X1 U277 ( .A(in_17bit_b[15]), .B(add_1_root_r112_carry_19_), .Y(
        add_1_root_r112_SUM_19_) );
  AND2X1 U278 ( .A(add_1_root_r112_carry_18_), .B(in_17bit_b[14]), .Y(
        add_1_root_r112_carry_19_) );
  XOR2X1 U279 ( .A(in_17bit_b[14]), .B(add_1_root_r112_carry_18_), .Y(
        add_1_root_r112_SUM_18_) );
  AND2X1 U280 ( .A(add_1_root_r112_carry_17_), .B(in_17bit_b[13]), .Y(
        add_1_root_r112_carry_18_) );
  XOR2X1 U281 ( .A(in_17bit_b[13]), .B(add_1_root_r112_carry_17_), .Y(
        add_1_root_r112_SUM_17_) );
  AND2X1 U282 ( .A(add_2_root_r119_carry_21_), .B(n39), .Y(
        add_2_root_r119_SUM_22_) );
  XOR2X1 U283 ( .A(n39), .B(add_2_root_r119_carry_21_), .Y(
        add_2_root_r119_SUM_21_) );
  AND2X1 U284 ( .A(in_17bit_b[1]), .B(in_17bit_b[0]), .Y(
        add_2_root_r119_carry_6_) );
  XOR2X1 U285 ( .A(in_17bit_b[0]), .B(in_17bit_b[1]), .Y(
        add_2_root_r119_SUM_5_) );
  AND2X1 U286 ( .A(add_1_root_r119_carry[22]), .B(n39), .Y(
        add_1_root_r119_SUM_23_) );
  XOR2X1 U287 ( .A(n39), .B(add_1_root_r119_carry[22]), .Y(
        add_1_root_r119_SUM_22_) );
  AND2X1 U288 ( .A(add_1_root_r119_carry[21]), .B(in_17bit_b[15]), .Y(
        add_1_root_r119_carry[22]) );
  XOR2X1 U289 ( .A(in_17bit_b[15]), .B(add_1_root_r119_carry[21]), .Y(
        add_1_root_r119_SUM_21_) );
  AND2X1 U290 ( .A(add_1_root_r119_carry[20]), .B(in_17bit_b[14]), .Y(
        add_1_root_r119_carry[21]) );
  XOR2X1 U291 ( .A(in_17bit_b[14]), .B(add_1_root_r119_carry[20]), .Y(
        add_1_root_r119_SUM_20_) );
  AND2X1 U292 ( .A(add_1_root_r119_A_6_), .B(in_17bit_b[0]), .Y(
        add_1_root_r119_carry[7]) );
  XOR2X1 U293 ( .A(in_17bit_b[0]), .B(add_1_root_r119_A_6_), .Y(
        add_1_root_r119_SUM_6_) );
  AND2X1 U294 ( .A(add_3_root_r119_carry_18_), .B(n39), .Y(
        add_1_root_r119_A_19_) );
  XOR2X1 U295 ( .A(n39), .B(add_3_root_r119_carry_18_), .Y(
        add_1_root_r119_A_18_) );
  AND2X1 U296 ( .A(in_17bit_b[1]), .B(in_17bit_b[0]), .Y(
        add_3_root_r119_carry_3_) );
  XOR2X1 U297 ( .A(in_17bit_b[0]), .B(in_17bit_b[1]), .Y(add_1_root_r119_A_2_)
         );
  AND2X1 U298 ( .A(add_2_root_r115_carry_19_), .B(n39), .Y(
        add_2_root_r115_SUM_20_) );
  XOR2X1 U299 ( .A(n39), .B(add_2_root_r115_carry_19_), .Y(
        add_2_root_r115_SUM_19_) );
  AND2X1 U300 ( .A(add_2_root_r115_carry_18_), .B(in_17bit_b[15]), .Y(
        add_2_root_r115_carry_19_) );
  XOR2X1 U301 ( .A(in_17bit_b[15]), .B(add_2_root_r115_carry_18_), .Y(
        add_2_root_r115_SUM_18_) );
  AND2X1 U302 ( .A(in_17bit_b[2]), .B(in_17bit_b[0]), .Y(
        add_2_root_r115_carry_4_) );
  XOR2X1 U303 ( .A(in_17bit_b[0]), .B(in_17bit_b[2]), .Y(
        add_2_root_r115_SUM_3_) );
  AND2X1 U304 ( .A(add_1_root_r115_carry_22_), .B(n39), .Y(
        add_1_root_r115_SUM_23_) );
  XOR2X1 U305 ( .A(n39), .B(add_1_root_r115_carry_22_), .Y(
        add_1_root_r115_SUM_22_) );
  AND2X1 U306 ( .A(add_1_root_r115_carry_21_), .B(in_17bit_b[15]), .Y(
        add_1_root_r115_carry_22_) );
  XOR2X1 U307 ( .A(in_17bit_b[15]), .B(add_1_root_r115_carry_21_), .Y(
        add_1_root_r115_SUM_21_) );
  AND2X1 U308 ( .A(in_17bit_b[2]), .B(in_17bit_b[0]), .Y(
        add_1_root_r115_carry_7_) );
  XOR2X1 U309 ( .A(in_17bit_b[0]), .B(in_17bit_b[2]), .Y(
        add_1_root_r115_SUM_6_) );
  XOR2X1 U310 ( .A(n18), .B(sub_add_54_b0_carry[16]), .Y(N29) );
  AND2X1 U311 ( .A(sub_add_54_b0_carry[15]), .B(n92), .Y(
        sub_add_54_b0_carry[16]) );
  XOR2X1 U312 ( .A(n92), .B(sub_add_54_b0_carry[15]), .Y(N28) );
  AND2X1 U313 ( .A(sub_add_54_b0_carry[14]), .B(n91), .Y(
        sub_add_54_b0_carry[15]) );
  XOR2X1 U314 ( .A(n91), .B(sub_add_54_b0_carry[14]), .Y(N27) );
  AND2X1 U315 ( .A(sub_add_54_b0_carry[13]), .B(n90), .Y(
        sub_add_54_b0_carry[14]) );
  XOR2X1 U316 ( .A(n90), .B(sub_add_54_b0_carry[13]), .Y(N26) );
  AND2X1 U317 ( .A(sub_add_54_b0_carry[12]), .B(n89), .Y(
        sub_add_54_b0_carry[13]) );
  XOR2X1 U318 ( .A(n89), .B(sub_add_54_b0_carry[12]), .Y(N25) );
  AND2X1 U319 ( .A(sub_add_54_b0_carry[11]), .B(n88), .Y(
        sub_add_54_b0_carry[12]) );
  XOR2X1 U320 ( .A(n88), .B(sub_add_54_b0_carry[11]), .Y(N24) );
  AND2X1 U321 ( .A(sub_add_54_b0_carry[10]), .B(n87), .Y(
        sub_add_54_b0_carry[11]) );
  XOR2X1 U322 ( .A(n87), .B(sub_add_54_b0_carry[10]), .Y(N23) );
  AND2X1 U323 ( .A(sub_add_54_b0_carry[9]), .B(n86), .Y(
        sub_add_54_b0_carry[10]) );
  XOR2X1 U324 ( .A(n86), .B(sub_add_54_b0_carry[9]), .Y(N22) );
  AND2X1 U325 ( .A(sub_add_54_b0_carry[8]), .B(n85), .Y(sub_add_54_b0_carry[9]) );
  XOR2X1 U326 ( .A(n85), .B(sub_add_54_b0_carry[8]), .Y(N21) );
  AND2X1 U327 ( .A(sub_add_54_b0_carry[7]), .B(n84), .Y(sub_add_54_b0_carry[8]) );
  XOR2X1 U328 ( .A(n84), .B(sub_add_54_b0_carry[7]), .Y(N20) );
  AND2X1 U329 ( .A(sub_add_54_b0_carry[6]), .B(n83), .Y(sub_add_54_b0_carry[7]) );
  XOR2X1 U330 ( .A(n83), .B(sub_add_54_b0_carry[6]), .Y(N19) );
  AND2X1 U331 ( .A(sub_add_54_b0_carry[5]), .B(n82), .Y(sub_add_54_b0_carry[6]) );
  XOR2X1 U332 ( .A(n82), .B(sub_add_54_b0_carry[5]), .Y(N18) );
  AND2X1 U333 ( .A(sub_add_54_b0_carry[4]), .B(n81), .Y(sub_add_54_b0_carry[5]) );
  XOR2X1 U334 ( .A(n81), .B(sub_add_54_b0_carry[4]), .Y(N17) );
  AND2X1 U335 ( .A(sub_add_54_b0_carry[3]), .B(n80), .Y(sub_add_54_b0_carry[4]) );
  XOR2X1 U336 ( .A(n80), .B(sub_add_54_b0_carry[3]), .Y(N16) );
  AND2X1 U337 ( .A(sub_add_54_b0_carry[2]), .B(n79), .Y(sub_add_54_b0_carry[3]) );
  XOR2X1 U338 ( .A(n79), .B(sub_add_54_b0_carry[2]), .Y(N15) );
  AND2X1 U339 ( .A(n77), .B(n78), .Y(sub_add_54_b0_carry[2]) );
  XOR2X1 U340 ( .A(n78), .B(n77), .Y(N14) );
  XOR2X1 U341 ( .A(n16), .B(sub_add_75_b0_carry[16]), .Y(N481) );
  AND2X1 U342 ( .A(sub_add_75_b0_carry[15]), .B(n12), .Y(
        sub_add_75_b0_carry[16]) );
  XOR2X1 U343 ( .A(n12), .B(sub_add_75_b0_carry[15]), .Y(N480) );
  AND2X1 U344 ( .A(sub_add_75_b0_carry[14]), .B(n13), .Y(
        sub_add_75_b0_carry[15]) );
  XOR2X1 U345 ( .A(n13), .B(sub_add_75_b0_carry[14]), .Y(N479) );
  AND2X1 U346 ( .A(sub_add_75_b0_carry[13]), .B(n14), .Y(
        sub_add_75_b0_carry[14]) );
  AND2X1 U347 ( .A(sub_add_75_b0_carry[12]), .B(n10), .Y(
        sub_add_75_b0_carry[13]) );
  XOR2X1 U348 ( .A(n10), .B(sub_add_75_b0_carry[12]), .Y(N477) );
  AND2X1 U349 ( .A(sub_add_75_b0_carry[11]), .B(n15), .Y(
        sub_add_75_b0_carry[12]) );
  AND2X1 U350 ( .A(sub_add_75_b0_carry[10]), .B(n11), .Y(
        sub_add_75_b0_carry[11]) );
  XOR2X1 U351 ( .A(n11), .B(sub_add_75_b0_carry[10]), .Y(N475) );
  AND2X1 U352 ( .A(n32), .B(n6), .Y(sub_add_75_b0_carry[10]) );
  AND2X1 U353 ( .A(in_17bit_b[0]), .B(in_17bit_b[4]), .Y(
        add_1_root_r112_carry_5_) );
endmodule


module multi16_6_DW01_add_0 ( A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, 
        A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, 
        A_4_, B_23_, B_22_, B_21_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, 
        B_14_, B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, 
        SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, 
        SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, 
        SUM_7_ );
  input A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_,
         A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, B_23_, B_22_,
         B_21_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_,
         B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_;
  output SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_,
         SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_,
         SUM_8_, SUM_7_;
  wire   n1, n2, n3, n4;
  wire   [23:7] carry;

  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry[7]), .CO(carry[8]), .S(SUM_7_)
         );
  ADDFX2 U1_21 ( .A(A_21_), .B(B_21_), .CI(carry[21]), .CO(carry[22]), .S(
        SUM_21_) );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry[20]), .CO(carry[21]), .S(
        SUM_20_) );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry[19]), .CO(carry[20]), .S(
        SUM_19_) );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry[18]), .CO(carry[19]), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry[17]), .CO(carry[18]), .S(
        SUM_17_) );
  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry[16]), .CO(carry[17]), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry[15]), .CO(carry[16]), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry[14]), .CO(carry[15]), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry[13]), .CO(carry[14]), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry[12]), .CO(carry[13]), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry[11]), .CO(carry[12]), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry[10]), .CO(carry[11]), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry[9]), .CO(carry[10]), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry[8]), .CO(carry[9]), .S(SUM_8_)
         );
  ADDFX2 U1_22 ( .A(A_22_), .B(B_22_), .CI(carry[22]), .CO(carry[23]), .S(
        SUM_22_) );
  AND2X2 U1 ( .A(A_4_), .B(B_4_), .Y(n1) );
  XOR2X1 U2 ( .A(B_23_), .B(carry[23]), .Y(SUM_23_) );
  OAI2BB1X1 U3 ( .A0N(n2), .A1N(A_6_), .B0(n3), .Y(carry[7]) );
  OAI21XL U4 ( .A0(A_6_), .A1(n2), .B0(B_6_), .Y(n3) );
  OAI2BB1X1 U5 ( .A0N(n1), .A1N(A_5_), .B0(n4), .Y(n2) );
  OAI21XL U6 ( .A0(A_5_), .A1(n1), .B0(B_5_), .Y(n4) );
endmodule


module multi16_6_DW01_add_4 ( A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, 
        A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, 
        B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, 
        B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, SUM_22_, SUM_21_, SUM_20_, 
        SUM_19_, SUM_18_, SUM_17_, SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, 
        SUM_11_, SUM_10_, SUM_9_, SUM_8_, SUM_7_ );
  input A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_,
         A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, B_20_, B_19_,
         B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, B_10_, B_9_,
         B_8_, B_7_, B_6_, B_5_;
  output SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_,
         SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_,
         SUM_7_;
  wire   carry_21_, carry_20_, carry_19_, carry_18_, carry_17_, carry_16_,
         carry_15_, carry_14_, carry_13_, carry_12_, carry_11_, carry_10_,
         carry_9_, carry_8_, carry_7_, n1;

  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry_16_), .CO(carry_17_), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry_15_), .CO(carry_16_), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry_14_), .CO(carry_15_), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry_13_), .CO(carry_14_), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry_12_), .CO(carry_13_), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry_11_), .CO(carry_12_), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry_10_), .CO(carry_11_), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry_9_), .CO(carry_10_), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry_8_), .CO(carry_9_), .S(SUM_8_)
         );
  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry_7_), .CO(carry_8_), .S(SUM_7_)
         );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry_20_), .CO(carry_21_), .S(
        SUM_20_) );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry_19_), .CO(carry_20_), .S(
        SUM_19_) );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry_18_), .CO(carry_19_), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry_17_), .CO(carry_18_), .S(
        SUM_17_) );
  ADDFX2 U1_21 ( .A(A_21_), .B(B_21_), .CI(carry_21_), .CO(SUM_22_), .S(
        SUM_21_) );
  OAI2BB1X1 U1 ( .A0N(A_6_), .A1N(B_6_), .B0(n1), .Y(carry_7_) );
  OAI211X1 U2 ( .A0(B_6_), .A1(A_6_), .B0(A_5_), .C0(B_5_), .Y(n1) );
endmodule


module multi16_6_DW01_add_6 ( A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, 
        A_16_, A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, 
        A_6_, A_5_, A_4_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, 
        B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, 
        SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, 
        SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, 
        SUM_7_ );
  input A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_,
         A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, B_20_,
         B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, B_10_,
         B_9_, B_8_, B_7_, B_6_, B_5_, B_4_;
  output SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_,
         SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_,
         SUM_8_, SUM_7_;
  wire   n1, n2, n3, n4, n5, n6;
  wire   [21:7] carry;

  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry[7]), .CO(carry[8]), .S(SUM_7_)
         );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry[18]), .CO(carry[19]), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry[17]), .CO(carry[18]), .S(
        SUM_17_) );
  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry[16]), .CO(carry[17]), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry[15]), .CO(carry[16]), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry[14]), .CO(carry[15]), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry[13]), .CO(carry[14]), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry[12]), .CO(carry[13]), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry[11]), .CO(carry[12]), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry[10]), .CO(carry[11]), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry[9]), .CO(carry[10]), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry[8]), .CO(carry[9]), .S(SUM_8_)
         );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry[19]), .CO(carry[20]), .S(
        SUM_19_) );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry[20]), .CO(carry[21]), .S(
        SUM_20_) );
  AND2X2 U1 ( .A(A_22_), .B(n2), .Y(n1) );
  AND2X2 U2 ( .A(A_21_), .B(carry[21]), .Y(n2) );
  AND2X2 U3 ( .A(A_4_), .B(B_4_), .Y(n3) );
  XOR2X1 U4 ( .A(A_23_), .B(n1), .Y(SUM_23_) );
  XOR2X1 U5 ( .A(A_21_), .B(carry[21]), .Y(SUM_21_) );
  XOR2X1 U6 ( .A(A_22_), .B(n2), .Y(SUM_22_) );
  OAI2BB1X1 U7 ( .A0N(n4), .A1N(A_6_), .B0(n5), .Y(carry[7]) );
  OAI21XL U8 ( .A0(A_6_), .A1(n4), .B0(B_6_), .Y(n5) );
  OAI2BB1X1 U9 ( .A0N(n3), .A1N(A_5_), .B0(n6), .Y(n4) );
  OAI21XL U10 ( .A0(A_5_), .A1(n3), .B0(B_5_), .Y(n6) );
endmodule


module multi16_6 ( in_17bit, in_8bit, out );
  input [16:0] in_17bit;
  input [7:0] in_8bit;
  output [16:0] out;
  wire   n254, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26,
         N27, N28, N29, N108, N109, N110, N111, N112, N113, N114, N115, N116,
         N117, N118, N119, N120, N121, N122, N123, N205, N206, N207, N208,
         N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, N219,
         N220, N221, N347, N348, N349, N350, N351, N352, N353, N354, N355,
         N356, N357, N358, N359, N360, N361, N362, N363, N446, N447, N448,
         N449, N450, N451, N452, N453, N454, N455, N456, N457, N458, N459,
         N460, N461, N462, N463, N477, N478, N479, N480,
         add_2_root_r119_carry_10_, add_2_root_r119_carry_11_,
         add_2_root_r119_carry_12_, add_2_root_r119_carry_13_,
         add_2_root_r119_carry_14_, add_2_root_r119_carry_15_,
         add_2_root_r119_carry_16_, add_2_root_r119_carry_17_,
         add_2_root_r119_carry_18_, add_2_root_r119_carry_19_,
         add_2_root_r119_carry_20_, add_2_root_r119_carry_21_,
         add_2_root_r119_carry_6_, add_2_root_r119_carry_7_,
         add_2_root_r119_carry_8_, add_2_root_r119_carry_9_,
         add_2_root_r119_SUM_5_, add_2_root_r119_SUM_6_,
         add_2_root_r119_SUM_7_, add_2_root_r119_SUM_8_,
         add_2_root_r119_SUM_9_, add_2_root_r119_SUM_10_,
         add_2_root_r119_SUM_11_, add_2_root_r119_SUM_12_,
         add_2_root_r119_SUM_13_, add_2_root_r119_SUM_14_,
         add_2_root_r119_SUM_15_, add_2_root_r119_SUM_16_,
         add_2_root_r119_SUM_17_, add_2_root_r119_SUM_18_,
         add_2_root_r119_SUM_19_, add_2_root_r119_SUM_20_,
         add_2_root_r119_SUM_21_, add_2_root_r119_SUM_22_,
         add_1_root_r119_SUM_6_, add_1_root_r119_SUM_7_,
         add_1_root_r119_SUM_8_, add_1_root_r119_SUM_9_,
         add_1_root_r119_SUM_10_, add_1_root_r119_SUM_11_,
         add_1_root_r119_SUM_12_, add_1_root_r119_SUM_13_,
         add_1_root_r119_SUM_14_, add_1_root_r119_SUM_15_,
         add_1_root_r119_SUM_16_, add_1_root_r119_SUM_17_,
         add_1_root_r119_SUM_18_, add_1_root_r119_SUM_19_,
         add_1_root_r119_SUM_20_, add_1_root_r119_SUM_21_,
         add_1_root_r119_SUM_22_, add_1_root_r119_SUM_23_,
         add_1_root_r119_A_2_, add_1_root_r119_A_3_, add_1_root_r119_A_4_,
         add_1_root_r119_A_5_, add_1_root_r119_A_6_, add_1_root_r119_A_7_,
         add_1_root_r119_A_8_, add_1_root_r119_A_9_, add_1_root_r119_A_10_,
         add_1_root_r119_A_11_, add_1_root_r119_A_12_, add_1_root_r119_A_13_,
         add_1_root_r119_A_14_, add_1_root_r119_A_15_, add_1_root_r119_A_16_,
         add_1_root_r119_A_17_, add_1_root_r119_A_18_, add_1_root_r119_A_19_,
         add_3_root_r119_carry_10_, add_3_root_r119_carry_11_,
         add_3_root_r119_carry_12_, add_3_root_r119_carry_13_,
         add_3_root_r119_carry_14_, add_3_root_r119_carry_15_,
         add_3_root_r119_carry_16_, add_3_root_r119_carry_17_,
         add_3_root_r119_carry_18_, add_3_root_r119_carry_3_,
         add_3_root_r119_carry_4_, add_3_root_r119_carry_5_,
         add_3_root_r119_carry_6_, add_3_root_r119_carry_7_,
         add_3_root_r119_carry_8_, add_3_root_r119_carry_9_,
         add_1_root_r112_carry_10_, add_1_root_r112_carry_11_,
         add_1_root_r112_carry_12_, add_1_root_r112_carry_13_,
         add_1_root_r112_carry_14_, add_1_root_r112_carry_15_,
         add_1_root_r112_carry_16_, add_1_root_r112_carry_17_,
         add_1_root_r112_carry_18_, add_1_root_r112_carry_19_,
         add_1_root_r112_carry_20_, add_1_root_r112_carry_5_,
         add_1_root_r112_carry_6_, add_1_root_r112_carry_7_,
         add_1_root_r112_carry_8_, add_1_root_r112_carry_9_,
         add_1_root_r112_SUM_1_, add_1_root_r112_SUM_2_,
         add_1_root_r112_SUM_3_, add_1_root_r112_SUM_4_,
         add_1_root_r112_SUM_5_, add_1_root_r112_SUM_6_,
         add_1_root_r112_SUM_7_, add_1_root_r112_SUM_8_,
         add_1_root_r112_SUM_9_, add_1_root_r112_SUM_10_,
         add_1_root_r112_SUM_11_, add_1_root_r112_SUM_12_,
         add_1_root_r112_SUM_13_, add_1_root_r112_SUM_14_,
         add_1_root_r112_SUM_15_, add_1_root_r112_SUM_16_,
         add_1_root_r112_SUM_17_, add_1_root_r112_SUM_18_,
         add_1_root_r112_SUM_19_, add_1_root_r112_SUM_20_,
         add_1_root_r112_SUM_21_, add_2_root_r115_carry_10_,
         add_2_root_r115_carry_11_, add_2_root_r115_carry_12_,
         add_2_root_r115_carry_13_, add_2_root_r115_carry_14_,
         add_2_root_r115_carry_15_, add_2_root_r115_carry_16_,
         add_2_root_r115_carry_17_, add_2_root_r115_carry_18_,
         add_2_root_r115_carry_19_, add_2_root_r115_carry_4_,
         add_2_root_r115_carry_5_, add_2_root_r115_carry_6_,
         add_2_root_r115_carry_7_, add_2_root_r115_carry_8_,
         add_2_root_r115_carry_9_, add_2_root_r115_SUM_3_,
         add_2_root_r115_SUM_4_, add_2_root_r115_SUM_5_,
         add_2_root_r115_SUM_6_, add_2_root_r115_SUM_7_,
         add_2_root_r115_SUM_8_, add_2_root_r115_SUM_9_,
         add_2_root_r115_SUM_10_, add_2_root_r115_SUM_11_,
         add_2_root_r115_SUM_12_, add_2_root_r115_SUM_13_,
         add_2_root_r115_SUM_14_, add_2_root_r115_SUM_15_,
         add_2_root_r115_SUM_16_, add_2_root_r115_SUM_17_,
         add_2_root_r115_SUM_18_, add_2_root_r115_SUM_19_,
         add_2_root_r115_SUM_20_, add_1_root_r115_carry_10_,
         add_1_root_r115_carry_11_, add_1_root_r115_carry_12_,
         add_1_root_r115_carry_13_, add_1_root_r115_carry_14_,
         add_1_root_r115_carry_15_, add_1_root_r115_carry_16_,
         add_1_root_r115_carry_17_, add_1_root_r115_carry_18_,
         add_1_root_r115_carry_19_, add_1_root_r115_carry_20_,
         add_1_root_r115_carry_21_, add_1_root_r115_carry_22_,
         add_1_root_r115_carry_7_, add_1_root_r115_carry_8_,
         add_1_root_r115_carry_9_, add_1_root_r115_SUM_6_,
         add_1_root_r115_SUM_7_, add_1_root_r115_SUM_8_,
         add_1_root_r115_SUM_9_, add_1_root_r115_SUM_10_,
         add_1_root_r115_SUM_11_, add_1_root_r115_SUM_12_,
         add_1_root_r115_SUM_13_, add_1_root_r115_SUM_14_,
         add_1_root_r115_SUM_15_, add_1_root_r115_SUM_16_,
         add_1_root_r115_SUM_17_, add_1_root_r115_SUM_18_,
         add_1_root_r115_SUM_19_, add_1_root_r115_SUM_20_,
         add_1_root_r115_SUM_21_, add_1_root_r115_SUM_22_,
         add_1_root_r115_SUM_23_, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n158, n160, n161, n162, n163, n164, n167, n168,
         n170, n171, n172, n173, n174, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253;
  wire   [16:0] in_17bit_b;
  wire   [23:8] neg_mul;
  wire   [15:10] sub_add_75_b0_carry;
  wire   [16:2] sub_add_54_b0_carry;
  wire   [22:7] add_1_root_r119_carry;

  multi16_6_DW01_add_0 add_0_root_r119 ( .A_22_(add_2_root_r119_SUM_22_), 
        .A_21_(add_2_root_r119_SUM_21_), .A_20_(add_2_root_r119_SUM_20_), 
        .A_19_(add_2_root_r119_SUM_19_), .A_18_(add_2_root_r119_SUM_18_), 
        .A_17_(add_2_root_r119_SUM_17_), .A_16_(add_2_root_r119_SUM_16_), 
        .A_15_(add_2_root_r119_SUM_15_), .A_14_(add_2_root_r119_SUM_14_), 
        .A_13_(add_2_root_r119_SUM_13_), .A_12_(add_2_root_r119_SUM_12_), 
        .A_11_(add_2_root_r119_SUM_11_), .A_10_(add_2_root_r119_SUM_10_), 
        .A_9_(add_2_root_r119_SUM_9_), .A_8_(add_2_root_r119_SUM_8_), .A_7_(
        add_2_root_r119_SUM_7_), .A_6_(add_2_root_r119_SUM_6_), .A_5_(
        add_2_root_r119_SUM_5_), .A_4_(in_17bit_b[0]), .B_23_(
        add_1_root_r119_SUM_23_), .B_22_(add_1_root_r119_SUM_22_), .B_21_(
        add_1_root_r119_SUM_21_), .B_20_(add_1_root_r119_SUM_20_), .B_19_(
        add_1_root_r119_SUM_19_), .B_18_(add_1_root_r119_SUM_18_), .B_17_(
        add_1_root_r119_SUM_17_), .B_16_(add_1_root_r119_SUM_16_), .B_15_(
        add_1_root_r119_SUM_15_), .B_14_(add_1_root_r119_SUM_14_), .B_13_(
        add_1_root_r119_SUM_13_), .B_12_(add_1_root_r119_SUM_12_), .B_11_(
        add_1_root_r119_SUM_11_), .B_10_(add_1_root_r119_SUM_10_), .B_9_(
        add_1_root_r119_SUM_9_), .B_8_(add_1_root_r119_SUM_8_), .B_7_(
        add_1_root_r119_SUM_7_), .B_6_(add_1_root_r119_SUM_6_), .B_5_(
        add_1_root_r119_A_5_), .B_4_(add_1_root_r119_A_4_), .SUM_23_(N363), 
        .SUM_22_(N362), .SUM_21_(N361), .SUM_20_(N360), .SUM_19_(N359), 
        .SUM_18_(N358), .SUM_17_(N357), .SUM_16_(N356), .SUM_15_(N355), 
        .SUM_14_(N354), .SUM_13_(N353), .SUM_12_(N352), .SUM_11_(N351), 
        .SUM_10_(N350), .SUM_9_(N349), .SUM_8_(N348), .SUM_7_(N347) );
  multi16_6_DW01_add_4 add_0_root_r112 ( .A_21_(n42), .A_20_(in_17bit_b[15]), 
        .A_19_(in_17bit_b[14]), .A_18_(in_17bit_b[13]), .A_17_(in_17bit_b[12]), 
        .A_16_(in_17bit_b[11]), .A_15_(in_17bit_b[10]), .A_14_(in_17bit_b[9]), 
        .A_13_(in_17bit_b[8]), .A_12_(in_17bit_b[7]), .A_11_(in_17bit_b[6]), 
        .A_10_(in_17bit_b[5]), .A_9_(in_17bit_b[4]), .A_8_(in_17bit_b[3]), 
        .A_7_(in_17bit_b[2]), .A_6_(in_17bit_b[1]), .A_5_(in_17bit_b[0]), 
        .B_21_(add_1_root_r112_SUM_21_), .B_20_(add_1_root_r112_SUM_20_), 
        .B_19_(add_1_root_r112_SUM_19_), .B_18_(add_1_root_r112_SUM_18_), 
        .B_17_(add_1_root_r112_SUM_17_), .B_16_(add_1_root_r112_SUM_16_), 
        .B_15_(add_1_root_r112_SUM_15_), .B_14_(add_1_root_r112_SUM_14_), 
        .B_13_(add_1_root_r112_SUM_13_), .B_12_(add_1_root_r112_SUM_12_), 
        .B_11_(add_1_root_r112_SUM_11_), .B_10_(add_1_root_r112_SUM_10_), 
        .B_9_(add_1_root_r112_SUM_9_), .B_8_(add_1_root_r112_SUM_8_), .B_7_(
        add_1_root_r112_SUM_7_), .B_6_(add_1_root_r112_SUM_6_), .B_5_(
        add_1_root_r112_SUM_5_), .SUM_22_(N123), .SUM_21_(N122), .SUM_20_(N121), .SUM_19_(N120), .SUM_18_(N119), .SUM_17_(N118), .SUM_16_(N117), .SUM_15_(
        N116), .SUM_14_(N115), .SUM_13_(N114), .SUM_12_(N113), .SUM_11_(N112), 
        .SUM_10_(N111), .SUM_9_(N110), .SUM_8_(N109), .SUM_7_(N108) );
  multi16_6_DW01_add_6 add_0_root_r115 ( .A_23_(add_1_root_r115_SUM_23_), 
        .A_22_(add_1_root_r115_SUM_22_), .A_21_(add_1_root_r115_SUM_21_), 
        .A_20_(add_1_root_r115_SUM_20_), .A_19_(add_1_root_r115_SUM_19_), 
        .A_18_(add_1_root_r115_SUM_18_), .A_17_(add_1_root_r115_SUM_17_), 
        .A_16_(add_1_root_r115_SUM_16_), .A_15_(add_1_root_r115_SUM_15_), 
        .A_14_(add_1_root_r115_SUM_14_), .A_13_(add_1_root_r115_SUM_13_), 
        .A_12_(add_1_root_r115_SUM_12_), .A_11_(add_1_root_r115_SUM_11_), 
        .A_10_(add_1_root_r115_SUM_10_), .A_9_(add_1_root_r115_SUM_9_), .A_8_(
        add_1_root_r115_SUM_8_), .A_7_(add_1_root_r115_SUM_7_), .A_6_(
        add_1_root_r115_SUM_6_), .A_5_(in_17bit_b[1]), .A_4_(in_17bit_b[0]), 
        .B_20_(add_2_root_r115_SUM_20_), .B_19_(add_2_root_r115_SUM_19_), 
        .B_18_(add_2_root_r115_SUM_18_), .B_17_(add_2_root_r115_SUM_17_), 
        .B_16_(add_2_root_r115_SUM_16_), .B_15_(add_2_root_r115_SUM_15_), 
        .B_14_(add_2_root_r115_SUM_14_), .B_13_(add_2_root_r115_SUM_13_), 
        .B_12_(add_2_root_r115_SUM_12_), .B_11_(add_2_root_r115_SUM_11_), 
        .B_10_(add_2_root_r115_SUM_10_), .B_9_(add_2_root_r115_SUM_9_), .B_8_(
        add_2_root_r115_SUM_8_), .B_7_(add_2_root_r115_SUM_7_), .B_6_(
        add_2_root_r115_SUM_6_), .B_5_(add_2_root_r115_SUM_5_), .B_4_(
        add_2_root_r115_SUM_4_), .SUM_23_(N221), .SUM_22_(N220), .SUM_21_(N219), .SUM_20_(N218), .SUM_19_(N217), .SUM_18_(N216), .SUM_17_(N215), .SUM_16_(
        N214), .SUM_15_(N213), .SUM_14_(N212), .SUM_13_(N211), .SUM_12_(N210), 
        .SUM_11_(N209), .SUM_10_(N208), .SUM_9_(N207), .SUM_8_(N206), .SUM_7_(
        N205) );
  TLATX1 neg_mul_reg_16_ ( .G(N446), .D(N456), .QN(n7) );
  TLATX1 neg_mul_reg_15_ ( .G(N446), .D(N455), .QN(n2) );
  TLATX1 neg_mul_reg_14_ ( .G(N446), .D(N454), .QN(n3) );
  TLATX1 neg_mul_reg_13_ ( .G(N446), .D(N453), .QN(n6) );
  TLATX1 neg_mul_reg_12_ ( .G(N446), .D(N452), .QN(n5) );
  TLATX1 neg_mul_reg_11_ ( .G(N446), .D(N451), .QN(n4) );
  TLATX1 neg_mul_reg_23_ ( .G(N446), .D(N463), .Q(neg_mul[23]), .QN(n1) );
  TLATX1 neg_mul_reg_22_ ( .G(N446), .D(N462), .Q(neg_mul[22]), .QN(n9) );
  TLATX1 neg_mul_reg_21_ ( .G(N446), .D(N461), .Q(neg_mul[21]), .QN(n13) );
  TLATX1 neg_mul_reg_20_ ( .G(N446), .D(N460), .Q(neg_mul[20]), .QN(n11) );
  TLATX1 neg_mul_reg_19_ ( .G(N446), .D(N459), .Q(neg_mul[19]), .QN(n12) );
  TLATX1 neg_mul_reg_18_ ( .G(N446), .D(N458), .QN(n15) );
  TLATX1 neg_mul_reg_17_ ( .G(N446), .D(N457), .QN(n14) );
  TLATX1 neg_mul_reg_9_ ( .G(N446), .D(N449), .Q(neg_mul[9]), .QN(n8) );
  TLATX1 neg_mul_reg_10_ ( .G(N446), .D(N450), .Q(neg_mul[10]), .QN(n10) );
  TLATX1 neg_mul_reg_8_ ( .G(N446), .D(N448), .Q(neg_mul[8]), .QN(n16) );
  TLATX1 neg_mul_reg_7_ ( .G(N446), .D(N447), .Q(out[0]) );
  XNOR2X2 U2 ( .A(n52), .B(n44), .Y(n78) );
  CLKINVX8 U3 ( .A(n46), .Y(n45) );
  AOI2BB2X1 U4 ( .B0(n60), .B1(n44), .A0N(n45), .A1N(neg_mul[8]), .Y(n61) );
  XNOR2X1 U5 ( .A(n52), .B(n44), .Y(n81) );
  INVX1 U6 ( .A(n71), .Y(n68) );
  OAI21XL U7 ( .A0(n44), .A1(n65), .B0(n64), .Y(n70) );
  NOR2X1 U8 ( .A(n52), .B(n67), .Y(n69) );
  BUFX4 U9 ( .A(n254), .Y(out[1]) );
  NOR2X2 U10 ( .A(n26), .B(n83), .Y(n84) );
  AOI2BB2X1 U11 ( .B0(n66), .B1(n44), .A0N(n45), .A1N(neg_mul[9]), .Y(n67) );
  NAND2X1 U12 ( .A(n44), .B(n8), .Y(n64) );
  AOI2BB2X1 U13 ( .B0(n74), .B1(n44), .A0N(n45), .A1N(neg_mul[10]), .Y(n75) );
  INVX8 U14 ( .A(n46), .Y(n44) );
  XNOR2X1 U15 ( .A(neg_mul[23]), .B(n40), .Y(n17) );
  NOR2X2 U16 ( .A(n25), .B(n81), .Y(n82) );
  INVXL U17 ( .A(n50), .Y(n49) );
  INVXL U18 ( .A(n50), .Y(n53) );
  NOR2BX1 U19 ( .AN(n50), .B(n75), .Y(n76) );
  NAND2X1 U20 ( .A(n44), .B(n10), .Y(n72) );
  AOI211X2 U21 ( .A0(n53), .A1(n63), .B0(n62), .C0(n39), .Y(n254) );
  XNOR2X1 U22 ( .A(n52), .B(n44), .Y(n85) );
  NOR2X2 U23 ( .A(n52), .B(n61), .Y(n62) );
  OAI21X1 U24 ( .A0(n44), .A1(n73), .B0(n72), .Y(n77) );
  INVX8 U25 ( .A(in_8bit[7]), .Y(n46) );
  NOR2X4 U26 ( .A(n79), .B(n78), .Y(n80) );
  OR2X4 U27 ( .A(n86), .B(n35), .Y(n24) );
  XNOR2X1 U28 ( .A(n52), .B(n44), .Y(n83) );
  INVX8 U29 ( .A(n50), .Y(n52) );
  INVX8 U30 ( .A(in_17bit[16]), .Y(n50) );
  INVX8 U31 ( .A(n86), .Y(n87) );
  XNOR2X4 U32 ( .A(n52), .B(n44), .Y(n86) );
  AOI22XL U33 ( .A0(N355), .A1(n249), .B0(n173), .B1(in_17bit_b[8]), .Y(n226)
         );
  AOI22XL U34 ( .A0(N356), .A1(n249), .B0(n173), .B1(in_17bit_b[9]), .Y(n229)
         );
  AOI22XL U35 ( .A0(N357), .A1(n249), .B0(n173), .B1(in_17bit_b[10]), .Y(n232)
         );
  AOI22XL U36 ( .A0(N358), .A1(n249), .B0(n173), .B1(in_17bit_b[11]), .Y(n235)
         );
  AOI22XL U37 ( .A0(N120), .A1(n246), .B0(N217), .B1(n250), .Y(n237) );
  AOI22XL U38 ( .A0(N359), .A1(n249), .B0(n173), .B1(in_17bit_b[12]), .Y(n238)
         );
  AOI22XL U39 ( .A0(N121), .A1(n246), .B0(N218), .B1(n250), .Y(n240) );
  AOI22XL U40 ( .A0(N360), .A1(n249), .B0(n173), .B1(in_17bit_b[13]), .Y(n241)
         );
  AOI22XL U41 ( .A0(N122), .A1(n246), .B0(N219), .B1(n250), .Y(n243) );
  AOI22XL U42 ( .A0(N361), .A1(n249), .B0(n173), .B1(in_17bit_b[14]), .Y(n244)
         );
  AOI22XL U43 ( .A0(N123), .A1(n246), .B0(N220), .B1(n250), .Y(n247) );
  AOI22XL U44 ( .A0(N362), .A1(n249), .B0(n173), .B1(in_17bit_b[15]), .Y(n248)
         );
  INVX1 U45 ( .A(n203), .Y(in_17bit_b[1]) );
  INVX1 U46 ( .A(n242), .Y(in_17bit_b[14]) );
  INVX1 U47 ( .A(n239), .Y(in_17bit_b[13]) );
  INVX1 U48 ( .A(n206), .Y(in_17bit_b[2]) );
  INVX1 U49 ( .A(n215), .Y(in_17bit_b[5]) );
  INVX1 U50 ( .A(n218), .Y(in_17bit_b[6]) );
  INVX1 U51 ( .A(n221), .Y(in_17bit_b[7]) );
  INVX1 U52 ( .A(n224), .Y(in_17bit_b[8]) );
  INVX1 U53 ( .A(n227), .Y(in_17bit_b[9]) );
  INVX1 U54 ( .A(n230), .Y(in_17bit_b[10]) );
  INVX1 U55 ( .A(n233), .Y(in_17bit_b[11]) );
  INVX1 U56 ( .A(n236), .Y(in_17bit_b[12]) );
  INVX1 U57 ( .A(n212), .Y(in_17bit_b[4]) );
  INVX1 U58 ( .A(n209), .Y(in_17bit_b[3]) );
  XNOR2X4 U59 ( .A(n19), .B(n3), .Y(out[7]) );
  NOR2X4 U60 ( .A(n27), .B(n85), .Y(n19) );
  AOI21X1 U61 ( .A0(n20), .A1(n21), .B0(n246), .Y(n199) );
  NOR4XL U62 ( .A(in_8bit[4]), .B(in_8bit[5]), .C(in_8bit[6]), .D(n45), .Y(n20) );
  NOR4X1 U63 ( .A(in_8bit[1]), .B(in_8bit[0]), .C(in_8bit[2]), .D(in_8bit[3]), 
        .Y(n21) );
  AND4X1 U64 ( .A(in_8bit[1]), .B(n45), .C(n194), .D(n43), .Y(n22) );
  ADDFX2 U65 ( .A(n42), .B(in_17bit_b[12]), .CI(add_1_root_r112_carry_16_), 
        .CO(add_1_root_r112_carry_17_), .S(add_1_root_r112_SUM_16_) );
  ADDFX2 U66 ( .A(add_1_root_r119_A_19_), .B(in_17bit_b[13]), .CI(
        add_1_root_r119_carry[19]), .CO(add_1_root_r119_carry[20]), .S(
        add_1_root_r119_SUM_19_) );
  ADDFX2 U67 ( .A(n42), .B(in_17bit_b[15]), .CI(add_3_root_r119_carry_17_), 
        .CO(add_3_root_r119_carry_18_), .S(add_1_root_r119_A_17_) );
  ADDFX2 U68 ( .A(n42), .B(in_17bit_b[14]), .CI(add_2_root_r115_carry_17_), 
        .CO(add_2_root_r115_carry_18_), .S(add_2_root_r115_SUM_17_) );
  ADDFX2 U69 ( .A(n42), .B(in_17bit_b[14]), .CI(add_1_root_r115_carry_20_), 
        .CO(add_1_root_r115_carry_21_), .S(add_1_root_r115_SUM_20_) );
  ADDFX2 U70 ( .A(n42), .B(in_17bit_b[15]), .CI(add_2_root_r119_carry_20_), 
        .CO(add_2_root_r119_carry_21_), .S(add_2_root_r119_SUM_20_) );
  INVX1 U71 ( .A(n56), .Y(n51) );
  ADDFX2 U72 ( .A(in_17bit_b[3]), .B(in_17bit_b[1]), .CI(
        add_2_root_r115_carry_4_), .CO(add_2_root_r115_carry_5_), .S(
        add_2_root_r115_SUM_4_) );
  ADDFX2 U73 ( .A(in_17bit_b[4]), .B(in_17bit_b[2]), .CI(
        add_2_root_r115_carry_5_), .CO(add_2_root_r115_carry_6_), .S(
        add_2_root_r115_SUM_5_) );
  ADDFX2 U74 ( .A(in_17bit_b[5]), .B(in_17bit_b[1]), .CI(
        add_1_root_r112_carry_5_), .CO(add_1_root_r112_carry_6_), .S(
        add_1_root_r112_SUM_5_) );
  ADDFX2 U75 ( .A(in_17bit_b[6]), .B(in_17bit_b[5]), .CI(
        add_3_root_r119_carry_7_), .CO(add_3_root_r119_carry_8_), .S(
        add_1_root_r119_A_7_) );
  ADDFX2 U76 ( .A(in_17bit_b[6]), .B(in_17bit_b[2]), .CI(
        add_1_root_r112_carry_6_), .CO(add_1_root_r112_carry_7_), .S(
        add_1_root_r112_SUM_6_) );
  ADDFX2 U77 ( .A(in_17bit_b[3]), .B(in_17bit_b[1]), .CI(
        add_1_root_r115_carry_7_), .CO(add_1_root_r115_carry_8_), .S(
        add_1_root_r115_SUM_7_) );
  ADDFX2 U78 ( .A(in_17bit_b[7]), .B(in_17bit_b[6]), .CI(
        add_3_root_r119_carry_8_), .CO(add_3_root_r119_carry_9_), .S(
        add_1_root_r119_A_8_) );
  ADDFX2 U79 ( .A(add_1_root_r119_A_7_), .B(in_17bit_b[1]), .CI(
        add_1_root_r119_carry[7]), .CO(add_1_root_r119_carry[8]), .S(
        add_1_root_r119_SUM_7_) );
  ADDFX2 U80 ( .A(in_17bit_b[2]), .B(in_17bit_b[1]), .CI(
        add_2_root_r119_carry_6_), .CO(add_2_root_r119_carry_7_), .S(
        add_2_root_r119_SUM_6_) );
  ADDFX2 U81 ( .A(in_17bit_b[4]), .B(in_17bit_b[2]), .CI(
        add_1_root_r115_carry_8_), .CO(add_1_root_r115_carry_9_), .S(
        add_1_root_r115_SUM_8_) );
  ADDFX2 U82 ( .A(in_17bit_b[8]), .B(in_17bit_b[7]), .CI(
        add_3_root_r119_carry_9_), .CO(add_3_root_r119_carry_10_), .S(
        add_1_root_r119_A_9_) );
  ADDFX2 U83 ( .A(add_1_root_r119_A_8_), .B(in_17bit_b[2]), .CI(
        add_1_root_r119_carry[8]), .CO(add_1_root_r119_carry[9]), .S(
        add_1_root_r119_SUM_8_) );
  ADDFX2 U84 ( .A(in_17bit_b[3]), .B(in_17bit_b[2]), .CI(
        add_2_root_r119_carry_7_), .CO(add_2_root_r119_carry_8_), .S(
        add_2_root_r119_SUM_7_) );
  ADDFX2 U85 ( .A(in_17bit_b[6]), .B(in_17bit_b[4]), .CI(
        add_2_root_r115_carry_7_), .CO(add_2_root_r115_carry_8_), .S(
        add_2_root_r115_SUM_7_) );
  ADDFX2 U86 ( .A(in_17bit_b[8]), .B(in_17bit_b[4]), .CI(
        add_1_root_r112_carry_8_), .CO(add_1_root_r112_carry_9_), .S(
        add_1_root_r112_SUM_8_) );
  ADDFX2 U87 ( .A(in_17bit_b[9]), .B(in_17bit_b[8]), .CI(
        add_3_root_r119_carry_10_), .CO(add_3_root_r119_carry_11_), .S(
        add_1_root_r119_A_10_) );
  ADDFX2 U88 ( .A(in_17bit_b[9]), .B(in_17bit_b[5]), .CI(
        add_1_root_r112_carry_9_), .CO(add_1_root_r112_carry_10_), .S(
        add_1_root_r112_SUM_9_) );
  ADDFX2 U89 ( .A(in_17bit_b[10]), .B(in_17bit_b[9]), .CI(
        add_3_root_r119_carry_11_), .CO(add_3_root_r119_carry_12_), .S(
        add_1_root_r119_A_11_) );
  ADDFX2 U90 ( .A(in_17bit_b[7]), .B(in_17bit_b[5]), .CI(
        add_2_root_r115_carry_8_), .CO(add_2_root_r115_carry_9_), .S(
        add_2_root_r115_SUM_8_) );
  ADDFX2 U91 ( .A(in_17bit_b[6]), .B(in_17bit_b[4]), .CI(
        add_1_root_r115_carry_10_), .CO(add_1_root_r115_carry_11_), .S(
        add_1_root_r115_SUM_10_) );
  ADDFX2 U92 ( .A(in_17bit_b[5]), .B(in_17bit_b[4]), .CI(
        add_2_root_r119_carry_9_), .CO(add_2_root_r119_carry_10_), .S(
        add_2_root_r119_SUM_9_) );
  ADDFX2 U93 ( .A(in_17bit_b[8]), .B(in_17bit_b[6]), .CI(
        add_2_root_r115_carry_9_), .CO(add_2_root_r115_carry_10_), .S(
        add_2_root_r115_SUM_9_) );
  ADDFX2 U94 ( .A(in_17bit_b[10]), .B(in_17bit_b[6]), .CI(
        add_1_root_r112_carry_10_), .CO(add_1_root_r112_carry_11_), .S(
        add_1_root_r112_SUM_10_) );
  ADDFX2 U95 ( .A(in_17bit_b[7]), .B(in_17bit_b[5]), .CI(
        add_1_root_r115_carry_11_), .CO(add_1_root_r115_carry_12_), .S(
        add_1_root_r115_SUM_11_) );
  ADDFX2 U96 ( .A(in_17bit_b[11]), .B(in_17bit_b[10]), .CI(
        add_3_root_r119_carry_12_), .CO(add_3_root_r119_carry_13_), .S(
        add_1_root_r119_A_12_) );
  ADDFX2 U97 ( .A(add_1_root_r119_A_11_), .B(in_17bit_b[5]), .CI(
        add_1_root_r119_carry[11]), .CO(add_1_root_r119_carry[12]), .S(
        add_1_root_r119_SUM_11_) );
  ADDFX2 U98 ( .A(in_17bit_b[6]), .B(in_17bit_b[5]), .CI(
        add_2_root_r119_carry_10_), .CO(add_2_root_r119_carry_11_), .S(
        add_2_root_r119_SUM_10_) );
  ADDFX2 U99 ( .A(in_17bit_b[9]), .B(in_17bit_b[7]), .CI(
        add_2_root_r115_carry_10_), .CO(add_2_root_r115_carry_11_), .S(
        add_2_root_r115_SUM_10_) );
  ADDFX2 U100 ( .A(in_17bit_b[11]), .B(in_17bit_b[7]), .CI(
        add_1_root_r112_carry_11_), .CO(add_1_root_r112_carry_12_), .S(
        add_1_root_r112_SUM_11_) );
  ADDFX2 U101 ( .A(in_17bit_b[8]), .B(in_17bit_b[6]), .CI(
        add_1_root_r115_carry_12_), .CO(add_1_root_r115_carry_13_), .S(
        add_1_root_r115_SUM_12_) );
  ADDFX2 U102 ( .A(in_17bit_b[12]), .B(in_17bit_b[11]), .CI(
        add_3_root_r119_carry_13_), .CO(add_3_root_r119_carry_14_), .S(
        add_1_root_r119_A_13_) );
  ADDFX2 U103 ( .A(add_1_root_r119_A_12_), .B(in_17bit_b[6]), .CI(
        add_1_root_r119_carry[12]), .CO(add_1_root_r119_carry[13]), .S(
        add_1_root_r119_SUM_12_) );
  ADDFX2 U104 ( .A(in_17bit_b[7]), .B(in_17bit_b[6]), .CI(
        add_2_root_r119_carry_11_), .CO(add_2_root_r119_carry_12_), .S(
        add_2_root_r119_SUM_11_) );
  ADDFX2 U105 ( .A(in_17bit_b[10]), .B(in_17bit_b[8]), .CI(
        add_2_root_r115_carry_11_), .CO(add_2_root_r115_carry_12_), .S(
        add_2_root_r115_SUM_11_) );
  ADDFX2 U106 ( .A(in_17bit_b[12]), .B(in_17bit_b[8]), .CI(
        add_1_root_r112_carry_12_), .CO(add_1_root_r112_carry_13_), .S(
        add_1_root_r112_SUM_12_) );
  ADDFX2 U107 ( .A(in_17bit_b[9]), .B(in_17bit_b[7]), .CI(
        add_1_root_r115_carry_13_), .CO(add_1_root_r115_carry_14_), .S(
        add_1_root_r115_SUM_13_) );
  ADDFX2 U108 ( .A(in_17bit_b[13]), .B(in_17bit_b[12]), .CI(
        add_3_root_r119_carry_14_), .CO(add_3_root_r119_carry_15_), .S(
        add_1_root_r119_A_14_) );
  ADDFX2 U109 ( .A(add_1_root_r119_A_13_), .B(in_17bit_b[7]), .CI(
        add_1_root_r119_carry[13]), .CO(add_1_root_r119_carry[14]), .S(
        add_1_root_r119_SUM_13_) );
  ADDFX2 U110 ( .A(in_17bit_b[8]), .B(in_17bit_b[7]), .CI(
        add_2_root_r119_carry_12_), .CO(add_2_root_r119_carry_13_), .S(
        add_2_root_r119_SUM_12_) );
  ADDFX2 U111 ( .A(in_17bit_b[11]), .B(in_17bit_b[9]), .CI(
        add_2_root_r115_carry_12_), .CO(add_2_root_r115_carry_13_), .S(
        add_2_root_r115_SUM_12_) );
  ADDFX2 U112 ( .A(in_17bit_b[13]), .B(in_17bit_b[9]), .CI(
        add_1_root_r112_carry_13_), .CO(add_1_root_r112_carry_14_), .S(
        add_1_root_r112_SUM_13_) );
  ADDFX2 U113 ( .A(in_17bit_b[10]), .B(in_17bit_b[8]), .CI(
        add_1_root_r115_carry_14_), .CO(add_1_root_r115_carry_15_), .S(
        add_1_root_r115_SUM_14_) );
  ADDFX2 U114 ( .A(in_17bit_b[14]), .B(in_17bit_b[13]), .CI(
        add_3_root_r119_carry_15_), .CO(add_3_root_r119_carry_16_), .S(
        add_1_root_r119_A_15_) );
  ADDFX2 U115 ( .A(add_1_root_r119_A_14_), .B(in_17bit_b[8]), .CI(
        add_1_root_r119_carry[14]), .CO(add_1_root_r119_carry[15]), .S(
        add_1_root_r119_SUM_14_) );
  ADDFX2 U116 ( .A(in_17bit_b[9]), .B(in_17bit_b[8]), .CI(
        add_2_root_r119_carry_13_), .CO(add_2_root_r119_carry_14_), .S(
        add_2_root_r119_SUM_13_) );
  ADDFX2 U117 ( .A(in_17bit_b[12]), .B(in_17bit_b[10]), .CI(
        add_2_root_r115_carry_13_), .CO(add_2_root_r115_carry_14_), .S(
        add_2_root_r115_SUM_13_) );
  ADDFX2 U118 ( .A(in_17bit_b[14]), .B(in_17bit_b[10]), .CI(
        add_1_root_r112_carry_14_), .CO(add_1_root_r112_carry_15_), .S(
        add_1_root_r112_SUM_14_) );
  ADDFX2 U119 ( .A(in_17bit_b[11]), .B(in_17bit_b[9]), .CI(
        add_1_root_r115_carry_15_), .CO(add_1_root_r115_carry_16_), .S(
        add_1_root_r115_SUM_15_) );
  ADDFX2 U120 ( .A(add_1_root_r119_A_15_), .B(in_17bit_b[9]), .CI(
        add_1_root_r119_carry[15]), .CO(add_1_root_r119_carry[16]), .S(
        add_1_root_r119_SUM_15_) );
  ADDFX2 U121 ( .A(in_17bit_b[3]), .B(in_17bit_b[2]), .CI(
        add_3_root_r119_carry_4_), .CO(add_3_root_r119_carry_5_), .S(
        add_1_root_r119_A_4_) );
  ADDFX2 U122 ( .A(in_17bit_b[2]), .B(in_17bit_b[1]), .CI(
        add_3_root_r119_carry_3_), .CO(add_3_root_r119_carry_4_), .S(
        add_1_root_r119_A_3_) );
  ADDFX2 U123 ( .A(in_17bit_b[10]), .B(in_17bit_b[9]), .CI(
        add_2_root_r119_carry_14_), .CO(add_2_root_r119_carry_15_), .S(
        add_2_root_r119_SUM_14_) );
  ADDFX2 U124 ( .A(in_17bit_b[13]), .B(in_17bit_b[11]), .CI(
        add_2_root_r115_carry_14_), .CO(add_2_root_r115_carry_15_), .S(
        add_2_root_r115_SUM_14_) );
  ADDFX2 U125 ( .A(in_17bit_b[15]), .B(in_17bit_b[11]), .CI(
        add_1_root_r112_carry_15_), .CO(add_1_root_r112_carry_16_), .S(
        add_1_root_r112_SUM_15_) );
  ADDFX2 U126 ( .A(in_17bit_b[12]), .B(in_17bit_b[10]), .CI(
        add_1_root_r115_carry_16_), .CO(add_1_root_r115_carry_17_), .S(
        add_1_root_r115_SUM_16_) );
  ADDFX2 U127 ( .A(add_1_root_r119_A_16_), .B(in_17bit_b[10]), .CI(
        add_1_root_r119_carry[16]), .CO(add_1_root_r119_carry[17]), .S(
        add_1_root_r119_SUM_16_) );
  ADDFX2 U128 ( .A(in_17bit_b[11]), .B(in_17bit_b[10]), .CI(
        add_2_root_r119_carry_15_), .CO(add_2_root_r119_carry_16_), .S(
        add_2_root_r119_SUM_15_) );
  ADDFX2 U129 ( .A(in_17bit_b[14]), .B(in_17bit_b[12]), .CI(
        add_2_root_r115_carry_15_), .CO(add_2_root_r115_carry_16_), .S(
        add_2_root_r115_SUM_15_) );
  ADDFX2 U130 ( .A(in_17bit_b[13]), .B(in_17bit_b[11]), .CI(
        add_1_root_r115_carry_17_), .CO(add_1_root_r115_carry_18_), .S(
        add_1_root_r115_SUM_17_) );
  ADDFX2 U131 ( .A(add_1_root_r119_A_17_), .B(in_17bit_b[11]), .CI(
        add_1_root_r119_carry[17]), .CO(add_1_root_r119_carry[18]), .S(
        add_1_root_r119_SUM_17_) );
  ADDFX2 U132 ( .A(in_17bit_b[12]), .B(in_17bit_b[11]), .CI(
        add_2_root_r119_carry_16_), .CO(add_2_root_r119_carry_17_), .S(
        add_2_root_r119_SUM_16_) );
  ADDFX2 U133 ( .A(in_17bit_b[14]), .B(in_17bit_b[12]), .CI(
        add_1_root_r115_carry_18_), .CO(add_1_root_r115_carry_19_), .S(
        add_1_root_r115_SUM_18_) );
  ADDFX2 U134 ( .A(add_1_root_r119_A_18_), .B(in_17bit_b[12]), .CI(
        add_1_root_r119_carry[18]), .CO(add_1_root_r119_carry[19]), .S(
        add_1_root_r119_SUM_18_) );
  ADDFX2 U135 ( .A(in_17bit_b[13]), .B(in_17bit_b[12]), .CI(
        add_2_root_r119_carry_17_), .CO(add_2_root_r119_carry_18_), .S(
        add_2_root_r119_SUM_17_) );
  ADDFX2 U136 ( .A(in_17bit_b[15]), .B(in_17bit_b[13]), .CI(
        add_2_root_r115_carry_16_), .CO(add_2_root_r115_carry_17_), .S(
        add_2_root_r115_SUM_16_) );
  ADDFX2 U137 ( .A(in_17bit_b[15]), .B(in_17bit_b[13]), .CI(
        add_1_root_r115_carry_19_), .CO(add_1_root_r115_carry_20_), .S(
        add_1_root_r115_SUM_19_) );
  ADDFX2 U138 ( .A(in_17bit_b[5]), .B(in_17bit_b[3]), .CI(
        add_2_root_r115_carry_6_), .CO(add_2_root_r115_carry_7_), .S(
        add_2_root_r115_SUM_6_) );
  ADDFX2 U139 ( .A(in_17bit_b[5]), .B(in_17bit_b[3]), .CI(
        add_1_root_r115_carry_9_), .CO(add_1_root_r115_carry_10_), .S(
        add_1_root_r115_SUM_9_) );
  ADDFX2 U140 ( .A(in_17bit_b[4]), .B(in_17bit_b[3]), .CI(
        add_2_root_r119_carry_8_), .CO(add_2_root_r119_carry_9_), .S(
        add_2_root_r119_SUM_8_) );
  ADDFX2 U141 ( .A(in_17bit_b[15]), .B(in_17bit_b[14]), .CI(
        add_3_root_r119_carry_16_), .CO(add_3_root_r119_carry_17_), .S(
        add_1_root_r119_A_16_) );
  ADDFX2 U142 ( .A(in_17bit_b[7]), .B(in_17bit_b[3]), .CI(
        add_1_root_r112_carry_7_), .CO(add_1_root_r112_carry_8_), .S(
        add_1_root_r112_SUM_7_) );
  ADDFX2 U143 ( .A(add_1_root_r119_A_9_), .B(in_17bit_b[3]), .CI(
        add_1_root_r119_carry[9]), .CO(add_1_root_r119_carry[10]), .S(
        add_1_root_r119_SUM_9_) );
  ADDFX2 U144 ( .A(add_1_root_r119_A_10_), .B(in_17bit_b[4]), .CI(
        add_1_root_r119_carry[10]), .CO(add_1_root_r119_carry[11]), .S(
        add_1_root_r119_SUM_10_) );
  ADDFX2 U145 ( .A(in_17bit_b[4]), .B(in_17bit_b[3]), .CI(
        add_3_root_r119_carry_5_), .CO(add_3_root_r119_carry_6_), .S(
        add_1_root_r119_A_5_) );
  ADDFX2 U146 ( .A(in_17bit_b[14]), .B(in_17bit_b[13]), .CI(
        add_2_root_r119_carry_18_), .CO(add_2_root_r119_carry_19_), .S(
        add_2_root_r119_SUM_18_) );
  ADDFX2 U147 ( .A(in_17bit_b[5]), .B(in_17bit_b[4]), .CI(
        add_3_root_r119_carry_6_), .CO(add_3_root_r119_carry_7_), .S(
        add_1_root_r119_A_6_) );
  ADDFX2 U148 ( .A(in_17bit_b[15]), .B(in_17bit_b[14]), .CI(
        add_2_root_r119_carry_19_), .CO(add_2_root_r119_carry_20_), .S(
        add_2_root_r119_SUM_19_) );
  BUFX3 U149 ( .A(in_17bit_b[16]), .Y(n42) );
  INVX1 U150 ( .A(n253), .Y(in_17bit_b[16]) );
  INVX1 U151 ( .A(n49), .Y(n54) );
  INVX1 U152 ( .A(n49), .Y(n55) );
  INVX1 U153 ( .A(n49), .Y(n56) );
  CLKINVX3 U154 ( .A(n200), .Y(in_17bit_b[0]) );
  INVX1 U155 ( .A(n173), .Y(n252) );
  NAND2XL U156 ( .A(N29), .B(n52), .Y(n253) );
  OAI21XL U157 ( .A0(n252), .A1(n253), .B0(n251), .Y(N463) );
  AOI22XL U158 ( .A0(N221), .A1(n250), .B0(N363), .B1(n249), .Y(n251) );
  CLKINVX3 U159 ( .A(n245), .Y(in_17bit_b[15]) );
  NAND2X1 U160 ( .A(n34), .B(in_8bit[1]), .Y(n88) );
  INVX1 U161 ( .A(in_8bit[0]), .Y(n43) );
  INVX1 U162 ( .A(in_8bit[2]), .Y(n47) );
  INVX1 U163 ( .A(in_8bit[5]), .Y(n48) );
  OAI21XL U164 ( .A0(n44), .A1(n59), .B0(n58), .Y(n63) );
  MXI2XL U165 ( .A(n1), .B(n17), .S0(n87), .Y(out[16]) );
  XOR2X4 U166 ( .A(n23), .B(n2), .Y(out[8]) );
  OR2X4 U167 ( .A(n86), .B(n29), .Y(n23) );
  XOR2X4 U168 ( .A(n24), .B(n7), .Y(out[9]) );
  NOR3X1 U169 ( .A(n47), .B(n174), .C(n43), .Y(n198) );
  AOI22XL U170 ( .A0(in_17bit[0]), .A1(n52), .B0(in_17bit[0]), .B1(n55), .Y(
        n200) );
  AOI22X1 U171 ( .A0(N27), .A1(n51), .B0(in_17bit[14]), .B1(n54), .Y(n242) );
  AOI22X1 U172 ( .A0(N28), .A1(n51), .B0(in_17bit[15]), .B1(n56), .Y(n245) );
  AOI22X1 U173 ( .A0(N26), .A1(n51), .B0(in_17bit[13]), .B1(n54), .Y(n239) );
  AOI22XL U174 ( .A0(N14), .A1(n52), .B0(in_17bit[1]), .B1(n54), .Y(n203) );
  AOI22XL U175 ( .A0(N15), .A1(n52), .B0(in_17bit[2]), .B1(n56), .Y(n206) );
  AOI22X1 U176 ( .A0(N16), .A1(n51), .B0(in_17bit[3]), .B1(n55), .Y(n209) );
  AOI22X1 U177 ( .A0(N17), .A1(n51), .B0(in_17bit[4]), .B1(n56), .Y(n212) );
  AOI22X1 U178 ( .A0(N18), .A1(n51), .B0(in_17bit[5]), .B1(n56), .Y(n215) );
  AOI22X1 U179 ( .A0(N19), .A1(n51), .B0(in_17bit[6]), .B1(n55), .Y(n218) );
  AOI22X1 U180 ( .A0(N20), .A1(n51), .B0(in_17bit[7]), .B1(n56), .Y(n221) );
  AOI22X1 U181 ( .A0(N21), .A1(n51), .B0(in_17bit[8]), .B1(n55), .Y(n224) );
  AOI22X1 U182 ( .A0(N23), .A1(n51), .B0(in_17bit[10]), .B1(n54), .Y(n230) );
  AOI22X1 U183 ( .A0(N24), .A1(n51), .B0(in_17bit[11]), .B1(n55), .Y(n233) );
  AOI22X1 U184 ( .A0(N25), .A1(n51), .B0(in_17bit[12]), .B1(n55), .Y(n236) );
  AOI22X1 U185 ( .A0(N22), .A1(n51), .B0(in_17bit[9]), .B1(n54), .Y(n227) );
  INVX1 U186 ( .A(n57), .Y(n79) );
  NAND2BX1 U187 ( .AN(n71), .B(n10), .Y(n57) );
  NAND2X1 U188 ( .A(n39), .B(n8), .Y(n71) );
  AND2X2 U189 ( .A(n79), .B(n4), .Y(n25) );
  AND2X2 U190 ( .A(n25), .B(n5), .Y(n26) );
  AND2X2 U191 ( .A(n26), .B(n6), .Y(n27) );
  NOR2X1 U192 ( .A(in_8bit[0]), .B(n94), .Y(n28) );
  AND2X2 U193 ( .A(n27), .B(n3), .Y(n29) );
  AOI21X1 U194 ( .A0(n93), .A1(n22), .B0(n31), .Y(n30) );
  INVX1 U195 ( .A(n30), .Y(n249) );
  AND2X2 U196 ( .A(n28), .B(n36), .Y(n31) );
  AOI21X1 U197 ( .A0(n36), .A1(n22), .B0(n33), .Y(n32) );
  INVX1 U198 ( .A(n32), .Y(n250) );
  AND2X2 U199 ( .A(n28), .B(n93), .Y(n33) );
  OAI2BB1X1 U200 ( .A0N(n197), .A1N(n34), .B0(n95), .Y(n173) );
  NAND3BX1 U201 ( .AN(n94), .B(n198), .C(in_8bit[5]), .Y(n95) );
  AND3X1 U202 ( .A(n45), .B(n89), .C(n48), .Y(n34) );
  NOR2XL U203 ( .A(n44), .B(n89), .Y(n90) );
  AND2X2 U204 ( .A(n29), .B(n2), .Y(n35) );
  INVX1 U205 ( .A(in_17bit[8]), .Y(n161) );
  INVX1 U206 ( .A(in_17bit[9]), .Y(n162) );
  INVX1 U207 ( .A(in_17bit[10]), .Y(n163) );
  INVX1 U208 ( .A(in_17bit[11]), .Y(n164) );
  INVX1 U209 ( .A(in_17bit[12]), .Y(n167) );
  INVX1 U210 ( .A(in_17bit[13]), .Y(n168) );
  INVX1 U211 ( .A(in_17bit[14]), .Y(n170) );
  INVX1 U212 ( .A(in_17bit[15]), .Y(n171) );
  INVX1 U213 ( .A(in_17bit[1]), .Y(n97) );
  INVX1 U214 ( .A(in_17bit[2]), .Y(n98) );
  INVX1 U215 ( .A(in_17bit[3]), .Y(n99) );
  INVX1 U216 ( .A(in_17bit[4]), .Y(n100) );
  INVX1 U217 ( .A(in_17bit[5]), .Y(n101) );
  INVX1 U218 ( .A(in_17bit[6]), .Y(n158) );
  INVX1 U219 ( .A(in_17bit[7]), .Y(n160) );
  INVX1 U220 ( .A(in_17bit[0]), .Y(n96) );
  AND3X2 U221 ( .A(in_8bit[2]), .B(n174), .C(in_8bit[5]), .Y(n36) );
  NAND2X1 U222 ( .A(n202), .B(n201), .Y(N447) );
  AOI22X1 U223 ( .A0(N108), .A1(n246), .B0(N205), .B1(n250), .Y(n201) );
  AOI22X1 U224 ( .A0(N347), .A1(n249), .B0(n173), .B1(in_17bit_b[0]), .Y(n202)
         );
  NAND2X1 U225 ( .A(n205), .B(n204), .Y(N448) );
  AOI22X1 U226 ( .A0(N109), .A1(n246), .B0(N206), .B1(n250), .Y(n204) );
  AOI22X1 U227 ( .A0(N348), .A1(n249), .B0(n173), .B1(n172), .Y(n205) );
  INVX1 U228 ( .A(n203), .Y(n172) );
  NAND2X1 U229 ( .A(n208), .B(n207), .Y(N449) );
  AOI22X1 U230 ( .A0(N110), .A1(n246), .B0(N207), .B1(n250), .Y(n207) );
  AOI22X1 U231 ( .A0(N349), .A1(n249), .B0(n173), .B1(in_17bit_b[2]), .Y(n208)
         );
  NAND2X1 U232 ( .A(n211), .B(n210), .Y(N450) );
  AOI22X1 U233 ( .A0(N111), .A1(n246), .B0(N208), .B1(n250), .Y(n210) );
  AOI22X1 U234 ( .A0(N350), .A1(n249), .B0(n173), .B1(in_17bit_b[3]), .Y(n211)
         );
  NAND2X1 U235 ( .A(n214), .B(n213), .Y(N451) );
  AOI22X1 U236 ( .A0(N112), .A1(n246), .B0(N209), .B1(n250), .Y(n213) );
  AOI22X1 U237 ( .A0(N351), .A1(n249), .B0(n173), .B1(in_17bit_b[4]), .Y(n214)
         );
  NAND2X1 U238 ( .A(n217), .B(n216), .Y(N452) );
  AOI22X1 U239 ( .A0(N113), .A1(n246), .B0(N210), .B1(n250), .Y(n216) );
  AOI22X1 U240 ( .A0(N352), .A1(n249), .B0(n173), .B1(in_17bit_b[5]), .Y(n217)
         );
  NAND2X1 U241 ( .A(n220), .B(n219), .Y(N453) );
  AOI22X1 U242 ( .A0(N114), .A1(n246), .B0(N211), .B1(n250), .Y(n219) );
  AOI22X1 U243 ( .A0(N353), .A1(n249), .B0(n173), .B1(in_17bit_b[6]), .Y(n220)
         );
  NAND2X1 U244 ( .A(n223), .B(n222), .Y(N454) );
  AOI22X1 U245 ( .A0(N115), .A1(n246), .B0(N212), .B1(n250), .Y(n222) );
  AOI22X1 U246 ( .A0(N354), .A1(n249), .B0(n173), .B1(in_17bit_b[7]), .Y(n223)
         );
  NAND2X1 U247 ( .A(n226), .B(n225), .Y(N455) );
  AOI22X1 U248 ( .A0(N116), .A1(n246), .B0(N213), .B1(n250), .Y(n225) );
  NAND2X1 U249 ( .A(n229), .B(n228), .Y(N456) );
  AOI22X1 U250 ( .A0(N117), .A1(n246), .B0(N214), .B1(n250), .Y(n228) );
  NAND2X1 U251 ( .A(n232), .B(n231), .Y(N457) );
  AOI22X1 U252 ( .A0(N118), .A1(n246), .B0(N215), .B1(n250), .Y(n231) );
  NAND2X1 U253 ( .A(n235), .B(n234), .Y(N458) );
  AOI22X1 U254 ( .A0(N119), .A1(n246), .B0(N216), .B1(n250), .Y(n234) );
  NAND2X1 U255 ( .A(n238), .B(n237), .Y(N459) );
  NAND2X1 U256 ( .A(n241), .B(n240), .Y(N460) );
  NAND2X1 U257 ( .A(n244), .B(n243), .Y(N461) );
  NAND2X1 U258 ( .A(n248), .B(n247), .Y(N462) );
  XNOR2X1 U259 ( .A(n15), .B(sub_add_75_b0_carry[11]), .Y(n37) );
  XNOR2X1 U260 ( .A(n14), .B(sub_add_75_b0_carry[10]), .Y(n38) );
  INVX1 U261 ( .A(n73), .Y(n74) );
  INVX1 U262 ( .A(n65), .Y(n66) );
  INVX1 U263 ( .A(n59), .Y(n60) );
  NAND2X2 U264 ( .A(n44), .B(n16), .Y(n58) );
  MX2X2 U265 ( .A(neg_mul[19]), .B(N477), .S0(n87), .Y(out[12]) );
  MX2X2 U266 ( .A(neg_mul[20]), .B(N478), .S0(n87), .Y(out[13]) );
  MX2X1 U267 ( .A(neg_mul[21]), .B(N479), .S0(n87), .Y(out[14]) );
  MX2X1 U268 ( .A(neg_mul[22]), .B(N480), .S0(n87), .Y(out[15]) );
  NAND4BBX1 U269 ( .AN(n249), .BN(n250), .C(n199), .D(n252), .Y(N446) );
  NOR4BX1 U270 ( .AN(n196), .B(n43), .C(in_8bit[1]), .D(in_8bit[2]), .Y(n197)
         );
  NOR2X1 U271 ( .A(in_8bit[6]), .B(in_8bit[3]), .Y(n196) );
  NOR2X1 U272 ( .A(out[0]), .B(neg_mul[8]), .Y(n39) );
  NAND4BXL U273 ( .AN(n45), .B(in_8bit[6]), .C(in_8bit[1]), .D(in_8bit[4]), 
        .Y(n94) );
  NAND2BX1 U274 ( .AN(n39), .B(neg_mul[9]), .Y(n65) );
  NAND2X1 U275 ( .A(out[0]), .B(neg_mul[8]), .Y(n59) );
  NAND2X1 U276 ( .A(neg_mul[10]), .B(n71), .Y(n73) );
  NAND2X1 U277 ( .A(n92), .B(n91), .Y(n246) );
  NAND3BX1 U278 ( .AN(n88), .B(n198), .C(in_8bit[6]), .Y(n92) );
  NAND3X1 U279 ( .A(n197), .B(in_8bit[5]), .C(n90), .Y(n91) );
  INVX1 U280 ( .A(n195), .Y(n93) );
  NAND3BX1 U281 ( .AN(in_8bit[5]), .B(n47), .C(in_8bit[3]), .Y(n195) );
  NOR2X1 U282 ( .A(in_8bit[6]), .B(in_8bit[4]), .Y(n194) );
  NAND2X1 U283 ( .A(sub_add_75_b0_carry[15]), .B(n9), .Y(n40) );
  INVX1 U284 ( .A(in_8bit[4]), .Y(n89) );
  INVX1 U285 ( .A(in_8bit[3]), .Y(n174) );
  AOI211X4 U286 ( .A0(n52), .A1(n77), .B0(n76), .C0(n79), .Y(out[3]) );
  AOI211X4 U287 ( .A0(n52), .A1(n70), .B0(n69), .C0(n68), .Y(out[2]) );
  XNOR2X4 U288 ( .A(n80), .B(n4), .Y(out[4]) );
  XNOR2X4 U289 ( .A(n82), .B(n5), .Y(out[5]) );
  XNOR2X4 U290 ( .A(n84), .B(n6), .Y(out[6]) );
  MXI2X4 U291 ( .A(n14), .B(n38), .S0(n87), .Y(out[10]) );
  MXI2X4 U292 ( .A(n15), .B(n37), .S0(n87), .Y(out[11]) );
  AND2X1 U293 ( .A(add_1_root_r112_carry_20_), .B(n42), .Y(
        add_1_root_r112_SUM_21_) );
  XOR2X1 U294 ( .A(n42), .B(add_1_root_r112_carry_20_), .Y(
        add_1_root_r112_SUM_20_) );
  AND2X1 U295 ( .A(add_1_root_r112_carry_19_), .B(in_17bit_b[15]), .Y(
        add_1_root_r112_carry_20_) );
  XOR2X1 U296 ( .A(in_17bit_b[15]), .B(add_1_root_r112_carry_19_), .Y(
        add_1_root_r112_SUM_19_) );
  AND2X1 U297 ( .A(add_1_root_r112_carry_18_), .B(in_17bit_b[14]), .Y(
        add_1_root_r112_carry_19_) );
  XOR2X1 U298 ( .A(in_17bit_b[14]), .B(add_1_root_r112_carry_18_), .Y(
        add_1_root_r112_SUM_18_) );
  AND2X1 U299 ( .A(add_1_root_r112_carry_17_), .B(in_17bit_b[13]), .Y(
        add_1_root_r112_carry_18_) );
  XOR2X1 U300 ( .A(in_17bit_b[13]), .B(add_1_root_r112_carry_17_), .Y(
        add_1_root_r112_SUM_17_) );
  AND2X1 U301 ( .A(add_2_root_r119_carry_21_), .B(n42), .Y(
        add_2_root_r119_SUM_22_) );
  XOR2X1 U302 ( .A(n42), .B(add_2_root_r119_carry_21_), .Y(
        add_2_root_r119_SUM_21_) );
  AND2X1 U303 ( .A(in_17bit_b[1]), .B(in_17bit_b[0]), .Y(
        add_2_root_r119_carry_6_) );
  XOR2X1 U304 ( .A(in_17bit_b[0]), .B(in_17bit_b[1]), .Y(
        add_2_root_r119_SUM_5_) );
  AND2X1 U305 ( .A(add_1_root_r119_carry[22]), .B(n42), .Y(
        add_1_root_r119_SUM_23_) );
  XOR2X1 U306 ( .A(n42), .B(add_1_root_r119_carry[22]), .Y(
        add_1_root_r119_SUM_22_) );
  AND2X1 U307 ( .A(add_1_root_r119_carry[21]), .B(in_17bit_b[15]), .Y(
        add_1_root_r119_carry[22]) );
  XOR2X1 U308 ( .A(in_17bit_b[15]), .B(add_1_root_r119_carry[21]), .Y(
        add_1_root_r119_SUM_21_) );
  AND2X1 U309 ( .A(add_1_root_r119_carry[20]), .B(in_17bit_b[14]), .Y(
        add_1_root_r119_carry[21]) );
  XOR2X1 U310 ( .A(in_17bit_b[14]), .B(add_1_root_r119_carry[20]), .Y(
        add_1_root_r119_SUM_20_) );
  AND2X1 U311 ( .A(add_1_root_r119_A_6_), .B(in_17bit_b[0]), .Y(
        add_1_root_r119_carry[7]) );
  XOR2X1 U312 ( .A(in_17bit_b[0]), .B(add_1_root_r119_A_6_), .Y(
        add_1_root_r119_SUM_6_) );
  AND2X1 U313 ( .A(add_3_root_r119_carry_18_), .B(n42), .Y(
        add_1_root_r119_A_19_) );
  XOR2X1 U314 ( .A(n42), .B(add_3_root_r119_carry_18_), .Y(
        add_1_root_r119_A_18_) );
  AND2X1 U315 ( .A(in_17bit_b[1]), .B(in_17bit_b[0]), .Y(
        add_3_root_r119_carry_3_) );
  XOR2X1 U316 ( .A(in_17bit_b[0]), .B(in_17bit_b[1]), .Y(add_1_root_r119_A_2_)
         );
  AND2X1 U317 ( .A(add_2_root_r115_carry_19_), .B(n42), .Y(
        add_2_root_r115_SUM_20_) );
  XOR2X1 U318 ( .A(n42), .B(add_2_root_r115_carry_19_), .Y(
        add_2_root_r115_SUM_19_) );
  AND2X1 U319 ( .A(add_2_root_r115_carry_18_), .B(in_17bit_b[15]), .Y(
        add_2_root_r115_carry_19_) );
  XOR2X1 U320 ( .A(in_17bit_b[15]), .B(add_2_root_r115_carry_18_), .Y(
        add_2_root_r115_SUM_18_) );
  AND2X1 U321 ( .A(in_17bit_b[2]), .B(in_17bit_b[0]), .Y(
        add_2_root_r115_carry_4_) );
  XOR2X1 U322 ( .A(in_17bit_b[0]), .B(in_17bit_b[2]), .Y(
        add_2_root_r115_SUM_3_) );
  AND2X1 U323 ( .A(add_1_root_r115_carry_22_), .B(n42), .Y(
        add_1_root_r115_SUM_23_) );
  XOR2X1 U324 ( .A(n42), .B(add_1_root_r115_carry_22_), .Y(
        add_1_root_r115_SUM_22_) );
  AND2X1 U325 ( .A(add_1_root_r115_carry_21_), .B(in_17bit_b[15]), .Y(
        add_1_root_r115_carry_22_) );
  XOR2X1 U326 ( .A(in_17bit_b[15]), .B(add_1_root_r115_carry_21_), .Y(
        add_1_root_r115_SUM_21_) );
  AND2X1 U327 ( .A(in_17bit_b[2]), .B(in_17bit_b[0]), .Y(
        add_1_root_r115_carry_7_) );
  XOR2X1 U328 ( .A(in_17bit_b[0]), .B(in_17bit_b[2]), .Y(
        add_1_root_r115_SUM_6_) );
  XOR2X1 U329 ( .A(n54), .B(sub_add_54_b0_carry[16]), .Y(N29) );
  AND2X1 U330 ( .A(sub_add_54_b0_carry[15]), .B(n171), .Y(
        sub_add_54_b0_carry[16]) );
  XOR2X1 U331 ( .A(n171), .B(sub_add_54_b0_carry[15]), .Y(N28) );
  AND2X1 U332 ( .A(sub_add_54_b0_carry[14]), .B(n170), .Y(
        sub_add_54_b0_carry[15]) );
  XOR2X1 U333 ( .A(n170), .B(sub_add_54_b0_carry[14]), .Y(N27) );
  AND2X1 U334 ( .A(sub_add_54_b0_carry[13]), .B(n168), .Y(
        sub_add_54_b0_carry[14]) );
  XOR2X1 U335 ( .A(n168), .B(sub_add_54_b0_carry[13]), .Y(N26) );
  AND2X1 U336 ( .A(sub_add_54_b0_carry[12]), .B(n167), .Y(
        sub_add_54_b0_carry[13]) );
  XOR2X1 U337 ( .A(n167), .B(sub_add_54_b0_carry[12]), .Y(N25) );
  AND2X1 U338 ( .A(sub_add_54_b0_carry[11]), .B(n164), .Y(
        sub_add_54_b0_carry[12]) );
  XOR2X1 U339 ( .A(n164), .B(sub_add_54_b0_carry[11]), .Y(N24) );
  AND2X1 U340 ( .A(sub_add_54_b0_carry[10]), .B(n163), .Y(
        sub_add_54_b0_carry[11]) );
  XOR2X1 U341 ( .A(n163), .B(sub_add_54_b0_carry[10]), .Y(N23) );
  AND2X1 U342 ( .A(sub_add_54_b0_carry[9]), .B(n162), .Y(
        sub_add_54_b0_carry[10]) );
  XOR2X1 U343 ( .A(n162), .B(sub_add_54_b0_carry[9]), .Y(N22) );
  AND2X1 U344 ( .A(sub_add_54_b0_carry[8]), .B(n161), .Y(
        sub_add_54_b0_carry[9]) );
  XOR2X1 U345 ( .A(n161), .B(sub_add_54_b0_carry[8]), .Y(N21) );
  AND2X1 U346 ( .A(sub_add_54_b0_carry[7]), .B(n160), .Y(
        sub_add_54_b0_carry[8]) );
  XOR2X1 U347 ( .A(n160), .B(sub_add_54_b0_carry[7]), .Y(N20) );
  AND2X1 U348 ( .A(sub_add_54_b0_carry[6]), .B(n158), .Y(
        sub_add_54_b0_carry[7]) );
  XOR2X1 U349 ( .A(n158), .B(sub_add_54_b0_carry[6]), .Y(N19) );
  AND2X1 U350 ( .A(sub_add_54_b0_carry[5]), .B(n101), .Y(
        sub_add_54_b0_carry[6]) );
  XOR2X1 U351 ( .A(n101), .B(sub_add_54_b0_carry[5]), .Y(N18) );
  AND2X1 U352 ( .A(sub_add_54_b0_carry[4]), .B(n100), .Y(
        sub_add_54_b0_carry[5]) );
  XOR2X1 U353 ( .A(n100), .B(sub_add_54_b0_carry[4]), .Y(N17) );
  AND2X1 U354 ( .A(sub_add_54_b0_carry[3]), .B(n99), .Y(sub_add_54_b0_carry[4]) );
  XOR2X1 U355 ( .A(n99), .B(sub_add_54_b0_carry[3]), .Y(N16) );
  AND2X1 U356 ( .A(sub_add_54_b0_carry[2]), .B(n98), .Y(sub_add_54_b0_carry[3]) );
  XOR2X1 U357 ( .A(n98), .B(sub_add_54_b0_carry[2]), .Y(N15) );
  AND2X1 U358 ( .A(n96), .B(n97), .Y(sub_add_54_b0_carry[2]) );
  XOR2X1 U359 ( .A(n97), .B(n96), .Y(N14) );
  XOR2X1 U360 ( .A(n9), .B(sub_add_75_b0_carry[15]), .Y(N480) );
  AND2X1 U361 ( .A(sub_add_75_b0_carry[14]), .B(n13), .Y(
        sub_add_75_b0_carry[15]) );
  XOR2X1 U362 ( .A(n13), .B(sub_add_75_b0_carry[14]), .Y(N479) );
  AND2X1 U363 ( .A(sub_add_75_b0_carry[13]), .B(n11), .Y(
        sub_add_75_b0_carry[14]) );
  XOR2X1 U364 ( .A(n11), .B(sub_add_75_b0_carry[13]), .Y(N478) );
  AND2X1 U365 ( .A(sub_add_75_b0_carry[12]), .B(n12), .Y(
        sub_add_75_b0_carry[13]) );
  XOR2X1 U366 ( .A(n12), .B(sub_add_75_b0_carry[12]), .Y(N477) );
  AND2X1 U367 ( .A(sub_add_75_b0_carry[11]), .B(n15), .Y(
        sub_add_75_b0_carry[12]) );
  AND2X1 U368 ( .A(sub_add_75_b0_carry[10]), .B(n14), .Y(
        sub_add_75_b0_carry[11]) );
  AND2X1 U369 ( .A(n35), .B(n7), .Y(sub_add_75_b0_carry[10]) );
  AND2X1 U370 ( .A(in_17bit_b[0]), .B(in_17bit_b[4]), .Y(
        add_1_root_r112_carry_5_) );
endmodule


module multi16_5_DW01_add_0 ( A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, 
        A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, 
        A_4_, B_23_, B_22_, B_21_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, 
        B_14_, B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, 
        SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, 
        SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, 
        SUM_7_ );
  input A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_,
         A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, B_23_, B_22_,
         B_21_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_,
         B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_;
  output SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_,
         SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_,
         SUM_8_, SUM_7_;
  wire   n1, n2, n3, n4;
  wire   [23:7] carry;

  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry[7]), .CO(carry[8]), .S(SUM_7_)
         );
  ADDFX2 U1_21 ( .A(A_21_), .B(B_21_), .CI(carry[21]), .CO(carry[22]), .S(
        SUM_21_) );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry[20]), .CO(carry[21]), .S(
        SUM_20_) );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry[19]), .CO(carry[20]), .S(
        SUM_19_) );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry[18]), .CO(carry[19]), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry[17]), .CO(carry[18]), .S(
        SUM_17_) );
  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry[16]), .CO(carry[17]), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry[15]), .CO(carry[16]), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry[14]), .CO(carry[15]), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry[13]), .CO(carry[14]), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry[12]), .CO(carry[13]), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry[11]), .CO(carry[12]), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry[10]), .CO(carry[11]), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry[9]), .CO(carry[10]), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry[8]), .CO(carry[9]), .S(SUM_8_)
         );
  ADDFX2 U1_22 ( .A(A_22_), .B(B_22_), .CI(carry[22]), .CO(carry[23]), .S(
        SUM_22_) );
  AND2X2 U1 ( .A(A_4_), .B(B_4_), .Y(n1) );
  XOR2X1 U2 ( .A(B_23_), .B(carry[23]), .Y(SUM_23_) );
  OAI2BB1X1 U3 ( .A0N(n2), .A1N(A_6_), .B0(n3), .Y(carry[7]) );
  OAI21XL U4 ( .A0(A_6_), .A1(n2), .B0(B_6_), .Y(n3) );
  OAI2BB1X1 U5 ( .A0N(n1), .A1N(A_5_), .B0(n4), .Y(n2) );
  OAI21XL U6 ( .A0(A_5_), .A1(n1), .B0(B_5_), .Y(n4) );
endmodule


module multi16_5_DW01_add_4 ( A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, 
        A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, 
        B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, 
        B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, SUM_22_, SUM_21_, SUM_20_, 
        SUM_19_, SUM_18_, SUM_17_, SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, 
        SUM_11_, SUM_10_, SUM_9_, SUM_8_, SUM_7_ );
  input A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_,
         A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, B_20_, B_19_,
         B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, B_10_, B_9_,
         B_8_, B_7_, B_6_, B_5_;
  output SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_,
         SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_,
         SUM_7_;
  wire   carry_21_, carry_20_, carry_19_, carry_18_, carry_17_, carry_16_,
         carry_15_, carry_14_, carry_13_, carry_12_, carry_11_, carry_10_,
         carry_9_, carry_8_, carry_7_, n1;

  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry_16_), .CO(carry_17_), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry_15_), .CO(carry_16_), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry_14_), .CO(carry_15_), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry_13_), .CO(carry_14_), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry_12_), .CO(carry_13_), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry_11_), .CO(carry_12_), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry_10_), .CO(carry_11_), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry_9_), .CO(carry_10_), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry_8_), .CO(carry_9_), .S(SUM_8_)
         );
  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry_7_), .CO(carry_8_), .S(SUM_7_)
         );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry_20_), .CO(carry_21_), .S(
        SUM_20_) );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry_19_), .CO(carry_20_), .S(
        SUM_19_) );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry_18_), .CO(carry_19_), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry_17_), .CO(carry_18_), .S(
        SUM_17_) );
  ADDFX2 U1_21 ( .A(A_21_), .B(B_21_), .CI(carry_21_), .CO(SUM_22_), .S(
        SUM_21_) );
  OAI2BB1X1 U1 ( .A0N(A_6_), .A1N(B_6_), .B0(n1), .Y(carry_7_) );
  OAI211X1 U2 ( .A0(B_6_), .A1(A_6_), .B0(A_5_), .C0(B_5_), .Y(n1) );
endmodule


module multi16_5_DW01_add_6 ( A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, 
        A_16_, A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, 
        A_6_, A_5_, A_4_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, 
        B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, 
        SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, 
        SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, 
        SUM_7_ );
  input A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_,
         A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, B_20_,
         B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, B_10_,
         B_9_, B_8_, B_7_, B_6_, B_5_, B_4_;
  output SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_,
         SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_,
         SUM_8_, SUM_7_;
  wire   n1, n2, n3, n4, n5, n6;
  wire   [21:7] carry;

  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry[7]), .CO(carry[8]), .S(SUM_7_)
         );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry[18]), .CO(carry[19]), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry[17]), .CO(carry[18]), .S(
        SUM_17_) );
  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry[16]), .CO(carry[17]), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry[15]), .CO(carry[16]), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry[14]), .CO(carry[15]), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry[13]), .CO(carry[14]), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry[12]), .CO(carry[13]), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry[11]), .CO(carry[12]), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry[10]), .CO(carry[11]), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry[9]), .CO(carry[10]), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry[8]), .CO(carry[9]), .S(SUM_8_)
         );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry[19]), .CO(carry[20]), .S(
        SUM_19_) );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry[20]), .CO(carry[21]), .S(
        SUM_20_) );
  AND2X2 U1 ( .A(A_22_), .B(n2), .Y(n1) );
  AND2X2 U2 ( .A(A_21_), .B(carry[21]), .Y(n2) );
  XOR2X1 U3 ( .A(A_23_), .B(n1), .Y(SUM_23_) );
  AND2X2 U4 ( .A(A_4_), .B(B_4_), .Y(n3) );
  XOR2X1 U5 ( .A(A_21_), .B(carry[21]), .Y(SUM_21_) );
  XOR2X1 U6 ( .A(A_22_), .B(n2), .Y(SUM_22_) );
  OAI2BB1X1 U7 ( .A0N(n4), .A1N(A_6_), .B0(n5), .Y(carry[7]) );
  OAI21XL U8 ( .A0(A_6_), .A1(n4), .B0(B_6_), .Y(n5) );
  OAI2BB1X1 U9 ( .A0N(n3), .A1N(A_5_), .B0(n6), .Y(n4) );
  OAI21XL U10 ( .A0(A_5_), .A1(n3), .B0(B_5_), .Y(n6) );
endmodule


module multi16_5 ( in_17bit, in_8bit, out );
  input [16:0] in_17bit;
  input [7:0] in_8bit;
  output [16:0] out;
  wire   n267, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26,
         N27, N28, N29, N108, N109, N110, N111, N112, N113, N114, N115, N116,
         N117, N118, N119, N120, N121, N122, N123, N205, N206, N207, N208,
         N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, N219,
         N220, N221, N347, N348, N349, N350, N351, N352, N353, N354, N355,
         N356, N357, N358, N359, N360, N361, N362, N363, N446, N447, N448,
         N449, N450, N451, N452, N453, N454, N455, N456, N457, N458, N459,
         N460, N461, N462, N463, N479, N480, N481, add_2_root_r119_carry_10_,
         add_2_root_r119_carry_11_, add_2_root_r119_carry_12_,
         add_2_root_r119_carry_13_, add_2_root_r119_carry_14_,
         add_2_root_r119_carry_15_, add_2_root_r119_carry_16_,
         add_2_root_r119_carry_17_, add_2_root_r119_carry_18_,
         add_2_root_r119_carry_19_, add_2_root_r119_carry_20_,
         add_2_root_r119_carry_21_, add_2_root_r119_carry_6_,
         add_2_root_r119_carry_7_, add_2_root_r119_carry_8_,
         add_2_root_r119_carry_9_, add_2_root_r119_SUM_5_,
         add_2_root_r119_SUM_6_, add_2_root_r119_SUM_7_,
         add_2_root_r119_SUM_8_, add_2_root_r119_SUM_9_,
         add_2_root_r119_SUM_10_, add_2_root_r119_SUM_11_,
         add_2_root_r119_SUM_12_, add_2_root_r119_SUM_13_,
         add_2_root_r119_SUM_14_, add_2_root_r119_SUM_15_,
         add_2_root_r119_SUM_16_, add_2_root_r119_SUM_17_,
         add_2_root_r119_SUM_18_, add_2_root_r119_SUM_19_,
         add_2_root_r119_SUM_20_, add_2_root_r119_SUM_21_,
         add_2_root_r119_SUM_22_, add_1_root_r119_SUM_6_,
         add_1_root_r119_SUM_7_, add_1_root_r119_SUM_8_,
         add_1_root_r119_SUM_9_, add_1_root_r119_SUM_10_,
         add_1_root_r119_SUM_11_, add_1_root_r119_SUM_12_,
         add_1_root_r119_SUM_13_, add_1_root_r119_SUM_14_,
         add_1_root_r119_SUM_15_, add_1_root_r119_SUM_16_,
         add_1_root_r119_SUM_17_, add_1_root_r119_SUM_18_,
         add_1_root_r119_SUM_19_, add_1_root_r119_SUM_20_,
         add_1_root_r119_SUM_21_, add_1_root_r119_SUM_22_,
         add_1_root_r119_SUM_23_, add_1_root_r119_A_2_, add_1_root_r119_A_3_,
         add_1_root_r119_A_4_, add_1_root_r119_A_5_, add_1_root_r119_A_6_,
         add_1_root_r119_A_7_, add_1_root_r119_A_8_, add_1_root_r119_A_9_,
         add_1_root_r119_A_10_, add_1_root_r119_A_11_, add_1_root_r119_A_12_,
         add_1_root_r119_A_13_, add_1_root_r119_A_14_, add_1_root_r119_A_15_,
         add_1_root_r119_A_16_, add_1_root_r119_A_17_, add_1_root_r119_A_18_,
         add_1_root_r119_A_19_, add_3_root_r119_carry_10_,
         add_3_root_r119_carry_11_, add_3_root_r119_carry_12_,
         add_3_root_r119_carry_13_, add_3_root_r119_carry_14_,
         add_3_root_r119_carry_15_, add_3_root_r119_carry_16_,
         add_3_root_r119_carry_17_, add_3_root_r119_carry_18_,
         add_3_root_r119_carry_3_, add_3_root_r119_carry_4_,
         add_3_root_r119_carry_5_, add_3_root_r119_carry_6_,
         add_3_root_r119_carry_7_, add_3_root_r119_carry_8_,
         add_3_root_r119_carry_9_, add_1_root_r112_carry_10_,
         add_1_root_r112_carry_11_, add_1_root_r112_carry_12_,
         add_1_root_r112_carry_13_, add_1_root_r112_carry_14_,
         add_1_root_r112_carry_15_, add_1_root_r112_carry_16_,
         add_1_root_r112_carry_17_, add_1_root_r112_carry_18_,
         add_1_root_r112_carry_19_, add_1_root_r112_carry_20_,
         add_1_root_r112_carry_5_, add_1_root_r112_carry_6_,
         add_1_root_r112_carry_7_, add_1_root_r112_carry_8_,
         add_1_root_r112_carry_9_, add_1_root_r112_SUM_1_,
         add_1_root_r112_SUM_2_, add_1_root_r112_SUM_3_,
         add_1_root_r112_SUM_4_, add_1_root_r112_SUM_5_,
         add_1_root_r112_SUM_6_, add_1_root_r112_SUM_7_,
         add_1_root_r112_SUM_8_, add_1_root_r112_SUM_9_,
         add_1_root_r112_SUM_10_, add_1_root_r112_SUM_11_,
         add_1_root_r112_SUM_12_, add_1_root_r112_SUM_13_,
         add_1_root_r112_SUM_14_, add_1_root_r112_SUM_15_,
         add_1_root_r112_SUM_16_, add_1_root_r112_SUM_17_,
         add_1_root_r112_SUM_18_, add_1_root_r112_SUM_19_,
         add_1_root_r112_SUM_20_, add_1_root_r112_SUM_21_,
         add_2_root_r115_carry_10_, add_2_root_r115_carry_11_,
         add_2_root_r115_carry_12_, add_2_root_r115_carry_13_,
         add_2_root_r115_carry_14_, add_2_root_r115_carry_15_,
         add_2_root_r115_carry_16_, add_2_root_r115_carry_17_,
         add_2_root_r115_carry_18_, add_2_root_r115_carry_19_,
         add_2_root_r115_carry_4_, add_2_root_r115_carry_5_,
         add_2_root_r115_carry_6_, add_2_root_r115_carry_7_,
         add_2_root_r115_carry_8_, add_2_root_r115_carry_9_,
         add_2_root_r115_SUM_3_, add_2_root_r115_SUM_4_,
         add_2_root_r115_SUM_5_, add_2_root_r115_SUM_6_,
         add_2_root_r115_SUM_7_, add_2_root_r115_SUM_8_,
         add_2_root_r115_SUM_9_, add_2_root_r115_SUM_10_,
         add_2_root_r115_SUM_11_, add_2_root_r115_SUM_12_,
         add_2_root_r115_SUM_13_, add_2_root_r115_SUM_14_,
         add_2_root_r115_SUM_15_, add_2_root_r115_SUM_16_,
         add_2_root_r115_SUM_17_, add_2_root_r115_SUM_18_,
         add_2_root_r115_SUM_19_, add_2_root_r115_SUM_20_,
         add_1_root_r115_carry_10_, add_1_root_r115_carry_11_,
         add_1_root_r115_carry_12_, add_1_root_r115_carry_13_,
         add_1_root_r115_carry_14_, add_1_root_r115_carry_15_,
         add_1_root_r115_carry_16_, add_1_root_r115_carry_17_,
         add_1_root_r115_carry_18_, add_1_root_r115_carry_19_,
         add_1_root_r115_carry_20_, add_1_root_r115_carry_21_,
         add_1_root_r115_carry_22_, add_1_root_r115_carry_7_,
         add_1_root_r115_carry_8_, add_1_root_r115_carry_9_,
         add_1_root_r115_SUM_6_, add_1_root_r115_SUM_7_,
         add_1_root_r115_SUM_8_, add_1_root_r115_SUM_9_,
         add_1_root_r115_SUM_10_, add_1_root_r115_SUM_11_,
         add_1_root_r115_SUM_12_, add_1_root_r115_SUM_13_,
         add_1_root_r115_SUM_14_, add_1_root_r115_SUM_15_,
         add_1_root_r115_SUM_16_, add_1_root_r115_SUM_17_,
         add_1_root_r115_SUM_18_, add_1_root_r115_SUM_19_,
         add_1_root_r115_SUM_20_, add_1_root_r115_SUM_21_,
         add_1_root_r115_SUM_22_, add_1_root_r115_SUM_23_, n2, n3, n4, n5, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n158, n160, n163,
         n164, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266;
  wire   [16:0] in_17bit_b;
  wire   [23:8] neg_mul;
  wire   [16:10] sub_add_75_b0_carry;
  wire   [15:2] sub_add_54_b0_carry;
  wire   [22:7] add_1_root_r119_carry;

  multi16_5_DW01_add_0 add_0_root_r119 ( .A_22_(add_2_root_r119_SUM_22_), 
        .A_21_(add_2_root_r119_SUM_21_), .A_20_(add_2_root_r119_SUM_20_), 
        .A_19_(add_2_root_r119_SUM_19_), .A_18_(add_2_root_r119_SUM_18_), 
        .A_17_(add_2_root_r119_SUM_17_), .A_16_(add_2_root_r119_SUM_16_), 
        .A_15_(add_2_root_r119_SUM_15_), .A_14_(add_2_root_r119_SUM_14_), 
        .A_13_(add_2_root_r119_SUM_13_), .A_12_(add_2_root_r119_SUM_12_), 
        .A_11_(add_2_root_r119_SUM_11_), .A_10_(add_2_root_r119_SUM_10_), 
        .A_9_(add_2_root_r119_SUM_9_), .A_8_(add_2_root_r119_SUM_8_), .A_7_(
        add_2_root_r119_SUM_7_), .A_6_(add_2_root_r119_SUM_6_), .A_5_(
        add_2_root_r119_SUM_5_), .A_4_(in_17bit_b[0]), .B_23_(
        add_1_root_r119_SUM_23_), .B_22_(add_1_root_r119_SUM_22_), .B_21_(
        add_1_root_r119_SUM_21_), .B_20_(add_1_root_r119_SUM_20_), .B_19_(
        add_1_root_r119_SUM_19_), .B_18_(add_1_root_r119_SUM_18_), .B_17_(
        add_1_root_r119_SUM_17_), .B_16_(add_1_root_r119_SUM_16_), .B_15_(
        add_1_root_r119_SUM_15_), .B_14_(add_1_root_r119_SUM_14_), .B_13_(
        add_1_root_r119_SUM_13_), .B_12_(add_1_root_r119_SUM_12_), .B_11_(
        add_1_root_r119_SUM_11_), .B_10_(add_1_root_r119_SUM_10_), .B_9_(
        add_1_root_r119_SUM_9_), .B_8_(add_1_root_r119_SUM_8_), .B_7_(
        add_1_root_r119_SUM_7_), .B_6_(add_1_root_r119_SUM_6_), .B_5_(
        add_1_root_r119_A_5_), .B_4_(add_1_root_r119_A_4_), .SUM_23_(N363), 
        .SUM_22_(N362), .SUM_21_(N361), .SUM_20_(N360), .SUM_19_(N359), 
        .SUM_18_(N358), .SUM_17_(N357), .SUM_16_(N356), .SUM_15_(N355), 
        .SUM_14_(N354), .SUM_13_(N353), .SUM_12_(N352), .SUM_11_(N351), 
        .SUM_10_(N350), .SUM_9_(N349), .SUM_8_(N348), .SUM_7_(N347) );
  multi16_5_DW01_add_4 add_0_root_r112 ( .A_21_(n38), .A_20_(in_17bit_b[15]), 
        .A_19_(in_17bit_b[14]), .A_18_(in_17bit_b[13]), .A_17_(in_17bit_b[12]), 
        .A_16_(in_17bit_b[11]), .A_15_(in_17bit_b[10]), .A_14_(in_17bit_b[9]), 
        .A_13_(in_17bit_b[8]), .A_12_(in_17bit_b[7]), .A_11_(in_17bit_b[6]), 
        .A_10_(in_17bit_b[5]), .A_9_(in_17bit_b[4]), .A_8_(in_17bit_b[3]), 
        .A_7_(in_17bit_b[2]), .A_6_(in_17bit_b[1]), .A_5_(in_17bit_b[0]), 
        .B_21_(add_1_root_r112_SUM_21_), .B_20_(add_1_root_r112_SUM_20_), 
        .B_19_(add_1_root_r112_SUM_19_), .B_18_(add_1_root_r112_SUM_18_), 
        .B_17_(add_1_root_r112_SUM_17_), .B_16_(add_1_root_r112_SUM_16_), 
        .B_15_(add_1_root_r112_SUM_15_), .B_14_(add_1_root_r112_SUM_14_), 
        .B_13_(add_1_root_r112_SUM_13_), .B_12_(add_1_root_r112_SUM_12_), 
        .B_11_(add_1_root_r112_SUM_11_), .B_10_(add_1_root_r112_SUM_10_), 
        .B_9_(add_1_root_r112_SUM_9_), .B_8_(add_1_root_r112_SUM_8_), .B_7_(
        add_1_root_r112_SUM_7_), .B_6_(add_1_root_r112_SUM_6_), .B_5_(
        add_1_root_r112_SUM_5_), .SUM_22_(N123), .SUM_21_(N122), .SUM_20_(N121), .SUM_19_(N120), .SUM_18_(N119), .SUM_17_(N118), .SUM_16_(N117), .SUM_15_(
        N116), .SUM_14_(N115), .SUM_13_(N114), .SUM_12_(N113), .SUM_11_(N112), 
        .SUM_10_(N111), .SUM_9_(N110), .SUM_8_(N109), .SUM_7_(N108) );
  multi16_5_DW01_add_6 add_0_root_r115 ( .A_23_(add_1_root_r115_SUM_23_), 
        .A_22_(add_1_root_r115_SUM_22_), .A_21_(add_1_root_r115_SUM_21_), 
        .A_20_(add_1_root_r115_SUM_20_), .A_19_(add_1_root_r115_SUM_19_), 
        .A_18_(add_1_root_r115_SUM_18_), .A_17_(add_1_root_r115_SUM_17_), 
        .A_16_(add_1_root_r115_SUM_16_), .A_15_(add_1_root_r115_SUM_15_), 
        .A_14_(add_1_root_r115_SUM_14_), .A_13_(add_1_root_r115_SUM_13_), 
        .A_12_(add_1_root_r115_SUM_12_), .A_11_(add_1_root_r115_SUM_11_), 
        .A_10_(add_1_root_r115_SUM_10_), .A_9_(add_1_root_r115_SUM_9_), .A_8_(
        add_1_root_r115_SUM_8_), .A_7_(add_1_root_r115_SUM_7_), .A_6_(
        add_1_root_r115_SUM_6_), .A_5_(in_17bit_b[1]), .A_4_(in_17bit_b[0]), 
        .B_20_(add_2_root_r115_SUM_20_), .B_19_(add_2_root_r115_SUM_19_), 
        .B_18_(add_2_root_r115_SUM_18_), .B_17_(add_2_root_r115_SUM_17_), 
        .B_16_(add_2_root_r115_SUM_16_), .B_15_(add_2_root_r115_SUM_15_), 
        .B_14_(add_2_root_r115_SUM_14_), .B_13_(add_2_root_r115_SUM_13_), 
        .B_12_(add_2_root_r115_SUM_12_), .B_11_(add_2_root_r115_SUM_11_), 
        .B_10_(add_2_root_r115_SUM_10_), .B_9_(add_2_root_r115_SUM_9_), .B_8_(
        add_2_root_r115_SUM_8_), .B_7_(add_2_root_r115_SUM_7_), .B_6_(
        add_2_root_r115_SUM_6_), .B_5_(add_2_root_r115_SUM_5_), .B_4_(
        add_2_root_r115_SUM_4_), .SUM_23_(N221), .SUM_22_(N220), .SUM_21_(N219), .SUM_20_(N218), .SUM_19_(N217), .SUM_18_(N216), .SUM_17_(N215), .SUM_16_(
        N214), .SUM_15_(N213), .SUM_14_(N212), .SUM_13_(N211), .SUM_12_(N210), 
        .SUM_11_(N209), .SUM_10_(N208), .SUM_9_(N207), .SUM_8_(N206), .SUM_7_(
        N205) );
  TLATX1 neg_mul_reg_16_ ( .G(N446), .D(N456), .QN(n8) );
  TLATX1 neg_mul_reg_15_ ( .G(N446), .D(N455), .QN(n5) );
  TLATX1 neg_mul_reg_14_ ( .G(N446), .D(N454), .QN(n7) );
  TLATX1 neg_mul_reg_13_ ( .G(N446), .D(N453), .QN(n6) );
  TLATX1 neg_mul_reg_12_ ( .G(N446), .D(N452), .Q(neg_mul[12]), .QN(n20) );
  TLATX1 neg_mul_reg_11_ ( .G(N446), .D(N451), .Q(n4), .QN(n13) );
  TLATX1 neg_mul_reg_23_ ( .G(N446), .D(N463), .Q(neg_mul[23]), .QN(n19) );
  TLATX1 neg_mul_reg_22_ ( .G(N446), .D(N462), .Q(neg_mul[22]), .QN(n11) );
  TLATX1 neg_mul_reg_21_ ( .G(N446), .D(N461), .Q(neg_mul[21]), .QN(n12) );
  TLATX1 neg_mul_reg_20_ ( .G(N446), .D(N460), .QN(n17) );
  TLATX1 neg_mul_reg_19_ ( .G(N446), .D(N459), .QN(n16) );
  TLATX1 neg_mul_reg_18_ ( .G(N446), .D(N458), .QN(n15) );
  TLATX1 neg_mul_reg_17_ ( .G(N446), .D(N457), .QN(n14) );
  TLATX1 neg_mul_reg_9_ ( .G(N446), .D(N449), .Q(neg_mul[9]), .QN(n10) );
  TLATX1 neg_mul_reg_10_ ( .G(N446), .D(N450), .Q(neg_mul[10]), .QN(n9) );
  TLATX1 neg_mul_reg_8_ ( .G(N446), .D(N448), .Q(neg_mul[8]), .QN(n18) );
  TLATX1 neg_mul_reg_7_ ( .G(N446), .D(N447), .Q(out[0]) );
  NOR2X2 U2 ( .A(n49), .B(n66), .Y(n68) );
  NAND4BX1 U3 ( .AN(n44), .B(n39), .C(in_8bit[1]), .D(in_8bit[4]), .Y(n98) );
  OAI21X4 U4 ( .A0(n3), .A1(n72), .B0(n71), .Y(n76) );
  OAI21X2 U5 ( .A0(n3), .A1(n64), .B0(n63), .Y(n69) );
  OAI21X2 U6 ( .A0(n3), .A1(n58), .B0(n57), .Y(n62) );
  MXI2X4 U7 ( .A(n15), .B(n31), .S0(n87), .Y(out[11]) );
  NAND2X2 U8 ( .A(n2), .B(n10), .Y(n63) );
  INVX8 U9 ( .A(in_8bit[7]), .Y(n45) );
  AOI2BB2X2 U10 ( .B0(n73), .B1(n3), .A0N(n44), .A1N(neg_mul[10]), .Y(n74) );
  AOI2BB2X2 U11 ( .B0(n65), .B1(n3), .A0N(n44), .A1N(neg_mul[9]), .Y(n66) );
  AOI2BB2X2 U12 ( .B0(n59), .B1(n3), .A0N(n44), .A1N(neg_mul[8]), .Y(n60) );
  CLKINVX4 U13 ( .A(n45), .Y(n44) );
  INVX4 U14 ( .A(n45), .Y(n43) );
  BUFX8 U15 ( .A(n267), .Y(out[3]) );
  AOI211X2 U16 ( .A0(n53), .A1(n76), .B0(n75), .C0(n78), .Y(n267) );
  NOR2X2 U17 ( .A(n53), .B(n74), .Y(n75) );
  MXI2X2 U18 ( .A(n16), .B(n33), .S0(n37), .Y(out[12]) );
  NOR2X2 U19 ( .A(n27), .B(n81), .Y(n82) );
  XNOR2X2 U20 ( .A(n24), .B(n5), .Y(out[8]) );
  BUFX3 U21 ( .A(n43), .Y(n2) );
  BUFX16 U22 ( .A(n43), .Y(n3) );
  BUFX12 U23 ( .A(n51), .Y(n22) );
  INVXL U24 ( .A(in_8bit[5]), .Y(n47) );
  BUFX3 U25 ( .A(n50), .Y(n21) );
  CLKINVX3 U26 ( .A(n22), .Y(n48) );
  INVX1 U27 ( .A(n22), .Y(n52) );
  NOR2BX2 U28 ( .AN(n22), .B(n60), .Y(n61) );
  XNOR2X1 U29 ( .A(n49), .B(n3), .Y(n83) );
  XOR2X4 U30 ( .A(n80), .B(neg_mul[12]), .Y(out[5]) );
  NAND2X2 U31 ( .A(n2), .B(n18), .Y(n57) );
  INVX8 U32 ( .A(n22), .Y(n49) );
  CLKINVX4 U33 ( .A(n22), .Y(n50) );
  NOR2X4 U34 ( .A(n28), .B(n83), .Y(n84) );
  INVXL U35 ( .A(n50), .Y(n54) );
  INVX8 U36 ( .A(n22), .Y(n53) );
  NOR2X4 U37 ( .A(n78), .B(n77), .Y(n23) );
  XNOR2X4 U38 ( .A(n21), .B(n3), .Y(n79) );
  NOR2X4 U39 ( .A(n26), .B(n79), .Y(n80) );
  INVX4 U40 ( .A(in_17bit[16]), .Y(n51) );
  INVX8 U41 ( .A(n86), .Y(n87) );
  NOR2X4 U42 ( .A(n86), .B(n30), .Y(n85) );
  XNOR2X4 U43 ( .A(n48), .B(n3), .Y(n86) );
  NAND2X2 U44 ( .A(n2), .B(n9), .Y(n71) );
  AOI211X4 U45 ( .A0(n53), .A1(n69), .B0(n68), .C0(n67), .Y(out[2]) );
  XOR2X2 U46 ( .A(n49), .B(n45), .Y(n77) );
  INVX1 U47 ( .A(n216), .Y(in_17bit_b[1]) );
  INVX1 U48 ( .A(n255), .Y(in_17bit_b[14]) );
  INVX1 U49 ( .A(n252), .Y(in_17bit_b[13]) );
  INVX1 U50 ( .A(n219), .Y(in_17bit_b[2]) );
  INVX1 U51 ( .A(n228), .Y(in_17bit_b[5]) );
  INVX1 U52 ( .A(n231), .Y(in_17bit_b[6]) );
  INVX1 U53 ( .A(n234), .Y(in_17bit_b[7]) );
  INVX1 U54 ( .A(n240), .Y(in_17bit_b[9]) );
  INVX1 U55 ( .A(n237), .Y(in_17bit_b[8]) );
  INVX1 U56 ( .A(n243), .Y(in_17bit_b[10]) );
  INVX1 U57 ( .A(n246), .Y(in_17bit_b[11]) );
  INVX1 U58 ( .A(n249), .Y(in_17bit_b[12]) );
  INVX1 U59 ( .A(n225), .Y(in_17bit_b[4]) );
  INVX1 U60 ( .A(n222), .Y(in_17bit_b[3]) );
  XOR2X4 U61 ( .A(n23), .B(n4), .Y(out[4]) );
  NOR2X2 U62 ( .A(n86), .B(n29), .Y(n24) );
  NAND4XL U63 ( .A(in_8bit[1]), .B(n44), .C(n203), .D(n183), .Y(n204) );
  OR4XL U64 ( .A(in_8bit[4]), .B(in_8bit[5]), .C(n39), .D(n44), .Y(n209) );
  INVX4 U65 ( .A(n77), .Y(n37) );
  NAND3X1 U66 ( .A(in_8bit[2]), .B(n42), .C(in_8bit[5]), .Y(n205) );
  NAND3BX1 U67 ( .AN(in_8bit[5]), .B(n46), .C(in_8bit[3]), .Y(n206) );
  NAND3X1 U68 ( .A(n3), .B(n41), .C(n47), .Y(n97) );
  INVX1 U69 ( .A(n40), .Y(n39) );
  OAI21XL U70 ( .A0(n265), .A1(n266), .B0(n264), .Y(N463) );
  AOI22X1 U71 ( .A0(N221), .A1(n263), .B0(N363), .B1(n262), .Y(n264) );
  INVX1 U72 ( .A(n182), .Y(n265) );
  ADDFX2 U73 ( .A(n38), .B(in_17bit_b[12]), .CI(add_1_root_r112_carry_16_), 
        .CO(add_1_root_r112_carry_17_), .S(add_1_root_r112_SUM_16_) );
  ADDFX2 U74 ( .A(add_1_root_r119_A_19_), .B(in_17bit_b[13]), .CI(
        add_1_root_r119_carry[19]), .CO(add_1_root_r119_carry[20]), .S(
        add_1_root_r119_SUM_19_) );
  ADDFX2 U75 ( .A(n38), .B(in_17bit_b[15]), .CI(add_3_root_r119_carry_17_), 
        .CO(add_3_root_r119_carry_18_), .S(add_1_root_r119_A_17_) );
  ADDFX2 U76 ( .A(n38), .B(in_17bit_b[14]), .CI(add_2_root_r115_carry_17_), 
        .CO(add_2_root_r115_carry_18_), .S(add_2_root_r115_SUM_17_) );
  ADDFX2 U77 ( .A(n38), .B(in_17bit_b[14]), .CI(add_1_root_r115_carry_20_), 
        .CO(add_1_root_r115_carry_21_), .S(add_1_root_r115_SUM_20_) );
  ADDFX2 U78 ( .A(n38), .B(in_17bit_b[15]), .CI(add_2_root_r119_carry_20_), 
        .CO(add_2_root_r119_carry_21_), .S(add_2_root_r119_SUM_20_) );
  INVX1 U79 ( .A(n52), .Y(n55) );
  ADDFX2 U80 ( .A(in_17bit_b[3]), .B(in_17bit_b[1]), .CI(
        add_2_root_r115_carry_4_), .CO(add_2_root_r115_carry_5_), .S(
        add_2_root_r115_SUM_4_) );
  ADDFX2 U81 ( .A(in_17bit_b[4]), .B(in_17bit_b[2]), .CI(
        add_2_root_r115_carry_5_), .CO(add_2_root_r115_carry_6_), .S(
        add_2_root_r115_SUM_5_) );
  ADDFX2 U82 ( .A(in_17bit_b[5]), .B(in_17bit_b[1]), .CI(
        add_1_root_r112_carry_5_), .CO(add_1_root_r112_carry_6_), .S(
        add_1_root_r112_SUM_5_) );
  ADDFX2 U83 ( .A(in_17bit_b[6]), .B(in_17bit_b[5]), .CI(
        add_3_root_r119_carry_7_), .CO(add_3_root_r119_carry_8_), .S(
        add_1_root_r119_A_7_) );
  ADDFX2 U84 ( .A(in_17bit_b[6]), .B(in_17bit_b[2]), .CI(
        add_1_root_r112_carry_6_), .CO(add_1_root_r112_carry_7_), .S(
        add_1_root_r112_SUM_6_) );
  ADDFX2 U85 ( .A(in_17bit_b[3]), .B(in_17bit_b[1]), .CI(
        add_1_root_r115_carry_7_), .CO(add_1_root_r115_carry_8_), .S(
        add_1_root_r115_SUM_7_) );
  ADDFX2 U86 ( .A(in_17bit_b[7]), .B(in_17bit_b[6]), .CI(
        add_3_root_r119_carry_8_), .CO(add_3_root_r119_carry_9_), .S(
        add_1_root_r119_A_8_) );
  ADDFX2 U87 ( .A(add_1_root_r119_A_7_), .B(in_17bit_b[1]), .CI(
        add_1_root_r119_carry[7]), .CO(add_1_root_r119_carry[8]), .S(
        add_1_root_r119_SUM_7_) );
  ADDFX2 U88 ( .A(in_17bit_b[2]), .B(in_17bit_b[1]), .CI(
        add_2_root_r119_carry_6_), .CO(add_2_root_r119_carry_7_), .S(
        add_2_root_r119_SUM_6_) );
  ADDFX2 U89 ( .A(in_17bit_b[4]), .B(in_17bit_b[2]), .CI(
        add_1_root_r115_carry_8_), .CO(add_1_root_r115_carry_9_), .S(
        add_1_root_r115_SUM_8_) );
  ADDFX2 U90 ( .A(in_17bit_b[8]), .B(in_17bit_b[7]), .CI(
        add_3_root_r119_carry_9_), .CO(add_3_root_r119_carry_10_), .S(
        add_1_root_r119_A_9_) );
  ADDFX2 U91 ( .A(add_1_root_r119_A_8_), .B(in_17bit_b[2]), .CI(
        add_1_root_r119_carry[8]), .CO(add_1_root_r119_carry[9]), .S(
        add_1_root_r119_SUM_8_) );
  ADDFX2 U92 ( .A(in_17bit_b[3]), .B(in_17bit_b[2]), .CI(
        add_2_root_r119_carry_7_), .CO(add_2_root_r119_carry_8_), .S(
        add_2_root_r119_SUM_7_) );
  ADDFX2 U93 ( .A(in_17bit_b[9]), .B(in_17bit_b[8]), .CI(
        add_3_root_r119_carry_10_), .CO(add_3_root_r119_carry_11_), .S(
        add_1_root_r119_A_10_) );
  ADDFX2 U94 ( .A(in_17bit_b[7]), .B(in_17bit_b[5]), .CI(
        add_2_root_r115_carry_8_), .CO(add_2_root_r115_carry_9_), .S(
        add_2_root_r115_SUM_8_) );
  ADDFX2 U95 ( .A(in_17bit_b[6]), .B(in_17bit_b[4]), .CI(
        add_1_root_r115_carry_10_), .CO(add_1_root_r115_carry_11_), .S(
        add_1_root_r115_SUM_10_) );
  ADDFX2 U96 ( .A(in_17bit_b[10]), .B(in_17bit_b[9]), .CI(
        add_3_root_r119_carry_11_), .CO(add_3_root_r119_carry_12_), .S(
        add_1_root_r119_A_11_) );
  ADDFX2 U97 ( .A(in_17bit_b[6]), .B(in_17bit_b[4]), .CI(
        add_2_root_r115_carry_7_), .CO(add_2_root_r115_carry_8_), .S(
        add_2_root_r115_SUM_7_) );
  ADDFX2 U98 ( .A(in_17bit_b[9]), .B(in_17bit_b[5]), .CI(
        add_1_root_r112_carry_9_), .CO(add_1_root_r112_carry_10_), .S(
        add_1_root_r112_SUM_9_) );
  ADDFX2 U99 ( .A(in_17bit_b[8]), .B(in_17bit_b[6]), .CI(
        add_2_root_r115_carry_9_), .CO(add_2_root_r115_carry_10_), .S(
        add_2_root_r115_SUM_9_) );
  ADDFX2 U100 ( .A(in_17bit_b[10]), .B(in_17bit_b[6]), .CI(
        add_1_root_r112_carry_10_), .CO(add_1_root_r112_carry_11_), .S(
        add_1_root_r112_SUM_10_) );
  ADDFX2 U101 ( .A(in_17bit_b[7]), .B(in_17bit_b[5]), .CI(
        add_1_root_r115_carry_11_), .CO(add_1_root_r115_carry_12_), .S(
        add_1_root_r115_SUM_11_) );
  ADDFX2 U102 ( .A(in_17bit_b[11]), .B(in_17bit_b[10]), .CI(
        add_3_root_r119_carry_12_), .CO(add_3_root_r119_carry_13_), .S(
        add_1_root_r119_A_12_) );
  ADDFX2 U103 ( .A(add_1_root_r119_A_11_), .B(in_17bit_b[5]), .CI(
        add_1_root_r119_carry[11]), .CO(add_1_root_r119_carry[12]), .S(
        add_1_root_r119_SUM_11_) );
  ADDFX2 U104 ( .A(in_17bit_b[6]), .B(in_17bit_b[5]), .CI(
        add_2_root_r119_carry_10_), .CO(add_2_root_r119_carry_11_), .S(
        add_2_root_r119_SUM_10_) );
  ADDFX2 U105 ( .A(in_17bit_b[9]), .B(in_17bit_b[7]), .CI(
        add_2_root_r115_carry_10_), .CO(add_2_root_r115_carry_11_), .S(
        add_2_root_r115_SUM_10_) );
  ADDFX2 U106 ( .A(in_17bit_b[11]), .B(in_17bit_b[7]), .CI(
        add_1_root_r112_carry_11_), .CO(add_1_root_r112_carry_12_), .S(
        add_1_root_r112_SUM_11_) );
  ADDFX2 U107 ( .A(in_17bit_b[8]), .B(in_17bit_b[6]), .CI(
        add_1_root_r115_carry_12_), .CO(add_1_root_r115_carry_13_), .S(
        add_1_root_r115_SUM_12_) );
  ADDFX2 U108 ( .A(in_17bit_b[12]), .B(in_17bit_b[11]), .CI(
        add_3_root_r119_carry_13_), .CO(add_3_root_r119_carry_14_), .S(
        add_1_root_r119_A_13_) );
  ADDFX2 U109 ( .A(add_1_root_r119_A_12_), .B(in_17bit_b[6]), .CI(
        add_1_root_r119_carry[12]), .CO(add_1_root_r119_carry[13]), .S(
        add_1_root_r119_SUM_12_) );
  ADDFX2 U110 ( .A(in_17bit_b[7]), .B(in_17bit_b[6]), .CI(
        add_2_root_r119_carry_11_), .CO(add_2_root_r119_carry_12_), .S(
        add_2_root_r119_SUM_11_) );
  ADDFX2 U111 ( .A(in_17bit_b[10]), .B(in_17bit_b[8]), .CI(
        add_2_root_r115_carry_11_), .CO(add_2_root_r115_carry_12_), .S(
        add_2_root_r115_SUM_11_) );
  ADDFX2 U112 ( .A(in_17bit_b[12]), .B(in_17bit_b[8]), .CI(
        add_1_root_r112_carry_12_), .CO(add_1_root_r112_carry_13_), .S(
        add_1_root_r112_SUM_12_) );
  ADDFX2 U113 ( .A(in_17bit_b[9]), .B(in_17bit_b[7]), .CI(
        add_1_root_r115_carry_13_), .CO(add_1_root_r115_carry_14_), .S(
        add_1_root_r115_SUM_13_) );
  ADDFX2 U114 ( .A(in_17bit_b[13]), .B(in_17bit_b[12]), .CI(
        add_3_root_r119_carry_14_), .CO(add_3_root_r119_carry_15_), .S(
        add_1_root_r119_A_14_) );
  ADDFX2 U115 ( .A(add_1_root_r119_A_13_), .B(in_17bit_b[7]), .CI(
        add_1_root_r119_carry[13]), .CO(add_1_root_r119_carry[14]), .S(
        add_1_root_r119_SUM_13_) );
  ADDFX2 U116 ( .A(in_17bit_b[8]), .B(in_17bit_b[7]), .CI(
        add_2_root_r119_carry_12_), .CO(add_2_root_r119_carry_13_), .S(
        add_2_root_r119_SUM_12_) );
  ADDFX2 U117 ( .A(in_17bit_b[11]), .B(in_17bit_b[9]), .CI(
        add_2_root_r115_carry_12_), .CO(add_2_root_r115_carry_13_), .S(
        add_2_root_r115_SUM_12_) );
  ADDFX2 U118 ( .A(in_17bit_b[13]), .B(in_17bit_b[9]), .CI(
        add_1_root_r112_carry_13_), .CO(add_1_root_r112_carry_14_), .S(
        add_1_root_r112_SUM_13_) );
  ADDFX2 U119 ( .A(in_17bit_b[10]), .B(in_17bit_b[8]), .CI(
        add_1_root_r115_carry_14_), .CO(add_1_root_r115_carry_15_), .S(
        add_1_root_r115_SUM_14_) );
  ADDFX2 U120 ( .A(in_17bit_b[14]), .B(in_17bit_b[13]), .CI(
        add_3_root_r119_carry_15_), .CO(add_3_root_r119_carry_16_), .S(
        add_1_root_r119_A_15_) );
  ADDFX2 U121 ( .A(add_1_root_r119_A_14_), .B(in_17bit_b[8]), .CI(
        add_1_root_r119_carry[14]), .CO(add_1_root_r119_carry[15]), .S(
        add_1_root_r119_SUM_14_) );
  ADDFX2 U122 ( .A(in_17bit_b[3]), .B(in_17bit_b[2]), .CI(
        add_3_root_r119_carry_4_), .CO(add_3_root_r119_carry_5_), .S(
        add_1_root_r119_A_4_) );
  ADDFX2 U123 ( .A(in_17bit_b[2]), .B(in_17bit_b[1]), .CI(
        add_3_root_r119_carry_3_), .CO(add_3_root_r119_carry_4_), .S(
        add_1_root_r119_A_3_) );
  ADDFX2 U124 ( .A(in_17bit_b[9]), .B(in_17bit_b[8]), .CI(
        add_2_root_r119_carry_13_), .CO(add_2_root_r119_carry_14_), .S(
        add_2_root_r119_SUM_13_) );
  ADDFX2 U125 ( .A(in_17bit_b[12]), .B(in_17bit_b[10]), .CI(
        add_2_root_r115_carry_13_), .CO(add_2_root_r115_carry_14_), .S(
        add_2_root_r115_SUM_13_) );
  ADDFX2 U126 ( .A(in_17bit_b[11]), .B(in_17bit_b[9]), .CI(
        add_1_root_r115_carry_15_), .CO(add_1_root_r115_carry_16_), .S(
        add_1_root_r115_SUM_15_) );
  ADDFX2 U127 ( .A(add_1_root_r119_A_15_), .B(in_17bit_b[9]), .CI(
        add_1_root_r119_carry[15]), .CO(add_1_root_r119_carry[16]), .S(
        add_1_root_r119_SUM_15_) );
  ADDFX2 U128 ( .A(in_17bit_b[10]), .B(in_17bit_b[9]), .CI(
        add_2_root_r119_carry_14_), .CO(add_2_root_r119_carry_15_), .S(
        add_2_root_r119_SUM_14_) );
  ADDFX2 U129 ( .A(in_17bit_b[13]), .B(in_17bit_b[11]), .CI(
        add_2_root_r115_carry_14_), .CO(add_2_root_r115_carry_15_), .S(
        add_2_root_r115_SUM_14_) );
  ADDFX2 U130 ( .A(in_17bit_b[15]), .B(in_17bit_b[11]), .CI(
        add_1_root_r112_carry_15_), .CO(add_1_root_r112_carry_16_), .S(
        add_1_root_r112_SUM_15_) );
  ADDFX2 U131 ( .A(in_17bit_b[12]), .B(in_17bit_b[10]), .CI(
        add_1_root_r115_carry_16_), .CO(add_1_root_r115_carry_17_), .S(
        add_1_root_r115_SUM_16_) );
  ADDFX2 U132 ( .A(add_1_root_r119_A_16_), .B(in_17bit_b[10]), .CI(
        add_1_root_r119_carry[16]), .CO(add_1_root_r119_carry[17]), .S(
        add_1_root_r119_SUM_16_) );
  ADDFX2 U133 ( .A(in_17bit_b[11]), .B(in_17bit_b[10]), .CI(
        add_2_root_r119_carry_15_), .CO(add_2_root_r119_carry_16_), .S(
        add_2_root_r119_SUM_15_) );
  ADDFX2 U134 ( .A(in_17bit_b[14]), .B(in_17bit_b[12]), .CI(
        add_2_root_r115_carry_15_), .CO(add_2_root_r115_carry_16_), .S(
        add_2_root_r115_SUM_15_) );
  ADDFX2 U135 ( .A(in_17bit_b[13]), .B(in_17bit_b[11]), .CI(
        add_1_root_r115_carry_17_), .CO(add_1_root_r115_carry_18_), .S(
        add_1_root_r115_SUM_17_) );
  ADDFX2 U136 ( .A(in_17bit_b[12]), .B(in_17bit_b[11]), .CI(
        add_2_root_r119_carry_16_), .CO(add_2_root_r119_carry_17_), .S(
        add_2_root_r119_SUM_16_) );
  ADDFX2 U137 ( .A(in_17bit_b[15]), .B(in_17bit_b[13]), .CI(
        add_2_root_r115_carry_16_), .CO(add_2_root_r115_carry_17_), .S(
        add_2_root_r115_SUM_16_) );
  ADDFX2 U138 ( .A(in_17bit_b[14]), .B(in_17bit_b[12]), .CI(
        add_1_root_r115_carry_18_), .CO(add_1_root_r115_carry_19_), .S(
        add_1_root_r115_SUM_18_) );
  ADDFX2 U139 ( .A(add_1_root_r119_A_18_), .B(in_17bit_b[12]), .CI(
        add_1_root_r119_carry[18]), .CO(add_1_root_r119_carry[19]), .S(
        add_1_root_r119_SUM_18_) );
  ADDFX2 U140 ( .A(in_17bit_b[13]), .B(in_17bit_b[12]), .CI(
        add_2_root_r119_carry_17_), .CO(add_2_root_r119_carry_18_), .S(
        add_2_root_r119_SUM_17_) );
  ADDFX2 U141 ( .A(in_17bit_b[14]), .B(in_17bit_b[13]), .CI(
        add_2_root_r119_carry_18_), .CO(add_2_root_r119_carry_19_), .S(
        add_2_root_r119_SUM_18_) );
  ADDFX2 U142 ( .A(in_17bit_b[5]), .B(in_17bit_b[3]), .CI(
        add_2_root_r115_carry_6_), .CO(add_2_root_r115_carry_7_), .S(
        add_2_root_r115_SUM_6_) );
  ADDFX2 U143 ( .A(in_17bit_b[7]), .B(in_17bit_b[3]), .CI(
        add_1_root_r112_carry_7_), .CO(add_1_root_r112_carry_8_), .S(
        add_1_root_r112_SUM_7_) );
  ADDFX2 U144 ( .A(in_17bit_b[8]), .B(in_17bit_b[4]), .CI(
        add_1_root_r112_carry_8_), .CO(add_1_root_r112_carry_9_), .S(
        add_1_root_r112_SUM_8_) );
  ADDFX2 U145 ( .A(in_17bit_b[5]), .B(in_17bit_b[3]), .CI(
        add_1_root_r115_carry_9_), .CO(add_1_root_r115_carry_10_), .S(
        add_1_root_r115_SUM_9_) );
  ADDFX2 U146 ( .A(in_17bit_b[4]), .B(in_17bit_b[3]), .CI(
        add_2_root_r119_carry_8_), .CO(add_2_root_r119_carry_9_), .S(
        add_2_root_r119_SUM_8_) );
  ADDFX2 U147 ( .A(add_1_root_r119_A_10_), .B(in_17bit_b[4]), .CI(
        add_1_root_r119_carry[10]), .CO(add_1_root_r119_carry[11]), .S(
        add_1_root_r119_SUM_10_) );
  ADDFX2 U148 ( .A(in_17bit_b[5]), .B(in_17bit_b[4]), .CI(
        add_2_root_r119_carry_9_), .CO(add_2_root_r119_carry_10_), .S(
        add_2_root_r119_SUM_9_) );
  ADDFX2 U149 ( .A(in_17bit_b[14]), .B(in_17bit_b[10]), .CI(
        add_1_root_r112_carry_14_), .CO(add_1_root_r112_carry_15_), .S(
        add_1_root_r112_SUM_14_) );
  ADDFX2 U150 ( .A(add_1_root_r119_A_17_), .B(in_17bit_b[11]), .CI(
        add_1_root_r119_carry[17]), .CO(add_1_root_r119_carry[18]), .S(
        add_1_root_r119_SUM_17_) );
  ADDFX2 U151 ( .A(in_17bit_b[15]), .B(in_17bit_b[14]), .CI(
        add_3_root_r119_carry_16_), .CO(add_3_root_r119_carry_17_), .S(
        add_1_root_r119_A_16_) );
  ADDFX2 U152 ( .A(add_1_root_r119_A_9_), .B(in_17bit_b[3]), .CI(
        add_1_root_r119_carry[9]), .CO(add_1_root_r119_carry[10]), .S(
        add_1_root_r119_SUM_9_) );
  ADDFX2 U153 ( .A(in_17bit_b[5]), .B(in_17bit_b[4]), .CI(
        add_3_root_r119_carry_6_), .CO(add_3_root_r119_carry_7_), .S(
        add_1_root_r119_A_6_) );
  ADDFX2 U154 ( .A(in_17bit_b[15]), .B(in_17bit_b[13]), .CI(
        add_1_root_r115_carry_19_), .CO(add_1_root_r115_carry_20_), .S(
        add_1_root_r115_SUM_19_) );
  ADDFX2 U155 ( .A(in_17bit_b[4]), .B(in_17bit_b[3]), .CI(
        add_3_root_r119_carry_5_), .CO(add_3_root_r119_carry_6_), .S(
        add_1_root_r119_A_5_) );
  ADDFX2 U156 ( .A(in_17bit_b[15]), .B(in_17bit_b[14]), .CI(
        add_2_root_r119_carry_19_), .CO(add_2_root_r119_carry_20_), .S(
        add_2_root_r119_SUM_19_) );
  INVX1 U157 ( .A(n211), .Y(n88) );
  BUFX3 U158 ( .A(in_17bit_b[16]), .Y(n38) );
  INVX1 U159 ( .A(n266), .Y(in_17bit_b[16]) );
  INVX1 U160 ( .A(in_8bit[2]), .Y(n46) );
  INVX1 U161 ( .A(in_8bit[3]), .Y(n42) );
  INVX1 U162 ( .A(in_8bit[6]), .Y(n40) );
  INVX1 U163 ( .A(in_8bit[4]), .Y(n41) );
  XNOR2X1 U164 ( .A(n55), .B(n25), .Y(N29) );
  NAND2X1 U165 ( .A(sub_add_54_b0_carry[15]), .B(n180), .Y(n25) );
  CLKINVX3 U166 ( .A(n213), .Y(in_17bit_b[0]) );
  NOR3X1 U167 ( .A(n46), .B(n42), .C(n183), .Y(n211) );
  NAND4BXL U168 ( .AN(n44), .B(in_8bit[4]), .C(in_8bit[5]), .D(n210), .Y(n89)
         );
  CLKINVX3 U169 ( .A(n258), .Y(in_17bit_b[15]) );
  OR2X2 U170 ( .A(n93), .B(n92), .Y(n262) );
  NOR2X1 U171 ( .A(n94), .B(n205), .Y(n92) );
  NOR2X1 U172 ( .A(n206), .B(n204), .Y(n93) );
  OR2X2 U173 ( .A(n96), .B(n95), .Y(n263) );
  NOR2X1 U174 ( .A(n94), .B(n206), .Y(n95) );
  NOR2X1 U175 ( .A(n205), .B(n204), .Y(n96) );
  OAI2BB1X1 U176 ( .A0N(n210), .A1N(n100), .B0(n99), .Y(n182) );
  INVX1 U177 ( .A(n97), .Y(n100) );
  NAND3BX1 U178 ( .AN(n98), .B(n211), .C(in_8bit[5]), .Y(n99) );
  NAND2X1 U179 ( .A(n215), .B(n214), .Y(N447) );
  AOI22X1 U180 ( .A0(N108), .A1(n259), .B0(N205), .B1(n263), .Y(n214) );
  AOI22X1 U181 ( .A0(N347), .A1(n262), .B0(n182), .B1(in_17bit_b[0]), .Y(n215)
         );
  NAND2X1 U182 ( .A(n218), .B(n217), .Y(N448) );
  AOI22X1 U183 ( .A0(N109), .A1(n259), .B0(N206), .B1(n263), .Y(n217) );
  AOI22X1 U184 ( .A0(N348), .A1(n262), .B0(n182), .B1(n181), .Y(n218) );
  INVX1 U185 ( .A(n216), .Y(n181) );
  NAND2X1 U186 ( .A(n221), .B(n220), .Y(N449) );
  AOI22X1 U187 ( .A0(N110), .A1(n259), .B0(N207), .B1(n263), .Y(n220) );
  AOI22X1 U188 ( .A0(N349), .A1(n262), .B0(n182), .B1(in_17bit_b[2]), .Y(n221)
         );
  NAND2X1 U189 ( .A(n224), .B(n223), .Y(N450) );
  AOI22X1 U190 ( .A0(N111), .A1(n259), .B0(N208), .B1(n263), .Y(n223) );
  AOI22X1 U191 ( .A0(N350), .A1(n262), .B0(n182), .B1(in_17bit_b[3]), .Y(n224)
         );
  NAND2X1 U192 ( .A(n227), .B(n226), .Y(N451) );
  AOI22X1 U193 ( .A0(N112), .A1(n259), .B0(N209), .B1(n263), .Y(n226) );
  AOI22X1 U194 ( .A0(N351), .A1(n262), .B0(n182), .B1(in_17bit_b[4]), .Y(n227)
         );
  NAND2X1 U195 ( .A(n230), .B(n229), .Y(N452) );
  AOI22X1 U196 ( .A0(N113), .A1(n259), .B0(N210), .B1(n263), .Y(n229) );
  AOI22X1 U197 ( .A0(N352), .A1(n262), .B0(n182), .B1(in_17bit_b[5]), .Y(n230)
         );
  NAND2X1 U198 ( .A(n233), .B(n232), .Y(N453) );
  AOI22X1 U199 ( .A0(N114), .A1(n259), .B0(N211), .B1(n263), .Y(n232) );
  AOI22X1 U200 ( .A0(N353), .A1(n262), .B0(n182), .B1(in_17bit_b[6]), .Y(n233)
         );
  NAND2X1 U201 ( .A(n236), .B(n235), .Y(N454) );
  AOI22X1 U202 ( .A0(N115), .A1(n259), .B0(N212), .B1(n263), .Y(n235) );
  AOI22X1 U203 ( .A0(N354), .A1(n262), .B0(n182), .B1(in_17bit_b[7]), .Y(n236)
         );
  NAND2X1 U204 ( .A(n239), .B(n238), .Y(N455) );
  AOI22X1 U205 ( .A0(N116), .A1(n259), .B0(N213), .B1(n263), .Y(n238) );
  AOI22X1 U206 ( .A0(N355), .A1(n262), .B0(n182), .B1(in_17bit_b[8]), .Y(n239)
         );
  NAND2X1 U207 ( .A(n242), .B(n241), .Y(N456) );
  AOI22X1 U208 ( .A0(N117), .A1(n259), .B0(N214), .B1(n263), .Y(n241) );
  AOI22X1 U209 ( .A0(N356), .A1(n262), .B0(n182), .B1(in_17bit_b[9]), .Y(n242)
         );
  NAND2X1 U210 ( .A(n245), .B(n244), .Y(N457) );
  AOI22X1 U211 ( .A0(N118), .A1(n259), .B0(N215), .B1(n263), .Y(n244) );
  AOI22X1 U212 ( .A0(N357), .A1(n262), .B0(n182), .B1(in_17bit_b[10]), .Y(n245) );
  NAND2X1 U213 ( .A(n248), .B(n247), .Y(N458) );
  AOI22X1 U214 ( .A0(N119), .A1(n259), .B0(N216), .B1(n263), .Y(n247) );
  AOI22X1 U215 ( .A0(N358), .A1(n262), .B0(n182), .B1(in_17bit_b[11]), .Y(n248) );
  NAND2X1 U216 ( .A(n251), .B(n250), .Y(N459) );
  AOI22X1 U217 ( .A0(N120), .A1(n259), .B0(N217), .B1(n263), .Y(n250) );
  AOI22X1 U218 ( .A0(N359), .A1(n262), .B0(n182), .B1(in_17bit_b[12]), .Y(n251) );
  NAND2X1 U219 ( .A(n254), .B(n253), .Y(N460) );
  AOI22X1 U220 ( .A0(N121), .A1(n259), .B0(N218), .B1(n263), .Y(n253) );
  AOI22X1 U221 ( .A0(N360), .A1(n262), .B0(n182), .B1(in_17bit_b[13]), .Y(n254) );
  NAND2X1 U222 ( .A(n257), .B(n256), .Y(N461) );
  AOI22X1 U223 ( .A0(N122), .A1(n259), .B0(N219), .B1(n263), .Y(n256) );
  AOI22X1 U224 ( .A0(N361), .A1(n262), .B0(n182), .B1(in_17bit_b[14]), .Y(n257) );
  NAND2X1 U225 ( .A(n261), .B(n260), .Y(N462) );
  AOI22X1 U226 ( .A0(N123), .A1(n259), .B0(N220), .B1(n263), .Y(n260) );
  AOI22X1 U227 ( .A0(N362), .A1(n262), .B0(n182), .B1(in_17bit_b[15]), .Y(n261) );
  INVX1 U228 ( .A(n70), .Y(n67) );
  XNOR2X1 U229 ( .A(n49), .B(n3), .Y(n81) );
  NAND4BBX1 U230 ( .AN(n262), .BN(n263), .C(n212), .D(n265), .Y(N446) );
  AOI2BB1X1 U231 ( .A0N(n209), .A1N(n208), .B0(n259), .Y(n212) );
  NOR2X1 U232 ( .A(n39), .B(in_8bit[4]), .Y(n203) );
  NOR4BX1 U233 ( .AN(n207), .B(n183), .C(in_8bit[1]), .D(in_8bit[2]), .Y(n210)
         );
  NOR2X1 U234 ( .A(n39), .B(in_8bit[3]), .Y(n207) );
  INVXL U235 ( .A(in_8bit[0]), .Y(n183) );
  AOI22X1 U236 ( .A0(N28), .A1(n52), .B0(in_17bit[15]), .B1(n54), .Y(n258) );
  AOI22X1 U237 ( .A0(N17), .A1(n52), .B0(in_17bit[4]), .B1(n54), .Y(n225) );
  AOI22X1 U238 ( .A0(N18), .A1(n52), .B0(in_17bit[5]), .B1(n55), .Y(n228) );
  AOI22X1 U239 ( .A0(N19), .A1(n52), .B0(in_17bit[6]), .B1(n54), .Y(n231) );
  AOI22X1 U240 ( .A0(N16), .A1(n52), .B0(in_17bit[3]), .B1(n54), .Y(n222) );
  AOI22X1 U241 ( .A0(N27), .A1(n52), .B0(in_17bit[14]), .B1(n55), .Y(n255) );
  AOI22X1 U242 ( .A0(N26), .A1(n52), .B0(in_17bit[13]), .B1(n54), .Y(n252) );
  AOI22X1 U243 ( .A0(N20), .A1(n52), .B0(in_17bit[7]), .B1(n54), .Y(n234) );
  AOI22X1 U244 ( .A0(N21), .A1(n52), .B0(in_17bit[8]), .B1(n55), .Y(n237) );
  AOI22X1 U245 ( .A0(N22), .A1(n52), .B0(in_17bit[9]), .B1(n55), .Y(n240) );
  AOI22X1 U246 ( .A0(N23), .A1(n52), .B0(in_17bit[10]), .B1(n54), .Y(n243) );
  AOI22X1 U247 ( .A0(N24), .A1(n52), .B0(in_17bit[11]), .B1(n55), .Y(n246) );
  AOI22X1 U248 ( .A0(N25), .A1(n52), .B0(in_17bit[12]), .B1(n54), .Y(n249) );
  INVX1 U249 ( .A(n56), .Y(n78) );
  NAND2BX1 U250 ( .AN(n70), .B(n9), .Y(n56) );
  NAND2X1 U251 ( .A(n35), .B(n10), .Y(n70) );
  AND2X2 U252 ( .A(n78), .B(n13), .Y(n26) );
  AND2X2 U253 ( .A(n26), .B(n20), .Y(n27) );
  AND2X2 U254 ( .A(n27), .B(n6), .Y(n28) );
  OR2XL U255 ( .A(n98), .B(in_8bit[0]), .Y(n94) );
  AND2X2 U256 ( .A(n28), .B(n7), .Y(n29) );
  OAI2BB1X1 U257 ( .A0N(n91), .A1N(n90), .B0(n89), .Y(n259) );
  NOR2X1 U258 ( .A(n40), .B(n88), .Y(n91) );
  NOR2BX1 U259 ( .AN(in_8bit[1]), .B(n97), .Y(n90) );
  AND2X2 U260 ( .A(n29), .B(n5), .Y(n30) );
  INVX1 U261 ( .A(in_17bit[13]), .Y(n178) );
  INVX1 U262 ( .A(in_17bit[3]), .Y(n163) );
  INVX1 U263 ( .A(in_17bit[4]), .Y(n164) );
  INVX1 U264 ( .A(in_17bit[5]), .Y(n170) );
  INVX1 U265 ( .A(in_17bit[6]), .Y(n171) );
  INVX1 U266 ( .A(in_17bit[7]), .Y(n172) );
  INVX1 U267 ( .A(in_17bit[8]), .Y(n173) );
  INVX1 U268 ( .A(in_17bit[9]), .Y(n174) );
  INVX1 U269 ( .A(in_17bit[10]), .Y(n175) );
  INVX1 U270 ( .A(in_17bit[11]), .Y(n176) );
  INVX1 U271 ( .A(in_17bit[12]), .Y(n177) );
  INVX1 U272 ( .A(in_17bit[14]), .Y(n179) );
  INVX1 U273 ( .A(in_17bit[15]), .Y(n180) );
  INVX1 U274 ( .A(in_17bit[1]), .Y(n158) );
  INVX1 U275 ( .A(in_17bit[2]), .Y(n160) );
  INVX1 U276 ( .A(in_17bit[0]), .Y(n101) );
  XNOR2X1 U277 ( .A(n15), .B(sub_add_75_b0_carry[11]), .Y(n31) );
  XNOR2X1 U278 ( .A(n14), .B(sub_add_75_b0_carry[10]), .Y(n32) );
  XNOR2X1 U279 ( .A(n16), .B(sub_add_75_b0_carry[12]), .Y(n33) );
  XNOR2X1 U280 ( .A(n17), .B(sub_add_75_b0_carry[13]), .Y(n34) );
  MX2X1 U281 ( .A(neg_mul[21]), .B(N479), .S0(n37), .Y(out[14]) );
  MX2X1 U282 ( .A(neg_mul[22]), .B(N480), .S0(n37), .Y(out[15]) );
  INVX1 U283 ( .A(n64), .Y(n65) );
  INVX1 U284 ( .A(n58), .Y(n59) );
  INVX1 U285 ( .A(n72), .Y(n73) );
  MX2X1 U286 ( .A(neg_mul[23]), .B(N481), .S0(n37), .Y(out[16]) );
  NOR2X1 U287 ( .A(out[0]), .B(neg_mul[8]), .Y(n35) );
  NAND2BX1 U288 ( .AN(n35), .B(neg_mul[9]), .Y(n64) );
  NAND2X1 U289 ( .A(out[0]), .B(neg_mul[8]), .Y(n58) );
  NAND2X1 U290 ( .A(neg_mul[10]), .B(n70), .Y(n72) );
  AOI211X4 U291 ( .A0(n49), .A1(n62), .B0(n61), .C0(n35), .Y(out[1]) );
  NAND2XL U292 ( .A(N29), .B(n49), .Y(n266) );
  AOI22XL U293 ( .A0(N15), .A1(n21), .B0(in_17bit[2]), .B1(n54), .Y(n219) );
  AOI22XL U294 ( .A0(N14), .A1(n52), .B0(in_17bit[1]), .B1(n55), .Y(n216) );
  AOI22XL U295 ( .A0(in_17bit[0]), .A1(n50), .B0(in_17bit[0]), .B1(n55), .Y(
        n213) );
  OR4X1 U296 ( .A(in_8bit[1]), .B(in_8bit[0]), .C(in_8bit[2]), .D(in_8bit[3]), 
        .Y(n208) );
  XNOR2X4 U297 ( .A(n82), .B(n6), .Y(out[6]) );
  XNOR2X4 U298 ( .A(n84), .B(n7), .Y(out[7]) );
  XNOR2X4 U299 ( .A(n85), .B(n8), .Y(out[9]) );
  MXI2X4 U300 ( .A(n14), .B(n32), .S0(n87), .Y(out[10]) );
  MXI2X4 U301 ( .A(n17), .B(n34), .S0(n37), .Y(out[13]) );
  AND2X1 U302 ( .A(add_1_root_r112_carry_20_), .B(n38), .Y(
        add_1_root_r112_SUM_21_) );
  XOR2X1 U303 ( .A(n38), .B(add_1_root_r112_carry_20_), .Y(
        add_1_root_r112_SUM_20_) );
  AND2X1 U304 ( .A(add_1_root_r112_carry_19_), .B(in_17bit_b[15]), .Y(
        add_1_root_r112_carry_20_) );
  XOR2X1 U305 ( .A(in_17bit_b[15]), .B(add_1_root_r112_carry_19_), .Y(
        add_1_root_r112_SUM_19_) );
  AND2X1 U306 ( .A(add_1_root_r112_carry_18_), .B(in_17bit_b[14]), .Y(
        add_1_root_r112_carry_19_) );
  XOR2X1 U307 ( .A(in_17bit_b[14]), .B(add_1_root_r112_carry_18_), .Y(
        add_1_root_r112_SUM_18_) );
  AND2X1 U308 ( .A(add_1_root_r112_carry_17_), .B(in_17bit_b[13]), .Y(
        add_1_root_r112_carry_18_) );
  XOR2X1 U309 ( .A(in_17bit_b[13]), .B(add_1_root_r112_carry_17_), .Y(
        add_1_root_r112_SUM_17_) );
  AND2X1 U310 ( .A(add_2_root_r119_carry_21_), .B(n38), .Y(
        add_2_root_r119_SUM_22_) );
  XOR2X1 U311 ( .A(n38), .B(add_2_root_r119_carry_21_), .Y(
        add_2_root_r119_SUM_21_) );
  AND2X1 U312 ( .A(in_17bit_b[1]), .B(in_17bit_b[0]), .Y(
        add_2_root_r119_carry_6_) );
  XOR2X1 U313 ( .A(in_17bit_b[0]), .B(in_17bit_b[1]), .Y(
        add_2_root_r119_SUM_5_) );
  AND2X1 U314 ( .A(add_1_root_r119_carry[22]), .B(n38), .Y(
        add_1_root_r119_SUM_23_) );
  XOR2X1 U315 ( .A(n38), .B(add_1_root_r119_carry[22]), .Y(
        add_1_root_r119_SUM_22_) );
  AND2X1 U316 ( .A(add_1_root_r119_carry[21]), .B(in_17bit_b[15]), .Y(
        add_1_root_r119_carry[22]) );
  XOR2X1 U317 ( .A(in_17bit_b[15]), .B(add_1_root_r119_carry[21]), .Y(
        add_1_root_r119_SUM_21_) );
  AND2X1 U318 ( .A(add_1_root_r119_carry[20]), .B(in_17bit_b[14]), .Y(
        add_1_root_r119_carry[21]) );
  XOR2X1 U319 ( .A(in_17bit_b[14]), .B(add_1_root_r119_carry[20]), .Y(
        add_1_root_r119_SUM_20_) );
  AND2X1 U320 ( .A(add_1_root_r119_A_6_), .B(in_17bit_b[0]), .Y(
        add_1_root_r119_carry[7]) );
  XOR2X1 U321 ( .A(in_17bit_b[0]), .B(add_1_root_r119_A_6_), .Y(
        add_1_root_r119_SUM_6_) );
  AND2X1 U322 ( .A(add_3_root_r119_carry_18_), .B(n38), .Y(
        add_1_root_r119_A_19_) );
  XOR2X1 U323 ( .A(n38), .B(add_3_root_r119_carry_18_), .Y(
        add_1_root_r119_A_18_) );
  AND2X1 U324 ( .A(in_17bit_b[1]), .B(in_17bit_b[0]), .Y(
        add_3_root_r119_carry_3_) );
  XOR2X1 U325 ( .A(in_17bit_b[0]), .B(in_17bit_b[1]), .Y(add_1_root_r119_A_2_)
         );
  AND2X1 U326 ( .A(add_2_root_r115_carry_19_), .B(n38), .Y(
        add_2_root_r115_SUM_20_) );
  XOR2X1 U327 ( .A(n38), .B(add_2_root_r115_carry_19_), .Y(
        add_2_root_r115_SUM_19_) );
  AND2X1 U328 ( .A(add_2_root_r115_carry_18_), .B(in_17bit_b[15]), .Y(
        add_2_root_r115_carry_19_) );
  XOR2X1 U329 ( .A(in_17bit_b[15]), .B(add_2_root_r115_carry_18_), .Y(
        add_2_root_r115_SUM_18_) );
  AND2X1 U330 ( .A(in_17bit_b[2]), .B(in_17bit_b[0]), .Y(
        add_2_root_r115_carry_4_) );
  XOR2X1 U331 ( .A(in_17bit_b[0]), .B(in_17bit_b[2]), .Y(
        add_2_root_r115_SUM_3_) );
  AND2X1 U332 ( .A(add_1_root_r115_carry_22_), .B(n38), .Y(
        add_1_root_r115_SUM_23_) );
  XOR2X1 U333 ( .A(n38), .B(add_1_root_r115_carry_22_), .Y(
        add_1_root_r115_SUM_22_) );
  AND2X1 U334 ( .A(add_1_root_r115_carry_21_), .B(in_17bit_b[15]), .Y(
        add_1_root_r115_carry_22_) );
  XOR2X1 U335 ( .A(in_17bit_b[15]), .B(add_1_root_r115_carry_21_), .Y(
        add_1_root_r115_SUM_21_) );
  AND2X1 U336 ( .A(in_17bit_b[2]), .B(in_17bit_b[0]), .Y(
        add_1_root_r115_carry_7_) );
  XOR2X1 U337 ( .A(in_17bit_b[0]), .B(in_17bit_b[2]), .Y(
        add_1_root_r115_SUM_6_) );
  XOR2X1 U338 ( .A(n180), .B(sub_add_54_b0_carry[15]), .Y(N28) );
  AND2X1 U339 ( .A(sub_add_54_b0_carry[14]), .B(n179), .Y(
        sub_add_54_b0_carry[15]) );
  XOR2X1 U340 ( .A(n179), .B(sub_add_54_b0_carry[14]), .Y(N27) );
  AND2X1 U341 ( .A(sub_add_54_b0_carry[13]), .B(n178), .Y(
        sub_add_54_b0_carry[14]) );
  XOR2X1 U342 ( .A(n178), .B(sub_add_54_b0_carry[13]), .Y(N26) );
  AND2X1 U343 ( .A(sub_add_54_b0_carry[12]), .B(n177), .Y(
        sub_add_54_b0_carry[13]) );
  XOR2X1 U344 ( .A(n177), .B(sub_add_54_b0_carry[12]), .Y(N25) );
  AND2X1 U345 ( .A(sub_add_54_b0_carry[11]), .B(n176), .Y(
        sub_add_54_b0_carry[12]) );
  XOR2X1 U346 ( .A(n176), .B(sub_add_54_b0_carry[11]), .Y(N24) );
  AND2X1 U347 ( .A(sub_add_54_b0_carry[10]), .B(n175), .Y(
        sub_add_54_b0_carry[11]) );
  XOR2X1 U348 ( .A(n175), .B(sub_add_54_b0_carry[10]), .Y(N23) );
  AND2X1 U349 ( .A(sub_add_54_b0_carry[9]), .B(n174), .Y(
        sub_add_54_b0_carry[10]) );
  XOR2X1 U350 ( .A(n174), .B(sub_add_54_b0_carry[9]), .Y(N22) );
  AND2X1 U351 ( .A(sub_add_54_b0_carry[8]), .B(n173), .Y(
        sub_add_54_b0_carry[9]) );
  XOR2X1 U352 ( .A(n173), .B(sub_add_54_b0_carry[8]), .Y(N21) );
  AND2X1 U353 ( .A(sub_add_54_b0_carry[7]), .B(n172), .Y(
        sub_add_54_b0_carry[8]) );
  XOR2X1 U354 ( .A(n172), .B(sub_add_54_b0_carry[7]), .Y(N20) );
  AND2X1 U355 ( .A(sub_add_54_b0_carry[6]), .B(n171), .Y(
        sub_add_54_b0_carry[7]) );
  XOR2X1 U356 ( .A(n171), .B(sub_add_54_b0_carry[6]), .Y(N19) );
  AND2X1 U357 ( .A(sub_add_54_b0_carry[5]), .B(n170), .Y(
        sub_add_54_b0_carry[6]) );
  XOR2X1 U358 ( .A(n170), .B(sub_add_54_b0_carry[5]), .Y(N18) );
  AND2X1 U359 ( .A(sub_add_54_b0_carry[4]), .B(n164), .Y(
        sub_add_54_b0_carry[5]) );
  XOR2X1 U360 ( .A(n164), .B(sub_add_54_b0_carry[4]), .Y(N17) );
  AND2X1 U361 ( .A(sub_add_54_b0_carry[3]), .B(n163), .Y(
        sub_add_54_b0_carry[4]) );
  XOR2X1 U362 ( .A(n163), .B(sub_add_54_b0_carry[3]), .Y(N16) );
  AND2X1 U363 ( .A(sub_add_54_b0_carry[2]), .B(n160), .Y(
        sub_add_54_b0_carry[3]) );
  XOR2X1 U364 ( .A(n160), .B(sub_add_54_b0_carry[2]), .Y(N15) );
  AND2X1 U365 ( .A(n101), .B(n158), .Y(sub_add_54_b0_carry[2]) );
  XOR2X1 U366 ( .A(n158), .B(n101), .Y(N14) );
  XOR2X1 U367 ( .A(n19), .B(sub_add_75_b0_carry[16]), .Y(N481) );
  AND2X1 U368 ( .A(sub_add_75_b0_carry[15]), .B(n11), .Y(
        sub_add_75_b0_carry[16]) );
  XOR2X1 U369 ( .A(n11), .B(sub_add_75_b0_carry[15]), .Y(N480) );
  AND2X1 U370 ( .A(sub_add_75_b0_carry[14]), .B(n12), .Y(
        sub_add_75_b0_carry[15]) );
  XOR2X1 U371 ( .A(n12), .B(sub_add_75_b0_carry[14]), .Y(N479) );
  AND2X1 U372 ( .A(sub_add_75_b0_carry[13]), .B(n17), .Y(
        sub_add_75_b0_carry[14]) );
  AND2X1 U373 ( .A(sub_add_75_b0_carry[12]), .B(n16), .Y(
        sub_add_75_b0_carry[13]) );
  AND2X1 U374 ( .A(sub_add_75_b0_carry[11]), .B(n15), .Y(
        sub_add_75_b0_carry[12]) );
  AND2X1 U375 ( .A(sub_add_75_b0_carry[10]), .B(n14), .Y(
        sub_add_75_b0_carry[11]) );
  AND2X1 U376 ( .A(n30), .B(n8), .Y(sub_add_75_b0_carry[10]) );
  AND2X1 U377 ( .A(in_17bit_b[0]), .B(in_17bit_b[4]), .Y(
        add_1_root_r112_carry_5_) );
endmodule


module multi16_4_DW01_add_0 ( A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, 
        A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, 
        A_4_, B_23_, B_22_, B_21_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, 
        B_14_, B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, 
        SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, 
        SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, 
        SUM_7_ );
  input A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_,
         A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, B_23_, B_22_,
         B_21_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_,
         B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_;
  output SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_,
         SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_,
         SUM_8_, SUM_7_;
  wire   n1, n2, n3, n4;
  wire   [23:7] carry;

  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry[7]), .CO(carry[8]), .S(SUM_7_)
         );
  ADDFX2 U1_21 ( .A(A_21_), .B(B_21_), .CI(carry[21]), .CO(carry[22]), .S(
        SUM_21_) );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry[20]), .CO(carry[21]), .S(
        SUM_20_) );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry[19]), .CO(carry[20]), .S(
        SUM_19_) );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry[18]), .CO(carry[19]), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry[17]), .CO(carry[18]), .S(
        SUM_17_) );
  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry[16]), .CO(carry[17]), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry[15]), .CO(carry[16]), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry[14]), .CO(carry[15]), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry[13]), .CO(carry[14]), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry[12]), .CO(carry[13]), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry[11]), .CO(carry[12]), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry[10]), .CO(carry[11]), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry[9]), .CO(carry[10]), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry[8]), .CO(carry[9]), .S(SUM_8_)
         );
  ADDFX2 U1_22 ( .A(A_22_), .B(B_22_), .CI(carry[22]), .CO(carry[23]), .S(
        SUM_22_) );
  AND2X2 U1 ( .A(A_4_), .B(B_4_), .Y(n1) );
  XOR2X1 U2 ( .A(B_23_), .B(carry[23]), .Y(SUM_23_) );
  OAI2BB1X1 U3 ( .A0N(n2), .A1N(A_6_), .B0(n3), .Y(carry[7]) );
  OAI21XL U4 ( .A0(A_6_), .A1(n2), .B0(B_6_), .Y(n3) );
  OAI2BB1X1 U5 ( .A0N(n1), .A1N(A_5_), .B0(n4), .Y(n2) );
  OAI21XL U6 ( .A0(A_5_), .A1(n1), .B0(B_5_), .Y(n4) );
endmodule


module multi16_4_DW01_add_4 ( A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, 
        A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, 
        B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, 
        B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, SUM_22_, SUM_21_, SUM_20_, 
        SUM_19_, SUM_18_, SUM_17_, SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, 
        SUM_11_, SUM_10_, SUM_9_, SUM_8_, SUM_7_ );
  input A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_,
         A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, B_20_, B_19_,
         B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, B_10_, B_9_,
         B_8_, B_7_, B_6_, B_5_;
  output SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_,
         SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_,
         SUM_7_;
  wire   carry_21_, carry_20_, carry_19_, carry_18_, carry_17_, carry_16_,
         carry_15_, carry_14_, carry_13_, carry_12_, carry_11_, carry_10_,
         carry_9_, carry_8_, carry_7_, n1;

  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry_16_), .CO(carry_17_), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry_15_), .CO(carry_16_), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry_14_), .CO(carry_15_), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry_13_), .CO(carry_14_), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry_12_), .CO(carry_13_), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry_11_), .CO(carry_12_), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry_10_), .CO(carry_11_), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry_9_), .CO(carry_10_), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry_8_), .CO(carry_9_), .S(SUM_8_)
         );
  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry_7_), .CO(carry_8_), .S(SUM_7_)
         );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry_20_), .CO(carry_21_), .S(
        SUM_20_) );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry_19_), .CO(carry_20_), .S(
        SUM_19_) );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry_18_), .CO(carry_19_), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry_17_), .CO(carry_18_), .S(
        SUM_17_) );
  ADDFX2 U1_21 ( .A(A_21_), .B(B_21_), .CI(carry_21_), .CO(SUM_22_), .S(
        SUM_21_) );
  OAI2BB1X1 U1 ( .A0N(A_6_), .A1N(B_6_), .B0(n1), .Y(carry_7_) );
  OAI211X1 U2 ( .A0(B_6_), .A1(A_6_), .B0(A_5_), .C0(B_5_), .Y(n1) );
endmodule


module multi16_4_DW01_add_6 ( A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, 
        A_16_, A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, 
        A_6_, A_5_, A_4_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, 
        B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, 
        SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, 
        SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, 
        SUM_7_ );
  input A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_,
         A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, B_20_,
         B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, B_10_,
         B_9_, B_8_, B_7_, B_6_, B_5_, B_4_;
  output SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_,
         SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_,
         SUM_8_, SUM_7_;
  wire   n1, n2, n3, n4, n5, n6;
  wire   [21:7] carry;

  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry[7]), .CO(carry[8]), .S(SUM_7_)
         );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry[18]), .CO(carry[19]), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry[17]), .CO(carry[18]), .S(
        SUM_17_) );
  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry[16]), .CO(carry[17]), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry[15]), .CO(carry[16]), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry[14]), .CO(carry[15]), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry[13]), .CO(carry[14]), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry[12]), .CO(carry[13]), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry[11]), .CO(carry[12]), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry[10]), .CO(carry[11]), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry[9]), .CO(carry[10]), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry[8]), .CO(carry[9]), .S(SUM_8_)
         );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry[19]), .CO(carry[20]), .S(
        SUM_19_) );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry[20]), .CO(carry[21]), .S(
        SUM_20_) );
  AND2X2 U1 ( .A(A_22_), .B(n2), .Y(n1) );
  AND2X2 U2 ( .A(A_21_), .B(carry[21]), .Y(n2) );
  XOR2X1 U3 ( .A(A_23_), .B(n1), .Y(SUM_23_) );
  XOR2X1 U4 ( .A(A_21_), .B(carry[21]), .Y(SUM_21_) );
  XOR2X1 U5 ( .A(A_22_), .B(n2), .Y(SUM_22_) );
  AND2X2 U6 ( .A(A_4_), .B(B_4_), .Y(n3) );
  OAI2BB1X1 U7 ( .A0N(n4), .A1N(A_6_), .B0(n5), .Y(carry[7]) );
  OAI21XL U8 ( .A0(A_6_), .A1(n4), .B0(B_6_), .Y(n5) );
  OAI2BB1X1 U9 ( .A0N(n3), .A1N(A_5_), .B0(n6), .Y(n4) );
  OAI21XL U10 ( .A0(A_5_), .A1(n3), .B0(B_5_), .Y(n6) );
endmodule


module multi16_4 ( in_17bit, in_8bit, out );
  input [16:0] in_17bit;
  input [7:0] in_8bit;
  output [16:0] out;
  wire   n257, n258, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24,
         N25, N26, N27, N28, N29, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, N205, N206,
         N207, N208, N209, N210, N211, N212, N213, N214, N215, N216, N217,
         N218, N219, N220, N221, N347, N348, N349, N350, N351, N352, N353,
         N354, N355, N356, N357, N358, N359, N360, N361, N362, N363, N446,
         N447, N448, N449, N450, N451, N452, N453, N454, N455, N456, N457,
         N458, N459, N460, N461, N462, N463, N476, N477, N478, N479, N480,
         add_2_root_r119_carry_10_, add_2_root_r119_carry_11_,
         add_2_root_r119_carry_12_, add_2_root_r119_carry_13_,
         add_2_root_r119_carry_14_, add_2_root_r119_carry_15_,
         add_2_root_r119_carry_16_, add_2_root_r119_carry_17_,
         add_2_root_r119_carry_18_, add_2_root_r119_carry_19_,
         add_2_root_r119_carry_20_, add_2_root_r119_carry_21_,
         add_2_root_r119_carry_6_, add_2_root_r119_carry_7_,
         add_2_root_r119_carry_8_, add_2_root_r119_carry_9_,
         add_2_root_r119_SUM_5_, add_2_root_r119_SUM_6_,
         add_2_root_r119_SUM_7_, add_2_root_r119_SUM_8_,
         add_2_root_r119_SUM_9_, add_2_root_r119_SUM_10_,
         add_2_root_r119_SUM_11_, add_2_root_r119_SUM_12_,
         add_2_root_r119_SUM_13_, add_2_root_r119_SUM_14_,
         add_2_root_r119_SUM_15_, add_2_root_r119_SUM_16_,
         add_2_root_r119_SUM_17_, add_2_root_r119_SUM_18_,
         add_2_root_r119_SUM_19_, add_2_root_r119_SUM_20_,
         add_2_root_r119_SUM_21_, add_2_root_r119_SUM_22_,
         add_1_root_r119_SUM_6_, add_1_root_r119_SUM_7_,
         add_1_root_r119_SUM_8_, add_1_root_r119_SUM_9_,
         add_1_root_r119_SUM_10_, add_1_root_r119_SUM_11_,
         add_1_root_r119_SUM_12_, add_1_root_r119_SUM_13_,
         add_1_root_r119_SUM_14_, add_1_root_r119_SUM_15_,
         add_1_root_r119_SUM_16_, add_1_root_r119_SUM_17_,
         add_1_root_r119_SUM_18_, add_1_root_r119_SUM_19_,
         add_1_root_r119_SUM_20_, add_1_root_r119_SUM_21_,
         add_1_root_r119_SUM_22_, add_1_root_r119_SUM_23_,
         add_1_root_r119_A_2_, add_1_root_r119_A_3_, add_1_root_r119_A_4_,
         add_1_root_r119_A_5_, add_1_root_r119_A_6_, add_1_root_r119_A_7_,
         add_1_root_r119_A_8_, add_1_root_r119_A_9_, add_1_root_r119_A_10_,
         add_1_root_r119_A_11_, add_1_root_r119_A_12_, add_1_root_r119_A_13_,
         add_1_root_r119_A_14_, add_1_root_r119_A_15_, add_1_root_r119_A_16_,
         add_1_root_r119_A_17_, add_1_root_r119_A_18_, add_1_root_r119_A_19_,
         add_3_root_r119_carry_10_, add_3_root_r119_carry_11_,
         add_3_root_r119_carry_12_, add_3_root_r119_carry_13_,
         add_3_root_r119_carry_14_, add_3_root_r119_carry_15_,
         add_3_root_r119_carry_16_, add_3_root_r119_carry_17_,
         add_3_root_r119_carry_18_, add_3_root_r119_carry_3_,
         add_3_root_r119_carry_4_, add_3_root_r119_carry_5_,
         add_3_root_r119_carry_6_, add_3_root_r119_carry_7_,
         add_3_root_r119_carry_8_, add_3_root_r119_carry_9_,
         add_1_root_r112_carry_10_, add_1_root_r112_carry_11_,
         add_1_root_r112_carry_12_, add_1_root_r112_carry_13_,
         add_1_root_r112_carry_14_, add_1_root_r112_carry_15_,
         add_1_root_r112_carry_16_, add_1_root_r112_carry_17_,
         add_1_root_r112_carry_18_, add_1_root_r112_carry_19_,
         add_1_root_r112_carry_20_, add_1_root_r112_carry_5_,
         add_1_root_r112_carry_6_, add_1_root_r112_carry_7_,
         add_1_root_r112_carry_8_, add_1_root_r112_carry_9_,
         add_1_root_r112_SUM_1_, add_1_root_r112_SUM_2_,
         add_1_root_r112_SUM_3_, add_1_root_r112_SUM_4_,
         add_1_root_r112_SUM_5_, add_1_root_r112_SUM_6_,
         add_1_root_r112_SUM_7_, add_1_root_r112_SUM_8_,
         add_1_root_r112_SUM_9_, add_1_root_r112_SUM_10_,
         add_1_root_r112_SUM_11_, add_1_root_r112_SUM_12_,
         add_1_root_r112_SUM_13_, add_1_root_r112_SUM_14_,
         add_1_root_r112_SUM_15_, add_1_root_r112_SUM_16_,
         add_1_root_r112_SUM_17_, add_1_root_r112_SUM_18_,
         add_1_root_r112_SUM_19_, add_1_root_r112_SUM_20_,
         add_1_root_r112_SUM_21_, add_2_root_r115_carry_10_,
         add_2_root_r115_carry_11_, add_2_root_r115_carry_12_,
         add_2_root_r115_carry_13_, add_2_root_r115_carry_14_,
         add_2_root_r115_carry_15_, add_2_root_r115_carry_16_,
         add_2_root_r115_carry_17_, add_2_root_r115_carry_18_,
         add_2_root_r115_carry_19_, add_2_root_r115_carry_4_,
         add_2_root_r115_carry_5_, add_2_root_r115_carry_6_,
         add_2_root_r115_carry_7_, add_2_root_r115_carry_8_,
         add_2_root_r115_carry_9_, add_2_root_r115_SUM_3_,
         add_2_root_r115_SUM_4_, add_2_root_r115_SUM_5_,
         add_2_root_r115_SUM_6_, add_2_root_r115_SUM_7_,
         add_2_root_r115_SUM_8_, add_2_root_r115_SUM_9_,
         add_2_root_r115_SUM_10_, add_2_root_r115_SUM_11_,
         add_2_root_r115_SUM_12_, add_2_root_r115_SUM_13_,
         add_2_root_r115_SUM_14_, add_2_root_r115_SUM_15_,
         add_2_root_r115_SUM_16_, add_2_root_r115_SUM_17_,
         add_2_root_r115_SUM_18_, add_2_root_r115_SUM_19_,
         add_2_root_r115_SUM_20_, add_1_root_r115_carry_10_,
         add_1_root_r115_carry_11_, add_1_root_r115_carry_12_,
         add_1_root_r115_carry_13_, add_1_root_r115_carry_14_,
         add_1_root_r115_carry_15_, add_1_root_r115_carry_16_,
         add_1_root_r115_carry_17_, add_1_root_r115_carry_18_,
         add_1_root_r115_carry_19_, add_1_root_r115_carry_20_,
         add_1_root_r115_carry_21_, add_1_root_r115_carry_22_,
         add_1_root_r115_carry_7_, add_1_root_r115_carry_8_,
         add_1_root_r115_carry_9_, add_1_root_r115_SUM_6_,
         add_1_root_r115_SUM_7_, add_1_root_r115_SUM_8_,
         add_1_root_r115_SUM_9_, add_1_root_r115_SUM_10_,
         add_1_root_r115_SUM_11_, add_1_root_r115_SUM_12_,
         add_1_root_r115_SUM_13_, add_1_root_r115_SUM_14_,
         add_1_root_r115_SUM_15_, add_1_root_r115_SUM_16_,
         add_1_root_r115_SUM_17_, add_1_root_r115_SUM_18_,
         add_1_root_r115_SUM_19_, add_1_root_r115_SUM_20_,
         add_1_root_r115_SUM_21_, add_1_root_r115_SUM_22_,
         add_1_root_r115_SUM_23_, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n158, n160, n163, n164, n167, n168, n170, n171,
         n172, n173, n174, n175, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256;
  wire   [16:0] in_17bit_b;
  wire   [23:8] neg_mul;
  wire   [15:10] sub_add_75_b0_carry;
  wire   [15:2] sub_add_54_b0_carry;
  wire   [22:7] add_1_root_r119_carry;

  multi16_4_DW01_add_0 add_0_root_r119 ( .A_22_(add_2_root_r119_SUM_22_), 
        .A_21_(add_2_root_r119_SUM_21_), .A_20_(add_2_root_r119_SUM_20_), 
        .A_19_(add_2_root_r119_SUM_19_), .A_18_(add_2_root_r119_SUM_18_), 
        .A_17_(add_2_root_r119_SUM_17_), .A_16_(add_2_root_r119_SUM_16_), 
        .A_15_(add_2_root_r119_SUM_15_), .A_14_(add_2_root_r119_SUM_14_), 
        .A_13_(add_2_root_r119_SUM_13_), .A_12_(add_2_root_r119_SUM_12_), 
        .A_11_(add_2_root_r119_SUM_11_), .A_10_(add_2_root_r119_SUM_10_), 
        .A_9_(add_2_root_r119_SUM_9_), .A_8_(add_2_root_r119_SUM_8_), .A_7_(
        add_2_root_r119_SUM_7_), .A_6_(add_2_root_r119_SUM_6_), .A_5_(
        add_2_root_r119_SUM_5_), .A_4_(in_17bit_b[0]), .B_23_(
        add_1_root_r119_SUM_23_), .B_22_(add_1_root_r119_SUM_22_), .B_21_(
        add_1_root_r119_SUM_21_), .B_20_(add_1_root_r119_SUM_20_), .B_19_(
        add_1_root_r119_SUM_19_), .B_18_(add_1_root_r119_SUM_18_), .B_17_(
        add_1_root_r119_SUM_17_), .B_16_(add_1_root_r119_SUM_16_), .B_15_(
        add_1_root_r119_SUM_15_), .B_14_(add_1_root_r119_SUM_14_), .B_13_(
        add_1_root_r119_SUM_13_), .B_12_(add_1_root_r119_SUM_12_), .B_11_(
        add_1_root_r119_SUM_11_), .B_10_(add_1_root_r119_SUM_10_), .B_9_(
        add_1_root_r119_SUM_9_), .B_8_(add_1_root_r119_SUM_8_), .B_7_(
        add_1_root_r119_SUM_7_), .B_6_(add_1_root_r119_SUM_6_), .B_5_(
        add_1_root_r119_A_5_), .B_4_(add_1_root_r119_A_4_), .SUM_23_(N363), 
        .SUM_22_(N362), .SUM_21_(N361), .SUM_20_(N360), .SUM_19_(N359), 
        .SUM_18_(N358), .SUM_17_(N357), .SUM_16_(N356), .SUM_15_(N355), 
        .SUM_14_(N354), .SUM_13_(N353), .SUM_12_(N352), .SUM_11_(N351), 
        .SUM_10_(N350), .SUM_9_(N349), .SUM_8_(N348), .SUM_7_(N347) );
  multi16_4_DW01_add_4 add_0_root_r112 ( .A_21_(n44), .A_20_(in_17bit_b[15]), 
        .A_19_(in_17bit_b[14]), .A_18_(in_17bit_b[13]), .A_17_(in_17bit_b[12]), 
        .A_16_(in_17bit_b[11]), .A_15_(in_17bit_b[10]), .A_14_(in_17bit_b[9]), 
        .A_13_(in_17bit_b[8]), .A_12_(in_17bit_b[7]), .A_11_(in_17bit_b[6]), 
        .A_10_(in_17bit_b[5]), .A_9_(in_17bit_b[4]), .A_8_(in_17bit_b[3]), 
        .A_7_(in_17bit_b[2]), .A_6_(in_17bit_b[1]), .A_5_(in_17bit_b[0]), 
        .B_21_(add_1_root_r112_SUM_21_), .B_20_(add_1_root_r112_SUM_20_), 
        .B_19_(add_1_root_r112_SUM_19_), .B_18_(add_1_root_r112_SUM_18_), 
        .B_17_(add_1_root_r112_SUM_17_), .B_16_(add_1_root_r112_SUM_16_), 
        .B_15_(add_1_root_r112_SUM_15_), .B_14_(add_1_root_r112_SUM_14_), 
        .B_13_(add_1_root_r112_SUM_13_), .B_12_(add_1_root_r112_SUM_12_), 
        .B_11_(add_1_root_r112_SUM_11_), .B_10_(add_1_root_r112_SUM_10_), 
        .B_9_(add_1_root_r112_SUM_9_), .B_8_(add_1_root_r112_SUM_8_), .B_7_(
        add_1_root_r112_SUM_7_), .B_6_(add_1_root_r112_SUM_6_), .B_5_(
        add_1_root_r112_SUM_5_), .SUM_22_(N123), .SUM_21_(N122), .SUM_20_(N121), .SUM_19_(N120), .SUM_18_(N119), .SUM_17_(N118), .SUM_16_(N117), .SUM_15_(
        N116), .SUM_14_(N115), .SUM_13_(N114), .SUM_12_(N113), .SUM_11_(N112), 
        .SUM_10_(N111), .SUM_9_(N110), .SUM_8_(N109), .SUM_7_(N108) );
  multi16_4_DW01_add_6 add_0_root_r115 ( .A_23_(add_1_root_r115_SUM_23_), 
        .A_22_(add_1_root_r115_SUM_22_), .A_21_(add_1_root_r115_SUM_21_), 
        .A_20_(add_1_root_r115_SUM_20_), .A_19_(add_1_root_r115_SUM_19_), 
        .A_18_(add_1_root_r115_SUM_18_), .A_17_(add_1_root_r115_SUM_17_), 
        .A_16_(add_1_root_r115_SUM_16_), .A_15_(add_1_root_r115_SUM_15_), 
        .A_14_(add_1_root_r115_SUM_14_), .A_13_(add_1_root_r115_SUM_13_), 
        .A_12_(add_1_root_r115_SUM_12_), .A_11_(add_1_root_r115_SUM_11_), 
        .A_10_(add_1_root_r115_SUM_10_), .A_9_(add_1_root_r115_SUM_9_), .A_8_(
        add_1_root_r115_SUM_8_), .A_7_(add_1_root_r115_SUM_7_), .A_6_(
        add_1_root_r115_SUM_6_), .A_5_(in_17bit_b[1]), .A_4_(in_17bit_b[0]), 
        .B_20_(add_2_root_r115_SUM_20_), .B_19_(add_2_root_r115_SUM_19_), 
        .B_18_(add_2_root_r115_SUM_18_), .B_17_(add_2_root_r115_SUM_17_), 
        .B_16_(add_2_root_r115_SUM_16_), .B_15_(add_2_root_r115_SUM_15_), 
        .B_14_(add_2_root_r115_SUM_14_), .B_13_(add_2_root_r115_SUM_13_), 
        .B_12_(add_2_root_r115_SUM_12_), .B_11_(add_2_root_r115_SUM_11_), 
        .B_10_(add_2_root_r115_SUM_10_), .B_9_(add_2_root_r115_SUM_9_), .B_8_(
        add_2_root_r115_SUM_8_), .B_7_(add_2_root_r115_SUM_7_), .B_6_(
        add_2_root_r115_SUM_6_), .B_5_(add_2_root_r115_SUM_5_), .B_4_(
        add_2_root_r115_SUM_4_), .SUM_23_(N221), .SUM_22_(N220), .SUM_21_(N219), .SUM_20_(N218), .SUM_19_(N217), .SUM_18_(N216), .SUM_17_(N215), .SUM_16_(
        N214), .SUM_15_(N213), .SUM_14_(N212), .SUM_13_(N211), .SUM_12_(N210), 
        .SUM_11_(N209), .SUM_10_(N208), .SUM_9_(N207), .SUM_8_(N206), .SUM_7_(
        N205) );
  TLATX1 neg_mul_reg_16_ ( .G(N446), .D(N456), .QN(n9) );
  TLATX1 neg_mul_reg_15_ ( .G(N446), .D(N455), .QN(n8) );
  TLATX1 neg_mul_reg_14_ ( .G(N446), .D(N454), .Q(neg_mul[14]), .QN(n2) );
  TLATX1 neg_mul_reg_13_ ( .G(N446), .D(N453), .QN(n7) );
  TLATX1 neg_mul_reg_12_ ( .G(N446), .D(N452), .QN(n6) );
  TLATX1 neg_mul_reg_11_ ( .G(N446), .D(N451), .QN(n5) );
  TLATX1 neg_mul_reg_9_ ( .G(N446), .D(N449), .QN(n4) );
  TLATX1 neg_mul_reg_23_ ( .G(N446), .D(N463), .Q(neg_mul[23]), .QN(n3) );
  TLATX1 neg_mul_reg_22_ ( .G(N446), .D(N462), .Q(neg_mul[22]), .QN(n10) );
  TLATX1 neg_mul_reg_21_ ( .G(N446), .D(N461), .Q(neg_mul[21]), .QN(n14) );
  TLATX1 neg_mul_reg_20_ ( .G(N446), .D(N460), .Q(neg_mul[20]), .QN(n12) );
  TLATX1 neg_mul_reg_19_ ( .G(N446), .D(N459), .Q(neg_mul[19]), .QN(n13) );
  TLATX1 neg_mul_reg_18_ ( .G(N446), .D(N458), .Q(neg_mul[18]), .QN(n11) );
  TLATX1 neg_mul_reg_17_ ( .G(N446), .D(N457), .QN(n16) );
  TLATX1 neg_mul_reg_10_ ( .G(N446), .D(N450), .Q(neg_mul[10]), .QN(n15) );
  TLATX1 neg_mul_reg_8_ ( .G(N446), .D(N448), .Q(neg_mul[8]), .QN(n17) );
  TLATX1 neg_mul_reg_7_ ( .G(N446), .D(N447), .Q(out[0]) );
  CLKINVX8 U2 ( .A(n19), .Y(out[1]) );
  BUFX8 U3 ( .A(n257), .Y(out[13]) );
  MX2X2 U4 ( .A(N478), .B(neg_mul[20]), .S0(n81), .Y(n257) );
  NAND2X2 U5 ( .A(n43), .B(n17), .Y(n58) );
  XNOR2X4 U6 ( .A(n40), .B(n43), .Y(n81) );
  MX2X2 U7 ( .A(neg_mul[18]), .B(N476), .S0(n82), .Y(out[11]) );
  INVX1 U8 ( .A(n92), .Y(n88) );
  BUFX8 U9 ( .A(in_8bit[7]), .Y(n43) );
  INVXL U10 ( .A(n39), .Y(n54) );
  XNOR2X1 U11 ( .A(neg_mul[23]), .B(n37), .Y(n18) );
  CLKINVX8 U12 ( .A(in_17bit[16]), .Y(n51) );
  CLKINVX8 U13 ( .A(in_17bit[16]), .Y(n50) );
  NOR2X4 U14 ( .A(n36), .B(n64), .Y(n65) );
  INVXL U15 ( .A(n49), .Y(n56) );
  INVXL U16 ( .A(n49), .Y(n55) );
  INVX8 U17 ( .A(n50), .Y(n39) );
  AOI2BB2X1 U18 ( .B0(n69), .B1(n43), .A0N(n43), .A1N(neg_mul[10]), .Y(n70) );
  INVX8 U19 ( .A(n81), .Y(n82) );
  MX2X2 U20 ( .A(neg_mul[19]), .B(N477), .S0(n82), .Y(out[12]) );
  XNOR2X2 U21 ( .A(n53), .B(n43), .Y(n73) );
  NOR2X4 U22 ( .A(n30), .B(n78), .Y(n24) );
  NOR2X4 U23 ( .A(n74), .B(n78), .Y(n75) );
  XNOR2X4 U24 ( .A(n39), .B(n43), .Y(n64) );
  INVX8 U25 ( .A(n51), .Y(n53) );
  INVX4 U26 ( .A(n258), .Y(n19) );
  AOI211X2 U27 ( .A0(n40), .A1(n63), .B0(n62), .C0(n36), .Y(n258) );
  NOR2X2 U28 ( .A(n39), .B(n61), .Y(n62) );
  INVX8 U29 ( .A(n51), .Y(n40) );
  XOR2X4 U30 ( .A(n27), .B(n9), .Y(out[9]) );
  OR2X4 U31 ( .A(n34), .B(n80), .Y(n27) );
  XNOR2X4 U32 ( .A(n53), .B(n43), .Y(n78) );
  NAND2X2 U33 ( .A(n24), .B(n2), .Y(n22) );
  NAND2X4 U34 ( .A(n21), .B(neg_mul[14]), .Y(n23) );
  NAND2X4 U35 ( .A(n22), .B(n23), .Y(out[7]) );
  CLKINVX4 U36 ( .A(n24), .Y(n21) );
  AND3X1 U37 ( .A(in_8bit[2]), .B(n48), .C(n47), .Y(n33) );
  INVX1 U38 ( .A(n206), .Y(in_17bit_b[1]) );
  INVX1 U39 ( .A(n245), .Y(in_17bit_b[14]) );
  INVX1 U40 ( .A(n242), .Y(in_17bit_b[13]) );
  INVX1 U41 ( .A(n209), .Y(in_17bit_b[2]) );
  INVX1 U42 ( .A(n218), .Y(in_17bit_b[5]) );
  INVX1 U43 ( .A(n221), .Y(in_17bit_b[6]) );
  INVX1 U44 ( .A(n224), .Y(in_17bit_b[7]) );
  INVX1 U45 ( .A(n227), .Y(in_17bit_b[8]) );
  INVX1 U46 ( .A(n230), .Y(in_17bit_b[9]) );
  INVX1 U47 ( .A(n233), .Y(in_17bit_b[10]) );
  INVX1 U48 ( .A(n236), .Y(in_17bit_b[11]) );
  INVX1 U49 ( .A(n239), .Y(in_17bit_b[12]) );
  INVX1 U50 ( .A(n215), .Y(in_17bit_b[4]) );
  INVX1 U51 ( .A(n212), .Y(in_17bit_b[3]) );
  NAND2XL U52 ( .A(n43), .B(n15), .Y(n67) );
  INVX1 U53 ( .A(n56), .Y(n52) );
  OAI21XL U54 ( .A0(n255), .A1(n256), .B0(n254), .Y(N463) );
  AOI22X1 U55 ( .A0(N221), .A1(n42), .B0(N363), .B1(n41), .Y(n254) );
  INVX1 U56 ( .A(n174), .Y(n255) );
  NAND3BX1 U57 ( .AN(n47), .B(n45), .C(n43), .Y(n91) );
  ADDFX2 U58 ( .A(n44), .B(in_17bit_b[12]), .CI(add_1_root_r112_carry_16_), 
        .CO(add_1_root_r112_carry_17_), .S(add_1_root_r112_SUM_16_) );
  ADDFX2 U59 ( .A(add_1_root_r119_A_19_), .B(in_17bit_b[13]), .CI(
        add_1_root_r119_carry[19]), .CO(add_1_root_r119_carry[20]), .S(
        add_1_root_r119_SUM_19_) );
  ADDFX2 U60 ( .A(n44), .B(in_17bit_b[15]), .CI(add_3_root_r119_carry_17_), 
        .CO(add_3_root_r119_carry_18_), .S(add_1_root_r119_A_17_) );
  ADDFX2 U61 ( .A(n44), .B(in_17bit_b[14]), .CI(add_2_root_r115_carry_17_), 
        .CO(add_2_root_r115_carry_18_), .S(add_2_root_r115_SUM_17_) );
  ADDFX2 U62 ( .A(n44), .B(in_17bit_b[14]), .CI(add_1_root_r115_carry_20_), 
        .CO(add_1_root_r115_carry_21_), .S(add_1_root_r115_SUM_20_) );
  ADDFX2 U63 ( .A(n44), .B(in_17bit_b[15]), .CI(add_2_root_r119_carry_20_), 
        .CO(add_2_root_r119_carry_21_), .S(add_2_root_r119_SUM_20_) );
  ADDFX2 U64 ( .A(in_17bit_b[3]), .B(in_17bit_b[1]), .CI(
        add_2_root_r115_carry_4_), .CO(add_2_root_r115_carry_5_), .S(
        add_2_root_r115_SUM_4_) );
  ADDFX2 U65 ( .A(in_17bit_b[4]), .B(in_17bit_b[2]), .CI(
        add_2_root_r115_carry_5_), .CO(add_2_root_r115_carry_6_), .S(
        add_2_root_r115_SUM_5_) );
  ADDFX2 U66 ( .A(in_17bit_b[5]), .B(in_17bit_b[1]), .CI(
        add_1_root_r112_carry_5_), .CO(add_1_root_r112_carry_6_), .S(
        add_1_root_r112_SUM_5_) );
  ADDFX2 U67 ( .A(in_17bit_b[6]), .B(in_17bit_b[5]), .CI(
        add_3_root_r119_carry_7_), .CO(add_3_root_r119_carry_8_), .S(
        add_1_root_r119_A_7_) );
  ADDFX2 U68 ( .A(in_17bit_b[6]), .B(in_17bit_b[2]), .CI(
        add_1_root_r112_carry_6_), .CO(add_1_root_r112_carry_7_), .S(
        add_1_root_r112_SUM_6_) );
  ADDFX2 U69 ( .A(in_17bit_b[3]), .B(in_17bit_b[1]), .CI(
        add_1_root_r115_carry_7_), .CO(add_1_root_r115_carry_8_), .S(
        add_1_root_r115_SUM_7_) );
  ADDFX2 U70 ( .A(in_17bit_b[7]), .B(in_17bit_b[6]), .CI(
        add_3_root_r119_carry_8_), .CO(add_3_root_r119_carry_9_), .S(
        add_1_root_r119_A_8_) );
  ADDFX2 U71 ( .A(add_1_root_r119_A_7_), .B(in_17bit_b[1]), .CI(
        add_1_root_r119_carry[7]), .CO(add_1_root_r119_carry[8]), .S(
        add_1_root_r119_SUM_7_) );
  ADDFX2 U72 ( .A(in_17bit_b[2]), .B(in_17bit_b[1]), .CI(
        add_2_root_r119_carry_6_), .CO(add_2_root_r119_carry_7_), .S(
        add_2_root_r119_SUM_6_) );
  ADDFX2 U73 ( .A(in_17bit_b[4]), .B(in_17bit_b[2]), .CI(
        add_1_root_r115_carry_8_), .CO(add_1_root_r115_carry_9_), .S(
        add_1_root_r115_SUM_8_) );
  ADDFX2 U74 ( .A(in_17bit_b[8]), .B(in_17bit_b[7]), .CI(
        add_3_root_r119_carry_9_), .CO(add_3_root_r119_carry_10_), .S(
        add_1_root_r119_A_9_) );
  ADDFX2 U75 ( .A(add_1_root_r119_A_8_), .B(in_17bit_b[2]), .CI(
        add_1_root_r119_carry[8]), .CO(add_1_root_r119_carry[9]), .S(
        add_1_root_r119_SUM_8_) );
  ADDFX2 U76 ( .A(in_17bit_b[3]), .B(in_17bit_b[2]), .CI(
        add_2_root_r119_carry_7_), .CO(add_2_root_r119_carry_8_), .S(
        add_2_root_r119_SUM_7_) );
  ADDFX2 U77 ( .A(in_17bit_b[6]), .B(in_17bit_b[4]), .CI(
        add_2_root_r115_carry_7_), .CO(add_2_root_r115_carry_8_), .S(
        add_2_root_r115_SUM_7_) );
  ADDFX2 U78 ( .A(in_17bit_b[8]), .B(in_17bit_b[4]), .CI(
        add_1_root_r112_carry_8_), .CO(add_1_root_r112_carry_9_), .S(
        add_1_root_r112_SUM_8_) );
  ADDFX2 U79 ( .A(in_17bit_b[9]), .B(in_17bit_b[8]), .CI(
        add_3_root_r119_carry_10_), .CO(add_3_root_r119_carry_11_), .S(
        add_1_root_r119_A_10_) );
  ADDFX2 U80 ( .A(in_17bit_b[6]), .B(in_17bit_b[4]), .CI(
        add_1_root_r115_carry_10_), .CO(add_1_root_r115_carry_11_), .S(
        add_1_root_r115_SUM_10_) );
  ADDFX2 U81 ( .A(in_17bit_b[10]), .B(in_17bit_b[9]), .CI(
        add_3_root_r119_carry_11_), .CO(add_3_root_r119_carry_12_), .S(
        add_1_root_r119_A_11_) );
  ADDFX2 U82 ( .A(in_17bit_b[7]), .B(in_17bit_b[5]), .CI(
        add_2_root_r115_carry_8_), .CO(add_2_root_r115_carry_9_), .S(
        add_2_root_r115_SUM_8_) );
  ADDFX2 U83 ( .A(in_17bit_b[9]), .B(in_17bit_b[5]), .CI(
        add_1_root_r112_carry_9_), .CO(add_1_root_r112_carry_10_), .S(
        add_1_root_r112_SUM_9_) );
  ADDFX2 U84 ( .A(add_1_root_r119_A_10_), .B(in_17bit_b[4]), .CI(
        add_1_root_r119_carry[10]), .CO(add_1_root_r119_carry[11]), .S(
        add_1_root_r119_SUM_10_) );
  ADDFX2 U85 ( .A(in_17bit_b[5]), .B(in_17bit_b[4]), .CI(
        add_2_root_r119_carry_9_), .CO(add_2_root_r119_carry_10_), .S(
        add_2_root_r119_SUM_9_) );
  ADDFX2 U86 ( .A(in_17bit_b[8]), .B(in_17bit_b[6]), .CI(
        add_2_root_r115_carry_9_), .CO(add_2_root_r115_carry_10_), .S(
        add_2_root_r115_SUM_9_) );
  ADDFX2 U87 ( .A(in_17bit_b[10]), .B(in_17bit_b[6]), .CI(
        add_1_root_r112_carry_10_), .CO(add_1_root_r112_carry_11_), .S(
        add_1_root_r112_SUM_10_) );
  ADDFX2 U88 ( .A(in_17bit_b[7]), .B(in_17bit_b[5]), .CI(
        add_1_root_r115_carry_11_), .CO(add_1_root_r115_carry_12_), .S(
        add_1_root_r115_SUM_11_) );
  ADDFX2 U89 ( .A(in_17bit_b[11]), .B(in_17bit_b[10]), .CI(
        add_3_root_r119_carry_12_), .CO(add_3_root_r119_carry_13_), .S(
        add_1_root_r119_A_12_) );
  ADDFX2 U90 ( .A(add_1_root_r119_A_11_), .B(in_17bit_b[5]), .CI(
        add_1_root_r119_carry[11]), .CO(add_1_root_r119_carry[12]), .S(
        add_1_root_r119_SUM_11_) );
  ADDFX2 U91 ( .A(in_17bit_b[6]), .B(in_17bit_b[5]), .CI(
        add_2_root_r119_carry_10_), .CO(add_2_root_r119_carry_11_), .S(
        add_2_root_r119_SUM_10_) );
  ADDFX2 U92 ( .A(in_17bit_b[9]), .B(in_17bit_b[7]), .CI(
        add_2_root_r115_carry_10_), .CO(add_2_root_r115_carry_11_), .S(
        add_2_root_r115_SUM_10_) );
  ADDFX2 U93 ( .A(in_17bit_b[11]), .B(in_17bit_b[7]), .CI(
        add_1_root_r112_carry_11_), .CO(add_1_root_r112_carry_12_), .S(
        add_1_root_r112_SUM_11_) );
  ADDFX2 U94 ( .A(in_17bit_b[8]), .B(in_17bit_b[6]), .CI(
        add_1_root_r115_carry_12_), .CO(add_1_root_r115_carry_13_), .S(
        add_1_root_r115_SUM_12_) );
  ADDFX2 U95 ( .A(in_17bit_b[12]), .B(in_17bit_b[11]), .CI(
        add_3_root_r119_carry_13_), .CO(add_3_root_r119_carry_14_), .S(
        add_1_root_r119_A_13_) );
  ADDFX2 U96 ( .A(add_1_root_r119_A_12_), .B(in_17bit_b[6]), .CI(
        add_1_root_r119_carry[12]), .CO(add_1_root_r119_carry[13]), .S(
        add_1_root_r119_SUM_12_) );
  ADDFX2 U97 ( .A(in_17bit_b[7]), .B(in_17bit_b[6]), .CI(
        add_2_root_r119_carry_11_), .CO(add_2_root_r119_carry_12_), .S(
        add_2_root_r119_SUM_11_) );
  ADDFX2 U98 ( .A(in_17bit_b[10]), .B(in_17bit_b[8]), .CI(
        add_2_root_r115_carry_11_), .CO(add_2_root_r115_carry_12_), .S(
        add_2_root_r115_SUM_11_) );
  ADDFX2 U99 ( .A(in_17bit_b[12]), .B(in_17bit_b[8]), .CI(
        add_1_root_r112_carry_12_), .CO(add_1_root_r112_carry_13_), .S(
        add_1_root_r112_SUM_12_) );
  ADDFX2 U100 ( .A(in_17bit_b[9]), .B(in_17bit_b[7]), .CI(
        add_1_root_r115_carry_13_), .CO(add_1_root_r115_carry_14_), .S(
        add_1_root_r115_SUM_13_) );
  ADDFX2 U101 ( .A(in_17bit_b[13]), .B(in_17bit_b[12]), .CI(
        add_3_root_r119_carry_14_), .CO(add_3_root_r119_carry_15_), .S(
        add_1_root_r119_A_14_) );
  ADDFX2 U102 ( .A(add_1_root_r119_A_13_), .B(in_17bit_b[7]), .CI(
        add_1_root_r119_carry[13]), .CO(add_1_root_r119_carry[14]), .S(
        add_1_root_r119_SUM_13_) );
  ADDFX2 U103 ( .A(in_17bit_b[8]), .B(in_17bit_b[7]), .CI(
        add_2_root_r119_carry_12_), .CO(add_2_root_r119_carry_13_), .S(
        add_2_root_r119_SUM_12_) );
  ADDFX2 U104 ( .A(in_17bit_b[11]), .B(in_17bit_b[9]), .CI(
        add_2_root_r115_carry_12_), .CO(add_2_root_r115_carry_13_), .S(
        add_2_root_r115_SUM_12_) );
  ADDFX2 U105 ( .A(in_17bit_b[13]), .B(in_17bit_b[9]), .CI(
        add_1_root_r112_carry_13_), .CO(add_1_root_r112_carry_14_), .S(
        add_1_root_r112_SUM_13_) );
  ADDFX2 U106 ( .A(in_17bit_b[10]), .B(in_17bit_b[8]), .CI(
        add_1_root_r115_carry_14_), .CO(add_1_root_r115_carry_15_), .S(
        add_1_root_r115_SUM_14_) );
  ADDFX2 U107 ( .A(in_17bit_b[14]), .B(in_17bit_b[13]), .CI(
        add_3_root_r119_carry_15_), .CO(add_3_root_r119_carry_16_), .S(
        add_1_root_r119_A_15_) );
  ADDFX2 U108 ( .A(add_1_root_r119_A_14_), .B(in_17bit_b[8]), .CI(
        add_1_root_r119_carry[14]), .CO(add_1_root_r119_carry[15]), .S(
        add_1_root_r119_SUM_14_) );
  ADDFX2 U109 ( .A(in_17bit_b[3]), .B(in_17bit_b[2]), .CI(
        add_3_root_r119_carry_4_), .CO(add_3_root_r119_carry_5_), .S(
        add_1_root_r119_A_4_) );
  ADDFX2 U110 ( .A(in_17bit_b[2]), .B(in_17bit_b[1]), .CI(
        add_3_root_r119_carry_3_), .CO(add_3_root_r119_carry_4_), .S(
        add_1_root_r119_A_3_) );
  ADDFX2 U111 ( .A(in_17bit_b[9]), .B(in_17bit_b[8]), .CI(
        add_2_root_r119_carry_13_), .CO(add_2_root_r119_carry_14_), .S(
        add_2_root_r119_SUM_13_) );
  ADDFX2 U112 ( .A(in_17bit_b[12]), .B(in_17bit_b[10]), .CI(
        add_2_root_r115_carry_13_), .CO(add_2_root_r115_carry_14_), .S(
        add_2_root_r115_SUM_13_) );
  ADDFX2 U113 ( .A(in_17bit_b[14]), .B(in_17bit_b[10]), .CI(
        add_1_root_r112_carry_14_), .CO(add_1_root_r112_carry_15_), .S(
        add_1_root_r112_SUM_14_) );
  ADDFX2 U114 ( .A(in_17bit_b[11]), .B(in_17bit_b[9]), .CI(
        add_1_root_r115_carry_15_), .CO(add_1_root_r115_carry_16_), .S(
        add_1_root_r115_SUM_15_) );
  ADDFX2 U115 ( .A(add_1_root_r119_A_15_), .B(in_17bit_b[9]), .CI(
        add_1_root_r119_carry[15]), .CO(add_1_root_r119_carry[16]), .S(
        add_1_root_r119_SUM_15_) );
  ADDFX2 U116 ( .A(in_17bit_b[10]), .B(in_17bit_b[9]), .CI(
        add_2_root_r119_carry_14_), .CO(add_2_root_r119_carry_15_), .S(
        add_2_root_r119_SUM_14_) );
  ADDFX2 U117 ( .A(in_17bit_b[13]), .B(in_17bit_b[11]), .CI(
        add_2_root_r115_carry_14_), .CO(add_2_root_r115_carry_15_), .S(
        add_2_root_r115_SUM_14_) );
  ADDFX2 U118 ( .A(in_17bit_b[15]), .B(in_17bit_b[11]), .CI(
        add_1_root_r112_carry_15_), .CO(add_1_root_r112_carry_16_), .S(
        add_1_root_r112_SUM_15_) );
  ADDFX2 U119 ( .A(in_17bit_b[12]), .B(in_17bit_b[10]), .CI(
        add_1_root_r115_carry_16_), .CO(add_1_root_r115_carry_17_), .S(
        add_1_root_r115_SUM_16_) );
  ADDFX2 U120 ( .A(add_1_root_r119_A_16_), .B(in_17bit_b[10]), .CI(
        add_1_root_r119_carry[16]), .CO(add_1_root_r119_carry[17]), .S(
        add_1_root_r119_SUM_16_) );
  ADDFX2 U121 ( .A(in_17bit_b[11]), .B(in_17bit_b[10]), .CI(
        add_2_root_r119_carry_15_), .CO(add_2_root_r119_carry_16_), .S(
        add_2_root_r119_SUM_15_) );
  ADDFX2 U122 ( .A(in_17bit_b[14]), .B(in_17bit_b[12]), .CI(
        add_2_root_r115_carry_15_), .CO(add_2_root_r115_carry_16_), .S(
        add_2_root_r115_SUM_15_) );
  ADDFX2 U123 ( .A(in_17bit_b[13]), .B(in_17bit_b[11]), .CI(
        add_1_root_r115_carry_17_), .CO(add_1_root_r115_carry_18_), .S(
        add_1_root_r115_SUM_17_) );
  ADDFX2 U124 ( .A(add_1_root_r119_A_17_), .B(in_17bit_b[11]), .CI(
        add_1_root_r119_carry[17]), .CO(add_1_root_r119_carry[18]), .S(
        add_1_root_r119_SUM_17_) );
  ADDFX2 U125 ( .A(in_17bit_b[12]), .B(in_17bit_b[11]), .CI(
        add_2_root_r119_carry_16_), .CO(add_2_root_r119_carry_17_), .S(
        add_2_root_r119_SUM_16_) );
  ADDFX2 U126 ( .A(in_17bit_b[14]), .B(in_17bit_b[12]), .CI(
        add_1_root_r115_carry_18_), .CO(add_1_root_r115_carry_19_), .S(
        add_1_root_r115_SUM_18_) );
  ADDFX2 U127 ( .A(add_1_root_r119_A_18_), .B(in_17bit_b[12]), .CI(
        add_1_root_r119_carry[18]), .CO(add_1_root_r119_carry[19]), .S(
        add_1_root_r119_SUM_18_) );
  ADDFX2 U128 ( .A(in_17bit_b[15]), .B(in_17bit_b[14]), .CI(
        add_3_root_r119_carry_16_), .CO(add_3_root_r119_carry_17_), .S(
        add_1_root_r119_A_16_) );
  ADDFX2 U129 ( .A(in_17bit_b[7]), .B(in_17bit_b[3]), .CI(
        add_1_root_r112_carry_7_), .CO(add_1_root_r112_carry_8_), .S(
        add_1_root_r112_SUM_7_) );
  ADDFX2 U130 ( .A(add_1_root_r119_A_9_), .B(in_17bit_b[3]), .CI(
        add_1_root_r119_carry[9]), .CO(add_1_root_r119_carry[10]), .S(
        add_1_root_r119_SUM_9_) );
  ADDFX2 U131 ( .A(in_17bit_b[4]), .B(in_17bit_b[3]), .CI(
        add_2_root_r119_carry_8_), .CO(add_2_root_r119_carry_9_), .S(
        add_2_root_r119_SUM_8_) );
  ADDFX2 U132 ( .A(in_17bit_b[5]), .B(in_17bit_b[3]), .CI(
        add_1_root_r115_carry_9_), .CO(add_1_root_r115_carry_10_), .S(
        add_1_root_r115_SUM_9_) );
  ADDFX2 U133 ( .A(in_17bit_b[5]), .B(in_17bit_b[4]), .CI(
        add_3_root_r119_carry_6_), .CO(add_3_root_r119_carry_7_), .S(
        add_1_root_r119_A_6_) );
  ADDFX2 U134 ( .A(in_17bit_b[15]), .B(in_17bit_b[13]), .CI(
        add_2_root_r115_carry_16_), .CO(add_2_root_r115_carry_17_), .S(
        add_2_root_r115_SUM_16_) );
  ADDFX2 U135 ( .A(in_17bit_b[13]), .B(in_17bit_b[12]), .CI(
        add_2_root_r119_carry_17_), .CO(add_2_root_r119_carry_18_), .S(
        add_2_root_r119_SUM_17_) );
  ADDFX2 U136 ( .A(in_17bit_b[5]), .B(in_17bit_b[3]), .CI(
        add_2_root_r115_carry_6_), .CO(add_2_root_r115_carry_7_), .S(
        add_2_root_r115_SUM_6_) );
  ADDFX2 U137 ( .A(in_17bit_b[4]), .B(in_17bit_b[3]), .CI(
        add_3_root_r119_carry_5_), .CO(add_3_root_r119_carry_6_), .S(
        add_1_root_r119_A_5_) );
  ADDFX2 U138 ( .A(in_17bit_b[15]), .B(in_17bit_b[13]), .CI(
        add_1_root_r115_carry_19_), .CO(add_1_root_r115_carry_20_), .S(
        add_1_root_r115_SUM_19_) );
  ADDFX2 U139 ( .A(in_17bit_b[14]), .B(in_17bit_b[13]), .CI(
        add_2_root_r119_carry_18_), .CO(add_2_root_r119_carry_19_), .S(
        add_2_root_r119_SUM_18_) );
  ADDFX2 U140 ( .A(in_17bit_b[15]), .B(in_17bit_b[14]), .CI(
        add_2_root_r119_carry_19_), .CO(add_2_root_r119_carry_20_), .S(
        add_2_root_r119_SUM_19_) );
  INVX1 U141 ( .A(n201), .Y(n83) );
  BUFX3 U142 ( .A(in_17bit_b[16]), .Y(n44) );
  INVX1 U143 ( .A(n256), .Y(in_17bit_b[16]) );
  NAND2X1 U144 ( .A(n247), .B(n246), .Y(N461) );
  AOI22X1 U145 ( .A0(N122), .A1(n249), .B0(N219), .B1(n42), .Y(n246) );
  AOI22X1 U146 ( .A0(N361), .A1(n41), .B0(n174), .B1(in_17bit_b[14]), .Y(n247)
         );
  NAND2X1 U147 ( .A(n251), .B(n250), .Y(N462) );
  AOI22X1 U148 ( .A0(N123), .A1(n249), .B0(N220), .B1(n42), .Y(n250) );
  AOI22X1 U149 ( .A0(N362), .A1(n41), .B0(n174), .B1(in_17bit_b[15]), .Y(n251)
         );
  BUFX3 U150 ( .A(in_8bit[5]), .Y(n47) );
  INVX1 U151 ( .A(in_8bit[0]), .Y(n46) );
  INVX1 U152 ( .A(in_8bit[3]), .Y(n48) );
  INVX1 U153 ( .A(n54), .Y(n49) );
  INVX1 U154 ( .A(in_8bit[4]), .Y(n45) );
  XNOR2X1 U155 ( .A(n56), .B(n25), .Y(N29) );
  NAND2X1 U156 ( .A(sub_add_54_b0_carry[15]), .B(n172), .Y(n25) );
  CLKINVX3 U157 ( .A(n203), .Y(in_17bit_b[0]) );
  NOR3X1 U158 ( .A(n175), .B(n48), .C(n46), .Y(n201) );
  NAND4BXL U159 ( .AN(n43), .B(in_8bit[4]), .C(n47), .D(n200), .Y(n85) );
  NAND3BX1 U160 ( .AN(n47), .B(n175), .C(in_8bit[3]), .Y(n196) );
  CLKINVX3 U161 ( .A(n248), .Y(in_17bit_b[15]) );
  BUFX3 U162 ( .A(n252), .Y(n41) );
  OAI2BB1X1 U163 ( .A0N(n26), .A1N(n33), .B0(n89), .Y(n252) );
  NAND2BX1 U164 ( .AN(n196), .B(n32), .Y(n89) );
  BUFX3 U165 ( .A(n253), .Y(n42) );
  OAI2BB1X1 U166 ( .A0N(n33), .A1N(n32), .B0(n90), .Y(n253) );
  NAND2BX1 U167 ( .AN(n196), .B(n26), .Y(n90) );
  OAI2BB1X1 U168 ( .A0N(n87), .A1N(n86), .B0(n85), .Y(n249) );
  NOR2BX1 U169 ( .AN(in_8bit[1]), .B(n91), .Y(n86) );
  NOR2X1 U170 ( .A(n84), .B(n83), .Y(n87) );
  OAI2BB1X1 U171 ( .A0N(n200), .A1N(n94), .B0(n93), .Y(n174) );
  INVX1 U172 ( .A(n91), .Y(n94) );
  NAND3BX1 U173 ( .AN(n92), .B(n201), .C(n47), .Y(n93) );
  AND2X2 U174 ( .A(n88), .B(n46), .Y(n26) );
  NAND2X1 U175 ( .A(n205), .B(n204), .Y(N447) );
  AOI22X1 U176 ( .A0(N108), .A1(n249), .B0(N205), .B1(n42), .Y(n204) );
  AOI22X1 U177 ( .A0(N347), .A1(n41), .B0(n174), .B1(in_17bit_b[0]), .Y(n205)
         );
  NAND2X1 U178 ( .A(n208), .B(n207), .Y(N448) );
  AOI22X1 U179 ( .A0(N109), .A1(n249), .B0(N206), .B1(n42), .Y(n207) );
  AOI22X1 U180 ( .A0(N348), .A1(n41), .B0(n174), .B1(n173), .Y(n208) );
  INVX1 U181 ( .A(n206), .Y(n173) );
  NAND2X1 U182 ( .A(n211), .B(n210), .Y(N449) );
  AOI22X1 U183 ( .A0(N110), .A1(n249), .B0(N207), .B1(n42), .Y(n210) );
  AOI22X1 U184 ( .A0(N349), .A1(n41), .B0(n174), .B1(in_17bit_b[2]), .Y(n211)
         );
  NAND2X1 U185 ( .A(n214), .B(n213), .Y(N450) );
  AOI22X1 U186 ( .A0(N111), .A1(n249), .B0(N208), .B1(n42), .Y(n213) );
  AOI22X1 U187 ( .A0(N350), .A1(n41), .B0(n174), .B1(in_17bit_b[3]), .Y(n214)
         );
  NAND2X1 U188 ( .A(n217), .B(n216), .Y(N451) );
  AOI22X1 U189 ( .A0(N112), .A1(n249), .B0(N209), .B1(n42), .Y(n216) );
  AOI22X1 U190 ( .A0(N351), .A1(n41), .B0(n174), .B1(in_17bit_b[4]), .Y(n217)
         );
  NAND2X1 U191 ( .A(n220), .B(n219), .Y(N452) );
  AOI22X1 U192 ( .A0(N113), .A1(n249), .B0(N210), .B1(n42), .Y(n219) );
  AOI22X1 U193 ( .A0(N352), .A1(n41), .B0(n174), .B1(in_17bit_b[5]), .Y(n220)
         );
  NAND2X1 U194 ( .A(n223), .B(n222), .Y(N453) );
  AOI22X1 U195 ( .A0(N114), .A1(n249), .B0(N211), .B1(n42), .Y(n222) );
  AOI22X1 U196 ( .A0(N353), .A1(n41), .B0(n174), .B1(in_17bit_b[6]), .Y(n223)
         );
  NAND2X1 U197 ( .A(n226), .B(n225), .Y(N454) );
  AOI22X1 U198 ( .A0(N115), .A1(n249), .B0(N212), .B1(n42), .Y(n225) );
  AOI22X1 U199 ( .A0(N354), .A1(n41), .B0(n174), .B1(in_17bit_b[7]), .Y(n226)
         );
  NAND2X1 U200 ( .A(n229), .B(n228), .Y(N455) );
  AOI22X1 U201 ( .A0(N116), .A1(n249), .B0(N213), .B1(n42), .Y(n228) );
  AOI22X1 U202 ( .A0(N355), .A1(n41), .B0(n174), .B1(in_17bit_b[8]), .Y(n229)
         );
  NAND2X1 U203 ( .A(n232), .B(n231), .Y(N456) );
  AOI22X1 U204 ( .A0(N117), .A1(n249), .B0(N214), .B1(n42), .Y(n231) );
  AOI22X1 U205 ( .A0(N356), .A1(n41), .B0(n174), .B1(in_17bit_b[9]), .Y(n232)
         );
  NAND2X1 U206 ( .A(n235), .B(n234), .Y(N457) );
  AOI22X1 U207 ( .A0(N118), .A1(n249), .B0(N215), .B1(n42), .Y(n234) );
  AOI22X1 U208 ( .A0(N357), .A1(n41), .B0(n174), .B1(in_17bit_b[10]), .Y(n235)
         );
  NAND2X1 U209 ( .A(n238), .B(n237), .Y(N458) );
  AOI22X1 U210 ( .A0(N119), .A1(n249), .B0(N216), .B1(n42), .Y(n237) );
  AOI22X1 U211 ( .A0(N358), .A1(n41), .B0(n174), .B1(in_17bit_b[11]), .Y(n238)
         );
  NAND2X1 U212 ( .A(n241), .B(n240), .Y(N459) );
  AOI22X1 U213 ( .A0(N120), .A1(n249), .B0(N217), .B1(n42), .Y(n240) );
  AOI22X1 U214 ( .A0(N359), .A1(n41), .B0(n174), .B1(in_17bit_b[12]), .Y(n241)
         );
  NAND2X1 U215 ( .A(n244), .B(n243), .Y(N460) );
  AOI22X1 U216 ( .A0(N121), .A1(n249), .B0(N218), .B1(n42), .Y(n243) );
  AOI22X1 U217 ( .A0(N360), .A1(n41), .B0(n174), .B1(in_17bit_b[13]), .Y(n244)
         );
  OAI21XL U218 ( .A0(n43), .A1(n59), .B0(n58), .Y(n63) );
  OAI21XL U219 ( .A0(n43), .A1(n68), .B0(n67), .Y(n72) );
  MXI2XL U220 ( .A(n3), .B(n18), .S0(n82), .Y(out[16]) );
  NOR4BXL U221 ( .AN(n197), .B(n46), .C(in_8bit[1]), .D(in_8bit[2]), .Y(n200)
         );
  INVXL U222 ( .A(in_8bit[2]), .Y(n175) );
  NAND4BBX1 U223 ( .AN(n41), .BN(n42), .C(n202), .D(n255), .Y(N446) );
  AOI2BB1X1 U224 ( .A0N(n199), .A1N(n198), .B0(n249), .Y(n202) );
  OR4X1 U225 ( .A(in_8bit[1]), .B(in_8bit[0]), .C(in_8bit[2]), .D(in_8bit[3]), 
        .Y(n198) );
  AOI22X1 U226 ( .A0(N27), .A1(n52), .B0(in_17bit[14]), .B1(n54), .Y(n245) );
  AOI22X1 U227 ( .A0(N28), .A1(n52), .B0(in_17bit[15]), .B1(n54), .Y(n248) );
  AOI22X1 U228 ( .A0(N16), .A1(n52), .B0(in_17bit[3]), .B1(n55), .Y(n212) );
  AOI22X1 U229 ( .A0(N17), .A1(n52), .B0(in_17bit[4]), .B1(n55), .Y(n215) );
  AOI22X1 U230 ( .A0(N18), .A1(n52), .B0(in_17bit[5]), .B1(n54), .Y(n218) );
  AOI22X1 U231 ( .A0(N19), .A1(n52), .B0(in_17bit[6]), .B1(n56), .Y(n221) );
  AOI22X1 U232 ( .A0(N20), .A1(n52), .B0(in_17bit[7]), .B1(n54), .Y(n224) );
  AOI22X1 U233 ( .A0(N21), .A1(n52), .B0(in_17bit[8]), .B1(n56), .Y(n227) );
  AOI22X1 U234 ( .A0(N22), .A1(n52), .B0(in_17bit[9]), .B1(n56), .Y(n230) );
  AOI22X1 U235 ( .A0(N23), .A1(n52), .B0(in_17bit[10]), .B1(n55), .Y(n233) );
  AOI22X1 U236 ( .A0(N24), .A1(n52), .B0(in_17bit[11]), .B1(n55), .Y(n236) );
  AOI22X1 U237 ( .A0(N25), .A1(n52), .B0(in_17bit[12]), .B1(n55), .Y(n239) );
  AOI22X1 U238 ( .A0(N26), .A1(n52), .B0(in_17bit[13]), .B1(n54), .Y(n242) );
  INVXL U239 ( .A(in_8bit[6]), .Y(n84) );
  INVX1 U240 ( .A(n57), .Y(n74) );
  NAND2BX1 U241 ( .AN(n66), .B(n15), .Y(n57) );
  AND2X2 U242 ( .A(n74), .B(n5), .Y(n28) );
  AND2X2 U243 ( .A(n28), .B(n6), .Y(n29) );
  AND2X2 U244 ( .A(n29), .B(n7), .Y(n30) );
  AND2X2 U245 ( .A(n30), .B(n2), .Y(n31) );
  AND4X1 U246 ( .A(in_8bit[1]), .B(n43), .C(n195), .D(n46), .Y(n32) );
  NAND2X1 U247 ( .A(n36), .B(n4), .Y(n66) );
  AND2X2 U248 ( .A(n31), .B(n8), .Y(n34) );
  INVX1 U249 ( .A(in_17bit[4]), .Y(n99) );
  INVX1 U250 ( .A(in_17bit[5]), .Y(n100) );
  INVX1 U251 ( .A(in_17bit[6]), .Y(n101) );
  INVX1 U252 ( .A(in_17bit[7]), .Y(n158) );
  INVX1 U253 ( .A(in_17bit[8]), .Y(n160) );
  INVX1 U254 ( .A(in_17bit[9]), .Y(n163) );
  INVX1 U255 ( .A(in_17bit[10]), .Y(n164) );
  INVX1 U256 ( .A(in_17bit[11]), .Y(n167) );
  INVX1 U257 ( .A(in_17bit[12]), .Y(n168) );
  INVX1 U258 ( .A(in_17bit[13]), .Y(n170) );
  INVX1 U259 ( .A(in_17bit[14]), .Y(n171) );
  INVX1 U260 ( .A(in_17bit[15]), .Y(n172) );
  INVX1 U261 ( .A(in_17bit[2]), .Y(n97) );
  INVX1 U262 ( .A(in_17bit[3]), .Y(n98) );
  INVX1 U263 ( .A(in_17bit[1]), .Y(n96) );
  INVX1 U264 ( .A(in_17bit[0]), .Y(n95) );
  XNOR2X1 U265 ( .A(n16), .B(sub_add_75_b0_carry[10]), .Y(n35) );
  MX2X1 U266 ( .A(neg_mul[21]), .B(N479), .S0(n82), .Y(out[14]) );
  MX2X1 U267 ( .A(neg_mul[22]), .B(N480), .S0(n82), .Y(out[15]) );
  INVX1 U268 ( .A(n68), .Y(n69) );
  AOI2BB2X1 U269 ( .B0(n60), .B1(n43), .A0N(n43), .A1N(neg_mul[8]), .Y(n61) );
  INVX1 U270 ( .A(n59), .Y(n60) );
  NOR2X1 U271 ( .A(out[0]), .B(neg_mul[8]), .Y(n36) );
  NAND2X1 U272 ( .A(out[0]), .B(neg_mul[8]), .Y(n59) );
  NAND2X1 U273 ( .A(neg_mul[10]), .B(n66), .Y(n68) );
  NAND2X1 U274 ( .A(sub_add_75_b0_carry[15]), .B(n10), .Y(n37) );
  NOR2X2 U275 ( .A(n53), .B(n70), .Y(n71) );
  NAND2XL U276 ( .A(N29), .B(n40), .Y(n256) );
  AOI22XL U277 ( .A0(N14), .A1(n40), .B0(in_17bit[1]), .B1(n56), .Y(n206) );
  AOI22XL U278 ( .A0(N15), .A1(n40), .B0(in_17bit[2]), .B1(n55), .Y(n209) );
  AOI22XL U279 ( .A0(in_17bit[0]), .A1(n40), .B0(in_17bit[0]), .B1(n56), .Y(
        n203) );
  OR4X1 U280 ( .A(in_8bit[4]), .B(n47), .C(in_8bit[6]), .D(n43), .Y(n199) );
  NOR2XL U281 ( .A(in_8bit[6]), .B(in_8bit[3]), .Y(n197) );
  NOR2XL U282 ( .A(in_8bit[6]), .B(in_8bit[4]), .Y(n195) );
  NAND4BXL U283 ( .AN(n43), .B(in_8bit[4]), .C(in_8bit[6]), .D(in_8bit[1]), 
        .Y(n92) );
  AOI211X4 U284 ( .A0(n53), .A1(n72), .B0(n71), .C0(n74), .Y(out[3]) );
  XNOR2X4 U285 ( .A(n65), .B(n4), .Y(out[2]) );
  XNOR2X4 U286 ( .A(n75), .B(n5), .Y(out[4]) );
  NOR2X4 U287 ( .A(n28), .B(n73), .Y(n76) );
  XNOR2X4 U288 ( .A(n76), .B(n6), .Y(out[5]) );
  XNOR2X4 U289 ( .A(n40), .B(n43), .Y(n80) );
  NOR2X4 U290 ( .A(n29), .B(n80), .Y(n77) );
  XNOR2X4 U291 ( .A(n77), .B(n7), .Y(out[6]) );
  NOR2X4 U292 ( .A(n31), .B(n80), .Y(n79) );
  XNOR2X4 U293 ( .A(n79), .B(n8), .Y(out[8]) );
  MXI2X4 U294 ( .A(n16), .B(n35), .S0(n82), .Y(out[10]) );
  AND2X1 U295 ( .A(add_1_root_r112_carry_20_), .B(n44), .Y(
        add_1_root_r112_SUM_21_) );
  XOR2X1 U296 ( .A(n44), .B(add_1_root_r112_carry_20_), .Y(
        add_1_root_r112_SUM_20_) );
  AND2X1 U297 ( .A(add_1_root_r112_carry_19_), .B(in_17bit_b[15]), .Y(
        add_1_root_r112_carry_20_) );
  XOR2X1 U298 ( .A(in_17bit_b[15]), .B(add_1_root_r112_carry_19_), .Y(
        add_1_root_r112_SUM_19_) );
  AND2X1 U299 ( .A(add_1_root_r112_carry_18_), .B(in_17bit_b[14]), .Y(
        add_1_root_r112_carry_19_) );
  XOR2X1 U300 ( .A(in_17bit_b[14]), .B(add_1_root_r112_carry_18_), .Y(
        add_1_root_r112_SUM_18_) );
  AND2X1 U301 ( .A(add_1_root_r112_carry_17_), .B(in_17bit_b[13]), .Y(
        add_1_root_r112_carry_18_) );
  XOR2X1 U302 ( .A(in_17bit_b[13]), .B(add_1_root_r112_carry_17_), .Y(
        add_1_root_r112_SUM_17_) );
  AND2X1 U303 ( .A(add_2_root_r119_carry_21_), .B(n44), .Y(
        add_2_root_r119_SUM_22_) );
  XOR2X1 U304 ( .A(n44), .B(add_2_root_r119_carry_21_), .Y(
        add_2_root_r119_SUM_21_) );
  AND2X1 U305 ( .A(in_17bit_b[1]), .B(in_17bit_b[0]), .Y(
        add_2_root_r119_carry_6_) );
  XOR2X1 U306 ( .A(in_17bit_b[0]), .B(in_17bit_b[1]), .Y(
        add_2_root_r119_SUM_5_) );
  AND2X1 U307 ( .A(add_1_root_r119_carry[22]), .B(n44), .Y(
        add_1_root_r119_SUM_23_) );
  XOR2X1 U308 ( .A(n44), .B(add_1_root_r119_carry[22]), .Y(
        add_1_root_r119_SUM_22_) );
  AND2X1 U309 ( .A(add_1_root_r119_carry[21]), .B(in_17bit_b[15]), .Y(
        add_1_root_r119_carry[22]) );
  XOR2X1 U310 ( .A(in_17bit_b[15]), .B(add_1_root_r119_carry[21]), .Y(
        add_1_root_r119_SUM_21_) );
  AND2X1 U311 ( .A(add_1_root_r119_carry[20]), .B(in_17bit_b[14]), .Y(
        add_1_root_r119_carry[21]) );
  XOR2X1 U312 ( .A(in_17bit_b[14]), .B(add_1_root_r119_carry[20]), .Y(
        add_1_root_r119_SUM_20_) );
  AND2X1 U313 ( .A(add_1_root_r119_A_6_), .B(in_17bit_b[0]), .Y(
        add_1_root_r119_carry[7]) );
  XOR2X1 U314 ( .A(in_17bit_b[0]), .B(add_1_root_r119_A_6_), .Y(
        add_1_root_r119_SUM_6_) );
  AND2X1 U315 ( .A(add_3_root_r119_carry_18_), .B(n44), .Y(
        add_1_root_r119_A_19_) );
  XOR2X1 U316 ( .A(n44), .B(add_3_root_r119_carry_18_), .Y(
        add_1_root_r119_A_18_) );
  AND2X1 U317 ( .A(in_17bit_b[1]), .B(in_17bit_b[0]), .Y(
        add_3_root_r119_carry_3_) );
  XOR2X1 U318 ( .A(in_17bit_b[0]), .B(in_17bit_b[1]), .Y(add_1_root_r119_A_2_)
         );
  AND2X1 U319 ( .A(add_2_root_r115_carry_19_), .B(n44), .Y(
        add_2_root_r115_SUM_20_) );
  XOR2X1 U320 ( .A(n44), .B(add_2_root_r115_carry_19_), .Y(
        add_2_root_r115_SUM_19_) );
  AND2X1 U321 ( .A(add_2_root_r115_carry_18_), .B(in_17bit_b[15]), .Y(
        add_2_root_r115_carry_19_) );
  XOR2X1 U322 ( .A(in_17bit_b[15]), .B(add_2_root_r115_carry_18_), .Y(
        add_2_root_r115_SUM_18_) );
  AND2X1 U323 ( .A(in_17bit_b[2]), .B(in_17bit_b[0]), .Y(
        add_2_root_r115_carry_4_) );
  XOR2X1 U324 ( .A(in_17bit_b[0]), .B(in_17bit_b[2]), .Y(
        add_2_root_r115_SUM_3_) );
  AND2X1 U325 ( .A(add_1_root_r115_carry_22_), .B(n44), .Y(
        add_1_root_r115_SUM_23_) );
  XOR2X1 U326 ( .A(n44), .B(add_1_root_r115_carry_22_), .Y(
        add_1_root_r115_SUM_22_) );
  AND2X1 U327 ( .A(add_1_root_r115_carry_21_), .B(in_17bit_b[15]), .Y(
        add_1_root_r115_carry_22_) );
  XOR2X1 U328 ( .A(in_17bit_b[15]), .B(add_1_root_r115_carry_21_), .Y(
        add_1_root_r115_SUM_21_) );
  AND2X1 U329 ( .A(in_17bit_b[2]), .B(in_17bit_b[0]), .Y(
        add_1_root_r115_carry_7_) );
  XOR2X1 U330 ( .A(in_17bit_b[0]), .B(in_17bit_b[2]), .Y(
        add_1_root_r115_SUM_6_) );
  XOR2X1 U331 ( .A(n172), .B(sub_add_54_b0_carry[15]), .Y(N28) );
  AND2X1 U332 ( .A(sub_add_54_b0_carry[14]), .B(n171), .Y(
        sub_add_54_b0_carry[15]) );
  XOR2X1 U333 ( .A(n171), .B(sub_add_54_b0_carry[14]), .Y(N27) );
  AND2X1 U334 ( .A(sub_add_54_b0_carry[13]), .B(n170), .Y(
        sub_add_54_b0_carry[14]) );
  XOR2X1 U335 ( .A(n170), .B(sub_add_54_b0_carry[13]), .Y(N26) );
  AND2X1 U336 ( .A(sub_add_54_b0_carry[12]), .B(n168), .Y(
        sub_add_54_b0_carry[13]) );
  XOR2X1 U337 ( .A(n168), .B(sub_add_54_b0_carry[12]), .Y(N25) );
  AND2X1 U338 ( .A(sub_add_54_b0_carry[11]), .B(n167), .Y(
        sub_add_54_b0_carry[12]) );
  XOR2X1 U339 ( .A(n167), .B(sub_add_54_b0_carry[11]), .Y(N24) );
  AND2X1 U340 ( .A(sub_add_54_b0_carry[10]), .B(n164), .Y(
        sub_add_54_b0_carry[11]) );
  XOR2X1 U341 ( .A(n164), .B(sub_add_54_b0_carry[10]), .Y(N23) );
  AND2X1 U342 ( .A(sub_add_54_b0_carry[9]), .B(n163), .Y(
        sub_add_54_b0_carry[10]) );
  XOR2X1 U343 ( .A(n163), .B(sub_add_54_b0_carry[9]), .Y(N22) );
  AND2X1 U344 ( .A(sub_add_54_b0_carry[8]), .B(n160), .Y(
        sub_add_54_b0_carry[9]) );
  XOR2X1 U345 ( .A(n160), .B(sub_add_54_b0_carry[8]), .Y(N21) );
  AND2X1 U346 ( .A(sub_add_54_b0_carry[7]), .B(n158), .Y(
        sub_add_54_b0_carry[8]) );
  XOR2X1 U347 ( .A(n158), .B(sub_add_54_b0_carry[7]), .Y(N20) );
  AND2X1 U348 ( .A(sub_add_54_b0_carry[6]), .B(n101), .Y(
        sub_add_54_b0_carry[7]) );
  XOR2X1 U349 ( .A(n101), .B(sub_add_54_b0_carry[6]), .Y(N19) );
  AND2X1 U350 ( .A(sub_add_54_b0_carry[5]), .B(n100), .Y(
        sub_add_54_b0_carry[6]) );
  XOR2X1 U351 ( .A(n100), .B(sub_add_54_b0_carry[5]), .Y(N18) );
  AND2X1 U352 ( .A(sub_add_54_b0_carry[4]), .B(n99), .Y(sub_add_54_b0_carry[5]) );
  XOR2X1 U353 ( .A(n99), .B(sub_add_54_b0_carry[4]), .Y(N17) );
  AND2X1 U354 ( .A(sub_add_54_b0_carry[3]), .B(n98), .Y(sub_add_54_b0_carry[4]) );
  XOR2X1 U355 ( .A(n98), .B(sub_add_54_b0_carry[3]), .Y(N16) );
  AND2X1 U356 ( .A(sub_add_54_b0_carry[2]), .B(n97), .Y(sub_add_54_b0_carry[3]) );
  XOR2X1 U357 ( .A(n97), .B(sub_add_54_b0_carry[2]), .Y(N15) );
  AND2X1 U358 ( .A(n95), .B(n96), .Y(sub_add_54_b0_carry[2]) );
  XOR2X1 U359 ( .A(n96), .B(n95), .Y(N14) );
  XOR2X1 U360 ( .A(n10), .B(sub_add_75_b0_carry[15]), .Y(N480) );
  AND2X1 U361 ( .A(sub_add_75_b0_carry[14]), .B(n14), .Y(
        sub_add_75_b0_carry[15]) );
  XOR2X1 U362 ( .A(n14), .B(sub_add_75_b0_carry[14]), .Y(N479) );
  AND2X1 U363 ( .A(sub_add_75_b0_carry[13]), .B(n12), .Y(
        sub_add_75_b0_carry[14]) );
  XOR2X1 U364 ( .A(n12), .B(sub_add_75_b0_carry[13]), .Y(N478) );
  AND2X1 U365 ( .A(sub_add_75_b0_carry[12]), .B(n13), .Y(
        sub_add_75_b0_carry[13]) );
  XOR2X1 U366 ( .A(n13), .B(sub_add_75_b0_carry[12]), .Y(N477) );
  AND2X1 U367 ( .A(sub_add_75_b0_carry[11]), .B(n11), .Y(
        sub_add_75_b0_carry[12]) );
  XOR2X1 U368 ( .A(n11), .B(sub_add_75_b0_carry[11]), .Y(N476) );
  AND2X1 U369 ( .A(sub_add_75_b0_carry[10]), .B(n16), .Y(
        sub_add_75_b0_carry[11]) );
  AND2X1 U370 ( .A(n34), .B(n9), .Y(sub_add_75_b0_carry[10]) );
  AND2X1 U371 ( .A(in_17bit_b[0]), .B(in_17bit_b[4]), .Y(
        add_1_root_r112_carry_5_) );
endmodule


module multi16_3_DW01_add_0 ( A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, 
        A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, 
        A_4_, B_23_, B_22_, B_21_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, 
        B_14_, B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, 
        SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, 
        SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, 
        SUM_7_ );
  input A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_,
         A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, B_23_, B_22_,
         B_21_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_,
         B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_;
  output SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_,
         SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_,
         SUM_8_, SUM_7_;
  wire   n1, n2, n3, n4;
  wire   [23:7] carry;

  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry[7]), .CO(carry[8]), .S(SUM_7_)
         );
  ADDFX2 U1_21 ( .A(A_21_), .B(B_21_), .CI(carry[21]), .CO(carry[22]), .S(
        SUM_21_) );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry[20]), .CO(carry[21]), .S(
        SUM_20_) );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry[19]), .CO(carry[20]), .S(
        SUM_19_) );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry[18]), .CO(carry[19]), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry[17]), .CO(carry[18]), .S(
        SUM_17_) );
  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry[16]), .CO(carry[17]), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry[15]), .CO(carry[16]), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry[14]), .CO(carry[15]), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry[13]), .CO(carry[14]), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry[12]), .CO(carry[13]), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry[11]), .CO(carry[12]), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry[10]), .CO(carry[11]), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry[9]), .CO(carry[10]), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry[8]), .CO(carry[9]), .S(SUM_8_)
         );
  ADDFX2 U1_22 ( .A(A_22_), .B(B_22_), .CI(carry[22]), .CO(carry[23]), .S(
        SUM_22_) );
  AND2X2 U1 ( .A(A_4_), .B(B_4_), .Y(n1) );
  XOR2X1 U2 ( .A(B_23_), .B(carry[23]), .Y(SUM_23_) );
  OAI2BB1X1 U3 ( .A0N(n2), .A1N(A_6_), .B0(n3), .Y(carry[7]) );
  OAI21XL U4 ( .A0(A_6_), .A1(n2), .B0(B_6_), .Y(n3) );
  OAI2BB1X1 U5 ( .A0N(n1), .A1N(A_5_), .B0(n4), .Y(n2) );
  OAI21XL U6 ( .A0(A_5_), .A1(n1), .B0(B_5_), .Y(n4) );
endmodule


module multi16_3_DW01_add_4 ( A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, 
        A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, 
        B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, 
        B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, SUM_22_, SUM_21_, SUM_20_, 
        SUM_19_, SUM_18_, SUM_17_, SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, 
        SUM_11_, SUM_10_, SUM_9_, SUM_8_, SUM_7_ );
  input A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_,
         A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, B_20_, B_19_,
         B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, B_10_, B_9_,
         B_8_, B_7_, B_6_, B_5_;
  output SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_,
         SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_,
         SUM_7_;
  wire   carry_21_, carry_20_, carry_19_, carry_18_, carry_17_, carry_16_,
         carry_15_, carry_14_, carry_13_, carry_12_, carry_11_, carry_10_,
         carry_9_, carry_8_, carry_7_, n1;

  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry_16_), .CO(carry_17_), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry_15_), .CO(carry_16_), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry_14_), .CO(carry_15_), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry_13_), .CO(carry_14_), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry_12_), .CO(carry_13_), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry_11_), .CO(carry_12_), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry_10_), .CO(carry_11_), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry_9_), .CO(carry_10_), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry_8_), .CO(carry_9_), .S(SUM_8_)
         );
  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry_7_), .CO(carry_8_), .S(SUM_7_)
         );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry_20_), .CO(carry_21_), .S(
        SUM_20_) );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry_19_), .CO(carry_20_), .S(
        SUM_19_) );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry_18_), .CO(carry_19_), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry_17_), .CO(carry_18_), .S(
        SUM_17_) );
  ADDFX2 U1_21 ( .A(A_21_), .B(B_21_), .CI(carry_21_), .CO(SUM_22_), .S(
        SUM_21_) );
  OAI2BB1X1 U1 ( .A0N(A_6_), .A1N(B_6_), .B0(n1), .Y(carry_7_) );
  OAI211X1 U2 ( .A0(B_6_), .A1(A_6_), .B0(A_5_), .C0(B_5_), .Y(n1) );
endmodule


module multi16_3_DW01_add_6 ( A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, 
        A_16_, A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, 
        A_6_, A_5_, A_4_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, 
        B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, 
        SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, 
        SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, 
        SUM_7_ );
  input A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_,
         A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, B_20_,
         B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, B_10_,
         B_9_, B_8_, B_7_, B_6_, B_5_, B_4_;
  output SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_,
         SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_,
         SUM_8_, SUM_7_;
  wire   n1, n2, n3, n4, n5, n6;
  wire   [21:7] carry;

  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry[7]), .CO(carry[8]), .S(SUM_7_)
         );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry[18]), .CO(carry[19]), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry[17]), .CO(carry[18]), .S(
        SUM_17_) );
  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry[16]), .CO(carry[17]), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry[15]), .CO(carry[16]), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry[14]), .CO(carry[15]), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry[13]), .CO(carry[14]), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry[12]), .CO(carry[13]), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry[11]), .CO(carry[12]), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry[10]), .CO(carry[11]), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry[9]), .CO(carry[10]), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry[8]), .CO(carry[9]), .S(SUM_8_)
         );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry[19]), .CO(carry[20]), .S(
        SUM_19_) );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry[20]), .CO(carry[21]), .S(
        SUM_20_) );
  AND2X2 U1 ( .A(A_22_), .B(n2), .Y(n1) );
  AND2X2 U2 ( .A(A_21_), .B(carry[21]), .Y(n2) );
  AND2X2 U3 ( .A(A_4_), .B(B_4_), .Y(n3) );
  XOR2X1 U4 ( .A(A_23_), .B(n1), .Y(SUM_23_) );
  XOR2X1 U5 ( .A(A_21_), .B(carry[21]), .Y(SUM_21_) );
  XOR2X1 U6 ( .A(A_22_), .B(n2), .Y(SUM_22_) );
  OAI2BB1X1 U7 ( .A0N(n4), .A1N(A_6_), .B0(n5), .Y(carry[7]) );
  OAI21XL U8 ( .A0(A_6_), .A1(n4), .B0(B_6_), .Y(n5) );
  OAI2BB1X1 U9 ( .A0N(n3), .A1N(A_5_), .B0(n6), .Y(n4) );
  OAI21XL U10 ( .A0(A_5_), .A1(n3), .B0(B_5_), .Y(n6) );
endmodule


module multi16_3 ( in_17bit, in_8bit, out );
  input [16:0] in_17bit;
  input [7:0] in_8bit;
  output [16:0] out;
  wire   N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27,
         N28, N29, N108, N109, N110, N111, N112, N113, N114, N115, N116, N117,
         N118, N119, N120, N121, N122, N123, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220,
         N221, N347, N348, N349, N350, N351, N352, N353, N354, N355, N356,
         N357, N358, N359, N360, N361, N362, N363, N446, N447, N448, N449,
         N450, N451, N452, N453, N454, N455, N456, N457, N458, N459, N460,
         N461, N462, N463, N476, N477, N478, N479, N480, N481,
         add_2_root_r119_carry_10_, add_2_root_r119_carry_11_,
         add_2_root_r119_carry_12_, add_2_root_r119_carry_13_,
         add_2_root_r119_carry_14_, add_2_root_r119_carry_15_,
         add_2_root_r119_carry_16_, add_2_root_r119_carry_17_,
         add_2_root_r119_carry_18_, add_2_root_r119_carry_19_,
         add_2_root_r119_carry_20_, add_2_root_r119_carry_21_,
         add_2_root_r119_carry_6_, add_2_root_r119_carry_7_,
         add_2_root_r119_carry_8_, add_2_root_r119_carry_9_,
         add_2_root_r119_SUM_5_, add_2_root_r119_SUM_6_,
         add_2_root_r119_SUM_7_, add_2_root_r119_SUM_8_,
         add_2_root_r119_SUM_9_, add_2_root_r119_SUM_10_,
         add_2_root_r119_SUM_11_, add_2_root_r119_SUM_12_,
         add_2_root_r119_SUM_13_, add_2_root_r119_SUM_14_,
         add_2_root_r119_SUM_15_, add_2_root_r119_SUM_16_,
         add_2_root_r119_SUM_17_, add_2_root_r119_SUM_18_,
         add_2_root_r119_SUM_19_, add_2_root_r119_SUM_20_,
         add_2_root_r119_SUM_21_, add_2_root_r119_SUM_22_,
         add_1_root_r119_SUM_6_, add_1_root_r119_SUM_7_,
         add_1_root_r119_SUM_8_, add_1_root_r119_SUM_9_,
         add_1_root_r119_SUM_10_, add_1_root_r119_SUM_11_,
         add_1_root_r119_SUM_12_, add_1_root_r119_SUM_13_,
         add_1_root_r119_SUM_14_, add_1_root_r119_SUM_15_,
         add_1_root_r119_SUM_16_, add_1_root_r119_SUM_17_,
         add_1_root_r119_SUM_18_, add_1_root_r119_SUM_19_,
         add_1_root_r119_SUM_20_, add_1_root_r119_SUM_21_,
         add_1_root_r119_SUM_22_, add_1_root_r119_SUM_23_,
         add_1_root_r119_A_2_, add_1_root_r119_A_3_, add_1_root_r119_A_4_,
         add_1_root_r119_A_5_, add_1_root_r119_A_6_, add_1_root_r119_A_7_,
         add_1_root_r119_A_8_, add_1_root_r119_A_9_, add_1_root_r119_A_10_,
         add_1_root_r119_A_11_, add_1_root_r119_A_12_, add_1_root_r119_A_13_,
         add_1_root_r119_A_14_, add_1_root_r119_A_15_, add_1_root_r119_A_16_,
         add_1_root_r119_A_17_, add_1_root_r119_A_18_, add_1_root_r119_A_19_,
         add_3_root_r119_carry_10_, add_3_root_r119_carry_11_,
         add_3_root_r119_carry_12_, add_3_root_r119_carry_13_,
         add_3_root_r119_carry_14_, add_3_root_r119_carry_15_,
         add_3_root_r119_carry_16_, add_3_root_r119_carry_17_,
         add_3_root_r119_carry_18_, add_3_root_r119_carry_3_,
         add_3_root_r119_carry_4_, add_3_root_r119_carry_5_,
         add_3_root_r119_carry_6_, add_3_root_r119_carry_7_,
         add_3_root_r119_carry_8_, add_3_root_r119_carry_9_,
         add_1_root_r112_carry_10_, add_1_root_r112_carry_11_,
         add_1_root_r112_carry_12_, add_1_root_r112_carry_13_,
         add_1_root_r112_carry_14_, add_1_root_r112_carry_15_,
         add_1_root_r112_carry_16_, add_1_root_r112_carry_17_,
         add_1_root_r112_carry_18_, add_1_root_r112_carry_19_,
         add_1_root_r112_carry_20_, add_1_root_r112_carry_5_,
         add_1_root_r112_carry_6_, add_1_root_r112_carry_7_,
         add_1_root_r112_carry_8_, add_1_root_r112_carry_9_,
         add_1_root_r112_SUM_1_, add_1_root_r112_SUM_2_,
         add_1_root_r112_SUM_3_, add_1_root_r112_SUM_4_,
         add_1_root_r112_SUM_5_, add_1_root_r112_SUM_6_,
         add_1_root_r112_SUM_7_, add_1_root_r112_SUM_8_,
         add_1_root_r112_SUM_9_, add_1_root_r112_SUM_10_,
         add_1_root_r112_SUM_11_, add_1_root_r112_SUM_12_,
         add_1_root_r112_SUM_13_, add_1_root_r112_SUM_14_,
         add_1_root_r112_SUM_15_, add_1_root_r112_SUM_16_,
         add_1_root_r112_SUM_17_, add_1_root_r112_SUM_18_,
         add_1_root_r112_SUM_19_, add_1_root_r112_SUM_20_,
         add_1_root_r112_SUM_21_, add_2_root_r115_carry_10_,
         add_2_root_r115_carry_11_, add_2_root_r115_carry_12_,
         add_2_root_r115_carry_13_, add_2_root_r115_carry_14_,
         add_2_root_r115_carry_15_, add_2_root_r115_carry_16_,
         add_2_root_r115_carry_17_, add_2_root_r115_carry_18_,
         add_2_root_r115_carry_19_, add_2_root_r115_carry_4_,
         add_2_root_r115_carry_5_, add_2_root_r115_carry_6_,
         add_2_root_r115_carry_7_, add_2_root_r115_carry_8_,
         add_2_root_r115_carry_9_, add_2_root_r115_SUM_3_,
         add_2_root_r115_SUM_4_, add_2_root_r115_SUM_5_,
         add_2_root_r115_SUM_6_, add_2_root_r115_SUM_7_,
         add_2_root_r115_SUM_8_, add_2_root_r115_SUM_9_,
         add_2_root_r115_SUM_10_, add_2_root_r115_SUM_11_,
         add_2_root_r115_SUM_12_, add_2_root_r115_SUM_13_,
         add_2_root_r115_SUM_14_, add_2_root_r115_SUM_15_,
         add_2_root_r115_SUM_16_, add_2_root_r115_SUM_17_,
         add_2_root_r115_SUM_18_, add_2_root_r115_SUM_19_,
         add_2_root_r115_SUM_20_, add_1_root_r115_carry_10_,
         add_1_root_r115_carry_11_, add_1_root_r115_carry_12_,
         add_1_root_r115_carry_13_, add_1_root_r115_carry_14_,
         add_1_root_r115_carry_15_, add_1_root_r115_carry_16_,
         add_1_root_r115_carry_17_, add_1_root_r115_carry_18_,
         add_1_root_r115_carry_19_, add_1_root_r115_carry_20_,
         add_1_root_r115_carry_21_, add_1_root_r115_carry_22_,
         add_1_root_r115_carry_7_, add_1_root_r115_carry_8_,
         add_1_root_r115_carry_9_, add_1_root_r115_SUM_6_,
         add_1_root_r115_SUM_7_, add_1_root_r115_SUM_8_,
         add_1_root_r115_SUM_9_, add_1_root_r115_SUM_10_,
         add_1_root_r115_SUM_11_, add_1_root_r115_SUM_12_,
         add_1_root_r115_SUM_13_, add_1_root_r115_SUM_14_,
         add_1_root_r115_SUM_15_, add_1_root_r115_SUM_16_,
         add_1_root_r115_SUM_17_, add_1_root_r115_SUM_18_,
         add_1_root_r115_SUM_19_, add_1_root_r115_SUM_20_,
         add_1_root_r115_SUM_21_, add_1_root_r115_SUM_22_,
         add_1_root_r115_SUM_23_, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n158, n160, n161, n162, n163, n164, n168,
         n170, n171, n172, n173, n174, n175, n176, n177, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257;
  wire   [16:0] in_17bit_b;
  wire   [23:8] neg_mul;
  wire   [16:10] sub_add_75_b0_carry;
  wire   [16:2] sub_add_54_b0_carry;
  wire   [22:7] add_1_root_r119_carry;

  multi16_3_DW01_add_0 add_0_root_r119 ( .A_22_(add_2_root_r119_SUM_22_), 
        .A_21_(add_2_root_r119_SUM_21_), .A_20_(add_2_root_r119_SUM_20_), 
        .A_19_(add_2_root_r119_SUM_19_), .A_18_(add_2_root_r119_SUM_18_), 
        .A_17_(add_2_root_r119_SUM_17_), .A_16_(add_2_root_r119_SUM_16_), 
        .A_15_(add_2_root_r119_SUM_15_), .A_14_(add_2_root_r119_SUM_14_), 
        .A_13_(add_2_root_r119_SUM_13_), .A_12_(add_2_root_r119_SUM_12_), 
        .A_11_(add_2_root_r119_SUM_11_), .A_10_(add_2_root_r119_SUM_10_), 
        .A_9_(add_2_root_r119_SUM_9_), .A_8_(add_2_root_r119_SUM_8_), .A_7_(
        add_2_root_r119_SUM_7_), .A_6_(add_2_root_r119_SUM_6_), .A_5_(
        add_2_root_r119_SUM_5_), .A_4_(in_17bit_b[0]), .B_23_(
        add_1_root_r119_SUM_23_), .B_22_(add_1_root_r119_SUM_22_), .B_21_(
        add_1_root_r119_SUM_21_), .B_20_(add_1_root_r119_SUM_20_), .B_19_(
        add_1_root_r119_SUM_19_), .B_18_(add_1_root_r119_SUM_18_), .B_17_(
        add_1_root_r119_SUM_17_), .B_16_(add_1_root_r119_SUM_16_), .B_15_(
        add_1_root_r119_SUM_15_), .B_14_(add_1_root_r119_SUM_14_), .B_13_(
        add_1_root_r119_SUM_13_), .B_12_(add_1_root_r119_SUM_12_), .B_11_(
        add_1_root_r119_SUM_11_), .B_10_(add_1_root_r119_SUM_10_), .B_9_(
        add_1_root_r119_SUM_9_), .B_8_(add_1_root_r119_SUM_8_), .B_7_(
        add_1_root_r119_SUM_7_), .B_6_(add_1_root_r119_SUM_6_), .B_5_(
        add_1_root_r119_A_5_), .B_4_(add_1_root_r119_A_4_), .SUM_23_(N363), 
        .SUM_22_(N362), .SUM_21_(N361), .SUM_20_(N360), .SUM_19_(N359), 
        .SUM_18_(N358), .SUM_17_(N357), .SUM_16_(N356), .SUM_15_(N355), 
        .SUM_14_(N354), .SUM_13_(N353), .SUM_12_(N352), .SUM_11_(N351), 
        .SUM_10_(N350), .SUM_9_(N349), .SUM_8_(N348), .SUM_7_(N347) );
  multi16_3_DW01_add_4 add_0_root_r112 ( .A_21_(n31), .A_20_(in_17bit_b[15]), 
        .A_19_(in_17bit_b[14]), .A_18_(in_17bit_b[13]), .A_17_(in_17bit_b[12]), 
        .A_16_(in_17bit_b[11]), .A_15_(in_17bit_b[10]), .A_14_(in_17bit_b[9]), 
        .A_13_(in_17bit_b[8]), .A_12_(in_17bit_b[7]), .A_11_(in_17bit_b[6]), 
        .A_10_(in_17bit_b[5]), .A_9_(in_17bit_b[4]), .A_8_(in_17bit_b[3]), 
        .A_7_(in_17bit_b[2]), .A_6_(in_17bit_b[1]), .A_5_(in_17bit_b[0]), 
        .B_21_(add_1_root_r112_SUM_21_), .B_20_(add_1_root_r112_SUM_20_), 
        .B_19_(add_1_root_r112_SUM_19_), .B_18_(add_1_root_r112_SUM_18_), 
        .B_17_(add_1_root_r112_SUM_17_), .B_16_(add_1_root_r112_SUM_16_), 
        .B_15_(add_1_root_r112_SUM_15_), .B_14_(add_1_root_r112_SUM_14_), 
        .B_13_(add_1_root_r112_SUM_13_), .B_12_(add_1_root_r112_SUM_12_), 
        .B_11_(add_1_root_r112_SUM_11_), .B_10_(add_1_root_r112_SUM_10_), 
        .B_9_(add_1_root_r112_SUM_9_), .B_8_(add_1_root_r112_SUM_8_), .B_7_(
        add_1_root_r112_SUM_7_), .B_6_(add_1_root_r112_SUM_6_), .B_5_(
        add_1_root_r112_SUM_5_), .SUM_22_(N123), .SUM_21_(N122), .SUM_20_(N121), .SUM_19_(N120), .SUM_18_(N119), .SUM_17_(N118), .SUM_16_(N117), .SUM_15_(
        N116), .SUM_14_(N115), .SUM_13_(N114), .SUM_12_(N113), .SUM_11_(N112), 
        .SUM_10_(N111), .SUM_9_(N110), .SUM_8_(N109), .SUM_7_(N108) );
  multi16_3_DW01_add_6 add_0_root_r115 ( .A_23_(add_1_root_r115_SUM_23_), 
        .A_22_(add_1_root_r115_SUM_22_), .A_21_(add_1_root_r115_SUM_21_), 
        .A_20_(add_1_root_r115_SUM_20_), .A_19_(add_1_root_r115_SUM_19_), 
        .A_18_(add_1_root_r115_SUM_18_), .A_17_(add_1_root_r115_SUM_17_), 
        .A_16_(add_1_root_r115_SUM_16_), .A_15_(add_1_root_r115_SUM_15_), 
        .A_14_(add_1_root_r115_SUM_14_), .A_13_(add_1_root_r115_SUM_13_), 
        .A_12_(add_1_root_r115_SUM_12_), .A_11_(add_1_root_r115_SUM_11_), 
        .A_10_(add_1_root_r115_SUM_10_), .A_9_(add_1_root_r115_SUM_9_), .A_8_(
        add_1_root_r115_SUM_8_), .A_7_(add_1_root_r115_SUM_7_), .A_6_(
        add_1_root_r115_SUM_6_), .A_5_(in_17bit_b[1]), .A_4_(in_17bit_b[0]), 
        .B_20_(add_2_root_r115_SUM_20_), .B_19_(add_2_root_r115_SUM_19_), 
        .B_18_(add_2_root_r115_SUM_18_), .B_17_(add_2_root_r115_SUM_17_), 
        .B_16_(add_2_root_r115_SUM_16_), .B_15_(add_2_root_r115_SUM_15_), 
        .B_14_(add_2_root_r115_SUM_14_), .B_13_(add_2_root_r115_SUM_13_), 
        .B_12_(add_2_root_r115_SUM_12_), .B_11_(add_2_root_r115_SUM_11_), 
        .B_10_(add_2_root_r115_SUM_10_), .B_9_(add_2_root_r115_SUM_9_), .B_8_(
        add_2_root_r115_SUM_8_), .B_7_(add_2_root_r115_SUM_7_), .B_6_(
        add_2_root_r115_SUM_6_), .B_5_(add_2_root_r115_SUM_5_), .B_4_(
        add_2_root_r115_SUM_4_), .SUM_23_(N221), .SUM_22_(N220), .SUM_21_(N219), .SUM_20_(N218), .SUM_19_(N217), .SUM_18_(N216), .SUM_17_(N215), .SUM_16_(
        N214), .SUM_15_(N213), .SUM_14_(N212), .SUM_13_(N211), .SUM_12_(N210), 
        .SUM_11_(N209), .SUM_10_(N208), .SUM_9_(N207), .SUM_8_(N206), .SUM_7_(
        N205) );
  TLATX1 neg_mul_reg_16_ ( .G(N446), .D(N456), .QN(n5) );
  TLATX1 neg_mul_reg_15_ ( .G(N446), .D(N455), .QN(n4) );
  TLATX1 neg_mul_reg_14_ ( .G(N446), .D(N454), .QN(n3) );
  TLATX1 neg_mul_reg_11_ ( .G(N446), .D(N451), .QN(n2) );
  TLATX1 neg_mul_reg_9_ ( .G(N446), .D(N449), .Q(neg_mul[9]), .QN(n16) );
  TLATX1 neg_mul_reg_23_ ( .G(N446), .D(N463), .Q(neg_mul[23]), .QN(n15) );
  TLATX1 neg_mul_reg_22_ ( .G(N446), .D(N462), .Q(neg_mul[22]), .QN(n8) );
  TLATX1 neg_mul_reg_21_ ( .G(N446), .D(N461), .Q(neg_mul[21]), .QN(n9) );
  TLATX1 neg_mul_reg_20_ ( .G(N446), .D(N460), .Q(neg_mul[20]), .QN(n10) );
  TLATX1 neg_mul_reg_19_ ( .G(N446), .D(N459), .Q(neg_mul[19]), .QN(n12) );
  TLATX1 neg_mul_reg_18_ ( .G(N446), .D(N458), .Q(neg_mul[18]), .QN(n11) );
  TLATX1 neg_mul_reg_17_ ( .G(N446), .D(N457), .QN(n13) );
  TLATX1 neg_mul_reg_13_ ( .G(N446), .D(N453), .Q(neg_mul[13]), .QN(n7) );
  TLATX1 neg_mul_reg_12_ ( .G(N446), .D(N452), .Q(neg_mul[12]), .QN(n6) );
  TLATX1 neg_mul_reg_10_ ( .G(N446), .D(N450), .Q(neg_mul[10]), .QN(n1) );
  TLATX1 neg_mul_reg_8_ ( .G(N446), .D(N448), .Q(neg_mul[8]), .QN(n14) );
  TLATX1 neg_mul_reg_7_ ( .G(N446), .D(N447), .Q(out[0]) );
  MX2X2 U2 ( .A(neg_mul[21]), .B(N479), .S0(n17), .Y(out[14]) );
  MX2X2 U3 ( .A(neg_mul[22]), .B(N480), .S0(n17), .Y(out[15]) );
  OAI21X4 U4 ( .A0(n55), .A1(n50), .B0(n54), .Y(n56) );
  CLKINVX8 U5 ( .A(n42), .Y(n50) );
  INVX8 U6 ( .A(n51), .Y(n45) );
  INVX4 U7 ( .A(n42), .Y(n51) );
  INVX3 U8 ( .A(in_17bit[16]), .Y(n43) );
  AOI2BB2X4 U9 ( .B0(n39), .B1(n14), .A0N(n40), .A1N(n53), .Y(n55) );
  AOI2BB2X4 U10 ( .B0(n52), .B1(n39), .A0N(n40), .A1N(neg_mul[8]), .Y(n57) );
  AOI2BB2X4 U11 ( .B0(n39), .B1(n1), .A0N(n40), .A1N(n63), .Y(n65) );
  AOI2BB2X2 U12 ( .B0(n39), .B1(n6), .A0N(n39), .A1N(n72), .Y(n73) );
  CLKINVX20 U13 ( .A(n41), .Y(n39) );
  CLKINVX1 U14 ( .A(n51), .Y(n44) );
  OAI21X4 U15 ( .A0(n80), .A1(n49), .B0(n79), .Y(n81) );
  INVX4 U16 ( .A(n45), .Y(n49) );
  AOI2BB1X4 U17 ( .A0N(n18), .A1N(n82), .B0(n81), .Y(out[6]) );
  AOI2BB2X1 U18 ( .B0(n39), .B1(n7), .A0N(n40), .A1N(n78), .Y(n80) );
  MX2X2 U19 ( .A(neg_mul[18]), .B(N476), .S0(n88), .Y(out[11]) );
  CLKINVX3 U20 ( .A(in_8bit[7]), .Y(n41) );
  INVX1 U21 ( .A(n97), .Y(n93) );
  INVX4 U22 ( .A(n50), .Y(n18) );
  AOI22X1 U23 ( .A0(N27), .A1(n44), .B0(in_17bit[14]), .B1(n48), .Y(n246) );
  CLKINVX1 U24 ( .A(n83), .Y(n17) );
  NOR2X4 U25 ( .A(n68), .B(n83), .Y(n69) );
  AOI2BB1X4 U26 ( .A0N(n18), .A1N(n75), .B0(n74), .Y(out[5]) );
  NOR2X2 U27 ( .A(n87), .B(n26), .Y(n19) );
  XOR2X4 U28 ( .A(n50), .B(n39), .Y(n83) );
  NOR2BX4 U29 ( .AN(n54), .B(n58), .Y(n60) );
  XOR2X4 U30 ( .A(n60), .B(neg_mul[9]), .Y(out[2]) );
  CLKINVX8 U31 ( .A(n41), .Y(n40) );
  AOI2BB2X2 U32 ( .B0(n71), .B1(n39), .A0N(n39), .A1N(neg_mul[12]), .Y(n75) );
  AOI2BB1X4 U33 ( .A0N(n18), .A1N(n67), .B0(n66), .Y(out[3]) );
  OAI21X4 U34 ( .A0(n73), .A1(n49), .B0(n76), .Y(n74) );
  XNOR2X4 U35 ( .A(n42), .B(n39), .Y(n87) );
  NOR2X2 U36 ( .A(n84), .B(n58), .Y(n85) );
  XNOR2X4 U37 ( .A(n19), .B(n5), .Y(out[9]) );
  INVX8 U38 ( .A(n87), .Y(n88) );
  OAI21X2 U39 ( .A0(n65), .A1(n50), .B0(n64), .Y(n66) );
  INVX8 U40 ( .A(n43), .Y(n42) );
  INVXL U41 ( .A(n44), .Y(n48) );
  INVXL U42 ( .A(n44), .Y(n47) );
  INVX1 U43 ( .A(n207), .Y(in_17bit_b[1]) );
  INVX1 U44 ( .A(n246), .Y(in_17bit_b[14]) );
  INVX1 U45 ( .A(n243), .Y(in_17bit_b[13]) );
  INVX1 U46 ( .A(n210), .Y(in_17bit_b[2]) );
  INVX1 U47 ( .A(n219), .Y(in_17bit_b[5]) );
  INVX1 U48 ( .A(n222), .Y(in_17bit_b[6]) );
  INVX1 U49 ( .A(n225), .Y(in_17bit_b[7]) );
  INVX1 U50 ( .A(n228), .Y(in_17bit_b[8]) );
  INVX1 U51 ( .A(n231), .Y(in_17bit_b[9]) );
  INVX1 U52 ( .A(n234), .Y(in_17bit_b[10]) );
  INVX1 U53 ( .A(n237), .Y(in_17bit_b[11]) );
  INVX1 U54 ( .A(n240), .Y(in_17bit_b[12]) );
  INVX1 U55 ( .A(n216), .Y(in_17bit_b[4]) );
  INVX1 U56 ( .A(n213), .Y(in_17bit_b[3]) );
  INVXL U57 ( .A(in_8bit[0]), .Y(n37) );
  INVXL U58 ( .A(in_8bit[4]), .Y(n36) );
  AOI2BB1X4 U59 ( .A0N(n45), .A1N(n57), .B0(n56), .Y(out[1]) );
  AOI21X1 U60 ( .A0(n20), .A1(n21), .B0(n250), .Y(n203) );
  NOR4XL U61 ( .A(in_8bit[4]), .B(n32), .C(in_8bit[6]), .D(n39), .Y(n20) );
  NOR4XL U62 ( .A(n38), .B(in_8bit[0]), .C(in_8bit[2]), .D(in_8bit[3]), .Y(n21) );
  AND4X1 U63 ( .A(n38), .B(n39), .C(n197), .D(n37), .Y(n22) );
  INVX1 U64 ( .A(n44), .Y(n46) );
  BUFX3 U65 ( .A(in_8bit[1]), .Y(n38) );
  NAND2X1 U66 ( .A(n23), .B(n38), .Y(n89) );
  INVX1 U67 ( .A(n33), .Y(n32) );
  INVX1 U68 ( .A(in_8bit[3]), .Y(n35) );
  NOR3X1 U69 ( .A(n34), .B(n35), .C(n37), .Y(n202) );
  NAND3X1 U70 ( .A(in_8bit[2]), .B(n35), .C(n32), .Y(n198) );
  ADDFX2 U71 ( .A(n31), .B(in_17bit_b[12]), .CI(add_1_root_r112_carry_16_), 
        .CO(add_1_root_r112_carry_17_), .S(add_1_root_r112_SUM_16_) );
  ADDFX2 U72 ( .A(add_1_root_r119_A_19_), .B(in_17bit_b[13]), .CI(
        add_1_root_r119_carry[19]), .CO(add_1_root_r119_carry[20]), .S(
        add_1_root_r119_SUM_19_) );
  ADDFX2 U73 ( .A(n31), .B(in_17bit_b[15]), .CI(add_3_root_r119_carry_17_), 
        .CO(add_3_root_r119_carry_18_), .S(add_1_root_r119_A_17_) );
  ADDFX2 U74 ( .A(n31), .B(in_17bit_b[14]), .CI(add_2_root_r115_carry_17_), 
        .CO(add_2_root_r115_carry_18_), .S(add_2_root_r115_SUM_17_) );
  ADDFX2 U75 ( .A(n31), .B(in_17bit_b[14]), .CI(add_1_root_r115_carry_20_), 
        .CO(add_1_root_r115_carry_21_), .S(add_1_root_r115_SUM_20_) );
  ADDFX2 U76 ( .A(n31), .B(in_17bit_b[15]), .CI(add_2_root_r119_carry_20_), 
        .CO(add_2_root_r119_carry_21_), .S(add_2_root_r119_SUM_20_) );
  AND3X1 U77 ( .A(n39), .B(n36), .C(n33), .Y(n23) );
  NOR2XL U78 ( .A(n39), .B(n36), .Y(n90) );
  ADDFX2 U79 ( .A(in_17bit_b[3]), .B(in_17bit_b[1]), .CI(
        add_2_root_r115_carry_4_), .CO(add_2_root_r115_carry_5_), .S(
        add_2_root_r115_SUM_4_) );
  ADDFX2 U80 ( .A(in_17bit_b[4]), .B(in_17bit_b[2]), .CI(
        add_2_root_r115_carry_5_), .CO(add_2_root_r115_carry_6_), .S(
        add_2_root_r115_SUM_5_) );
  ADDFX2 U81 ( .A(in_17bit_b[5]), .B(in_17bit_b[1]), .CI(
        add_1_root_r112_carry_5_), .CO(add_1_root_r112_carry_6_), .S(
        add_1_root_r112_SUM_5_) );
  ADDFX2 U82 ( .A(in_17bit_b[6]), .B(in_17bit_b[5]), .CI(
        add_3_root_r119_carry_7_), .CO(add_3_root_r119_carry_8_), .S(
        add_1_root_r119_A_7_) );
  ADDFX2 U83 ( .A(in_17bit_b[6]), .B(in_17bit_b[2]), .CI(
        add_1_root_r112_carry_6_), .CO(add_1_root_r112_carry_7_), .S(
        add_1_root_r112_SUM_6_) );
  ADDFX2 U84 ( .A(in_17bit_b[3]), .B(in_17bit_b[1]), .CI(
        add_1_root_r115_carry_7_), .CO(add_1_root_r115_carry_8_), .S(
        add_1_root_r115_SUM_7_) );
  ADDFX2 U85 ( .A(in_17bit_b[7]), .B(in_17bit_b[6]), .CI(
        add_3_root_r119_carry_8_), .CO(add_3_root_r119_carry_9_), .S(
        add_1_root_r119_A_8_) );
  ADDFX2 U86 ( .A(add_1_root_r119_A_7_), .B(in_17bit_b[1]), .CI(
        add_1_root_r119_carry[7]), .CO(add_1_root_r119_carry[8]), .S(
        add_1_root_r119_SUM_7_) );
  ADDFX2 U87 ( .A(in_17bit_b[2]), .B(in_17bit_b[1]), .CI(
        add_2_root_r119_carry_6_), .CO(add_2_root_r119_carry_7_), .S(
        add_2_root_r119_SUM_6_) );
  ADDFX2 U88 ( .A(in_17bit_b[4]), .B(in_17bit_b[2]), .CI(
        add_1_root_r115_carry_8_), .CO(add_1_root_r115_carry_9_), .S(
        add_1_root_r115_SUM_8_) );
  ADDFX2 U89 ( .A(in_17bit_b[8]), .B(in_17bit_b[7]), .CI(
        add_3_root_r119_carry_9_), .CO(add_3_root_r119_carry_10_), .S(
        add_1_root_r119_A_9_) );
  ADDFX2 U90 ( .A(add_1_root_r119_A_8_), .B(in_17bit_b[2]), .CI(
        add_1_root_r119_carry[8]), .CO(add_1_root_r119_carry[9]), .S(
        add_1_root_r119_SUM_8_) );
  ADDFX2 U91 ( .A(in_17bit_b[3]), .B(in_17bit_b[2]), .CI(
        add_2_root_r119_carry_7_), .CO(add_2_root_r119_carry_8_), .S(
        add_2_root_r119_SUM_7_) );
  ADDFX2 U92 ( .A(in_17bit_b[6]), .B(in_17bit_b[4]), .CI(
        add_2_root_r115_carry_7_), .CO(add_2_root_r115_carry_8_), .S(
        add_2_root_r115_SUM_7_) );
  ADDFX2 U93 ( .A(in_17bit_b[8]), .B(in_17bit_b[4]), .CI(
        add_1_root_r112_carry_8_), .CO(add_1_root_r112_carry_9_), .S(
        add_1_root_r112_SUM_8_) );
  ADDFX2 U94 ( .A(in_17bit_b[9]), .B(in_17bit_b[8]), .CI(
        add_3_root_r119_carry_10_), .CO(add_3_root_r119_carry_11_), .S(
        add_1_root_r119_A_10_) );
  ADDFX2 U95 ( .A(in_17bit_b[7]), .B(in_17bit_b[5]), .CI(
        add_2_root_r115_carry_8_), .CO(add_2_root_r115_carry_9_), .S(
        add_2_root_r115_SUM_8_) );
  ADDFX2 U96 ( .A(in_17bit_b[9]), .B(in_17bit_b[5]), .CI(
        add_1_root_r112_carry_9_), .CO(add_1_root_r112_carry_10_), .S(
        add_1_root_r112_SUM_9_) );
  ADDFX2 U97 ( .A(in_17bit_b[10]), .B(in_17bit_b[9]), .CI(
        add_3_root_r119_carry_11_), .CO(add_3_root_r119_carry_12_), .S(
        add_1_root_r119_A_11_) );
  ADDFX2 U98 ( .A(add_1_root_r119_A_10_), .B(in_17bit_b[4]), .CI(
        add_1_root_r119_carry[10]), .CO(add_1_root_r119_carry[11]), .S(
        add_1_root_r119_SUM_10_) );
  ADDFX2 U99 ( .A(in_17bit_b[8]), .B(in_17bit_b[6]), .CI(
        add_2_root_r115_carry_9_), .CO(add_2_root_r115_carry_10_), .S(
        add_2_root_r115_SUM_9_) );
  ADDFX2 U100 ( .A(in_17bit_b[10]), .B(in_17bit_b[6]), .CI(
        add_1_root_r112_carry_10_), .CO(add_1_root_r112_carry_11_), .S(
        add_1_root_r112_SUM_10_) );
  ADDFX2 U101 ( .A(in_17bit_b[7]), .B(in_17bit_b[5]), .CI(
        add_1_root_r115_carry_11_), .CO(add_1_root_r115_carry_12_), .S(
        add_1_root_r115_SUM_11_) );
  ADDFX2 U102 ( .A(in_17bit_b[11]), .B(in_17bit_b[10]), .CI(
        add_3_root_r119_carry_12_), .CO(add_3_root_r119_carry_13_), .S(
        add_1_root_r119_A_12_) );
  ADDFX2 U103 ( .A(add_1_root_r119_A_11_), .B(in_17bit_b[5]), .CI(
        add_1_root_r119_carry[11]), .CO(add_1_root_r119_carry[12]), .S(
        add_1_root_r119_SUM_11_) );
  ADDFX2 U104 ( .A(in_17bit_b[6]), .B(in_17bit_b[5]), .CI(
        add_2_root_r119_carry_10_), .CO(add_2_root_r119_carry_11_), .S(
        add_2_root_r119_SUM_10_) );
  ADDFX2 U105 ( .A(in_17bit_b[9]), .B(in_17bit_b[7]), .CI(
        add_2_root_r115_carry_10_), .CO(add_2_root_r115_carry_11_), .S(
        add_2_root_r115_SUM_10_) );
  ADDFX2 U106 ( .A(in_17bit_b[11]), .B(in_17bit_b[7]), .CI(
        add_1_root_r112_carry_11_), .CO(add_1_root_r112_carry_12_), .S(
        add_1_root_r112_SUM_11_) );
  ADDFX2 U107 ( .A(in_17bit_b[8]), .B(in_17bit_b[6]), .CI(
        add_1_root_r115_carry_12_), .CO(add_1_root_r115_carry_13_), .S(
        add_1_root_r115_SUM_12_) );
  ADDFX2 U108 ( .A(in_17bit_b[12]), .B(in_17bit_b[11]), .CI(
        add_3_root_r119_carry_13_), .CO(add_3_root_r119_carry_14_), .S(
        add_1_root_r119_A_13_) );
  ADDFX2 U109 ( .A(add_1_root_r119_A_12_), .B(in_17bit_b[6]), .CI(
        add_1_root_r119_carry[12]), .CO(add_1_root_r119_carry[13]), .S(
        add_1_root_r119_SUM_12_) );
  ADDFX2 U110 ( .A(in_17bit_b[7]), .B(in_17bit_b[6]), .CI(
        add_2_root_r119_carry_11_), .CO(add_2_root_r119_carry_12_), .S(
        add_2_root_r119_SUM_11_) );
  ADDFX2 U111 ( .A(in_17bit_b[10]), .B(in_17bit_b[8]), .CI(
        add_2_root_r115_carry_11_), .CO(add_2_root_r115_carry_12_), .S(
        add_2_root_r115_SUM_11_) );
  ADDFX2 U112 ( .A(in_17bit_b[12]), .B(in_17bit_b[8]), .CI(
        add_1_root_r112_carry_12_), .CO(add_1_root_r112_carry_13_), .S(
        add_1_root_r112_SUM_12_) );
  ADDFX2 U113 ( .A(in_17bit_b[9]), .B(in_17bit_b[7]), .CI(
        add_1_root_r115_carry_13_), .CO(add_1_root_r115_carry_14_), .S(
        add_1_root_r115_SUM_13_) );
  ADDFX2 U114 ( .A(in_17bit_b[13]), .B(in_17bit_b[12]), .CI(
        add_3_root_r119_carry_14_), .CO(add_3_root_r119_carry_15_), .S(
        add_1_root_r119_A_14_) );
  ADDFX2 U115 ( .A(add_1_root_r119_A_13_), .B(in_17bit_b[7]), .CI(
        add_1_root_r119_carry[13]), .CO(add_1_root_r119_carry[14]), .S(
        add_1_root_r119_SUM_13_) );
  ADDFX2 U116 ( .A(in_17bit_b[8]), .B(in_17bit_b[7]), .CI(
        add_2_root_r119_carry_12_), .CO(add_2_root_r119_carry_13_), .S(
        add_2_root_r119_SUM_12_) );
  ADDFX2 U117 ( .A(in_17bit_b[11]), .B(in_17bit_b[9]), .CI(
        add_2_root_r115_carry_12_), .CO(add_2_root_r115_carry_13_), .S(
        add_2_root_r115_SUM_12_) );
  ADDFX2 U118 ( .A(in_17bit_b[13]), .B(in_17bit_b[9]), .CI(
        add_1_root_r112_carry_13_), .CO(add_1_root_r112_carry_14_), .S(
        add_1_root_r112_SUM_13_) );
  ADDFX2 U119 ( .A(in_17bit_b[10]), .B(in_17bit_b[8]), .CI(
        add_1_root_r115_carry_14_), .CO(add_1_root_r115_carry_15_), .S(
        add_1_root_r115_SUM_14_) );
  ADDFX2 U120 ( .A(in_17bit_b[14]), .B(in_17bit_b[13]), .CI(
        add_3_root_r119_carry_15_), .CO(add_3_root_r119_carry_16_), .S(
        add_1_root_r119_A_15_) );
  ADDFX2 U121 ( .A(add_1_root_r119_A_14_), .B(in_17bit_b[8]), .CI(
        add_1_root_r119_carry[14]), .CO(add_1_root_r119_carry[15]), .S(
        add_1_root_r119_SUM_14_) );
  ADDFX2 U122 ( .A(in_17bit_b[9]), .B(in_17bit_b[8]), .CI(
        add_2_root_r119_carry_13_), .CO(add_2_root_r119_carry_14_), .S(
        add_2_root_r119_SUM_13_) );
  ADDFX2 U123 ( .A(in_17bit_b[12]), .B(in_17bit_b[10]), .CI(
        add_2_root_r115_carry_13_), .CO(add_2_root_r115_carry_14_), .S(
        add_2_root_r115_SUM_13_) );
  ADDFX2 U124 ( .A(in_17bit_b[14]), .B(in_17bit_b[10]), .CI(
        add_1_root_r112_carry_14_), .CO(add_1_root_r112_carry_15_), .S(
        add_1_root_r112_SUM_14_) );
  ADDFX2 U125 ( .A(in_17bit_b[11]), .B(in_17bit_b[9]), .CI(
        add_1_root_r115_carry_15_), .CO(add_1_root_r115_carry_16_), .S(
        add_1_root_r115_SUM_15_) );
  ADDFX2 U126 ( .A(add_1_root_r119_A_15_), .B(in_17bit_b[9]), .CI(
        add_1_root_r119_carry[15]), .CO(add_1_root_r119_carry[16]), .S(
        add_1_root_r119_SUM_15_) );
  ADDFX2 U127 ( .A(in_17bit_b[3]), .B(in_17bit_b[2]), .CI(
        add_3_root_r119_carry_4_), .CO(add_3_root_r119_carry_5_), .S(
        add_1_root_r119_A_4_) );
  ADDFX2 U128 ( .A(in_17bit_b[2]), .B(in_17bit_b[1]), .CI(
        add_3_root_r119_carry_3_), .CO(add_3_root_r119_carry_4_), .S(
        add_1_root_r119_A_3_) );
  ADDFX2 U129 ( .A(in_17bit_b[10]), .B(in_17bit_b[9]), .CI(
        add_2_root_r119_carry_14_), .CO(add_2_root_r119_carry_15_), .S(
        add_2_root_r119_SUM_14_) );
  ADDFX2 U130 ( .A(in_17bit_b[13]), .B(in_17bit_b[11]), .CI(
        add_2_root_r115_carry_14_), .CO(add_2_root_r115_carry_15_), .S(
        add_2_root_r115_SUM_14_) );
  ADDFX2 U131 ( .A(in_17bit_b[15]), .B(in_17bit_b[11]), .CI(
        add_1_root_r112_carry_15_), .CO(add_1_root_r112_carry_16_), .S(
        add_1_root_r112_SUM_15_) );
  ADDFX2 U132 ( .A(in_17bit_b[12]), .B(in_17bit_b[10]), .CI(
        add_1_root_r115_carry_16_), .CO(add_1_root_r115_carry_17_), .S(
        add_1_root_r115_SUM_16_) );
  ADDFX2 U133 ( .A(add_1_root_r119_A_16_), .B(in_17bit_b[10]), .CI(
        add_1_root_r119_carry[16]), .CO(add_1_root_r119_carry[17]), .S(
        add_1_root_r119_SUM_16_) );
  ADDFX2 U134 ( .A(in_17bit_b[11]), .B(in_17bit_b[10]), .CI(
        add_2_root_r119_carry_15_), .CO(add_2_root_r119_carry_16_), .S(
        add_2_root_r119_SUM_15_) );
  ADDFX2 U135 ( .A(in_17bit_b[14]), .B(in_17bit_b[12]), .CI(
        add_2_root_r115_carry_15_), .CO(add_2_root_r115_carry_16_), .S(
        add_2_root_r115_SUM_15_) );
  ADDFX2 U136 ( .A(in_17bit_b[13]), .B(in_17bit_b[11]), .CI(
        add_1_root_r115_carry_17_), .CO(add_1_root_r115_carry_18_), .S(
        add_1_root_r115_SUM_17_) );
  ADDFX2 U137 ( .A(add_1_root_r119_A_17_), .B(in_17bit_b[11]), .CI(
        add_1_root_r119_carry[17]), .CO(add_1_root_r119_carry[18]), .S(
        add_1_root_r119_SUM_17_) );
  ADDFX2 U138 ( .A(in_17bit_b[12]), .B(in_17bit_b[11]), .CI(
        add_2_root_r119_carry_16_), .CO(add_2_root_r119_carry_17_), .S(
        add_2_root_r119_SUM_16_) );
  ADDFX2 U139 ( .A(in_17bit_b[15]), .B(in_17bit_b[13]), .CI(
        add_2_root_r115_carry_16_), .CO(add_2_root_r115_carry_17_), .S(
        add_2_root_r115_SUM_16_) );
  ADDFX2 U140 ( .A(add_1_root_r119_A_18_), .B(in_17bit_b[12]), .CI(
        add_1_root_r119_carry[18]), .CO(add_1_root_r119_carry[19]), .S(
        add_1_root_r119_SUM_18_) );
  ADDFX2 U141 ( .A(in_17bit_b[13]), .B(in_17bit_b[12]), .CI(
        add_2_root_r119_carry_17_), .CO(add_2_root_r119_carry_18_), .S(
        add_2_root_r119_SUM_17_) );
  ADDFX2 U142 ( .A(in_17bit_b[15]), .B(in_17bit_b[13]), .CI(
        add_1_root_r115_carry_19_), .CO(add_1_root_r115_carry_20_), .S(
        add_1_root_r115_SUM_19_) );
  ADDFX2 U143 ( .A(in_17bit_b[7]), .B(in_17bit_b[3]), .CI(
        add_1_root_r112_carry_7_), .CO(add_1_root_r112_carry_8_), .S(
        add_1_root_r112_SUM_7_) );
  ADDFX2 U144 ( .A(in_17bit_b[4]), .B(in_17bit_b[3]), .CI(
        add_2_root_r119_carry_8_), .CO(add_2_root_r119_carry_9_), .S(
        add_2_root_r119_SUM_8_) );
  ADDFX2 U145 ( .A(in_17bit_b[5]), .B(in_17bit_b[4]), .CI(
        add_2_root_r119_carry_9_), .CO(add_2_root_r119_carry_10_), .S(
        add_2_root_r119_SUM_9_) );
  ADDFX2 U146 ( .A(in_17bit_b[14]), .B(in_17bit_b[13]), .CI(
        add_2_root_r119_carry_18_), .CO(add_2_root_r119_carry_19_), .S(
        add_2_root_r119_SUM_18_) );
  ADDFX2 U147 ( .A(in_17bit_b[5]), .B(in_17bit_b[3]), .CI(
        add_2_root_r115_carry_6_), .CO(add_2_root_r115_carry_7_), .S(
        add_2_root_r115_SUM_6_) );
  ADDFX2 U148 ( .A(in_17bit_b[5]), .B(in_17bit_b[3]), .CI(
        add_1_root_r115_carry_9_), .CO(add_1_root_r115_carry_10_), .S(
        add_1_root_r115_SUM_9_) );
  ADDFX2 U149 ( .A(add_1_root_r119_A_9_), .B(in_17bit_b[3]), .CI(
        add_1_root_r119_carry[9]), .CO(add_1_root_r119_carry[10]), .S(
        add_1_root_r119_SUM_9_) );
  ADDFX2 U150 ( .A(in_17bit_b[6]), .B(in_17bit_b[4]), .CI(
        add_1_root_r115_carry_10_), .CO(add_1_root_r115_carry_11_), .S(
        add_1_root_r115_SUM_10_) );
  ADDFX2 U151 ( .A(in_17bit_b[14]), .B(in_17bit_b[12]), .CI(
        add_1_root_r115_carry_18_), .CO(add_1_root_r115_carry_19_), .S(
        add_1_root_r115_SUM_18_) );
  ADDFX2 U152 ( .A(in_17bit_b[15]), .B(in_17bit_b[14]), .CI(
        add_3_root_r119_carry_16_), .CO(add_3_root_r119_carry_17_), .S(
        add_1_root_r119_A_16_) );
  ADDFX2 U153 ( .A(in_17bit_b[4]), .B(in_17bit_b[3]), .CI(
        add_3_root_r119_carry_5_), .CO(add_3_root_r119_carry_6_), .S(
        add_1_root_r119_A_5_) );
  ADDFX2 U154 ( .A(in_17bit_b[5]), .B(in_17bit_b[4]), .CI(
        add_3_root_r119_carry_6_), .CO(add_3_root_r119_carry_7_), .S(
        add_1_root_r119_A_6_) );
  ADDFX2 U155 ( .A(in_17bit_b[15]), .B(in_17bit_b[14]), .CI(
        add_2_root_r119_carry_19_), .CO(add_2_root_r119_carry_20_), .S(
        add_2_root_r119_SUM_19_) );
  BUFX3 U156 ( .A(in_17bit_b[16]), .Y(n31) );
  INVX1 U157 ( .A(n257), .Y(in_17bit_b[16]) );
  INVX1 U158 ( .A(n199), .Y(n96) );
  NAND3BX1 U159 ( .AN(n32), .B(n34), .C(in_8bit[3]), .Y(n199) );
  INVXL U160 ( .A(in_8bit[5]), .Y(n33) );
  CLKINVX3 U161 ( .A(n204), .Y(in_17bit_b[0]) );
  INVX1 U162 ( .A(n177), .Y(n256) );
  NAND2XL U163 ( .A(N29), .B(n18), .Y(n257) );
  INVX1 U164 ( .A(n64), .Y(n68) );
  INVX1 U165 ( .A(n79), .Y(n84) );
  OAI21XL U166 ( .A0(n256), .A1(n257), .B0(n255), .Y(N463) );
  AOI22X1 U167 ( .A0(N221), .A1(n30), .B0(N363), .B1(n29), .Y(n255) );
  CLKINVX3 U168 ( .A(n249), .Y(in_17bit_b[15]) );
  INVX1 U169 ( .A(in_8bit[2]), .Y(n34) );
  AOI22XL U170 ( .A0(N28), .A1(n44), .B0(in_17bit[15]), .B1(n46), .Y(n249) );
  AOI22XL U171 ( .A0(N16), .A1(n44), .B0(in_17bit[3]), .B1(n47), .Y(n213) );
  AOI22XL U172 ( .A0(N17), .A1(n44), .B0(in_17bit[4]), .B1(n46), .Y(n216) );
  AOI22XL U173 ( .A0(N18), .A1(n44), .B0(in_17bit[5]), .B1(n48), .Y(n219) );
  AOI22XL U174 ( .A0(N19), .A1(n44), .B0(in_17bit[6]), .B1(n47), .Y(n222) );
  AOI22XL U175 ( .A0(N20), .A1(n44), .B0(in_17bit[7]), .B1(n46), .Y(n225) );
  AOI22XL U176 ( .A0(N21), .A1(n44), .B0(in_17bit[8]), .B1(n47), .Y(n228) );
  AOI22XL U177 ( .A0(N22), .A1(n44), .B0(in_17bit[9]), .B1(n46), .Y(n231) );
  AOI22XL U178 ( .A0(N23), .A1(n44), .B0(in_17bit[10]), .B1(n46), .Y(n234) );
  AOI22XL U179 ( .A0(N24), .A1(n44), .B0(in_17bit[11]), .B1(n48), .Y(n237) );
  AOI22XL U180 ( .A0(N25), .A1(n44), .B0(in_17bit[12]), .B1(n47), .Y(n240) );
  AOI22XL U181 ( .A0(N26), .A1(n44), .B0(in_17bit[13]), .B1(n47), .Y(n243) );
  AOI22XL U182 ( .A0(in_17bit[0]), .A1(n18), .B0(in_17bit[0]), .B1(n48), .Y(
        n204) );
  AOI22XL U183 ( .A0(N14), .A1(n18), .B0(in_17bit[1]), .B1(n48), .Y(n207) );
  AOI22XL U184 ( .A0(N15), .A1(n18), .B0(in_17bit[2]), .B1(n47), .Y(n210) );
  NAND2BX1 U185 ( .AN(n70), .B(n6), .Y(n76) );
  INVX1 U186 ( .A(n54), .Y(n59) );
  AND2X2 U187 ( .A(n84), .B(n3), .Y(n24) );
  BUFX3 U188 ( .A(n253), .Y(n29) );
  OAI2BB1X1 U189 ( .A0N(n96), .A1N(n22), .B0(n94), .Y(n253) );
  NAND2BX1 U190 ( .AN(n198), .B(n25), .Y(n94) );
  BUFX3 U191 ( .A(n254), .Y(n30) );
  OAI2BB1X1 U192 ( .A0N(n25), .A1N(n96), .B0(n95), .Y(n254) );
  NAND2BX1 U193 ( .AN(n198), .B(n22), .Y(n95) );
  NAND2BX1 U194 ( .AN(n61), .B(n1), .Y(n64) );
  NAND2X1 U195 ( .A(n68), .B(n2), .Y(n70) );
  NAND2BX1 U196 ( .AN(n76), .B(n7), .Y(n79) );
  OAI2BB1X1 U197 ( .A0N(n201), .A1N(n23), .B0(n98), .Y(n177) );
  NAND3BX1 U198 ( .AN(n97), .B(n202), .C(n32), .Y(n98) );
  AND2X2 U199 ( .A(n93), .B(n37), .Y(n25) );
  NAND2X1 U200 ( .A(n59), .B(n16), .Y(n61) );
  AND2X2 U201 ( .A(n24), .B(n4), .Y(n26) );
  INVX1 U202 ( .A(in_17bit[0]), .Y(n99) );
  INVX1 U203 ( .A(in_17bit[13]), .Y(n173) );
  INVX1 U204 ( .A(in_17bit[1]), .Y(n100) );
  INVX1 U205 ( .A(in_17bit[2]), .Y(n101) );
  INVX1 U206 ( .A(in_17bit[3]), .Y(n158) );
  INVX1 U207 ( .A(in_17bit[4]), .Y(n160) );
  INVX1 U208 ( .A(in_17bit[5]), .Y(n161) );
  INVX1 U209 ( .A(in_17bit[6]), .Y(n162) );
  INVX1 U210 ( .A(in_17bit[7]), .Y(n163) );
  INVX1 U211 ( .A(in_17bit[8]), .Y(n164) );
  INVX1 U212 ( .A(in_17bit[9]), .Y(n168) );
  INVX1 U213 ( .A(in_17bit[10]), .Y(n170) );
  INVX1 U214 ( .A(in_17bit[11]), .Y(n171) );
  INVX1 U215 ( .A(in_17bit[12]), .Y(n172) );
  INVX1 U216 ( .A(in_17bit[14]), .Y(n174) );
  INVX1 U217 ( .A(in_17bit[15]), .Y(n175) );
  NAND2X1 U218 ( .A(n206), .B(n205), .Y(N447) );
  AOI22X1 U219 ( .A0(N108), .A1(n250), .B0(N205), .B1(n30), .Y(n205) );
  AOI22X1 U220 ( .A0(N347), .A1(n29), .B0(n177), .B1(in_17bit_b[0]), .Y(n206)
         );
  NAND2X1 U221 ( .A(n209), .B(n208), .Y(N448) );
  AOI22X1 U222 ( .A0(N109), .A1(n250), .B0(N206), .B1(n30), .Y(n208) );
  AOI22X1 U223 ( .A0(N348), .A1(n29), .B0(n177), .B1(n176), .Y(n209) );
  INVX1 U224 ( .A(n207), .Y(n176) );
  NAND2X1 U225 ( .A(n212), .B(n211), .Y(N449) );
  AOI22X1 U226 ( .A0(N110), .A1(n250), .B0(N207), .B1(n30), .Y(n211) );
  AOI22X1 U227 ( .A0(N349), .A1(n29), .B0(n177), .B1(in_17bit_b[2]), .Y(n212)
         );
  NAND2X1 U228 ( .A(n215), .B(n214), .Y(N450) );
  AOI22X1 U229 ( .A0(N111), .A1(n250), .B0(N208), .B1(n30), .Y(n214) );
  AOI22X1 U230 ( .A0(N350), .A1(n29), .B0(n177), .B1(in_17bit_b[3]), .Y(n215)
         );
  NAND2X1 U231 ( .A(n218), .B(n217), .Y(N451) );
  AOI22X1 U232 ( .A0(N112), .A1(n250), .B0(N209), .B1(n30), .Y(n217) );
  AOI22X1 U233 ( .A0(N351), .A1(n29), .B0(n177), .B1(in_17bit_b[4]), .Y(n218)
         );
  NAND2X1 U234 ( .A(n221), .B(n220), .Y(N452) );
  AOI22X1 U235 ( .A0(N113), .A1(n250), .B0(N210), .B1(n30), .Y(n220) );
  AOI22X1 U236 ( .A0(N352), .A1(n29), .B0(n177), .B1(in_17bit_b[5]), .Y(n221)
         );
  NAND2X1 U237 ( .A(n224), .B(n223), .Y(N453) );
  AOI22X1 U238 ( .A0(N114), .A1(n250), .B0(N211), .B1(n30), .Y(n223) );
  AOI22X1 U239 ( .A0(N353), .A1(n29), .B0(n177), .B1(in_17bit_b[6]), .Y(n224)
         );
  NAND2X1 U240 ( .A(n227), .B(n226), .Y(N454) );
  AOI22X1 U241 ( .A0(N115), .A1(n250), .B0(N212), .B1(n30), .Y(n226) );
  AOI22X1 U242 ( .A0(N354), .A1(n29), .B0(n177), .B1(in_17bit_b[7]), .Y(n227)
         );
  NAND2X1 U243 ( .A(n230), .B(n229), .Y(N455) );
  AOI22X1 U244 ( .A0(N116), .A1(n250), .B0(N213), .B1(n30), .Y(n229) );
  AOI22X1 U245 ( .A0(N355), .A1(n29), .B0(n177), .B1(in_17bit_b[8]), .Y(n230)
         );
  NAND2X1 U246 ( .A(n233), .B(n232), .Y(N456) );
  AOI22X1 U247 ( .A0(N117), .A1(n250), .B0(N214), .B1(n30), .Y(n232) );
  AOI22X1 U248 ( .A0(N356), .A1(n29), .B0(n177), .B1(in_17bit_b[9]), .Y(n233)
         );
  NAND2X1 U249 ( .A(n236), .B(n235), .Y(N457) );
  AOI22X1 U250 ( .A0(N118), .A1(n250), .B0(N215), .B1(n30), .Y(n235) );
  AOI22X1 U251 ( .A0(N357), .A1(n29), .B0(n177), .B1(in_17bit_b[10]), .Y(n236)
         );
  NAND2X1 U252 ( .A(n239), .B(n238), .Y(N458) );
  AOI22X1 U253 ( .A0(N119), .A1(n250), .B0(N216), .B1(n30), .Y(n238) );
  AOI22X1 U254 ( .A0(N358), .A1(n29), .B0(n177), .B1(in_17bit_b[11]), .Y(n239)
         );
  NAND2X1 U255 ( .A(n242), .B(n241), .Y(N459) );
  AOI22X1 U256 ( .A0(N120), .A1(n250), .B0(N217), .B1(n30), .Y(n241) );
  AOI22X1 U257 ( .A0(N359), .A1(n29), .B0(n177), .B1(in_17bit_b[12]), .Y(n242)
         );
  NAND2X1 U258 ( .A(n245), .B(n244), .Y(N460) );
  AOI22X1 U259 ( .A0(N121), .A1(n250), .B0(N218), .B1(n30), .Y(n244) );
  AOI22X1 U260 ( .A0(N360), .A1(n29), .B0(n177), .B1(in_17bit_b[13]), .Y(n245)
         );
  NAND2X1 U261 ( .A(n248), .B(n247), .Y(N461) );
  AOI22X1 U262 ( .A0(N122), .A1(n250), .B0(N219), .B1(n30), .Y(n247) );
  AOI22X1 U263 ( .A0(N361), .A1(n29), .B0(n177), .B1(in_17bit_b[14]), .Y(n248)
         );
  NAND2X1 U264 ( .A(n252), .B(n251), .Y(N462) );
  AOI22X1 U265 ( .A0(N123), .A1(n250), .B0(N220), .B1(n30), .Y(n251) );
  AOI22X1 U266 ( .A0(N362), .A1(n29), .B0(n177), .B1(in_17bit_b[15]), .Y(n252)
         );
  INVX1 U267 ( .A(n63), .Y(n62) );
  XNOR2X1 U268 ( .A(n13), .B(sub_add_75_b0_carry[10]), .Y(n27) );
  MX2X2 U269 ( .A(neg_mul[19]), .B(N477), .S0(n88), .Y(out[12]) );
  MX2X4 U270 ( .A(neg_mul[20]), .B(N478), .S0(n88), .Y(out[13]) );
  INVX1 U271 ( .A(n53), .Y(n52) );
  INVX1 U272 ( .A(n72), .Y(n71) );
  AOI2BB2X1 U273 ( .B0(n77), .B1(n39), .A0N(n40), .A1N(neg_mul[13]), .Y(n82)
         );
  INVX1 U274 ( .A(n78), .Y(n77) );
  MX2X1 U275 ( .A(neg_mul[23]), .B(N481), .S0(n17), .Y(out[16]) );
  NAND4BBX1 U276 ( .AN(n29), .BN(n30), .C(n203), .D(n256), .Y(N446) );
  NOR4BX1 U277 ( .AN(n200), .B(n37), .C(n38), .D(in_8bit[2]), .Y(n201) );
  NOR2X1 U278 ( .A(in_8bit[6]), .B(in_8bit[3]), .Y(n200) );
  NAND4BXL U279 ( .AN(n40), .B(n38), .C(in_8bit[4]), .D(in_8bit[6]), .Y(n97)
         );
  NAND2X1 U280 ( .A(n92), .B(n91), .Y(n250) );
  NAND3BX1 U281 ( .AN(n89), .B(n202), .C(in_8bit[6]), .Y(n92) );
  NAND3X1 U282 ( .A(n201), .B(n32), .C(n90), .Y(n91) );
  NOR2X1 U283 ( .A(in_8bit[6]), .B(in_8bit[4]), .Y(n197) );
  NAND2X1 U284 ( .A(neg_mul[13]), .B(n76), .Y(n78) );
  NAND2X1 U285 ( .A(out[0]), .B(neg_mul[8]), .Y(n53) );
  NAND2X1 U286 ( .A(neg_mul[12]), .B(n70), .Y(n72) );
  NAND2X1 U287 ( .A(neg_mul[10]), .B(n61), .Y(n63) );
  OR2X2 U288 ( .A(out[0]), .B(neg_mul[8]), .Y(n54) );
  XNOR2X4 U289 ( .A(n42), .B(n39), .Y(n58) );
  AOI2BB2X4 U290 ( .B0(n62), .B1(n39), .A0N(n40), .A1N(neg_mul[10]), .Y(n67)
         );
  XNOR2X4 U291 ( .A(n69), .B(n2), .Y(out[4]) );
  XNOR2X4 U292 ( .A(n85), .B(n3), .Y(out[7]) );
  NOR2X4 U293 ( .A(n87), .B(n24), .Y(n86) );
  XNOR2X4 U294 ( .A(n86), .B(n4), .Y(out[8]) );
  MXI2X4 U295 ( .A(n13), .B(n27), .S0(n88), .Y(out[10]) );
  AND2X1 U296 ( .A(add_1_root_r112_carry_20_), .B(n31), .Y(
        add_1_root_r112_SUM_21_) );
  XOR2X1 U297 ( .A(n31), .B(add_1_root_r112_carry_20_), .Y(
        add_1_root_r112_SUM_20_) );
  AND2X1 U298 ( .A(add_1_root_r112_carry_19_), .B(in_17bit_b[15]), .Y(
        add_1_root_r112_carry_20_) );
  XOR2X1 U299 ( .A(in_17bit_b[15]), .B(add_1_root_r112_carry_19_), .Y(
        add_1_root_r112_SUM_19_) );
  AND2X1 U300 ( .A(add_1_root_r112_carry_18_), .B(in_17bit_b[14]), .Y(
        add_1_root_r112_carry_19_) );
  XOR2X1 U301 ( .A(in_17bit_b[14]), .B(add_1_root_r112_carry_18_), .Y(
        add_1_root_r112_SUM_18_) );
  AND2X1 U302 ( .A(add_1_root_r112_carry_17_), .B(in_17bit_b[13]), .Y(
        add_1_root_r112_carry_18_) );
  XOR2X1 U303 ( .A(in_17bit_b[13]), .B(add_1_root_r112_carry_17_), .Y(
        add_1_root_r112_SUM_17_) );
  AND2X1 U304 ( .A(add_2_root_r119_carry_21_), .B(n31), .Y(
        add_2_root_r119_SUM_22_) );
  XOR2X1 U305 ( .A(n31), .B(add_2_root_r119_carry_21_), .Y(
        add_2_root_r119_SUM_21_) );
  AND2X1 U306 ( .A(in_17bit_b[1]), .B(in_17bit_b[0]), .Y(
        add_2_root_r119_carry_6_) );
  XOR2X1 U307 ( .A(in_17bit_b[0]), .B(in_17bit_b[1]), .Y(
        add_2_root_r119_SUM_5_) );
  AND2X1 U308 ( .A(add_1_root_r119_carry[22]), .B(n31), .Y(
        add_1_root_r119_SUM_23_) );
  XOR2X1 U309 ( .A(n31), .B(add_1_root_r119_carry[22]), .Y(
        add_1_root_r119_SUM_22_) );
  AND2X1 U310 ( .A(add_1_root_r119_carry[21]), .B(in_17bit_b[15]), .Y(
        add_1_root_r119_carry[22]) );
  XOR2X1 U311 ( .A(in_17bit_b[15]), .B(add_1_root_r119_carry[21]), .Y(
        add_1_root_r119_SUM_21_) );
  AND2X1 U312 ( .A(add_1_root_r119_carry[20]), .B(in_17bit_b[14]), .Y(
        add_1_root_r119_carry[21]) );
  XOR2X1 U313 ( .A(in_17bit_b[14]), .B(add_1_root_r119_carry[20]), .Y(
        add_1_root_r119_SUM_20_) );
  AND2X1 U314 ( .A(add_1_root_r119_A_6_), .B(in_17bit_b[0]), .Y(
        add_1_root_r119_carry[7]) );
  XOR2X1 U315 ( .A(in_17bit_b[0]), .B(add_1_root_r119_A_6_), .Y(
        add_1_root_r119_SUM_6_) );
  AND2X1 U316 ( .A(add_3_root_r119_carry_18_), .B(n31), .Y(
        add_1_root_r119_A_19_) );
  XOR2X1 U317 ( .A(n31), .B(add_3_root_r119_carry_18_), .Y(
        add_1_root_r119_A_18_) );
  AND2X1 U318 ( .A(in_17bit_b[1]), .B(in_17bit_b[0]), .Y(
        add_3_root_r119_carry_3_) );
  XOR2X1 U319 ( .A(in_17bit_b[0]), .B(in_17bit_b[1]), .Y(add_1_root_r119_A_2_)
         );
  AND2X1 U320 ( .A(add_2_root_r115_carry_19_), .B(n31), .Y(
        add_2_root_r115_SUM_20_) );
  XOR2X1 U321 ( .A(n31), .B(add_2_root_r115_carry_19_), .Y(
        add_2_root_r115_SUM_19_) );
  AND2X1 U322 ( .A(add_2_root_r115_carry_18_), .B(in_17bit_b[15]), .Y(
        add_2_root_r115_carry_19_) );
  XOR2X1 U323 ( .A(in_17bit_b[15]), .B(add_2_root_r115_carry_18_), .Y(
        add_2_root_r115_SUM_18_) );
  AND2X1 U324 ( .A(in_17bit_b[2]), .B(in_17bit_b[0]), .Y(
        add_2_root_r115_carry_4_) );
  XOR2X1 U325 ( .A(in_17bit_b[0]), .B(in_17bit_b[2]), .Y(
        add_2_root_r115_SUM_3_) );
  AND2X1 U326 ( .A(add_1_root_r115_carry_22_), .B(n31), .Y(
        add_1_root_r115_SUM_23_) );
  XOR2X1 U327 ( .A(n31), .B(add_1_root_r115_carry_22_), .Y(
        add_1_root_r115_SUM_22_) );
  AND2X1 U328 ( .A(add_1_root_r115_carry_21_), .B(in_17bit_b[15]), .Y(
        add_1_root_r115_carry_22_) );
  XOR2X1 U329 ( .A(in_17bit_b[15]), .B(add_1_root_r115_carry_21_), .Y(
        add_1_root_r115_SUM_21_) );
  AND2X1 U330 ( .A(in_17bit_b[2]), .B(in_17bit_b[0]), .Y(
        add_1_root_r115_carry_7_) );
  XOR2X1 U331 ( .A(in_17bit_b[0]), .B(in_17bit_b[2]), .Y(
        add_1_root_r115_SUM_6_) );
  XOR2X1 U332 ( .A(n51), .B(sub_add_54_b0_carry[16]), .Y(N29) );
  AND2X1 U333 ( .A(sub_add_54_b0_carry[15]), .B(n175), .Y(
        sub_add_54_b0_carry[16]) );
  XOR2X1 U334 ( .A(n175), .B(sub_add_54_b0_carry[15]), .Y(N28) );
  AND2X1 U335 ( .A(sub_add_54_b0_carry[14]), .B(n174), .Y(
        sub_add_54_b0_carry[15]) );
  XOR2X1 U336 ( .A(n174), .B(sub_add_54_b0_carry[14]), .Y(N27) );
  AND2X1 U337 ( .A(sub_add_54_b0_carry[13]), .B(n173), .Y(
        sub_add_54_b0_carry[14]) );
  XOR2X1 U338 ( .A(n173), .B(sub_add_54_b0_carry[13]), .Y(N26) );
  AND2X1 U339 ( .A(sub_add_54_b0_carry[12]), .B(n172), .Y(
        sub_add_54_b0_carry[13]) );
  XOR2X1 U340 ( .A(n172), .B(sub_add_54_b0_carry[12]), .Y(N25) );
  AND2X1 U341 ( .A(sub_add_54_b0_carry[11]), .B(n171), .Y(
        sub_add_54_b0_carry[12]) );
  XOR2X1 U342 ( .A(n171), .B(sub_add_54_b0_carry[11]), .Y(N24) );
  AND2X1 U343 ( .A(sub_add_54_b0_carry[10]), .B(n170), .Y(
        sub_add_54_b0_carry[11]) );
  XOR2X1 U344 ( .A(n170), .B(sub_add_54_b0_carry[10]), .Y(N23) );
  AND2X1 U345 ( .A(sub_add_54_b0_carry[9]), .B(n168), .Y(
        sub_add_54_b0_carry[10]) );
  XOR2X1 U346 ( .A(n168), .B(sub_add_54_b0_carry[9]), .Y(N22) );
  AND2X1 U347 ( .A(sub_add_54_b0_carry[8]), .B(n164), .Y(
        sub_add_54_b0_carry[9]) );
  XOR2X1 U348 ( .A(n164), .B(sub_add_54_b0_carry[8]), .Y(N21) );
  AND2X1 U349 ( .A(sub_add_54_b0_carry[7]), .B(n163), .Y(
        sub_add_54_b0_carry[8]) );
  XOR2X1 U350 ( .A(n163), .B(sub_add_54_b0_carry[7]), .Y(N20) );
  AND2X1 U351 ( .A(sub_add_54_b0_carry[6]), .B(n162), .Y(
        sub_add_54_b0_carry[7]) );
  XOR2X1 U352 ( .A(n162), .B(sub_add_54_b0_carry[6]), .Y(N19) );
  AND2X1 U353 ( .A(sub_add_54_b0_carry[5]), .B(n161), .Y(
        sub_add_54_b0_carry[6]) );
  XOR2X1 U354 ( .A(n161), .B(sub_add_54_b0_carry[5]), .Y(N18) );
  AND2X1 U355 ( .A(sub_add_54_b0_carry[4]), .B(n160), .Y(
        sub_add_54_b0_carry[5]) );
  XOR2X1 U356 ( .A(n160), .B(sub_add_54_b0_carry[4]), .Y(N17) );
  AND2X1 U357 ( .A(sub_add_54_b0_carry[3]), .B(n158), .Y(
        sub_add_54_b0_carry[4]) );
  XOR2X1 U358 ( .A(n158), .B(sub_add_54_b0_carry[3]), .Y(N16) );
  AND2X1 U359 ( .A(sub_add_54_b0_carry[2]), .B(n101), .Y(
        sub_add_54_b0_carry[3]) );
  XOR2X1 U360 ( .A(n101), .B(sub_add_54_b0_carry[2]), .Y(N15) );
  AND2X1 U361 ( .A(n99), .B(n100), .Y(sub_add_54_b0_carry[2]) );
  XOR2X1 U362 ( .A(n100), .B(n99), .Y(N14) );
  XOR2X1 U363 ( .A(n15), .B(sub_add_75_b0_carry[16]), .Y(N481) );
  AND2X1 U364 ( .A(sub_add_75_b0_carry[15]), .B(n8), .Y(
        sub_add_75_b0_carry[16]) );
  XOR2X1 U365 ( .A(n8), .B(sub_add_75_b0_carry[15]), .Y(N480) );
  AND2X1 U366 ( .A(sub_add_75_b0_carry[14]), .B(n9), .Y(
        sub_add_75_b0_carry[15]) );
  XOR2X1 U367 ( .A(n9), .B(sub_add_75_b0_carry[14]), .Y(N479) );
  AND2X1 U368 ( .A(sub_add_75_b0_carry[13]), .B(n10), .Y(
        sub_add_75_b0_carry[14]) );
  XOR2X1 U369 ( .A(n10), .B(sub_add_75_b0_carry[13]), .Y(N478) );
  AND2X1 U370 ( .A(sub_add_75_b0_carry[12]), .B(n12), .Y(
        sub_add_75_b0_carry[13]) );
  XOR2X1 U371 ( .A(n12), .B(sub_add_75_b0_carry[12]), .Y(N477) );
  AND2X1 U372 ( .A(sub_add_75_b0_carry[11]), .B(n11), .Y(
        sub_add_75_b0_carry[12]) );
  XOR2X1 U373 ( .A(n11), .B(sub_add_75_b0_carry[11]), .Y(N476) );
  AND2X1 U374 ( .A(sub_add_75_b0_carry[10]), .B(n13), .Y(
        sub_add_75_b0_carry[11]) );
  AND2X1 U375 ( .A(n26), .B(n5), .Y(sub_add_75_b0_carry[10]) );
  AND2X1 U376 ( .A(in_17bit_b[0]), .B(in_17bit_b[4]), .Y(
        add_1_root_r112_carry_5_) );
endmodule


module multi16_2_DW01_add_0 ( A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, 
        A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, 
        A_4_, B_23_, B_22_, B_21_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, 
        B_14_, B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, 
        SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, 
        SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, 
        SUM_7_ );
  input A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_,
         A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, B_23_, B_22_,
         B_21_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_,
         B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_;
  output SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_,
         SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_,
         SUM_8_, SUM_7_;
  wire   n1, n2, n3, n4;
  wire   [23:7] carry;

  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry[7]), .CO(carry[8]), .S(SUM_7_)
         );
  ADDFX2 U1_21 ( .A(A_21_), .B(B_21_), .CI(carry[21]), .CO(carry[22]), .S(
        SUM_21_) );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry[20]), .CO(carry[21]), .S(
        SUM_20_) );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry[19]), .CO(carry[20]), .S(
        SUM_19_) );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry[18]), .CO(carry[19]), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry[17]), .CO(carry[18]), .S(
        SUM_17_) );
  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry[16]), .CO(carry[17]), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry[15]), .CO(carry[16]), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry[14]), .CO(carry[15]), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry[13]), .CO(carry[14]), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry[12]), .CO(carry[13]), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry[11]), .CO(carry[12]), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry[10]), .CO(carry[11]), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry[9]), .CO(carry[10]), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry[8]), .CO(carry[9]), .S(SUM_8_)
         );
  ADDFX2 U1_22 ( .A(A_22_), .B(B_22_), .CI(carry[22]), .CO(carry[23]), .S(
        SUM_22_) );
  AND2X2 U1 ( .A(A_4_), .B(B_4_), .Y(n1) );
  XOR2X1 U2 ( .A(B_23_), .B(carry[23]), .Y(SUM_23_) );
  OAI2BB1X1 U3 ( .A0N(n2), .A1N(A_6_), .B0(n3), .Y(carry[7]) );
  OAI21XL U4 ( .A0(A_6_), .A1(n2), .B0(B_6_), .Y(n3) );
  OAI2BB1X1 U5 ( .A0N(n1), .A1N(A_5_), .B0(n4), .Y(n2) );
  OAI21XL U6 ( .A0(A_5_), .A1(n1), .B0(B_5_), .Y(n4) );
endmodule


module multi16_2_DW01_add_4 ( A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, 
        A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, 
        B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, 
        B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, SUM_22_, SUM_21_, SUM_20_, 
        SUM_19_, SUM_18_, SUM_17_, SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, 
        SUM_11_, SUM_10_, SUM_9_, SUM_8_, SUM_7_ );
  input A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_,
         A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, B_20_, B_19_,
         B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, B_10_, B_9_,
         B_8_, B_7_, B_6_, B_5_;
  output SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_,
         SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_,
         SUM_7_;
  wire   carry_21_, carry_20_, carry_19_, carry_18_, carry_17_, carry_16_,
         carry_15_, carry_14_, carry_13_, carry_12_, carry_11_, carry_10_,
         carry_9_, carry_8_, carry_7_, n1;

  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry_16_), .CO(carry_17_), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry_15_), .CO(carry_16_), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry_14_), .CO(carry_15_), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry_13_), .CO(carry_14_), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry_12_), .CO(carry_13_), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry_11_), .CO(carry_12_), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry_10_), .CO(carry_11_), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry_9_), .CO(carry_10_), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry_8_), .CO(carry_9_), .S(SUM_8_)
         );
  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry_7_), .CO(carry_8_), .S(SUM_7_)
         );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry_20_), .CO(carry_21_), .S(
        SUM_20_) );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry_19_), .CO(carry_20_), .S(
        SUM_19_) );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry_18_), .CO(carry_19_), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry_17_), .CO(carry_18_), .S(
        SUM_17_) );
  ADDFX2 U1_21 ( .A(A_21_), .B(B_21_), .CI(carry_21_), .CO(SUM_22_), .S(
        SUM_21_) );
  OAI2BB1X1 U1 ( .A0N(A_6_), .A1N(B_6_), .B0(n1), .Y(carry_7_) );
  OAI211X1 U2 ( .A0(B_6_), .A1(A_6_), .B0(A_5_), .C0(B_5_), .Y(n1) );
endmodule


module multi16_2_DW01_add_6 ( A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, 
        A_16_, A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, 
        A_6_, A_5_, A_4_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, 
        B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, 
        SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, 
        SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, 
        SUM_7_ );
  input A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_,
         A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, B_20_,
         B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, B_10_,
         B_9_, B_8_, B_7_, B_6_, B_5_, B_4_;
  output SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_,
         SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_,
         SUM_8_, SUM_7_;
  wire   n1, n2, n3, n4, n5, n6;
  wire   [21:7] carry;

  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry[7]), .CO(carry[8]), .S(SUM_7_)
         );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry[18]), .CO(carry[19]), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry[17]), .CO(carry[18]), .S(
        SUM_17_) );
  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry[16]), .CO(carry[17]), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry[15]), .CO(carry[16]), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry[14]), .CO(carry[15]), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry[13]), .CO(carry[14]), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry[12]), .CO(carry[13]), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry[11]), .CO(carry[12]), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry[10]), .CO(carry[11]), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry[9]), .CO(carry[10]), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry[8]), .CO(carry[9]), .S(SUM_8_)
         );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry[19]), .CO(carry[20]), .S(
        SUM_19_) );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry[20]), .CO(carry[21]), .S(
        SUM_20_) );
  AND2X2 U1 ( .A(A_22_), .B(n2), .Y(n1) );
  AND2X2 U2 ( .A(A_21_), .B(carry[21]), .Y(n2) );
  AND2X2 U3 ( .A(A_4_), .B(B_4_), .Y(n3) );
  XOR2X1 U4 ( .A(A_23_), .B(n1), .Y(SUM_23_) );
  XOR2X1 U5 ( .A(A_21_), .B(carry[21]), .Y(SUM_21_) );
  XOR2X1 U6 ( .A(A_22_), .B(n2), .Y(SUM_22_) );
  OAI2BB1X1 U7 ( .A0N(n4), .A1N(A_6_), .B0(n5), .Y(carry[7]) );
  OAI21XL U8 ( .A0(A_6_), .A1(n4), .B0(B_6_), .Y(n5) );
  OAI2BB1X1 U9 ( .A0N(n3), .A1N(A_5_), .B0(n6), .Y(n4) );
  OAI21XL U10 ( .A0(A_5_), .A1(n3), .B0(B_5_), .Y(n6) );
endmodule


module multi16_2 ( in_17bit, in_8bit, out );
  input [16:0] in_17bit;
  input [7:0] in_8bit;
  output [16:0] out;
  wire   n262, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26,
         N27, N28, N29, N108, N109, N110, N111, N112, N113, N114, N115, N116,
         N117, N118, N119, N120, N121, N122, N123, N205, N206, N207, N208,
         N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, N219,
         N220, N221, N347, N348, N349, N350, N351, N352, N353, N354, N355,
         N356, N357, N358, N359, N360, N361, N362, N363, N446, N447, N448,
         N449, N450, N451, N452, N453, N454, N455, N456, N457, N458, N459,
         N460, N461, N462, N463, N478, N479, N480, N481,
         add_2_root_r119_carry_10_, add_2_root_r119_carry_11_,
         add_2_root_r119_carry_12_, add_2_root_r119_carry_13_,
         add_2_root_r119_carry_14_, add_2_root_r119_carry_15_,
         add_2_root_r119_carry_16_, add_2_root_r119_carry_17_,
         add_2_root_r119_carry_18_, add_2_root_r119_carry_19_,
         add_2_root_r119_carry_20_, add_2_root_r119_carry_21_,
         add_2_root_r119_carry_6_, add_2_root_r119_carry_7_,
         add_2_root_r119_carry_8_, add_2_root_r119_carry_9_,
         add_2_root_r119_SUM_5_, add_2_root_r119_SUM_6_,
         add_2_root_r119_SUM_7_, add_2_root_r119_SUM_8_,
         add_2_root_r119_SUM_9_, add_2_root_r119_SUM_10_,
         add_2_root_r119_SUM_11_, add_2_root_r119_SUM_12_,
         add_2_root_r119_SUM_13_, add_2_root_r119_SUM_14_,
         add_2_root_r119_SUM_15_, add_2_root_r119_SUM_16_,
         add_2_root_r119_SUM_17_, add_2_root_r119_SUM_18_,
         add_2_root_r119_SUM_19_, add_2_root_r119_SUM_20_,
         add_2_root_r119_SUM_21_, add_2_root_r119_SUM_22_,
         add_1_root_r119_SUM_6_, add_1_root_r119_SUM_7_,
         add_1_root_r119_SUM_8_, add_1_root_r119_SUM_9_,
         add_1_root_r119_SUM_10_, add_1_root_r119_SUM_11_,
         add_1_root_r119_SUM_12_, add_1_root_r119_SUM_13_,
         add_1_root_r119_SUM_14_, add_1_root_r119_SUM_15_,
         add_1_root_r119_SUM_16_, add_1_root_r119_SUM_17_,
         add_1_root_r119_SUM_18_, add_1_root_r119_SUM_19_,
         add_1_root_r119_SUM_20_, add_1_root_r119_SUM_21_,
         add_1_root_r119_SUM_22_, add_1_root_r119_SUM_23_,
         add_1_root_r119_A_2_, add_1_root_r119_A_3_, add_1_root_r119_A_4_,
         add_1_root_r119_A_5_, add_1_root_r119_A_6_, add_1_root_r119_A_7_,
         add_1_root_r119_A_8_, add_1_root_r119_A_9_, add_1_root_r119_A_10_,
         add_1_root_r119_A_11_, add_1_root_r119_A_12_, add_1_root_r119_A_13_,
         add_1_root_r119_A_14_, add_1_root_r119_A_15_, add_1_root_r119_A_16_,
         add_1_root_r119_A_17_, add_1_root_r119_A_18_, add_1_root_r119_A_19_,
         add_3_root_r119_carry_10_, add_3_root_r119_carry_11_,
         add_3_root_r119_carry_12_, add_3_root_r119_carry_13_,
         add_3_root_r119_carry_14_, add_3_root_r119_carry_15_,
         add_3_root_r119_carry_16_, add_3_root_r119_carry_17_,
         add_3_root_r119_carry_18_, add_3_root_r119_carry_3_,
         add_3_root_r119_carry_4_, add_3_root_r119_carry_5_,
         add_3_root_r119_carry_6_, add_3_root_r119_carry_7_,
         add_3_root_r119_carry_8_, add_3_root_r119_carry_9_,
         add_1_root_r112_carry_10_, add_1_root_r112_carry_11_,
         add_1_root_r112_carry_12_, add_1_root_r112_carry_13_,
         add_1_root_r112_carry_14_, add_1_root_r112_carry_15_,
         add_1_root_r112_carry_16_, add_1_root_r112_carry_17_,
         add_1_root_r112_carry_18_, add_1_root_r112_carry_19_,
         add_1_root_r112_carry_20_, add_1_root_r112_carry_5_,
         add_1_root_r112_carry_6_, add_1_root_r112_carry_7_,
         add_1_root_r112_carry_8_, add_1_root_r112_carry_9_,
         add_1_root_r112_SUM_1_, add_1_root_r112_SUM_2_,
         add_1_root_r112_SUM_3_, add_1_root_r112_SUM_4_,
         add_1_root_r112_SUM_5_, add_1_root_r112_SUM_6_,
         add_1_root_r112_SUM_7_, add_1_root_r112_SUM_8_,
         add_1_root_r112_SUM_9_, add_1_root_r112_SUM_10_,
         add_1_root_r112_SUM_11_, add_1_root_r112_SUM_12_,
         add_1_root_r112_SUM_13_, add_1_root_r112_SUM_14_,
         add_1_root_r112_SUM_15_, add_1_root_r112_SUM_16_,
         add_1_root_r112_SUM_17_, add_1_root_r112_SUM_18_,
         add_1_root_r112_SUM_19_, add_1_root_r112_SUM_20_,
         add_1_root_r112_SUM_21_, add_2_root_r115_carry_10_,
         add_2_root_r115_carry_11_, add_2_root_r115_carry_12_,
         add_2_root_r115_carry_13_, add_2_root_r115_carry_14_,
         add_2_root_r115_carry_15_, add_2_root_r115_carry_16_,
         add_2_root_r115_carry_17_, add_2_root_r115_carry_18_,
         add_2_root_r115_carry_19_, add_2_root_r115_carry_4_,
         add_2_root_r115_carry_5_, add_2_root_r115_carry_6_,
         add_2_root_r115_carry_7_, add_2_root_r115_carry_8_,
         add_2_root_r115_carry_9_, add_2_root_r115_SUM_3_,
         add_2_root_r115_SUM_4_, add_2_root_r115_SUM_5_,
         add_2_root_r115_SUM_6_, add_2_root_r115_SUM_7_,
         add_2_root_r115_SUM_8_, add_2_root_r115_SUM_9_,
         add_2_root_r115_SUM_10_, add_2_root_r115_SUM_11_,
         add_2_root_r115_SUM_12_, add_2_root_r115_SUM_13_,
         add_2_root_r115_SUM_14_, add_2_root_r115_SUM_15_,
         add_2_root_r115_SUM_16_, add_2_root_r115_SUM_17_,
         add_2_root_r115_SUM_18_, add_2_root_r115_SUM_19_,
         add_2_root_r115_SUM_20_, add_1_root_r115_carry_10_,
         add_1_root_r115_carry_11_, add_1_root_r115_carry_12_,
         add_1_root_r115_carry_13_, add_1_root_r115_carry_14_,
         add_1_root_r115_carry_15_, add_1_root_r115_carry_16_,
         add_1_root_r115_carry_17_, add_1_root_r115_carry_18_,
         add_1_root_r115_carry_19_, add_1_root_r115_carry_20_,
         add_1_root_r115_carry_21_, add_1_root_r115_carry_22_,
         add_1_root_r115_carry_7_, add_1_root_r115_carry_8_,
         add_1_root_r115_carry_9_, add_1_root_r115_SUM_6_,
         add_1_root_r115_SUM_7_, add_1_root_r115_SUM_8_,
         add_1_root_r115_SUM_9_, add_1_root_r115_SUM_10_,
         add_1_root_r115_SUM_11_, add_1_root_r115_SUM_12_,
         add_1_root_r115_SUM_13_, add_1_root_r115_SUM_14_,
         add_1_root_r115_SUM_15_, add_1_root_r115_SUM_16_,
         add_1_root_r115_SUM_17_, add_1_root_r115_SUM_18_,
         add_1_root_r115_SUM_19_, add_1_root_r115_SUM_20_,
         add_1_root_r115_SUM_21_, add_1_root_r115_SUM_22_,
         add_1_root_r115_SUM_23_, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n158, n160, n161, n162, n163, n164, n168, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261;
  wire   [16:0] in_17bit_b;
  wire   [23:8] neg_mul;
  wire   [16:10] sub_add_75_b0_carry;
  wire   [15:2] sub_add_54_b0_carry;
  wire   [22:7] add_1_root_r119_carry;

  multi16_2_DW01_add_0 add_0_root_r119 ( .A_22_(add_2_root_r119_SUM_22_), 
        .A_21_(add_2_root_r119_SUM_21_), .A_20_(add_2_root_r119_SUM_20_), 
        .A_19_(add_2_root_r119_SUM_19_), .A_18_(add_2_root_r119_SUM_18_), 
        .A_17_(add_2_root_r119_SUM_17_), .A_16_(add_2_root_r119_SUM_16_), 
        .A_15_(add_2_root_r119_SUM_15_), .A_14_(add_2_root_r119_SUM_14_), 
        .A_13_(add_2_root_r119_SUM_13_), .A_12_(add_2_root_r119_SUM_12_), 
        .A_11_(add_2_root_r119_SUM_11_), .A_10_(add_2_root_r119_SUM_10_), 
        .A_9_(add_2_root_r119_SUM_9_), .A_8_(add_2_root_r119_SUM_8_), .A_7_(
        add_2_root_r119_SUM_7_), .A_6_(add_2_root_r119_SUM_6_), .A_5_(
        add_2_root_r119_SUM_5_), .A_4_(in_17bit_b[0]), .B_23_(
        add_1_root_r119_SUM_23_), .B_22_(add_1_root_r119_SUM_22_), .B_21_(
        add_1_root_r119_SUM_21_), .B_20_(add_1_root_r119_SUM_20_), .B_19_(
        add_1_root_r119_SUM_19_), .B_18_(add_1_root_r119_SUM_18_), .B_17_(
        add_1_root_r119_SUM_17_), .B_16_(add_1_root_r119_SUM_16_), .B_15_(
        add_1_root_r119_SUM_15_), .B_14_(add_1_root_r119_SUM_14_), .B_13_(
        add_1_root_r119_SUM_13_), .B_12_(add_1_root_r119_SUM_12_), .B_11_(
        add_1_root_r119_SUM_11_), .B_10_(add_1_root_r119_SUM_10_), .B_9_(
        add_1_root_r119_SUM_9_), .B_8_(add_1_root_r119_SUM_8_), .B_7_(
        add_1_root_r119_SUM_7_), .B_6_(add_1_root_r119_SUM_6_), .B_5_(
        add_1_root_r119_A_5_), .B_4_(add_1_root_r119_A_4_), .SUM_23_(N363), 
        .SUM_22_(N362), .SUM_21_(N361), .SUM_20_(N360), .SUM_19_(N359), 
        .SUM_18_(N358), .SUM_17_(N357), .SUM_16_(N356), .SUM_15_(N355), 
        .SUM_14_(N354), .SUM_13_(N353), .SUM_12_(N352), .SUM_11_(N351), 
        .SUM_10_(N350), .SUM_9_(N349), .SUM_8_(N348), .SUM_7_(N347) );
  multi16_2_DW01_add_4 add_0_root_r112 ( .A_21_(n44), .A_20_(in_17bit_b[15]), 
        .A_19_(in_17bit_b[14]), .A_18_(in_17bit_b[13]), .A_17_(in_17bit_b[12]), 
        .A_16_(in_17bit_b[11]), .A_15_(in_17bit_b[10]), .A_14_(in_17bit_b[9]), 
        .A_13_(in_17bit_b[8]), .A_12_(in_17bit_b[7]), .A_11_(in_17bit_b[6]), 
        .A_10_(in_17bit_b[5]), .A_9_(in_17bit_b[4]), .A_8_(in_17bit_b[3]), 
        .A_7_(in_17bit_b[2]), .A_6_(in_17bit_b[1]), .A_5_(in_17bit_b[0]), 
        .B_21_(add_1_root_r112_SUM_21_), .B_20_(add_1_root_r112_SUM_20_), 
        .B_19_(add_1_root_r112_SUM_19_), .B_18_(add_1_root_r112_SUM_18_), 
        .B_17_(add_1_root_r112_SUM_17_), .B_16_(add_1_root_r112_SUM_16_), 
        .B_15_(add_1_root_r112_SUM_15_), .B_14_(add_1_root_r112_SUM_14_), 
        .B_13_(add_1_root_r112_SUM_13_), .B_12_(add_1_root_r112_SUM_12_), 
        .B_11_(add_1_root_r112_SUM_11_), .B_10_(add_1_root_r112_SUM_10_), 
        .B_9_(add_1_root_r112_SUM_9_), .B_8_(add_1_root_r112_SUM_8_), .B_7_(
        add_1_root_r112_SUM_7_), .B_6_(add_1_root_r112_SUM_6_), .B_5_(
        add_1_root_r112_SUM_5_), .SUM_22_(N123), .SUM_21_(N122), .SUM_20_(N121), .SUM_19_(N120), .SUM_18_(N119), .SUM_17_(N118), .SUM_16_(N117), .SUM_15_(
        N116), .SUM_14_(N115), .SUM_13_(N114), .SUM_12_(N113), .SUM_11_(N112), 
        .SUM_10_(N111), .SUM_9_(N110), .SUM_8_(N109), .SUM_7_(N108) );
  multi16_2_DW01_add_6 add_0_root_r115 ( .A_23_(add_1_root_r115_SUM_23_), 
        .A_22_(add_1_root_r115_SUM_22_), .A_21_(add_1_root_r115_SUM_21_), 
        .A_20_(add_1_root_r115_SUM_20_), .A_19_(add_1_root_r115_SUM_19_), 
        .A_18_(add_1_root_r115_SUM_18_), .A_17_(add_1_root_r115_SUM_17_), 
        .A_16_(add_1_root_r115_SUM_16_), .A_15_(add_1_root_r115_SUM_15_), 
        .A_14_(add_1_root_r115_SUM_14_), .A_13_(add_1_root_r115_SUM_13_), 
        .A_12_(add_1_root_r115_SUM_12_), .A_11_(add_1_root_r115_SUM_11_), 
        .A_10_(add_1_root_r115_SUM_10_), .A_9_(add_1_root_r115_SUM_9_), .A_8_(
        add_1_root_r115_SUM_8_), .A_7_(add_1_root_r115_SUM_7_), .A_6_(
        add_1_root_r115_SUM_6_), .A_5_(in_17bit_b[1]), .A_4_(in_17bit_b[0]), 
        .B_20_(add_2_root_r115_SUM_20_), .B_19_(add_2_root_r115_SUM_19_), 
        .B_18_(add_2_root_r115_SUM_18_), .B_17_(add_2_root_r115_SUM_17_), 
        .B_16_(add_2_root_r115_SUM_16_), .B_15_(add_2_root_r115_SUM_15_), 
        .B_14_(add_2_root_r115_SUM_14_), .B_13_(add_2_root_r115_SUM_13_), 
        .B_12_(add_2_root_r115_SUM_12_), .B_11_(add_2_root_r115_SUM_11_), 
        .B_10_(add_2_root_r115_SUM_10_), .B_9_(add_2_root_r115_SUM_9_), .B_8_(
        add_2_root_r115_SUM_8_), .B_7_(add_2_root_r115_SUM_7_), .B_6_(
        add_2_root_r115_SUM_6_), .B_5_(add_2_root_r115_SUM_5_), .B_4_(
        add_2_root_r115_SUM_4_), .SUM_23_(N221), .SUM_22_(N220), .SUM_21_(N219), .SUM_20_(N218), .SUM_19_(N217), .SUM_18_(N216), .SUM_17_(N215), .SUM_16_(
        N214), .SUM_15_(N213), .SUM_14_(N212), .SUM_13_(N211), .SUM_12_(N210), 
        .SUM_11_(N209), .SUM_10_(N208), .SUM_9_(N207), .SUM_8_(N206), .SUM_7_(
        N205) );
  TLATX1 neg_mul_reg_16_ ( .G(N446), .D(N456), .QN(n6) );
  TLATX1 neg_mul_reg_15_ ( .G(N446), .D(N455), .Q(n2), .QN(n13) );
  TLATX1 neg_mul_reg_14_ ( .G(N446), .D(N454), .QN(n5) );
  TLATX1 neg_mul_reg_13_ ( .G(N446), .D(N453), .Q(neg_mul[13]), .QN(n3) );
  TLATX1 neg_mul_reg_12_ ( .G(N446), .D(N452), .QN(n4) );
  TLATX1 neg_mul_reg_11_ ( .G(N446), .D(N451), .Q(neg_mul[11]), .QN(n18) );
  TLATX1 neg_mul_reg_23_ ( .G(N446), .D(N463), .Q(neg_mul[23]), .QN(n17) );
  TLATX1 neg_mul_reg_22_ ( .G(N446), .D(N462), .Q(neg_mul[22]), .QN(n11) );
  TLATX1 neg_mul_reg_21_ ( .G(N446), .D(N461), .Q(neg_mul[21]), .QN(n12) );
  TLATX1 neg_mul_reg_20_ ( .G(N446), .D(N460), .Q(neg_mul[20]), .QN(n9) );
  TLATX1 neg_mul_reg_19_ ( .G(N446), .D(N459), .Q(neg_mul[19]), .QN(n10) );
  TLATX1 neg_mul_reg_18_ ( .G(N446), .D(N458), .QN(n15) );
  TLATX1 neg_mul_reg_17_ ( .G(N446), .D(N457), .QN(n14) );
  TLATX1 neg_mul_reg_9_ ( .G(N446), .D(N449), .Q(neg_mul[9]), .QN(n8) );
  TLATX1 neg_mul_reg_10_ ( .G(N446), .D(N450), .Q(neg_mul[10]), .QN(n7) );
  TLATX1 neg_mul_reg_8_ ( .G(N446), .D(N448), .Q(neg_mul[8]), .QN(n16) );
  TLATX1 neg_mul_reg_7_ ( .G(N446), .D(N447), .Q(out[0]) );
  OAI21X4 U2 ( .A0(n80), .A1(n61), .B0(n79), .Y(n81) );
  MXI2X4 U3 ( .A(n15), .B(n40), .S0(n92), .Y(out[11]) );
  AOI2BB2X1 U4 ( .B0(n77), .B1(n51), .A0N(n52), .A1N(neg_mul[10]), .Y(n82) );
  INVX3 U5 ( .A(n53), .Y(n52) );
  INVX12 U6 ( .A(n86), .Y(n92) );
  CLKINVX3 U7 ( .A(n55), .Y(n62) );
  INVX4 U8 ( .A(n58), .Y(n61) );
  NAND2X2 U9 ( .A(n55), .B(n51), .Y(n22) );
  CLKINVX8 U10 ( .A(n56), .Y(n55) );
  OAI21X4 U11 ( .A0(n67), .A1(n62), .B0(n66), .Y(n68) );
  AOI2BB2X2 U12 ( .B0(n51), .B1(n7), .A0N(n52), .A1N(n78), .Y(n80) );
  AOI2BB2X2 U13 ( .B0(n51), .B1(n8), .A0N(n52), .A1N(n72), .Y(n73) );
  INVX20 U14 ( .A(n53), .Y(n51) );
  BUFX4 U15 ( .A(n262), .Y(out[12]) );
  AOI2BB2X2 U16 ( .B0(n51), .B1(n16), .A0N(n51), .A1N(n65), .Y(n67) );
  MXI2X4 U17 ( .A(n14), .B(n39), .S0(n92), .Y(out[10]) );
  NAND2X2 U18 ( .A(n20), .B(n21), .Y(n23) );
  CLKINVX3 U19 ( .A(n58), .Y(n20) );
  MX2X1 U20 ( .A(n25), .B(neg_mul[19]), .S0(n86), .Y(n262) );
  INVX2 U21 ( .A(in_8bit[7]), .Y(n53) );
  INVX1 U22 ( .A(n101), .Y(n97) );
  XOR2X4 U23 ( .A(n85), .B(neg_mul[11]), .Y(out[4]) );
  OR2X2 U24 ( .A(n86), .B(n38), .Y(n32) );
  INVX3 U25 ( .A(n51), .Y(n19) );
  AOI2BB2X1 U26 ( .B0(n71), .B1(n51), .A0N(n52), .A1N(neg_mul[9]), .Y(n75) );
  NAND2X4 U27 ( .A(n23), .B(n22), .Y(n88) );
  CLKINVX8 U28 ( .A(in_17bit[16]), .Y(n56) );
  XOR2X4 U29 ( .A(n58), .B(n19), .Y(n86) );
  INVXL U30 ( .A(n56), .Y(n54) );
  INVX1 U31 ( .A(n51), .Y(n21) );
  AOI2BB2X1 U32 ( .B0(n64), .B1(n51), .A0N(n52), .A1N(neg_mul[8]), .Y(n69) );
  XOR2X4 U33 ( .A(n89), .B(neg_mul[13]), .Y(out[6]) );
  XOR2X4 U34 ( .A(n32), .B(n6), .Y(out[9]) );
  XNOR2X2 U35 ( .A(n58), .B(n51), .Y(n83) );
  MX2X4 U36 ( .A(neg_mul[20]), .B(N478), .S0(n92), .Y(out[13]) );
  NOR2X2 U37 ( .A(n86), .B(n36), .Y(n24) );
  XNOR2X1 U38 ( .A(n55), .B(n51), .Y(n90) );
  INVX8 U39 ( .A(n56), .Y(n58) );
  NOR2X4 U40 ( .A(n35), .B(n90), .Y(n91) );
  NOR2X4 U41 ( .A(n84), .B(n83), .Y(n85) );
  NOR2X4 U42 ( .A(n34), .B(n88), .Y(n89) );
  INVX1 U43 ( .A(n211), .Y(in_17bit_b[1]) );
  INVX1 U44 ( .A(n250), .Y(in_17bit_b[14]) );
  INVX1 U45 ( .A(n247), .Y(in_17bit_b[13]) );
  INVX1 U46 ( .A(n214), .Y(in_17bit_b[2]) );
  INVX1 U47 ( .A(n223), .Y(in_17bit_b[5]) );
  INVX1 U48 ( .A(n226), .Y(in_17bit_b[6]) );
  INVX1 U49 ( .A(n232), .Y(in_17bit_b[8]) );
  INVX1 U50 ( .A(n235), .Y(in_17bit_b[9]) );
  INVX1 U51 ( .A(n229), .Y(in_17bit_b[7]) );
  INVX1 U52 ( .A(n238), .Y(in_17bit_b[10]) );
  INVX1 U53 ( .A(n241), .Y(in_17bit_b[11]) );
  INVX1 U54 ( .A(n244), .Y(in_17bit_b[12]) );
  INVX1 U55 ( .A(n220), .Y(in_17bit_b[4]) );
  INVX1 U56 ( .A(n217), .Y(in_17bit_b[3]) );
  INVXL U57 ( .A(in_8bit[0]), .Y(n49) );
  INVXL U58 ( .A(in_8bit[4]), .Y(n48) );
  XOR2X4 U59 ( .A(n24), .B(n2), .Y(out[8]) );
  XOR2X1 U60 ( .A(n10), .B(sub_add_75_b0_carry[12]), .Y(n25) );
  AOI21X1 U61 ( .A0(n27), .A1(n28), .B0(n254), .Y(n207) );
  NOR4XL U62 ( .A(in_8bit[4]), .B(in_8bit[5]), .C(in_8bit[6]), .D(n51), .Y(n27) );
  NOR4XL U63 ( .A(n50), .B(in_8bit[0]), .C(in_8bit[2]), .D(in_8bit[3]), .Y(n28) );
  AND4X1 U64 ( .A(n50), .B(n51), .C(n201), .D(n49), .Y(n29) );
  INVX1 U65 ( .A(n63), .Y(n57) );
  BUFX3 U66 ( .A(in_8bit[1]), .Y(n50) );
  NAND2X1 U67 ( .A(n30), .B(n50), .Y(n93) );
  INVX1 U68 ( .A(in_8bit[3]), .Y(n47) );
  NOR3X1 U69 ( .A(n46), .B(n47), .C(n49), .Y(n206) );
  NAND3X1 U70 ( .A(in_8bit[2]), .B(n47), .C(in_8bit[5]), .Y(n202) );
  ADDFX2 U71 ( .A(n44), .B(in_17bit_b[12]), .CI(add_1_root_r112_carry_16_), 
        .CO(add_1_root_r112_carry_17_), .S(add_1_root_r112_SUM_16_) );
  ADDFX2 U72 ( .A(add_1_root_r119_A_19_), .B(in_17bit_b[13]), .CI(
        add_1_root_r119_carry[19]), .CO(add_1_root_r119_carry[20]), .S(
        add_1_root_r119_SUM_19_) );
  ADDFX2 U73 ( .A(n44), .B(in_17bit_b[15]), .CI(add_3_root_r119_carry_17_), 
        .CO(add_3_root_r119_carry_18_), .S(add_1_root_r119_A_17_) );
  ADDFX2 U74 ( .A(n44), .B(in_17bit_b[14]), .CI(add_2_root_r115_carry_17_), 
        .CO(add_2_root_r115_carry_18_), .S(add_2_root_r115_SUM_17_) );
  ADDFX2 U75 ( .A(n44), .B(in_17bit_b[14]), .CI(add_1_root_r115_carry_20_), 
        .CO(add_1_root_r115_carry_21_), .S(add_1_root_r115_SUM_20_) );
  ADDFX2 U76 ( .A(n44), .B(in_17bit_b[15]), .CI(add_2_root_r119_carry_20_), 
        .CO(add_2_root_r119_carry_21_), .S(add_2_root_r119_SUM_20_) );
  AND3X1 U77 ( .A(n51), .B(n48), .C(n45), .Y(n30) );
  NOR2XL U78 ( .A(n51), .B(n48), .Y(n94) );
  ADDFX2 U79 ( .A(in_17bit_b[3]), .B(in_17bit_b[1]), .CI(
        add_2_root_r115_carry_4_), .CO(add_2_root_r115_carry_5_), .S(
        add_2_root_r115_SUM_4_) );
  ADDFX2 U80 ( .A(in_17bit_b[4]), .B(in_17bit_b[2]), .CI(
        add_2_root_r115_carry_5_), .CO(add_2_root_r115_carry_6_), .S(
        add_2_root_r115_SUM_5_) );
  ADDFX2 U81 ( .A(in_17bit_b[5]), .B(in_17bit_b[1]), .CI(
        add_1_root_r112_carry_5_), .CO(add_1_root_r112_carry_6_), .S(
        add_1_root_r112_SUM_5_) );
  ADDFX2 U82 ( .A(in_17bit_b[6]), .B(in_17bit_b[5]), .CI(
        add_3_root_r119_carry_7_), .CO(add_3_root_r119_carry_8_), .S(
        add_1_root_r119_A_7_) );
  ADDFX2 U83 ( .A(in_17bit_b[6]), .B(in_17bit_b[2]), .CI(
        add_1_root_r112_carry_6_), .CO(add_1_root_r112_carry_7_), .S(
        add_1_root_r112_SUM_6_) );
  ADDFX2 U84 ( .A(in_17bit_b[3]), .B(in_17bit_b[1]), .CI(
        add_1_root_r115_carry_7_), .CO(add_1_root_r115_carry_8_), .S(
        add_1_root_r115_SUM_7_) );
  ADDFX2 U85 ( .A(in_17bit_b[7]), .B(in_17bit_b[6]), .CI(
        add_3_root_r119_carry_8_), .CO(add_3_root_r119_carry_9_), .S(
        add_1_root_r119_A_8_) );
  ADDFX2 U86 ( .A(add_1_root_r119_A_7_), .B(in_17bit_b[1]), .CI(
        add_1_root_r119_carry[7]), .CO(add_1_root_r119_carry[8]), .S(
        add_1_root_r119_SUM_7_) );
  ADDFX2 U87 ( .A(in_17bit_b[2]), .B(in_17bit_b[1]), .CI(
        add_2_root_r119_carry_6_), .CO(add_2_root_r119_carry_7_), .S(
        add_2_root_r119_SUM_6_) );
  ADDFX2 U88 ( .A(in_17bit_b[4]), .B(in_17bit_b[2]), .CI(
        add_1_root_r115_carry_8_), .CO(add_1_root_r115_carry_9_), .S(
        add_1_root_r115_SUM_8_) );
  ADDFX2 U89 ( .A(in_17bit_b[8]), .B(in_17bit_b[7]), .CI(
        add_3_root_r119_carry_9_), .CO(add_3_root_r119_carry_10_), .S(
        add_1_root_r119_A_9_) );
  ADDFX2 U90 ( .A(add_1_root_r119_A_8_), .B(in_17bit_b[2]), .CI(
        add_1_root_r119_carry[8]), .CO(add_1_root_r119_carry[9]), .S(
        add_1_root_r119_SUM_8_) );
  ADDFX2 U91 ( .A(in_17bit_b[3]), .B(in_17bit_b[2]), .CI(
        add_2_root_r119_carry_7_), .CO(add_2_root_r119_carry_8_), .S(
        add_2_root_r119_SUM_7_) );
  ADDFX2 U92 ( .A(in_17bit_b[6]), .B(in_17bit_b[4]), .CI(
        add_2_root_r115_carry_7_), .CO(add_2_root_r115_carry_8_), .S(
        add_2_root_r115_SUM_7_) );
  ADDFX2 U93 ( .A(in_17bit_b[8]), .B(in_17bit_b[4]), .CI(
        add_1_root_r112_carry_8_), .CO(add_1_root_r112_carry_9_), .S(
        add_1_root_r112_SUM_8_) );
  ADDFX2 U94 ( .A(in_17bit_b[9]), .B(in_17bit_b[8]), .CI(
        add_3_root_r119_carry_10_), .CO(add_3_root_r119_carry_11_), .S(
        add_1_root_r119_A_10_) );
  ADDFX2 U95 ( .A(in_17bit_b[7]), .B(in_17bit_b[5]), .CI(
        add_2_root_r115_carry_8_), .CO(add_2_root_r115_carry_9_), .S(
        add_2_root_r115_SUM_8_) );
  ADDFX2 U96 ( .A(in_17bit_b[9]), .B(in_17bit_b[5]), .CI(
        add_1_root_r112_carry_9_), .CO(add_1_root_r112_carry_10_), .S(
        add_1_root_r112_SUM_9_) );
  ADDFX2 U97 ( .A(in_17bit_b[6]), .B(in_17bit_b[4]), .CI(
        add_1_root_r115_carry_10_), .CO(add_1_root_r115_carry_11_), .S(
        add_1_root_r115_SUM_10_) );
  ADDFX2 U98 ( .A(in_17bit_b[10]), .B(in_17bit_b[9]), .CI(
        add_3_root_r119_carry_11_), .CO(add_3_root_r119_carry_12_), .S(
        add_1_root_r119_A_11_) );
  ADDFX2 U99 ( .A(add_1_root_r119_A_10_), .B(in_17bit_b[4]), .CI(
        add_1_root_r119_carry[10]), .CO(add_1_root_r119_carry[11]), .S(
        add_1_root_r119_SUM_10_) );
  ADDFX2 U100 ( .A(in_17bit_b[5]), .B(in_17bit_b[4]), .CI(
        add_2_root_r119_carry_9_), .CO(add_2_root_r119_carry_10_), .S(
        add_2_root_r119_SUM_9_) );
  ADDFX2 U101 ( .A(in_17bit_b[8]), .B(in_17bit_b[6]), .CI(
        add_2_root_r115_carry_9_), .CO(add_2_root_r115_carry_10_), .S(
        add_2_root_r115_SUM_9_) );
  ADDFX2 U102 ( .A(in_17bit_b[10]), .B(in_17bit_b[6]), .CI(
        add_1_root_r112_carry_10_), .CO(add_1_root_r112_carry_11_), .S(
        add_1_root_r112_SUM_10_) );
  ADDFX2 U103 ( .A(in_17bit_b[7]), .B(in_17bit_b[5]), .CI(
        add_1_root_r115_carry_11_), .CO(add_1_root_r115_carry_12_), .S(
        add_1_root_r115_SUM_11_) );
  ADDFX2 U104 ( .A(in_17bit_b[11]), .B(in_17bit_b[10]), .CI(
        add_3_root_r119_carry_12_), .CO(add_3_root_r119_carry_13_), .S(
        add_1_root_r119_A_12_) );
  ADDFX2 U105 ( .A(add_1_root_r119_A_11_), .B(in_17bit_b[5]), .CI(
        add_1_root_r119_carry[11]), .CO(add_1_root_r119_carry[12]), .S(
        add_1_root_r119_SUM_11_) );
  ADDFX2 U106 ( .A(in_17bit_b[6]), .B(in_17bit_b[5]), .CI(
        add_2_root_r119_carry_10_), .CO(add_2_root_r119_carry_11_), .S(
        add_2_root_r119_SUM_10_) );
  ADDFX2 U107 ( .A(in_17bit_b[9]), .B(in_17bit_b[7]), .CI(
        add_2_root_r115_carry_10_), .CO(add_2_root_r115_carry_11_), .S(
        add_2_root_r115_SUM_10_) );
  ADDFX2 U108 ( .A(in_17bit_b[11]), .B(in_17bit_b[7]), .CI(
        add_1_root_r112_carry_11_), .CO(add_1_root_r112_carry_12_), .S(
        add_1_root_r112_SUM_11_) );
  ADDFX2 U109 ( .A(in_17bit_b[8]), .B(in_17bit_b[6]), .CI(
        add_1_root_r115_carry_12_), .CO(add_1_root_r115_carry_13_), .S(
        add_1_root_r115_SUM_12_) );
  ADDFX2 U110 ( .A(in_17bit_b[12]), .B(in_17bit_b[11]), .CI(
        add_3_root_r119_carry_13_), .CO(add_3_root_r119_carry_14_), .S(
        add_1_root_r119_A_13_) );
  ADDFX2 U111 ( .A(add_1_root_r119_A_12_), .B(in_17bit_b[6]), .CI(
        add_1_root_r119_carry[12]), .CO(add_1_root_r119_carry[13]), .S(
        add_1_root_r119_SUM_12_) );
  ADDFX2 U112 ( .A(in_17bit_b[7]), .B(in_17bit_b[6]), .CI(
        add_2_root_r119_carry_11_), .CO(add_2_root_r119_carry_12_), .S(
        add_2_root_r119_SUM_11_) );
  ADDFX2 U113 ( .A(in_17bit_b[10]), .B(in_17bit_b[8]), .CI(
        add_2_root_r115_carry_11_), .CO(add_2_root_r115_carry_12_), .S(
        add_2_root_r115_SUM_11_) );
  ADDFX2 U114 ( .A(in_17bit_b[12]), .B(in_17bit_b[8]), .CI(
        add_1_root_r112_carry_12_), .CO(add_1_root_r112_carry_13_), .S(
        add_1_root_r112_SUM_12_) );
  ADDFX2 U115 ( .A(in_17bit_b[9]), .B(in_17bit_b[7]), .CI(
        add_1_root_r115_carry_13_), .CO(add_1_root_r115_carry_14_), .S(
        add_1_root_r115_SUM_13_) );
  ADDFX2 U116 ( .A(in_17bit_b[13]), .B(in_17bit_b[12]), .CI(
        add_3_root_r119_carry_14_), .CO(add_3_root_r119_carry_15_), .S(
        add_1_root_r119_A_14_) );
  ADDFX2 U117 ( .A(add_1_root_r119_A_13_), .B(in_17bit_b[7]), .CI(
        add_1_root_r119_carry[13]), .CO(add_1_root_r119_carry[14]), .S(
        add_1_root_r119_SUM_13_) );
  ADDFX2 U118 ( .A(in_17bit_b[8]), .B(in_17bit_b[7]), .CI(
        add_2_root_r119_carry_12_), .CO(add_2_root_r119_carry_13_), .S(
        add_2_root_r119_SUM_12_) );
  ADDFX2 U119 ( .A(in_17bit_b[11]), .B(in_17bit_b[9]), .CI(
        add_2_root_r115_carry_12_), .CO(add_2_root_r115_carry_13_), .S(
        add_2_root_r115_SUM_12_) );
  ADDFX2 U120 ( .A(in_17bit_b[13]), .B(in_17bit_b[9]), .CI(
        add_1_root_r112_carry_13_), .CO(add_1_root_r112_carry_14_), .S(
        add_1_root_r112_SUM_13_) );
  ADDFX2 U121 ( .A(in_17bit_b[10]), .B(in_17bit_b[8]), .CI(
        add_1_root_r115_carry_14_), .CO(add_1_root_r115_carry_15_), .S(
        add_1_root_r115_SUM_14_) );
  ADDFX2 U122 ( .A(add_1_root_r119_A_14_), .B(in_17bit_b[8]), .CI(
        add_1_root_r119_carry[14]), .CO(add_1_root_r119_carry[15]), .S(
        add_1_root_r119_SUM_14_) );
  ADDFX2 U123 ( .A(in_17bit_b[9]), .B(in_17bit_b[8]), .CI(
        add_2_root_r119_carry_13_), .CO(add_2_root_r119_carry_14_), .S(
        add_2_root_r119_SUM_13_) );
  ADDFX2 U124 ( .A(in_17bit_b[12]), .B(in_17bit_b[10]), .CI(
        add_2_root_r115_carry_13_), .CO(add_2_root_r115_carry_14_), .S(
        add_2_root_r115_SUM_13_) );
  ADDFX2 U125 ( .A(in_17bit_b[14]), .B(in_17bit_b[10]), .CI(
        add_1_root_r112_carry_14_), .CO(add_1_root_r112_carry_15_), .S(
        add_1_root_r112_SUM_14_) );
  ADDFX2 U126 ( .A(in_17bit_b[11]), .B(in_17bit_b[9]), .CI(
        add_1_root_r115_carry_15_), .CO(add_1_root_r115_carry_16_), .S(
        add_1_root_r115_SUM_15_) );
  ADDFX2 U127 ( .A(add_1_root_r119_A_15_), .B(in_17bit_b[9]), .CI(
        add_1_root_r119_carry[15]), .CO(add_1_root_r119_carry[16]), .S(
        add_1_root_r119_SUM_15_) );
  ADDFX2 U128 ( .A(in_17bit_b[10]), .B(in_17bit_b[9]), .CI(
        add_2_root_r119_carry_14_), .CO(add_2_root_r119_carry_15_), .S(
        add_2_root_r119_SUM_14_) );
  ADDFX2 U129 ( .A(in_17bit_b[13]), .B(in_17bit_b[11]), .CI(
        add_2_root_r115_carry_14_), .CO(add_2_root_r115_carry_15_), .S(
        add_2_root_r115_SUM_14_) );
  ADDFX2 U130 ( .A(in_17bit_b[15]), .B(in_17bit_b[11]), .CI(
        add_1_root_r112_carry_15_), .CO(add_1_root_r112_carry_16_), .S(
        add_1_root_r112_SUM_15_) );
  ADDFX2 U131 ( .A(in_17bit_b[12]), .B(in_17bit_b[10]), .CI(
        add_1_root_r115_carry_16_), .CO(add_1_root_r115_carry_17_), .S(
        add_1_root_r115_SUM_16_) );
  ADDFX2 U132 ( .A(add_1_root_r119_A_16_), .B(in_17bit_b[10]), .CI(
        add_1_root_r119_carry[16]), .CO(add_1_root_r119_carry[17]), .S(
        add_1_root_r119_SUM_16_) );
  ADDFX2 U133 ( .A(in_17bit_b[11]), .B(in_17bit_b[10]), .CI(
        add_2_root_r119_carry_15_), .CO(add_2_root_r119_carry_16_), .S(
        add_2_root_r119_SUM_15_) );
  ADDFX2 U134 ( .A(in_17bit_b[14]), .B(in_17bit_b[12]), .CI(
        add_2_root_r115_carry_15_), .CO(add_2_root_r115_carry_16_), .S(
        add_2_root_r115_SUM_15_) );
  ADDFX2 U135 ( .A(in_17bit_b[13]), .B(in_17bit_b[11]), .CI(
        add_1_root_r115_carry_17_), .CO(add_1_root_r115_carry_18_), .S(
        add_1_root_r115_SUM_17_) );
  ADDFX2 U136 ( .A(add_1_root_r119_A_17_), .B(in_17bit_b[11]), .CI(
        add_1_root_r119_carry[17]), .CO(add_1_root_r119_carry[18]), .S(
        add_1_root_r119_SUM_17_) );
  ADDFX2 U137 ( .A(in_17bit_b[12]), .B(in_17bit_b[11]), .CI(
        add_2_root_r119_carry_16_), .CO(add_2_root_r119_carry_17_), .S(
        add_2_root_r119_SUM_16_) );
  ADDFX2 U138 ( .A(in_17bit_b[14]), .B(in_17bit_b[12]), .CI(
        add_1_root_r115_carry_18_), .CO(add_1_root_r115_carry_19_), .S(
        add_1_root_r115_SUM_18_) );
  ADDFX2 U139 ( .A(in_17bit_b[5]), .B(in_17bit_b[3]), .CI(
        add_2_root_r115_carry_6_), .CO(add_2_root_r115_carry_7_), .S(
        add_2_root_r115_SUM_6_) );
  ADDFX2 U140 ( .A(add_1_root_r119_A_9_), .B(in_17bit_b[3]), .CI(
        add_1_root_r119_carry[9]), .CO(add_1_root_r119_carry[10]), .S(
        add_1_root_r119_SUM_9_) );
  ADDFX2 U141 ( .A(in_17bit_b[13]), .B(in_17bit_b[12]), .CI(
        add_2_root_r119_carry_17_), .CO(add_2_root_r119_carry_18_), .S(
        add_2_root_r119_SUM_17_) );
  ADDFX2 U142 ( .A(in_17bit_b[7]), .B(in_17bit_b[3]), .CI(
        add_1_root_r112_carry_7_), .CO(add_1_root_r112_carry_8_), .S(
        add_1_root_r112_SUM_7_) );
  ADDFX2 U143 ( .A(in_17bit_b[14]), .B(in_17bit_b[13]), .CI(
        add_3_root_r119_carry_15_), .CO(add_3_root_r119_carry_16_), .S(
        add_1_root_r119_A_15_) );
  ADDFX2 U144 ( .A(in_17bit_b[3]), .B(in_17bit_b[2]), .CI(
        add_3_root_r119_carry_4_), .CO(add_3_root_r119_carry_5_), .S(
        add_1_root_r119_A_4_) );
  ADDFX2 U145 ( .A(in_17bit_b[2]), .B(in_17bit_b[1]), .CI(
        add_3_root_r119_carry_3_), .CO(add_3_root_r119_carry_4_), .S(
        add_1_root_r119_A_3_) );
  ADDFX2 U146 ( .A(in_17bit_b[5]), .B(in_17bit_b[3]), .CI(
        add_1_root_r115_carry_9_), .CO(add_1_root_r115_carry_10_), .S(
        add_1_root_r115_SUM_9_) );
  ADDFX2 U147 ( .A(in_17bit_b[15]), .B(in_17bit_b[14]), .CI(
        add_3_root_r119_carry_16_), .CO(add_3_root_r119_carry_17_), .S(
        add_1_root_r119_A_16_) );
  ADDFX2 U148 ( .A(in_17bit_b[4]), .B(in_17bit_b[3]), .CI(
        add_3_root_r119_carry_5_), .CO(add_3_root_r119_carry_6_), .S(
        add_1_root_r119_A_5_) );
  ADDFX2 U149 ( .A(in_17bit_b[15]), .B(in_17bit_b[13]), .CI(
        add_2_root_r115_carry_16_), .CO(add_2_root_r115_carry_17_), .S(
        add_2_root_r115_SUM_16_) );
  ADDFX2 U150 ( .A(add_1_root_r119_A_18_), .B(in_17bit_b[12]), .CI(
        add_1_root_r119_carry[18]), .CO(add_1_root_r119_carry[19]), .S(
        add_1_root_r119_SUM_18_) );
  ADDFX2 U151 ( .A(in_17bit_b[15]), .B(in_17bit_b[13]), .CI(
        add_1_root_r115_carry_19_), .CO(add_1_root_r115_carry_20_), .S(
        add_1_root_r115_SUM_19_) );
  ADDFX2 U152 ( .A(in_17bit_b[4]), .B(in_17bit_b[3]), .CI(
        add_2_root_r119_carry_8_), .CO(add_2_root_r119_carry_9_), .S(
        add_2_root_r119_SUM_8_) );
  ADDFX2 U153 ( .A(in_17bit_b[5]), .B(in_17bit_b[4]), .CI(
        add_3_root_r119_carry_6_), .CO(add_3_root_r119_carry_7_), .S(
        add_1_root_r119_A_6_) );
  ADDFX2 U154 ( .A(in_17bit_b[14]), .B(in_17bit_b[13]), .CI(
        add_2_root_r119_carry_18_), .CO(add_2_root_r119_carry_19_), .S(
        add_2_root_r119_SUM_18_) );
  ADDFX2 U155 ( .A(in_17bit_b[15]), .B(in_17bit_b[14]), .CI(
        add_2_root_r119_carry_19_), .CO(add_2_root_r119_carry_20_), .S(
        add_2_root_r119_SUM_19_) );
  BUFX3 U156 ( .A(in_17bit_b[16]), .Y(n44) );
  INVX1 U157 ( .A(n261), .Y(in_17bit_b[16]) );
  INVX1 U158 ( .A(n203), .Y(n100) );
  NAND3BX1 U159 ( .AN(in_8bit[5]), .B(n46), .C(in_8bit[3]), .Y(n203) );
  INVX1 U160 ( .A(n54), .Y(n59) );
  INVX1 U161 ( .A(in_8bit[5]), .Y(n45) );
  INVX1 U162 ( .A(n54), .Y(n63) );
  INVX1 U163 ( .A(n54), .Y(n60) );
  XNOR2X1 U164 ( .A(n63), .B(n31), .Y(N29) );
  NAND2X1 U165 ( .A(sub_add_54_b0_carry[15]), .B(n179), .Y(n31) );
  CLKINVX3 U166 ( .A(n208), .Y(in_17bit_b[0]) );
  OAI21XL U167 ( .A0(n260), .A1(n261), .B0(n259), .Y(N463) );
  AOI22X1 U168 ( .A0(N221), .A1(n43), .B0(N363), .B1(n42), .Y(n259) );
  INVX1 U169 ( .A(n181), .Y(n260) );
  INVX1 U170 ( .A(n79), .Y(n84) );
  CLKINVX3 U171 ( .A(n253), .Y(in_17bit_b[15]) );
  INVX1 U172 ( .A(in_8bit[2]), .Y(n46) );
  AOI22X1 U173 ( .A0(N27), .A1(n57), .B0(in_17bit[14]), .B1(n60), .Y(n250) );
  AOI22X1 U174 ( .A0(N28), .A1(n57), .B0(in_17bit[15]), .B1(n59), .Y(n253) );
  AOI22X1 U175 ( .A0(N17), .A1(n57), .B0(in_17bit[4]), .B1(n63), .Y(n220) );
  AOI22X1 U176 ( .A0(N18), .A1(n57), .B0(in_17bit[5]), .B1(n60), .Y(n223) );
  AOI22X1 U177 ( .A0(N19), .A1(n57), .B0(in_17bit[6]), .B1(n59), .Y(n226) );
  AOI22X1 U178 ( .A0(N20), .A1(n57), .B0(in_17bit[7]), .B1(n63), .Y(n229) );
  AOI22X1 U179 ( .A0(N21), .A1(n57), .B0(in_17bit[8]), .B1(n60), .Y(n232) );
  AOI22X1 U180 ( .A0(N22), .A1(n57), .B0(in_17bit[9]), .B1(n60), .Y(n235) );
  AOI22X1 U181 ( .A0(N23), .A1(n57), .B0(in_17bit[10]), .B1(n63), .Y(n238) );
  AOI22X1 U182 ( .A0(N24), .A1(n57), .B0(in_17bit[11]), .B1(n59), .Y(n241) );
  AOI22X1 U183 ( .A0(N25), .A1(n57), .B0(in_17bit[12]), .B1(n59), .Y(n244) );
  AOI22X1 U184 ( .A0(N26), .A1(n57), .B0(in_17bit[13]), .B1(n63), .Y(n247) );
  AOI22X1 U185 ( .A0(N15), .A1(n57), .B0(in_17bit[2]), .B1(n59), .Y(n214) );
  NAND2X1 U186 ( .A(n70), .B(n8), .Y(n76) );
  AND2X2 U187 ( .A(n84), .B(n18), .Y(n33) );
  AND2X2 U188 ( .A(n33), .B(n4), .Y(n34) );
  AND2X2 U189 ( .A(n34), .B(n3), .Y(n35) );
  AND2X2 U190 ( .A(n35), .B(n5), .Y(n36) );
  BUFX3 U191 ( .A(n257), .Y(n42) );
  OAI2BB1X1 U192 ( .A0N(n100), .A1N(n29), .B0(n98), .Y(n257) );
  NAND2BX1 U193 ( .AN(n202), .B(n37), .Y(n98) );
  BUFX3 U194 ( .A(n258), .Y(n43) );
  OAI2BB1X1 U195 ( .A0N(n37), .A1N(n100), .B0(n99), .Y(n258) );
  NAND2BX1 U196 ( .AN(n202), .B(n29), .Y(n99) );
  NAND2BX1 U197 ( .AN(n76), .B(n7), .Y(n79) );
  INVX1 U198 ( .A(n66), .Y(n70) );
  OAI2BB1X1 U199 ( .A0N(n205), .A1N(n30), .B0(n158), .Y(n181) );
  NAND3BX1 U200 ( .AN(n101), .B(n206), .C(in_8bit[5]), .Y(n158) );
  AND2X2 U201 ( .A(n97), .B(n49), .Y(n37) );
  AND2X2 U202 ( .A(n36), .B(n13), .Y(n38) );
  INVX1 U203 ( .A(in_17bit[4]), .Y(n164) );
  INVX1 U204 ( .A(in_17bit[5]), .Y(n168) );
  INVX1 U205 ( .A(in_17bit[6]), .Y(n170) );
  INVX1 U206 ( .A(in_17bit[7]), .Y(n171) );
  INVX1 U207 ( .A(in_17bit[8]), .Y(n172) );
  INVX1 U208 ( .A(in_17bit[9]), .Y(n173) );
  INVX1 U209 ( .A(in_17bit[10]), .Y(n174) );
  INVX1 U210 ( .A(in_17bit[11]), .Y(n175) );
  INVX1 U211 ( .A(in_17bit[12]), .Y(n176) );
  INVX1 U212 ( .A(in_17bit[13]), .Y(n177) );
  INVX1 U213 ( .A(in_17bit[14]), .Y(n178) );
  INVX1 U214 ( .A(in_17bit[15]), .Y(n179) );
  INVX1 U215 ( .A(in_17bit[2]), .Y(n162) );
  INVX1 U216 ( .A(in_17bit[3]), .Y(n163) );
  INVX1 U217 ( .A(in_17bit[1]), .Y(n161) );
  INVX1 U218 ( .A(in_17bit[0]), .Y(n160) );
  NAND2X1 U219 ( .A(n210), .B(n209), .Y(N447) );
  AOI22X1 U220 ( .A0(N108), .A1(n254), .B0(N205), .B1(n43), .Y(n209) );
  AOI22X1 U221 ( .A0(N347), .A1(n42), .B0(n181), .B1(in_17bit_b[0]), .Y(n210)
         );
  NAND2X1 U222 ( .A(n213), .B(n212), .Y(N448) );
  AOI22X1 U223 ( .A0(N109), .A1(n254), .B0(N206), .B1(n43), .Y(n212) );
  AOI22X1 U224 ( .A0(N348), .A1(n42), .B0(n181), .B1(n180), .Y(n213) );
  INVX1 U225 ( .A(n211), .Y(n180) );
  NAND2X1 U226 ( .A(n216), .B(n215), .Y(N449) );
  AOI22X1 U227 ( .A0(N110), .A1(n254), .B0(N207), .B1(n43), .Y(n215) );
  AOI22X1 U228 ( .A0(N349), .A1(n42), .B0(n181), .B1(in_17bit_b[2]), .Y(n216)
         );
  NAND2X1 U229 ( .A(n219), .B(n218), .Y(N450) );
  AOI22X1 U230 ( .A0(N111), .A1(n254), .B0(N208), .B1(n43), .Y(n218) );
  AOI22X1 U231 ( .A0(N350), .A1(n42), .B0(n181), .B1(in_17bit_b[3]), .Y(n219)
         );
  NAND2X1 U232 ( .A(n222), .B(n221), .Y(N451) );
  AOI22X1 U233 ( .A0(N112), .A1(n254), .B0(N209), .B1(n43), .Y(n221) );
  AOI22X1 U234 ( .A0(N351), .A1(n42), .B0(n181), .B1(in_17bit_b[4]), .Y(n222)
         );
  NAND2X1 U235 ( .A(n225), .B(n224), .Y(N452) );
  AOI22X1 U236 ( .A0(N113), .A1(n254), .B0(N210), .B1(n43), .Y(n224) );
  AOI22X1 U237 ( .A0(N352), .A1(n42), .B0(n181), .B1(in_17bit_b[5]), .Y(n225)
         );
  NAND2X1 U238 ( .A(n228), .B(n227), .Y(N453) );
  AOI22X1 U239 ( .A0(N114), .A1(n254), .B0(N211), .B1(n43), .Y(n227) );
  AOI22X1 U240 ( .A0(N353), .A1(n42), .B0(n181), .B1(in_17bit_b[6]), .Y(n228)
         );
  NAND2X1 U241 ( .A(n231), .B(n230), .Y(N454) );
  AOI22X1 U242 ( .A0(N115), .A1(n254), .B0(N212), .B1(n43), .Y(n230) );
  AOI22X1 U243 ( .A0(N354), .A1(n42), .B0(n181), .B1(in_17bit_b[7]), .Y(n231)
         );
  NAND2X1 U244 ( .A(n234), .B(n233), .Y(N455) );
  AOI22X1 U245 ( .A0(N116), .A1(n254), .B0(N213), .B1(n43), .Y(n233) );
  AOI22X1 U246 ( .A0(N355), .A1(n42), .B0(n181), .B1(in_17bit_b[8]), .Y(n234)
         );
  NAND2X1 U247 ( .A(n237), .B(n236), .Y(N456) );
  AOI22X1 U248 ( .A0(N117), .A1(n254), .B0(N214), .B1(n43), .Y(n236) );
  AOI22X1 U249 ( .A0(N356), .A1(n42), .B0(n181), .B1(in_17bit_b[9]), .Y(n237)
         );
  NAND2X1 U250 ( .A(n240), .B(n239), .Y(N457) );
  AOI22X1 U251 ( .A0(N118), .A1(n254), .B0(N215), .B1(n43), .Y(n239) );
  AOI22X1 U252 ( .A0(N357), .A1(n42), .B0(n181), .B1(in_17bit_b[10]), .Y(n240)
         );
  NAND2X1 U253 ( .A(n243), .B(n242), .Y(N458) );
  AOI22X1 U254 ( .A0(N119), .A1(n254), .B0(N216), .B1(n43), .Y(n242) );
  AOI22X1 U255 ( .A0(N358), .A1(n42), .B0(n181), .B1(in_17bit_b[11]), .Y(n243)
         );
  NAND2X1 U256 ( .A(n246), .B(n245), .Y(N459) );
  AOI22X1 U257 ( .A0(N120), .A1(n254), .B0(N217), .B1(n43), .Y(n245) );
  AOI22X1 U258 ( .A0(N359), .A1(n42), .B0(n181), .B1(in_17bit_b[12]), .Y(n246)
         );
  NAND2X1 U259 ( .A(n249), .B(n248), .Y(N460) );
  AOI22X1 U260 ( .A0(N121), .A1(n254), .B0(N218), .B1(n43), .Y(n248) );
  AOI22X1 U261 ( .A0(N360), .A1(n42), .B0(n181), .B1(in_17bit_b[13]), .Y(n249)
         );
  NAND2X1 U262 ( .A(n252), .B(n251), .Y(N461) );
  AOI22X1 U263 ( .A0(N122), .A1(n254), .B0(N219), .B1(n43), .Y(n251) );
  AOI22X1 U264 ( .A0(N361), .A1(n42), .B0(n181), .B1(in_17bit_b[14]), .Y(n252)
         );
  NAND2X1 U265 ( .A(n256), .B(n255), .Y(N462) );
  AOI22X1 U266 ( .A0(N123), .A1(n254), .B0(N220), .B1(n43), .Y(n255) );
  AOI22X1 U267 ( .A0(N362), .A1(n42), .B0(n181), .B1(in_17bit_b[15]), .Y(n256)
         );
  MX2X1 U268 ( .A(neg_mul[21]), .B(N479), .S0(n92), .Y(out[14]) );
  INVX1 U269 ( .A(n65), .Y(n64) );
  XNOR2X1 U270 ( .A(n14), .B(sub_add_75_b0_carry[10]), .Y(n39) );
  XNOR2X1 U271 ( .A(n15), .B(sub_add_75_b0_carry[11]), .Y(n40) );
  INVX1 U272 ( .A(n72), .Y(n71) );
  INVX1 U273 ( .A(n78), .Y(n77) );
  MX2X1 U274 ( .A(neg_mul[22]), .B(N480), .S0(n92), .Y(out[15]) );
  MX2X1 U275 ( .A(neg_mul[23]), .B(N481), .S0(n92), .Y(out[16]) );
  NAND4BBX1 U276 ( .AN(n42), .BN(n43), .C(n207), .D(n260), .Y(N446) );
  NOR4BX1 U277 ( .AN(n204), .B(n49), .C(n50), .D(in_8bit[2]), .Y(n205) );
  NOR2X1 U278 ( .A(in_8bit[6]), .B(in_8bit[3]), .Y(n204) );
  NAND4BXL U279 ( .AN(n52), .B(n50), .C(in_8bit[4]), .D(in_8bit[6]), .Y(n101)
         );
  NAND2X1 U280 ( .A(n96), .B(n95), .Y(n254) );
  NAND3BX1 U281 ( .AN(n93), .B(n206), .C(in_8bit[6]), .Y(n96) );
  NAND3X1 U282 ( .A(n205), .B(in_8bit[5]), .C(n94), .Y(n95) );
  NOR2X1 U283 ( .A(in_8bit[6]), .B(in_8bit[4]), .Y(n201) );
  NAND2BX1 U284 ( .AN(n70), .B(neg_mul[9]), .Y(n72) );
  NAND2X1 U285 ( .A(neg_mul[10]), .B(n76), .Y(n78) );
  NAND2X1 U286 ( .A(out[0]), .B(neg_mul[8]), .Y(n65) );
  OR2X2 U287 ( .A(out[0]), .B(neg_mul[8]), .Y(n66) );
  NAND2XL U288 ( .A(N29), .B(n54), .Y(n261) );
  AOI22XL U289 ( .A0(N16), .A1(n54), .B0(in_17bit[3]), .B1(n59), .Y(n217) );
  AOI22XL U290 ( .A0(in_17bit[0]), .A1(n54), .B0(in_17bit[0]), .B1(n60), .Y(
        n208) );
  AOI22XL U291 ( .A0(N14), .A1(n54), .B0(in_17bit[1]), .B1(n60), .Y(n211) );
  AOI2BB1X4 U292 ( .A0N(n55), .A1N(n69), .B0(n68), .Y(out[1]) );
  OAI21X4 U293 ( .A0(n73), .A1(n61), .B0(n76), .Y(n74) );
  AOI2BB1X4 U294 ( .A0N(n55), .A1N(n75), .B0(n74), .Y(out[2]) );
  AOI2BB1X4 U295 ( .A0N(n55), .A1N(n82), .B0(n81), .Y(out[3]) );
  NOR2X4 U296 ( .A(n33), .B(n86), .Y(n87) );
  XNOR2X4 U297 ( .A(n87), .B(n4), .Y(out[5]) );
  XNOR2X4 U298 ( .A(n91), .B(n5), .Y(out[7]) );
  AND2X1 U299 ( .A(add_1_root_r112_carry_20_), .B(n44), .Y(
        add_1_root_r112_SUM_21_) );
  XOR2X1 U300 ( .A(n44), .B(add_1_root_r112_carry_20_), .Y(
        add_1_root_r112_SUM_20_) );
  AND2X1 U301 ( .A(add_1_root_r112_carry_19_), .B(in_17bit_b[15]), .Y(
        add_1_root_r112_carry_20_) );
  XOR2X1 U302 ( .A(in_17bit_b[15]), .B(add_1_root_r112_carry_19_), .Y(
        add_1_root_r112_SUM_19_) );
  AND2X1 U303 ( .A(add_1_root_r112_carry_18_), .B(in_17bit_b[14]), .Y(
        add_1_root_r112_carry_19_) );
  XOR2X1 U304 ( .A(in_17bit_b[14]), .B(add_1_root_r112_carry_18_), .Y(
        add_1_root_r112_SUM_18_) );
  AND2X1 U305 ( .A(add_1_root_r112_carry_17_), .B(in_17bit_b[13]), .Y(
        add_1_root_r112_carry_18_) );
  XOR2X1 U306 ( .A(in_17bit_b[13]), .B(add_1_root_r112_carry_17_), .Y(
        add_1_root_r112_SUM_17_) );
  AND2X1 U307 ( .A(add_2_root_r119_carry_21_), .B(n44), .Y(
        add_2_root_r119_SUM_22_) );
  XOR2X1 U308 ( .A(n44), .B(add_2_root_r119_carry_21_), .Y(
        add_2_root_r119_SUM_21_) );
  AND2X1 U309 ( .A(in_17bit_b[1]), .B(in_17bit_b[0]), .Y(
        add_2_root_r119_carry_6_) );
  XOR2X1 U310 ( .A(in_17bit_b[0]), .B(in_17bit_b[1]), .Y(
        add_2_root_r119_SUM_5_) );
  AND2X1 U311 ( .A(add_1_root_r119_carry[22]), .B(n44), .Y(
        add_1_root_r119_SUM_23_) );
  XOR2X1 U312 ( .A(n44), .B(add_1_root_r119_carry[22]), .Y(
        add_1_root_r119_SUM_22_) );
  AND2X1 U313 ( .A(add_1_root_r119_carry[21]), .B(in_17bit_b[15]), .Y(
        add_1_root_r119_carry[22]) );
  XOR2X1 U314 ( .A(in_17bit_b[15]), .B(add_1_root_r119_carry[21]), .Y(
        add_1_root_r119_SUM_21_) );
  AND2X1 U315 ( .A(add_1_root_r119_carry[20]), .B(in_17bit_b[14]), .Y(
        add_1_root_r119_carry[21]) );
  XOR2X1 U316 ( .A(in_17bit_b[14]), .B(add_1_root_r119_carry[20]), .Y(
        add_1_root_r119_SUM_20_) );
  AND2X1 U317 ( .A(add_1_root_r119_A_6_), .B(in_17bit_b[0]), .Y(
        add_1_root_r119_carry[7]) );
  XOR2X1 U318 ( .A(in_17bit_b[0]), .B(add_1_root_r119_A_6_), .Y(
        add_1_root_r119_SUM_6_) );
  AND2X1 U319 ( .A(add_3_root_r119_carry_18_), .B(n44), .Y(
        add_1_root_r119_A_19_) );
  XOR2X1 U320 ( .A(n44), .B(add_3_root_r119_carry_18_), .Y(
        add_1_root_r119_A_18_) );
  AND2X1 U321 ( .A(in_17bit_b[1]), .B(in_17bit_b[0]), .Y(
        add_3_root_r119_carry_3_) );
  XOR2X1 U322 ( .A(in_17bit_b[0]), .B(in_17bit_b[1]), .Y(add_1_root_r119_A_2_)
         );
  AND2X1 U323 ( .A(add_2_root_r115_carry_19_), .B(n44), .Y(
        add_2_root_r115_SUM_20_) );
  XOR2X1 U324 ( .A(n44), .B(add_2_root_r115_carry_19_), .Y(
        add_2_root_r115_SUM_19_) );
  AND2X1 U325 ( .A(add_2_root_r115_carry_18_), .B(in_17bit_b[15]), .Y(
        add_2_root_r115_carry_19_) );
  XOR2X1 U326 ( .A(in_17bit_b[15]), .B(add_2_root_r115_carry_18_), .Y(
        add_2_root_r115_SUM_18_) );
  AND2X1 U327 ( .A(in_17bit_b[2]), .B(in_17bit_b[0]), .Y(
        add_2_root_r115_carry_4_) );
  XOR2X1 U328 ( .A(in_17bit_b[0]), .B(in_17bit_b[2]), .Y(
        add_2_root_r115_SUM_3_) );
  AND2X1 U329 ( .A(add_1_root_r115_carry_22_), .B(n44), .Y(
        add_1_root_r115_SUM_23_) );
  XOR2X1 U330 ( .A(n44), .B(add_1_root_r115_carry_22_), .Y(
        add_1_root_r115_SUM_22_) );
  AND2X1 U331 ( .A(add_1_root_r115_carry_21_), .B(in_17bit_b[15]), .Y(
        add_1_root_r115_carry_22_) );
  XOR2X1 U332 ( .A(in_17bit_b[15]), .B(add_1_root_r115_carry_21_), .Y(
        add_1_root_r115_SUM_21_) );
  AND2X1 U333 ( .A(in_17bit_b[2]), .B(in_17bit_b[0]), .Y(
        add_1_root_r115_carry_7_) );
  XOR2X1 U334 ( .A(in_17bit_b[0]), .B(in_17bit_b[2]), .Y(
        add_1_root_r115_SUM_6_) );
  XOR2X1 U335 ( .A(n179), .B(sub_add_54_b0_carry[15]), .Y(N28) );
  AND2X1 U336 ( .A(sub_add_54_b0_carry[14]), .B(n178), .Y(
        sub_add_54_b0_carry[15]) );
  XOR2X1 U337 ( .A(n178), .B(sub_add_54_b0_carry[14]), .Y(N27) );
  AND2X1 U338 ( .A(sub_add_54_b0_carry[13]), .B(n177), .Y(
        sub_add_54_b0_carry[14]) );
  XOR2X1 U339 ( .A(n177), .B(sub_add_54_b0_carry[13]), .Y(N26) );
  AND2X1 U340 ( .A(sub_add_54_b0_carry[12]), .B(n176), .Y(
        sub_add_54_b0_carry[13]) );
  XOR2X1 U341 ( .A(n176), .B(sub_add_54_b0_carry[12]), .Y(N25) );
  AND2X1 U342 ( .A(sub_add_54_b0_carry[11]), .B(n175), .Y(
        sub_add_54_b0_carry[12]) );
  XOR2X1 U343 ( .A(n175), .B(sub_add_54_b0_carry[11]), .Y(N24) );
  AND2X1 U344 ( .A(sub_add_54_b0_carry[10]), .B(n174), .Y(
        sub_add_54_b0_carry[11]) );
  XOR2X1 U345 ( .A(n174), .B(sub_add_54_b0_carry[10]), .Y(N23) );
  AND2X1 U346 ( .A(sub_add_54_b0_carry[9]), .B(n173), .Y(
        sub_add_54_b0_carry[10]) );
  XOR2X1 U347 ( .A(n173), .B(sub_add_54_b0_carry[9]), .Y(N22) );
  AND2X1 U348 ( .A(sub_add_54_b0_carry[8]), .B(n172), .Y(
        sub_add_54_b0_carry[9]) );
  XOR2X1 U349 ( .A(n172), .B(sub_add_54_b0_carry[8]), .Y(N21) );
  AND2X1 U350 ( .A(sub_add_54_b0_carry[7]), .B(n171), .Y(
        sub_add_54_b0_carry[8]) );
  XOR2X1 U351 ( .A(n171), .B(sub_add_54_b0_carry[7]), .Y(N20) );
  AND2X1 U352 ( .A(sub_add_54_b0_carry[6]), .B(n170), .Y(
        sub_add_54_b0_carry[7]) );
  XOR2X1 U353 ( .A(n170), .B(sub_add_54_b0_carry[6]), .Y(N19) );
  AND2X1 U354 ( .A(sub_add_54_b0_carry[5]), .B(n168), .Y(
        sub_add_54_b0_carry[6]) );
  XOR2X1 U355 ( .A(n168), .B(sub_add_54_b0_carry[5]), .Y(N18) );
  AND2X1 U356 ( .A(sub_add_54_b0_carry[4]), .B(n164), .Y(
        sub_add_54_b0_carry[5]) );
  XOR2X1 U357 ( .A(n164), .B(sub_add_54_b0_carry[4]), .Y(N17) );
  AND2X1 U358 ( .A(sub_add_54_b0_carry[3]), .B(n163), .Y(
        sub_add_54_b0_carry[4]) );
  XOR2X1 U359 ( .A(n163), .B(sub_add_54_b0_carry[3]), .Y(N16) );
  AND2X1 U360 ( .A(sub_add_54_b0_carry[2]), .B(n162), .Y(
        sub_add_54_b0_carry[3]) );
  XOR2X1 U361 ( .A(n162), .B(sub_add_54_b0_carry[2]), .Y(N15) );
  AND2X1 U362 ( .A(n160), .B(n161), .Y(sub_add_54_b0_carry[2]) );
  XOR2X1 U363 ( .A(n161), .B(n160), .Y(N14) );
  XOR2X1 U364 ( .A(n17), .B(sub_add_75_b0_carry[16]), .Y(N481) );
  AND2X1 U365 ( .A(sub_add_75_b0_carry[15]), .B(n11), .Y(
        sub_add_75_b0_carry[16]) );
  XOR2X1 U366 ( .A(n11), .B(sub_add_75_b0_carry[15]), .Y(N480) );
  AND2X1 U367 ( .A(sub_add_75_b0_carry[14]), .B(n12), .Y(
        sub_add_75_b0_carry[15]) );
  XOR2X1 U368 ( .A(n12), .B(sub_add_75_b0_carry[14]), .Y(N479) );
  AND2X1 U369 ( .A(sub_add_75_b0_carry[13]), .B(n9), .Y(
        sub_add_75_b0_carry[14]) );
  XOR2X1 U370 ( .A(n9), .B(sub_add_75_b0_carry[13]), .Y(N478) );
  AND2X1 U371 ( .A(sub_add_75_b0_carry[12]), .B(n10), .Y(
        sub_add_75_b0_carry[13]) );
  AND2X1 U372 ( .A(sub_add_75_b0_carry[11]), .B(n15), .Y(
        sub_add_75_b0_carry[12]) );
  AND2X1 U373 ( .A(sub_add_75_b0_carry[10]), .B(n14), .Y(
        sub_add_75_b0_carry[11]) );
  AND2X1 U374 ( .A(n38), .B(n6), .Y(sub_add_75_b0_carry[10]) );
  AND2X1 U375 ( .A(in_17bit_b[0]), .B(in_17bit_b[4]), .Y(
        add_1_root_r112_carry_5_) );
endmodule


module multi16_1_DW01_add_0 ( A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, 
        A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, 
        A_4_, B_23_, B_22_, B_21_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, 
        B_14_, B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, 
        SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, 
        SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, 
        SUM_7_ );
  input A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_,
         A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, B_23_, B_22_,
         B_21_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_,
         B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_;
  output SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_,
         SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_,
         SUM_8_, SUM_7_;
  wire   n1, n2, n3, n4;
  wire   [23:7] carry;

  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry[7]), .CO(carry[8]), .S(SUM_7_)
         );
  ADDFX2 U1_21 ( .A(A_21_), .B(B_21_), .CI(carry[21]), .CO(carry[22]), .S(
        SUM_21_) );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry[20]), .CO(carry[21]), .S(
        SUM_20_) );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry[19]), .CO(carry[20]), .S(
        SUM_19_) );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry[18]), .CO(carry[19]), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry[17]), .CO(carry[18]), .S(
        SUM_17_) );
  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry[16]), .CO(carry[17]), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry[15]), .CO(carry[16]), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry[14]), .CO(carry[15]), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry[13]), .CO(carry[14]), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry[12]), .CO(carry[13]), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry[11]), .CO(carry[12]), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry[10]), .CO(carry[11]), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry[9]), .CO(carry[10]), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry[8]), .CO(carry[9]), .S(SUM_8_)
         );
  ADDFX2 U1_22 ( .A(A_22_), .B(B_22_), .CI(carry[22]), .CO(carry[23]), .S(
        SUM_22_) );
  AND2X2 U1 ( .A(A_4_), .B(B_4_), .Y(n1) );
  XOR2X1 U2 ( .A(B_23_), .B(carry[23]), .Y(SUM_23_) );
  OAI2BB1X1 U3 ( .A0N(n2), .A1N(A_6_), .B0(n3), .Y(carry[7]) );
  OAI21XL U4 ( .A0(A_6_), .A1(n2), .B0(B_6_), .Y(n3) );
  OAI2BB1X1 U5 ( .A0N(n1), .A1N(A_5_), .B0(n4), .Y(n2) );
  OAI21XL U6 ( .A0(A_5_), .A1(n1), .B0(B_5_), .Y(n4) );
endmodule


module multi16_1_DW01_add_4 ( A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, 
        A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, 
        B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, 
        B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, SUM_22_, SUM_21_, SUM_20_, 
        SUM_19_, SUM_18_, SUM_17_, SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, 
        SUM_11_, SUM_10_, SUM_9_, SUM_8_, SUM_7_ );
  input A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_,
         A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, B_20_, B_19_,
         B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, B_10_, B_9_,
         B_8_, B_7_, B_6_, B_5_;
  output SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_,
         SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_,
         SUM_7_;
  wire   carry_21_, carry_20_, carry_19_, carry_18_, carry_17_, carry_16_,
         carry_15_, carry_14_, carry_13_, carry_12_, carry_11_, carry_10_,
         carry_9_, carry_8_, carry_7_, n1;

  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry_16_), .CO(carry_17_), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry_15_), .CO(carry_16_), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry_14_), .CO(carry_15_), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry_13_), .CO(carry_14_), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry_12_), .CO(carry_13_), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry_11_), .CO(carry_12_), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry_10_), .CO(carry_11_), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry_9_), .CO(carry_10_), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry_8_), .CO(carry_9_), .S(SUM_8_)
         );
  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry_7_), .CO(carry_8_), .S(SUM_7_)
         );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry_20_), .CO(carry_21_), .S(
        SUM_20_) );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry_19_), .CO(carry_20_), .S(
        SUM_19_) );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry_18_), .CO(carry_19_), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry_17_), .CO(carry_18_), .S(
        SUM_17_) );
  ADDFX2 U1_21 ( .A(A_21_), .B(B_21_), .CI(carry_21_), .CO(SUM_22_), .S(
        SUM_21_) );
  OAI2BB1X1 U1 ( .A0N(A_6_), .A1N(B_6_), .B0(n1), .Y(carry_7_) );
  OAI211X1 U2 ( .A0(B_6_), .A1(A_6_), .B0(A_5_), .C0(B_5_), .Y(n1) );
endmodule


module multi16_1_DW01_add_6 ( A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, 
        A_16_, A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, 
        A_6_, A_5_, A_4_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, 
        B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, 
        SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, 
        SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, 
        SUM_7_ );
  input A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_,
         A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, B_20_,
         B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, B_10_,
         B_9_, B_8_, B_7_, B_6_, B_5_, B_4_;
  output SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_,
         SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_,
         SUM_8_, SUM_7_;
  wire   n1, n2, n3, n4, n5, n6;
  wire   [21:7] carry;

  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry[7]), .CO(carry[8]), .S(SUM_7_)
         );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry[18]), .CO(carry[19]), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry[17]), .CO(carry[18]), .S(
        SUM_17_) );
  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry[16]), .CO(carry[17]), .S(
        SUM_16_) );
  ADDFX2 U1_15 ( .A(A_15_), .B(B_15_), .CI(carry[15]), .CO(carry[16]), .S(
        SUM_15_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry[14]), .CO(carry[15]), .S(
        SUM_14_) );
  ADDFX2 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry[13]), .CO(carry[14]), .S(
        SUM_13_) );
  ADDFX2 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry[12]), .CO(carry[13]), .S(
        SUM_12_) );
  ADDFX2 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry[11]), .CO(carry[12]), .S(
        SUM_11_) );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry[10]), .CO(carry[11]), .S(
        SUM_10_) );
  ADDFX2 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry[9]), .CO(carry[10]), .S(SUM_9_)
         );
  ADDFX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry[8]), .CO(carry[9]), .S(SUM_8_)
         );
  ADDFX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry[19]), .CO(carry[20]), .S(
        SUM_19_) );
  ADDFX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry[20]), .CO(carry[21]), .S(
        SUM_20_) );
  AND2X2 U1 ( .A(A_22_), .B(n2), .Y(n1) );
  AND2X2 U2 ( .A(A_21_), .B(carry[21]), .Y(n2) );
  XOR2X1 U3 ( .A(A_23_), .B(n1), .Y(SUM_23_) );
  XOR2X1 U4 ( .A(A_21_), .B(carry[21]), .Y(SUM_21_) );
  XOR2X1 U5 ( .A(A_22_), .B(n2), .Y(SUM_22_) );
  AND2X2 U6 ( .A(A_4_), .B(B_4_), .Y(n3) );
  OAI2BB1X1 U7 ( .A0N(n4), .A1N(A_6_), .B0(n5), .Y(carry[7]) );
  OAI21XL U8 ( .A0(A_6_), .A1(n4), .B0(B_6_), .Y(n5) );
  OAI2BB1X1 U9 ( .A0N(n3), .A1N(A_5_), .B0(n6), .Y(n4) );
  OAI21XL U10 ( .A0(A_5_), .A1(n3), .B0(B_5_), .Y(n6) );
endmodule


module multi16_1 ( in_17bit, in_8bit, out );
  input [16:0] in_17bit;
  input [7:0] in_8bit;
  output [16:0] out;
  wire   n262, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26,
         N27, N28, N29, N108, N109, N110, N111, N112, N113, N114, N115, N116,
         N117, N118, N119, N120, N121, N122, N123, N205, N206, N207, N208,
         N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, N219,
         N220, N221, N347, N348, N349, N350, N351, N352, N353, N354, N355,
         N356, N357, N358, N359, N360, N361, N362, N363, N446, N447, N448,
         N449, N450, N451, N452, N453, N454, N455, N456, N457, N458, N459,
         N460, N461, N462, N463, N477, N478, N479, N480,
         add_2_root_r119_carry_10_, add_2_root_r119_carry_11_,
         add_2_root_r119_carry_12_, add_2_root_r119_carry_13_,
         add_2_root_r119_carry_14_, add_2_root_r119_carry_15_,
         add_2_root_r119_carry_16_, add_2_root_r119_carry_17_,
         add_2_root_r119_carry_18_, add_2_root_r119_carry_19_,
         add_2_root_r119_carry_20_, add_2_root_r119_carry_21_,
         add_2_root_r119_carry_6_, add_2_root_r119_carry_7_,
         add_2_root_r119_carry_8_, add_2_root_r119_carry_9_,
         add_2_root_r119_SUM_5_, add_2_root_r119_SUM_6_,
         add_2_root_r119_SUM_7_, add_2_root_r119_SUM_8_,
         add_2_root_r119_SUM_9_, add_2_root_r119_SUM_10_,
         add_2_root_r119_SUM_11_, add_2_root_r119_SUM_12_,
         add_2_root_r119_SUM_13_, add_2_root_r119_SUM_14_,
         add_2_root_r119_SUM_15_, add_2_root_r119_SUM_16_,
         add_2_root_r119_SUM_17_, add_2_root_r119_SUM_18_,
         add_2_root_r119_SUM_19_, add_2_root_r119_SUM_20_,
         add_2_root_r119_SUM_21_, add_2_root_r119_SUM_22_,
         add_1_root_r119_SUM_6_, add_1_root_r119_SUM_7_,
         add_1_root_r119_SUM_8_, add_1_root_r119_SUM_9_,
         add_1_root_r119_SUM_10_, add_1_root_r119_SUM_11_,
         add_1_root_r119_SUM_12_, add_1_root_r119_SUM_13_,
         add_1_root_r119_SUM_14_, add_1_root_r119_SUM_15_,
         add_1_root_r119_SUM_16_, add_1_root_r119_SUM_17_,
         add_1_root_r119_SUM_18_, add_1_root_r119_SUM_19_,
         add_1_root_r119_SUM_20_, add_1_root_r119_SUM_21_,
         add_1_root_r119_SUM_22_, add_1_root_r119_SUM_23_,
         add_1_root_r119_A_2_, add_1_root_r119_A_3_, add_1_root_r119_A_4_,
         add_1_root_r119_A_5_, add_1_root_r119_A_6_, add_1_root_r119_A_7_,
         add_1_root_r119_A_8_, add_1_root_r119_A_9_, add_1_root_r119_A_10_,
         add_1_root_r119_A_11_, add_1_root_r119_A_12_, add_1_root_r119_A_13_,
         add_1_root_r119_A_14_, add_1_root_r119_A_15_, add_1_root_r119_A_16_,
         add_1_root_r119_A_17_, add_1_root_r119_A_18_, add_1_root_r119_A_19_,
         add_3_root_r119_carry_10_, add_3_root_r119_carry_11_,
         add_3_root_r119_carry_12_, add_3_root_r119_carry_13_,
         add_3_root_r119_carry_14_, add_3_root_r119_carry_15_,
         add_3_root_r119_carry_16_, add_3_root_r119_carry_17_,
         add_3_root_r119_carry_18_, add_3_root_r119_carry_3_,
         add_3_root_r119_carry_4_, add_3_root_r119_carry_5_,
         add_3_root_r119_carry_6_, add_3_root_r119_carry_7_,
         add_3_root_r119_carry_8_, add_3_root_r119_carry_9_,
         add_1_root_r112_carry_10_, add_1_root_r112_carry_11_,
         add_1_root_r112_carry_12_, add_1_root_r112_carry_13_,
         add_1_root_r112_carry_14_, add_1_root_r112_carry_15_,
         add_1_root_r112_carry_16_, add_1_root_r112_carry_17_,
         add_1_root_r112_carry_18_, add_1_root_r112_carry_19_,
         add_1_root_r112_carry_20_, add_1_root_r112_carry_5_,
         add_1_root_r112_carry_6_, add_1_root_r112_carry_7_,
         add_1_root_r112_carry_8_, add_1_root_r112_carry_9_,
         add_1_root_r112_SUM_1_, add_1_root_r112_SUM_2_,
         add_1_root_r112_SUM_3_, add_1_root_r112_SUM_4_,
         add_1_root_r112_SUM_5_, add_1_root_r112_SUM_6_,
         add_1_root_r112_SUM_7_, add_1_root_r112_SUM_8_,
         add_1_root_r112_SUM_9_, add_1_root_r112_SUM_10_,
         add_1_root_r112_SUM_11_, add_1_root_r112_SUM_12_,
         add_1_root_r112_SUM_13_, add_1_root_r112_SUM_14_,
         add_1_root_r112_SUM_15_, add_1_root_r112_SUM_16_,
         add_1_root_r112_SUM_17_, add_1_root_r112_SUM_18_,
         add_1_root_r112_SUM_19_, add_1_root_r112_SUM_20_,
         add_1_root_r112_SUM_21_, add_2_root_r115_carry_10_,
         add_2_root_r115_carry_11_, add_2_root_r115_carry_12_,
         add_2_root_r115_carry_13_, add_2_root_r115_carry_14_,
         add_2_root_r115_carry_15_, add_2_root_r115_carry_16_,
         add_2_root_r115_carry_17_, add_2_root_r115_carry_18_,
         add_2_root_r115_carry_19_, add_2_root_r115_carry_4_,
         add_2_root_r115_carry_5_, add_2_root_r115_carry_6_,
         add_2_root_r115_carry_7_, add_2_root_r115_carry_8_,
         add_2_root_r115_carry_9_, add_2_root_r115_SUM_3_,
         add_2_root_r115_SUM_4_, add_2_root_r115_SUM_5_,
         add_2_root_r115_SUM_6_, add_2_root_r115_SUM_7_,
         add_2_root_r115_SUM_8_, add_2_root_r115_SUM_9_,
         add_2_root_r115_SUM_10_, add_2_root_r115_SUM_11_,
         add_2_root_r115_SUM_12_, add_2_root_r115_SUM_13_,
         add_2_root_r115_SUM_14_, add_2_root_r115_SUM_15_,
         add_2_root_r115_SUM_16_, add_2_root_r115_SUM_17_,
         add_2_root_r115_SUM_18_, add_2_root_r115_SUM_19_,
         add_2_root_r115_SUM_20_, add_1_root_r115_carry_10_,
         add_1_root_r115_carry_11_, add_1_root_r115_carry_12_,
         add_1_root_r115_carry_13_, add_1_root_r115_carry_14_,
         add_1_root_r115_carry_15_, add_1_root_r115_carry_16_,
         add_1_root_r115_carry_17_, add_1_root_r115_carry_18_,
         add_1_root_r115_carry_19_, add_1_root_r115_carry_20_,
         add_1_root_r115_carry_21_, add_1_root_r115_carry_22_,
         add_1_root_r115_carry_7_, add_1_root_r115_carry_8_,
         add_1_root_r115_carry_9_, add_1_root_r115_SUM_6_,
         add_1_root_r115_SUM_7_, add_1_root_r115_SUM_8_,
         add_1_root_r115_SUM_9_, add_1_root_r115_SUM_10_,
         add_1_root_r115_SUM_11_, add_1_root_r115_SUM_12_,
         add_1_root_r115_SUM_13_, add_1_root_r115_SUM_14_,
         add_1_root_r115_SUM_15_, add_1_root_r115_SUM_16_,
         add_1_root_r115_SUM_17_, add_1_root_r115_SUM_18_,
         add_1_root_r115_SUM_19_, add_1_root_r115_SUM_20_,
         add_1_root_r115_SUM_21_, add_1_root_r115_SUM_22_,
         add_1_root_r115_SUM_23_, n1, n2, n3, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n158, n160, n163, n164, n167, n168, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261;
  wire   [16:0] in_17bit_b;
  wire   [23:8] neg_mul;
  wire   [15:10] sub_add_75_b0_carry;
  wire   [16:2] sub_add_54_b0_carry;
  wire   [22:7] add_1_root_r119_carry;

  multi16_1_DW01_add_0 add_0_root_r119 ( .A_22_(add_2_root_r119_SUM_22_), 
        .A_21_(add_2_root_r119_SUM_21_), .A_20_(add_2_root_r119_SUM_20_), 
        .A_19_(add_2_root_r119_SUM_19_), .A_18_(add_2_root_r119_SUM_18_), 
        .A_17_(add_2_root_r119_SUM_17_), .A_16_(add_2_root_r119_SUM_16_), 
        .A_15_(add_2_root_r119_SUM_15_), .A_14_(add_2_root_r119_SUM_14_), 
        .A_13_(add_2_root_r119_SUM_13_), .A_12_(add_2_root_r119_SUM_12_), 
        .A_11_(add_2_root_r119_SUM_11_), .A_10_(add_2_root_r119_SUM_10_), 
        .A_9_(add_2_root_r119_SUM_9_), .A_8_(add_2_root_r119_SUM_8_), .A_7_(
        add_2_root_r119_SUM_7_), .A_6_(add_2_root_r119_SUM_6_), .A_5_(
        add_2_root_r119_SUM_5_), .A_4_(in_17bit_b[0]), .B_23_(
        add_1_root_r119_SUM_23_), .B_22_(add_1_root_r119_SUM_22_), .B_21_(
        add_1_root_r119_SUM_21_), .B_20_(add_1_root_r119_SUM_20_), .B_19_(
        add_1_root_r119_SUM_19_), .B_18_(add_1_root_r119_SUM_18_), .B_17_(
        add_1_root_r119_SUM_17_), .B_16_(add_1_root_r119_SUM_16_), .B_15_(
        add_1_root_r119_SUM_15_), .B_14_(add_1_root_r119_SUM_14_), .B_13_(
        add_1_root_r119_SUM_13_), .B_12_(add_1_root_r119_SUM_12_), .B_11_(
        add_1_root_r119_SUM_11_), .B_10_(add_1_root_r119_SUM_10_), .B_9_(
        add_1_root_r119_SUM_9_), .B_8_(add_1_root_r119_SUM_8_), .B_7_(
        add_1_root_r119_SUM_7_), .B_6_(add_1_root_r119_SUM_6_), .B_5_(
        add_1_root_r119_A_5_), .B_4_(add_1_root_r119_A_4_), .SUM_23_(N363), 
        .SUM_22_(N362), .SUM_21_(N361), .SUM_20_(N360), .SUM_19_(N359), 
        .SUM_18_(N358), .SUM_17_(N357), .SUM_16_(N356), .SUM_15_(N355), 
        .SUM_14_(N354), .SUM_13_(N353), .SUM_12_(N352), .SUM_11_(N351), 
        .SUM_10_(N350), .SUM_9_(N349), .SUM_8_(N348), .SUM_7_(N347) );
  multi16_1_DW01_add_4 add_0_root_r112 ( .A_21_(n41), .A_20_(in_17bit_b[15]), 
        .A_19_(in_17bit_b[14]), .A_18_(in_17bit_b[13]), .A_17_(in_17bit_b[12]), 
        .A_16_(in_17bit_b[11]), .A_15_(in_17bit_b[10]), .A_14_(in_17bit_b[9]), 
        .A_13_(in_17bit_b[8]), .A_12_(in_17bit_b[7]), .A_11_(in_17bit_b[6]), 
        .A_10_(in_17bit_b[5]), .A_9_(in_17bit_b[4]), .A_8_(in_17bit_b[3]), 
        .A_7_(in_17bit_b[2]), .A_6_(in_17bit_b[1]), .A_5_(in_17bit_b[0]), 
        .B_21_(add_1_root_r112_SUM_21_), .B_20_(add_1_root_r112_SUM_20_), 
        .B_19_(add_1_root_r112_SUM_19_), .B_18_(add_1_root_r112_SUM_18_), 
        .B_17_(add_1_root_r112_SUM_17_), .B_16_(add_1_root_r112_SUM_16_), 
        .B_15_(add_1_root_r112_SUM_15_), .B_14_(add_1_root_r112_SUM_14_), 
        .B_13_(add_1_root_r112_SUM_13_), .B_12_(add_1_root_r112_SUM_12_), 
        .B_11_(add_1_root_r112_SUM_11_), .B_10_(add_1_root_r112_SUM_10_), 
        .B_9_(add_1_root_r112_SUM_9_), .B_8_(add_1_root_r112_SUM_8_), .B_7_(
        add_1_root_r112_SUM_7_), .B_6_(add_1_root_r112_SUM_6_), .B_5_(
        add_1_root_r112_SUM_5_), .SUM_22_(N123), .SUM_21_(N122), .SUM_20_(N121), .SUM_19_(N120), .SUM_18_(N119), .SUM_17_(N118), .SUM_16_(N117), .SUM_15_(
        N116), .SUM_14_(N115), .SUM_13_(N114), .SUM_12_(N113), .SUM_11_(N112), 
        .SUM_10_(N111), .SUM_9_(N110), .SUM_8_(N109), .SUM_7_(N108) );
  multi16_1_DW01_add_6 add_0_root_r115 ( .A_23_(add_1_root_r115_SUM_23_), 
        .A_22_(add_1_root_r115_SUM_22_), .A_21_(add_1_root_r115_SUM_21_), 
        .A_20_(add_1_root_r115_SUM_20_), .A_19_(add_1_root_r115_SUM_19_), 
        .A_18_(add_1_root_r115_SUM_18_), .A_17_(add_1_root_r115_SUM_17_), 
        .A_16_(add_1_root_r115_SUM_16_), .A_15_(add_1_root_r115_SUM_15_), 
        .A_14_(add_1_root_r115_SUM_14_), .A_13_(add_1_root_r115_SUM_13_), 
        .A_12_(add_1_root_r115_SUM_12_), .A_11_(add_1_root_r115_SUM_11_), 
        .A_10_(add_1_root_r115_SUM_10_), .A_9_(add_1_root_r115_SUM_9_), .A_8_(
        add_1_root_r115_SUM_8_), .A_7_(add_1_root_r115_SUM_7_), .A_6_(
        add_1_root_r115_SUM_6_), .A_5_(in_17bit_b[1]), .A_4_(in_17bit_b[0]), 
        .B_20_(add_2_root_r115_SUM_20_), .B_19_(add_2_root_r115_SUM_19_), 
        .B_18_(add_2_root_r115_SUM_18_), .B_17_(add_2_root_r115_SUM_17_), 
        .B_16_(add_2_root_r115_SUM_16_), .B_15_(add_2_root_r115_SUM_15_), 
        .B_14_(add_2_root_r115_SUM_14_), .B_13_(add_2_root_r115_SUM_13_), 
        .B_12_(add_2_root_r115_SUM_12_), .B_11_(add_2_root_r115_SUM_11_), 
        .B_10_(add_2_root_r115_SUM_10_), .B_9_(add_2_root_r115_SUM_9_), .B_8_(
        add_2_root_r115_SUM_8_), .B_7_(add_2_root_r115_SUM_7_), .B_6_(
        add_2_root_r115_SUM_6_), .B_5_(add_2_root_r115_SUM_5_), .B_4_(
        add_2_root_r115_SUM_4_), .SUM_23_(N221), .SUM_22_(N220), .SUM_21_(N219), .SUM_20_(N218), .SUM_19_(N217), .SUM_18_(N216), .SUM_17_(N215), .SUM_16_(
        N214), .SUM_15_(N213), .SUM_14_(N212), .SUM_13_(N211), .SUM_12_(N210), 
        .SUM_11_(N209), .SUM_10_(N208), .SUM_9_(N207), .SUM_8_(N206), .SUM_7_(
        N205) );
  TLATX1 neg_mul_reg_16_ ( .G(N446), .D(N456), .QN(n10) );
  TLATX1 neg_mul_reg_15_ ( .G(N446), .D(N455), .QN(n8) );
  TLATX1 neg_mul_reg_14_ ( .G(N446), .D(N454), .Q(neg_mul[14]), .QN(n6) );
  TLATX1 neg_mul_reg_13_ ( .G(N446), .D(N453), .Q(neg_mul[13]), .QN(n20) );
  TLATX1 neg_mul_reg_12_ ( .G(N446), .D(N452), .QN(n9) );
  TLATX1 neg_mul_reg_11_ ( .G(N446), .D(N451), .Q(neg_mul[11]), .QN(n5) );
  TLATX1 neg_mul_reg_23_ ( .G(N446), .D(N463), .Q(neg_mul[23]), .QN(n7) );
  TLATX1 neg_mul_reg_22_ ( .G(N446), .D(N462), .Q(neg_mul[22]), .QN(n13) );
  TLATX1 neg_mul_reg_21_ ( .G(N446), .D(N461), .Q(neg_mul[21]), .QN(n14) );
  TLATX1 neg_mul_reg_20_ ( .G(N446), .D(N460), .Q(neg_mul[20]), .QN(n15) );
  TLATX1 neg_mul_reg_19_ ( .G(N446), .D(N459), .Q(neg_mul[19]), .QN(n16) );
  TLATX1 neg_mul_reg_18_ ( .G(N446), .D(N458), .QN(n18) );
  TLATX1 neg_mul_reg_17_ ( .G(N446), .D(N457), .QN(n17) );
  TLATX1 neg_mul_reg_9_ ( .G(N446), .D(N449), .Q(neg_mul[9]), .QN(n12) );
  TLATX1 neg_mul_reg_10_ ( .G(N446), .D(N450), .Q(neg_mul[10]), .QN(n11) );
  TLATX1 neg_mul_reg_8_ ( .G(N446), .D(N448), .Q(neg_mul[8]), .QN(n19) );
  TLATX1 neg_mul_reg_7_ ( .G(N446), .D(N447), .Q(out[0]) );
  BUFX8 U2 ( .A(n82), .Y(n3) );
  XNOR2X4 U3 ( .A(n22), .B(n42), .Y(n82) );
  NOR2BX4 U4 ( .AN(n1), .B(n3), .Y(n81) );
  CLKINVX20 U5 ( .A(n80), .Y(n1) );
  NOR2X2 U6 ( .A(n28), .B(n84), .Y(n85) );
  XNOR2X2 U7 ( .A(n22), .B(n42), .Y(n84) );
  XOR2X4 U8 ( .A(n83), .B(n2), .Y(out[5]) );
  CLKINVX20 U9 ( .A(n9), .Y(n2) );
  MXI2X1 U10 ( .A(n18), .B(n35), .S0(n87), .Y(n262) );
  INVX8 U11 ( .A(n86), .Y(n87) );
  MXI2X2 U12 ( .A(n17), .B(n34), .S0(n87), .Y(out[10]) );
  BUFX3 U13 ( .A(n262), .Y(out[11]) );
  AOI211X4 U14 ( .A0(n72), .A1(n22), .B0(n71), .C0(n70), .Y(out[2]) );
  CLKINVX8 U15 ( .A(n44), .Y(n42) );
  INVX4 U16 ( .A(in_8bit[7]), .Y(n44) );
  MX2X1 U17 ( .A(neg_mul[21]), .B(N479), .S0(n87), .Y(out[14]) );
  NAND2X1 U18 ( .A(n42), .B(n12), .Y(n66) );
  MX2X1 U19 ( .A(neg_mul[22]), .B(N480), .S0(n87), .Y(out[15]) );
  OAI21XL U20 ( .A0(n42), .A1(n75), .B0(n74), .Y(n79) );
  NAND2X1 U21 ( .A(n42), .B(n11), .Y(n74) );
  INVX1 U22 ( .A(n97), .Y(n93) );
  CLKINVX3 U23 ( .A(n58), .Y(n54) );
  CLKINVX3 U24 ( .A(n44), .Y(n43) );
  XNOR2X1 U25 ( .A(neg_mul[23]), .B(n37), .Y(n21) );
  NOR2X4 U26 ( .A(n22), .B(n77), .Y(n78) );
  XOR2X4 U27 ( .A(n81), .B(neg_mul[11]), .Y(out[4]) );
  OAI21X2 U28 ( .A0(n42), .A1(n61), .B0(n60), .Y(n65) );
  XOR2X4 U29 ( .A(n85), .B(neg_mul[13]), .Y(out[6]) );
  INVX1 U30 ( .A(n52), .Y(n51) );
  NOR2X2 U31 ( .A(n22), .B(n69), .Y(n71) );
  XOR2X4 U32 ( .A(n23), .B(neg_mul[14]), .Y(out[7]) );
  NOR2X2 U33 ( .A(n22), .B(n63), .Y(n64) );
  BUFX20 U34 ( .A(in_17bit[16]), .Y(n22) );
  AOI211X2 U35 ( .A0(n55), .A1(n65), .B0(n64), .C0(n36), .Y(out[1]) );
  INVXL U36 ( .A(in_17bit[16]), .Y(n52) );
  INVX4 U37 ( .A(n58), .Y(n55) );
  CLKINVX8 U38 ( .A(n22), .Y(n58) );
  NOR2X4 U39 ( .A(n27), .B(n3), .Y(n83) );
  NOR2X4 U40 ( .A(n86), .B(n33), .Y(n24) );
  XNOR2X4 U41 ( .A(n22), .B(n42), .Y(n86) );
  XNOR2X4 U42 ( .A(n24), .B(n10), .Y(out[9]) );
  AOI2BB2X1 U43 ( .B0(n68), .B1(n42), .A0N(n43), .A1N(neg_mul[9]), .Y(n69) );
  AOI2BB2X1 U44 ( .B0(n62), .B1(n42), .A0N(n43), .A1N(neg_mul[8]), .Y(n63) );
  NAND2X1 U45 ( .A(n42), .B(n19), .Y(n60) );
  AOI2BB2X1 U46 ( .B0(n76), .B1(n42), .A0N(n43), .A1N(neg_mul[10]), .Y(n77) );
  MX2X4 U47 ( .A(neg_mul[19]), .B(N477), .S0(n87), .Y(out[12]) );
  MX2X4 U48 ( .A(neg_mul[20]), .B(N478), .S0(n87), .Y(out[13]) );
  AND3X1 U49 ( .A(in_8bit[2]), .B(n49), .C(n47), .Y(n32) );
  INVX1 U50 ( .A(n211), .Y(in_17bit_b[1]) );
  INVX1 U51 ( .A(n250), .Y(in_17bit_b[14]) );
  INVX1 U52 ( .A(n247), .Y(in_17bit_b[13]) );
  INVX1 U53 ( .A(n214), .Y(in_17bit_b[2]) );
  INVX1 U54 ( .A(n223), .Y(in_17bit_b[5]) );
  INVX1 U55 ( .A(n226), .Y(in_17bit_b[6]) );
  INVX1 U56 ( .A(n229), .Y(in_17bit_b[7]) );
  INVX1 U57 ( .A(n232), .Y(in_17bit_b[8]) );
  INVX1 U58 ( .A(n235), .Y(in_17bit_b[9]) );
  INVX1 U59 ( .A(n238), .Y(in_17bit_b[10]) );
  INVX1 U60 ( .A(n241), .Y(in_17bit_b[11]) );
  INVX1 U61 ( .A(n244), .Y(in_17bit_b[12]) );
  INVX1 U62 ( .A(n220), .Y(in_17bit_b[4]) );
  INVX1 U63 ( .A(n217), .Y(in_17bit_b[3]) );
  NOR2X4 U64 ( .A(n29), .B(n3), .Y(n23) );
  OAI21XL U65 ( .A0(n42), .A1(n67), .B0(n66), .Y(n72) );
  NAND3XL U66 ( .A(n43), .B(n45), .C(n48), .Y(n96) );
  INVX1 U67 ( .A(n48), .Y(n47) );
  INVX1 U68 ( .A(n179), .Y(n260) );
  OAI21XL U69 ( .A0(n260), .A1(n261), .B0(n259), .Y(N463) );
  AOI22X1 U70 ( .A0(N221), .A1(n40), .B0(N363), .B1(n39), .Y(n259) );
  ADDFX2 U71 ( .A(n41), .B(in_17bit_b[12]), .CI(add_1_root_r112_carry_16_), 
        .CO(add_1_root_r112_carry_17_), .S(add_1_root_r112_SUM_16_) );
  ADDFX2 U72 ( .A(add_1_root_r119_A_19_), .B(in_17bit_b[13]), .CI(
        add_1_root_r119_carry[19]), .CO(add_1_root_r119_carry[20]), .S(
        add_1_root_r119_SUM_19_) );
  ADDFX2 U73 ( .A(n41), .B(in_17bit_b[15]), .CI(add_3_root_r119_carry_17_), 
        .CO(add_3_root_r119_carry_18_), .S(add_1_root_r119_A_17_) );
  ADDFX2 U74 ( .A(n41), .B(in_17bit_b[14]), .CI(add_2_root_r115_carry_17_), 
        .CO(add_2_root_r115_carry_18_), .S(add_2_root_r115_SUM_17_) );
  ADDFX2 U75 ( .A(n41), .B(in_17bit_b[14]), .CI(add_1_root_r115_carry_20_), 
        .CO(add_1_root_r115_carry_21_), .S(add_1_root_r115_SUM_20_) );
  ADDFX2 U76 ( .A(n41), .B(in_17bit_b[15]), .CI(add_2_root_r119_carry_20_), 
        .CO(add_2_root_r119_carry_21_), .S(add_2_root_r119_SUM_20_) );
  ADDFX2 U77 ( .A(in_17bit_b[3]), .B(in_17bit_b[1]), .CI(
        add_2_root_r115_carry_4_), .CO(add_2_root_r115_carry_5_), .S(
        add_2_root_r115_SUM_4_) );
  ADDFX2 U78 ( .A(in_17bit_b[4]), .B(in_17bit_b[2]), .CI(
        add_2_root_r115_carry_5_), .CO(add_2_root_r115_carry_6_), .S(
        add_2_root_r115_SUM_5_) );
  ADDFX2 U79 ( .A(in_17bit_b[5]), .B(in_17bit_b[1]), .CI(
        add_1_root_r112_carry_5_), .CO(add_1_root_r112_carry_6_), .S(
        add_1_root_r112_SUM_5_) );
  ADDFX2 U80 ( .A(in_17bit_b[6]), .B(in_17bit_b[5]), .CI(
        add_3_root_r119_carry_7_), .CO(add_3_root_r119_carry_8_), .S(
        add_1_root_r119_A_7_) );
  ADDFX2 U81 ( .A(in_17bit_b[6]), .B(in_17bit_b[2]), .CI(
        add_1_root_r112_carry_6_), .CO(add_1_root_r112_carry_7_), .S(
        add_1_root_r112_SUM_6_) );
  ADDFX2 U82 ( .A(in_17bit_b[3]), .B(in_17bit_b[1]), .CI(
        add_1_root_r115_carry_7_), .CO(add_1_root_r115_carry_8_), .S(
        add_1_root_r115_SUM_7_) );
  ADDFX2 U83 ( .A(in_17bit_b[7]), .B(in_17bit_b[6]), .CI(
        add_3_root_r119_carry_8_), .CO(add_3_root_r119_carry_9_), .S(
        add_1_root_r119_A_8_) );
  ADDFX2 U84 ( .A(add_1_root_r119_A_7_), .B(in_17bit_b[1]), .CI(
        add_1_root_r119_carry[7]), .CO(add_1_root_r119_carry[8]), .S(
        add_1_root_r119_SUM_7_) );
  ADDFX2 U85 ( .A(in_17bit_b[2]), .B(in_17bit_b[1]), .CI(
        add_2_root_r119_carry_6_), .CO(add_2_root_r119_carry_7_), .S(
        add_2_root_r119_SUM_6_) );
  ADDFX2 U86 ( .A(in_17bit_b[4]), .B(in_17bit_b[2]), .CI(
        add_1_root_r115_carry_8_), .CO(add_1_root_r115_carry_9_), .S(
        add_1_root_r115_SUM_8_) );
  ADDFX2 U87 ( .A(in_17bit_b[8]), .B(in_17bit_b[7]), .CI(
        add_3_root_r119_carry_9_), .CO(add_3_root_r119_carry_10_), .S(
        add_1_root_r119_A_9_) );
  ADDFX2 U88 ( .A(add_1_root_r119_A_8_), .B(in_17bit_b[2]), .CI(
        add_1_root_r119_carry[8]), .CO(add_1_root_r119_carry[9]), .S(
        add_1_root_r119_SUM_8_) );
  ADDFX2 U89 ( .A(in_17bit_b[3]), .B(in_17bit_b[2]), .CI(
        add_2_root_r119_carry_7_), .CO(add_2_root_r119_carry_8_), .S(
        add_2_root_r119_SUM_7_) );
  ADDFX2 U90 ( .A(in_17bit_b[6]), .B(in_17bit_b[4]), .CI(
        add_2_root_r115_carry_7_), .CO(add_2_root_r115_carry_8_), .S(
        add_2_root_r115_SUM_7_) );
  ADDFX2 U91 ( .A(in_17bit_b[8]), .B(in_17bit_b[4]), .CI(
        add_1_root_r112_carry_8_), .CO(add_1_root_r112_carry_9_), .S(
        add_1_root_r112_SUM_8_) );
  ADDFX2 U92 ( .A(in_17bit_b[9]), .B(in_17bit_b[8]), .CI(
        add_3_root_r119_carry_10_), .CO(add_3_root_r119_carry_11_), .S(
        add_1_root_r119_A_10_) );
  ADDFX2 U93 ( .A(in_17bit_b[7]), .B(in_17bit_b[5]), .CI(
        add_2_root_r115_carry_8_), .CO(add_2_root_r115_carry_9_), .S(
        add_2_root_r115_SUM_8_) );
  ADDFX2 U94 ( .A(in_17bit_b[9]), .B(in_17bit_b[5]), .CI(
        add_1_root_r112_carry_9_), .CO(add_1_root_r112_carry_10_), .S(
        add_1_root_r112_SUM_9_) );
  ADDFX2 U95 ( .A(in_17bit_b[6]), .B(in_17bit_b[4]), .CI(
        add_1_root_r115_carry_10_), .CO(add_1_root_r115_carry_11_), .S(
        add_1_root_r115_SUM_10_) );
  ADDFX2 U96 ( .A(add_1_root_r119_A_10_), .B(in_17bit_b[4]), .CI(
        add_1_root_r119_carry[10]), .CO(add_1_root_r119_carry[11]), .S(
        add_1_root_r119_SUM_10_) );
  ADDFX2 U97 ( .A(in_17bit_b[5]), .B(in_17bit_b[4]), .CI(
        add_2_root_r119_carry_9_), .CO(add_2_root_r119_carry_10_), .S(
        add_2_root_r119_SUM_9_) );
  ADDFX2 U98 ( .A(in_17bit_b[8]), .B(in_17bit_b[6]), .CI(
        add_2_root_r115_carry_9_), .CO(add_2_root_r115_carry_10_), .S(
        add_2_root_r115_SUM_9_) );
  ADDFX2 U99 ( .A(in_17bit_b[10]), .B(in_17bit_b[6]), .CI(
        add_1_root_r112_carry_10_), .CO(add_1_root_r112_carry_11_), .S(
        add_1_root_r112_SUM_10_) );
  ADDFX2 U100 ( .A(in_17bit_b[7]), .B(in_17bit_b[5]), .CI(
        add_1_root_r115_carry_11_), .CO(add_1_root_r115_carry_12_), .S(
        add_1_root_r115_SUM_11_) );
  ADDFX2 U101 ( .A(in_17bit_b[11]), .B(in_17bit_b[10]), .CI(
        add_3_root_r119_carry_12_), .CO(add_3_root_r119_carry_13_), .S(
        add_1_root_r119_A_12_) );
  ADDFX2 U102 ( .A(add_1_root_r119_A_11_), .B(in_17bit_b[5]), .CI(
        add_1_root_r119_carry[11]), .CO(add_1_root_r119_carry[12]), .S(
        add_1_root_r119_SUM_11_) );
  ADDFX2 U103 ( .A(in_17bit_b[6]), .B(in_17bit_b[5]), .CI(
        add_2_root_r119_carry_10_), .CO(add_2_root_r119_carry_11_), .S(
        add_2_root_r119_SUM_10_) );
  ADDFX2 U104 ( .A(in_17bit_b[9]), .B(in_17bit_b[7]), .CI(
        add_2_root_r115_carry_10_), .CO(add_2_root_r115_carry_11_), .S(
        add_2_root_r115_SUM_10_) );
  ADDFX2 U105 ( .A(in_17bit_b[11]), .B(in_17bit_b[7]), .CI(
        add_1_root_r112_carry_11_), .CO(add_1_root_r112_carry_12_), .S(
        add_1_root_r112_SUM_11_) );
  ADDFX2 U106 ( .A(in_17bit_b[8]), .B(in_17bit_b[6]), .CI(
        add_1_root_r115_carry_12_), .CO(add_1_root_r115_carry_13_), .S(
        add_1_root_r115_SUM_12_) );
  ADDFX2 U107 ( .A(in_17bit_b[12]), .B(in_17bit_b[11]), .CI(
        add_3_root_r119_carry_13_), .CO(add_3_root_r119_carry_14_), .S(
        add_1_root_r119_A_13_) );
  ADDFX2 U108 ( .A(add_1_root_r119_A_12_), .B(in_17bit_b[6]), .CI(
        add_1_root_r119_carry[12]), .CO(add_1_root_r119_carry[13]), .S(
        add_1_root_r119_SUM_12_) );
  ADDFX2 U109 ( .A(in_17bit_b[7]), .B(in_17bit_b[6]), .CI(
        add_2_root_r119_carry_11_), .CO(add_2_root_r119_carry_12_), .S(
        add_2_root_r119_SUM_11_) );
  ADDFX2 U110 ( .A(in_17bit_b[10]), .B(in_17bit_b[8]), .CI(
        add_2_root_r115_carry_11_), .CO(add_2_root_r115_carry_12_), .S(
        add_2_root_r115_SUM_11_) );
  ADDFX2 U111 ( .A(in_17bit_b[12]), .B(in_17bit_b[8]), .CI(
        add_1_root_r112_carry_12_), .CO(add_1_root_r112_carry_13_), .S(
        add_1_root_r112_SUM_12_) );
  ADDFX2 U112 ( .A(in_17bit_b[9]), .B(in_17bit_b[7]), .CI(
        add_1_root_r115_carry_13_), .CO(add_1_root_r115_carry_14_), .S(
        add_1_root_r115_SUM_13_) );
  ADDFX2 U113 ( .A(in_17bit_b[13]), .B(in_17bit_b[12]), .CI(
        add_3_root_r119_carry_14_), .CO(add_3_root_r119_carry_15_), .S(
        add_1_root_r119_A_14_) );
  ADDFX2 U114 ( .A(add_1_root_r119_A_13_), .B(in_17bit_b[7]), .CI(
        add_1_root_r119_carry[13]), .CO(add_1_root_r119_carry[14]), .S(
        add_1_root_r119_SUM_13_) );
  ADDFX2 U115 ( .A(in_17bit_b[8]), .B(in_17bit_b[7]), .CI(
        add_2_root_r119_carry_12_), .CO(add_2_root_r119_carry_13_), .S(
        add_2_root_r119_SUM_12_) );
  ADDFX2 U116 ( .A(in_17bit_b[11]), .B(in_17bit_b[9]), .CI(
        add_2_root_r115_carry_12_), .CO(add_2_root_r115_carry_13_), .S(
        add_2_root_r115_SUM_12_) );
  ADDFX2 U117 ( .A(in_17bit_b[13]), .B(in_17bit_b[9]), .CI(
        add_1_root_r112_carry_13_), .CO(add_1_root_r112_carry_14_), .S(
        add_1_root_r112_SUM_13_) );
  ADDFX2 U118 ( .A(in_17bit_b[10]), .B(in_17bit_b[8]), .CI(
        add_1_root_r115_carry_14_), .CO(add_1_root_r115_carry_15_), .S(
        add_1_root_r115_SUM_14_) );
  ADDFX2 U119 ( .A(in_17bit_b[14]), .B(in_17bit_b[13]), .CI(
        add_3_root_r119_carry_15_), .CO(add_3_root_r119_carry_16_), .S(
        add_1_root_r119_A_15_) );
  ADDFX2 U120 ( .A(add_1_root_r119_A_14_), .B(in_17bit_b[8]), .CI(
        add_1_root_r119_carry[14]), .CO(add_1_root_r119_carry[15]), .S(
        add_1_root_r119_SUM_14_) );
  ADDFX2 U121 ( .A(in_17bit_b[9]), .B(in_17bit_b[8]), .CI(
        add_2_root_r119_carry_13_), .CO(add_2_root_r119_carry_14_), .S(
        add_2_root_r119_SUM_13_) );
  ADDFX2 U122 ( .A(in_17bit_b[12]), .B(in_17bit_b[10]), .CI(
        add_2_root_r115_carry_13_), .CO(add_2_root_r115_carry_14_), .S(
        add_2_root_r115_SUM_13_) );
  ADDFX2 U123 ( .A(in_17bit_b[14]), .B(in_17bit_b[10]), .CI(
        add_1_root_r112_carry_14_), .CO(add_1_root_r112_carry_15_), .S(
        add_1_root_r112_SUM_14_) );
  ADDFX2 U124 ( .A(in_17bit_b[11]), .B(in_17bit_b[9]), .CI(
        add_1_root_r115_carry_15_), .CO(add_1_root_r115_carry_16_), .S(
        add_1_root_r115_SUM_15_) );
  ADDFX2 U125 ( .A(add_1_root_r119_A_15_), .B(in_17bit_b[9]), .CI(
        add_1_root_r119_carry[15]), .CO(add_1_root_r119_carry[16]), .S(
        add_1_root_r119_SUM_15_) );
  ADDFX2 U126 ( .A(in_17bit_b[10]), .B(in_17bit_b[9]), .CI(
        add_2_root_r119_carry_14_), .CO(add_2_root_r119_carry_15_), .S(
        add_2_root_r119_SUM_14_) );
  ADDFX2 U127 ( .A(in_17bit_b[13]), .B(in_17bit_b[11]), .CI(
        add_2_root_r115_carry_14_), .CO(add_2_root_r115_carry_15_), .S(
        add_2_root_r115_SUM_14_) );
  ADDFX2 U128 ( .A(in_17bit_b[15]), .B(in_17bit_b[11]), .CI(
        add_1_root_r112_carry_15_), .CO(add_1_root_r112_carry_16_), .S(
        add_1_root_r112_SUM_15_) );
  ADDFX2 U129 ( .A(in_17bit_b[12]), .B(in_17bit_b[10]), .CI(
        add_1_root_r115_carry_16_), .CO(add_1_root_r115_carry_17_), .S(
        add_1_root_r115_SUM_16_) );
  ADDFX2 U130 ( .A(add_1_root_r119_A_16_), .B(in_17bit_b[10]), .CI(
        add_1_root_r119_carry[16]), .CO(add_1_root_r119_carry[17]), .S(
        add_1_root_r119_SUM_16_) );
  ADDFX2 U131 ( .A(in_17bit_b[11]), .B(in_17bit_b[10]), .CI(
        add_2_root_r119_carry_15_), .CO(add_2_root_r119_carry_16_), .S(
        add_2_root_r119_SUM_15_) );
  ADDFX2 U132 ( .A(in_17bit_b[14]), .B(in_17bit_b[12]), .CI(
        add_2_root_r115_carry_15_), .CO(add_2_root_r115_carry_16_), .S(
        add_2_root_r115_SUM_15_) );
  ADDFX2 U133 ( .A(in_17bit_b[13]), .B(in_17bit_b[11]), .CI(
        add_1_root_r115_carry_17_), .CO(add_1_root_r115_carry_18_), .S(
        add_1_root_r115_SUM_17_) );
  ADDFX2 U134 ( .A(add_1_root_r119_A_17_), .B(in_17bit_b[11]), .CI(
        add_1_root_r119_carry[17]), .CO(add_1_root_r119_carry[18]), .S(
        add_1_root_r119_SUM_17_) );
  ADDFX2 U135 ( .A(in_17bit_b[12]), .B(in_17bit_b[11]), .CI(
        add_2_root_r119_carry_16_), .CO(add_2_root_r119_carry_17_), .S(
        add_2_root_r119_SUM_16_) );
  ADDFX2 U136 ( .A(in_17bit_b[14]), .B(in_17bit_b[12]), .CI(
        add_1_root_r115_carry_18_), .CO(add_1_root_r115_carry_19_), .S(
        add_1_root_r115_SUM_18_) );
  ADDFX2 U137 ( .A(add_1_root_r119_A_18_), .B(in_17bit_b[12]), .CI(
        add_1_root_r119_carry[18]), .CO(add_1_root_r119_carry[19]), .S(
        add_1_root_r119_SUM_18_) );
  ADDFX2 U138 ( .A(in_17bit_b[15]), .B(in_17bit_b[14]), .CI(
        add_3_root_r119_carry_16_), .CO(add_3_root_r119_carry_17_), .S(
        add_1_root_r119_A_16_) );
  ADDFX2 U139 ( .A(in_17bit_b[13]), .B(in_17bit_b[12]), .CI(
        add_2_root_r119_carry_17_), .CO(add_2_root_r119_carry_18_), .S(
        add_2_root_r119_SUM_17_) );
  ADDFX2 U140 ( .A(in_17bit_b[5]), .B(in_17bit_b[3]), .CI(
        add_2_root_r115_carry_6_), .CO(add_2_root_r115_carry_7_), .S(
        add_2_root_r115_SUM_6_) );
  ADDFX2 U141 ( .A(in_17bit_b[7]), .B(in_17bit_b[3]), .CI(
        add_1_root_r112_carry_7_), .CO(add_1_root_r112_carry_8_), .S(
        add_1_root_r112_SUM_7_) );
  ADDFX2 U142 ( .A(in_17bit_b[10]), .B(in_17bit_b[9]), .CI(
        add_3_root_r119_carry_11_), .CO(add_3_root_r119_carry_12_), .S(
        add_1_root_r119_A_11_) );
  ADDFX2 U143 ( .A(in_17bit_b[15]), .B(in_17bit_b[13]), .CI(
        add_1_root_r115_carry_19_), .CO(add_1_root_r115_carry_20_), .S(
        add_1_root_r115_SUM_19_) );
  ADDFX2 U144 ( .A(in_17bit_b[14]), .B(in_17bit_b[13]), .CI(
        add_2_root_r119_carry_18_), .CO(add_2_root_r119_carry_19_), .S(
        add_2_root_r119_SUM_18_) );
  ADDFX2 U145 ( .A(add_1_root_r119_A_9_), .B(in_17bit_b[3]), .CI(
        add_1_root_r119_carry[9]), .CO(add_1_root_r119_carry[10]), .S(
        add_1_root_r119_SUM_9_) );
  ADDFX2 U146 ( .A(in_17bit_b[4]), .B(in_17bit_b[3]), .CI(
        add_2_root_r119_carry_8_), .CO(add_2_root_r119_carry_9_), .S(
        add_2_root_r119_SUM_8_) );
  ADDFX2 U147 ( .A(in_17bit_b[3]), .B(in_17bit_b[2]), .CI(
        add_3_root_r119_carry_4_), .CO(add_3_root_r119_carry_5_), .S(
        add_1_root_r119_A_4_) );
  ADDFX2 U148 ( .A(in_17bit_b[2]), .B(in_17bit_b[1]), .CI(
        add_3_root_r119_carry_3_), .CO(add_3_root_r119_carry_4_), .S(
        add_1_root_r119_A_3_) );
  ADDFX2 U149 ( .A(in_17bit_b[15]), .B(in_17bit_b[13]), .CI(
        add_2_root_r115_carry_16_), .CO(add_2_root_r115_carry_17_), .S(
        add_2_root_r115_SUM_16_) );
  ADDFX2 U150 ( .A(in_17bit_b[5]), .B(in_17bit_b[3]), .CI(
        add_1_root_r115_carry_9_), .CO(add_1_root_r115_carry_10_), .S(
        add_1_root_r115_SUM_9_) );
  ADDFX2 U151 ( .A(in_17bit_b[5]), .B(in_17bit_b[4]), .CI(
        add_3_root_r119_carry_6_), .CO(add_3_root_r119_carry_7_), .S(
        add_1_root_r119_A_6_) );
  ADDFX2 U152 ( .A(in_17bit_b[4]), .B(in_17bit_b[3]), .CI(
        add_3_root_r119_carry_5_), .CO(add_3_root_r119_carry_6_), .S(
        add_1_root_r119_A_5_) );
  ADDFX2 U153 ( .A(in_17bit_b[15]), .B(in_17bit_b[14]), .CI(
        add_2_root_r119_carry_19_), .CO(add_2_root_r119_carry_20_), .S(
        add_2_root_r119_SUM_19_) );
  BUFX3 U154 ( .A(in_17bit_b[16]), .Y(n41) );
  INVX1 U155 ( .A(n261), .Y(in_17bit_b[16]) );
  NAND2X1 U156 ( .A(n252), .B(n251), .Y(N461) );
  AOI22X1 U157 ( .A0(N122), .A1(n254), .B0(N219), .B1(n40), .Y(n251) );
  AOI22X1 U158 ( .A0(N361), .A1(n39), .B0(n179), .B1(in_17bit_b[14]), .Y(n252)
         );
  NAND2X1 U159 ( .A(n256), .B(n255), .Y(N462) );
  AOI22X1 U160 ( .A0(N123), .A1(n254), .B0(N220), .B1(n40), .Y(n255) );
  AOI22X1 U161 ( .A0(N362), .A1(n39), .B0(n179), .B1(in_17bit_b[15]), .Y(n256)
         );
  INVX1 U162 ( .A(in_8bit[0]), .Y(n46) );
  INVX1 U163 ( .A(in_8bit[4]), .Y(n45) );
  INVX1 U164 ( .A(n51), .Y(n57) );
  INVX1 U165 ( .A(n51), .Y(n56) );
  INVX1 U166 ( .A(in_8bit[3]), .Y(n49) );
  INVX1 U167 ( .A(in_8bit[5]), .Y(n48) );
  NOR3X1 U168 ( .A(n180), .B(n49), .C(n46), .Y(n206) );
  CLKINVX3 U169 ( .A(n208), .Y(in_17bit_b[0]) );
  NAND3BX1 U170 ( .AN(n47), .B(n180), .C(in_8bit[3]), .Y(n201) );
  NAND3X1 U171 ( .A(n205), .B(n47), .C(n89), .Y(n90) );
  NOR2XL U172 ( .A(n42), .B(n45), .Y(n89) );
  NAND2XL U173 ( .A(N29), .B(n50), .Y(n261) );
  CLKINVX3 U174 ( .A(n253), .Y(in_17bit_b[15]) );
  BUFX3 U175 ( .A(n257), .Y(n39) );
  OAI2BB1X1 U176 ( .A0N(n25), .A1N(n32), .B0(n94), .Y(n257) );
  NAND2BX1 U177 ( .AN(n201), .B(n31), .Y(n94) );
  BUFX3 U178 ( .A(n258), .Y(n40) );
  OAI2BB1X1 U179 ( .A0N(n32), .A1N(n31), .B0(n95), .Y(n258) );
  NAND2BX1 U180 ( .AN(n201), .B(n25), .Y(n95) );
  OAI2BB1X1 U181 ( .A0N(n92), .A1N(n91), .B0(n90), .Y(n254) );
  NOR2BX1 U182 ( .AN(in_8bit[1]), .B(n96), .Y(n91) );
  NOR2BX1 U183 ( .AN(n206), .B(n88), .Y(n92) );
  OAI2BB1X1 U184 ( .A0N(n205), .A1N(n99), .B0(n98), .Y(n179) );
  INVX1 U185 ( .A(n96), .Y(n99) );
  NAND3BX1 U186 ( .AN(n97), .B(n206), .C(n47), .Y(n98) );
  AND2X2 U187 ( .A(n93), .B(n46), .Y(n25) );
  NAND2X1 U188 ( .A(n210), .B(n209), .Y(N447) );
  AOI22X1 U189 ( .A0(N108), .A1(n254), .B0(N205), .B1(n40), .Y(n209) );
  AOI22X1 U190 ( .A0(N347), .A1(n39), .B0(n179), .B1(in_17bit_b[0]), .Y(n210)
         );
  NAND2X1 U191 ( .A(n213), .B(n212), .Y(N448) );
  AOI22X1 U192 ( .A0(N109), .A1(n254), .B0(N206), .B1(n40), .Y(n212) );
  AOI22X1 U193 ( .A0(N348), .A1(n39), .B0(n179), .B1(n178), .Y(n213) );
  INVX1 U194 ( .A(n211), .Y(n178) );
  NAND2X1 U195 ( .A(n216), .B(n215), .Y(N449) );
  AOI22X1 U196 ( .A0(N110), .A1(n254), .B0(N207), .B1(n40), .Y(n215) );
  AOI22X1 U197 ( .A0(N349), .A1(n39), .B0(n179), .B1(in_17bit_b[2]), .Y(n216)
         );
  NAND2X1 U198 ( .A(n219), .B(n218), .Y(N450) );
  AOI22X1 U199 ( .A0(N111), .A1(n254), .B0(N208), .B1(n40), .Y(n218) );
  AOI22X1 U200 ( .A0(N350), .A1(n39), .B0(n179), .B1(in_17bit_b[3]), .Y(n219)
         );
  NAND2X1 U201 ( .A(n222), .B(n221), .Y(N451) );
  AOI22X1 U202 ( .A0(N112), .A1(n254), .B0(N209), .B1(n40), .Y(n221) );
  AOI22X1 U203 ( .A0(N351), .A1(n39), .B0(n179), .B1(in_17bit_b[4]), .Y(n222)
         );
  NAND2X1 U204 ( .A(n225), .B(n224), .Y(N452) );
  AOI22X1 U205 ( .A0(N113), .A1(n254), .B0(N210), .B1(n40), .Y(n224) );
  AOI22X1 U206 ( .A0(N352), .A1(n39), .B0(n179), .B1(in_17bit_b[5]), .Y(n225)
         );
  NAND2X1 U207 ( .A(n228), .B(n227), .Y(N453) );
  AOI22X1 U208 ( .A0(N114), .A1(n254), .B0(N211), .B1(n40), .Y(n227) );
  AOI22X1 U209 ( .A0(N353), .A1(n39), .B0(n179), .B1(in_17bit_b[6]), .Y(n228)
         );
  NAND2X1 U210 ( .A(n231), .B(n230), .Y(N454) );
  AOI22X1 U211 ( .A0(N115), .A1(n254), .B0(N212), .B1(n40), .Y(n230) );
  AOI22X1 U212 ( .A0(N354), .A1(n39), .B0(n179), .B1(in_17bit_b[7]), .Y(n231)
         );
  NAND2X1 U213 ( .A(n234), .B(n233), .Y(N455) );
  AOI22X1 U214 ( .A0(N116), .A1(n254), .B0(N213), .B1(n40), .Y(n233) );
  AOI22X1 U215 ( .A0(N355), .A1(n39), .B0(n179), .B1(in_17bit_b[8]), .Y(n234)
         );
  NAND2X1 U216 ( .A(n237), .B(n236), .Y(N456) );
  AOI22X1 U217 ( .A0(N117), .A1(n254), .B0(N214), .B1(n40), .Y(n236) );
  AOI22X1 U218 ( .A0(N356), .A1(n39), .B0(n179), .B1(in_17bit_b[9]), .Y(n237)
         );
  NAND2X1 U219 ( .A(n240), .B(n239), .Y(N457) );
  AOI22X1 U220 ( .A0(N118), .A1(n254), .B0(N215), .B1(n40), .Y(n239) );
  AOI22X1 U221 ( .A0(N357), .A1(n39), .B0(n179), .B1(in_17bit_b[10]), .Y(n240)
         );
  NAND2X1 U222 ( .A(n243), .B(n242), .Y(N458) );
  AOI22X1 U223 ( .A0(N119), .A1(n254), .B0(N216), .B1(n40), .Y(n242) );
  AOI22X1 U224 ( .A0(N358), .A1(n39), .B0(n179), .B1(in_17bit_b[11]), .Y(n243)
         );
  NAND2X1 U225 ( .A(n246), .B(n245), .Y(N459) );
  AOI22X1 U226 ( .A0(N120), .A1(n254), .B0(N217), .B1(n40), .Y(n245) );
  AOI22X1 U227 ( .A0(N359), .A1(n39), .B0(n179), .B1(in_17bit_b[12]), .Y(n246)
         );
  NAND2X1 U228 ( .A(n249), .B(n248), .Y(N460) );
  AOI22X1 U229 ( .A0(N121), .A1(n254), .B0(N218), .B1(n40), .Y(n248) );
  AOI22X1 U230 ( .A0(N360), .A1(n39), .B0(n179), .B1(in_17bit_b[13]), .Y(n249)
         );
  INVX1 U231 ( .A(n73), .Y(n70) );
  MXI2XL U232 ( .A(n7), .B(n21), .S0(n87), .Y(out[16]) );
  XOR2X4 U233 ( .A(n26), .B(n8), .Y(out[8]) );
  OR2X2 U234 ( .A(n86), .B(n30), .Y(n26) );
  NOR4BXL U235 ( .AN(n202), .B(n46), .C(in_8bit[1]), .D(in_8bit[2]), .Y(n205)
         );
  INVXL U236 ( .A(in_8bit[2]), .Y(n180) );
  NAND4BBX1 U237 ( .AN(n39), .BN(n40), .C(n207), .D(n260), .Y(N446) );
  AOI2BB1X1 U238 ( .A0N(n204), .A1N(n203), .B0(n254), .Y(n207) );
  OR4X1 U239 ( .A(in_8bit[1]), .B(in_8bit[0]), .C(in_8bit[2]), .D(in_8bit[3]), 
        .Y(n203) );
  AOI22XL U240 ( .A0(in_17bit[0]), .A1(n54), .B0(in_17bit[0]), .B1(n57), .Y(
        n208) );
  AOI22XL U241 ( .A0(N14), .A1(n54), .B0(in_17bit[1]), .B1(n57), .Y(n211) );
  AOI22XL U242 ( .A0(N15), .A1(n54), .B0(in_17bit[2]), .B1(n56), .Y(n214) );
  AOI22X1 U243 ( .A0(N27), .A1(n51), .B0(in_17bit[14]), .B1(n57), .Y(n250) );
  AOI22X1 U244 ( .A0(N28), .A1(n51), .B0(in_17bit[15]), .B1(n56), .Y(n253) );
  AOI22X1 U245 ( .A0(N16), .A1(n51), .B0(in_17bit[3]), .B1(n56), .Y(n217) );
  AOI22X1 U246 ( .A0(N17), .A1(n51), .B0(in_17bit[4]), .B1(n53), .Y(n220) );
  AOI22X1 U247 ( .A0(N18), .A1(n51), .B0(in_17bit[5]), .B1(n57), .Y(n223) );
  AOI22X1 U248 ( .A0(N19), .A1(n51), .B0(in_17bit[6]), .B1(n52), .Y(n226) );
  AOI22X1 U249 ( .A0(N26), .A1(n51), .B0(in_17bit[13]), .B1(n56), .Y(n247) );
  AOI22X1 U250 ( .A0(N20), .A1(n51), .B0(in_17bit[7]), .B1(n57), .Y(n229) );
  AOI22X1 U251 ( .A0(N21), .A1(n51), .B0(in_17bit[8]), .B1(n56), .Y(n232) );
  AOI22X1 U252 ( .A0(N22), .A1(n51), .B0(in_17bit[9]), .B1(n53), .Y(n235) );
  AOI22X1 U253 ( .A0(N23), .A1(n51), .B0(in_17bit[10]), .B1(n52), .Y(n238) );
  AOI22X1 U254 ( .A0(N24), .A1(n51), .B0(in_17bit[11]), .B1(n53), .Y(n241) );
  AOI22X1 U255 ( .A0(N25), .A1(n51), .B0(in_17bit[12]), .B1(n53), .Y(n244) );
  INVXL U256 ( .A(in_8bit[6]), .Y(n88) );
  INVX1 U257 ( .A(n59), .Y(n80) );
  NAND2BX1 U258 ( .AN(n73), .B(n11), .Y(n59) );
  NAND2X1 U259 ( .A(n36), .B(n12), .Y(n73) );
  AND2X2 U260 ( .A(n80), .B(n5), .Y(n27) );
  AND2X2 U261 ( .A(n27), .B(n9), .Y(n28) );
  AND2X2 U262 ( .A(n28), .B(n20), .Y(n29) );
  AND2X2 U263 ( .A(n29), .B(n6), .Y(n30) );
  AND4X1 U264 ( .A(in_8bit[1]), .B(n43), .C(n200), .D(n46), .Y(n31) );
  AND2X2 U265 ( .A(n30), .B(n8), .Y(n33) );
  INVX1 U266 ( .A(in_17bit[0]), .Y(n100) );
  INVX1 U267 ( .A(in_17bit[13]), .Y(n175) );
  INVX1 U268 ( .A(in_17bit[1]), .Y(n101) );
  INVX1 U269 ( .A(in_17bit[2]), .Y(n158) );
  INVX1 U270 ( .A(in_17bit[3]), .Y(n160) );
  INVX1 U271 ( .A(in_17bit[4]), .Y(n163) );
  INVX1 U272 ( .A(in_17bit[5]), .Y(n164) );
  INVX1 U273 ( .A(in_17bit[6]), .Y(n167) );
  INVX1 U274 ( .A(in_17bit[7]), .Y(n168) );
  INVX1 U275 ( .A(in_17bit[8]), .Y(n170) );
  INVX1 U276 ( .A(in_17bit[9]), .Y(n171) );
  INVX1 U277 ( .A(in_17bit[10]), .Y(n172) );
  INVX1 U278 ( .A(in_17bit[11]), .Y(n173) );
  INVX1 U279 ( .A(in_17bit[12]), .Y(n174) );
  INVX1 U280 ( .A(in_17bit[14]), .Y(n176) );
  INVX1 U281 ( .A(in_17bit[15]), .Y(n177) );
  INVXL U282 ( .A(n51), .Y(n53) );
  XNOR2X1 U283 ( .A(n17), .B(sub_add_75_b0_carry[10]), .Y(n34) );
  INVX1 U284 ( .A(n75), .Y(n76) );
  INVX1 U285 ( .A(n67), .Y(n68) );
  INVX1 U286 ( .A(n61), .Y(n62) );
  XNOR2X1 U287 ( .A(n18), .B(sub_add_75_b0_carry[11]), .Y(n35) );
  NOR2X1 U288 ( .A(out[0]), .B(neg_mul[8]), .Y(n36) );
  NAND2BX1 U289 ( .AN(n36), .B(neg_mul[9]), .Y(n67) );
  NAND2X1 U290 ( .A(out[0]), .B(neg_mul[8]), .Y(n61) );
  NAND2X1 U291 ( .A(neg_mul[10]), .B(n73), .Y(n75) );
  NAND2X1 U292 ( .A(sub_add_75_b0_carry[15]), .B(n13), .Y(n37) );
  INVXL U293 ( .A(n52), .Y(n50) );
  AOI211X4 U294 ( .A0(n22), .A1(n79), .B0(n78), .C0(n80), .Y(out[3]) );
  OR4X1 U295 ( .A(in_8bit[4]), .B(n47), .C(in_8bit[6]), .D(n43), .Y(n204) );
  NOR2XL U296 ( .A(in_8bit[6]), .B(in_8bit[3]), .Y(n202) );
  NOR2XL U297 ( .A(in_8bit[6]), .B(in_8bit[4]), .Y(n200) );
  NAND4BXL U298 ( .AN(n43), .B(in_8bit[4]), .C(in_8bit[1]), .D(in_8bit[6]), 
        .Y(n97) );
  AND2X1 U299 ( .A(add_1_root_r112_carry_20_), .B(n41), .Y(
        add_1_root_r112_SUM_21_) );
  XOR2X1 U300 ( .A(n41), .B(add_1_root_r112_carry_20_), .Y(
        add_1_root_r112_SUM_20_) );
  AND2X1 U301 ( .A(add_1_root_r112_carry_19_), .B(in_17bit_b[15]), .Y(
        add_1_root_r112_carry_20_) );
  XOR2X1 U302 ( .A(in_17bit_b[15]), .B(add_1_root_r112_carry_19_), .Y(
        add_1_root_r112_SUM_19_) );
  AND2X1 U303 ( .A(add_1_root_r112_carry_18_), .B(in_17bit_b[14]), .Y(
        add_1_root_r112_carry_19_) );
  XOR2X1 U304 ( .A(in_17bit_b[14]), .B(add_1_root_r112_carry_18_), .Y(
        add_1_root_r112_SUM_18_) );
  AND2X1 U305 ( .A(add_1_root_r112_carry_17_), .B(in_17bit_b[13]), .Y(
        add_1_root_r112_carry_18_) );
  XOR2X1 U306 ( .A(in_17bit_b[13]), .B(add_1_root_r112_carry_17_), .Y(
        add_1_root_r112_SUM_17_) );
  AND2X1 U307 ( .A(add_2_root_r119_carry_21_), .B(n41), .Y(
        add_2_root_r119_SUM_22_) );
  XOR2X1 U308 ( .A(n41), .B(add_2_root_r119_carry_21_), .Y(
        add_2_root_r119_SUM_21_) );
  AND2X1 U309 ( .A(in_17bit_b[1]), .B(in_17bit_b[0]), .Y(
        add_2_root_r119_carry_6_) );
  XOR2X1 U310 ( .A(in_17bit_b[0]), .B(in_17bit_b[1]), .Y(
        add_2_root_r119_SUM_5_) );
  AND2X1 U311 ( .A(add_1_root_r119_carry[22]), .B(n41), .Y(
        add_1_root_r119_SUM_23_) );
  XOR2X1 U312 ( .A(n41), .B(add_1_root_r119_carry[22]), .Y(
        add_1_root_r119_SUM_22_) );
  AND2X1 U313 ( .A(add_1_root_r119_carry[21]), .B(in_17bit_b[15]), .Y(
        add_1_root_r119_carry[22]) );
  XOR2X1 U314 ( .A(in_17bit_b[15]), .B(add_1_root_r119_carry[21]), .Y(
        add_1_root_r119_SUM_21_) );
  AND2X1 U315 ( .A(add_1_root_r119_carry[20]), .B(in_17bit_b[14]), .Y(
        add_1_root_r119_carry[21]) );
  XOR2X1 U316 ( .A(in_17bit_b[14]), .B(add_1_root_r119_carry[20]), .Y(
        add_1_root_r119_SUM_20_) );
  AND2X1 U317 ( .A(add_1_root_r119_A_6_), .B(in_17bit_b[0]), .Y(
        add_1_root_r119_carry[7]) );
  XOR2X1 U318 ( .A(in_17bit_b[0]), .B(add_1_root_r119_A_6_), .Y(
        add_1_root_r119_SUM_6_) );
  AND2X1 U319 ( .A(add_3_root_r119_carry_18_), .B(n41), .Y(
        add_1_root_r119_A_19_) );
  XOR2X1 U320 ( .A(n41), .B(add_3_root_r119_carry_18_), .Y(
        add_1_root_r119_A_18_) );
  AND2X1 U321 ( .A(in_17bit_b[1]), .B(in_17bit_b[0]), .Y(
        add_3_root_r119_carry_3_) );
  XOR2X1 U322 ( .A(in_17bit_b[0]), .B(in_17bit_b[1]), .Y(add_1_root_r119_A_2_)
         );
  AND2X1 U323 ( .A(add_2_root_r115_carry_19_), .B(n41), .Y(
        add_2_root_r115_SUM_20_) );
  XOR2X1 U324 ( .A(n41), .B(add_2_root_r115_carry_19_), .Y(
        add_2_root_r115_SUM_19_) );
  AND2X1 U325 ( .A(add_2_root_r115_carry_18_), .B(in_17bit_b[15]), .Y(
        add_2_root_r115_carry_19_) );
  XOR2X1 U326 ( .A(in_17bit_b[15]), .B(add_2_root_r115_carry_18_), .Y(
        add_2_root_r115_SUM_18_) );
  AND2X1 U327 ( .A(in_17bit_b[2]), .B(in_17bit_b[0]), .Y(
        add_2_root_r115_carry_4_) );
  XOR2X1 U328 ( .A(in_17bit_b[0]), .B(in_17bit_b[2]), .Y(
        add_2_root_r115_SUM_3_) );
  AND2X1 U329 ( .A(add_1_root_r115_carry_22_), .B(n41), .Y(
        add_1_root_r115_SUM_23_) );
  XOR2X1 U330 ( .A(n41), .B(add_1_root_r115_carry_22_), .Y(
        add_1_root_r115_SUM_22_) );
  AND2X1 U331 ( .A(add_1_root_r115_carry_21_), .B(in_17bit_b[15]), .Y(
        add_1_root_r115_carry_22_) );
  XOR2X1 U332 ( .A(in_17bit_b[15]), .B(add_1_root_r115_carry_21_), .Y(
        add_1_root_r115_SUM_21_) );
  AND2X1 U333 ( .A(in_17bit_b[2]), .B(in_17bit_b[0]), .Y(
        add_1_root_r115_carry_7_) );
  XOR2X1 U334 ( .A(in_17bit_b[0]), .B(in_17bit_b[2]), .Y(
        add_1_root_r115_SUM_6_) );
  XOR2X1 U335 ( .A(n52), .B(sub_add_54_b0_carry[16]), .Y(N29) );
  AND2X1 U336 ( .A(sub_add_54_b0_carry[15]), .B(n177), .Y(
        sub_add_54_b0_carry[16]) );
  XOR2X1 U337 ( .A(n177), .B(sub_add_54_b0_carry[15]), .Y(N28) );
  AND2X1 U338 ( .A(sub_add_54_b0_carry[14]), .B(n176), .Y(
        sub_add_54_b0_carry[15]) );
  XOR2X1 U339 ( .A(n176), .B(sub_add_54_b0_carry[14]), .Y(N27) );
  AND2X1 U340 ( .A(sub_add_54_b0_carry[13]), .B(n175), .Y(
        sub_add_54_b0_carry[14]) );
  XOR2X1 U341 ( .A(n175), .B(sub_add_54_b0_carry[13]), .Y(N26) );
  AND2X1 U342 ( .A(sub_add_54_b0_carry[12]), .B(n174), .Y(
        sub_add_54_b0_carry[13]) );
  XOR2X1 U343 ( .A(n174), .B(sub_add_54_b0_carry[12]), .Y(N25) );
  AND2X1 U344 ( .A(sub_add_54_b0_carry[11]), .B(n173), .Y(
        sub_add_54_b0_carry[12]) );
  XOR2X1 U345 ( .A(n173), .B(sub_add_54_b0_carry[11]), .Y(N24) );
  AND2X1 U346 ( .A(sub_add_54_b0_carry[10]), .B(n172), .Y(
        sub_add_54_b0_carry[11]) );
  XOR2X1 U347 ( .A(n172), .B(sub_add_54_b0_carry[10]), .Y(N23) );
  AND2X1 U348 ( .A(sub_add_54_b0_carry[9]), .B(n171), .Y(
        sub_add_54_b0_carry[10]) );
  XOR2X1 U349 ( .A(n171), .B(sub_add_54_b0_carry[9]), .Y(N22) );
  AND2X1 U350 ( .A(sub_add_54_b0_carry[8]), .B(n170), .Y(
        sub_add_54_b0_carry[9]) );
  XOR2X1 U351 ( .A(n170), .B(sub_add_54_b0_carry[8]), .Y(N21) );
  AND2X1 U352 ( .A(sub_add_54_b0_carry[7]), .B(n168), .Y(
        sub_add_54_b0_carry[8]) );
  XOR2X1 U353 ( .A(n168), .B(sub_add_54_b0_carry[7]), .Y(N20) );
  AND2X1 U354 ( .A(sub_add_54_b0_carry[6]), .B(n167), .Y(
        sub_add_54_b0_carry[7]) );
  XOR2X1 U355 ( .A(n167), .B(sub_add_54_b0_carry[6]), .Y(N19) );
  AND2X1 U356 ( .A(sub_add_54_b0_carry[5]), .B(n164), .Y(
        sub_add_54_b0_carry[6]) );
  XOR2X1 U357 ( .A(n164), .B(sub_add_54_b0_carry[5]), .Y(N18) );
  AND2X1 U358 ( .A(sub_add_54_b0_carry[4]), .B(n163), .Y(
        sub_add_54_b0_carry[5]) );
  XOR2X1 U359 ( .A(n163), .B(sub_add_54_b0_carry[4]), .Y(N17) );
  AND2X1 U360 ( .A(sub_add_54_b0_carry[3]), .B(n160), .Y(
        sub_add_54_b0_carry[4]) );
  XOR2X1 U361 ( .A(n160), .B(sub_add_54_b0_carry[3]), .Y(N16) );
  AND2X1 U362 ( .A(sub_add_54_b0_carry[2]), .B(n158), .Y(
        sub_add_54_b0_carry[3]) );
  XOR2X1 U363 ( .A(n158), .B(sub_add_54_b0_carry[2]), .Y(N15) );
  AND2X1 U364 ( .A(n100), .B(n101), .Y(sub_add_54_b0_carry[2]) );
  XOR2X1 U365 ( .A(n101), .B(n100), .Y(N14) );
  XOR2X1 U366 ( .A(n13), .B(sub_add_75_b0_carry[15]), .Y(N480) );
  AND2X1 U367 ( .A(sub_add_75_b0_carry[14]), .B(n14), .Y(
        sub_add_75_b0_carry[15]) );
  XOR2X1 U368 ( .A(n14), .B(sub_add_75_b0_carry[14]), .Y(N479) );
  AND2X1 U369 ( .A(sub_add_75_b0_carry[13]), .B(n15), .Y(
        sub_add_75_b0_carry[14]) );
  XOR2X1 U370 ( .A(n15), .B(sub_add_75_b0_carry[13]), .Y(N478) );
  AND2X1 U371 ( .A(sub_add_75_b0_carry[12]), .B(n16), .Y(
        sub_add_75_b0_carry[13]) );
  XOR2X1 U372 ( .A(n16), .B(sub_add_75_b0_carry[12]), .Y(N477) );
  AND2X1 U373 ( .A(sub_add_75_b0_carry[11]), .B(n18), .Y(
        sub_add_75_b0_carry[12]) );
  AND2X1 U374 ( .A(sub_add_75_b0_carry[10]), .B(n17), .Y(
        sub_add_75_b0_carry[11]) );
  AND2X1 U375 ( .A(n33), .B(n10), .Y(sub_add_75_b0_carry[10]) );
  AND2X1 U376 ( .A(in_17bit_b[0]), .B(in_17bit_b[4]), .Y(
        add_1_root_r112_carry_5_) );
endmodule


module butterfly_DW01_sub_14 ( A, B, DIFF );
  input [16:0] A;
  input [16:0] B;
  output [16:0] DIFF;
  wire   n152, n153, n1, n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151;

  NOR2XL U3 ( .A(n99), .B(n100), .Y(n94) );
  CLKBUFX2 U4 ( .A(A[14]), .Y(n31) );
  INVX2 U5 ( .A(n31), .Y(n109) );
  INVX8 U6 ( .A(n88), .Y(n141) );
  XNOR2X4 U7 ( .A(n116), .B(n1), .Y(DIFF[14]) );
  AND2X1 U8 ( .A(n92), .B(n106), .Y(n1) );
  NAND4X4 U9 ( .A(n30), .B(n91), .C(n94), .D(n95), .Y(n78) );
  XOR2X2 U10 ( .A(n60), .B(n61), .Y(DIFF[3]) );
  INVX4 U11 ( .A(n89), .Y(n42) );
  AOI22X4 U12 ( .A0(n18), .A1(n109), .B0(n110), .B1(n106), .Y(n101) );
  AOI21X4 U13 ( .A0(n101), .A1(n102), .B0(n103), .Y(n77) );
  INVX2 U14 ( .A(n17), .Y(n18) );
  OAI21X2 U15 ( .A0(n8), .A1(n34), .B0(n15), .Y(n22) );
  INVXL U16 ( .A(n46), .Y(n48) );
  CLKINVX2 U17 ( .A(n39), .Y(n20) );
  NAND2X2 U18 ( .A(n35), .B(n40), .Y(n132) );
  NAND2BX2 U19 ( .AN(A[1]), .B(B[1]), .Y(n146) );
  NAND4X1 U20 ( .A(n62), .B(n146), .C(n65), .D(n75), .Y(n100) );
  NAND2BX1 U21 ( .AN(B[7]), .B(A[7]), .Y(n89) );
  NAND2BX2 U22 ( .AN(B[4]), .B(A[4]), .Y(n57) );
  BUFX3 U23 ( .A(B[4]), .Y(n21) );
  INVX1 U24 ( .A(n137), .Y(n11) );
  XNOR2X1 U25 ( .A(n63), .B(n29), .Y(DIFF[2]) );
  INVX4 U26 ( .A(n23), .Y(DIFF[6]) );
  XNOR2X2 U27 ( .A(n32), .B(n7), .Y(DIFF[9]) );
  OAI2BB1X1 U28 ( .A0N(n20), .A1N(n36), .B0(n40), .Y(n32) );
  INVX1 U29 ( .A(n35), .Y(n33) );
  XNOR2X2 U30 ( .A(n138), .B(n26), .Y(DIFF[10]) );
  OAI21X2 U31 ( .A0(n8), .A1(n34), .B0(n15), .Y(n138) );
  NAND2X1 U32 ( .A(n124), .B(n96), .Y(n128) );
  CLKINVX4 U33 ( .A(n152), .Y(n2) );
  INVX8 U34 ( .A(n2), .Y(DIFF[8]) );
  XOR2X1 U35 ( .A(n19), .B(n37), .Y(n152) );
  AND2X2 U36 ( .A(n93), .B(n105), .Y(n4) );
  INVX8 U37 ( .A(n124), .Y(n39) );
  NAND2XL U38 ( .A(n89), .B(n88), .Y(n87) );
  INVX3 U39 ( .A(n44), .Y(n49) );
  INVXL U40 ( .A(n122), .Y(n13) );
  NOR2BXL U41 ( .AN(n134), .B(n123), .Y(n137) );
  OAI2BB1X1 U42 ( .A0N(n44), .A1N(n45), .B0(n46), .Y(n41) );
  CLKINVX3 U43 ( .A(n83), .Y(n95) );
  INVXL U44 ( .A(n110), .Y(n5) );
  NAND2BX1 U45 ( .AN(A[10]), .B(B[10]), .Y(n133) );
  DLY1X1 U46 ( .A(n106), .Y(n6) );
  INVX4 U47 ( .A(n145), .Y(n43) );
  NOR2BX4 U48 ( .AN(B[12]), .B(A[12]), .Y(n121) );
  OR2X2 U49 ( .A(n33), .B(n34), .Y(n7) );
  CLKINVX8 U50 ( .A(n99), .Y(n85) );
  CLKINVX3 U51 ( .A(n150), .Y(n64) );
  NAND2BX2 U52 ( .AN(B[1]), .B(A[1]), .Y(n70) );
  OAI21X4 U53 ( .A0(n82), .A1(n83), .B0(n84), .Y(n81) );
  AOI21X2 U54 ( .A0(n85), .A1(n86), .B0(n87), .Y(n82) );
  AND2X1 U55 ( .A(n92), .B(n90), .Y(n113) );
  INVX8 U56 ( .A(n90), .Y(n110) );
  BUFX4 U57 ( .A(n35), .Y(n15) );
  OAI2BB1X4 U58 ( .A0N(n113), .A1N(n112), .B0(n6), .Y(n111) );
  NAND2BX4 U59 ( .AN(A[12]), .B(B[12]), .Y(n93) );
  NAND2XL U60 ( .A(n124), .B(n96), .Y(n119) );
  AOI21X4 U61 ( .A0(n36), .A1(n20), .B0(n38), .Y(n8) );
  INVXL U62 ( .A(n135), .Y(n139) );
  BUFX8 U63 ( .A(A[10]), .Y(n9) );
  XOR2X4 U64 ( .A(n45), .B(n47), .Y(n153) );
  NAND2X4 U65 ( .A(n56), .B(n57), .Y(n53) );
  NOR2X4 U66 ( .A(n42), .B(n141), .Y(n10) );
  NAND3X4 U67 ( .A(n131), .B(n132), .C(n133), .Y(n130) );
  XNOR2X4 U68 ( .A(n136), .B(n11), .Y(DIFF[11]) );
  XNOR2X4 U69 ( .A(n111), .B(n12), .Y(DIFF[15]) );
  NAND2XL U70 ( .A(n104), .B(n91), .Y(n12) );
  OAI2BB1X4 U71 ( .A0N(n22), .A1N(n13), .B0(n135), .Y(n136) );
  NAND2X4 U72 ( .A(n14), .B(n130), .Y(n125) );
  AND2X4 U73 ( .A(n134), .B(n135), .Y(n14) );
  XNOR2X4 U74 ( .A(n76), .B(n16), .Y(DIFF[16]) );
  XOR2X4 U75 ( .A(B[16]), .B(A[16]), .Y(n16) );
  INVX8 U76 ( .A(n96), .Y(n34) );
  NAND2BX4 U77 ( .AN(A[9]), .B(B[9]), .Y(n96) );
  NAND2X4 U78 ( .A(n46), .B(n52), .Y(n143) );
  NAND2X4 U79 ( .A(n126), .B(n125), .Y(n84) );
  NAND2BX1 U80 ( .AN(A[11]), .B(B[11]), .Y(n126) );
  AND3X4 U81 ( .A(n93), .B(n90), .C(n92), .Y(n30) );
  NAND2BX1 U82 ( .AN(A[9]), .B(B[9]), .Y(n131) );
  INVX8 U83 ( .A(n151), .Y(n51) );
  INVXL U84 ( .A(B[14]), .Y(n17) );
  OAI2BB1X4 U85 ( .A0N(n85), .A1N(n58), .B0(n10), .Y(n19) );
  NAND2BX2 U86 ( .AN(A[2]), .B(B[2]), .Y(n62) );
  NAND2BXL U87 ( .AN(B[2]), .B(A[2]), .Y(n150) );
  INVX8 U88 ( .A(n98), .Y(n123) );
  XNOR2X2 U89 ( .A(n117), .B(n25), .Y(DIFF[13]) );
  NAND2BX4 U90 ( .AN(B[10]), .B(n9), .Y(n135) );
  NOR2X4 U91 ( .A(n42), .B(n141), .Y(n140) );
  INVX4 U92 ( .A(n91), .Y(n108) );
  NAND2BX4 U93 ( .AN(B[3]), .B(A[3]), .Y(n66) );
  NAND2BX4 U94 ( .AN(B[12]), .B(A[12]), .Y(n105) );
  NOR3X4 U95 ( .A(n121), .B(n122), .C(n123), .Y(n120) );
  NAND4X2 U96 ( .A(n114), .B(n107), .C(n105), .D(n115), .Y(n112) );
  XOR2X2 U97 ( .A(n53), .B(n54), .Y(DIFF[5]) );
  OAI21X4 U98 ( .A0(n50), .A1(n51), .B0(n52), .Y(n45) );
  INVX4 U99 ( .A(n53), .Y(n50) );
  OAI21X4 U100 ( .A0(n142), .A1(n143), .B0(n144), .Y(n88) );
  NOR2X4 U101 ( .A(n43), .B(n49), .Y(n144) );
  NAND4BX2 U102 ( .AN(n39), .B(n96), .C(n97), .D(n98), .Y(n83) );
  NAND3X4 U103 ( .A(n114), .B(n105), .C(n115), .Y(n117) );
  NAND3X4 U104 ( .A(n125), .B(n93), .C(n126), .Y(n114) );
  NAND3BX4 U105 ( .AN(n119), .B(n19), .C(n120), .Y(n115) );
  XNOR2X4 U106 ( .A(n41), .B(n27), .Y(DIFF[7]) );
  NAND2BX4 U107 ( .AN(A[5]), .B(B[5]), .Y(n151) );
  XOR2X4 U108 ( .A(n127), .B(n4), .Y(DIFF[12]) );
  OAI21X2 U109 ( .A0(n128), .A1(n129), .B0(n84), .Y(n127) );
  OR2X4 U110 ( .A(n118), .B(n110), .Y(n25) );
  INVX4 U111 ( .A(n107), .Y(n118) );
  CLKINVX4 U112 ( .A(n153), .Y(n23) );
  AOI21X4 U113 ( .A0(n117), .A1(n5), .B0(n118), .Y(n116) );
  INVX8 U114 ( .A(n97), .Y(n122) );
  NAND2BX4 U115 ( .AN(B[5]), .B(A[5]), .Y(n52) );
  NAND2BX4 U116 ( .AN(A[3]), .B(B[3]), .Y(n65) );
  NAND2BX4 U117 ( .AN(B[13]), .B(A[13]), .Y(n107) );
  OR2XL U118 ( .A(n42), .B(n43), .Y(n27) );
  NAND2X2 U119 ( .A(n62), .B(n65), .Y(n148) );
  OAI2BB1X4 U120 ( .A0N(n85), .A1N(n58), .B0(n140), .Y(n36) );
  OR2X2 U121 ( .A(n139), .B(n122), .Y(n26) );
  INVX4 U122 ( .A(n146), .Y(n69) );
  NAND2X2 U123 ( .A(n58), .B(n59), .Y(n56) );
  NOR2X2 U124 ( .A(n51), .B(n57), .Y(n142) );
  XNOR2X1 U125 ( .A(n58), .B(n28), .Y(DIFF[4]) );
  NAND2XL U126 ( .A(n57), .B(n59), .Y(n28) );
  OR2XL U127 ( .A(n64), .B(n67), .Y(n29) );
  AOI21XL U128 ( .A0(n62), .A1(n63), .B0(n64), .Y(n61) );
  NOR2XL U129 ( .A(n73), .B(n69), .Y(n72) );
  INVXL U130 ( .A(n70), .Y(n73) );
  OAI21XL U131 ( .A0(n68), .A1(n69), .B0(n70), .Y(n63) );
  NAND2BX2 U132 ( .AN(B[15]), .B(A[15]), .Y(n104) );
  NAND2BX4 U133 ( .AN(B[6]), .B(A[6]), .Y(n46) );
  NAND2XL U134 ( .A(n75), .B(n74), .Y(DIFF[0]) );
  NAND2BXL U135 ( .AN(n75), .B(n74), .Y(n71) );
  INVX1 U136 ( .A(n104), .Y(n103) );
  NOR2XL U137 ( .A(n38), .B(n39), .Y(n37) );
  INVXL U138 ( .A(n40), .Y(n38) );
  NOR2XL U139 ( .A(n48), .B(n49), .Y(n47) );
  INVX1 U140 ( .A(n62), .Y(n67) );
  INVX1 U141 ( .A(n52), .Y(n55) );
  XOR2X1 U142 ( .A(n71), .B(n72), .Y(DIFF[1]) );
  NAND2X1 U143 ( .A(n65), .B(n66), .Y(n60) );
  INVX1 U144 ( .A(n71), .Y(n68) );
  NAND2BX4 U145 ( .AN(n86), .B(n100), .Y(n58) );
  NAND2BX2 U146 ( .AN(A[4]), .B(n21), .Y(n59) );
  NOR2X2 U147 ( .A(n64), .B(n149), .Y(n147) );
  OAI21X2 U148 ( .A0(n69), .A1(n74), .B0(n70), .Y(n149) );
  NAND2BX2 U149 ( .AN(B[11]), .B(A[11]), .Y(n134) );
  NAND2BX1 U150 ( .AN(B[0]), .B(A[0]), .Y(n74) );
  NAND2BX1 U151 ( .AN(A[0]), .B(B[0]), .Y(n75) );
  NOR2XL U152 ( .A(n55), .B(n51), .Y(n54) );
  NAND3XL U153 ( .A(n98), .B(n97), .C(n36), .Y(n129) );
  NAND4BX2 U154 ( .AN(n51), .B(n145), .C(n44), .D(n59), .Y(n99) );
  NAND3X4 U155 ( .A(n77), .B(n78), .C(n79), .Y(n76) );
  NAND2BX4 U156 ( .AN(n80), .B(n81), .Y(n79) );
  NAND4X2 U157 ( .A(n92), .B(n91), .C(n90), .D(n93), .Y(n80) );
  AOI31X2 U158 ( .A0(n105), .A1(n106), .A2(n107), .B0(n108), .Y(n102) );
  NAND2BX4 U159 ( .AN(A[15]), .B(B[15]), .Y(n91) );
  NAND2BX4 U160 ( .AN(B[14]), .B(A[14]), .Y(n106) );
  NAND2BX4 U161 ( .AN(A[14]), .B(B[14]), .Y(n92) );
  NAND2BX4 U162 ( .AN(A[13]), .B(B[13]), .Y(n90) );
  NAND2BX4 U163 ( .AN(A[11]), .B(B[11]), .Y(n98) );
  NAND2BX4 U164 ( .AN(A[10]), .B(B[10]), .Y(n97) );
  NAND2BX4 U165 ( .AN(B[9]), .B(A[9]), .Y(n35) );
  NAND2BX4 U166 ( .AN(B[8]), .B(A[8]), .Y(n40) );
  NAND2BX4 U167 ( .AN(A[8]), .B(B[8]), .Y(n124) );
  OAI21X4 U168 ( .A0(n147), .A1(n148), .B0(n66), .Y(n86) );
  NAND2BX4 U169 ( .AN(A[7]), .B(B[7]), .Y(n145) );
  NAND2BX4 U170 ( .AN(A[6]), .B(B[6]), .Y(n44) );
endmodule


module butterfly_DW01_add_21 ( A, B, SUM );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  wire   n159, n160, n161, n162, n163, n164, n165, n1, n3, n4, n5, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158;

  INVX4 U2 ( .A(n109), .Y(n1) );
  CLKINVX8 U3 ( .A(n11), .Y(n109) );
  OAI21X1 U4 ( .A0(n136), .A1(n137), .B0(n99), .Y(n135) );
  NAND2BX4 U5 ( .AN(n14), .B(n18), .Y(n99) );
  BUFX20 U6 ( .A(n45), .Y(SUM[11]) );
  INVX3 U7 ( .A(n62), .Y(n61) );
  INVX4 U8 ( .A(n134), .Y(n132) );
  NAND2X2 U9 ( .A(n142), .B(n144), .Y(n26) );
  CLKBUFX3 U10 ( .A(n54), .Y(n3) );
  CLKINVX4 U11 ( .A(n60), .Y(n153) );
  CLKINVX2 U12 ( .A(n53), .Y(n10) );
  OR2X2 U13 ( .A(A[12]), .B(B[12]), .Y(n107) );
  AOI21X2 U14 ( .A0(n32), .A1(n31), .B0(n101), .Y(n97) );
  NOR2X2 U15 ( .A(n12), .B(n112), .Y(n122) );
  OAI21X2 U16 ( .A0(n112), .A1(n117), .B0(n125), .Y(n124) );
  NAND2X2 U17 ( .A(B[2]), .B(A[2]), .Y(n82) );
  OR2X4 U18 ( .A(A[2]), .B(B[2]), .Y(n85) );
  XOR2X4 U19 ( .A(n74), .B(n75), .Y(SUM[4]) );
  BUFX20 U20 ( .A(n163), .Y(SUM[6]) );
  XOR2X4 U21 ( .A(n65), .B(n66), .Y(n163) );
  BUFX20 U22 ( .A(n162), .Y(SUM[7]) );
  NAND2X4 U23 ( .A(n42), .B(n43), .Y(n162) );
  NAND3X2 U24 ( .A(n20), .B(n67), .C(n152), .Y(n150) );
  NAND2X2 U25 ( .A(B[0]), .B(A[0]), .Y(n91) );
  INVXL U26 ( .A(n70), .Y(n25) );
  CLKINVX3 U27 ( .A(n69), .Y(n20) );
  OAI21X2 U28 ( .A0(n90), .A1(n91), .B0(n88), .Y(n158) );
  CLKINVX3 U29 ( .A(n154), .Y(n31) );
  CLKINVX3 U30 ( .A(n142), .Y(n141) );
  NAND2X2 U31 ( .A(n52), .B(n56), .Y(n139) );
  INVX1 U32 ( .A(n117), .Y(n127) );
  OR2X2 U33 ( .A(A[3]), .B(B[3]), .Y(n155) );
  OAI21X2 U34 ( .A0(n46), .A1(n154), .B0(n73), .Y(n71) );
  BUFX12 U35 ( .A(n159), .Y(SUM[15]) );
  OR2X2 U36 ( .A(n29), .B(n30), .Y(n58) );
  NOR2X1 U37 ( .A(n24), .B(n63), .Y(n29) );
  NOR2BX1 U38 ( .AN(n88), .B(n90), .Y(n89) );
  INVX1 U39 ( .A(n24), .Y(n65) );
  NOR2BX1 U40 ( .AN(n56), .B(n57), .Y(n55) );
  XOR2X1 U41 ( .A(n22), .B(n51), .Y(n161) );
  INVX1 U42 ( .A(n146), .Y(n39) );
  NAND2X1 U43 ( .A(n58), .B(n41), .Y(n42) );
  NAND2X2 U44 ( .A(n40), .B(n59), .Y(n43) );
  INVX1 U45 ( .A(n59), .Y(n41) );
  INVX4 U46 ( .A(B[11]), .Y(n4) );
  INVX4 U47 ( .A(n4), .Y(n5) );
  INVX4 U48 ( .A(n61), .Y(n27) );
  BUFX3 U49 ( .A(n164), .Y(SUM[5]) );
  AND2X2 U50 ( .A(n120), .B(n9), .Y(n7) );
  INVX1 U51 ( .A(n154), .Y(n74) );
  CLKINVX3 U52 ( .A(n100), .Y(n154) );
  NAND2X1 U53 ( .A(n110), .B(n143), .Y(n8) );
  NOR2BX1 U54 ( .AN(n117), .B(n12), .Y(n128) );
  NOR2X2 U55 ( .A(n12), .B(n120), .Y(n119) );
  CLKINVX3 U56 ( .A(n12), .Y(n104) );
  NOR2BX1 U57 ( .AN(n70), .B(n69), .Y(n72) );
  NOR3BX2 U58 ( .AN(n107), .B(n1), .C(n14), .Y(n131) );
  INVXL U59 ( .A(n147), .Y(n22) );
  NAND2X2 U60 ( .A(B[9]), .B(A[9]), .Y(n52) );
  NAND2X4 U61 ( .A(B[10]), .B(A[10]), .Y(n142) );
  OR2X4 U62 ( .A(A[12]), .B(B[12]), .Y(n9) );
  NAND2X2 U63 ( .A(B[12]), .B(A[12]), .Y(n120) );
  CLKINVX8 U64 ( .A(n106), .Y(n112) );
  BUFX2 U65 ( .A(B[14]), .Y(n21) );
  NOR2X4 U66 ( .A(A[10]), .B(B[10]), .Y(n11) );
  NOR2X4 U67 ( .A(A[13]), .B(B[13]), .Y(n12) );
  NAND3X2 U68 ( .A(n13), .B(n54), .C(n131), .Y(n130) );
  AND2X1 U69 ( .A(n111), .B(n108), .Y(n13) );
  OAI2BB1X1 U70 ( .A0N(n139), .A1N(n138), .B0(n140), .Y(n18) );
  NOR2X2 U71 ( .A(B[11]), .B(A[11]), .Y(n14) );
  NAND2X1 U72 ( .A(n109), .B(n145), .Y(n144) );
  NAND2X4 U73 ( .A(n93), .B(n94), .Y(n92) );
  BUFX20 U74 ( .A(n160), .Y(SUM[14]) );
  NAND3XL U75 ( .A(n110), .B(n109), .C(n54), .Y(n137) );
  INVX4 U76 ( .A(n111), .Y(n57) );
  XNOR2X4 U77 ( .A(n121), .B(n15), .Y(n159) );
  AND2X2 U78 ( .A(n115), .B(n105), .Y(n15) );
  XOR2X2 U79 ( .A(n123), .B(n128), .Y(SUM[13]) );
  NAND2X4 U80 ( .A(n28), .B(n99), .Y(n96) );
  AOI2BB1X4 U81 ( .A0N(n68), .A1N(n69), .B0(n25), .Y(n24) );
  XNOR2X4 U82 ( .A(n126), .B(n16), .Y(n160) );
  AND2X1 U83 ( .A(n106), .B(n125), .Y(n16) );
  NOR2BX4 U84 ( .AN(n17), .B(n127), .Y(n126) );
  NAND2X4 U85 ( .A(n123), .B(n104), .Y(n17) );
  AOI21X4 U86 ( .A0(n5), .A1(A[11]), .B0(n141), .Y(n140) );
  INVXL U87 ( .A(n102), .Y(n101) );
  CLKBUFX2 U88 ( .A(n64), .Y(n19) );
  INVX2 U89 ( .A(n115), .Y(n114) );
  NOR2X4 U90 ( .A(n113), .B(n114), .Y(n93) );
  INVX8 U91 ( .A(n151), .Y(n69) );
  NAND4X2 U92 ( .A(n104), .B(n105), .C(n106), .D(n9), .Y(n95) );
  AOI21X4 U93 ( .A0(n116), .A1(n117), .B0(n118), .Y(n113) );
  NAND2X1 U94 ( .A(B[14]), .B(A[14]), .Y(n125) );
  INVX8 U95 ( .A(n50), .Y(n147) );
  BUFX4 U96 ( .A(A[1]), .Y(n23) );
  NAND4BX2 U97 ( .AN(n57), .B(n10), .C(n109), .D(n110), .Y(n98) );
  XNOR2X4 U98 ( .A(n26), .B(n8), .Y(n45) );
  NAND2X4 U99 ( .A(n148), .B(n56), .Y(n50) );
  NOR2BX4 U100 ( .AN(n82), .B(n158), .Y(n156) );
  NOR2BX4 U101 ( .AN(n64), .B(n153), .Y(n149) );
  NAND2X2 U102 ( .A(B[5]), .B(A[5]), .Y(n70) );
  AOI21X4 U103 ( .A0(A[14]), .A1(n21), .B0(n119), .Y(n116) );
  NOR2BX1 U104 ( .AN(n73), .B(n46), .Y(n75) );
  NAND2X4 U105 ( .A(n70), .B(n73), .Y(n152) );
  NAND2X2 U106 ( .A(B[6]), .B(A[6]), .Y(n64) );
  INVX8 U107 ( .A(n108), .Y(n53) );
  INVX1 U108 ( .A(n67), .Y(n63) );
  NAND2X2 U109 ( .A(B[7]), .B(A[7]), .Y(n60) );
  NAND2X2 U110 ( .A(B[1]), .B(n23), .Y(n88) );
  NAND2X2 U111 ( .A(n9), .B(n110), .Y(n133) );
  OAI2BB1X2 U112 ( .A0N(n86), .A1N(n87), .B0(n88), .Y(n83) );
  NAND2BX4 U113 ( .AN(n95), .B(n96), .Y(n94) );
  NOR2X4 U114 ( .A(A[4]), .B(B[4]), .Y(n46) );
  NOR2X4 U115 ( .A(n53), .B(n11), .Y(n138) );
  NAND2X4 U116 ( .A(B[13]), .B(A[13]), .Y(n117) );
  OAI21X4 U117 ( .A0(n132), .A1(n133), .B0(n120), .Y(n129) );
  INVX8 U118 ( .A(n38), .Y(SUM[10]) );
  XOR2X4 U119 ( .A(n145), .B(n39), .Y(n38) );
  OR2X4 U120 ( .A(n97), .B(n98), .Y(n28) );
  XOR2X2 U121 ( .A(n3), .B(n55), .Y(SUM[8]) );
  NAND2X4 U122 ( .A(B[8]), .B(A[8]), .Y(n56) );
  INVXL U123 ( .A(n19), .Y(n30) );
  INVX4 U124 ( .A(n58), .Y(n40) );
  OR2X4 U125 ( .A(B[7]), .B(A[7]), .Y(n62) );
  NAND2X4 U126 ( .A(n32), .B(n31), .Y(n33) );
  NAND2X4 U127 ( .A(n33), .B(n102), .Y(n54) );
  CLKINVX8 U128 ( .A(n103), .Y(n32) );
  NAND4BBX4 U129 ( .AN(n69), .BN(n46), .C(n62), .D(n67), .Y(n103) );
  BUFX3 U130 ( .A(n165), .Y(SUM[0]) );
  BUFX4 U131 ( .A(n161), .Y(SUM[9]) );
  NAND2X4 U132 ( .A(B[4]), .B(A[4]), .Y(n73) );
  XOR2X4 U133 ( .A(n135), .B(n7), .Y(SUM[12]) );
  XOR2X1 U134 ( .A(n76), .B(n77), .Y(SUM[3]) );
  OAI21XL U135 ( .A0(n80), .A1(n81), .B0(n82), .Y(n76) );
  NOR2BX1 U136 ( .AN(n78), .B(n79), .Y(n77) );
  INVXL U137 ( .A(n83), .Y(n80) );
  NAND2X2 U138 ( .A(n106), .B(n105), .Y(n118) );
  NOR2XL U139 ( .A(A[0]), .B(B[0]), .Y(n44) );
  NAND2X4 U140 ( .A(n54), .B(n111), .Y(n148) );
  OAI21X4 U141 ( .A0(n147), .A1(n53), .B0(n52), .Y(n145) );
  INVX2 U142 ( .A(n71), .Y(n68) );
  INVX4 U143 ( .A(n86), .Y(n90) );
  NAND2X1 U144 ( .A(B[3]), .B(A[3]), .Y(n78) );
  NAND2XL U145 ( .A(B[15]), .B(A[15]), .Y(n115) );
  INVXL U146 ( .A(n91), .Y(n87) );
  NOR2BX1 U147 ( .AN(n91), .B(n44), .Y(n165) );
  AOI21X2 U148 ( .A0(n123), .A1(n122), .B0(n124), .Y(n121) );
  NOR2BX1 U149 ( .AN(n19), .B(n63), .Y(n66) );
  XOR2X1 U150 ( .A(n71), .B(n72), .Y(n164) );
  NOR2BX1 U151 ( .AN(n60), .B(n61), .Y(n59) );
  XOR2X1 U152 ( .A(n83), .B(n84), .Y(SUM[2]) );
  NOR2BX1 U153 ( .AN(n82), .B(n81), .Y(n84) );
  INVX1 U154 ( .A(n85), .Y(n81) );
  XOR2X1 U155 ( .A(n87), .B(n89), .Y(SUM[1]) );
  INVXL U156 ( .A(n155), .Y(n79) );
  XNOR3X4 U157 ( .A(B[16]), .B(A[16]), .C(n92), .Y(n47) );
  INVX8 U158 ( .A(n47), .Y(SUM[16]) );
  NOR2BXL U159 ( .AN(n142), .B(n11), .Y(n146) );
  NAND2XL U160 ( .A(A[11]), .B(n5), .Y(n143) );
  NAND2XL U161 ( .A(n111), .B(n10), .Y(n136) );
  NOR2BXL U162 ( .AN(n52), .B(n53), .Y(n51) );
  OR2X4 U163 ( .A(A[15]), .B(B[15]), .Y(n105) );
  OR2X4 U164 ( .A(B[14]), .B(A[14]), .Y(n106) );
  NAND2BX4 U165 ( .AN(n129), .B(n130), .Y(n123) );
  OAI2BB1X4 U166 ( .A0N(n139), .A1N(n138), .B0(n140), .Y(n134) );
  OR2X4 U167 ( .A(B[11]), .B(A[11]), .Y(n110) );
  OR2X4 U168 ( .A(A[9]), .B(B[9]), .Y(n108) );
  OR2X4 U169 ( .A(A[8]), .B(B[8]), .Y(n111) );
  OAI2BB1X4 U170 ( .A0N(n149), .A1N(n150), .B0(n27), .Y(n102) );
  OR2X4 U171 ( .A(B[6]), .B(A[6]), .Y(n67) );
  OR2X4 U172 ( .A(B[5]), .B(A[5]), .Y(n151) );
  OAI21X4 U173 ( .A0(n156), .A1(n157), .B0(n78), .Y(n100) );
  NAND2X4 U174 ( .A(n85), .B(n155), .Y(n157) );
  OR2X4 U175 ( .A(A[1]), .B(B[1]), .Y(n86) );
endmodule


module butterfly_DW01_sub_36 ( A, B, DIFF );
  input [16:0] A;
  input [16:0] B;
  output [16:0] DIFF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191;

  CLKINVX3 U3 ( .A(n103), .Y(n86) );
  AOI21X1 U4 ( .A0(n88), .A1(n87), .B0(n86), .Y(n120) );
  CLKINVX3 U5 ( .A(n132), .Y(n114) );
  BUFX4 U6 ( .A(n109), .Y(n12) );
  NAND2BX4 U7 ( .AN(B[13]), .B(A[13]), .Y(n87) );
  INVX4 U8 ( .A(n123), .Y(n89) );
  NOR2X1 U9 ( .A(n80), .B(n81), .Y(n76) );
  AND3X2 U10 ( .A(n73), .B(n74), .C(n75), .Y(n72) );
  INVX4 U11 ( .A(n191), .Y(n54) );
  INVX4 U12 ( .A(n95), .Y(n22) );
  AOI21X4 U13 ( .A0(n153), .A1(B[10]), .B0(n154), .Y(n151) );
  CLKINVX3 U14 ( .A(n113), .Y(n119) );
  NAND2X2 U15 ( .A(n123), .B(n103), .Y(n113) );
  AOI21X4 U16 ( .A0(n151), .A1(n140), .B0(n152), .Y(n150) );
  NAND3X2 U17 ( .A(n161), .B(n174), .C(n38), .Y(n183) );
  NOR2X2 U18 ( .A(n89), .B(n90), .Y(n1) );
  INVX4 U19 ( .A(n87), .Y(n2) );
  OR2X4 U20 ( .A(n1), .B(n2), .Y(n129) );
  NAND2BX4 U21 ( .AN(n129), .B(n130), .Y(n128) );
  AOI21X1 U22 ( .A0(n21), .A1(n142), .B0(n168), .Y(n167) );
  INVX3 U23 ( .A(n144), .Y(n168) );
  NAND2BX4 U24 ( .AN(A[10]), .B(B[10]), .Y(n142) );
  XOR2X2 U25 ( .A(n40), .B(n48), .Y(DIFF[4]) );
  XNOR2X2 U26 ( .A(B[16]), .B(A[16]), .Y(n69) );
  NAND2BX4 U27 ( .AN(A[14]), .B(B[14]), .Y(n103) );
  XNOR2X4 U28 ( .A(n148), .B(n17), .Y(DIFF[12]) );
  AOI21X2 U29 ( .A0(n119), .A1(n137), .B0(n120), .Y(n118) );
  INVX2 U30 ( .A(n143), .Y(n164) );
  NAND2X2 U31 ( .A(n155), .B(n156), .Y(n141) );
  NAND2BX1 U32 ( .AN(A[9]), .B(B[9]), .Y(n140) );
  CLKINVX3 U33 ( .A(n141), .Y(n154) );
  CLKINVX3 U34 ( .A(n142), .Y(n115) );
  NAND2BX1 U35 ( .AN(A[7]), .B(B[7]), .Y(n159) );
  INVX1 U36 ( .A(A[5]), .Y(n8) );
  NAND3X1 U37 ( .A(n121), .B(n122), .C(n119), .Y(n117) );
  CLKINVX3 U38 ( .A(n74), .Y(n106) );
  NAND2BX2 U39 ( .AN(B[14]), .B(A[14]), .Y(n88) );
  CLKINVX3 U40 ( .A(n155), .Y(n21) );
  NOR3BX2 U41 ( .AN(n35), .B(n162), .C(n24), .Y(n169) );
  AND2X2 U42 ( .A(n123), .B(n87), .Y(n18) );
  OAI21XL U43 ( .A0(n91), .A1(n79), .B0(n92), .Y(n71) );
  NAND2BX1 U44 ( .AN(A[7]), .B(B[7]), .Y(n35) );
  NAND2BX1 U45 ( .AN(A[0]), .B(B[0]), .Y(n67) );
  NOR2X1 U46 ( .A(n49), .B(n47), .Y(n48) );
  INVX2 U47 ( .A(n90), .Y(n137) );
  NOR2X4 U48 ( .A(n116), .B(n124), .Y(n121) );
  CLKINVX3 U49 ( .A(n38), .Y(n34) );
  INVX1 U50 ( .A(n43), .Y(n47) );
  NAND2BX1 U51 ( .AN(A[11]), .B(B[11]), .Y(n145) );
  CLKINVX3 U52 ( .A(n145), .Y(n124) );
  NAND3X1 U53 ( .A(n146), .B(n147), .C(n109), .Y(n135) );
  NAND2X2 U54 ( .A(n135), .B(n136), .Y(n134) );
  NOR2X1 U55 ( .A(n115), .B(n116), .Y(n147) );
  NAND2X4 U56 ( .A(n55), .B(n52), .Y(n188) );
  XNOR2X4 U57 ( .A(n3), .B(n176), .Y(DIFF[10]) );
  AND3X4 U58 ( .A(n177), .B(n178), .C(n179), .Y(n3) );
  NAND2X2 U59 ( .A(n61), .B(n66), .Y(n190) );
  NAND2BX1 U60 ( .AN(A[11]), .B(B[11]), .Y(n132) );
  NOR2X1 U61 ( .A(n112), .B(n113), .Y(n111) );
  NOR2X2 U62 ( .A(n114), .B(n112), .Y(n146) );
  NOR3X2 U63 ( .A(n124), .B(n89), .C(n116), .Y(n131) );
  NAND2BX2 U64 ( .AN(B[3]), .B(A[3]), .Y(n56) );
  XNOR2X4 U65 ( .A(n163), .B(n4), .Y(DIFF[11]) );
  OR2X2 U66 ( .A(n164), .B(n165), .Y(n4) );
  NAND2X4 U67 ( .A(n54), .B(n55), .Y(n100) );
  NAND2X1 U68 ( .A(n95), .B(n94), .Y(n112) );
  BUFX3 U69 ( .A(n27), .Y(n5) );
  NAND4BX2 U70 ( .AN(n158), .B(n38), .C(n159), .D(n40), .Y(n27) );
  NAND4BX4 U71 ( .AN(n34), .B(n6), .C(n175), .D(n174), .Y(n170) );
  AND2X2 U72 ( .A(n94), .B(n161), .Y(n6) );
  NAND4BX2 U73 ( .AN(n173), .B(n7), .C(n174), .D(n40), .Y(n171) );
  AND2X2 U74 ( .A(n38), .B(n39), .Y(n7) );
  NAND2BX2 U75 ( .AN(B[6]), .B(A[6]), .Y(n162) );
  NAND2BX2 U76 ( .AN(B[10]), .B(A[10]), .Y(n144) );
  AOI21X4 U77 ( .A0(n180), .A1(n181), .B0(n21), .Y(n179) );
  NOR3X4 U78 ( .A(n22), .B(n24), .C(n184), .Y(n180) );
  NAND4X2 U79 ( .A(n52), .B(n65), .C(n55), .D(n67), .Y(n81) );
  INVX12 U80 ( .A(n156), .Y(n25) );
  OAI2BB1X2 U81 ( .A0N(n8), .A1N(B[5]), .B0(n39), .Y(n158) );
  NAND2X4 U82 ( .A(n30), .B(n35), .Y(n97) );
  INVX3 U83 ( .A(n174), .Y(n42) );
  NAND2X1 U84 ( .A(n32), .B(n33), .Y(n37) );
  AOI21X4 U85 ( .A0(n157), .A1(n9), .B0(n25), .Y(n172) );
  NAND2X2 U86 ( .A(n117), .B(n118), .Y(n107) );
  NAND2X1 U87 ( .A(n38), .B(n94), .Y(n185) );
  NOR2X2 U88 ( .A(n24), .B(n25), .Y(n15) );
  NAND3X2 U89 ( .A(n12), .B(n110), .C(n111), .Y(n108) );
  AOI21X4 U90 ( .A0(n127), .A1(n12), .B0(n128), .Y(n126) );
  NOR3BX2 U91 ( .AN(n132), .B(n133), .C(n112), .Y(n127) );
  NOR2X4 U92 ( .A(n11), .B(n34), .Y(n31) );
  NAND2X1 U93 ( .A(n39), .B(n40), .Y(n10) );
  NAND4X4 U94 ( .A(n174), .B(n160), .C(n38), .D(n161), .Y(n98) );
  NAND2BX1 U95 ( .AN(A[7]), .B(B[7]), .Y(n160) );
  NAND2BX4 U96 ( .AN(n107), .B(n108), .Y(n105) );
  AND4X2 U97 ( .A(n95), .B(n9), .C(n142), .D(n96), .Y(n149) );
  INVX2 U98 ( .A(n80), .Y(n70) );
  NAND4BX2 U99 ( .AN(n89), .B(n102), .C(n103), .D(n104), .Y(n80) );
  NAND2X2 U100 ( .A(n143), .B(n144), .Y(n152) );
  NAND2X2 U101 ( .A(n143), .B(n144), .Y(n138) );
  INVX8 U102 ( .A(n102), .Y(n116) );
  NAND3BX1 U103 ( .AN(n185), .B(n40), .C(n186), .Y(n177) );
  NAND2BX4 U104 ( .AN(B[1]), .B(A[1]), .Y(n61) );
  NAND4BX4 U105 ( .AN(n169), .B(n170), .C(n171), .D(n172), .Y(n20) );
  NAND2BX4 U106 ( .AN(B[5]), .B(A[5]), .Y(n44) );
  NAND2BX2 U107 ( .AN(A[1]), .B(B[1]), .Y(n65) );
  NAND2BXL U108 ( .AN(A[1]), .B(B[1]), .Y(n189) );
  NAND2BX2 U109 ( .AN(B[15]), .B(A[15]), .Y(n74) );
  NAND2BX2 U110 ( .AN(n26), .B(n5), .Y(n23) );
  INVX2 U111 ( .A(n159), .Y(n187) );
  NOR2X2 U112 ( .A(n115), .B(n168), .Y(n176) );
  NAND2XL U113 ( .A(n35), .B(n36), .Y(n28) );
  NAND3X4 U114 ( .A(n97), .B(n36), .C(n98), .Y(n26) );
  NAND4BX4 U115 ( .AN(n157), .B(n97), .C(n98), .D(n27), .Y(n109) );
  INVX2 U116 ( .A(n61), .Y(n64) );
  OAI21X2 U117 ( .A0(n59), .A1(n60), .B0(n61), .Y(n53) );
  NAND2BX1 U118 ( .AN(A[7]), .B(B[7]), .Y(n99) );
  NAND2BX4 U119 ( .AN(B[8]), .B(A[8]), .Y(n156) );
  OR2X4 U120 ( .A(n21), .B(n22), .Y(n13) );
  INVX8 U121 ( .A(n24), .Y(n9) );
  INVX4 U122 ( .A(n36), .Y(n157) );
  NAND2X2 U123 ( .A(n36), .B(n162), .Y(n182) );
  NAND2BX4 U124 ( .AN(B[7]), .B(A[7]), .Y(n36) );
  NAND4XL U125 ( .A(n96), .B(n9), .C(n142), .D(n95), .Y(n79) );
  INVX8 U126 ( .A(n94), .Y(n24) );
  XNOR2X4 U127 ( .A(n105), .B(n16), .Y(DIFF[15]) );
  XOR2X4 U128 ( .A(n68), .B(n69), .Y(DIFF[16]) );
  NAND2BX4 U129 ( .AN(A[2]), .B(B[2]), .Y(n52) );
  INVX2 U130 ( .A(n52), .Y(n58) );
  NAND3X2 U131 ( .A(n174), .B(n39), .C(n40), .Y(n33) );
  INVX4 U132 ( .A(n41), .Y(n32) );
  OAI21X4 U133 ( .A0(n42), .A1(n43), .B0(n44), .Y(n41) );
  NAND4X4 U134 ( .A(n100), .B(n81), .C(n101), .D(n56), .Y(n40) );
  NAND2BX4 U135 ( .AN(A[13]), .B(B[13]), .Y(n123) );
  NAND2BX4 U136 ( .AN(B[11]), .B(A[11]), .Y(n143) );
  NOR3BX2 U137 ( .AN(n95), .B(n158), .C(n187), .Y(n186) );
  NAND2BX4 U138 ( .AN(B[4]), .B(A[4]), .Y(n43) );
  NAND2X2 U139 ( .A(n94), .B(n99), .Y(n173) );
  NAND3X2 U140 ( .A(n140), .B(n141), .C(n142), .Y(n139) );
  NOR2X4 U141 ( .A(n30), .B(n31), .Y(n29) );
  NAND2BX2 U142 ( .AN(A[15]), .B(B[15]), .Y(n104) );
  OAI2BB1X4 U143 ( .A0N(n166), .A1N(n20), .B0(n167), .Y(n163) );
  NAND2BX4 U144 ( .AN(B[12]), .B(A[12]), .Y(n90) );
  INVX4 U145 ( .A(n162), .Y(n30) );
  AND2X4 U146 ( .A(n10), .B(n43), .Y(n46) );
  NAND2BX4 U147 ( .AN(A[4]), .B(B[4]), .Y(n39) );
  XOR2X4 U148 ( .A(n45), .B(n46), .Y(DIFF[5]) );
  AND2X4 U149 ( .A(n32), .B(n33), .Y(n11) );
  NOR2X1 U150 ( .A(n64), .B(n60), .Y(n63) );
  NOR3X1 U151 ( .A(n114), .B(n115), .C(n116), .Y(n110) );
  XNOR2X4 U152 ( .A(n20), .B(n13), .Y(DIFF[9]) );
  XNOR2X4 U153 ( .A(n37), .B(n14), .Y(DIFF[6]) );
  OR2X4 U154 ( .A(n30), .B(n34), .Y(n14) );
  XOR2X4 U155 ( .A(n23), .B(n15), .Y(DIFF[8]) );
  INVX2 U156 ( .A(n62), .Y(n59) );
  NOR2X1 U157 ( .A(n85), .B(n86), .Y(n84) );
  XOR2X1 U158 ( .A(n50), .B(n51), .Y(DIFF[3]) );
  AOI21X1 U159 ( .A0(n52), .A1(n53), .B0(n54), .Y(n51) );
  OR2X4 U160 ( .A(n85), .B(n106), .Y(n16) );
  XOR2X1 U161 ( .A(n62), .B(n63), .Y(DIFF[1]) );
  AND2X1 U162 ( .A(n102), .B(n90), .Y(n17) );
  NAND2BXL U163 ( .AN(A[11]), .B(B[11]), .Y(n96) );
  NAND2BXL U164 ( .AN(B[0]), .B(A[0]), .Y(n66) );
  INVXL U165 ( .A(A[10]), .Y(n153) );
  NOR2X1 U166 ( .A(n115), .B(n22), .Y(n166) );
  INVXL U167 ( .A(n93), .Y(n92) );
  NAND2X1 U168 ( .A(n76), .B(n77), .Y(n75) );
  NOR2X1 U169 ( .A(n78), .B(n79), .Y(n77) );
  NAND2XL U170 ( .A(n174), .B(n44), .Y(n45) );
  NAND2XL U171 ( .A(n25), .B(n95), .Y(n178) );
  NAND2XL U172 ( .A(n103), .B(n88), .Y(n125) );
  NAND2BX2 U173 ( .AN(n182), .B(n183), .Y(n181) );
  AOI21X2 U174 ( .A0(n121), .A1(n122), .B0(n137), .Y(n136) );
  NAND2X2 U175 ( .A(n131), .B(n122), .Y(n130) );
  INVXL U176 ( .A(n39), .Y(n49) );
  NAND4XL U177 ( .A(n99), .B(n39), .C(n174), .D(n38), .Y(n78) );
  NAND2X1 U178 ( .A(n66), .B(n67), .Y(DIFF[0]) );
  INVX1 U179 ( .A(n65), .Y(n60) );
  INVX1 U180 ( .A(n104), .Y(n85) );
  AOI2BB1XL U181 ( .A0N(n19), .A1N(n78), .B0(n26), .Y(n91) );
  AND3X1 U182 ( .A(n56), .B(n100), .C(n101), .Y(n19) );
  XOR2X2 U183 ( .A(n53), .B(n57), .Y(DIFF[2]) );
  NOR2XL U184 ( .A(n54), .B(n58), .Y(n57) );
  NAND2XL U185 ( .A(n55), .B(n56), .Y(n50) );
  NAND3XL U186 ( .A(n102), .B(n123), .C(n142), .Y(n133) );
  NAND2BX1 U187 ( .AN(n67), .B(n66), .Y(n62) );
  OAI21X1 U188 ( .A0(n82), .A1(n83), .B0(n84), .Y(n73) );
  NAND2X1 U189 ( .A(n87), .B(n88), .Y(n83) );
  NOR2XL U190 ( .A(n89), .B(n90), .Y(n82) );
  OAI2BB1X2 U191 ( .A0N(n70), .A1N(n71), .B0(n72), .Y(n68) );
  NOR2BX1 U192 ( .AN(B[11]), .B(A[11]), .Y(n165) );
  NAND2BX4 U193 ( .AN(A[5]), .B(B[5]), .Y(n174) );
  NAND2BXL U194 ( .AN(A[7]), .B(B[7]), .Y(n175) );
  NOR2BX1 U195 ( .AN(B[7]), .B(A[7]), .Y(n184) );
  NAND2BX1 U196 ( .AN(B[2]), .B(A[2]), .Y(n191) );
  XOR2X4 U197 ( .A(n28), .B(n29), .Y(DIFF[7]) );
  XOR2X4 U198 ( .A(n125), .B(n126), .Y(DIFF[14]) );
  XOR2X4 U199 ( .A(n134), .B(n18), .Y(DIFF[13]) );
  NAND2BX4 U200 ( .AN(n138), .B(n139), .Y(n122) );
  AOI21X4 U201 ( .A0(n149), .A1(n109), .B0(n93), .Y(n148) );
  NOR2X4 U202 ( .A(n150), .B(n124), .Y(n93) );
  NAND2BX4 U203 ( .AN(A[12]), .B(B[12]), .Y(n102) );
  NAND2BX4 U204 ( .AN(B[9]), .B(A[9]), .Y(n155) );
  NAND2X4 U205 ( .A(n44), .B(n43), .Y(n161) );
  NAND2BX4 U206 ( .AN(A[9]), .B(B[9]), .Y(n95) );
  NAND3BX4 U207 ( .AN(n188), .B(n189), .C(n190), .Y(n101) );
  NAND2BX4 U208 ( .AN(A[3]), .B(B[3]), .Y(n55) );
  NAND2BX4 U209 ( .AN(A[8]), .B(B[8]), .Y(n94) );
  NAND2BX4 U210 ( .AN(A[6]), .B(B[6]), .Y(n38) );
endmodule


module butterfly_DW01_add_43 ( A, B, SUM );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177;

  AND2X4 U2 ( .A(n34), .B(n148), .Y(n26) );
  OAI21X2 U3 ( .A0(n113), .A1(n98), .B0(n99), .Y(n109) );
  CLKINVX3 U4 ( .A(n36), .Y(n166) );
  NAND2X2 U5 ( .A(n158), .B(n133), .Y(n155) );
  INVXL U6 ( .A(n139), .Y(n1) );
  INVX8 U7 ( .A(n44), .Y(n139) );
  NAND2X2 U8 ( .A(n148), .B(n51), .Y(n163) );
  NAND3BX4 U9 ( .AN(n166), .B(n170), .C(n35), .Y(n169) );
  OAI21X2 U10 ( .A0(n175), .A1(n176), .B0(n164), .Y(n170) );
  OAI21X4 U11 ( .A0(n55), .A1(n19), .B0(n20), .Y(n52) );
  INVX4 U12 ( .A(n6), .Y(n43) );
  INVX8 U13 ( .A(n101), .Y(n140) );
  NOR2BX1 U14 ( .AN(n73), .B(n29), .Y(n75) );
  NOR2BX2 U15 ( .AN(n98), .B(n96), .Y(n129) );
  INVX4 U16 ( .A(n114), .Y(n96) );
  NOR2BX2 U17 ( .AN(n99), .B(n113), .Y(n120) );
  NAND2X2 U18 ( .A(B[0]), .B(A[0]), .Y(n81) );
  NAND2BX2 U19 ( .AN(n38), .B(n39), .Y(n37) );
  INVX1 U20 ( .A(n33), .Y(n167) );
  OR2X2 U21 ( .A(A[3]), .B(B[3]), .Y(n71) );
  NOR2X2 U22 ( .A(n52), .B(n53), .Y(n49) );
  INVX1 U23 ( .A(n54), .Y(n53) );
  AND2X2 U24 ( .A(B[7]), .B(A[7]), .Y(n6) );
  CLKINVX3 U25 ( .A(n92), .Y(n113) );
  OAI2BB1X1 U26 ( .A0N(n76), .A1N(n77), .B0(n78), .Y(n74) );
  INVX4 U27 ( .A(n148), .Y(n42) );
  INVX1 U28 ( .A(n136), .Y(n157) );
  OAI21X1 U29 ( .A0(n89), .A1(n90), .B0(n91), .Y(n88) );
  NOR2X1 U30 ( .A(n94), .B(n95), .Y(n89) );
  OAI21XL U31 ( .A0(n105), .A1(n100), .B0(n106), .Y(n102) );
  INVX1 U32 ( .A(n107), .Y(n87) );
  XOR2X1 U33 ( .A(n77), .B(n79), .Y(SUM[1]) );
  NAND2X1 U34 ( .A(n23), .B(n64), .Y(n14) );
  BUFX8 U35 ( .A(n24), .Y(n2) );
  BUFX8 U36 ( .A(n24), .Y(n3) );
  AND2X2 U37 ( .A(n91), .B(n93), .Y(n4) );
  AND2X1 U38 ( .A(n138), .B(n133), .Y(n5) );
  INVX1 U39 ( .A(n47), .Y(n46) );
  XOR2X4 U40 ( .A(n7), .B(n8), .Y(SUM[7]) );
  OR2X4 U41 ( .A(n45), .B(n46), .Y(n7) );
  AND2X1 U42 ( .A(n43), .B(n44), .Y(n8) );
  NAND4X4 U43 ( .A(n92), .B(n116), .C(n115), .D(n114), .Y(n112) );
  NAND2XL U44 ( .A(n92), .B(n93), .Y(n90) );
  INVX8 U45 ( .A(n116), .Y(n121) );
  OR2X2 U46 ( .A(A[11]), .B(B[11]), .Y(n27) );
  NAND3X2 U47 ( .A(A[5]), .B(B[5]), .C(n3), .Y(n165) );
  NAND2X4 U48 ( .A(n9), .B(n10), .Y(n16) );
  OR3X4 U49 ( .A(n150), .B(n151), .C(n20), .Y(n9) );
  AND3X4 U50 ( .A(n47), .B(n165), .C(n43), .Y(n10) );
  BUFX12 U51 ( .A(n57), .Y(n20) );
  INVX8 U52 ( .A(n51), .Y(n151) );
  NAND3BX4 U53 ( .AN(n11), .B(n161), .C(n162), .Y(n159) );
  OR2X2 U54 ( .A(n166), .B(n167), .Y(n11) );
  OAI2BB1X2 U55 ( .A0N(n145), .A1N(n135), .B0(n136), .Y(n104) );
  NAND3X1 U56 ( .A(n28), .B(n138), .C(n26), .Y(n107) );
  NAND4BX2 U57 ( .AN(n163), .B(n12), .C(n22), .D(n63), .Y(n162) );
  AND2X2 U58 ( .A(n44), .B(n3), .Y(n12) );
  NAND2X2 U59 ( .A(A[10]), .B(B[10]), .Y(n133) );
  NAND2X2 U60 ( .A(n101), .B(n136), .Y(n117) );
  NAND2XL U61 ( .A(n47), .B(n3), .Y(n62) );
  OAI21X2 U62 ( .A0(n72), .A1(n29), .B0(n73), .Y(n68) );
  INVX4 U63 ( .A(n74), .Y(n72) );
  NOR2X1 U64 ( .A(A[2]), .B(B[2]), .Y(n29) );
  INVX8 U65 ( .A(n63), .Y(n55) );
  NAND2X2 U66 ( .A(n58), .B(n59), .Y(n48) );
  NOR2BX2 U67 ( .AN(n114), .B(n117), .Y(n125) );
  NAND2X4 U68 ( .A(n27), .B(n138), .Y(n17) );
  NAND3BX1 U69 ( .AN(n20), .B(n2), .C(n51), .Y(n154) );
  NAND3X4 U70 ( .A(n138), .B(n34), .C(n146), .Y(n135) );
  AND2X1 U71 ( .A(n54), .B(n51), .Y(n21) );
  NAND2XL U72 ( .A(n51), .B(n3), .Y(n50) );
  OR2X4 U73 ( .A(n151), .B(n55), .Y(n13) );
  NOR2X4 U74 ( .A(n139), .B(n140), .Y(n137) );
  NAND2X4 U75 ( .A(n22), .B(n63), .Y(n66) );
  INVX4 U76 ( .A(n17), .Y(n18) );
  NAND2X4 U77 ( .A(A[8]), .B(B[8]), .Y(n36) );
  NAND2X2 U78 ( .A(n39), .B(n1), .Y(n106) );
  INVX4 U79 ( .A(n38), .Y(n164) );
  NAND3X2 U80 ( .A(n35), .B(n36), .C(n37), .Y(n31) );
  NAND2BX4 U81 ( .AN(n13), .B(n149), .Y(n100) );
  OR2X4 U82 ( .A(A[9]), .B(B[9]), .Y(n34) );
  NAND2X4 U83 ( .A(n16), .B(n164), .Y(n161) );
  NAND2X4 U84 ( .A(n159), .B(n160), .Y(n158) );
  AND2X2 U85 ( .A(n34), .B(n138), .Y(n160) );
  NAND3BX4 U86 ( .AN(n171), .B(n172), .C(n22), .Y(n35) );
  NOR3X4 U87 ( .A(n42), .B(n151), .C(n55), .Y(n172) );
  NAND3BX2 U88 ( .AN(n46), .B(n177), .C(n43), .Y(n176) );
  OAI21X1 U89 ( .A0(n96), .A1(n97), .B0(n98), .Y(n95) );
  NAND2X4 U90 ( .A(n115), .B(n114), .Y(n122) );
  AOI21X2 U91 ( .A0(n125), .A1(n118), .B0(n126), .Y(n124) );
  NAND4BX2 U92 ( .AN(n117), .B(n92), .C(n114), .D(n118), .Y(n110) );
  CLKINVX8 U93 ( .A(n127), .Y(n115) );
  INVX1 U94 ( .A(B[2]), .Y(n174) );
  NAND4BX4 U95 ( .AN(n109), .B(n110), .C(n111), .D(n112), .Y(n108) );
  NAND2X2 U96 ( .A(B[4]), .B(A[4]), .Y(n57) );
  AND2X2 U97 ( .A(n20), .B(n19), .Y(n23) );
  OR2X4 U98 ( .A(A[15]), .B(B[15]), .Y(n93) );
  INVX4 U99 ( .A(n2), .Y(n150) );
  OAI2BB1X2 U100 ( .A0N(n14), .A1N(n15), .B0(n54), .Y(n61) );
  AND2X1 U101 ( .A(n63), .B(n51), .Y(n15) );
  XOR2X2 U102 ( .A(n74), .B(n75), .Y(SUM[2]) );
  XOR2X2 U103 ( .A(n22), .B(n67), .Y(SUM[4]) );
  NAND2X2 U104 ( .A(B[1]), .B(A[1]), .Y(n78) );
  XOR2X4 U105 ( .A(n108), .B(n4), .Y(SUM[15]) );
  NAND2X4 U106 ( .A(B[9]), .B(A[9]), .Y(n33) );
  NAND2X4 U107 ( .A(n106), .B(n141), .Y(n40) );
  NOR2X2 U108 ( .A(n60), .B(n55), .Y(n59) );
  XOR2X4 U109 ( .A(n82), .B(n83), .Y(SUM[16]) );
  OAI21X4 U110 ( .A0(n84), .A1(n85), .B0(n86), .Y(n82) );
  XOR2X4 U111 ( .A(n168), .B(n5), .Y(SUM[10]) );
  XOR2X4 U112 ( .A(n155), .B(n156), .Y(SUM[11]) );
  NAND2X2 U113 ( .A(n43), .B(n47), .Y(n152) );
  NAND2X2 U114 ( .A(B[6]), .B(A[6]), .Y(n47) );
  NAND2X2 U115 ( .A(n148), .B(n44), .Y(n38) );
  XNOR2X4 U116 ( .A(n61), .B(n62), .Y(SUM[6]) );
  INVX4 U117 ( .A(n76), .Y(n80) );
  OR2X4 U118 ( .A(A[4]), .B(B[4]), .Y(n63) );
  AOI21X2 U119 ( .A0(n48), .A1(n49), .B0(n50), .Y(n45) );
  OAI21X2 U120 ( .A0(A[2]), .A1(B[2]), .B0(n71), .Y(n60) );
  NOR2X2 U121 ( .A(n139), .B(n150), .Y(n149) );
  NAND3X4 U122 ( .A(n133), .B(n134), .C(n135), .Y(n118) );
  NAND2X4 U123 ( .A(B[12]), .B(A[12]), .Y(n97) );
  OR2X4 U124 ( .A(B[1]), .B(A[1]), .Y(n76) );
  NAND3X4 U125 ( .A(n18), .B(n137), .C(n26), .Y(n127) );
  OR2X4 U126 ( .A(B[10]), .B(A[10]), .Y(n138) );
  CLKBUFX8 U127 ( .A(n56), .Y(n19) );
  NAND3X1 U128 ( .A(A[5]), .B(B[5]), .C(n2), .Y(n153) );
  NAND3X1 U129 ( .A(A[5]), .B(B[5]), .C(n2), .Y(n177) );
  OR2X4 U130 ( .A(B[6]), .B(A[6]), .Y(n24) );
  NOR2BX1 U131 ( .AN(n97), .B(n140), .Y(n143) );
  NOR2BX1 U132 ( .AN(n20), .B(n55), .Y(n67) );
  OAI2BB1X4 U133 ( .A0N(n34), .A1N(n169), .B0(n33), .Y(n168) );
  INVX1 U134 ( .A(n97), .Y(n132) );
  INVX4 U135 ( .A(n40), .Y(n144) );
  INVX1 U136 ( .A(n98), .Y(n126) );
  NAND2BX4 U137 ( .AN(n60), .B(n58), .Y(n64) );
  OAI211X2 U138 ( .A0(n121), .A1(n122), .B0(n124), .C0(n123), .Y(n119) );
  AND2X1 U139 ( .A(n33), .B(n34), .Y(n32) );
  NAND2BX4 U140 ( .AN(n100), .B(n22), .Y(n141) );
  XOR2X4 U141 ( .A(n65), .B(n21), .Y(SUM[5]) );
  NAND2X4 U142 ( .A(n19), .B(n64), .Y(n22) );
  AND2X1 U143 ( .A(n19), .B(n64), .Y(n105) );
  INVXL U144 ( .A(n99), .Y(n94) );
  NAND2XL U145 ( .A(B[3]), .B(A[3]), .Y(n56) );
  AND2X1 U146 ( .A(n133), .B(n147), .Y(n145) );
  NAND2XL U147 ( .A(B[15]), .B(A[15]), .Y(n91) );
  NOR2BX1 U148 ( .AN(n81), .B(n25), .Y(SUM[0]) );
  NOR2XL U149 ( .A(A[0]), .B(B[0]), .Y(n25) );
  INVX1 U150 ( .A(n117), .Y(n131) );
  NAND3BXL U151 ( .AN(n97), .B(n92), .C(n114), .Y(n111) );
  NAND2XL U152 ( .A(n44), .B(n3), .Y(n171) );
  AOI21X2 U153 ( .A0(n131), .A1(n118), .B0(n132), .Y(n130) );
  NOR2BXL U154 ( .AN(n36), .B(n42), .Y(n41) );
  NOR3X2 U155 ( .A(n151), .B(n150), .C(n20), .Y(n175) );
  NAND2BXL U156 ( .AN(n97), .B(n114), .Y(n123) );
  XOR2X2 U157 ( .A(n68), .B(n69), .Y(SUM[3]) );
  NOR2BX1 U158 ( .AN(n19), .B(n70), .Y(n69) );
  INVX1 U159 ( .A(n71), .Y(n70) );
  NAND4BXL U160 ( .AN(n96), .B(n101), .C(n92), .D(n93), .Y(n85) );
  INVX1 U161 ( .A(n81), .Y(n77) );
  INVXL U162 ( .A(n104), .Y(n103) );
  INVX1 U163 ( .A(n88), .Y(n86) );
  INVX1 U164 ( .A(n20), .Y(n30) );
  OAI2BB1X1 U165 ( .A0N(B[9]), .A1N(A[9]), .B0(n36), .Y(n146) );
  INVXL U166 ( .A(A[2]), .Y(n173) );
  NAND2X1 U167 ( .A(B[13]), .B(A[13]), .Y(n98) );
  NAND2XL U168 ( .A(B[14]), .B(A[14]), .Y(n99) );
  OR2XL U169 ( .A(A[11]), .B(B[11]), .Y(n28) );
  NAND2XL U170 ( .A(B[2]), .B(A[2]), .Y(n73) );
  XOR2X1 U171 ( .A(B[16]), .B(A[16]), .Y(n83) );
  AOI21X1 U172 ( .A0(n87), .A1(n102), .B0(n103), .Y(n84) );
  NAND2X1 U173 ( .A(B[5]), .B(A[5]), .Y(n54) );
  OAI21X2 U174 ( .A0(n121), .A1(n127), .B0(n130), .Y(n128) );
  AOI21X2 U175 ( .A0(B[11]), .A1(A[11]), .B0(n157), .Y(n156) );
  NAND2XL U176 ( .A(B[11]), .B(A[11]), .Y(n134) );
  NAND2XL U177 ( .A(B[11]), .B(A[11]), .Y(n147) );
  OR2X2 U178 ( .A(A[11]), .B(B[11]), .Y(n136) );
  NAND2BX4 U179 ( .AN(n30), .B(n66), .Y(n65) );
  NOR2BX1 U180 ( .AN(n78), .B(n80), .Y(n79) );
  XOR2X4 U181 ( .A(n31), .B(n32), .Y(SUM[9]) );
  XOR2X4 U182 ( .A(n40), .B(n41), .Y(SUM[8]) );
  XOR2X4 U183 ( .A(n119), .B(n120), .Y(SUM[14]) );
  OR2X4 U184 ( .A(A[14]), .B(B[14]), .Y(n92) );
  XOR2X4 U185 ( .A(n128), .B(n129), .Y(SUM[13]) );
  OR2X4 U186 ( .A(A[13]), .B(B[13]), .Y(n114) );
  NAND2BX4 U187 ( .AN(n39), .B(n141), .Y(n116) );
  XOR2X4 U188 ( .A(n142), .B(n143), .Y(SUM[12]) );
  OR2X4 U189 ( .A(A[12]), .B(B[12]), .Y(n101) );
  OAI21X4 U190 ( .A0(n144), .A1(n107), .B0(n104), .Y(n142) );
  NAND3BX4 U191 ( .AN(n152), .B(n153), .C(n154), .Y(n39) );
  OAI221X2 U192 ( .A0(n80), .A1(n81), .B0(n173), .B1(n174), .C0(n78), .Y(n58)
         );
  OR2X4 U193 ( .A(B[7]), .B(A[7]), .Y(n44) );
  OR2X4 U194 ( .A(B[8]), .B(A[8]), .Y(n148) );
  OR2X4 U195 ( .A(A[5]), .B(B[5]), .Y(n51) );
endmodule


module butterfly_DW01_sub_38 ( A, B, DIFF );
  input [16:0] A;
  input [16:0] B;
  output [16:0] DIFF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191;

  OAI21X1 U3 ( .A0(n94), .A1(n33), .B0(n113), .Y(n106) );
  NAND2BX1 U4 ( .AN(B[3]), .B(A[3]), .Y(n71) );
  NAND3X2 U5 ( .A(n144), .B(n104), .C(n145), .Y(n17) );
  NAND2X4 U6 ( .A(n165), .B(n164), .Y(n113) );
  NAND2BX4 U7 ( .AN(A[3]), .B(B[3]), .Y(n70) );
  CLKINVX3 U8 ( .A(n147), .Y(n155) );
  NAND3X4 U9 ( .A(n6), .B(n29), .C(n67), .Y(n95) );
  NAND2X4 U10 ( .A(n54), .B(n55), .Y(n50) );
  INVX8 U11 ( .A(n26), .Y(n27) );
  XOR2X4 U12 ( .A(n60), .B(n61), .Y(DIFF[5]) );
  OAI21X4 U13 ( .A0(n178), .A1(n1), .B0(n35), .Y(n181) );
  INVX4 U14 ( .A(n102), .Y(n125) );
  NAND2X4 U15 ( .A(n105), .B(n151), .Y(n150) );
  CLKINVX8 U16 ( .A(n129), .Y(n161) );
  NAND3X4 U17 ( .A(n36), .B(n112), .C(n162), .Y(n129) );
  NAND3BX4 U18 ( .AN(n37), .B(n1), .C(n28), .Y(n34) );
  NAND2BX1 U19 ( .AN(A[10]), .B(B[10]), .Y(n162) );
  CLKINVX3 U20 ( .A(n36), .Y(n178) );
  NAND3X4 U21 ( .A(n147), .B(n148), .C(n149), .Y(n140) );
  BUFX8 U22 ( .A(n38), .Y(n1) );
  INVX4 U23 ( .A(n1), .Y(n42) );
  NAND2X4 U24 ( .A(n35), .B(n1), .Y(n148) );
  INVX8 U25 ( .A(n49), .Y(n52) );
  NAND2BX4 U26 ( .AN(B[6]), .B(A[6]), .Y(n49) );
  NAND3X2 U27 ( .A(n138), .B(n139), .C(n140), .Y(n124) );
  INVX1 U28 ( .A(B[7]), .Y(n166) );
  INVX2 U29 ( .A(n62), .Y(n59) );
  OAI2BB1X2 U30 ( .A0N(n135), .A1N(n124), .B0(n136), .Y(n134) );
  NOR2X2 U31 ( .A(n103), .B(n141), .Y(n135) );
  NAND2X2 U32 ( .A(n111), .B(n161), .Y(n153) );
  NOR2BX1 U33 ( .AN(n139), .B(n174), .Y(n173) );
  NAND2BX2 U34 ( .AN(B[8]), .B(A[8]), .Y(n38) );
  INVX1 U35 ( .A(n101), .Y(n126) );
  INVX1 U36 ( .A(B[11]), .Y(n151) );
  NAND3X1 U37 ( .A(n138), .B(n139), .C(n140), .Y(n146) );
  NAND4X1 U38 ( .A(n161), .B(n111), .C(n105), .D(n40), .Y(n145) );
  AOI2BB1X2 U39 ( .A0N(n10), .A1N(n166), .B0(n167), .Y(n164) );
  INVX1 U40 ( .A(n104), .Y(n137) );
  INVX4 U41 ( .A(n40), .Y(n26) );
  INVX1 U42 ( .A(n112), .Y(n41) );
  INVX1 U43 ( .A(n109), .Y(n108) );
  OAI21XL U44 ( .A0(n96), .A1(n97), .B0(n98), .Y(n88) );
  CLKINVX3 U45 ( .A(n53), .Y(n48) );
  INVX1 U46 ( .A(n116), .Y(n46) );
  INVX1 U47 ( .A(n7), .Y(n54) );
  AND2X2 U48 ( .A(n89), .B(n100), .Y(n12) );
  NOR2X1 U49 ( .A(n45), .B(n46), .Y(n44) );
  NAND4BX1 U50 ( .AN(n41), .B(n36), .C(n110), .D(n111), .Y(n93) );
  INVX2 U51 ( .A(n105), .Y(n143) );
  OAI2BB1X4 U52 ( .A0N(B[11]), .A1N(n2), .B0(n154), .Y(n109) );
  CLKINVX20 U53 ( .A(A[11]), .Y(n2) );
  BUFX3 U54 ( .A(n76), .Y(n25) );
  AOI21X1 U55 ( .A0(n137), .A1(n130), .B0(n125), .Y(n136) );
  NAND2BX2 U56 ( .AN(B[13]), .B(A[13]), .Y(n102) );
  NAND2BX2 U57 ( .AN(A[9]), .B(B[9]), .Y(n147) );
  NAND2BX4 U58 ( .AN(B[14]), .B(A[14]), .Y(n101) );
  NAND2BX1 U59 ( .AN(B[15]), .B(A[15]), .Y(n89) );
  OAI2BB1X1 U60 ( .A0N(n58), .A1N(n186), .B0(n62), .Y(n7) );
  INVX4 U61 ( .A(n3), .Y(n4) );
  NAND2X1 U62 ( .A(n116), .B(n186), .Y(n169) );
  INVX2 U63 ( .A(n186), .Y(n3) );
  INVX4 U64 ( .A(n123), .Y(n141) );
  NAND2BXL U65 ( .AN(A[10]), .B(B[10]), .Y(n149) );
  NAND2X2 U66 ( .A(n123), .B(n146), .Y(n144) );
  OAI21X4 U67 ( .A0(n160), .A1(A[10]), .B0(n148), .Y(n156) );
  CLKINVX3 U68 ( .A(n183), .Y(n45) );
  NOR2X1 U69 ( .A(n175), .B(n35), .Y(n174) );
  NAND3X2 U70 ( .A(n4), .B(n56), .C(n57), .Y(n55) );
  NAND2X4 U71 ( .A(n82), .B(n80), .Y(n5) );
  CLKINVX4 U72 ( .A(n5), .Y(n6) );
  BUFX8 U73 ( .A(n70), .Y(n29) );
  BUFX1 U74 ( .A(n95), .Y(n13) );
  NAND2BX4 U75 ( .AN(B[10]), .B(A[10]), .Y(n139) );
  XNOR2X4 U76 ( .A(n170), .B(n8), .Y(DIFF[11]) );
  NAND2XL U77 ( .A(n111), .B(n138), .Y(n8) );
  AND2X2 U78 ( .A(n35), .B(n36), .Y(n31) );
  INVX1 U79 ( .A(A[7]), .Y(n9) );
  INVX4 U80 ( .A(n9), .Y(n10) );
  NAND2BX2 U81 ( .AN(A[2]), .B(B[2]), .Y(n67) );
  NAND2X1 U82 ( .A(n185), .B(n184), .Y(n16) );
  NAND4X2 U83 ( .A(n32), .B(n11), .C(n112), .D(n57), .Y(n39) );
  AND2X2 U84 ( .A(n56), .B(n53), .Y(n11) );
  NAND2XL U85 ( .A(n111), .B(n105), .Y(n127) );
  BUFX8 U86 ( .A(n39), .Y(n28) );
  NAND2BX4 U87 ( .AN(B[11]), .B(A[11]), .Y(n138) );
  NAND2BX4 U88 ( .AN(B[4]), .B(A[4]), .Y(n187) );
  INVX8 U89 ( .A(n130), .Y(n103) );
  OAI21X2 U90 ( .A0(n85), .A1(n86), .B0(n87), .Y(n83) );
  NAND2BX1 U91 ( .AN(B[1]), .B(A[1]), .Y(n76) );
  XOR2X4 U92 ( .A(n117), .B(n12), .Y(DIFF[15]) );
  XOR2X1 U93 ( .A(n57), .B(n63), .Y(DIFF[4]) );
  NAND2X2 U94 ( .A(n53), .B(n56), .Y(n168) );
  NAND2BX4 U95 ( .AN(A[6]), .B(B[6]), .Y(n53) );
  NAND2X1 U96 ( .A(n25), .B(n81), .Y(n190) );
  AND2X2 U97 ( .A(n116), .B(n186), .Y(n32) );
  AND3X4 U98 ( .A(n71), .B(n95), .C(n114), .Y(n14) );
  NAND3BX4 U99 ( .AN(n127), .B(n128), .C(n27), .Y(n119) );
  NOR2X2 U100 ( .A(n58), .B(n64), .Y(n63) );
  XNOR2X4 U101 ( .A(n177), .B(n15), .Y(DIFF[10]) );
  OR2X1 U102 ( .A(n175), .B(n158), .Y(n15) );
  NAND4BX4 U103 ( .AN(n118), .B(n119), .C(n120), .D(n121), .Y(n117) );
  INVX4 U104 ( .A(n31), .Y(n21) );
  XOR2X4 U105 ( .A(n17), .B(n18), .Y(DIFF[13]) );
  AND2X1 U106 ( .A(n102), .B(n130), .Y(n18) );
  NOR2X1 U107 ( .A(n104), .B(n122), .Y(n118) );
  OAI21X4 U108 ( .A0(n155), .A1(n156), .B0(n157), .Y(n154) );
  NOR2X4 U109 ( .A(n158), .B(n159), .Y(n157) );
  NOR2X4 U110 ( .A(n59), .B(n52), .Y(n185) );
  NOR2X4 U111 ( .A(n134), .B(n133), .Y(n132) );
  NAND3BX2 U112 ( .AN(n122), .B(n123), .C(n124), .Y(n121) );
  XNOR2X4 U113 ( .A(n152), .B(n19), .Y(DIFF[12]) );
  OR2X2 U114 ( .A(n143), .B(n137), .Y(n19) );
  NAND2BX4 U115 ( .AN(B[12]), .B(A[12]), .Y(n104) );
  NAND2XL U116 ( .A(n110), .B(n36), .Y(n171) );
  NAND2BX4 U117 ( .AN(A[8]), .B(B[8]), .Y(n112) );
  NOR2X2 U118 ( .A(n86), .B(n13), .Y(n91) );
  OAI2BB1X4 U119 ( .A0N(n57), .A1N(n163), .B0(n113), .Y(n40) );
  NAND2XL U120 ( .A(n99), .B(n101), .Y(n131) );
  AND2X1 U121 ( .A(n99), .B(n100), .Y(n98) );
  NAND4BX2 U122 ( .AN(n103), .B(n105), .C(n99), .D(n100), .Y(n86) );
  NOR2X4 U123 ( .A(n24), .B(n45), .Y(n184) );
  NAND2X2 U124 ( .A(n91), .B(n92), .Y(n90) );
  NOR3BX4 U125 ( .AN(n28), .B(n37), .C(n42), .Y(n172) );
  OAI21X4 U126 ( .A0(n155), .A1(n28), .B0(n179), .Y(n177) );
  OAI21X4 U127 ( .A0(n47), .A1(n48), .B0(n49), .Y(n43) );
  XOR2X4 U128 ( .A(n50), .B(n51), .Y(DIFF[6]) );
  AND3X4 U129 ( .A(n182), .B(B[6]), .C(n183), .Y(n167) );
  NAND2BX2 U130 ( .AN(A[10]), .B(B[10]), .Y(n110) );
  CLKINVX4 U131 ( .A(n138), .Y(n159) );
  AND2X4 U132 ( .A(n58), .B(n186), .Y(n24) );
  NAND2X1 U133 ( .A(n101), .B(n102), .Y(n97) );
  AOI31X2 U134 ( .A0(n16), .A1(n36), .A2(n180), .B0(n181), .Y(n179) );
  NOR2X2 U135 ( .A(n167), .B(n176), .Y(n180) );
  INVX4 U136 ( .A(n50), .Y(n47) );
  NAND2X2 U137 ( .A(n111), .B(n130), .Y(n142) );
  NAND2BX4 U138 ( .AN(A[11]), .B(B[11]), .Y(n111) );
  NAND2BX4 U139 ( .AN(B[9]), .B(A[9]), .Y(n35) );
  NAND2BX4 U140 ( .AN(A[7]), .B(B[7]), .Y(n116) );
  OAI21X4 U141 ( .A0(n10), .A1(n166), .B0(n112), .Y(n176) );
  NAND2BX2 U142 ( .AN(B[2]), .B(A[2]), .Y(n191) );
  NOR3BX4 U143 ( .AN(n165), .B(n176), .C(n167), .Y(n37) );
  OAI21X4 U144 ( .A0(n153), .A1(n26), .B0(n109), .Y(n152) );
  NAND2BX4 U145 ( .AN(B[5]), .B(A[5]), .Y(n62) );
  NOR4X2 U146 ( .A(n26), .B(n142), .C(n143), .D(n129), .Y(n133) );
  NAND2BX4 U147 ( .AN(A[15]), .B(B[15]), .Y(n100) );
  NAND2BX4 U148 ( .AN(A[12]), .B(B[12]), .Y(n105) );
  NAND2BX4 U149 ( .AN(B[7]), .B(A[7]), .Y(n183) );
  NAND2X2 U150 ( .A(n34), .B(n21), .Y(n22) );
  NAND2X4 U151 ( .A(n20), .B(n31), .Y(n23) );
  NAND2X4 U152 ( .A(n23), .B(n22), .Y(DIFF[9]) );
  INVX4 U153 ( .A(n34), .Y(n20) );
  INVX4 U154 ( .A(n187), .Y(n58) );
  NAND2BX4 U155 ( .AN(A[5]), .B(B[5]), .Y(n186) );
  NAND2BX2 U156 ( .AN(A[1]), .B(B[1]), .Y(n189) );
  NAND2BX2 U157 ( .AN(A[1]), .B(B[1]), .Y(n80) );
  NAND2X4 U158 ( .A(n14), .B(n115), .Y(n57) );
  NAND3BX4 U159 ( .AN(n188), .B(n189), .C(n190), .Y(n115) );
  AOI21X2 U160 ( .A0(n56), .A1(n57), .B0(n58), .Y(n61) );
  NAND2BX4 U161 ( .AN(A[9]), .B(B[9]), .Y(n36) );
  INVX4 U162 ( .A(n110), .Y(n175) );
  OAI21X4 U163 ( .A0(n171), .A1(n172), .B0(n173), .Y(n170) );
  NAND2BX4 U164 ( .AN(A[4]), .B(B[4]), .Y(n56) );
  INVX4 U165 ( .A(n139), .Y(n158) );
  CLKINVX3 U166 ( .A(n80), .Y(n75) );
  NAND2BX4 U167 ( .AN(A[13]), .B(B[13]), .Y(n130) );
  NOR2X1 U168 ( .A(n52), .B(n48), .Y(n51) );
  NAND2X2 U169 ( .A(n69), .B(n29), .Y(n114) );
  NOR2X2 U170 ( .A(n122), .B(n129), .Y(n128) );
  XOR2X1 U171 ( .A(n68), .B(n72), .Y(DIFF[2]) );
  AOI21X1 U172 ( .A0(n125), .A1(n99), .B0(n126), .Y(n120) );
  NOR2X1 U173 ( .A(n79), .B(n75), .Y(n78) );
  XNOR2X4 U174 ( .A(n27), .B(n30), .Y(DIFF[8]) );
  OR2X4 U175 ( .A(n41), .B(n42), .Y(n30) );
  INVXL U176 ( .A(n93), .Y(n107) );
  NAND2X4 U177 ( .A(n130), .B(n99), .Y(n122) );
  NOR2X2 U178 ( .A(n168), .B(n169), .Y(n163) );
  NAND2XL U179 ( .A(n29), .B(n71), .Y(n65) );
  AOI21XL U180 ( .A0(n67), .A1(n68), .B0(n69), .Y(n66) );
  AND3X4 U181 ( .A(n88), .B(n89), .C(n90), .Y(n87) );
  INVXL U182 ( .A(n56), .Y(n64) );
  INVXL U183 ( .A(B[10]), .Y(n160) );
  INVXL U184 ( .A(n25), .Y(n79) );
  INVX2 U185 ( .A(n191), .Y(n69) );
  NOR2X1 U186 ( .A(n93), .B(n94), .Y(n92) );
  NOR2X1 U187 ( .A(n69), .B(n73), .Y(n72) );
  INVX1 U188 ( .A(n67), .Y(n73) );
  XOR2X1 U189 ( .A(n65), .B(n66), .Y(DIFF[3]) );
  NOR2XL U190 ( .A(n103), .B(n104), .Y(n96) );
  INVXL U191 ( .A(A[6]), .Y(n182) );
  OAI21X2 U192 ( .A0(n74), .A1(n75), .B0(n25), .Y(n68) );
  INVX1 U193 ( .A(n77), .Y(n74) );
  XOR2X2 U194 ( .A(n77), .B(n78), .Y(DIFF[1]) );
  AND3X1 U195 ( .A(n114), .B(n71), .C(n115), .Y(n33) );
  XOR2X2 U196 ( .A(n84), .B(n83), .Y(DIFF[16]) );
  XNOR2X1 U197 ( .A(B[16]), .B(A[16]), .Y(n84) );
  AOI21X1 U198 ( .A0(n106), .A1(n107), .B0(n108), .Y(n85) );
  NAND2X1 U199 ( .A(n81), .B(n82), .Y(DIFF[0]) );
  NAND2BX1 U200 ( .AN(n82), .B(n81), .Y(n77) );
  NAND2BX1 U201 ( .AN(B[0]), .B(A[0]), .Y(n81) );
  NAND2BX1 U202 ( .AN(A[0]), .B(B[0]), .Y(n82) );
  NAND2X2 U203 ( .A(n29), .B(n67), .Y(n188) );
  NAND4BXL U204 ( .AN(n46), .B(n4), .C(n53), .D(n56), .Y(n94) );
  NAND2XL U205 ( .A(n4), .B(n62), .Y(n60) );
  XOR2X4 U206 ( .A(n43), .B(n44), .Y(DIFF[7]) );
  XOR2X4 U207 ( .A(n132), .B(n131), .Y(DIFF[14]) );
  NAND2BX4 U208 ( .AN(A[14]), .B(B[14]), .Y(n99) );
  OAI2BB1X4 U209 ( .A0N(A[11]), .A1N(n105), .B0(n150), .Y(n123) );
  NAND2X4 U210 ( .A(n184), .B(n185), .Y(n165) );
endmodule


module butterfly_DW01_add_52 ( A, B, SUM );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  wire   n147, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146;

  NAND3X1 U2 ( .A(n33), .B(n88), .C(n89), .Y(n87) );
  INVX4 U3 ( .A(n85), .Y(n115) );
  INVX1 U4 ( .A(n46), .Y(n1) );
  INVX4 U5 ( .A(n39), .Y(n46) );
  BUFX2 U6 ( .A(B[9]), .Y(n5) );
  NOR2X1 U7 ( .A(A[13]), .B(B[13]), .Y(n98) );
  AOI21X4 U8 ( .A0(n108), .A1(n83), .B0(n109), .Y(n107) );
  INVX2 U9 ( .A(n108), .Y(n114) );
  NAND2BX4 U10 ( .AN(n111), .B(n83), .Y(n105) );
  XOR2X4 U11 ( .A(n59), .B(n60), .Y(SUM[3]) );
  BUFX8 U12 ( .A(n128), .Y(n2) );
  NAND2XL U13 ( .A(B[10]), .B(A[10]), .Y(n128) );
  INVX1 U14 ( .A(n91), .Y(n62) );
  NAND3BX1 U15 ( .AN(n90), .B(n91), .C(n92), .Y(n86) );
  NAND2X1 U16 ( .A(B[0]), .B(A[0]), .Y(n71) );
  OR2X2 U17 ( .A(A[7]), .B(B[7]), .Y(n43) );
  CLKINVX3 U18 ( .A(n88), .Y(n133) );
  INVX1 U19 ( .A(n32), .Y(n27) );
  NAND2X2 U20 ( .A(n122), .B(n123), .Y(n120) );
  NAND2X2 U21 ( .A(n122), .B(n123), .Y(n124) );
  NOR2BX1 U22 ( .AN(n49), .B(n48), .Y(n51) );
  NAND2X2 U23 ( .A(n14), .B(n15), .Y(SUM[8]) );
  NAND2X1 U24 ( .A(n12), .B(n36), .Y(n15) );
  INVX4 U25 ( .A(n77), .Y(n3) );
  CLKINVX3 U26 ( .A(n3), .Y(n4) );
  NOR2X1 U27 ( .A(n24), .B(n145), .Y(n141) );
  NOR2X2 U28 ( .A(A[1]), .B(B[1]), .Y(n145) );
  OR2X2 U29 ( .A(A[1]), .B(B[1]), .Y(n67) );
  INVX2 U30 ( .A(n52), .Y(n48) );
  NAND2X1 U31 ( .A(n84), .B(n97), .Y(n6) );
  NAND2X2 U32 ( .A(B[11]), .B(A[11]), .Y(n126) );
  NAND3X2 U33 ( .A(n83), .B(n84), .C(n85), .Y(n79) );
  OR2X4 U34 ( .A(n76), .B(n77), .Y(n10) );
  NAND2X1 U35 ( .A(B[6]), .B(A[6]), .Y(n42) );
  INVX3 U36 ( .A(n33), .Y(n146) );
  XNOR2X4 U37 ( .A(n104), .B(n6), .Y(SUM[15]) );
  NAND3X4 U38 ( .A(n88), .B(n5), .C(A[9]), .Y(n127) );
  AOI21X4 U39 ( .A0(n1), .A1(n40), .B0(n41), .Y(n38) );
  NAND2X2 U40 ( .A(B[2]), .B(A[2]), .Y(n64) );
  NAND2XL U41 ( .A(n33), .B(n34), .Y(n20) );
  CLKINVX8 U42 ( .A(n147), .Y(n16) );
  OR2X2 U43 ( .A(A[3]), .B(B[3]), .Y(n91) );
  AOI21X2 U44 ( .A0(n86), .A1(n138), .B0(n87), .Y(n76) );
  NAND4X2 U45 ( .A(n25), .B(n88), .C(n33), .D(n89), .Y(n93) );
  CLKINVX2 U46 ( .A(n84), .Y(n103) );
  NOR2X4 U47 ( .A(n102), .B(n103), .Y(n94) );
  XOR2X2 U48 ( .A(n40), .B(n45), .Y(SUM[6]) );
  NAND2X1 U49 ( .A(A[12]), .B(B[12]), .Y(n99) );
  NAND2X2 U50 ( .A(B[12]), .B(A[12]), .Y(n116) );
  NAND2X4 U51 ( .A(B[1]), .B(A[1]), .Y(n69) );
  XOR2X4 U52 ( .A(n37), .B(n38), .Y(n147) );
  INVX2 U53 ( .A(n83), .Y(n102) );
  OAI211X2 U54 ( .A0(n98), .A1(n99), .B0(n100), .C0(n101), .Y(n95) );
  INVX4 U55 ( .A(n134), .Y(n132) );
  OAI2BB1X1 U56 ( .A0N(B[11]), .A1N(A[11]), .B0(n82), .Y(n7) );
  CLKINVX20 U57 ( .A(n7), .Y(n131) );
  AOI21X1 U58 ( .A0(n138), .A1(n30), .B0(n31), .Y(n28) );
  NAND3BX4 U59 ( .AN(n54), .B(n52), .C(n39), .Y(n139) );
  BUFX8 U60 ( .A(A[4]), .Y(n8) );
  NOR2X4 U61 ( .A(n79), .B(n80), .Y(n78) );
  INVX8 U62 ( .A(n110), .Y(n117) );
  AOI21X4 U63 ( .A0(n94), .A1(n95), .B0(n96), .Y(n74) );
  OAI2BB1X4 U64 ( .A0N(n141), .A1N(n142), .B0(n143), .Y(n92) );
  NAND3X2 U65 ( .A(n30), .B(n32), .C(n29), .Y(n137) );
  NAND2X4 U66 ( .A(n55), .B(n56), .Y(n53) );
  NAND4X4 U67 ( .A(n125), .B(n2), .C(n126), .D(n127), .Y(n77) );
  AND2X4 U68 ( .A(n77), .B(n82), .Y(n11) );
  OAI21X4 U69 ( .A0(n47), .A1(n48), .B0(n49), .Y(n40) );
  NAND3BX4 U70 ( .AN(n32), .B(n33), .C(n88), .Y(n125) );
  AOI2BB2X4 U71 ( .B0(B[7]), .B1(A[7]), .A0N(n46), .A1N(n49), .Y(n140) );
  NOR2X4 U72 ( .A(A[2]), .B(B[2]), .Y(n24) );
  NOR2BXL U73 ( .AN(n64), .B(n24), .Y(n66) );
  NOR2BX4 U74 ( .AN(n2), .B(n133), .Y(n135) );
  NOR2X4 U75 ( .A(n11), .B(n117), .Y(n106) );
  NAND2X2 U76 ( .A(n129), .B(n43), .Y(n138) );
  AOI21X4 U77 ( .A0(n4), .A1(n82), .B0(n117), .Y(n113) );
  BUFX8 U78 ( .A(B[4]), .Y(n9) );
  OAI21X4 U79 ( .A0(n113), .A1(n111), .B0(n114), .Y(n112) );
  NAND2X4 U80 ( .A(B[5]), .B(A[5]), .Y(n49) );
  INVX4 U81 ( .A(n89), .Y(n31) );
  XOR2X4 U82 ( .A(n20), .B(n21), .Y(SUM[9]) );
  INVX4 U83 ( .A(n50), .Y(n47) );
  XOR2X4 U84 ( .A(n23), .B(n124), .Y(SUM[12]) );
  NAND2BX4 U85 ( .AN(n93), .B(n35), .Y(n110) );
  NAND2X4 U86 ( .A(n81), .B(n85), .Y(n111) );
  NAND2X4 U87 ( .A(n10), .B(n78), .Y(n75) );
  NAND2XL U88 ( .A(n13), .B(n35), .Y(n14) );
  INVXL U89 ( .A(n35), .Y(n12) );
  INVX1 U90 ( .A(n36), .Y(n13) );
  INVX8 U91 ( .A(n16), .Y(SUM[7]) );
  NAND4X2 U92 ( .A(n26), .B(n55), .C(n52), .D(n39), .Y(n90) );
  NAND2X2 U93 ( .A(A[3]), .B(B[3]), .Y(n61) );
  INVX1 U94 ( .A(n101), .Y(n109) );
  NOR2BX2 U95 ( .AN(n32), .B(n31), .Y(n36) );
  NAND2X4 U96 ( .A(n129), .B(n43), .Y(n29) );
  XOR2X1 U97 ( .A(n50), .B(n51), .Y(SUM[5]) );
  NOR2BX4 U98 ( .AN(n92), .B(n62), .Y(n56) );
  XNOR2X4 U99 ( .A(n134), .B(n18), .Y(SUM[10]) );
  CLKINVX20 U100 ( .A(n135), .Y(n18) );
  AND2X1 U101 ( .A(n116), .B(n81), .Y(n23) );
  INVX2 U102 ( .A(n97), .Y(n96) );
  AND2X1 U103 ( .A(n83), .B(n101), .Y(n19) );
  INVXL U104 ( .A(n55), .Y(n58) );
  NOR2BXL U105 ( .AN(n61), .B(n62), .Y(n60) );
  NOR2X2 U106 ( .A(n27), .B(n28), .Y(n21) );
  OAI2BB1XL U107 ( .A0N(n67), .A1N(n68), .B0(n69), .Y(n65) );
  INVXL U108 ( .A(n42), .Y(n41) );
  OR2X4 U109 ( .A(A[8]), .B(B[8]), .Y(n89) );
  NOR2BX1 U110 ( .AN(n71), .B(n22), .Y(SUM[0]) );
  NOR2XL U111 ( .A(A[0]), .B(B[0]), .Y(n22) );
  XOR2X1 U112 ( .A(n65), .B(n66), .Y(SUM[2]) );
  NAND2XL U113 ( .A(n85), .B(n100), .Y(n118) );
  INVX1 U114 ( .A(n116), .Y(n121) );
  NOR2X2 U115 ( .A(n31), .B(n146), .Y(n136) );
  NAND2X2 U116 ( .A(n81), .B(n82), .Y(n80) );
  XOR2X1 U117 ( .A(n56), .B(n57), .Y(SUM[4]) );
  NOR2BX1 U118 ( .AN(n54), .B(n58), .Y(n57) );
  NOR2BX1 U119 ( .AN(n42), .B(n46), .Y(n45) );
  OAI21XL U120 ( .A0(n63), .A1(n24), .B0(n64), .Y(n59) );
  INVX1 U121 ( .A(n65), .Y(n63) );
  XOR2X1 U122 ( .A(n68), .B(n70), .Y(SUM[1]) );
  NOR2BX1 U123 ( .AN(n69), .B(n145), .Y(n70) );
  NAND2X2 U124 ( .A(n53), .B(n54), .Y(n50) );
  NAND2X1 U125 ( .A(n71), .B(n69), .Y(n142) );
  NOR2BX2 U126 ( .AN(n64), .B(n144), .Y(n143) );
  INVX1 U127 ( .A(n61), .Y(n144) );
  INVX1 U128 ( .A(n71), .Y(n68) );
  OR2X4 U129 ( .A(A[11]), .B(B[11]), .Y(n25) );
  OR2X4 U130 ( .A(A[7]), .B(B[7]), .Y(n26) );
  NAND2XL U131 ( .A(n43), .B(n44), .Y(n37) );
  NAND2XL U132 ( .A(B[7]), .B(A[7]), .Y(n44) );
  NAND2X2 U133 ( .A(B[13]), .B(A[13]), .Y(n100) );
  NAND2X2 U134 ( .A(B[14]), .B(A[14]), .Y(n101) );
  NAND2X2 U135 ( .A(n9), .B(n8), .Y(n54) );
  NAND2X1 U136 ( .A(A[15]), .B(B[15]), .Y(n97) );
  NAND2X4 U137 ( .A(n74), .B(n75), .Y(n72) );
  NAND2XL U138 ( .A(n5), .B(A[9]), .Y(n34) );
  XOR2X4 U139 ( .A(n72), .B(n73), .Y(SUM[16]) );
  XOR2X4 U140 ( .A(B[16]), .B(A[16]), .Y(n73) );
  OR2X4 U141 ( .A(B[15]), .B(A[15]), .Y(n84) );
  OAI21X4 U142 ( .A0(n105), .A1(n106), .B0(n107), .Y(n104) );
  XOR2X4 U143 ( .A(n112), .B(n19), .Y(SUM[14]) );
  OR2X4 U144 ( .A(A[14]), .B(B[14]), .Y(n83) );
  OAI21X4 U145 ( .A0(n115), .A1(n116), .B0(n100), .Y(n108) );
  XOR2X4 U146 ( .A(n118), .B(n119), .Y(SUM[13]) );
  AOI21X4 U147 ( .A0(n120), .A1(n81), .B0(n121), .Y(n119) );
  OR2X4 U148 ( .A(A[13]), .B(B[13]), .Y(n85) );
  NAND2X4 U149 ( .A(n77), .B(n82), .Y(n123) );
  NAND2BX4 U150 ( .AN(n93), .B(n35), .Y(n122) );
  NAND2X4 U151 ( .A(n29), .B(n30), .Y(n35) );
  NAND2BX4 U152 ( .AN(n90), .B(n56), .Y(n30) );
  OR2X4 U153 ( .A(A[12]), .B(B[12]), .Y(n81) );
  XOR2X4 U154 ( .A(n130), .B(n131), .Y(SUM[11]) );
  OR2X4 U155 ( .A(A[11]), .B(B[11]), .Y(n82) );
  OAI21X4 U156 ( .A0(n132), .A1(n133), .B0(n2), .Y(n130) );
  OR2X4 U157 ( .A(A[10]), .B(B[10]), .Y(n88) );
  OAI2BB1X4 U158 ( .A0N(n136), .A1N(n137), .B0(n34), .Y(n134) );
  NAND3X4 U159 ( .A(n140), .B(n42), .C(n139), .Y(n129) );
  NAND2X4 U160 ( .A(B[8]), .B(A[8]), .Y(n32) );
  OR2X4 U161 ( .A(A[6]), .B(B[6]), .Y(n39) );
  OR2X4 U162 ( .A(A[5]), .B(B[5]), .Y(n52) );
  OR2X4 U163 ( .A(n8), .B(n9), .Y(n55) );
  OR2X4 U164 ( .A(A[9]), .B(B[9]), .Y(n33) );
endmodule


module butterfly_DW01_add_64 ( A, B, SUM );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  wire   n158, n159, n160, n1, n2, n3, n4, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157;

  XOR2X4 U2 ( .A(n35), .B(n30), .Y(SUM[9]) );
  NAND4BBX4 U3 ( .AN(n8), .BN(n116), .C(n36), .D(n85), .Y(n114) );
  INVX1 U4 ( .A(n97), .Y(n1) );
  CLKINVX3 U5 ( .A(n36), .Y(n2) );
  INVX4 U6 ( .A(n2), .Y(n3) );
  INVX8 U7 ( .A(n86), .Y(n96) );
  BUFX3 U8 ( .A(A[12]), .Y(n4) );
  NAND3X4 U9 ( .A(n29), .B(n94), .C(n95), .Y(n78) );
  INVX8 U10 ( .A(n57), .Y(n55) );
  INVX4 U11 ( .A(n51), .Y(n48) );
  OR2X4 U12 ( .A(A[1]), .B(n16), .Y(n70) );
  OAI21X4 U13 ( .A0(n42), .A1(n43), .B0(n44), .Y(n39) );
  BUFX3 U14 ( .A(n160), .Y(SUM[4]) );
  INVX8 U15 ( .A(n7), .Y(SUM[6]) );
  XOR2X2 U16 ( .A(n60), .B(n61), .Y(SUM[3]) );
  BUFX3 U17 ( .A(n159), .Y(SUM[5]) );
  OAI21X2 U18 ( .A0(n98), .A1(n93), .B0(n32), .Y(n94) );
  NAND2X2 U19 ( .A(B[13]), .B(A[13]), .Y(n90) );
  BUFX3 U20 ( .A(n99), .Y(n32) );
  INVX4 U21 ( .A(n80), .Y(n11) );
  BUFX3 U22 ( .A(B[1]), .Y(n16) );
  OR2X2 U23 ( .A(A[4]), .B(B[4]), .Y(n59) );
  INVX1 U24 ( .A(n70), .Y(n74) );
  INVX1 U25 ( .A(n59), .Y(n54) );
  XOR2X1 U26 ( .A(n51), .B(n52), .Y(n159) );
  NOR2BX1 U27 ( .AN(n50), .B(n49), .Y(n52) );
  INVX1 U28 ( .A(n22), .Y(n144) );
  NOR2X2 U29 ( .A(A[7]), .B(B[7]), .Y(n27) );
  XNOR2X4 U30 ( .A(n45), .B(n46), .Y(n7) );
  AND2X2 U31 ( .A(A[9]), .B(B[9]), .Y(n15) );
  BUFX3 U32 ( .A(B[12]), .Y(n18) );
  NOR2BX2 U33 ( .AN(n105), .B(n117), .Y(n131) );
  NAND4BX1 U34 ( .AN(n140), .B(n141), .C(n34), .D(n142), .Y(n8) );
  NAND2X4 U35 ( .A(B[8]), .B(A[8]), .Y(n135) );
  NAND2X1 U36 ( .A(B[14]), .B(A[14]), .Y(n89) );
  OAI21X4 U37 ( .A0(n82), .A1(n83), .B0(n84), .Y(n81) );
  XNOR2X4 U38 ( .A(n25), .B(n9), .Y(SUM[13]) );
  CLKINVX20 U39 ( .A(n26), .Y(n9) );
  OR2X2 U40 ( .A(A[7]), .B(B[7]), .Y(n41) );
  XNOR2X4 U41 ( .A(n10), .B(n130), .Y(SUM[12]) );
  AND2X1 U42 ( .A(n91), .B(n127), .Y(n10) );
  NAND2X2 U43 ( .A(B[10]), .B(A[10]), .Y(n110) );
  NAND2X1 U44 ( .A(n84), .B(n86), .Y(n111) );
  NAND4BX4 U45 ( .AN(n27), .B(n59), .C(n53), .D(n47), .Y(n93) );
  XNOR2X4 U46 ( .A(n76), .B(n12), .Y(SUM[16]) );
  XNOR2X4 U47 ( .A(B[16]), .B(A[16]), .Y(n12) );
  INVX1 U48 ( .A(A[11]), .Y(n106) );
  NOR2X2 U49 ( .A(A[11]), .B(B[11]), .Y(n140) );
  INVX1 U50 ( .A(B[11]), .Y(n107) );
  XNOR2X4 U51 ( .A(n13), .B(n111), .Y(SUM[15]) );
  NAND3X4 U52 ( .A(n113), .B(n112), .C(n114), .Y(n13) );
  NOR2BX2 U53 ( .AN(n135), .B(n38), .Y(n37) );
  NAND2X4 U54 ( .A(n109), .B(n110), .Y(n132) );
  BUFX1 U55 ( .A(A[5]), .Y(n21) );
  NAND3X2 U56 ( .A(n21), .B(B[5]), .C(n47), .Y(n154) );
  AND2X4 U57 ( .A(n80), .B(n91), .Y(n29) );
  NOR2X4 U58 ( .A(A[9]), .B(B[9]), .Y(n138) );
  NAND3X4 U59 ( .A(n129), .B(n128), .C(n127), .Y(n25) );
  NAND3BX2 U60 ( .AN(n117), .B(n105), .C(n91), .Y(n128) );
  NAND2X4 U61 ( .A(n14), .B(n15), .Y(n108) );
  OR2X4 U62 ( .A(B[10]), .B(A[10]), .Y(n14) );
  NAND4BX2 U63 ( .AN(n117), .B(n118), .C(n1), .D(n105), .Y(n113) );
  NAND2XL U64 ( .A(n109), .B(n110), .Y(n101) );
  NAND3BX2 U65 ( .AN(n11), .B(n36), .C(n91), .Y(n129) );
  CLKINVX8 U66 ( .A(n115), .Y(n80) );
  NAND2X2 U67 ( .A(B[11]), .B(A[11]), .Y(n134) );
  NAND2X4 U68 ( .A(n4), .B(n18), .Y(n126) );
  XNOR2X4 U69 ( .A(n121), .B(n17), .Y(SUM[14]) );
  AND2X1 U70 ( .A(n85), .B(n89), .Y(n17) );
  NOR2X4 U71 ( .A(n87), .B(n88), .Y(n82) );
  NAND2X2 U72 ( .A(n89), .B(n90), .Y(n88) );
  AOI21X2 U73 ( .A0(n80), .A1(n36), .B0(n131), .Y(n130) );
  NOR2X4 U74 ( .A(A[13]), .B(B[13]), .Y(n19) );
  INVX8 U75 ( .A(n116), .Y(n118) );
  AND2X1 U76 ( .A(n92), .B(n90), .Y(n26) );
  NAND2X2 U77 ( .A(n91), .B(n105), .Y(n104) );
  NAND2X1 U78 ( .A(n110), .B(n141), .Y(n149) );
  OAI2BB1X2 U79 ( .A0N(n145), .A1N(n146), .B0(n110), .Y(n143) );
  NAND2X4 U80 ( .A(n108), .B(n134), .Y(n133) );
  AOI21X2 U81 ( .A0(n119), .A1(n85), .B0(n120), .Y(n112) );
  NAND2X4 U82 ( .A(n91), .B(n92), .Y(n116) );
  NAND2X1 U83 ( .A(B[6]), .B(A[6]), .Y(n44) );
  NOR2X4 U84 ( .A(n19), .B(n126), .Y(n87) );
  INVX4 U85 ( .A(n81), .Y(n79) );
  NAND2X2 U86 ( .A(n85), .B(n86), .Y(n83) );
  NAND2X4 U87 ( .A(n118), .B(n105), .Y(n124) );
  CLKBUFXL U88 ( .A(B[4]), .Y(n20) );
  NAND4X4 U89 ( .A(n44), .B(n152), .C(n153), .D(n154), .Y(n139) );
  NAND4X2 U90 ( .A(n20), .B(A[4]), .C(n47), .D(n53), .Y(n152) );
  INVX8 U91 ( .A(n85), .Y(n97) );
  NOR2BX2 U92 ( .AN(n118), .B(n11), .Y(n122) );
  AOI21X4 U93 ( .A0(n122), .A1(n3), .B0(n123), .Y(n121) );
  OAI2BB1X1 U94 ( .A0N(B[11]), .A1N(A[11]), .B0(n105), .Y(n22) );
  XOR2X4 U95 ( .A(n143), .B(n144), .Y(SUM[11]) );
  OAI21X4 U96 ( .A0(n101), .A1(n102), .B0(n103), .Y(n77) );
  OAI21X4 U97 ( .A0(n19), .A1(n126), .B0(n90), .Y(n119) );
  NAND4X1 U98 ( .A(n33), .B(n135), .C(n147), .D(n148), .Y(n146) );
  OAI21X2 U99 ( .A0(n124), .A1(n117), .B0(n125), .Y(n123) );
  AOI21X4 U100 ( .A0(n35), .A1(n34), .B0(n151), .Y(n150) );
  NAND3BX4 U101 ( .AN(n38), .B(n57), .C(n155), .Y(n147) );
  INVX4 U102 ( .A(n142), .Y(n38) );
  NAND3X2 U103 ( .A(n147), .B(n135), .C(n148), .Y(n35) );
  NAND3X2 U104 ( .A(n142), .B(n41), .C(n139), .Y(n148) );
  NAND2X4 U105 ( .A(n62), .B(n100), .Y(n57) );
  NAND2X4 U106 ( .A(B[3]), .B(A[3]), .Y(n62) );
  XOR2X4 U107 ( .A(n39), .B(n40), .Y(SUM[7]) );
  NOR4X4 U108 ( .A(n104), .B(n96), .C(n97), .D(n19), .Y(n103) );
  BUFX12 U109 ( .A(n158), .Y(SUM[8]) );
  XOR2X2 U110 ( .A(n36), .B(n37), .Y(n158) );
  XOR2X4 U111 ( .A(n149), .B(n150), .Y(SUM[10]) );
  NOR2BX1 U112 ( .AN(n44), .B(n43), .Y(n46) );
  NOR2BX1 U113 ( .AN(n56), .B(n54), .Y(n58) );
  NOR2XL U114 ( .A(A[0]), .B(B[0]), .Y(n28) );
  OR2X4 U115 ( .A(B[6]), .B(A[6]), .Y(n47) );
  OAI21X4 U116 ( .A0(n55), .A1(n93), .B0(n99), .Y(n36) );
  CLKINVX3 U117 ( .A(n119), .Y(n125) );
  OAI21X4 U118 ( .A0(n54), .A1(n55), .B0(n56), .Y(n51) );
  OAI21XL U119 ( .A0(n106), .A1(n107), .B0(n108), .Y(n102) );
  OAI21X4 U120 ( .A0(n48), .A1(n49), .B0(n50), .Y(n45) );
  AND2X1 U121 ( .A(n34), .B(n141), .Y(n145) );
  INVXL U122 ( .A(n69), .Y(n65) );
  INVXL U123 ( .A(n75), .Y(n71) );
  INVX2 U124 ( .A(n45), .Y(n42) );
  NOR2X4 U125 ( .A(B[10]), .B(A[10]), .Y(n137) );
  NAND2X4 U126 ( .A(n31), .B(n156), .Y(n100) );
  AND2X1 U127 ( .A(n62), .B(n100), .Y(n98) );
  NOR2BX1 U128 ( .AN(n75), .B(n28), .Y(SUM[0]) );
  INVX1 U129 ( .A(n47), .Y(n43) );
  INVX1 U130 ( .A(n67), .Y(n64) );
  INVX1 U131 ( .A(n33), .Y(n151) );
  INVX1 U132 ( .A(n89), .Y(n120) );
  XOR2X1 U133 ( .A(n57), .B(n58), .Y(n160) );
  XOR2X1 U134 ( .A(n67), .B(n68), .Y(SUM[2]) );
  NOR2BX1 U135 ( .AN(n66), .B(n65), .Y(n68) );
  AND2X1 U136 ( .A(n33), .B(n34), .Y(n30) );
  INVX1 U137 ( .A(n93), .Y(n155) );
  XOR2X1 U138 ( .A(n71), .B(n73), .Y(SUM[1]) );
  NOR2BXL U139 ( .AN(n72), .B(n74), .Y(n73) );
  OAI2BB1X1 U140 ( .A0N(n70), .A1N(n71), .B0(n72), .Y(n67) );
  NOR2BX1 U141 ( .AN(n62), .B(n63), .Y(n61) );
  OAI21XL U142 ( .A0(n64), .A1(n65), .B0(n66), .Y(n60) );
  INVX1 U143 ( .A(n157), .Y(n63) );
  NAND2XL U144 ( .A(B[9]), .B(A[9]), .Y(n33) );
  NAND2X2 U145 ( .A(B[2]), .B(A[2]), .Y(n66) );
  NAND2X1 U146 ( .A(B[0]), .B(A[0]), .Y(n75) );
  NAND2X1 U147 ( .A(n16), .B(A[1]), .Y(n72) );
  NAND2XL U148 ( .A(B[15]), .B(A[15]), .Y(n84) );
  AND2X4 U149 ( .A(n69), .B(n157), .Y(n31) );
  NAND2XL U150 ( .A(B[4]), .B(A[4]), .Y(n56) );
  NAND2XL U151 ( .A(B[5]), .B(A[5]), .Y(n50) );
  NAND2XL U152 ( .A(n18), .B(n4), .Y(n127) );
  OR2X2 U153 ( .A(A[2]), .B(B[2]), .Y(n69) );
  NAND2X1 U154 ( .A(B[7]), .B(A[7]), .Y(n153) );
  AOI21XL U155 ( .A0(B[7]), .A1(A[7]), .B0(n27), .Y(n40) );
  NOR3X2 U156 ( .A(n96), .B(n97), .C(n19), .Y(n95) );
  CLKINVX3 U157 ( .A(n53), .Y(n49) );
  NAND3X4 U158 ( .A(n77), .B(n78), .C(n79), .Y(n76) );
  OR2X4 U159 ( .A(A[15]), .B(B[15]), .Y(n86) );
  OR2X4 U160 ( .A(B[14]), .B(A[14]), .Y(n85) );
  OR2X4 U161 ( .A(A[13]), .B(B[13]), .Y(n92) );
  NOR2X4 U162 ( .A(n132), .B(n133), .Y(n117) );
  NAND2BX4 U163 ( .AN(n135), .B(n136), .Y(n109) );
  NOR2X4 U164 ( .A(n137), .B(n138), .Y(n136) );
  NAND2X4 U165 ( .A(n139), .B(n41), .Y(n99) );
  NAND4BX4 U166 ( .AN(n140), .B(n141), .C(n34), .D(n142), .Y(n115) );
  OR2X4 U167 ( .A(B[12]), .B(A[12]), .Y(n91) );
  OR2X4 U168 ( .A(A[11]), .B(B[11]), .Y(n105) );
  OR2X4 U169 ( .A(A[5]), .B(B[5]), .Y(n53) );
  OAI211X2 U170 ( .A0(n74), .A1(n75), .B0(n72), .C0(n66), .Y(n156) );
  OR2X4 U171 ( .A(A[3]), .B(B[3]), .Y(n157) );
  OR2X4 U172 ( .A(A[8]), .B(B[8]), .Y(n142) );
  OR2X4 U173 ( .A(A[9]), .B(B[9]), .Y(n34) );
  OR2X4 U174 ( .A(A[10]), .B(B[10]), .Y(n141) );
endmodule


module butterfly_DW01_add_69 ( A, B, SUM );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179;

  OAI21X2 U2 ( .A0(A[11]), .A1(B[11]), .B0(n143), .Y(n151) );
  NAND2X2 U3 ( .A(n162), .B(n17), .Y(n161) );
  OAI2BB1X4 U4 ( .A0N(n118), .A1N(n110), .B0(n114), .Y(n116) );
  NAND2X2 U5 ( .A(B[10]), .B(A[10]), .Y(n139) );
  XOR2X2 U6 ( .A(n67), .B(n68), .Y(SUM[2]) );
  NAND2X2 U7 ( .A(n39), .B(n44), .Y(n48) );
  NAND3X2 U8 ( .A(A[1]), .B(n7), .C(n69), .Y(n57) );
  CLKINVX2 U9 ( .A(n93), .Y(n133) );
  AND2X2 U10 ( .A(n140), .B(n21), .Y(n15) );
  INVXL U11 ( .A(n22), .Y(n4) );
  AND2X2 U12 ( .A(n102), .B(n142), .Y(n16) );
  AND2X2 U13 ( .A(n45), .B(n1), .Y(n146) );
  NOR2X1 U14 ( .A(n44), .B(n105), .Y(n163) );
  OR3X2 U15 ( .A(n105), .B(n149), .C(n179), .Y(n160) );
  CLKINVX3 U16 ( .A(n171), .Y(n162) );
  NAND2X2 U17 ( .A(n101), .B(n102), .Y(n136) );
  NOR2BX2 U18 ( .AN(n17), .B(n93), .Y(n135) );
  AOI21X1 U19 ( .A0(n112), .A1(n85), .B0(n113), .Y(n111) );
  INVX1 U20 ( .A(n75), .Y(n71) );
  INVX1 U21 ( .A(n69), .Y(n65) );
  OAI2BB1X1 U22 ( .A0N(n70), .A1N(n71), .B0(n72), .Y(n67) );
  NOR2X2 U23 ( .A(n63), .B(n52), .Y(n51) );
  NAND2X1 U24 ( .A(B[9]), .B(A[9]), .Y(n140) );
  NAND3X2 U25 ( .A(n26), .B(n17), .C(n28), .Y(n23) );
  OR2X2 U26 ( .A(A[11]), .B(B[11]), .Y(n142) );
  NAND2BX1 U27 ( .AN(n102), .B(n120), .Y(n127) );
  NOR2BX1 U28 ( .AN(n120), .B(n93), .Y(n125) );
  INVX1 U29 ( .A(n115), .Y(n118) );
  NAND3BX1 U30 ( .AN(n63), .B(n104), .C(n19), .Y(n103) );
  OAI21XL U31 ( .A0(n82), .A1(n83), .B0(n84), .Y(n81) );
  NAND2X2 U32 ( .A(B[0]), .B(A[0]), .Y(n75) );
  NOR2BX1 U33 ( .AN(n66), .B(n65), .Y(n68) );
  NOR2BX1 U34 ( .AN(n92), .B(n98), .Y(n130) );
  NOR2BX2 U35 ( .AN(n56), .B(n63), .Y(n62) );
  INVX4 U36 ( .A(n54), .Y(n63) );
  NAND2X1 U37 ( .A(B[8]), .B(A[8]), .Y(n22) );
  NAND2X2 U38 ( .A(A[6]), .B(B[6]), .Y(n1) );
  INVXL U39 ( .A(n143), .Y(n154) );
  NOR2X1 U40 ( .A(n25), .B(n93), .Y(n129) );
  CLKINVX3 U41 ( .A(n6), .Y(n7) );
  NOR2XL U42 ( .A(n134), .B(n63), .Y(n169) );
  CLKBUFXL U43 ( .A(n28), .Y(n2) );
  NAND2XL U44 ( .A(n101), .B(n102), .Y(n100) );
  NAND2X1 U45 ( .A(n17), .B(n45), .Y(n35) );
  NAND2X4 U46 ( .A(B[7]), .B(A[7]), .Y(n45) );
  NOR3BX4 U47 ( .AN(n155), .B(n156), .C(n157), .Y(n153) );
  NAND2X4 U48 ( .A(n3), .B(n145), .Y(n28) );
  AND2X4 U49 ( .A(n144), .B(n146), .Y(n3) );
  NOR2BX2 U50 ( .AN(n139), .B(n154), .Y(n167) );
  NAND3BX4 U51 ( .AN(n4), .B(n23), .C(n24), .Y(n5) );
  XOR2X4 U52 ( .A(n5), .B(n15), .Y(SUM[9]) );
  NAND2X1 U53 ( .A(n41), .B(n42), .Y(n40) );
  INVX4 U54 ( .A(n42), .Y(n105) );
  NAND3BX2 U55 ( .AN(n147), .B(n42), .C(n148), .Y(n145) );
  NAND4BX2 U56 ( .AN(n25), .B(n26), .C(n17), .D(n27), .Y(n24) );
  XOR2X4 U57 ( .A(n27), .B(n59), .Y(SUM[4]) );
  AND2X1 U58 ( .A(n45), .B(n1), .Y(n176) );
  OAI21X4 U59 ( .A0(n64), .A1(n65), .B0(n66), .Y(n61) );
  NAND2X2 U60 ( .A(B[5]), .B(A[5]), .Y(n43) );
  OR2X4 U61 ( .A(A[5]), .B(B[5]), .Y(n41) );
  AOI21X4 U62 ( .A0(n135), .A1(n28), .B0(n136), .Y(n131) );
  NAND2X4 U63 ( .A(n172), .B(n69), .Y(n55) );
  OR2X4 U64 ( .A(A[12]), .B(B[12]), .Y(n120) );
  INVX2 U65 ( .A(n86), .Y(n96) );
  NAND2X2 U66 ( .A(B[11]), .B(A[11]), .Y(n102) );
  NOR2X1 U67 ( .A(A[5]), .B(B[5]), .Y(n147) );
  NOR2X4 U68 ( .A(n25), .B(n171), .Y(n170) );
  NAND2X4 U69 ( .A(n168), .B(n155), .Y(n166) );
  NAND3X4 U70 ( .A(n27), .B(n17), .C(n170), .Y(n155) );
  NAND2X2 U71 ( .A(B[14]), .B(A[14]), .Y(n89) );
  NOR2BX1 U72 ( .AN(n89), .B(n97), .Y(n117) );
  NAND3X4 U73 ( .A(n139), .B(n140), .C(n141), .Y(n138) );
  NAND3X2 U74 ( .A(A[8]), .B(B[8]), .C(n21), .Y(n141) );
  OR2X4 U75 ( .A(A[8]), .B(B[8]), .Y(n26) );
  NAND3BX1 U76 ( .AN(n128), .B(n169), .C(n129), .Y(n123) );
  INVX4 U77 ( .A(n17), .Y(n34) );
  OR2X2 U78 ( .A(A[5]), .B(B[5]), .Y(n20) );
  NOR2BX2 U79 ( .AN(n44), .B(n60), .Y(n59) );
  NOR2X4 U80 ( .A(n75), .B(n74), .Y(n172) );
  NOR2BX2 U81 ( .AN(n72), .B(n74), .Y(n73) );
  INVX3 U82 ( .A(n70), .Y(n74) );
  AOI21X4 U83 ( .A0(n38), .A1(n39), .B0(n40), .Y(n37) );
  AND2X4 U84 ( .A(n39), .B(n44), .Y(n14) );
  XOR2X4 U85 ( .A(n107), .B(n108), .Y(SUM[15]) );
  NAND2X1 U86 ( .A(B[1]), .B(A[1]), .Y(n72) );
  NAND2X2 U87 ( .A(B[2]), .B(A[2]), .Y(n58) );
  INVXL U88 ( .A(B[1]), .Y(n6) );
  XOR2X2 U89 ( .A(n71), .B(n73), .Y(SUM[1]) );
  NAND2X2 U90 ( .A(n142), .B(n143), .Y(n137) );
  OR2X4 U91 ( .A(A[10]), .B(B[10]), .Y(n143) );
  INVX2 U92 ( .A(n33), .Y(n32) );
  AND2X2 U93 ( .A(n55), .B(n56), .Y(n9) );
  OAI21X4 U94 ( .A0(n153), .A1(n154), .B0(n139), .Y(n152) );
  INVX8 U95 ( .A(n85), .Y(n97) );
  OR2X4 U96 ( .A(A[14]), .B(B[14]), .Y(n85) );
  OAI2BB1X2 U97 ( .A0N(n109), .A1N(n110), .B0(n111), .Y(n107) );
  OR2X2 U98 ( .A(A[9]), .B(B[9]), .Y(n10) );
  CLKINVX2 U99 ( .A(n53), .Y(n52) );
  NOR2BX4 U100 ( .AN(n1), .B(n37), .Y(n36) );
  NOR2X2 U101 ( .A(n115), .B(n97), .Y(n109) );
  NAND2X1 U102 ( .A(n120), .B(n119), .Y(n115) );
  OR2X2 U103 ( .A(A[8]), .B(B[8]), .Y(n11) );
  AOI31X2 U104 ( .A0(n2), .A1(n17), .A2(n125), .B0(n126), .Y(n124) );
  OAI2BB1X4 U105 ( .A0N(n8), .A1N(n9), .B0(n51), .Y(n39) );
  AND2X1 U106 ( .A(n57), .B(n58), .Y(n8) );
  NAND2X2 U107 ( .A(B[4]), .B(A[4]), .Y(n44) );
  AOI21X4 U108 ( .A0(n48), .A1(n41), .B0(n49), .Y(n47) );
  NAND2BX2 U109 ( .AN(n34), .B(n28), .Y(n33) );
  NAND2X2 U110 ( .A(n162), .B(n17), .Y(n177) );
  NAND3BX2 U111 ( .AN(n149), .B(n42), .C(B[5]), .Y(n144) );
  NAND4BX2 U112 ( .AN(n25), .B(n133), .C(n27), .D(n17), .Y(n132) );
  XOR2X2 U113 ( .A(n62), .B(n61), .Y(SUM[3]) );
  XOR2X4 U114 ( .A(n35), .B(n36), .Y(SUM[7]) );
  NAND3X2 U115 ( .A(n123), .B(n92), .C(n124), .Y(n121) );
  NAND2X2 U116 ( .A(n140), .B(n158), .Y(n157) );
  NAND2X2 U117 ( .A(n158), .B(n140), .Y(n173) );
  AOI21X2 U118 ( .A0(n159), .A1(n160), .B0(n161), .Y(n156) );
  AOI21X2 U119 ( .A0(n163), .A1(n164), .B0(n165), .Y(n159) );
  INVX4 U120 ( .A(n119), .Y(n91) );
  OR2X2 U121 ( .A(B[13]), .B(A[13]), .Y(n119) );
  OR2X1 U122 ( .A(A[3]), .B(B[3]), .Y(n54) );
  NAND4X2 U123 ( .A(n56), .B(n55), .C(n58), .D(n57), .Y(n104) );
  NOR2XL U124 ( .A(n91), .B(n98), .Y(n94) );
  NOR2BX2 U125 ( .AN(n90), .B(n91), .Y(n122) );
  XOR2X4 U126 ( .A(n50), .B(n14), .Y(SUM[5]) );
  XOR2X4 U127 ( .A(n47), .B(n46), .Y(SUM[6]) );
  NAND2X1 U128 ( .A(B[13]), .B(A[13]), .Y(n90) );
  OR2X4 U129 ( .A(A[2]), .B(B[2]), .Y(n69) );
  NAND2X4 U130 ( .A(B[12]), .B(A[12]), .Y(n92) );
  OAI21X2 U131 ( .A0(n98), .A1(n101), .B0(n127), .Y(n126) );
  OR2X4 U132 ( .A(A[7]), .B(B[7]), .Y(n17) );
  NAND2X4 U133 ( .A(n10), .B(n11), .Y(n171) );
  AND2X1 U134 ( .A(B[4]), .B(A[4]), .Y(n148) );
  NOR2X4 U135 ( .A(n134), .B(n63), .Y(n27) );
  OAI2BB1X1 U136 ( .A0N(n92), .A1N(n90), .B0(n119), .Y(n114) );
  INVXL U137 ( .A(n53), .Y(n60) );
  NAND2BX2 U138 ( .AN(n22), .B(n21), .Y(n158) );
  INVX4 U139 ( .A(n104), .Y(n134) );
  NOR2XL U140 ( .A(n96), .B(n97), .Y(n95) );
  AND2X2 U141 ( .A(n12), .B(n13), .Y(n19) );
  NOR2X1 U142 ( .A(n106), .B(n60), .Y(n12) );
  NOR2XL U143 ( .A(n34), .B(n105), .Y(n13) );
  INVX4 U144 ( .A(n120), .Y(n98) );
  NAND2XL U145 ( .A(n85), .B(n86), .Y(n83) );
  NAND2XL U146 ( .A(n89), .B(n90), .Y(n88) );
  INVX2 U147 ( .A(n67), .Y(n64) );
  AOI31X2 U148 ( .A0(n160), .A1(n175), .A2(n176), .B0(n177), .Y(n174) );
  NAND2XL U149 ( .A(n17), .B(n120), .Y(n128) );
  OR2X4 U150 ( .A(A[1]), .B(B[1]), .Y(n70) );
  XOR2X2 U151 ( .A(n76), .B(n77), .Y(SUM[16]) );
  OAI21X1 U152 ( .A0(n78), .A1(n79), .B0(n80), .Y(n76) );
  OR2XL U153 ( .A(A[15]), .B(B[15]), .Y(n86) );
  NOR2BX1 U154 ( .AN(n75), .B(n18), .Y(SUM[0]) );
  NOR2XL U155 ( .A(A[0]), .B(B[0]), .Y(n18) );
  INVX1 U156 ( .A(n114), .Y(n112) );
  NAND2X1 U157 ( .A(n94), .B(n95), .Y(n79) );
  NAND3BXL U158 ( .AN(n178), .B(n42), .C(n148), .Y(n175) );
  XOR2X4 U159 ( .A(n29), .B(n30), .Y(SUM[8]) );
  NAND2X1 U160 ( .A(n22), .B(n26), .Y(n30) );
  NAND2XL U161 ( .A(n42), .B(n1), .Y(n46) );
  NAND2X1 U162 ( .A(n43), .B(n41), .Y(n50) );
  NOR2X2 U163 ( .A(n173), .B(n174), .Y(n168) );
  NOR2XL U164 ( .A(n25), .B(n34), .Y(n31) );
  NOR2BX2 U165 ( .AN(n84), .B(n96), .Y(n108) );
  NOR2XL U166 ( .A(n91), .B(n92), .Y(n87) );
  NOR2X1 U167 ( .A(n87), .B(n88), .Y(n82) );
  INVXL U168 ( .A(n41), .Y(n106) );
  NOR2X1 U169 ( .A(n99), .B(n100), .Y(n78) );
  AOI21XL U170 ( .A0(n103), .A1(n33), .B0(n93), .Y(n99) );
  INVXL U171 ( .A(B[5]), .Y(n179) );
  NAND2XL U172 ( .A(n45), .B(n1), .Y(n165) );
  INVX1 U173 ( .A(n89), .Y(n113) );
  NAND2X2 U174 ( .A(n26), .B(n21), .Y(n150) );
  NAND2X1 U175 ( .A(B[3]), .B(A[3]), .Y(n56) );
  INVX1 U176 ( .A(A[5]), .Y(n149) );
  NAND2XL U177 ( .A(B[15]), .B(A[15]), .Y(n84) );
  XOR2X1 U178 ( .A(B[16]), .B(A[16]), .Y(n77) );
  INVX1 U179 ( .A(n81), .Y(n80) );
  OR2XL U180 ( .A(A[5]), .B(B[5]), .Y(n164) );
  NAND3X4 U181 ( .A(n53), .B(n42), .C(n20), .Y(n25) );
  AOI21X2 U182 ( .A0(n169), .A1(n31), .B0(n32), .Y(n29) );
  NAND2XL U183 ( .A(B[2]), .B(A[2]), .Y(n66) );
  NOR2XL U184 ( .A(A[5]), .B(B[5]), .Y(n178) );
  AND2X2 U185 ( .A(n43), .B(n44), .Y(n38) );
  CLKINVX3 U186 ( .A(n43), .Y(n49) );
  XOR2X4 U187 ( .A(n116), .B(n117), .Y(SUM[14]) );
  XOR2X4 U188 ( .A(n121), .B(n122), .Y(SUM[13]) );
  XOR2X4 U189 ( .A(n110), .B(n130), .Y(SUM[12]) );
  NAND2X4 U190 ( .A(n131), .B(n132), .Y(n110) );
  NAND2BX4 U191 ( .AN(n137), .B(n138), .Y(n101) );
  OR2X4 U192 ( .A(n150), .B(n151), .Y(n93) );
  XOR2X4 U193 ( .A(n152), .B(n16), .Y(SUM[11]) );
  XOR2X4 U194 ( .A(n166), .B(n167), .Y(SUM[10]) );
  OR2X4 U195 ( .A(A[4]), .B(B[4]), .Y(n53) );
  OR2X4 U196 ( .A(A[6]), .B(B[6]), .Y(n42) );
  OR2X4 U197 ( .A(A[9]), .B(B[9]), .Y(n21) );
endmodule


module butterfly_DW01_sub_68 ( A, B, DIFF );
  input [16:0] A;
  input [16:0] B;
  output [16:0] DIFF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213;

  AOI21X2 U3 ( .A0(n206), .A1(n3), .B0(n30), .Y(n202) );
  INVX8 U4 ( .A(n16), .Y(n30) );
  NAND2BX2 U5 ( .AN(B[4]), .B(A[4]), .Y(n3) );
  NAND2X1 U6 ( .A(n57), .B(n58), .Y(n56) );
  NAND2X4 U7 ( .A(n89), .B(n90), .Y(n57) );
  AND2X1 U8 ( .A(n119), .B(n130), .Y(n1) );
  INVX4 U9 ( .A(n130), .Y(n125) );
  NAND2BX4 U10 ( .AN(A[15]), .B(B[15]), .Y(n130) );
  INVX2 U11 ( .A(n28), .Y(n43) );
  NAND2X2 U12 ( .A(n162), .B(n163), .Y(n140) );
  NOR2X2 U13 ( .A(n168), .B(n169), .Y(n162) );
  NOR2X2 U14 ( .A(n29), .B(n30), .Y(n27) );
  NAND4BX2 U15 ( .AN(n78), .B(n166), .C(n80), .D(n81), .Y(n61) );
  NAND2BX2 U16 ( .AN(n97), .B(n96), .Y(n94) );
  INVX2 U17 ( .A(n23), .Y(n44) );
  NAND2X1 U18 ( .A(n90), .B(n60), .Y(n86) );
  NAND3X2 U19 ( .A(n109), .B(n32), .C(n183), .Y(n187) );
  NAND2BX1 U20 ( .AN(A[4]), .B(B[4]), .Y(n35) );
  NAND2X2 U21 ( .A(n60), .B(n59), .Y(n71) );
  OR2X2 U22 ( .A(B[9]), .B(n2), .Y(n40) );
  INVX1 U23 ( .A(A[9]), .Y(n2) );
  NAND2X2 U24 ( .A(n204), .B(n28), .Y(n22) );
  NAND2BX1 U25 ( .AN(B[15]), .B(A[15]), .Y(n119) );
  OAI21XL U26 ( .A0(n120), .A1(n121), .B0(n122), .Y(n117) );
  NAND2X2 U27 ( .A(n164), .B(n165), .Y(n58) );
  INVX4 U28 ( .A(n80), .Y(n77) );
  OAI21X2 U29 ( .A0(n92), .A1(n78), .B0(n93), .Y(n88) );
  CLKINVX3 U30 ( .A(n73), .Y(n89) );
  INVX1 U31 ( .A(n3), .Y(n84) );
  AOI21X2 U32 ( .A0(n199), .A1(n200), .B0(n201), .Y(n196) );
  NAND2BX1 U33 ( .AN(n182), .B(n15), .Y(n201) );
  AOI21X2 U34 ( .A0(n202), .A1(n203), .B0(n204), .Y(n200) );
  NOR2X1 U35 ( .A(n103), .B(n104), .Y(n99) );
  NAND2X1 U36 ( .A(n105), .B(n106), .Y(n104) );
  OAI2BB1X2 U37 ( .A0N(n171), .A1N(n153), .B0(n157), .Y(n102) );
  NOR2X1 U38 ( .A(n176), .B(n177), .Y(n171) );
  NAND2BX2 U39 ( .AN(A[0]), .B(B[0]), .Y(n97) );
  NAND2X1 U40 ( .A(n16), .B(n63), .Y(n62) );
  NOR2X1 U41 ( .A(n47), .B(n29), .Y(n46) );
  NOR2X1 U42 ( .A(n141), .B(n158), .Y(n152) );
  INVX1 U43 ( .A(A[5]), .Y(n189) );
  INVX4 U44 ( .A(n167), .Y(n78) );
  BUFX12 U45 ( .A(n37), .Y(n16) );
  NOR2X1 U46 ( .A(n77), .B(n78), .Y(n76) );
  AOI21X4 U47 ( .A0(n41), .A1(n144), .B0(n145), .Y(n143) );
  INVX2 U48 ( .A(n129), .Y(n120) );
  XOR2X4 U49 ( .A(n82), .B(n83), .Y(DIFF[5]) );
  NAND2BX2 U50 ( .AN(B[13]), .B(A[13]), .Y(n124) );
  NAND4BX2 U51 ( .AN(n43), .B(n39), .C(n157), .D(n170), .Y(n141) );
  AND2X2 U52 ( .A(n170), .B(n154), .Y(n7) );
  NAND2BXL U53 ( .AN(B[5]), .B(A[5]), .Y(n206) );
  NAND3XL U54 ( .A(n15), .B(n16), .C(n38), .Y(n33) );
  AOI21XL U55 ( .A0(n112), .A1(n61), .B0(n113), .Y(n107) );
  OAI21X2 U56 ( .A0(n48), .A1(n49), .B0(n50), .Y(n45) );
  AND3X1 U57 ( .A(n109), .B(n32), .C(n140), .Y(n14) );
  NAND3BX2 U58 ( .AN(n139), .B(n128), .C(n105), .Y(n133) );
  NAND2BX2 U59 ( .AN(A[6]), .B(B[6]), .Y(n37) );
  NAND2BX1 U60 ( .AN(A[10]), .B(B[10]), .Y(n170) );
  NAND2BXL U61 ( .AN(A[10]), .B(B[10]), .Y(n172) );
  INVX1 U62 ( .A(n31), .Y(n25) );
  NAND2BX1 U63 ( .AN(A[5]), .B(B[5]), .Y(n31) );
  INVX1 U64 ( .A(n97), .Y(n74) );
  NOR2X4 U65 ( .A(n70), .B(n71), .Y(n69) );
  NAND2BX4 U66 ( .AN(B[6]), .B(A[6]), .Y(n63) );
  NAND2XL U67 ( .A(n35), .B(n90), .Y(n169) );
  INVX1 U68 ( .A(n35), .Y(n190) );
  NAND2BX2 U69 ( .AN(B[8]), .B(A[8]), .Y(n23) );
  NAND3X4 U70 ( .A(n172), .B(n173), .C(n174), .Y(n153) );
  XOR2X4 U71 ( .A(n142), .B(n143), .Y(DIFF[14]) );
  INVX2 U72 ( .A(n111), .Y(n47) );
  INVX8 U73 ( .A(n32), .Y(n204) );
  NAND2BX4 U74 ( .AN(B[7]), .B(A[7]), .Y(n111) );
  NAND4BX1 U75 ( .AN(n25), .B(n27), .C(n26), .D(n28), .Y(n24) );
  NAND2BX2 U76 ( .AN(A[4]), .B(B[4]), .Y(n54) );
  NAND2BX4 U77 ( .AN(B[1]), .B(A[1]), .Y(n93) );
  NAND3X2 U78 ( .A(n67), .B(n68), .C(n69), .Y(n66) );
  XOR2X4 U79 ( .A(n11), .B(n12), .Y(DIFF[16]) );
  NAND2BX2 U80 ( .AN(A[8]), .B(B[8]), .Y(n28) );
  NAND2BX2 U81 ( .AN(B[11]), .B(A[11]), .Y(n155) );
  NAND2X2 U82 ( .A(n105), .B(n41), .Y(n161) );
  NAND2BX4 U83 ( .AN(A[9]), .B(B[9]), .Y(n39) );
  OAI21X1 U84 ( .A0(B[5]), .A1(n189), .B0(n4), .Y(n26) );
  NAND3X2 U85 ( .A(n22), .B(n23), .C(n24), .Y(n21) );
  INVX4 U86 ( .A(n15), .Y(n29) );
  NAND3BX4 U87 ( .AN(n207), .B(n208), .C(n209), .Y(n199) );
  INVX2 U88 ( .A(n63), .Y(n52) );
  INVX2 U89 ( .A(n53), .Y(n51) );
  OR2X1 U90 ( .A(n95), .B(n78), .Y(n8) );
  NAND2XL U91 ( .A(n128), .B(n121), .Y(n160) );
  NAND3X4 U92 ( .A(n121), .B(n154), .C(n155), .Y(n6) );
  XNOR2X4 U93 ( .A(n19), .B(n9), .Y(DIFF[4]) );
  NAND4BX4 U94 ( .AN(n85), .B(n58), .C(n61), .D(n60), .Y(n19) );
  NAND2X4 U95 ( .A(n63), .B(n111), .Y(n205) );
  NAND2BX4 U96 ( .AN(B[4]), .B(A[4]), .Y(n4) );
  NAND3X1 U97 ( .A(n59), .B(n60), .C(n61), .Y(n55) );
  NAND2X4 U98 ( .A(n156), .B(n121), .Y(n148) );
  OAI21X4 U99 ( .A0(n133), .A1(n14), .B0(n134), .Y(n132) );
  AOI21X2 U100 ( .A0(n135), .A1(n136), .B0(n137), .Y(n134) );
  OAI2BB1X2 U101 ( .A0N(A[9]), .A1N(n175), .B0(n23), .Y(n173) );
  AOI21X2 U102 ( .A0(n116), .A1(n117), .B0(n118), .Y(n115) );
  BUFX20 U103 ( .A(n36), .Y(n15) );
  NAND2BX4 U104 ( .AN(A[1]), .B(B[1]), .Y(n167) );
  NOR2X1 U105 ( .A(n138), .B(n139), .Y(n135) );
  NAND4BXL U106 ( .AN(n58), .B(n15), .C(n131), .D(n105), .Y(n114) );
  CLKINVX3 U107 ( .A(n141), .Y(n105) );
  XNOR2X2 U108 ( .A(n94), .B(n8), .Y(DIFF[1]) );
  AOI21X1 U109 ( .A0(n51), .A1(n16), .B0(n52), .Y(n50) );
  NAND3BX2 U110 ( .AN(n30), .B(n213), .C(n90), .Y(n207) );
  NAND2X1 U111 ( .A(n90), .B(n15), .Y(n194) );
  NAND2BX2 U112 ( .AN(A[3]), .B(B[3]), .Y(n90) );
  INVX2 U113 ( .A(n101), .Y(n106) );
  OAI21X2 U114 ( .A0(n114), .A1(n101), .B0(n115), .Y(n98) );
  NOR2XL U115 ( .A(n101), .B(n102), .Y(n100) );
  NAND4BX2 U116 ( .AN(n125), .B(n127), .C(n128), .D(n129), .Y(n101) );
  AOI21X4 U117 ( .A0(n152), .A1(n41), .B0(n13), .Y(n151) );
  AND2X2 U118 ( .A(n148), .B(n136), .Y(n13) );
  NAND2X2 U119 ( .A(n146), .B(n124), .Y(n145) );
  OAI21X4 U120 ( .A0(n179), .A1(n180), .B0(n154), .Y(n178) );
  NAND2X2 U121 ( .A(n181), .B(n172), .Y(n180) );
  NAND2BX2 U122 ( .AN(B[14]), .B(A[14]), .Y(n123) );
  NOR2X2 U123 ( .A(n77), .B(n78), .Y(n165) );
  AND2X4 U124 ( .A(n157), .B(n155), .Y(n5) );
  NAND2BX4 U125 ( .AN(A[11]), .B(B[11]), .Y(n157) );
  NAND2X4 U126 ( .A(n93), .B(n96), .Y(n81) );
  NAND2BX2 U127 ( .AN(B[10]), .B(A[10]), .Y(n154) );
  XOR2X4 U128 ( .A(n132), .B(n1), .Y(DIFF[15]) );
  NAND2XL U129 ( .A(n39), .B(n40), .Y(n17) );
  OAI21X1 U130 ( .A0(n126), .A1(n124), .B0(n123), .Y(n137) );
  AND2X2 U131 ( .A(n124), .B(n123), .Y(n122) );
  OR3X4 U132 ( .A(n98), .B(n99), .C(n100), .Y(n11) );
  NAND2BX4 U133 ( .AN(B[3]), .B(A[3]), .Y(n60) );
  NOR2X2 U134 ( .A(n120), .B(n138), .Y(n147) );
  NAND2BX4 U135 ( .AN(A[14]), .B(B[14]), .Y(n127) );
  AOI21X2 U136 ( .A0(n80), .A1(n88), .B0(n89), .Y(n87) );
  NAND2X2 U137 ( .A(n147), .B(n136), .Y(n146) );
  INVX4 U138 ( .A(n57), .Y(n85) );
  AOI31X2 U139 ( .A0(n184), .A1(n185), .A2(n186), .B0(n187), .Y(n179) );
  XOR2X4 U140 ( .A(n18), .B(n17), .Y(DIFF[9]) );
  AOI21X4 U141 ( .A0(n19), .A1(n20), .B0(n21), .Y(n18) );
  NAND2BX4 U142 ( .AN(A[7]), .B(B[7]), .Y(n36) );
  NAND2X1 U143 ( .A(n28), .B(n35), .Y(n34) );
  NAND2X2 U144 ( .A(n39), .B(n28), .Y(n182) );
  NAND2X1 U145 ( .A(n60), .B(n73), .Y(n191) );
  NAND2X1 U146 ( .A(n60), .B(n73), .Y(n210) );
  NAND2BX4 U147 ( .AN(B[2]), .B(A[2]), .Y(n73) );
  NOR2X1 U148 ( .A(n89), .B(n77), .Y(n91) );
  XNOR2X4 U149 ( .A(n10), .B(n62), .Y(DIFF[6]) );
  CLKINVX3 U150 ( .A(n148), .Y(n138) );
  NOR2XL U151 ( .A(n52), .B(n47), .Y(n110) );
  NAND2X2 U152 ( .A(n64), .B(n53), .Y(n10) );
  NAND3XL U153 ( .A(n54), .B(n16), .C(n38), .Y(n49) );
  NAND2X1 U154 ( .A(n129), .B(n127), .Y(n139) );
  INVXL U155 ( .A(n155), .Y(n177) );
  NAND2BX2 U156 ( .AN(n65), .B(n66), .Y(n64) );
  INVXL U157 ( .A(B[9]), .Y(n175) );
  NOR2XL U158 ( .A(n125), .B(n126), .Y(n116) );
  NAND2BX4 U159 ( .AN(n6), .B(n153), .Y(n136) );
  NOR2XL U160 ( .A(n43), .B(n44), .Y(n42) );
  XNOR2X4 U161 ( .A(n195), .B(n7), .Y(DIFF[10]) );
  OR2X2 U162 ( .A(n84), .B(n190), .Y(n9) );
  NOR2BXL U163 ( .AN(n60), .B(n85), .Y(n112) );
  XNOR2X1 U164 ( .A(B[16]), .B(A[16]), .Y(n12) );
  NAND2BXL U165 ( .AN(B[0]), .B(A[0]), .Y(n96) );
  XOR2X2 U166 ( .A(n88), .B(n91), .Y(DIFF[2]) );
  NAND2XL U167 ( .A(n109), .B(n110), .Y(n108) );
  INVX2 U168 ( .A(n183), .Y(n197) );
  INVX1 U169 ( .A(n113), .Y(n131) );
  NAND2X1 U170 ( .A(n16), .B(n15), .Y(n188) );
  NAND3BX1 U171 ( .AN(n191), .B(n192), .C(n193), .Y(n185) );
  NOR2X1 U172 ( .A(n30), .B(n194), .Y(n184) );
  NAND2XL U173 ( .A(n129), .B(n124), .Y(n150) );
  XNOR2X4 U174 ( .A(n159), .B(n160), .Y(DIFF[12]) );
  NOR2X2 U175 ( .A(n33), .B(n34), .Y(n20) );
  NAND2X1 U176 ( .A(n127), .B(n123), .Y(n142) );
  NOR2X1 U177 ( .A(n149), .B(n141), .Y(n144) );
  NAND2X2 U178 ( .A(n128), .B(n157), .Y(n156) );
  INVX1 U179 ( .A(n94), .Y(n92) );
  INVXL U180 ( .A(n93), .Y(n95) );
  NAND3XL U181 ( .A(n54), .B(n16), .C(n38), .Y(n113) );
  NAND2X2 U182 ( .A(n23), .B(n40), .Y(n198) );
  INVX1 U183 ( .A(n127), .Y(n126) );
  INVX1 U184 ( .A(n119), .Y(n118) );
  INVX1 U185 ( .A(n154), .Y(n176) );
  NAND3BXL U186 ( .AN(n74), .B(n167), .C(n80), .Y(n192) );
  XOR2X2 U187 ( .A(n86), .B(n87), .Y(DIFF[3]) );
  NAND2XL U188 ( .A(n38), .B(n53), .Y(n82) );
  AOI21X2 U189 ( .A0(n54), .A1(n19), .B0(n84), .Y(n83) );
  NOR2X2 U190 ( .A(n55), .B(n56), .Y(n48) );
  NAND3XL U191 ( .A(n167), .B(n80), .C(n81), .Y(n193) );
  NAND3BX2 U192 ( .AN(n210), .B(n211), .C(n212), .Y(n209) );
  NAND3BXL U193 ( .AN(n74), .B(n167), .C(n80), .Y(n211) );
  NAND3XL U194 ( .A(n167), .B(n80), .C(n81), .Y(n212) );
  INVXL U195 ( .A(n128), .Y(n158) );
  NAND2XL U196 ( .A(n129), .B(n128), .Y(n149) );
  NAND2X1 U197 ( .A(n182), .B(n183), .Y(n181) );
  NAND2XL U198 ( .A(n96), .B(n97), .Y(DIFF[0]) );
  AOI21XL U199 ( .A0(n72), .A1(B[3]), .B0(n73), .Y(n70) );
  INVXL U200 ( .A(A[3]), .Y(n72) );
  NAND4BXL U201 ( .AN(n78), .B(n79), .C(n80), .D(n81), .Y(n67) );
  NAND3BX1 U202 ( .AN(n74), .B(n75), .C(n76), .Y(n68) );
  NAND2BXL U203 ( .AN(A[4]), .B(B[4]), .Y(n213) );
  NAND2BX2 U204 ( .AN(A[5]), .B(B[5]), .Y(n38) );
  OAI21XL U205 ( .A0(n107), .A1(n108), .B0(n15), .Y(n103) );
  NAND3X1 U206 ( .A(n15), .B(n38), .C(n16), .Y(n168) );
  NAND2BXL U207 ( .AN(A[9]), .B(B[9]), .Y(n174) );
  NAND4BXL U208 ( .AN(n89), .B(n60), .C(n61), .D(n58), .Y(n163) );
  AOI21XL U209 ( .A0(B[5]), .A1(n189), .B0(n190), .Y(n186) );
  NAND2BXL U210 ( .AN(A[5]), .B(B[5]), .Y(n208) );
  NAND2BXL U211 ( .AN(A[5]), .B(B[5]), .Y(n203) );
  NAND2BX1 U212 ( .AN(B[5]), .B(A[5]), .Y(n53) );
  OAI2BB1X1 U213 ( .A0N(B[5]), .A1N(n189), .B0(n54), .Y(n65) );
  NAND2BXL U214 ( .AN(A[3]), .B(B[3]), .Y(n75) );
  NAND2BXL U215 ( .AN(A[3]), .B(B[3]), .Y(n79) );
  AOI21XL U216 ( .A0(n72), .A1(B[3]), .B0(n74), .Y(n164) );
  NAND2BXL U217 ( .AN(A[3]), .B(B[3]), .Y(n166) );
  XOR2X4 U218 ( .A(n41), .B(n42), .Y(DIFF[8]) );
  XOR2X4 U219 ( .A(n45), .B(n46), .Y(DIFF[7]) );
  XOR2X4 U220 ( .A(n150), .B(n151), .Y(DIFF[13]) );
  NAND2BX4 U221 ( .AN(A[13]), .B(B[13]), .Y(n129) );
  NAND2BX4 U222 ( .AN(B[12]), .B(A[12]), .Y(n121) );
  NAND2BX4 U223 ( .AN(A[12]), .B(B[12]), .Y(n128) );
  NAND2X4 U224 ( .A(n102), .B(n161), .Y(n159) );
  NAND3X4 U225 ( .A(n109), .B(n32), .C(n140), .Y(n41) );
  XOR2X4 U226 ( .A(n178), .B(n5), .Y(DIFF[11]) );
  NAND3BX4 U227 ( .AN(n188), .B(n31), .C(n26), .Y(n109) );
  NOR2X4 U228 ( .A(n196), .B(n197), .Y(n195) );
  NAND2X4 U229 ( .A(n198), .B(n39), .Y(n183) );
  NAND2X4 U230 ( .A(n205), .B(n15), .Y(n32) );
  NAND2BX4 U231 ( .AN(B[4]), .B(A[4]), .Y(n59) );
  NAND2BX4 U232 ( .AN(A[2]), .B(B[2]), .Y(n80) );
endmodule


module butterfly_DW01_add_94 ( A, B, SUM );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201;

  CLKINVX3 U2 ( .A(n106), .Y(n127) );
  NAND2X1 U3 ( .A(A[5]), .B(B[5]), .Y(n19) );
  NAND3BX4 U4 ( .AN(n10), .B(n182), .C(n183), .Y(n171) );
  CLKINVX8 U5 ( .A(n28), .Y(n166) );
  BUFX8 U6 ( .A(n163), .Y(n1) );
  NOR2X2 U7 ( .A(n135), .B(n136), .Y(n131) );
  INVX8 U8 ( .A(n117), .Y(n135) );
  NAND2X4 U9 ( .A(B[8]), .B(A[8]), .Y(n36) );
  NOR2X4 U10 ( .A(n167), .B(n168), .Y(n164) );
  OR2X4 U11 ( .A(A[11]), .B(B[11]), .Y(n113) );
  INVX1 U12 ( .A(n1), .Y(n181) );
  OAI21X2 U13 ( .A0(n161), .A1(n162), .B0(n1), .Y(n157) );
  INVX3 U14 ( .A(n15), .Y(n59) );
  NOR2X2 U15 ( .A(n19), .B(n20), .Y(n170) );
  INVX4 U16 ( .A(n174), .Y(n71) );
  CLKINVX3 U17 ( .A(n34), .Y(n29) );
  INVX1 U18 ( .A(A[4]), .Y(n56) );
  CLKINVX3 U19 ( .A(n169), .Y(n167) );
  OR2X2 U20 ( .A(A[2]), .B(B[2]), .Y(n194) );
  NAND2X2 U21 ( .A(n42), .B(n36), .Y(n31) );
  INVX1 U22 ( .A(n109), .Y(n151) );
  OAI21XL U23 ( .A0(n108), .A1(n109), .B0(n110), .Y(n107) );
  AND2X2 U24 ( .A(n137), .B(n115), .Y(n22) );
  INVX1 U25 ( .A(n110), .Y(n14) );
  OR2X2 U26 ( .A(A[14]), .B(B[14]), .Y(n105) );
  CLKINVX3 U27 ( .A(n195), .Y(n82) );
  BUFX3 U28 ( .A(n77), .Y(n15) );
  INVX4 U29 ( .A(n194), .Y(n84) );
  OAI21X2 U30 ( .A0(n43), .A1(n44), .B0(n45), .Y(n39) );
  NOR2X1 U31 ( .A(n52), .B(n53), .Y(n43) );
  NAND2X1 U32 ( .A(B[10]), .B(A[10]), .Y(n163) );
  CLKINVX3 U33 ( .A(n115), .Y(n146) );
  INVX4 U34 ( .A(n38), .Y(n150) );
  CLKINVX3 U35 ( .A(n113), .Y(n156) );
  NAND2X2 U36 ( .A(B[12]), .B(A[12]), .Y(n109) );
  NAND2X2 U37 ( .A(n120), .B(n6), .Y(n37) );
  NAND3X2 U38 ( .A(n31), .B(n32), .C(n33), .Y(n30) );
  XOR2X1 U39 ( .A(n89), .B(n91), .Y(SUM[1]) );
  NOR2X1 U40 ( .A(n75), .B(n76), .Y(n72) );
  AND2X2 U41 ( .A(n68), .B(n55), .Y(n24) );
  INVX4 U42 ( .A(n121), .Y(n42) );
  AND2X2 U43 ( .A(n188), .B(n189), .Y(n2) );
  NAND4BBX4 U44 ( .AN(n3), .BN(n170), .C(n171), .D(n36), .Y(n33) );
  NAND2X1 U45 ( .A(n41), .B(n49), .Y(n3) );
  AOI2BB2X2 U46 ( .B0(B[11]), .B1(A[11]), .A0N(n159), .A1N(n160), .Y(n158) );
  NOR2XL U47 ( .A(A[10]), .B(B[10]), .Y(n159) );
  NAND2XL U48 ( .A(A[9]), .B(B[9]), .Y(n160) );
  NAND2X2 U49 ( .A(B[9]), .B(A[9]), .Y(n27) );
  NOR2XL U50 ( .A(n170), .B(n198), .Y(n190) );
  NAND2X2 U51 ( .A(n137), .B(n21), .Y(n136) );
  NAND2X1 U52 ( .A(n174), .B(n121), .Y(n185) );
  NAND2XL U53 ( .A(n110), .B(n138), .Y(n147) );
  NAND2BXL U54 ( .AN(n109), .B(n138), .Y(n143) );
  CLKINVX4 U55 ( .A(n138), .Y(n108) );
  OAI21X4 U56 ( .A0(n4), .A1(n5), .B0(n27), .Y(n187) );
  OR2X2 U57 ( .A(n199), .B(n200), .Y(n4) );
  AND3X4 U58 ( .A(n2), .B(n190), .C(n191), .Y(n5) );
  NAND4BX4 U59 ( .AN(n185), .B(n32), .C(n186), .D(n78), .Y(n34) );
  XOR2X4 U60 ( .A(n78), .B(n79), .Y(SUM[4]) );
  NAND3BX2 U61 ( .AN(n185), .B(n186), .C(n78), .Y(n191) );
  NAND2BX2 U62 ( .AN(n59), .B(n60), .Y(n75) );
  OR2X2 U63 ( .A(n11), .B(n12), .Y(n61) );
  NOR2X2 U64 ( .A(n63), .B(n51), .Y(n11) );
  AND2X2 U65 ( .A(n1), .B(n169), .Y(n18) );
  NAND2BX1 U66 ( .AN(n27), .B(n169), .Y(n178) );
  NAND2X1 U67 ( .A(n22), .B(n99), .Y(n128) );
  NAND2BX1 U68 ( .AN(n51), .B(n50), .Y(n44) );
  NAND4X1 U69 ( .A(n9), .B(A[4]), .C(n183), .D(n182), .Y(n189) );
  OR2X2 U70 ( .A(A[5]), .B(B[5]), .Y(n182) );
  NOR2XL U71 ( .A(A[6]), .B(B[6]), .Y(n20) );
  OR2X2 U72 ( .A(A[6]), .B(B[6]), .Y(n183) );
  NOR2X2 U73 ( .A(n65), .B(n66), .Y(n63) );
  NAND2BX2 U74 ( .AN(n59), .B(n60), .Y(n65) );
  NAND2X1 U75 ( .A(n27), .B(n28), .Y(n26) );
  OAI21X1 U76 ( .A0(A[5]), .A1(B[5]), .B0(n64), .Y(n51) );
  INVX3 U77 ( .A(n50), .Y(n46) );
  OR2XL U78 ( .A(A[6]), .B(B[6]), .Y(n50) );
  CLKINVX3 U79 ( .A(n42), .Y(n6) );
  NAND2X2 U80 ( .A(B[7]), .B(A[7]), .Y(n41) );
  NAND2X1 U81 ( .A(A[4]), .B(n9), .Y(n10) );
  NAND2X2 U82 ( .A(n37), .B(n38), .Y(n35) );
  NOR2BX4 U83 ( .AN(n74), .B(n73), .Y(n79) );
  OAI21X2 U84 ( .A0(n72), .A1(n73), .B0(n74), .Y(n69) );
  AOI2BB1X4 U85 ( .A0N(n56), .A1N(n57), .B0(n58), .Y(n67) );
  AND2X4 U86 ( .A(n64), .B(n183), .Y(n172) );
  NOR2XL U87 ( .A(A[6]), .B(B[6]), .Y(n23) );
  OAI21X2 U88 ( .A0(n109), .A1(n133), .B0(n134), .Y(n132) );
  AOI21XL U89 ( .A0(n118), .A1(n37), .B0(n119), .Y(n116) );
  INVX8 U90 ( .A(n119), .Y(n99) );
  NAND2XL U91 ( .A(n169), .B(n28), .Y(n177) );
  OAI21X4 U92 ( .A0(A[14]), .A1(B[14]), .B0(n138), .Y(n133) );
  NAND2BX2 U93 ( .AN(n23), .B(n64), .Y(n197) );
  NAND2X1 U94 ( .A(B[5]), .B(A[5]), .Y(n47) );
  AOI2BB1X2 U95 ( .A0N(n46), .A1N(n47), .B0(n48), .Y(n45) );
  AOI21X4 U96 ( .A0(n120), .A1(n6), .B0(n150), .Y(n129) );
  OAI21XL U97 ( .A0(n122), .A1(n123), .B0(n124), .Y(n118) );
  OAI21X4 U98 ( .A0(n128), .A1(n7), .B0(n130), .Y(n125) );
  BUFX1 U99 ( .A(n129), .Y(n7) );
  NOR2X2 U100 ( .A(n131), .B(n132), .Y(n130) );
  OR2X1 U101 ( .A(A[15]), .B(B[15]), .Y(n106) );
  OR2X4 U102 ( .A(A[5]), .B(B[5]), .Y(n174) );
  XOR2X4 U103 ( .A(n39), .B(n40), .Y(SUM[7]) );
  NAND2X1 U104 ( .A(B[14]), .B(A[14]), .Y(n111) );
  NOR2X4 U105 ( .A(n42), .B(n71), .Y(n173) );
  INVX4 U106 ( .A(n197), .Y(n186) );
  AOI21X4 U107 ( .A0(n180), .A1(n33), .B0(n181), .Y(n179) );
  NAND2X4 U108 ( .A(n173), .B(n172), .Y(n112) );
  NAND2X2 U109 ( .A(B[13]), .B(A[13]), .Y(n110) );
  NAND2X4 U110 ( .A(n99), .B(n145), .Y(n144) );
  NAND2X1 U111 ( .A(n21), .B(n138), .Y(n142) );
  NAND3X4 U112 ( .A(A[2]), .B(B[2]), .C(n195), .Y(n68) );
  NOR2X4 U113 ( .A(n129), .B(n144), .Y(n13) );
  NAND2XL U114 ( .A(n41), .B(n49), .Y(n198) );
  OAI22X1 U115 ( .A0(A[9]), .A1(B[9]), .B0(A[10]), .B1(B[10]), .Y(n161) );
  NOR2BX1 U116 ( .AN(n109), .B(n146), .Y(n153) );
  OAI21X2 U117 ( .A0(n83), .A1(n84), .B0(n85), .Y(n80) );
  NOR2BX2 U118 ( .AN(n49), .B(n46), .Y(n62) );
  INVX4 U119 ( .A(n57), .Y(n9) );
  NAND3BX2 U120 ( .AN(n129), .B(n115), .C(n99), .Y(n149) );
  NOR2BX4 U121 ( .AN(n8), .B(n141), .Y(n140) );
  NOR2X4 U122 ( .A(n13), .B(n14), .Y(n8) );
  INVX3 U123 ( .A(B[4]), .Y(n57) );
  NOR2BX1 U124 ( .AN(n90), .B(n92), .Y(n91) );
  NAND2X1 U125 ( .A(n105), .B(n111), .Y(n139) );
  AND2X4 U126 ( .A(n115), .B(n113), .Y(n21) );
  NAND2X4 U127 ( .A(n28), .B(n32), .Y(n199) );
  NAND2XL U128 ( .A(n32), .B(n36), .Y(n16) );
  NOR2BX2 U129 ( .AN(n47), .B(n71), .Y(n70) );
  NOR2BX1 U130 ( .AN(n41), .B(n42), .Y(n40) );
  NAND2X2 U131 ( .A(n99), .B(n6), .Y(n155) );
  NAND2X2 U132 ( .A(n67), .B(n55), .Y(n66) );
  NOR2X4 U133 ( .A(n184), .B(n199), .Y(n180) );
  NAND2X2 U134 ( .A(n31), .B(n169), .Y(n184) );
  NOR2X2 U135 ( .A(n150), .B(n120), .Y(n154) );
  NAND4BX4 U136 ( .AN(n170), .B(n49), .C(n41), .D(n171), .Y(n120) );
  NOR2BX4 U137 ( .AN(n32), .B(n166), .Y(n165) );
  NAND3X4 U138 ( .A(n194), .B(n195), .C(n196), .Y(n55) );
  NOR2X2 U139 ( .A(A[11]), .B(B[11]), .Y(n168) );
  OAI2BB1X1 U140 ( .A0N(n110), .A1N(n111), .B0(n105), .Y(n134) );
  NAND2BX4 U141 ( .AN(n29), .B(n30), .Y(n25) );
  OAI22X4 U142 ( .A0(n155), .A1(n154), .B0(n156), .B1(n135), .Y(n152) );
  NAND2XL U143 ( .A(n68), .B(n55), .Y(n76) );
  INVX4 U144 ( .A(n68), .Y(n58) );
  OAI21X2 U145 ( .A0(n135), .A1(n142), .B0(n143), .Y(n141) );
  XOR2X2 U146 ( .A(n80), .B(n81), .Y(SUM[3]) );
  XNOR2X4 U147 ( .A(n25), .B(n26), .Y(SUM[9]) );
  INVX4 U148 ( .A(n133), .Y(n137) );
  NAND2X2 U149 ( .A(B[6]), .B(A[6]), .Y(n49) );
  AOI2BB1X1 U150 ( .A0N(n56), .A1N(n57), .B0(n58), .Y(n54) );
  NOR2X2 U151 ( .A(n108), .B(n146), .Y(n145) );
  OR2X4 U152 ( .A(A[8]), .B(B[8]), .Y(n32) );
  OR2X4 U153 ( .A(A[12]), .B(B[12]), .Y(n115) );
  XOR2X4 U154 ( .A(n125), .B(n126), .Y(SUM[15]) );
  XOR2X4 U155 ( .A(n175), .B(n176), .Y(SUM[11]) );
  OR2X4 U156 ( .A(A[9]), .B(B[9]), .Y(n28) );
  OR2X4 U157 ( .A(A[10]), .B(B[10]), .Y(n169) );
  XOR2X2 U158 ( .A(n86), .B(n87), .Y(SUM[2]) );
  NOR2BX2 U159 ( .AN(n85), .B(n84), .Y(n87) );
  INVX4 U160 ( .A(n64), .Y(n73) );
  OR2X4 U161 ( .A(A[7]), .B(B[7]), .Y(n121) );
  INVXL U162 ( .A(n47), .Y(n12) );
  XOR2X4 U163 ( .A(n61), .B(n62), .Y(SUM[6]) );
  XOR2X4 U164 ( .A(n69), .B(n70), .Y(SUM[5]) );
  NAND2X1 U165 ( .A(n9), .B(A[4]), .Y(n74) );
  OR2X4 U166 ( .A(A[4]), .B(B[4]), .Y(n64) );
  NAND2X1 U167 ( .A(n54), .B(n55), .Y(n53) );
  NAND2XL U168 ( .A(B[3]), .B(A[3]), .Y(n77) );
  INVX2 U169 ( .A(n86), .Y(n83) );
  INVXL U170 ( .A(n112), .Y(n124) );
  OR2X4 U171 ( .A(A[13]), .B(B[13]), .Y(n138) );
  XNOR2X4 U172 ( .A(n35), .B(n16), .Y(SUM[8]) );
  XNOR2X4 U173 ( .A(n17), .B(n147), .Y(SUM[13]) );
  NAND2X2 U174 ( .A(n148), .B(n149), .Y(n17) );
  NAND2BX4 U175 ( .AN(n112), .B(n78), .Y(n38) );
  NOR2BX1 U176 ( .AN(n111), .B(n107), .Y(n102) );
  INVXL U177 ( .A(n49), .Y(n48) );
  NOR2BXL U178 ( .AN(n15), .B(n82), .Y(n81) );
  OAI21X2 U179 ( .A0(n96), .A1(n97), .B0(n98), .Y(n94) );
  NOR2XL U180 ( .A(n116), .B(n117), .Y(n96) );
  NAND2X1 U181 ( .A(n100), .B(n113), .Y(n97) );
  INVX1 U182 ( .A(n101), .Y(n98) );
  AOI21X1 U183 ( .A0(n21), .A1(n117), .B0(n151), .Y(n148) );
  NOR2BX2 U184 ( .AN(n104), .B(n127), .Y(n126) );
  OAI21X1 U185 ( .A0(n102), .A1(n103), .B0(n104), .Y(n101) );
  NAND2XL U186 ( .A(n105), .B(n106), .Y(n103) );
  NAND4BXL U187 ( .AN(n108), .B(n115), .C(n105), .D(n106), .Y(n114) );
  NAND3X4 U188 ( .A(n24), .B(n60), .C(n15), .Y(n78) );
  OAI2BB1X1 U189 ( .A0N(n88), .A1N(n89), .B0(n90), .Y(n86) );
  NAND2XL U190 ( .A(n68), .B(n55), .Y(n123) );
  NAND2XL U191 ( .A(n60), .B(n15), .Y(n122) );
  NAND2XL U192 ( .A(B[15]), .B(A[15]), .Y(n104) );
  NAND2BXL U193 ( .AN(n59), .B(n60), .Y(n52) );
  XOR2X1 U194 ( .A(B[16]), .B(A[16]), .Y(n95) );
  INVX1 U195 ( .A(n93), .Y(n89) );
  AND2X2 U196 ( .A(n93), .B(n201), .Y(SUM[0]) );
  OR2X2 U197 ( .A(A[0]), .B(B[0]), .Y(n201) );
  NAND2X1 U198 ( .A(B[0]), .B(A[0]), .Y(n93) );
  NAND2XL U199 ( .A(B[1]), .B(A[1]), .Y(n90) );
  AND2X1 U200 ( .A(B[1]), .B(A[1]), .Y(n196) );
  OR2X2 U201 ( .A(A[1]), .B(B[1]), .Y(n88) );
  AOI21X2 U202 ( .A0(B[11]), .A1(A[11]), .B0(n156), .Y(n176) );
  NAND2XL U203 ( .A(B[2]), .B(A[2]), .Y(n85) );
  NAND2XL U204 ( .A(A[8]), .B(B[8]), .Y(n188) );
  AOI21XL U205 ( .A0(B[8]), .A1(A[8]), .B0(n121), .Y(n200) );
  NAND2XL U206 ( .A(B[8]), .B(A[8]), .Y(n162) );
  XOR2X4 U207 ( .A(n94), .B(n95), .Y(SUM[16]) );
  CLKINVX3 U208 ( .A(n114), .Y(n100) );
  XOR2X4 U209 ( .A(n140), .B(n139), .Y(SUM[14]) );
  XOR2X4 U210 ( .A(n152), .B(n153), .Y(SUM[12]) );
  NAND2BX4 U211 ( .AN(n157), .B(n158), .Y(n117) );
  NAND2X4 U212 ( .A(n164), .B(n165), .Y(n119) );
  OAI211X2 U213 ( .A0(n34), .A1(n177), .B0(n179), .C0(n178), .Y(n175) );
  XOR2X4 U214 ( .A(n187), .B(n18), .Y(SUM[10]) );
  NAND2X4 U215 ( .A(n192), .B(n193), .Y(n60) );
  NOR2X4 U216 ( .A(n82), .B(n84), .Y(n193) );
  NOR2X4 U217 ( .A(n92), .B(n93), .Y(n192) );
  CLKINVX3 U218 ( .A(n88), .Y(n92) );
  OR2X4 U219 ( .A(A[3]), .B(B[3]), .Y(n195) );
endmodule


module butterfly_DW01_sub_69 ( A, B, DIFF );
  input [16:0] A;
  input [16:0] B;
  output [16:0] DIFF;
  wire   n181, n1, n2, n3, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180;

  INVX3 U3 ( .A(n93), .Y(n79) );
  AOI21X4 U4 ( .A0(n99), .A1(n128), .B0(n129), .Y(n126) );
  NAND2X4 U5 ( .A(n1), .B(n152), .Y(n135) );
  AND3X4 U6 ( .A(n39), .B(n110), .C(n114), .Y(n1) );
  XOR2X2 U7 ( .A(n45), .B(n3), .Y(n2) );
  CLKINVX20 U8 ( .A(n2), .Y(DIFF[5]) );
  OR2X2 U9 ( .A(n46), .B(n43), .Y(n3) );
  AOI21X4 U10 ( .A0(n32), .A1(n30), .B0(n175), .Y(n168) );
  NOR2X4 U11 ( .A(n79), .B(n80), .Y(n77) );
  CLKINVX8 U12 ( .A(n35), .Y(n41) );
  AOI21X4 U13 ( .A0(n111), .A1(n112), .B0(n113), .Y(n104) );
  INVX2 U14 ( .A(n114), .Y(n113) );
  AOI21X2 U15 ( .A0(n115), .A1(n116), .B0(n41), .Y(n112) );
  AOI21X2 U16 ( .A0(n104), .A1(n105), .B0(n106), .Y(n95) );
  NOR2BX4 U17 ( .AN(n9), .B(n98), .Y(n97) );
  CLKBUFX8 U18 ( .A(n181), .Y(DIFF[3]) );
  INVX4 U19 ( .A(n49), .Y(n51) );
  NAND2BX1 U20 ( .AN(A[1]), .B(B[1]), .Y(n68) );
  NAND3BX2 U21 ( .AN(n161), .B(n29), .C(n28), .Y(n169) );
  INVX1 U22 ( .A(n31), .Y(n175) );
  XOR2X2 U23 ( .A(n26), .B(n27), .Y(DIFF[8]) );
  XOR2X1 U24 ( .A(n53), .B(n54), .Y(n181) );
  XOR2X1 U25 ( .A(n29), .B(n50), .Y(DIFF[4]) );
  OR2X2 U26 ( .A(n24), .B(n25), .Y(n5) );
  AND2X4 U27 ( .A(n108), .B(n32), .Y(n6) );
  INVX4 U28 ( .A(n109), .Y(n25) );
  AOI21XL U29 ( .A0(n28), .A1(n29), .B0(n30), .Y(n156) );
  NAND2X2 U30 ( .A(n29), .B(n49), .Y(n47) );
  CLKINVX3 U31 ( .A(n170), .Y(n28) );
  NAND4BX2 U32 ( .AN(n41), .B(n117), .C(n108), .D(n49), .Y(n170) );
  NAND3XL U33 ( .A(n150), .B(n151), .C(n135), .Y(n149) );
  NAND2BX2 U34 ( .AN(B[6]), .B(A[6]), .Y(n180) );
  NOR2X1 U35 ( .A(n165), .B(n25), .Y(n163) );
  NAND2X2 U36 ( .A(n58), .B(n55), .Y(n171) );
  AND2X1 U37 ( .A(n21), .B(n100), .Y(n157) );
  NAND3X1 U38 ( .A(n99), .B(n92), .C(n81), .Y(n98) );
  XNOR2X4 U39 ( .A(n20), .B(n7), .Y(DIFF[13]) );
  AND2X1 U40 ( .A(n86), .B(n82), .Y(n7) );
  AND2X2 U41 ( .A(n86), .B(n93), .Y(n9) );
  CLKINVX2 U42 ( .A(n86), .Y(n85) );
  NAND2BX4 U43 ( .AN(A[7]), .B(B[7]), .Y(n38) );
  NOR2BX4 U44 ( .AN(B[7]), .B(A[7]), .Y(n179) );
  NAND2BX2 U45 ( .AN(B[15]), .B(A[15]), .Y(n120) );
  NAND3X1 U46 ( .A(n102), .B(n103), .C(n100), .Y(n153) );
  INVX4 U47 ( .A(n102), .Y(n129) );
  NAND2XL U48 ( .A(n92), .B(n86), .Y(n141) );
  AOI21X2 U49 ( .A0(n125), .A1(n126), .B0(n127), .Y(n123) );
  NAND2X2 U50 ( .A(n82), .B(n83), .Y(n124) );
  INVX1 U51 ( .A(n130), .Y(n128) );
  NAND2BX2 U52 ( .AN(n130), .B(n147), .Y(n146) );
  NAND2XL U53 ( .A(n86), .B(n81), .Y(n122) );
  NOR2X2 U54 ( .A(n79), .B(n78), .Y(n119) );
  NAND3X4 U55 ( .A(n82), .B(n83), .C(n84), .Y(n76) );
  INVX3 U56 ( .A(A[9]), .Y(n159) );
  NAND2BXL U57 ( .AN(B[9]), .B(A[9]), .Y(n166) );
  NOR2X4 U58 ( .A(n25), .B(n127), .Y(n134) );
  NOR2X2 U59 ( .A(n25), .B(n127), .Y(n151) );
  NOR2X4 U60 ( .A(n178), .B(n179), .Y(n177) );
  NAND3BX2 U61 ( .AN(n145), .B(n146), .C(n100), .Y(n142) );
  NAND2BX1 U62 ( .AN(A[1]), .B(B[1]), .Y(n172) );
  OAI21X2 U63 ( .A0(n62), .A1(n63), .B0(n64), .Y(n56) );
  NAND2X2 U64 ( .A(n92), .B(n153), .Y(n148) );
  INVX1 U65 ( .A(n107), .Y(n165) );
  INVX8 U66 ( .A(n92), .Y(n127) );
  XNOR2X4 U67 ( .A(n71), .B(n8), .Y(DIFF[16]) );
  XOR2X4 U68 ( .A(B[16]), .B(A[16]), .Y(n8) );
  NAND2BX2 U69 ( .AN(B[8]), .B(A[8]), .Y(n31) );
  XNOR2X4 U70 ( .A(n154), .B(n155), .Y(DIFF[12]) );
  NAND2X2 U71 ( .A(n35), .B(n36), .Y(n15) );
  NOR2BX2 U72 ( .AN(B[5]), .B(A[5]), .Y(n178) );
  NAND2X4 U73 ( .A(n35), .B(n176), .Y(n17) );
  BUFX2 U74 ( .A(A[14]), .Y(n10) );
  NAND3X2 U75 ( .A(n39), .B(n114), .C(n110), .Y(n30) );
  AND2X2 U76 ( .A(n39), .B(n110), .Y(n105) );
  NOR2X4 U77 ( .A(n136), .B(n137), .Y(n133) );
  NAND4BX2 U78 ( .AN(n131), .B(n147), .C(n132), .D(n107), .Y(n125) );
  DLY1X1 U79 ( .A(n44), .Y(n14) );
  NOR2X2 U80 ( .A(n136), .B(n137), .Y(n150) );
  NOR2X2 U81 ( .A(n43), .B(n51), .Y(n111) );
  NAND2X2 U82 ( .A(n100), .B(n101), .Y(n96) );
  NAND2X2 U83 ( .A(n92), .B(n86), .Y(n91) );
  INVX4 U84 ( .A(n99), .Y(n136) );
  NAND4BX4 U85 ( .AN(n87), .B(n28), .C(n88), .D(n89), .Y(n73) );
  NOR2X4 U86 ( .A(n90), .B(n91), .Y(n89) );
  NAND4X2 U87 ( .A(n107), .B(n32), .C(n108), .D(n109), .Y(n106) );
  BUFX1 U88 ( .A(n84), .Y(n11) );
  CLKINVX3 U89 ( .A(n81), .Y(n80) );
  NAND2XL U90 ( .A(n84), .B(n81), .Y(n139) );
  AOI21X4 U91 ( .A0(n163), .A1(n23), .B0(n164), .Y(n162) );
  XNOR2X4 U92 ( .A(n12), .B(n162), .Y(DIFF[11]) );
  AND2X1 U93 ( .A(n102), .B(n158), .Y(n12) );
  XNOR2X4 U94 ( .A(n167), .B(n13), .Y(DIFF[10]) );
  AND2X1 U95 ( .A(n107), .B(n130), .Y(n13) );
  AND2X1 U96 ( .A(n146), .B(n102), .Y(n21) );
  NAND4BX2 U97 ( .AN(n41), .B(n117), .C(n49), .D(n29), .Y(n152) );
  NAND2BX2 U98 ( .AN(A[11]), .B(B[11]), .Y(n158) );
  NAND4BX2 U99 ( .AN(n161), .B(n109), .C(n99), .D(n107), .Y(n87) );
  AOI21X2 U100 ( .A0(n23), .A1(n109), .B0(n24), .Y(n167) );
  CLKINVX8 U101 ( .A(n160), .Y(n131) );
  NAND2X2 U102 ( .A(n85), .B(n84), .Y(n75) );
  AND2X4 U103 ( .A(n102), .B(n103), .Y(n101) );
  NAND2X1 U104 ( .A(n102), .B(n83), .Y(n145) );
  NAND2BX4 U105 ( .AN(A[11]), .B(B[11]), .Y(n147) );
  NOR3X4 U106 ( .A(n19), .B(n123), .C(n124), .Y(n121) );
  AND3X4 U107 ( .A(n133), .B(n134), .C(n135), .Y(n19) );
  NAND2BX4 U108 ( .AN(A[11]), .B(B[11]), .Y(n99) );
  NAND3X4 U109 ( .A(n72), .B(n73), .C(n74), .Y(n71) );
  NAND2BX4 U110 ( .AN(A[9]), .B(B[9]), .Y(n160) );
  NOR2BX1 U111 ( .AN(n59), .B(n22), .Y(n115) );
  NAND2BX4 U112 ( .AN(B[3]), .B(A[3]), .Y(n59) );
  INVX4 U113 ( .A(n180), .Y(n37) );
  NAND2X4 U114 ( .A(n6), .B(n107), .Y(n137) );
  NAND2X2 U115 ( .A(n81), .B(n93), .Y(n90) );
  OAI21X4 U116 ( .A0(n42), .A1(n43), .B0(n14), .Y(n36) );
  INVX4 U117 ( .A(n45), .Y(n42) );
  XOR2X4 U118 ( .A(n36), .B(n40), .Y(DIFF[6]) );
  AND3X4 U119 ( .A(n148), .B(n83), .C(n149), .Y(n20) );
  NAND2BX4 U120 ( .AN(A[5]), .B(B[5]), .Y(n117) );
  OAI21X2 U121 ( .A0(n156), .A1(n87), .B0(n157), .Y(n154) );
  NAND4BX2 U122 ( .AN(n137), .B(n135), .C(n109), .D(n99), .Y(n144) );
  NAND4X2 U123 ( .A(n55), .B(n68), .C(n58), .D(n70), .Y(n94) );
  AND2X4 U124 ( .A(n15), .B(n180), .Y(n34) );
  NAND2BX4 U125 ( .AN(A[6]), .B(B[6]), .Y(n35) );
  OR2X4 U126 ( .A(n96), .B(n95), .Y(n16) );
  NAND2X4 U127 ( .A(n16), .B(n97), .Y(n72) );
  NAND2BX4 U128 ( .AN(A[4]), .B(B[4]), .Y(n49) );
  OAI21X4 U129 ( .A0(B[9]), .A1(n159), .B0(n31), .Y(n132) );
  AOI21X1 U130 ( .A0(n28), .A1(n29), .B0(n30), .Y(n27) );
  OAI21X4 U131 ( .A0(n121), .A1(n122), .B0(n11), .Y(n118) );
  NAND2BX4 U132 ( .AN(A[7]), .B(B[7]), .Y(n108) );
  NAND2X4 U133 ( .A(n18), .B(n177), .Y(n110) );
  INVX4 U134 ( .A(n17), .Y(n18) );
  NAND2X4 U135 ( .A(n44), .B(n48), .Y(n176) );
  AND2X2 U136 ( .A(n57), .B(n58), .Y(n22) );
  OAI21X1 U137 ( .A0(n165), .A1(n166), .B0(n130), .Y(n164) );
  AOI31X2 U138 ( .A0(n75), .A1(n76), .A2(n77), .B0(n78), .Y(n74) );
  XNOR2X4 U139 ( .A(n23), .B(n5), .Y(DIFF[9]) );
  NAND2BX4 U140 ( .AN(A[9]), .B(B[9]), .Y(n109) );
  NAND2BX4 U141 ( .AN(B[13]), .B(A[13]), .Y(n82) );
  NAND2X4 U142 ( .A(n64), .B(n69), .Y(n173) );
  NAND2XL U143 ( .A(n69), .B(n70), .Y(DIFF[0]) );
  NAND2BXL U144 ( .AN(n70), .B(n69), .Y(n65) );
  NOR2XL U145 ( .A(n37), .B(n41), .Y(n40) );
  XNOR2X4 U146 ( .A(n138), .B(n139), .Y(DIFF[14]) );
  INVX1 U147 ( .A(n94), .Y(n88) );
  NAND2X2 U148 ( .A(n47), .B(n48), .Y(n45) );
  NAND2BX4 U149 ( .AN(n130), .B(n147), .Y(n103) );
  CLKINVX3 U150 ( .A(n144), .Y(n143) );
  NOR2X1 U151 ( .A(n51), .B(n52), .Y(n50) );
  INVXL U152 ( .A(n48), .Y(n52) );
  XOR2X1 U153 ( .A(n65), .B(n66), .Y(DIFF[1]) );
  NOR2X1 U154 ( .A(n67), .B(n63), .Y(n66) );
  INVX1 U155 ( .A(n64), .Y(n67) );
  INVXL U156 ( .A(n44), .Y(n46) );
  NAND2XL U157 ( .A(n31), .B(n32), .Y(n26) );
  INVX1 U158 ( .A(n65), .Y(n62) );
  INVX1 U159 ( .A(n117), .Y(n43) );
  INVX1 U160 ( .A(n68), .Y(n63) );
  INVX1 U161 ( .A(n166), .Y(n24) );
  NAND2XL U162 ( .A(n38), .B(n39), .Y(n33) );
  XOR2X1 U163 ( .A(n56), .B(n60), .Y(DIFF[2]) );
  NOR2XL U164 ( .A(n57), .B(n61), .Y(n60) );
  INVXL U165 ( .A(n55), .Y(n61) );
  NAND2XL U166 ( .A(n58), .B(n59), .Y(n53) );
  AOI21XL U167 ( .A0(n55), .A1(n56), .B0(n57), .Y(n54) );
  NAND2BX2 U168 ( .AN(B[2]), .B(A[2]), .Y(n174) );
  NAND2BX1 U169 ( .AN(B[0]), .B(A[0]), .Y(n69) );
  NAND2BX1 U170 ( .AN(A[0]), .B(B[0]), .Y(n70) );
  NAND2BX2 U171 ( .AN(B[7]), .B(A[7]), .Y(n39) );
  NAND2XL U172 ( .A(n83), .B(n92), .Y(n155) );
  XOR2X4 U173 ( .A(n33), .B(n34), .Y(DIFF[7]) );
  XOR2X4 U174 ( .A(n118), .B(n119), .Y(DIFF[15]) );
  CLKINVX3 U175 ( .A(n120), .Y(n78) );
  NAND2BX4 U176 ( .AN(A[15]), .B(B[15]), .Y(n93) );
  NAND2BX4 U177 ( .AN(A[14]), .B(B[14]), .Y(n81) );
  NAND2BX4 U178 ( .AN(B[14]), .B(n10), .Y(n84) );
  OAI21X4 U179 ( .A0(n140), .A1(n141), .B0(n82), .Y(n138) );
  NOR2X4 U180 ( .A(n142), .B(n143), .Y(n140) );
  NAND2BX4 U181 ( .AN(A[13]), .B(B[13]), .Y(n86) );
  NAND2BX4 U182 ( .AN(A[12]), .B(B[12]), .Y(n92) );
  NAND2BX4 U183 ( .AN(B[12]), .B(A[12]), .Y(n83) );
  NAND4BX4 U184 ( .AN(n131), .B(n158), .C(n132), .D(n107), .Y(n100) );
  NAND2BX4 U185 ( .AN(B[11]), .B(A[11]), .Y(n102) );
  NAND2X4 U186 ( .A(n168), .B(n169), .Y(n23) );
  NAND4BX4 U187 ( .AN(n22), .B(n94), .C(n116), .D(n59), .Y(n29) );
  NAND3BX4 U188 ( .AN(n171), .B(n172), .C(n173), .Y(n116) );
  NAND2BX4 U189 ( .AN(B[1]), .B(A[1]), .Y(n64) );
  NAND2BX4 U190 ( .AN(A[2]), .B(B[2]), .Y(n55) );
  NAND2BX4 U191 ( .AN(A[3]), .B(B[3]), .Y(n58) );
  CLKINVX3 U192 ( .A(n174), .Y(n57) );
  CLKINVX3 U193 ( .A(n32), .Y(n161) );
  NAND2BX4 U194 ( .AN(B[4]), .B(A[4]), .Y(n48) );
  NAND2BX4 U195 ( .AN(B[5]), .B(A[5]), .Y(n44) );
  NAND2X4 U196 ( .A(n37), .B(n38), .Y(n114) );
  NAND2BX4 U197 ( .AN(A[8]), .B(B[8]), .Y(n32) );
  NAND2BX4 U198 ( .AN(B[10]), .B(A[10]), .Y(n130) );
  NAND2BX4 U199 ( .AN(A[10]), .B(B[10]), .Y(n107) );
endmodule


module butterfly_DW01_sub_82 ( A, B, DIFF );
  input [16:0] A;
  input [16:0] B;
  output [16:0] DIFF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170;

  CLKINVX3 U3 ( .A(n26), .Y(n25) );
  AOI21X2 U4 ( .A0(n76), .A1(n77), .B0(n78), .Y(n71) );
  OAI21XL U5 ( .A0(n85), .A1(n113), .B0(n114), .Y(n100) );
  XOR2X4 U6 ( .A(n6), .B(n7), .Y(DIFF[9]) );
  NOR3X4 U7 ( .A(n18), .B(n46), .C(n160), .Y(n159) );
  INVX2 U8 ( .A(n161), .Y(n18) );
  INVX8 U9 ( .A(n19), .Y(n73) );
  NAND2X2 U10 ( .A(n103), .B(n104), .Y(n88) );
  AOI31X2 U11 ( .A0(n103), .A1(n104), .A2(n105), .B0(n106), .Y(n102) );
  NOR2X2 U12 ( .A(n130), .B(n107), .Y(n134) );
  INVX1 U13 ( .A(n80), .Y(n130) );
  NAND2BX4 U14 ( .AN(A[14]), .B(B[14]), .Y(n111) );
  INVX3 U15 ( .A(n29), .Y(n31) );
  AOI21X4 U16 ( .A0(n31), .A1(n26), .B0(n24), .Y(n168) );
  NAND2BX4 U17 ( .AN(A[8]), .B(B[8]), .Y(n161) );
  NOR2X2 U18 ( .A(n107), .B(n93), .Y(n105) );
  NOR2X1 U19 ( .A(n80), .B(n93), .Y(n106) );
  NAND2BX1 U20 ( .AN(A[1]), .B(B[1]), .Y(n64) );
  NAND2X1 U21 ( .A(n110), .B(n103), .Y(n121) );
  INVX1 U22 ( .A(A[3]), .Y(n167) );
  NAND2X1 U23 ( .A(n95), .B(n110), .Y(n124) );
  NOR2X2 U24 ( .A(n34), .B(n28), .Y(n158) );
  INVX4 U25 ( .A(n145), .Y(n28) );
  XOR2X2 U26 ( .A(n52), .B(n56), .Y(DIFF[2]) );
  INVXL U27 ( .A(n51), .Y(n57) );
  NOR2X1 U28 ( .A(n82), .B(n79), .Y(n126) );
  NAND2X2 U29 ( .A(n43), .B(n44), .Y(n38) );
  CLKINVX3 U30 ( .A(n150), .Y(n34) );
  OAI21X1 U31 ( .A0(n59), .A1(n60), .B0(n61), .Y(n52) );
  INVX1 U32 ( .A(n62), .Y(n59) );
  NAND2BX2 U33 ( .AN(A[3]), .B(B[3]), .Y(n54) );
  NAND2X1 U34 ( .A(n71), .B(n72), .Y(n70) );
  NOR2X1 U35 ( .A(n84), .B(n85), .Y(n76) );
  NOR2X2 U36 ( .A(n83), .B(n85), .Y(n116) );
  NAND2X2 U37 ( .A(n117), .B(n118), .Y(n115) );
  AND3X2 U38 ( .A(n13), .B(n14), .C(n15), .Y(n6) );
  INVX1 U39 ( .A(n12), .Y(n10) );
  NAND2BX2 U40 ( .AN(A[10]), .B(B[10]), .Y(n142) );
  NAND2X2 U41 ( .A(n135), .B(n88), .Y(n133) );
  XOR2X1 U42 ( .A(n62), .B(n63), .Y(DIFF[1]) );
  INVX1 U43 ( .A(n39), .Y(n48) );
  INVX1 U44 ( .A(n14), .Y(n17) );
  NOR2X1 U45 ( .A(n24), .B(n25), .Y(n23) );
  NOR2BX4 U46 ( .AN(B[7]), .B(A[7]), .Y(n147) );
  NOR2BX1 U47 ( .AN(n95), .B(n87), .Y(n127) );
  INVX3 U48 ( .A(n87), .Y(n74) );
  NAND2BX4 U49 ( .AN(n34), .B(n35), .Y(n32) );
  INVX8 U50 ( .A(n42), .Y(n46) );
  NAND2XL U51 ( .A(n142), .B(n141), .Y(n156) );
  NAND2BX2 U52 ( .AN(A[5]), .B(B[5]), .Y(n150) );
  NAND2X2 U53 ( .A(n33), .B(n39), .Y(n144) );
  NAND2BX1 U54 ( .AN(A[2]), .B(B[2]), .Y(n163) );
  NOR2X1 U55 ( .A(n37), .B(n34), .Y(n36) );
  XNOR2X4 U56 ( .A(n67), .B(n1), .Y(DIFF[16]) );
  XNOR2X1 U57 ( .A(B[16]), .B(A[16]), .Y(n1) );
  NOR2X2 U58 ( .A(n121), .B(n107), .Y(n119) );
  NAND2BX4 U59 ( .AN(B[12]), .B(A[12]), .Y(n80) );
  NAND3BX4 U60 ( .AN(n100), .B(n101), .C(n102), .Y(n97) );
  OAI21X4 U61 ( .A0(B[3]), .A1(n167), .B0(n58), .Y(n92) );
  OAI21X1 U62 ( .A0(n79), .A1(n80), .B0(n81), .Y(n77) );
  NOR2X4 U63 ( .A(n82), .B(n83), .Y(n81) );
  NAND2BX1 U64 ( .AN(B[14]), .B(A[14]), .Y(n114) );
  NAND2BX1 U65 ( .AN(A[0]), .B(B[0]), .Y(n66) );
  OAI21X2 U66 ( .A0(n79), .A1(n80), .B0(n113), .Y(n120) );
  NAND3X4 U67 ( .A(n163), .B(n164), .C(n165), .Y(n91) );
  AND3X4 U68 ( .A(n144), .B(n145), .C(n146), .Y(n9) );
  CLKINVX3 U69 ( .A(n20), .Y(n132) );
  NOR2BX4 U70 ( .AN(n150), .B(n147), .Y(n146) );
  NAND4X1 U71 ( .A(n170), .B(n150), .C(n145), .D(n144), .Y(n169) );
  XNOR2X4 U72 ( .A(n30), .B(n4), .Y(DIFF[6]) );
  NAND2BX2 U73 ( .AN(A[6]), .B(B[6]), .Y(n145) );
  NAND2BX2 U74 ( .AN(B[6]), .B(A[6]), .Y(n29) );
  INVXL U75 ( .A(n33), .Y(n37) );
  NAND2X4 U76 ( .A(n32), .B(n33), .Y(n30) );
  NAND2BX4 U77 ( .AN(B[5]), .B(A[5]), .Y(n33) );
  NAND2BX4 U78 ( .AN(n20), .B(n112), .Y(n108) );
  NAND2X4 U79 ( .A(n73), .B(n21), .Y(n112) );
  INVX8 U80 ( .A(n112), .Y(n122) );
  OAI21X4 U81 ( .A0(n122), .A1(n20), .B0(n74), .Y(n135) );
  NOR2X4 U82 ( .A(n45), .B(n46), .Y(n43) );
  XNOR2X4 U83 ( .A(n16), .B(n5), .Y(DIFF[8]) );
  INVX1 U84 ( .A(n64), .Y(n60) );
  NOR2BX1 U85 ( .AN(n61), .B(n60), .Y(n63) );
  NOR2X1 U86 ( .A(n93), .B(n87), .Y(n109) );
  NAND2BX2 U87 ( .AN(A[15]), .B(B[15]), .Y(n96) );
  NAND2BX1 U88 ( .AN(B[15]), .B(A[15]), .Y(n99) );
  NAND2X1 U89 ( .A(n95), .B(n96), .Y(n94) );
  NAND2BX2 U90 ( .AN(A[2]), .B(B[2]), .Y(n51) );
  INVX8 U91 ( .A(n95), .Y(n107) );
  NAND3X2 U92 ( .A(n108), .B(n95), .C(n109), .Y(n101) );
  NAND2BX4 U93 ( .AN(A[12]), .B(B[12]), .Y(n95) );
  AOI21X2 U94 ( .A0(n104), .A1(n119), .B0(n120), .Y(n118) );
  NAND4X2 U95 ( .A(n51), .B(n64), .C(n54), .D(n66), .Y(n75) );
  AOI21X2 U96 ( .A0(n51), .A1(n52), .B0(n53), .Y(n50) );
  NAND2BX2 U97 ( .AN(B[2]), .B(A[2]), .Y(n58) );
  AOI31X2 U98 ( .A0(n103), .A1(n95), .A2(n104), .B0(n130), .Y(n129) );
  NAND3X2 U99 ( .A(n137), .B(n2), .C(n139), .Y(n136) );
  NAND2BX2 U100 ( .AN(B[7]), .B(A[7]), .Y(n148) );
  NAND2BX4 U101 ( .AN(B[8]), .B(A[8]), .Y(n14) );
  INVX1 U102 ( .A(B[1]), .Y(n166) );
  NOR2BX1 U103 ( .AN(B[7]), .B(A[7]), .Y(n160) );
  INVX1 U104 ( .A(n54), .Y(n45) );
  NAND2X2 U105 ( .A(n12), .B(n14), .Y(n137) );
  CLKINVX4 U106 ( .A(n75), .Y(n41) );
  INVX2 U107 ( .A(n111), .Y(n85) );
  OAI21X2 U108 ( .A0(n122), .A1(n20), .B0(n123), .Y(n117) );
  NOR2X2 U109 ( .A(n124), .B(n87), .Y(n123) );
  NOR2X2 U110 ( .A(n93), .B(n94), .Y(n68) );
  AND2X4 U111 ( .A(n162), .B(n75), .Y(n3) );
  CLKINVX4 U112 ( .A(n96), .Y(n84) );
  NAND2BX4 U113 ( .AN(n92), .B(n91), .Y(n44) );
  XOR2X2 U114 ( .A(n35), .B(n36), .Y(DIFF[5]) );
  NAND3X4 U115 ( .A(n158), .B(n21), .C(n159), .Y(n15) );
  NAND3X4 U116 ( .A(n38), .B(n39), .C(n40), .Y(n35) );
  NAND2BX4 U117 ( .AN(B[4]), .B(A[4]), .Y(n39) );
  INVX4 U118 ( .A(n148), .Y(n24) );
  XOR2X2 U119 ( .A(n49), .B(n50), .Y(DIFF[3]) );
  NAND4BX2 U120 ( .AN(n149), .B(n42), .C(n150), .D(n145), .Y(n19) );
  OAI21X4 U121 ( .A0(n27), .A1(n28), .B0(n29), .Y(n22) );
  NAND2BX4 U122 ( .AN(B[9]), .B(A[9]), .Y(n12) );
  NAND2BX4 U123 ( .AN(A[9]), .B(B[9]), .Y(n138) );
  NAND4X1 U124 ( .A(n12), .B(n14), .C(n13), .D(n15), .Y(n154) );
  INVX4 U125 ( .A(n113), .Y(n82) );
  NAND2BX4 U126 ( .AN(B[13]), .B(A[13]), .Y(n113) );
  XOR2X2 U127 ( .A(n21), .B(n47), .Y(DIFF[4]) );
  INVX4 U128 ( .A(n3), .Y(n21) );
  OAI2BB1X4 U129 ( .A0N(n168), .A1N(n169), .B0(n161), .Y(n13) );
  XOR2X4 U130 ( .A(n125), .B(n126), .Y(DIFF[13]) );
  OAI2BB1X4 U131 ( .A0N(n127), .A1N(n128), .B0(n129), .Y(n125) );
  BUFX8 U132 ( .A(n138), .Y(n2) );
  NAND2BX4 U133 ( .AN(B[10]), .B(A[10]), .Y(n141) );
  NAND2BX2 U134 ( .AN(B[11]), .B(A[11]), .Y(n140) );
  NAND2X4 U135 ( .A(n110), .B(n111), .Y(n93) );
  INVX2 U136 ( .A(n30), .Y(n27) );
  NAND2X2 U137 ( .A(n54), .B(n44), .Y(n162) );
  NAND2XL U138 ( .A(n73), .B(n21), .Y(n131) );
  NOR2BXL U139 ( .AN(n142), .B(n11), .Y(n153) );
  AOI21X2 U140 ( .A0(n68), .A1(n69), .B0(n70), .Y(n67) );
  NAND2X2 U141 ( .A(n41), .B(n42), .Y(n40) );
  OR2XL U142 ( .A(n17), .B(n18), .Y(n5) );
  INVX4 U143 ( .A(n114), .Y(n83) );
  OR2X4 U144 ( .A(n31), .B(n28), .Y(n4) );
  NAND2XL U145 ( .A(n103), .B(n140), .Y(n152) );
  AOI21XL U146 ( .A0(n89), .A1(n73), .B0(n20), .Y(n86) );
  INVXL U147 ( .A(n92), .Y(n90) );
  NAND2XL U148 ( .A(n65), .B(n66), .Y(DIFF[0]) );
  NAND2X1 U149 ( .A(n131), .B(n132), .Y(n128) );
  XNOR2X4 U150 ( .A(n151), .B(n152), .Y(DIFF[11]) );
  XNOR2X4 U151 ( .A(n155), .B(n156), .Y(DIFF[10]) );
  OR2X2 U152 ( .A(n10), .B(n11), .Y(n7) );
  NAND3X1 U153 ( .A(n13), .B(n14), .C(n15), .Y(n157) );
  NOR2XL U154 ( .A(n46), .B(n48), .Y(n47) );
  OAI21X2 U155 ( .A0(n3), .A1(n19), .B0(n132), .Y(n16) );
  INVX1 U156 ( .A(n2), .Y(n11) );
  INVX1 U157 ( .A(n58), .Y(n53) );
  AOI21XL U158 ( .A0(n90), .A1(n91), .B0(n45), .Y(n89) );
  NOR2X2 U159 ( .A(n53), .B(n57), .Y(n56) );
  NAND4XL U160 ( .A(n41), .B(n73), .C(n74), .D(n68), .Y(n72) );
  NAND2BX1 U161 ( .AN(n66), .B(n65), .Y(n62) );
  NAND2X4 U162 ( .A(n8), .B(n136), .Y(n104) );
  AND2X4 U163 ( .A(n140), .B(n141), .Y(n8) );
  OR2X4 U164 ( .A(n143), .B(n9), .Y(n20) );
  NOR2BX1 U165 ( .AN(B[7]), .B(A[7]), .Y(n149) );
  NAND2BXL U166 ( .AN(B[0]), .B(A[0]), .Y(n65) );
  OAI2BB1X2 U167 ( .A0N(A[1]), .A1N(n166), .B0(n65), .Y(n164) );
  NAND2XL U168 ( .A(n54), .B(n55), .Y(n49) );
  NAND2BXL U169 ( .AN(B[3]), .B(A[3]), .Y(n55) );
  OAI21XL U170 ( .A0(n86), .A1(n87), .B0(n88), .Y(n69) );
  OAI21X1 U171 ( .A0(n147), .A1(n29), .B0(n148), .Y(n143) );
  NAND2BXL U172 ( .AN(A[10]), .B(B[10]), .Y(n139) );
  NAND2BX1 U173 ( .AN(A[7]), .B(B[7]), .Y(n26) );
  NAND2BXL U174 ( .AN(A[7]), .B(B[7]), .Y(n170) );
  NAND2BX1 U175 ( .AN(B[1]), .B(A[1]), .Y(n61) );
  NAND2BXL U176 ( .AN(A[1]), .B(B[1]), .Y(n165) );
  XOR2X4 U177 ( .A(n22), .B(n23), .Y(DIFF[7]) );
  XOR2X4 U178 ( .A(n97), .B(n98), .Y(DIFF[15]) );
  NOR2X4 U179 ( .A(n84), .B(n78), .Y(n98) );
  CLKINVX3 U180 ( .A(n99), .Y(n78) );
  XOR2X4 U181 ( .A(n115), .B(n116), .Y(DIFF[14]) );
  CLKINVX3 U182 ( .A(n110), .Y(n79) );
  NAND2BX4 U183 ( .AN(A[13]), .B(B[13]), .Y(n110) );
  XOR2X4 U184 ( .A(n133), .B(n134), .Y(DIFF[12]) );
  NAND4BX4 U185 ( .AN(n18), .B(n2), .C(n103), .D(n142), .Y(n87) );
  NAND2BX4 U186 ( .AN(A[11]), .B(B[11]), .Y(n103) );
  OAI2BB1X4 U187 ( .A0N(n153), .A1N(n154), .B0(n141), .Y(n151) );
  OAI2BB1X4 U188 ( .A0N(n2), .A1N(n157), .B0(n12), .Y(n155) );
  NAND2BX4 U189 ( .AN(A[4]), .B(B[4]), .Y(n42) );
endmodule


module butterfly_DW01_add_88 ( A, B, SUM );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  wire   n179, n180, n181, n182, n183, n184, n185, n1, n2, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178;

  INVX2 U2 ( .A(n70), .Y(n73) );
  XOR2X4 U3 ( .A(n75), .B(B[16]), .Y(n7) );
  NOR2X4 U4 ( .A(n121), .B(n138), .Y(n114) );
  NAND2X4 U5 ( .A(n127), .B(n87), .Y(n126) );
  NOR2X4 U6 ( .A(n83), .B(n82), .Y(n81) );
  XOR2X4 U7 ( .A(n32), .B(n33), .Y(SUM[8]) );
  BUFX8 U8 ( .A(n92), .Y(n1) );
  BUFX12 U9 ( .A(n92), .Y(n2) );
  NAND2X2 U10 ( .A(B[1]), .B(n9), .Y(n178) );
  BUFX8 U11 ( .A(A[1]), .Y(n9) );
  OAI21X4 U12 ( .A0(n79), .A1(n80), .B0(n81), .Y(n78) );
  AOI21X2 U13 ( .A0(n89), .A1(n90), .B0(n91), .Y(n80) );
  OAI21X4 U14 ( .A0(B[8]), .A1(A[8]), .B0(n2), .Y(n151) );
  DLY1X1 U15 ( .A(B[10]), .Y(n12) );
  AOI31X2 U16 ( .A0(n163), .A1(n164), .A2(n165), .B0(n166), .Y(n162) );
  OAI2BB1X2 U17 ( .A0N(n167), .A1N(n154), .B0(n94), .Y(n165) );
  XOR2X4 U18 ( .A(n28), .B(n29), .Y(n180) );
  NOR2BX2 U19 ( .AN(n30), .B(n31), .Y(n29) );
  BUFX16 U20 ( .A(n182), .Y(SUM[6]) );
  BUFX12 U21 ( .A(n183), .Y(SUM[4]) );
  BUFX16 U22 ( .A(n184), .Y(SUM[3]) );
  XOR2X2 U23 ( .A(n61), .B(n62), .Y(n184) );
  NAND3X2 U24 ( .A(A[12]), .B(B[12]), .C(n84), .Y(n118) );
  NAND3X1 U25 ( .A(n86), .B(n87), .C(n88), .Y(n82) );
  CLKINVX3 U26 ( .A(n112), .Y(n173) );
  INVX2 U27 ( .A(n99), .Y(n174) );
  NOR2BX2 U28 ( .AN(n119), .B(n138), .Y(n137) );
  NOR2BX1 U29 ( .AN(n120), .B(n142), .Y(n145) );
  OAI221XL U30 ( .A0(n73), .A1(n74), .B0(n176), .B1(n177), .C0(n178), .Y(n100)
         );
  CLKINVX3 U31 ( .A(n113), .Y(n135) );
  INVX1 U32 ( .A(A[2]), .Y(n176) );
  OAI21X2 U33 ( .A0(A[3]), .A1(B[3]), .B0(n69), .Y(n101) );
  INVX1 U34 ( .A(n37), .Y(n153) );
  CLKINVX3 U35 ( .A(n137), .Y(n8) );
  INVX1 U36 ( .A(n145), .Y(n15) );
  NOR2BX2 U37 ( .AN(n146), .B(n131), .Y(n147) );
  NAND2X1 U38 ( .A(n116), .B(n85), .Y(n122) );
  XOR2X1 U39 ( .A(n58), .B(n59), .Y(n183) );
  XOR2X2 U40 ( .A(n48), .B(n49), .Y(n182) );
  BUFX8 U41 ( .A(n181), .Y(SUM[7]) );
  NOR2BX1 U42 ( .AN(n37), .B(n41), .Y(n44) );
  NOR2BX1 U43 ( .AN(n34), .B(n35), .Y(n33) );
  BUFX8 U44 ( .A(n180), .Y(SUM[9]) );
  INVX4 U45 ( .A(n88), .Y(n131) );
  NOR2X1 U46 ( .A(A[3]), .B(B[3]), .Y(n6) );
  INVX3 U47 ( .A(n87), .Y(n138) );
  NOR2X4 U48 ( .A(n153), .B(n40), .Y(n172) );
  OAI2BB1X4 U49 ( .A0N(n172), .A1N(n154), .B0(n94), .Y(n171) );
  NAND2X2 U50 ( .A(n113), .B(n93), .Y(n152) );
  NAND2X1 U51 ( .A(A[10]), .B(B[10]), .Y(n158) );
  AOI21X2 U52 ( .A0(n30), .A1(n134), .B0(n135), .Y(n133) );
  NAND4X2 U53 ( .A(n37), .B(n154), .C(n36), .D(n102), .Y(n149) );
  NAND3X2 U54 ( .A(n103), .B(n104), .C(n105), .Y(n42) );
  NAND2X1 U55 ( .A(B[15]), .B(A[15]), .Y(n116) );
  AND2X4 U56 ( .A(n93), .B(n1), .Y(n24) );
  INVX8 U57 ( .A(n102), .Y(n40) );
  INVX2 U58 ( .A(n95), .Y(n41) );
  NAND3BX1 U59 ( .AN(n46), .B(n174), .C(n95), .Y(n112) );
  XNOR2X4 U60 ( .A(n136), .B(n8), .Y(SUM[14]) );
  NOR2X2 U61 ( .A(n153), .B(n40), .Y(n167) );
  NOR2BX2 U62 ( .AN(n161), .B(n162), .Y(n160) );
  XOR2X4 U63 ( .A(n43), .B(n44), .Y(n181) );
  INVX4 U64 ( .A(n53), .Y(n50) );
  NOR2BX1 U65 ( .AN(n57), .B(n55), .Y(n59) );
  OAI2BB1X2 U66 ( .A0N(n2), .A1N(n28), .B0(n30), .Y(n168) );
  OAI21X4 U67 ( .A0(n45), .A1(n46), .B0(n47), .Y(n43) );
  NAND2X2 U68 ( .A(n30), .B(n110), .Y(n109) );
  INVX8 U69 ( .A(n25), .Y(n30) );
  NAND2X1 U70 ( .A(n84), .B(n85), .Y(n83) );
  NAND3BX2 U71 ( .AN(n131), .B(n84), .C(n87), .Y(n130) );
  INVX4 U72 ( .A(n127), .Y(n141) );
  NAND4BX2 U73 ( .AN(n99), .B(n104), .C(n95), .D(n58), .Y(n36) );
  OAI2BB1X4 U74 ( .A0N(n114), .A1N(n115), .B0(n116), .Y(n111) );
  INVX4 U75 ( .A(n111), .Y(n77) );
  NAND3X4 U76 ( .A(n164), .B(n34), .C(n171), .Y(n28) );
  NAND3BX4 U77 ( .AN(n35), .B(n58), .C(n173), .Y(n164) );
  NAND2X2 U78 ( .A(n119), .B(n120), .Y(n117) );
  INVX2 U79 ( .A(n85), .Y(n121) );
  INVX4 U80 ( .A(n48), .Y(n45) );
  NOR2X4 U81 ( .A(n16), .B(n130), .Y(n124) );
  OAI2BB1X4 U82 ( .A0N(n139), .A1N(n140), .B0(n141), .Y(n136) );
  INVX8 U83 ( .A(n14), .Y(SUM[13]) );
  OAI21X4 U84 ( .A0(A[5]), .A1(B[5]), .B0(n60), .Y(n99) );
  NAND3BX1 U85 ( .AN(n106), .B(n107), .C(n108), .Y(n79) );
  NAND2X2 U86 ( .A(B[8]), .B(A[8]), .Y(n34) );
  CLKINVX2 U87 ( .A(n106), .Y(n10) );
  OR2X2 U88 ( .A(A[11]), .B(B[11]), .Y(n86) );
  OR2X4 U89 ( .A(A[11]), .B(B[11]), .Y(n113) );
  INVX8 U90 ( .A(n157), .Y(n106) );
  NAND2X4 U91 ( .A(n78), .B(n77), .Y(n76) );
  OAI221X2 U92 ( .A0(n73), .A1(n74), .B0(n176), .B1(n177), .C0(n178), .Y(n11)
         );
  NOR2BX1 U93 ( .AN(n100), .B(n101), .Y(n96) );
  NAND4X4 U94 ( .A(n10), .B(n148), .C(n108), .D(n129), .Y(n140) );
  NAND4BX2 U95 ( .AN(n51), .B(n105), .C(n104), .D(n95), .Y(n154) );
  OR2X4 U96 ( .A(A[10]), .B(B[10]), .Y(n13) );
  AND2X2 U97 ( .A(n13), .B(n2), .Y(n21) );
  OAI2BB1X4 U98 ( .A0N(n88), .A1N(n140), .B0(n146), .Y(n144) );
  BUFX20 U99 ( .A(n179), .Y(SUM[15]) );
  INVX4 U100 ( .A(n26), .Y(n27) );
  NOR2BX4 U101 ( .AN(n108), .B(n106), .Y(n26) );
  NAND2X4 U102 ( .A(B[7]), .B(A[7]), .Y(n37) );
  XOR2X4 U103 ( .A(n144), .B(n15), .Y(n14) );
  AND2X4 U104 ( .A(n128), .B(n129), .Y(n16) );
  NOR2X4 U105 ( .A(n27), .B(n132), .Y(n128) );
  XNOR2X4 U106 ( .A(n76), .B(n7), .Y(SUM[16]) );
  CLKINVX3 U107 ( .A(A[16]), .Y(n75) );
  NAND2X4 U108 ( .A(B[4]), .B(A[4]), .Y(n57) );
  BUFX3 U109 ( .A(n185), .Y(SUM[0]) );
  NAND3X2 U110 ( .A(n21), .B(n86), .C(n155), .Y(n148) );
  AND2X2 U111 ( .A(B[9]), .B(A[9]), .Y(n25) );
  INVXL U112 ( .A(n93), .Y(n170) );
  XOR2X4 U113 ( .A(n168), .B(n169), .Y(SUM[10]) );
  NAND2BX2 U114 ( .AN(n117), .B(n118), .Y(n115) );
  NAND2X2 U115 ( .A(A[11]), .B(B[11]), .Y(n108) );
  INVX2 U116 ( .A(B[2]), .Y(n177) );
  NOR2XL U117 ( .A(A[0]), .B(B[0]), .Y(n22) );
  NOR2X1 U118 ( .A(n131), .B(n142), .Y(n139) );
  NOR2BX2 U119 ( .AN(n161), .B(n170), .Y(n169) );
  XOR2X4 U120 ( .A(n140), .B(n147), .Y(SUM[12]) );
  INVX4 U121 ( .A(n103), .Y(n51) );
  OAI21X4 U122 ( .A0(n50), .A1(n51), .B0(n52), .Y(n48) );
  NOR2BXL U123 ( .AN(n66), .B(n65), .Y(n68) );
  INVXL U124 ( .A(n63), .Y(n97) );
  OAI2BB1X2 U125 ( .A0N(B[5]), .A1N(A[5]), .B0(n57), .Y(n105) );
  OR2X4 U126 ( .A(A[2]), .B(B[2]), .Y(n69) );
  NAND2XL U127 ( .A(B[8]), .B(A[8]), .Y(n110) );
  AND2X4 U128 ( .A(n133), .B(n24), .Y(n132) );
  INVXL U129 ( .A(n74), .Y(n71) );
  NOR2BX1 U130 ( .AN(n74), .B(n22), .Y(n185) );
  INVX1 U131 ( .A(n67), .Y(n64) );
  NOR2X1 U132 ( .A(n41), .B(n42), .Y(n39) );
  NAND3X1 U133 ( .A(n36), .B(n37), .C(n38), .Y(n32) );
  NAND2XL U134 ( .A(n86), .B(n108), .Y(n159) );
  NAND4BXL U135 ( .AN(n41), .B(n2), .C(n13), .D(n94), .Y(n91) );
  NAND2X2 U136 ( .A(n30), .B(n156), .Y(n155) );
  INVX4 U137 ( .A(n94), .Y(n35) );
  NOR2BXL U138 ( .AN(n47), .B(n46), .Y(n49) );
  XOR2X1 U139 ( .A(n53), .B(n54), .Y(SUM[5]) );
  NOR2BXL U140 ( .AN(n52), .B(n51), .Y(n54) );
  INVXL U141 ( .A(n2), .Y(n31) );
  NOR2BX1 U142 ( .AN(n63), .B(n6), .Y(n62) );
  OAI21XL U143 ( .A0(n64), .A1(n65), .B0(n66), .Y(n61) );
  XOR2X1 U144 ( .A(n67), .B(n68), .Y(SUM[2]) );
  XOR2X1 U145 ( .A(n71), .B(n72), .Y(SUM[1]) );
  NOR2BXL U146 ( .AN(n178), .B(n73), .Y(n72) );
  NAND2X4 U147 ( .A(n63), .B(n175), .Y(n58) );
  INVX1 U148 ( .A(n69), .Y(n65) );
  OAI21X1 U149 ( .A0(n96), .A1(n97), .B0(n98), .Y(n90) );
  NOR2XL U150 ( .A(n99), .B(n46), .Y(n98) );
  OAI2BB1X1 U151 ( .A0N(n70), .A1N(n71), .B0(n178), .Y(n67) );
  AND2X2 U152 ( .A(n23), .B(n37), .Y(n89) );
  AND2X1 U153 ( .A(n42), .B(n102), .Y(n23) );
  NAND2X2 U154 ( .A(B[3]), .B(A[3]), .Y(n63) );
  NAND2XL U155 ( .A(B[5]), .B(A[5]), .Y(n52) );
  NAND2XL U156 ( .A(B[6]), .B(A[6]), .Y(n47) );
  NAND2XL U157 ( .A(B[2]), .B(A[2]), .Y(n66) );
  NAND2X1 U158 ( .A(B[0]), .B(A[0]), .Y(n74) );
  NAND2X1 U159 ( .A(B[8]), .B(A[8]), .Y(n156) );
  NAND2X1 U160 ( .A(B[8]), .B(A[8]), .Y(n134) );
  INVX8 U161 ( .A(n84), .Y(n142) );
  NOR2XL U162 ( .A(n39), .B(n40), .Y(n38) );
  INVX8 U163 ( .A(n104), .Y(n46) );
  NAND2X2 U164 ( .A(B[14]), .B(A[14]), .Y(n119) );
  NAND2X2 U165 ( .A(B[13]), .B(A[13]), .Y(n120) );
  NAND2XL U166 ( .A(n93), .B(n2), .Y(n166) );
  NAND3XL U167 ( .A(n2), .B(n109), .C(n13), .Y(n107) );
  NAND2XL U168 ( .A(B[12]), .B(A[12]), .Y(n146) );
  NAND2XL U169 ( .A(A[12]), .B(B[12]), .Y(n143) );
  NAND2XL U170 ( .A(n12), .B(A[10]), .Y(n161) );
  OAI21X4 U171 ( .A0(n55), .A1(n56), .B0(n57), .Y(n53) );
  CLKINVX3 U172 ( .A(n58), .Y(n56) );
  CLKINVX3 U173 ( .A(n60), .Y(n55) );
  XOR2X4 U174 ( .A(n123), .B(n122), .Y(n179) );
  NOR2X4 U175 ( .A(n124), .B(n125), .Y(n123) );
  NAND2X4 U176 ( .A(n126), .B(n119), .Y(n125) );
  OR2X4 U177 ( .A(A[15]), .B(B[15]), .Y(n85) );
  OR2X4 U178 ( .A(A[14]), .B(B[14]), .Y(n87) );
  OAI21X4 U179 ( .A0(n142), .A1(n143), .B0(n120), .Y(n127) );
  OR2X4 U180 ( .A(B[13]), .B(A[13]), .Y(n84) );
  OR2X4 U181 ( .A(A[12]), .B(B[12]), .Y(n88) );
  NAND2X4 U182 ( .A(n149), .B(n150), .Y(n129) );
  NOR2X4 U183 ( .A(n152), .B(n151), .Y(n150) );
  NAND2BX4 U184 ( .AN(n158), .B(n113), .Y(n157) );
  XOR2X4 U185 ( .A(n160), .B(n159), .Y(SUM[11]) );
  AND2X2 U186 ( .A(n30), .B(n34), .Y(n163) );
  OR2X4 U187 ( .A(B[10]), .B(A[10]), .Y(n93) );
  OR2X4 U188 ( .A(A[5]), .B(B[5]), .Y(n103) );
  NAND3X4 U189 ( .A(A[6]), .B(B[6]), .C(n95), .Y(n102) );
  OR2X4 U190 ( .A(A[7]), .B(B[7]), .Y(n95) );
  OR2X4 U191 ( .A(A[4]), .B(B[4]), .Y(n60) );
  OR2X4 U192 ( .A(A[6]), .B(B[6]), .Y(n104) );
  NAND2BX4 U193 ( .AN(n101), .B(n11), .Y(n175) );
  OR2X4 U194 ( .A(n9), .B(B[1]), .Y(n70) );
  OR2X4 U195 ( .A(B[8]), .B(A[8]), .Y(n94) );
  OR2X4 U196 ( .A(A[9]), .B(B[9]), .Y(n92) );
endmodule


module butterfly_DW01_add_103 ( A, B, SUM );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207;

  NAND3BX1 U2 ( .AN(n130), .B(n131), .C(n158), .Y(n157) );
  NAND2X2 U3 ( .A(B[11]), .B(A[11]), .Y(n124) );
  NAND3X2 U4 ( .A(n171), .B(n172), .C(n40), .Y(n1) );
  NAND2X2 U5 ( .A(n151), .B(n111), .Y(n150) );
  NAND2X4 U6 ( .A(n27), .B(n70), .Y(n79) );
  INVX4 U7 ( .A(n26), .Y(n27) );
  NAND3X4 U8 ( .A(n35), .B(n81), .C(n80), .Y(n70) );
  NAND4BX4 U9 ( .AN(n159), .B(n124), .C(n169), .D(n149), .Y(n170) );
  CLKINVX4 U10 ( .A(n142), .Y(n2) );
  CLKINVX8 U11 ( .A(n2), .Y(n3) );
  CLKINVX8 U12 ( .A(n19), .Y(n20) );
  NAND2X4 U13 ( .A(n156), .B(n157), .Y(n153) );
  CLKINVX8 U14 ( .A(n120), .Y(n163) );
  INVX2 U15 ( .A(n115), .Y(n146) );
  INVX4 U16 ( .A(n85), .Y(n74) );
  INVXL U17 ( .A(A[5]), .Y(n22) );
  INVXL U18 ( .A(A[8]), .Y(n14) );
  INVXL U19 ( .A(B[8]), .Y(n15) );
  NAND2XL U20 ( .A(B[0]), .B(A[0]), .Y(n101) );
  INVX1 U21 ( .A(n101), .Y(n97) );
  OAI21X2 U22 ( .A0(n91), .A1(n92), .B0(n93), .Y(n88) );
  NAND2X1 U23 ( .A(B[2]), .B(A[2]), .Y(n93) );
  NAND2X1 U24 ( .A(B[4]), .B(A[4]), .Y(n72) );
  INVX1 U25 ( .A(n68), .Y(n87) );
  INVX1 U26 ( .A(n71), .Y(n78) );
  OAI21XL U27 ( .A0(n108), .A1(n109), .B0(n110), .Y(n107) );
  NOR2X1 U28 ( .A(n121), .B(n122), .Y(n104) );
  AOI21X1 U29 ( .A0(n145), .A1(n111), .B0(n146), .Y(n139) );
  CLKINVX3 U30 ( .A(n64), .Y(n10) );
  NOR2X2 U31 ( .A(n165), .B(n166), .Y(n164) );
  AOI2BB1X2 U32 ( .A0N(n163), .A1N(n124), .B0(n168), .Y(n167) );
  NAND2X1 U33 ( .A(B[14]), .B(A[14]), .Y(n115) );
  NOR2X2 U34 ( .A(n173), .B(n174), .Y(n172) );
  NOR2BX1 U35 ( .AN(n184), .B(n129), .Y(n199) );
  NOR2BX1 U36 ( .AN(n45), .B(n46), .Y(n44) );
  XOR2X1 U37 ( .A(n97), .B(n99), .Y(SUM[1]) );
  CLKINVX4 U38 ( .A(n76), .Y(n73) );
  AND2X2 U39 ( .A(n118), .B(n120), .Y(n4) );
  CLKINVX3 U40 ( .A(n56), .Y(n19) );
  AND2X2 U41 ( .A(n133), .B(n134), .Y(n5) );
  AND2X4 U42 ( .A(n8), .B(n6), .Y(n156) );
  OR2X2 U43 ( .A(n143), .B(n124), .Y(n6) );
  NAND4X2 U44 ( .A(n7), .B(n138), .C(n139), .D(n140), .Y(n136) );
  OR2X4 U45 ( .A(n149), .B(n150), .Y(n7) );
  NOR2X1 U46 ( .A(n196), .B(n197), .Y(n192) );
  INVX2 U47 ( .A(n1), .Y(n29) );
  NAND2X2 U48 ( .A(n159), .B(n151), .Y(n8) );
  NOR2BX1 U49 ( .AN(n116), .B(n117), .Y(n162) );
  OR2XL U50 ( .A(A[7]), .B(B[7]), .Y(n41) );
  AOI21X2 U51 ( .A0(B[7]), .A1(A[7]), .B0(n53), .Y(n64) );
  NAND2X2 U52 ( .A(n63), .B(n10), .Y(n11) );
  NAND2X4 U53 ( .A(n9), .B(n64), .Y(n12) );
  NAND2X4 U54 ( .A(n11), .B(n12), .Y(SUM[7]) );
  INVX4 U55 ( .A(n63), .Y(n9) );
  OAI2BB1X4 U56 ( .A0N(n65), .A1N(n66), .B0(n20), .Y(n63) );
  NAND2XL U57 ( .A(n135), .B(n177), .Y(n197) );
  NAND2X4 U58 ( .A(n50), .B(n190), .Y(n200) );
  INVX8 U59 ( .A(n196), .Y(n190) );
  XNOR2X4 U60 ( .A(n32), .B(n33), .Y(SUM[5]) );
  OAI2BB1X2 U61 ( .A0N(n96), .A1N(n97), .B0(n98), .Y(n94) );
  CLKINVX8 U62 ( .A(n61), .Y(n50) );
  OR2XL U63 ( .A(A[7]), .B(B[7]), .Y(n42) );
  INVX4 U64 ( .A(n143), .Y(n151) );
  AND2X4 U65 ( .A(n111), .B(n144), .Y(n24) );
  CLKINVX8 U66 ( .A(n178), .Y(n46) );
  CLKINVX8 U67 ( .A(n177), .Y(n129) );
  NAND2X1 U68 ( .A(n195), .B(n177), .Y(n194) );
  NOR2X4 U69 ( .A(n129), .B(n183), .Y(n182) );
  NOR2X1 U70 ( .A(A[9]), .B(B[9]), .Y(n185) );
  NAND4BX2 U71 ( .AN(n189), .B(n190), .C(n191), .D(n40), .Y(n188) );
  NAND2X4 U72 ( .A(n187), .B(n188), .Y(n16) );
  CLKINVX3 U73 ( .A(n144), .Y(n130) );
  BUFX3 U74 ( .A(n76), .Y(n13) );
  NAND2X4 U75 ( .A(n69), .B(n68), .Y(n26) );
  NAND2X1 U76 ( .A(n68), .B(n85), .Y(n173) );
  NAND2X1 U77 ( .A(n71), .B(n85), .Y(n32) );
  OAI2BB1X4 U78 ( .A0N(n14), .A1N(n15), .B0(n144), .Y(n176) );
  XOR2X4 U79 ( .A(n16), .B(n17), .Y(SUM[11]) );
  AND2X1 U80 ( .A(n124), .B(n144), .Y(n17) );
  NAND2X1 U81 ( .A(n177), .B(n178), .Y(n175) );
  NAND3XL U82 ( .A(n13), .B(n135), .C(n85), .Y(n189) );
  AND2X4 U83 ( .A(n72), .B(n79), .Y(n18) );
  NOR2X4 U84 ( .A(n18), .B(n74), .Y(n77) );
  NAND2X2 U85 ( .A(n45), .B(n184), .Y(n181) );
  NAND2XL U86 ( .A(A[6]), .B(B[6]), .Y(n56) );
  NAND3BXL U87 ( .AN(n90), .B(n132), .C(n5), .Y(n125) );
  OAI21X4 U88 ( .A0(n104), .A1(n105), .B0(n106), .Y(n102) );
  NAND2XL U89 ( .A(n123), .B(n124), .Y(n122) );
  XOR2X4 U90 ( .A(n37), .B(n75), .Y(SUM[6]) );
  NAND2X2 U91 ( .A(B[5]), .B(A[5]), .Y(n71) );
  INVX3 U92 ( .A(B[5]), .Y(n23) );
  OAI21X4 U93 ( .A0(n46), .A1(n49), .B0(n45), .Y(n195) );
  CLKINVX3 U94 ( .A(n57), .Y(n55) );
  OR2X1 U95 ( .A(A[15]), .B(B[15]), .Y(n112) );
  NOR2X2 U96 ( .A(A[11]), .B(B[11]), .Y(n183) );
  NOR2X2 U97 ( .A(A[5]), .B(B[5]), .Y(n204) );
  NAND2X4 U98 ( .A(n25), .B(n62), .Y(n58) );
  NAND2XL U99 ( .A(n20), .B(n13), .Y(n75) );
  INVX8 U100 ( .A(n123), .Y(n159) );
  NOR2X4 U101 ( .A(n163), .B(n169), .Y(n165) );
  NOR3X4 U102 ( .A(n73), .B(n22), .C(n23), .Y(n21) );
  NOR2X4 U103 ( .A(n77), .B(n78), .Y(n37) );
  NAND3X1 U104 ( .A(n24), .B(n141), .C(n131), .Y(n140) );
  NOR2X4 U105 ( .A(n3), .B(n130), .Y(n179) );
  OAI21X4 U106 ( .A0(n117), .A1(n118), .B0(n116), .Y(n145) );
  AOI21X4 U107 ( .A0(n50), .A1(n40), .B0(n51), .Y(n48) );
  OAI21X4 U108 ( .A0(n52), .A1(n53), .B0(n54), .Y(n51) );
  NAND2X2 U109 ( .A(n79), .B(n72), .Y(n33) );
  NOR3BX2 U110 ( .AN(n111), .B(n143), .C(n124), .Y(n147) );
  NOR2X2 U111 ( .A(n206), .B(n207), .Y(n82) );
  OR2X2 U112 ( .A(n60), .B(n61), .Y(n25) );
  NAND4X2 U113 ( .A(n41), .B(n68), .C(n85), .D(n13), .Y(n61) );
  XOR2X4 U114 ( .A(n88), .B(n89), .Y(SUM[3]) );
  NAND2X1 U115 ( .A(B[1]), .B(A[1]), .Y(n98) );
  OR2X2 U116 ( .A(B[2]), .B(A[2]), .Y(n38) );
  NOR2X1 U117 ( .A(B[2]), .B(A[2]), .Y(n207) );
  NAND2X2 U118 ( .A(B[2]), .B(A[2]), .Y(n81) );
  NAND2X1 U119 ( .A(A[13]), .B(B[13]), .Y(n116) );
  OAI21X2 U120 ( .A0(n143), .A1(n1), .B0(n155), .Y(n154) );
  NAND2X1 U121 ( .A(B[3]), .B(A[3]), .Y(n83) );
  OR2X2 U122 ( .A(A[3]), .B(B[3]), .Y(n69) );
  OR2X4 U123 ( .A(B[1]), .B(A[1]), .Y(n96) );
  NOR2X2 U124 ( .A(n3), .B(n143), .Y(n158) );
  NAND2X4 U125 ( .A(n131), .B(n179), .Y(n169) );
  INVX4 U126 ( .A(n128), .Y(n47) );
  OR2X4 U127 ( .A(A[8]), .B(B[8]), .Y(n128) );
  NAND2X4 U128 ( .A(n28), .B(n29), .Y(n30) );
  XOR2X4 U129 ( .A(n102), .B(n103), .Y(SUM[16]) );
  NOR3BX2 U130 ( .AN(n111), .B(n123), .C(n143), .Y(n148) );
  NOR2X2 U131 ( .A(n147), .B(n148), .Y(n138) );
  NAND2X4 U132 ( .A(n34), .B(n131), .Y(n202) );
  INVX8 U133 ( .A(n40), .Y(n60) );
  XOR2X4 U134 ( .A(n40), .B(n86), .Y(SUM[4]) );
  AND2X4 U135 ( .A(n69), .B(n132), .Y(n40) );
  NOR2X2 U136 ( .A(n3), .B(n143), .Y(n141) );
  NAND2X2 U137 ( .A(n194), .B(n184), .Y(n193) );
  NAND2X2 U138 ( .A(B[10]), .B(A[10]), .Y(n184) );
  OR3X4 U139 ( .A(n73), .B(n204), .C(n205), .Y(n57) );
  NAND2X2 U140 ( .A(B[9]), .B(A[9]), .Y(n45) );
  AOI21X2 U141 ( .A0(n131), .A1(n192), .B0(n193), .Y(n187) );
  OAI21X4 U142 ( .A0(n47), .A1(n48), .B0(n49), .Y(n43) );
  NAND2X4 U143 ( .A(B[12]), .B(A[12]), .Y(n118) );
  XNOR2X4 U144 ( .A(n152), .B(n31), .Y(SUM[14]) );
  NOR2X4 U145 ( .A(n153), .B(n154), .Y(n152) );
  NAND2X4 U146 ( .A(B[8]), .B(A[8]), .Y(n49) );
  NOR3X2 U147 ( .A(n55), .B(n19), .C(n21), .Y(n52) );
  NOR2X1 U148 ( .A(n87), .B(n129), .Y(n191) );
  NOR2X4 U149 ( .A(n176), .B(n175), .Y(n171) );
  NAND2BX4 U150 ( .AN(n53), .B(n131), .Y(n62) );
  NAND2X4 U151 ( .A(n30), .B(n164), .Y(n161) );
  INVXL U152 ( .A(n163), .Y(n28) );
  OAI21X2 U153 ( .A0(n163), .A1(n123), .B0(n167), .Y(n166) );
  NOR2X1 U154 ( .A(n117), .B(n118), .Y(n113) );
  INVX2 U155 ( .A(n160), .Y(n117) );
  NOR2BX1 U156 ( .AN(n49), .B(n47), .Y(n59) );
  NAND4X2 U157 ( .A(n42), .B(n177), .C(n178), .D(n128), .Y(n142) );
  AND2X2 U158 ( .A(n83), .B(n84), .Y(n35) );
  NOR2BX1 U159 ( .AN(n98), .B(n100), .Y(n99) );
  NOR2XL U160 ( .A(n74), .B(n87), .Y(n133) );
  XNOR2X4 U161 ( .A(n136), .B(n137), .Y(SUM[15]) );
  NAND2X1 U162 ( .A(n110), .B(n112), .Y(n137) );
  AND2X1 U163 ( .A(n111), .B(n115), .Y(n31) );
  NAND2XL U164 ( .A(n115), .B(n116), .Y(n114) );
  AND2X2 U165 ( .A(n190), .B(n135), .Y(n34) );
  NAND2X4 U166 ( .A(n178), .B(n128), .Y(n196) );
  NAND2X1 U167 ( .A(n36), .B(n67), .Y(n66) );
  AND2X2 U168 ( .A(n71), .B(n72), .Y(n36) );
  NOR2X2 U169 ( .A(n185), .B(n186), .Y(n180) );
  NAND2XL U170 ( .A(B[15]), .B(A[15]), .Y(n110) );
  NOR2BX1 U171 ( .AN(n101), .B(n39), .Y(SUM[0]) );
  NOR2XL U172 ( .A(A[0]), .B(B[0]), .Y(n39) );
  INVX1 U173 ( .A(n94), .Y(n91) );
  INVX1 U174 ( .A(n195), .Y(n201) );
  AOI21X1 U175 ( .A0(n125), .A1(n62), .B0(n119), .Y(n121) );
  NAND2X1 U176 ( .A(n126), .B(n127), .Y(n119) );
  NOR2XL U177 ( .A(n129), .B(n130), .Y(n126) );
  NOR2XL U178 ( .A(n47), .B(n46), .Y(n127) );
  INVX1 U179 ( .A(n145), .Y(n155) );
  NAND2XL U180 ( .A(n135), .B(n13), .Y(n174) );
  INVX1 U181 ( .A(n82), .Y(n80) );
  INVX1 U182 ( .A(n118), .Y(n168) );
  NAND4BX2 U183 ( .AN(n82), .B(n81), .C(n83), .D(n84), .Y(n132) );
  NOR2BX2 U184 ( .AN(n72), .B(n87), .Y(n86) );
  NAND4BXL U185 ( .AN(n117), .B(n120), .C(n112), .D(n111), .Y(n105) );
  INVX1 U186 ( .A(n107), .Y(n106) );
  INVX1 U187 ( .A(n69), .Y(n90) );
  NOR2X1 U188 ( .A(n113), .B(n114), .Y(n108) );
  NAND2XL U189 ( .A(n111), .B(n112), .Y(n109) );
  NAND3XL U190 ( .A(n68), .B(n69), .C(n70), .Y(n67) );
  NAND2XL U191 ( .A(B[7]), .B(A[7]), .Y(n203) );
  NAND3BX2 U192 ( .AN(n101), .B(n96), .C(n38), .Y(n84) );
  NAND2XL U193 ( .A(B[7]), .B(A[7]), .Y(n54) );
  NAND2XL U194 ( .A(B[4]), .B(A[4]), .Y(n205) );
  XNOR2X1 U195 ( .A(n94), .B(n95), .Y(SUM[2]) );
  NAND2XL U196 ( .A(A[8]), .B(B[8]), .Y(n186) );
  XOR2X1 U197 ( .A(B[16]), .B(A[16]), .Y(n103) );
  INVXL U198 ( .A(n96), .Y(n100) );
  NAND2XL U199 ( .A(A[1]), .B(B[1]), .Y(n206) );
  NOR2XL U200 ( .A(n53), .B(n73), .Y(n134) );
  NOR2XL U201 ( .A(n73), .B(n74), .Y(n65) );
  OR2X4 U202 ( .A(A[5]), .B(B[5]), .Y(n85) );
  NOR2XL U203 ( .A(B[2]), .B(A[2]), .Y(n92) );
  OAI21XL U204 ( .A0(B[2]), .A1(A[2]), .B0(n93), .Y(n95) );
  XOR2X4 U205 ( .A(n43), .B(n44), .Y(SUM[9]) );
  XOR2X4 U206 ( .A(n58), .B(n59), .Y(SUM[8]) );
  NOR2BX4 U207 ( .AN(n83), .B(n90), .Y(n89) );
  CLKINVX3 U208 ( .A(n135), .Y(n53) );
  NAND2X4 U209 ( .A(n120), .B(n160), .Y(n143) );
  OR2X4 U210 ( .A(A[14]), .B(B[14]), .Y(n111) );
  XOR2X4 U211 ( .A(n161), .B(n162), .Y(SUM[13]) );
  OR2X4 U212 ( .A(A[13]), .B(B[13]), .Y(n160) );
  XOR2X4 U213 ( .A(n170), .B(n4), .Y(SUM[12]) );
  OR2X4 U214 ( .A(B[12]), .B(A[12]), .Y(n120) );
  NAND3X4 U215 ( .A(n171), .B(n172), .C(n40), .Y(n149) );
  OAI21X4 U216 ( .A0(n180), .A1(n181), .B0(n182), .Y(n123) );
  OR2X4 U217 ( .A(B[11]), .B(A[11]), .Y(n144) );
  XOR2X4 U218 ( .A(n198), .B(n199), .Y(SUM[10]) );
  OR2X4 U219 ( .A(B[10]), .B(A[10]), .Y(n177) );
  OAI211X2 U220 ( .A0(n200), .A1(n60), .B0(n201), .C0(n202), .Y(n198) );
  NAND4BX4 U221 ( .AN(n21), .B(n203), .C(n57), .D(n20), .Y(n131) );
  OR2X4 U222 ( .A(A[7]), .B(B[7]), .Y(n135) );
  OR2X4 U223 ( .A(A[9]), .B(B[9]), .Y(n178) );
  OR2X4 U224 ( .A(B[6]), .B(A[6]), .Y(n76) );
  OR2X4 U225 ( .A(A[4]), .B(B[4]), .Y(n68) );
endmodule


module butterfly_DW01_sub_79 ( A, B, DIFF );
  input [16:0] A;
  input [16:0] B;
  output [16:0] DIFF;
  wire   n224, n225, n226, n227, n228, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n29, n30, n31, n32, n33, n34, n35, n36, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223;

  NAND2X2 U3 ( .A(n102), .B(n108), .Y(n105) );
  NAND2X1 U4 ( .A(n62), .B(n63), .Y(n60) );
  NOR2X4 U5 ( .A(n195), .B(n194), .Y(n193) );
  CLKINVX8 U6 ( .A(n175), .Y(n29) );
  NAND3X4 U7 ( .A(n120), .B(n121), .C(n122), .Y(n118) );
  NAND2XL U8 ( .A(n189), .B(n190), .Y(n182) );
  CLKINVX3 U9 ( .A(B[5]), .Y(n72) );
  NAND2BX4 U10 ( .AN(n107), .B(n123), .Y(n122) );
  NAND3X1 U11 ( .A(n83), .B(n56), .C(n90), .Y(n86) );
  NOR3X4 U12 ( .A(n98), .B(n99), .C(n100), .Y(n216) );
  BUFX20 U13 ( .A(n73), .Y(n56) );
  NAND2BX4 U14 ( .AN(B[6]), .B(A[6]), .Y(n76) );
  NAND2BX4 U15 ( .AN(n107), .B(n6), .Y(n223) );
  NAND4BX4 U16 ( .AN(n88), .B(n56), .C(n84), .D(n89), .Y(n87) );
  NOR2X4 U17 ( .A(n105), .B(n223), .Y(n222) );
  AOI21X4 U18 ( .A0(n175), .A1(n155), .B0(n176), .Y(n174) );
  AOI21X4 U19 ( .A0(n84), .A1(n89), .B0(n114), .Y(n113) );
  NOR2X2 U20 ( .A(n176), .B(n178), .Y(n177) );
  NAND2BX4 U21 ( .AN(B[3]), .B(A[3]), .Y(n80) );
  NAND4BX1 U22 ( .AN(n107), .B(n6), .C(n102), .D(n108), .Y(n81) );
  XOR2X4 U23 ( .A(n130), .B(n131), .Y(DIFF[16]) );
  NAND4XL U24 ( .A(n42), .B(n78), .C(n79), .D(n80), .Y(n67) );
  BUFX16 U25 ( .A(n228), .Y(DIFF[5]) );
  OAI2BB1X2 U26 ( .A0N(n6), .A1N(n118), .B0(n119), .Y(n116) );
  BUFX20 U27 ( .A(n226), .Y(DIFF[7]) );
  AND2X2 U28 ( .A(n56), .B(n83), .Y(n9) );
  INVX2 U29 ( .A(n200), .Y(n62) );
  NAND2BX2 U30 ( .AN(B[9]), .B(A[9]), .Y(n57) );
  NAND2BX1 U31 ( .AN(A[13]), .B(B[13]), .Y(n150) );
  NAND2BX1 U32 ( .AN(A[14]), .B(B[14]), .Y(n149) );
  NAND2BX1 U33 ( .AN(B[13]), .B(A[13]), .Y(n146) );
  NAND4BX1 U34 ( .AN(n154), .B(n149), .C(n155), .D(n150), .Y(n137) );
  NAND2BX1 U35 ( .AN(A[15]), .B(B[15]), .Y(n144) );
  INVX1 U36 ( .A(n58), .Y(n208) );
  NAND2BX1 U37 ( .AN(n129), .B(n100), .Y(n123) );
  NOR2X2 U38 ( .A(n99), .B(n111), .Y(n220) );
  NAND2X1 U39 ( .A(n103), .B(n104), .Y(n23) );
  OR3X2 U40 ( .A(n99), .B(n100), .C(n98), .Y(n16) );
  NAND2BX2 U41 ( .AN(B[5]), .B(A[5]), .Y(n91) );
  INVX1 U42 ( .A(n123), .Y(n24) );
  INVX4 U43 ( .A(n102), .Y(n109) );
  INVX1 U44 ( .A(n80), .Y(n117) );
  BUFX8 U45 ( .A(n69), .Y(n55) );
  NAND2BX2 U46 ( .AN(B[7]), .B(A[7]), .Y(n75) );
  CLKINVX3 U47 ( .A(n201), .Y(n19) );
  NOR2X1 U48 ( .A(n194), .B(n203), .Y(n202) );
  INVX1 U49 ( .A(n202), .Y(n20) );
  NAND2X1 U50 ( .A(n57), .B(n59), .Y(n199) );
  INVX1 U51 ( .A(n186), .Y(n194) );
  INVX1 U52 ( .A(n155), .Y(n178) );
  INVX1 U53 ( .A(n177), .Y(n30) );
  INVX1 U54 ( .A(n147), .Y(n176) );
  NAND2BX2 U55 ( .AN(n182), .B(n183), .Y(n156) );
  NAND3BX2 U56 ( .AN(n184), .B(n185), .C(n186), .Y(n183) );
  OAI2BB1X2 U57 ( .A0N(n187), .A1N(B[9]), .B0(n188), .Y(n185) );
  NAND4BXL U58 ( .AN(n137), .B(n138), .C(n139), .D(n140), .Y(n136) );
  NAND2BX1 U59 ( .AN(B[11]), .B(A[11]), .Y(n157) );
  XNOR2X4 U60 ( .A(n14), .B(n15), .Y(DIFF[9]) );
  INVX2 U61 ( .A(B[4]), .Y(n18) );
  AND2X2 U62 ( .A(n65), .B(n59), .Y(n2) );
  OR2X2 U63 ( .A(n105), .B(n106), .Y(n3) );
  NAND2BX2 U64 ( .AN(A[7]), .B(B[7]), .Y(n69) );
  AND2X4 U65 ( .A(n23), .B(n3), .Y(n95) );
  NAND3X1 U66 ( .A(n126), .B(n121), .C(n127), .Y(n124) );
  NAND2X2 U67 ( .A(n4), .B(n211), .Y(n204) );
  NAND3XL U68 ( .A(n75), .B(n76), .C(n77), .Y(n38) );
  NAND2X4 U69 ( .A(n55), .B(n9), .Y(n7) );
  NAND2X1 U70 ( .A(n70), .B(n71), .Y(n39) );
  NOR2X2 U71 ( .A(n172), .B(n45), .Y(n170) );
  BUFX20 U72 ( .A(n224), .Y(DIFF[13]) );
  NAND2X4 U73 ( .A(n215), .B(n214), .Y(n4) );
  NAND2BX4 U74 ( .AN(n5), .B(n102), .Y(n98) );
  INVX8 U75 ( .A(n101), .Y(n5) );
  INVX8 U76 ( .A(n5), .Y(n6) );
  NAND3X2 U77 ( .A(n8), .B(n4), .C(n10), .Y(n61) );
  INVX4 U78 ( .A(n7), .Y(n8) );
  AND2X2 U79 ( .A(n198), .B(n84), .Y(n10) );
  INVX8 U80 ( .A(n12), .Y(DIFF[14]) );
  OAI21X2 U81 ( .A0(n38), .A1(n39), .B0(n55), .Y(n68) );
  INVX1 U82 ( .A(n210), .Y(n114) );
  NAND2XL U83 ( .A(n139), .B(n55), .Y(n160) );
  AND2X4 U84 ( .A(n139), .B(n55), .Y(n46) );
  NAND2X2 U85 ( .A(n56), .B(n55), .Y(n179) );
  OAI21X2 U86 ( .A0(n88), .A1(n210), .B0(n91), .Y(n94) );
  INVX2 U87 ( .A(n83), .Y(n88) );
  XOR2X2 U88 ( .A(n4), .B(n41), .Y(n40) );
  NAND4X4 U89 ( .A(n70), .B(n209), .C(n77), .D(n11), .Y(n63) );
  AND2X4 U90 ( .A(n75), .B(n76), .Y(n11) );
  XOR2X4 U91 ( .A(n13), .B(n169), .Y(n12) );
  AND2X2 U92 ( .A(n145), .B(n149), .Y(n13) );
  AND3X4 U93 ( .A(n59), .B(n60), .C(n61), .Y(n14) );
  AND2X1 U94 ( .A(n57), .B(n58), .Y(n15) );
  NAND3X4 U95 ( .A(n157), .B(n147), .C(n156), .Y(n172) );
  NAND2X4 U96 ( .A(n166), .B(n145), .Y(n164) );
  OAI21X2 U97 ( .A0(n167), .A1(n168), .B0(n149), .Y(n166) );
  NAND2XL U98 ( .A(n56), .B(n76), .Y(n36) );
  NOR2X2 U99 ( .A(n200), .B(n208), .Y(n206) );
  NAND2BX2 U100 ( .AN(A[9]), .B(B[9]), .Y(n192) );
  BUFX20 U101 ( .A(n225), .Y(DIFF[12]) );
  NAND2X2 U102 ( .A(n201), .B(n20), .Y(n21) );
  NOR2BX2 U103 ( .AN(A[8]), .B(B[8]), .Y(n188) );
  XOR2X4 U104 ( .A(n173), .B(n174), .Y(n224) );
  NAND3X4 U105 ( .A(n204), .B(n57), .C(n205), .Y(n201) );
  AND3X2 U106 ( .A(n84), .B(n55), .C(n56), .Y(n44) );
  NAND2X2 U107 ( .A(n84), .B(n83), .Y(n97) );
  INVX2 U108 ( .A(n84), .Y(n115) );
  NOR2X4 U109 ( .A(n109), .B(n110), .Y(n104) );
  NAND2BX4 U110 ( .AN(A[1]), .B(B[1]), .Y(n163) );
  NOR2BX4 U111 ( .AN(n16), .B(n217), .Y(n96) );
  NAND2XL U112 ( .A(n83), .B(n91), .Y(n112) );
  NAND2BX2 U113 ( .AN(B[8]), .B(A[8]), .Y(n59) );
  NOR2X1 U114 ( .A(n208), .B(n59), .Y(n207) );
  NAND4X1 U115 ( .A(n84), .B(n56), .C(n55), .D(n83), .Y(n213) );
  NAND2X4 U116 ( .A(n31), .B(n32), .Y(n225) );
  NAND2X4 U117 ( .A(n29), .B(n177), .Y(n32) );
  OAI2BB1X4 U118 ( .A0N(B[5]), .A1N(n181), .B0(n84), .Y(n180) );
  AOI21X2 U119 ( .A0(n196), .A1(n61), .B0(n197), .Y(n195) );
  INVX8 U120 ( .A(n51), .Y(DIFF[3]) );
  INVX4 U121 ( .A(n18), .Y(n17) );
  AOI21X2 U122 ( .A0(n62), .A1(n63), .B0(n199), .Y(n196) );
  XOR2X4 U123 ( .A(n116), .B(n52), .Y(n51) );
  OAI2BB1X4 U124 ( .A0N(n218), .A1N(B[3]), .B0(n219), .Y(n82) );
  AND2X2 U125 ( .A(n81), .B(n82), .Y(n42) );
  NAND2BX1 U126 ( .AN(B[2]), .B(A[2]), .Y(n119) );
  NAND2XL U127 ( .A(n82), .B(n81), .Y(n161) );
  NAND2BX4 U128 ( .AN(B[10]), .B(A[10]), .Y(n186) );
  INVX4 U129 ( .A(n210), .Y(n74) );
  NAND3X2 U130 ( .A(n72), .B(A[5]), .C(n56), .Y(n209) );
  NAND4BBX4 U131 ( .AN(B[5]), .BN(n17), .C(n56), .D(A[4]), .Y(n77) );
  NAND3X4 U132 ( .A(n56), .B(A[5]), .C(n74), .Y(n70) );
  NAND3X2 U133 ( .A(n139), .B(n140), .C(n4), .Y(n33) );
  OR2X4 U134 ( .A(n114), .B(n115), .Y(n41) );
  NAND2BX1 U135 ( .AN(n107), .B(n6), .Y(n106) );
  CLKINVX8 U136 ( .A(n6), .Y(n110) );
  INVX8 U137 ( .A(n163), .Y(n99) );
  NAND2X2 U138 ( .A(n141), .B(n104), .Y(n78) );
  OR2X4 U139 ( .A(n117), .B(n109), .Y(n52) );
  NAND2BX2 U140 ( .AN(B[1]), .B(A[1]), .Y(n120) );
  NAND2X2 U141 ( .A(n175), .B(n30), .Y(n31) );
  NOR2X4 U142 ( .A(n93), .B(n94), .Y(n92) );
  AOI21X4 U143 ( .A0(n95), .A1(n96), .B0(n97), .Y(n93) );
  AND2X4 U144 ( .A(n127), .B(n54), .Y(n128) );
  NOR2X4 U145 ( .A(n216), .B(n217), .Y(n215) );
  INVX8 U146 ( .A(A[1]), .Y(n107) );
  BUFX20 U147 ( .A(n227), .Y(DIFF[6]) );
  NAND2BX4 U148 ( .AN(B[1]), .B(A[1]), .Y(n127) );
  AOI21X2 U149 ( .A0(n206), .A1(n63), .B0(n207), .Y(n205) );
  NAND2BX4 U150 ( .AN(A[9]), .B(B[9]), .Y(n58) );
  NAND2X4 U151 ( .A(n123), .B(n108), .Y(n121) );
  INVX8 U152 ( .A(B[1]), .Y(n108) );
  INVX4 U153 ( .A(n54), .Y(n53) );
  NAND2BX4 U154 ( .AN(A[1]), .B(B[1]), .Y(n54) );
  OAI2BB1X4 U155 ( .A0N(n66), .A1N(n67), .B0(n68), .Y(n64) );
  NAND2BX4 U156 ( .AN(B[12]), .B(A[12]), .Y(n147) );
  NAND4BX4 U157 ( .AN(n45), .B(n157), .C(n156), .D(n33), .Y(n175) );
  NAND2X4 U158 ( .A(n19), .B(n202), .Y(n22) );
  NAND2X4 U159 ( .A(n21), .B(n22), .Y(DIFF[10]) );
  NOR2X1 U160 ( .A(n53), .B(n111), .Y(n103) );
  NAND2X4 U161 ( .A(n123), .B(n25), .Y(n26) );
  NAND2X2 U162 ( .A(n24), .B(n128), .Y(n27) );
  NAND2X4 U163 ( .A(n26), .B(n27), .Y(DIFF[1]) );
  INVX3 U164 ( .A(n128), .Y(n25) );
  NAND2BX4 U165 ( .AN(B[4]), .B(A[4]), .Y(n210) );
  NAND2BX4 U166 ( .AN(A[5]), .B(B[5]), .Y(n83) );
  NAND2X2 U167 ( .A(n155), .B(n150), .Y(n171) );
  NAND2BX4 U168 ( .AN(A[12]), .B(B[12]), .Y(n155) );
  INVX20 U169 ( .A(n40), .Y(DIFF[4]) );
  NAND2BXL U170 ( .AN(B[14]), .B(A[14]), .Y(n145) );
  NAND2X2 U171 ( .A(n65), .B(n55), .Y(n200) );
  INVXL U172 ( .A(n78), .Y(n138) );
  NAND2BX1 U173 ( .AN(B[15]), .B(A[15]), .Y(n134) );
  AND4X4 U174 ( .A(n191), .B(n192), .C(n189), .D(n190), .Y(n139) );
  AND2X4 U175 ( .A(n63), .B(n46), .Y(n45) );
  XNOR2X4 U176 ( .A(n164), .B(n34), .Y(DIFF[15]) );
  OR2X4 U177 ( .A(n154), .B(n165), .Y(n34) );
  NAND2XL U178 ( .A(n198), .B(n58), .Y(n212) );
  XOR2X4 U179 ( .A(n35), .B(n85), .Y(n226) );
  AND3X4 U180 ( .A(n87), .B(n86), .C(n76), .Y(n35) );
  XOR2X4 U181 ( .A(n36), .B(n92), .Y(n227) );
  XNOR2X4 U182 ( .A(n193), .B(n43), .Y(DIFF[11]) );
  AOI21XL U183 ( .A0(n146), .A1(n147), .B0(n148), .Y(n142) );
  XOR2X4 U184 ( .A(n64), .B(n2), .Y(DIFF[8]) );
  NAND2XL U185 ( .A(n55), .B(n75), .Y(n85) );
  NOR2BX2 U186 ( .AN(n119), .B(n110), .Y(n125) );
  NAND2BX1 U187 ( .AN(n107), .B(n123), .Y(n126) );
  NAND2X1 U188 ( .A(n91), .B(n210), .Y(n90) );
  NOR2X2 U189 ( .A(n212), .B(n213), .Y(n211) );
  NAND2BX1 U190 ( .AN(A[8]), .B(B[8]), .Y(n191) );
  AND2X1 U191 ( .A(n189), .B(n157), .Y(n43) );
  AND2X2 U192 ( .A(n44), .B(n83), .Y(n66) );
  INVXL U193 ( .A(n190), .Y(n203) );
  INVX1 U194 ( .A(n134), .Y(n165) );
  NOR2BX1 U195 ( .AN(A[9]), .B(B[9]), .Y(n184) );
  INVX1 U196 ( .A(n146), .Y(n167) );
  OAI21XL U197 ( .A0(n161), .A1(n162), .B0(n140), .Y(n158) );
  NAND2BX1 U198 ( .AN(A[8]), .B(B[8]), .Y(n65) );
  NAND2BX1 U199 ( .AN(A[8]), .B(B[8]), .Y(n198) );
  NAND2X1 U200 ( .A(n149), .B(n150), .Y(n148) );
  OAI21XL U201 ( .A0(n151), .A1(n152), .B0(n153), .Y(n132) );
  NAND2XL U202 ( .A(n156), .B(n157), .Y(n152) );
  INVX1 U203 ( .A(n137), .Y(n153) );
  AOI21X1 U204 ( .A0(n158), .A1(n159), .B0(n160), .Y(n151) );
  INVX1 U205 ( .A(n144), .Y(n154) );
  NAND2X1 U206 ( .A(n150), .B(n146), .Y(n173) );
  INVXL U207 ( .A(n63), .Y(n159) );
  NAND2XL U208 ( .A(n190), .B(n58), .Y(n197) );
  INVX1 U209 ( .A(A[9]), .Y(n187) );
  AND3X2 U210 ( .A(n134), .B(n135), .C(n136), .Y(n133) );
  OAI21XL U211 ( .A0(n142), .A1(n143), .B0(n144), .Y(n135) );
  INVX1 U212 ( .A(n145), .Y(n143) );
  INVXL U213 ( .A(A[5]), .Y(n181) );
  XNOR2X1 U214 ( .A(B[16]), .B(A[16]), .Y(n131) );
  NAND2X1 U215 ( .A(n132), .B(n133), .Y(n130) );
  NAND2X1 U216 ( .A(n100), .B(n129), .Y(DIFF[0]) );
  INVX1 U217 ( .A(n129), .Y(n111) );
  NAND2BX1 U218 ( .AN(B[0]), .B(A[0]), .Y(n100) );
  NAND2BX1 U219 ( .AN(A[0]), .B(B[0]), .Y(n129) );
  NAND3XL U220 ( .A(n72), .B(A[5]), .C(n56), .Y(n71) );
  NOR2BX1 U221 ( .AN(A[2]), .B(B[2]), .Y(n219) );
  NAND2X4 U222 ( .A(n82), .B(n80), .Y(n217) );
  INVXL U223 ( .A(A[3]), .Y(n218) );
  NAND4BXL U224 ( .AN(n100), .B(n54), .C(n6), .D(n102), .Y(n79) );
  NAND2XL U225 ( .A(n79), .B(n80), .Y(n162) );
  NOR2XL U226 ( .A(n53), .B(n111), .Y(n141) );
  XOR2X4 U227 ( .A(n113), .B(n112), .Y(n228) );
  XOR2X4 U228 ( .A(n125), .B(n124), .Y(DIFF[2]) );
  NOR2X4 U229 ( .A(n167), .B(n168), .Y(n169) );
  AOI21X4 U230 ( .A0(n170), .A1(n33), .B0(n171), .Y(n168) );
  NOR2X4 U231 ( .A(n179), .B(n180), .Y(n140) );
  NAND2BX4 U232 ( .AN(A[11]), .B(B[11]), .Y(n189) );
  NAND2BX4 U233 ( .AN(A[10]), .B(B[10]), .Y(n190) );
  NAND2BX4 U234 ( .AN(A[6]), .B(B[6]), .Y(n73) );
  NAND2BX4 U235 ( .AN(A[4]), .B(n17), .Y(n84) );
  NAND2X4 U236 ( .A(n215), .B(n214), .Y(n89) );
  AOI21X4 U237 ( .A0(n220), .A1(n221), .B0(n222), .Y(n214) );
  NOR2X4 U238 ( .A(n109), .B(n110), .Y(n221) );
  NAND2BX4 U239 ( .AN(A[2]), .B(B[2]), .Y(n101) );
  NAND2BX4 U240 ( .AN(A[3]), .B(B[3]), .Y(n102) );
endmodule


module butterfly_DW01_add_114 ( A, B, SUM );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  wire   n223, n224, n225, n226, n227, n228, n229, n1, n3, n7, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n24, n25, n26,
         n27, n28, n29, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222;

  NAND2X2 U2 ( .A(B[10]), .B(A[10]), .Y(n187) );
  NOR2X2 U3 ( .A(n188), .B(n189), .Y(n183) );
  NOR2X2 U4 ( .A(n186), .B(n45), .Y(n185) );
  NAND2BX4 U5 ( .AN(A[5]), .B(n87), .Y(n18) );
  BUFX1 U6 ( .A(B[2]), .Y(n11) );
  BUFX3 U7 ( .A(A[11]), .Y(n1) );
  NOR2X2 U8 ( .A(n107), .B(n108), .Y(n106) );
  AOI21X4 U9 ( .A0(n109), .A1(n110), .B0(n111), .Y(n108) );
  NAND2X4 U10 ( .A(n99), .B(n100), .Y(n13) );
  NOR4X4 U11 ( .A(n74), .B(n73), .C(n75), .D(n76), .Y(n221) );
  NAND2X1 U12 ( .A(A[2]), .B(B[2]), .Y(n113) );
  NAND2X4 U13 ( .A(B[1]), .B(A[1]), .Y(n110) );
  NOR2X2 U14 ( .A(n75), .B(n77), .Y(n207) );
  INVX4 U15 ( .A(n33), .Y(n227) );
  NAND2X1 U16 ( .A(n71), .B(n72), .Y(n175) );
  NAND4BX2 U17 ( .AN(n73), .B(n176), .C(n177), .D(n178), .Y(n71) );
  BUFX20 U18 ( .A(n226), .Y(SUM[11]) );
  NAND2X2 U19 ( .A(n60), .B(n206), .Y(n195) );
  OAI21X4 U20 ( .A0(n214), .A1(n67), .B0(n215), .Y(n210) );
  NAND2BX1 U21 ( .AN(n159), .B(n160), .Y(n149) );
  AOI21X4 U22 ( .A0(n190), .A1(n19), .B0(n159), .Y(n181) );
  OAI21X4 U23 ( .A0(n192), .A1(n191), .B0(n72), .Y(n159) );
  AND2X2 U24 ( .A(n109), .B(n110), .Y(n40) );
  AND2X2 U25 ( .A(B[1]), .B(A[1]), .Y(n219) );
  BUFX4 U26 ( .A(n102), .Y(n3) );
  OAI22X2 U27 ( .A0(n205), .A1(n212), .B0(n72), .B1(n213), .Y(n211) );
  NAND4BX4 U28 ( .AN(n73), .B(n176), .C(n177), .D(n178), .Y(n205) );
  BUFX8 U29 ( .A(n223), .Y(SUM[15]) );
  NAND2X4 U30 ( .A(n62), .B(n63), .Y(n190) );
  BUFX20 U31 ( .A(n227), .Y(SUM[9]) );
  XOR2X4 U32 ( .A(n27), .B(n40), .Y(SUM[2]) );
  NAND2X2 U33 ( .A(n204), .B(n58), .Y(n196) );
  NAND4BX2 U34 ( .AN(n50), .B(n137), .C(n190), .D(n19), .Y(n172) );
  NAND2X2 U35 ( .A(B[11]), .B(n1), .Y(n141) );
  NOR2XL U36 ( .A(n157), .B(n141), .Y(n168) );
  CLKINVX3 U37 ( .A(n194), .Y(n29) );
  INVX4 U38 ( .A(n98), .Y(n15) );
  AOI2BB1X2 U39 ( .A0N(n173), .A1N(n142), .B0(n174), .Y(n171) );
  OAI21XL U40 ( .A0(n141), .A1(n173), .B0(n131), .Y(n174) );
  NOR2BX1 U41 ( .AN(n59), .B(n198), .Y(n206) );
  AOI2BB1X2 U42 ( .A0N(n198), .A1N(n199), .B0(n200), .Y(n197) );
  NOR2BX1 U43 ( .AN(n141), .B(n45), .Y(n194) );
  BUFX3 U44 ( .A(n16), .Y(n9) );
  INVX1 U45 ( .A(n153), .Y(n182) );
  CLKINVX3 U46 ( .A(n137), .Y(n173) );
  NAND2BX1 U47 ( .AN(n157), .B(n134), .Y(n158) );
  NOR2BX1 U48 ( .AN(n134), .B(n157), .Y(n152) );
  BUFX12 U49 ( .A(n61), .Y(n19) );
  OR2X2 U50 ( .A(A[7]), .B(B[7]), .Y(n81) );
  BUFX8 U51 ( .A(n135), .Y(n50) );
  NAND2X1 U52 ( .A(B[15]), .B(A[15]), .Y(n125) );
  OR2X2 U53 ( .A(A[14]), .B(B[14]), .Y(n134) );
  OR2X2 U54 ( .A(A[15]), .B(B[15]), .Y(n126) );
  INVX1 U55 ( .A(n113), .Y(n107) );
  AOI2BB1X2 U56 ( .A0N(n73), .A1N(n85), .B0(n86), .Y(n84) );
  XOR2X2 U57 ( .A(n118), .B(n119), .Y(SUM[16]) );
  INVX8 U58 ( .A(n203), .Y(n186) );
  XOR2X4 U59 ( .A(n38), .B(n37), .Y(SUM[10]) );
  AND2X2 U60 ( .A(n52), .B(n53), .Y(n7) );
  XNOR2X4 U61 ( .A(n61), .B(n105), .Y(SUM[4]) );
  OAI21X2 U62 ( .A0(A[1]), .A1(B[1]), .B0(n115), .Y(n109) );
  NAND2X2 U63 ( .A(B[3]), .B(A[3]), .Y(n97) );
  INVX1 U64 ( .A(n97), .Y(n12) );
  INVX1 U65 ( .A(n19), .Y(n14) );
  INVX3 U66 ( .A(n112), .Y(n111) );
  NAND4BBX2 U67 ( .AN(n186), .BN(n45), .C(n53), .D(n59), .Y(n135) );
  AND2X2 U68 ( .A(n114), .B(n97), .Y(n36) );
  NAND2XL U69 ( .A(n176), .B(n88), .Y(n191) );
  NAND2X2 U70 ( .A(n142), .B(n141), .Y(n153) );
  INVX4 U71 ( .A(n181), .Y(n20) );
  NAND2X4 U72 ( .A(n99), .B(n100), .Y(n94) );
  NAND2X2 U73 ( .A(n110), .B(n116), .Y(n26) );
  OAI2BB1X4 U74 ( .A0N(n19), .A1N(n10), .B0(n68), .Y(n65) );
  NAND2X2 U75 ( .A(n24), .B(n25), .Y(n10) );
  OAI21X4 U76 ( .A0(n82), .A1(n89), .B0(n85), .Y(n90) );
  OAI211X2 U77 ( .A0(n195), .A1(n14), .B0(n196), .C0(n197), .Y(n193) );
  NAND4BXL U78 ( .AN(n74), .B(n92), .C(n88), .D(n81), .Y(n147) );
  INVX4 U79 ( .A(n205), .Y(n58) );
  NAND3BX4 U80 ( .AN(n12), .B(n16), .C(n96), .Y(n95) );
  NAND2XL U81 ( .A(n85), .B(n93), .Y(n102) );
  NAND2X2 U82 ( .A(n52), .B(n187), .Y(n184) );
  OR3X4 U83 ( .A(n13), .B(n15), .C(n12), .Y(n61) );
  OR2X2 U84 ( .A(n72), .B(n157), .Y(n39) );
  NAND2X1 U85 ( .A(n113), .B(n112), .Y(n27) );
  INVX2 U86 ( .A(n61), .Y(n67) );
  NAND2XL U87 ( .A(n99), .B(n100), .Y(n146) );
  INVX8 U88 ( .A(n15), .Y(n16) );
  NOR2X2 U89 ( .A(n75), .B(n76), .Y(n209) );
  NAND2X4 U90 ( .A(n16), .B(n97), .Y(n104) );
  NAND3BX1 U91 ( .AN(n50), .B(n137), .C(n175), .Y(n170) );
  INVX8 U92 ( .A(n17), .Y(SUM[1]) );
  XOR2X4 U93 ( .A(n115), .B(n26), .Y(n17) );
  NAND2X1 U94 ( .A(n177), .B(n178), .Y(n192) );
  NAND4BX4 U95 ( .AN(n163), .B(n164), .C(n165), .D(n166), .Y(n161) );
  AOI2BB1X2 U96 ( .A0N(n39), .A1N(n50), .B0(n168), .Y(n164) );
  NAND3X4 U97 ( .A(n60), .B(n59), .C(n19), .Y(n55) );
  OR4X2 U98 ( .A(n73), .B(n74), .C(n75), .D(n77), .Y(n24) );
  NOR2X2 U99 ( .A(n69), .B(n70), .Y(n68) );
  BUFX20 U100 ( .A(n224), .Y(SUM[14]) );
  NAND4BBX2 U101 ( .AN(n50), .BN(n157), .C(n190), .D(n19), .Y(n165) );
  XOR2X4 U102 ( .A(n90), .B(n91), .Y(n229) );
  NOR2BX2 U103 ( .AN(n87), .B(n73), .Y(n91) );
  OR2X4 U104 ( .A(B[5]), .B(n18), .Y(n178) );
  NAND2X4 U105 ( .A(B[5]), .B(A[5]), .Y(n85) );
  NAND4X4 U106 ( .A(n116), .B(n115), .C(n114), .D(n112), .Y(n98) );
  NAND2XL U107 ( .A(n9), .B(n97), .Y(n145) );
  NAND2X4 U108 ( .A(A[7]), .B(B[7]), .Y(n72) );
  BUFX20 U109 ( .A(n229), .Y(SUM[6]) );
  NOR2X1 U110 ( .A(n142), .B(n157), .Y(n163) );
  NAND2X4 U111 ( .A(n137), .B(n138), .Y(n157) );
  NOR2X2 U112 ( .A(n157), .B(n50), .Y(n167) );
  NOR4X2 U113 ( .A(n73), .B(n74), .C(n75), .D(n77), .Y(n220) );
  NOR2X4 U114 ( .A(A[11]), .B(B[11]), .Y(n45) );
  NOR2X4 U115 ( .A(n95), .B(n94), .Y(n82) );
  NOR2X4 U116 ( .A(n74), .B(n73), .Y(n208) );
  OR4X2 U117 ( .A(n73), .B(n74), .C(n76), .D(n75), .Y(n25) );
  NAND2X1 U118 ( .A(n96), .B(n92), .Y(n105) );
  NOR2X4 U119 ( .A(n104), .B(n94), .Y(n103) );
  OR2X4 U120 ( .A(A[12]), .B(B[12]), .Y(n137) );
  AOI21X2 U121 ( .A0(n167), .A1(n58), .B0(n156), .Y(n166) );
  AOI21X1 U122 ( .A0(n152), .A1(n153), .B0(n154), .Y(n151) );
  NAND2XL U123 ( .A(n155), .B(n130), .Y(n154) );
  OAI21X2 U124 ( .A0(n133), .A1(n131), .B0(n132), .Y(n156) );
  NAND2X2 U125 ( .A(B[12]), .B(A[12]), .Y(n131) );
  NAND2X4 U126 ( .A(B[13]), .B(A[13]), .Y(n132) );
  INVX4 U127 ( .A(n59), .Y(n64) );
  OR2X4 U128 ( .A(A[13]), .B(B[13]), .Y(n138) );
  OAI21X2 U129 ( .A0(n220), .A1(n221), .B0(n222), .Y(n214) );
  NAND2X4 U130 ( .A(B[6]), .B(A[6]), .Y(n87) );
  INVX4 U131 ( .A(A[7]), .Y(n77) );
  OR2X4 U132 ( .A(A[9]), .B(B[9]), .Y(n53) );
  NAND2X4 U133 ( .A(B[9]), .B(A[9]), .Y(n52) );
  INVX4 U134 ( .A(B[7]), .Y(n76) );
  BUFX20 U135 ( .A(n228), .Y(SUM[8]) );
  NAND2X4 U136 ( .A(n20), .B(n21), .Y(n22) );
  NAND2X4 U137 ( .A(n22), .B(n182), .Y(n179) );
  INVX1 U138 ( .A(n50), .Y(n21) );
  BUFX20 U139 ( .A(n225), .Y(SUM[12]) );
  NOR2BX2 U140 ( .AN(n56), .B(n64), .Y(n66) );
  OAI21X2 U141 ( .A0(n198), .A1(n56), .B0(n201), .Y(n200) );
  AOI2BB1X2 U142 ( .A0N(n216), .A1N(n56), .B0(n217), .Y(n215) );
  NAND2X2 U143 ( .A(B[8]), .B(A[8]), .Y(n56) );
  INVX4 U144 ( .A(n138), .Y(n133) );
  INVX4 U145 ( .A(n53), .Y(n216) );
  NOR2XL U146 ( .A(n64), .B(n72), .Y(n54) );
  NAND2X1 U147 ( .A(n53), .B(n59), .Y(n213) );
  INVX8 U148 ( .A(n34), .Y(SUM[13]) );
  NAND2X4 U149 ( .A(n203), .B(n53), .Y(n198) );
  INVX8 U150 ( .A(n41), .Y(n226) );
  NAND2XL U151 ( .A(n132), .B(n138), .Y(n169) );
  NOR2X2 U152 ( .A(n216), .B(n64), .Y(n222) );
  INVX8 U153 ( .A(n42), .Y(n59) );
  AND2X4 U154 ( .A(n125), .B(n126), .Y(n28) );
  OAI2BB1X2 U155 ( .A0N(n149), .A1N(n150), .B0(n151), .Y(n148) );
  INVX2 U156 ( .A(n187), .Y(n202) );
  NAND2XL U157 ( .A(n134), .B(n126), .Y(n31) );
  XNOR2X4 U158 ( .A(n35), .B(n169), .Y(n34) );
  AND3X4 U159 ( .A(n170), .B(n171), .C(n172), .Y(n35) );
  NAND2XL U160 ( .A(n53), .B(n59), .Y(n212) );
  XNOR2X4 U161 ( .A(n51), .B(n7), .Y(n33) );
  XNOR2X4 U162 ( .A(n101), .B(n3), .Y(SUM[5]) );
  INVX8 U163 ( .A(n88), .Y(n73) );
  NOR2X4 U164 ( .A(A[8]), .B(B[8]), .Y(n42) );
  NOR2XL U165 ( .A(A[9]), .B(B[9]), .Y(n188) );
  NAND2XL U166 ( .A(A[8]), .B(B[8]), .Y(n189) );
  XOR2X4 U167 ( .A(n193), .B(n29), .Y(n41) );
  XNOR2X4 U168 ( .A(n106), .B(n36), .Y(SUM[3]) );
  NOR2BXL U169 ( .AN(n131), .B(n173), .Y(n180) );
  NAND2XL U170 ( .A(n131), .B(n132), .Y(n128) );
  OAI21X1 U171 ( .A0(n123), .A1(n124), .B0(n125), .Y(n122) );
  OR2X2 U172 ( .A(n31), .B(n32), .Y(n43) );
  NAND2XL U173 ( .A(n137), .B(n138), .Y(n32) );
  OR2X4 U174 ( .A(A[1]), .B(B[1]), .Y(n116) );
  NAND3BX4 U175 ( .AN(n44), .B(n11), .C(n114), .Y(n99) );
  NAND2XL U176 ( .A(B[14]), .B(A[14]), .Y(n130) );
  NAND2BX4 U177 ( .AN(n89), .B(n88), .Y(n83) );
  INVX1 U178 ( .A(n52), .Y(n217) );
  XNOR2X4 U179 ( .A(n161), .B(n162), .Y(n224) );
  INVX1 U180 ( .A(n72), .Y(n69) );
  NAND2BX1 U181 ( .AN(n72), .B(n59), .Y(n199) );
  AOI2BB1X1 U182 ( .A0N(n186), .A1N(n52), .B0(n202), .Y(n201) );
  INVXL U183 ( .A(n87), .Y(n86) );
  INVX1 U184 ( .A(n81), .Y(n80) );
  NOR2BX1 U185 ( .AN(n59), .B(n198), .Y(n204) );
  AND2X1 U186 ( .A(n203), .B(n187), .Y(n37) );
  OR2X4 U187 ( .A(n210), .B(n211), .Y(n38) );
  NAND2X1 U188 ( .A(n130), .B(n134), .Y(n162) );
  OAI21XL U189 ( .A0(n145), .A1(n146), .B0(n136), .Y(n143) );
  INVX1 U190 ( .A(n147), .Y(n136) );
  NAND2X1 U191 ( .A(n156), .B(n134), .Y(n155) );
  NOR2BXL U192 ( .AN(n134), .B(n133), .Y(n127) );
  NOR2X1 U193 ( .A(n139), .B(n140), .Y(n120) );
  NAND2XL U194 ( .A(n141), .B(n142), .Y(n140) );
  AOI21XL U195 ( .A0(n143), .A1(n144), .B0(n50), .Y(n139) );
  NOR2X1 U196 ( .A(n69), .B(n70), .Y(n144) );
  INVX1 U197 ( .A(n130), .Y(n129) );
  NOR2XL U198 ( .A(n50), .B(n158), .Y(n150) );
  INVX1 U199 ( .A(n122), .Y(n121) );
  INVX1 U200 ( .A(n126), .Y(n124) );
  AOI21X1 U201 ( .A0(n127), .A1(n128), .B0(n129), .Y(n123) );
  INVXL U202 ( .A(A[2]), .Y(n44) );
  XOR2X1 U203 ( .A(B[16]), .B(A[16]), .Y(n119) );
  OAI21XL U204 ( .A0(n120), .A1(n43), .B0(n121), .Y(n118) );
  INVX1 U205 ( .A(n117), .Y(n115) );
  AND2X2 U206 ( .A(n117), .B(n218), .Y(SUM[0]) );
  OR2X2 U207 ( .A(A[0]), .B(B[0]), .Y(n218) );
  NAND2X1 U208 ( .A(B[0]), .B(A[0]), .Y(n117) );
  NAND2X2 U209 ( .A(n93), .B(n92), .Y(n89) );
  INVX8 U210 ( .A(n93), .Y(n74) );
  INVX8 U211 ( .A(n92), .Y(n75) );
  NAND2XL U212 ( .A(n19), .B(n190), .Y(n160) );
  NAND4BX4 U213 ( .AN(n54), .B(n55), .C(n56), .D(n57), .Y(n51) );
  NAND2X4 U214 ( .A(n58), .B(n59), .Y(n57) );
  NAND2X4 U215 ( .A(n62), .B(n63), .Y(n60) );
  XOR2X4 U216 ( .A(n65), .B(n66), .Y(n228) );
  CLKINVX3 U217 ( .A(n71), .Y(n70) );
  XOR2X4 U218 ( .A(n78), .B(n79), .Y(SUM[7]) );
  NOR2BX4 U219 ( .AN(n72), .B(n80), .Y(n79) );
  OAI21X4 U220 ( .A0(n83), .A1(n82), .B0(n84), .Y(n78) );
  OAI21X4 U221 ( .A0(n103), .A1(n75), .B0(n96), .Y(n101) );
  XOR2X4 U222 ( .A(n148), .B(n28), .Y(n223) );
  XOR2X4 U223 ( .A(n179), .B(n180), .Y(n225) );
  OAI21X4 U224 ( .A0(n183), .A1(n184), .B0(n185), .Y(n142) );
  NAND2X4 U225 ( .A(n207), .B(n208), .Y(n63) );
  NAND2X4 U226 ( .A(n209), .B(n208), .Y(n62) );
  OR2X4 U227 ( .A(A[7]), .B(B[7]), .Y(n177) );
  NAND3X4 U228 ( .A(n87), .B(n96), .C(n85), .Y(n176) );
  NAND2X4 U229 ( .A(B[4]), .B(A[4]), .Y(n96) );
  NAND3X4 U230 ( .A(n112), .B(n114), .C(n219), .Y(n100) );
  OR2X4 U231 ( .A(B[2]), .B(A[2]), .Y(n112) );
  OR2X4 U232 ( .A(A[3]), .B(B[3]), .Y(n114) );
  OR2X4 U233 ( .A(B[4]), .B(A[4]), .Y(n92) );
  OR2X4 U234 ( .A(A[5]), .B(B[5]), .Y(n93) );
  OR2X4 U235 ( .A(A[6]), .B(B[6]), .Y(n88) );
  OR2X4 U236 ( .A(A[10]), .B(B[10]), .Y(n203) );
endmodule


module butterfly_DW01_add_108 ( A, B, SUM );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  wire   n162, n1, n2, n3, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161;

  NOR2XL U2 ( .A(n40), .B(n150), .Y(n146) );
  INVX1 U3 ( .A(B[9]), .Y(n11) );
  NOR2X4 U4 ( .A(n93), .B(n94), .Y(n88) );
  NOR2X1 U5 ( .A(n19), .B(n111), .Y(n108) );
  NOR2X4 U6 ( .A(n19), .B(n97), .Y(n93) );
  NAND3X4 U7 ( .A(n34), .B(n137), .C(n1), .Y(n122) );
  INVX3 U8 ( .A(n109), .Y(n114) );
  NAND2X4 U9 ( .A(n95), .B(n96), .Y(n94) );
  NAND2X4 U10 ( .A(n27), .B(n145), .Y(n30) );
  NOR2X4 U11 ( .A(n100), .B(n98), .Y(n102) );
  NAND3X2 U12 ( .A(n46), .B(n131), .C(n132), .Y(n130) );
  BUFX12 U13 ( .A(n162), .Y(SUM[9]) );
  NAND2X4 U14 ( .A(B[8]), .B(A[8]), .Y(n45) );
  OAI211X2 U15 ( .A0(n81), .A1(n82), .B0(n79), .C0(n74), .Y(n160) );
  CLKINVX3 U16 ( .A(n77), .Y(n81) );
  OR2X4 U17 ( .A(A[4]), .B(B[4]), .Y(n66) );
  NAND2X4 U18 ( .A(B[4]), .B(A[4]), .Y(n63) );
  BUFX4 U19 ( .A(n124), .Y(n1) );
  NOR2X2 U20 ( .A(n120), .B(n7), .Y(n141) );
  NAND3BX2 U21 ( .AN(n63), .B(n55), .C(n56), .Y(n154) );
  INVXL U22 ( .A(n55), .Y(n51) );
  INVX2 U23 ( .A(n125), .Y(n120) );
  AND2X2 U24 ( .A(n121), .B(n105), .Y(n123) );
  BUFX3 U25 ( .A(B[11]), .Y(n10) );
  BUFX3 U26 ( .A(A[11]), .Y(n14) );
  INVX1 U27 ( .A(n96), .Y(n113) );
  INVX1 U28 ( .A(n145), .Y(n28) );
  NAND2X1 U29 ( .A(B[0]), .B(A[0]), .Y(n82) );
  BUFX3 U30 ( .A(B[7]), .Y(n5) );
  NOR2X2 U31 ( .A(n133), .B(n134), .Y(n32) );
  XOR2X2 U32 ( .A(n67), .B(n68), .Y(SUM[3]) );
  NOR2BX1 U33 ( .AN(n69), .B(n70), .Y(n68) );
  NAND2X2 U34 ( .A(n43), .B(n44), .Y(n42) );
  NAND2X2 U35 ( .A(n2), .B(n128), .Y(n149) );
  INVX4 U36 ( .A(n131), .Y(n40) );
  AND2X2 U37 ( .A(n46), .B(n132), .Y(n2) );
  NOR2X4 U38 ( .A(A[7]), .B(B[7]), .Y(n159) );
  INVX4 U39 ( .A(n19), .Y(n106) );
  INVX3 U40 ( .A(n11), .Y(n12) );
  AOI21X1 U41 ( .A0(n10), .A1(n14), .B0(n7), .Y(n145) );
  XNOR2X4 U42 ( .A(n32), .B(n3), .Y(SUM[12]) );
  AND2X1 U43 ( .A(n97), .B(n105), .Y(n3) );
  NAND3X4 U44 ( .A(n13), .B(n137), .C(n1), .Y(n136) );
  CLKINVX8 U45 ( .A(n99), .Y(n157) );
  INVX2 U46 ( .A(n91), .Y(n111) );
  NAND2X1 U47 ( .A(A[9]), .B(B[9]), .Y(n39) );
  INVXL U48 ( .A(n40), .Y(n6) );
  NOR2X4 U49 ( .A(n40), .B(n120), .Y(n119) );
  NOR2X1 U50 ( .A(B[11]), .B(A[11]), .Y(n7) );
  XNOR2X4 U51 ( .A(n83), .B(n8), .Y(SUM[16]) );
  XNOR2X4 U52 ( .A(B[16]), .B(A[16]), .Y(n8) );
  NAND3BX4 U53 ( .AN(n150), .B(n121), .C(n105), .Y(n129) );
  INVX4 U54 ( .A(n152), .Y(n22) );
  NOR2BX1 U55 ( .AN(n39), .B(n40), .Y(n38) );
  NAND4BX4 U56 ( .AN(n9), .B(n15), .C(n119), .D(n157), .Y(n118) );
  NAND2X2 U57 ( .A(n105), .B(n121), .Y(n9) );
  INVXL U58 ( .A(n121), .Y(n135) );
  OAI21X4 U59 ( .A0(n61), .A1(n62), .B0(n63), .Y(n57) );
  INVX4 U60 ( .A(n64), .Y(n61) );
  INVX4 U61 ( .A(n125), .Y(n150) );
  AND2X2 U62 ( .A(n127), .B(n126), .Y(n13) );
  NOR2X4 U63 ( .A(n139), .B(n140), .Y(n138) );
  NOR3BX4 U64 ( .AN(n128), .B(n129), .C(n130), .Y(n116) );
  NAND2X1 U65 ( .A(B[6]), .B(A[6]), .Y(n52) );
  INVX1 U66 ( .A(n104), .Y(n134) );
  NOR2X4 U67 ( .A(B[9]), .B(A[9]), .Y(n139) );
  AOI21X2 U68 ( .A0(n6), .A1(n37), .B0(n153), .Y(n152) );
  OAI2BB1X4 U69 ( .A0N(n146), .A1N(n147), .B0(n126), .Y(n144) );
  NAND2BX2 U70 ( .AN(n99), .B(n64), .Y(n44) );
  NAND2BX2 U71 ( .AN(n49), .B(n128), .Y(n43) );
  NAND3X4 U72 ( .A(A[5]), .B(B[5]), .C(n55), .Y(n156) );
  NAND2X2 U73 ( .A(B[3]), .B(A[3]), .Y(n69) );
  INVX2 U74 ( .A(n66), .Y(n62) );
  AND2X2 U75 ( .A(n64), .B(n46), .Y(n15) );
  XOR2X2 U76 ( .A(n37), .B(n38), .Y(n162) );
  NAND2X1 U77 ( .A(A[11]), .B(B[11]), .Y(n124) );
  NOR2X2 U78 ( .A(n143), .B(n40), .Y(n142) );
  NAND2X1 U79 ( .A(n96), .B(n106), .Y(n115) );
  NAND2X2 U80 ( .A(B[10]), .B(A[10]), .Y(n126) );
  NAND2X4 U81 ( .A(n141), .B(n142), .Y(n100) );
  OAI2BB1X4 U82 ( .A0N(n43), .A1N(n31), .B0(n102), .Y(n85) );
  XNOR2X4 U83 ( .A(n107), .B(n16), .Y(SUM[15]) );
  AND2X2 U84 ( .A(n90), .B(n92), .Y(n16) );
  XOR2X4 U85 ( .A(n112), .B(n18), .Y(n17) );
  AND2X1 U86 ( .A(n91), .B(n95), .Y(n18) );
  XOR2X2 U87 ( .A(n57), .B(n59), .Y(SUM[5]) );
  XOR2X4 U88 ( .A(n47), .B(n48), .Y(SUM[7]) );
  NAND2X4 U89 ( .A(n91), .B(n92), .Y(n89) );
  NAND2BX4 U90 ( .AN(n45), .B(n138), .Y(n127) );
  NAND3X4 U91 ( .A(A[9]), .B(n12), .C(n125), .Y(n137) );
  AOI21X1 U92 ( .A0(n103), .A1(n69), .B0(n99), .Y(n101) );
  OAI21X1 U93 ( .A0(n111), .A1(n96), .B0(n95), .Y(n110) );
  NAND2X4 U94 ( .A(A[13]), .B(B[13]), .Y(n96) );
  NAND2X4 U95 ( .A(n25), .B(n90), .Y(n87) );
  NAND4X4 U96 ( .A(n36), .B(n105), .C(n92), .D(n106), .Y(n98) );
  NAND4X1 U97 ( .A(n39), .B(n45), .C(n149), .D(n148), .Y(n147) );
  NAND3BX4 U98 ( .AN(n143), .B(n64), .C(n157), .Y(n148) );
  NOR2X4 U99 ( .A(B[13]), .B(A[13]), .Y(n19) );
  XOR2X2 U100 ( .A(n64), .B(n65), .Y(SUM[4]) );
  NAND4X4 U101 ( .A(n52), .B(n154), .C(n155), .D(n156), .Y(n128) );
  NAND3X4 U102 ( .A(n148), .B(n45), .C(n149), .Y(n37) );
  NAND2X4 U103 ( .A(n122), .B(n123), .Y(n117) );
  AND2X4 U104 ( .A(n127), .B(n126), .Y(n34) );
  NOR2X2 U105 ( .A(n104), .B(n98), .Y(n84) );
  NOR2X2 U106 ( .A(B[10]), .B(A[10]), .Y(n140) );
  NAND2X4 U107 ( .A(n69), .B(n103), .Y(n64) );
  INVX8 U108 ( .A(n17), .Y(SUM[14]) );
  NAND3BX4 U109 ( .AN(n84), .B(n85), .C(n86), .Y(n83) );
  NAND2X4 U110 ( .A(n151), .B(n22), .Y(n23) );
  NAND2X1 U111 ( .A(n21), .B(n152), .Y(n24) );
  NAND2X4 U112 ( .A(n23), .B(n24), .Y(SUM[10]) );
  INVXL U113 ( .A(n151), .Y(n21) );
  OR2X4 U114 ( .A(n88), .B(n89), .Y(n25) );
  INVX4 U115 ( .A(n87), .Y(n86) );
  AND2X2 U116 ( .A(n44), .B(n43), .Y(n26) );
  NOR2X2 U117 ( .A(n26), .B(n100), .Y(n133) );
  XOR2X2 U118 ( .A(n53), .B(n54), .Y(SUM[6]) );
  OAI2BB1X4 U119 ( .A0N(n56), .A1N(n57), .B0(n58), .Y(n53) );
  XNOR2X4 U120 ( .A(n41), .B(n42), .Y(SUM[8]) );
  NAND2X2 U121 ( .A(n144), .B(n28), .Y(n29) );
  NAND2X4 U122 ( .A(n29), .B(n30), .Y(SUM[11]) );
  INVX4 U123 ( .A(n144), .Y(n27) );
  INVX2 U124 ( .A(n46), .Y(n143) );
  INVX1 U125 ( .A(n101), .Y(n31) );
  NOR2BX1 U126 ( .AN(n52), .B(n51), .Y(n54) );
  NAND2X4 U127 ( .A(n35), .B(n160), .Y(n103) );
  NAND2X2 U128 ( .A(A[12]), .B(B[12]), .Y(n97) );
  OR2X4 U129 ( .A(A[6]), .B(B[6]), .Y(n55) );
  AND2X4 U130 ( .A(n161), .B(n71), .Y(n35) );
  INVXL U131 ( .A(n161), .Y(n73) );
  OAI21X2 U132 ( .A0(n50), .A1(n51), .B0(n52), .Y(n47) );
  INVX2 U133 ( .A(n53), .Y(n50) );
  OR2X4 U134 ( .A(A[3]), .B(B[3]), .Y(n71) );
  NOR2BX1 U135 ( .AN(n82), .B(n33), .Y(SUM[0]) );
  NOR2XL U136 ( .A(A[0]), .B(B[0]), .Y(n33) );
  NAND2X1 U137 ( .A(n45), .B(n46), .Y(n41) );
  INVX1 U138 ( .A(n75), .Y(n72) );
  NAND2XL U139 ( .A(n126), .B(n125), .Y(n151) );
  INVXL U140 ( .A(n39), .Y(n153) );
  NOR2BX1 U141 ( .AN(n63), .B(n62), .Y(n65) );
  NOR2BX1 U142 ( .AN(n58), .B(n60), .Y(n59) );
  INVXL U143 ( .A(n56), .Y(n60) );
  OAI21XL U144 ( .A0(n72), .A1(n73), .B0(n74), .Y(n67) );
  INVX1 U145 ( .A(n71), .Y(n70) );
  XOR2X1 U146 ( .A(n75), .B(n76), .Y(SUM[2]) );
  NOR2BX1 U147 ( .AN(n74), .B(n73), .Y(n76) );
  XOR2X1 U148 ( .A(n78), .B(n80), .Y(SUM[1]) );
  NOR2BXL U149 ( .AN(n79), .B(n81), .Y(n80) );
  OAI2BB1X1 U150 ( .A0N(n77), .A1N(n78), .B0(n79), .Y(n75) );
  INVX1 U151 ( .A(n82), .Y(n78) );
  NOR2XL U152 ( .A(A[5]), .B(B[5]), .Y(n158) );
  NAND2X2 U153 ( .A(B[7]), .B(A[7]), .Y(n155) );
  OR2X2 U154 ( .A(B[14]), .B(A[14]), .Y(n36) );
  AOI21XL U155 ( .A0(n5), .A1(A[7]), .B0(n49), .Y(n48) );
  NAND2X2 U156 ( .A(B[2]), .B(A[2]), .Y(n74) );
  NAND2X1 U157 ( .A(B[1]), .B(A[1]), .Y(n79) );
  NAND2XL U158 ( .A(B[15]), .B(A[15]), .Y(n90) );
  NAND2XL U159 ( .A(B[5]), .B(A[5]), .Y(n58) );
  OR2X2 U160 ( .A(A[2]), .B(B[2]), .Y(n161) );
  AOI21X4 U161 ( .A0(n109), .A1(n108), .B0(n110), .Y(n107) );
  OR2X4 U162 ( .A(A[15]), .B(B[15]), .Y(n92) );
  AOI21X4 U163 ( .A0(n109), .A1(n106), .B0(n113), .Y(n112) );
  NAND2X4 U164 ( .A(B[14]), .B(A[14]), .Y(n95) );
  OR2X4 U165 ( .A(B[14]), .B(A[14]), .Y(n91) );
  XOR2X4 U166 ( .A(n114), .B(n115), .Y(SUM[13]) );
  NAND4BX4 U167 ( .AN(n116), .B(n117), .C(n118), .D(n97), .Y(n109) );
  OR2X4 U168 ( .A(A[12]), .B(B[12]), .Y(n105) );
  NAND2BX4 U169 ( .AN(n135), .B(n136), .Y(n104) );
  CLKINVX3 U170 ( .A(n132), .Y(n49) );
  OR2X4 U171 ( .A(B[11]), .B(A[11]), .Y(n121) );
  OR2X4 U172 ( .A(A[5]), .B(B[5]), .Y(n56) );
  OR2X4 U173 ( .A(A[7]), .B(B[7]), .Y(n132) );
  NAND4BBX4 U174 ( .AN(n158), .BN(n159), .C(n55), .D(n66), .Y(n99) );
  OR2X4 U175 ( .A(A[1]), .B(B[1]), .Y(n77) );
  OR2X4 U176 ( .A(A[8]), .B(B[8]), .Y(n46) );
  OR2X4 U177 ( .A(A[9]), .B(B[9]), .Y(n131) );
  OR2X4 U178 ( .A(B[10]), .B(A[10]), .Y(n125) );
endmodule


module butterfly_DW01_add_112 ( A, B, SUM );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216;

  OAI2BB1X4 U2 ( .A0N(n1), .A1N(n2), .B0(n182), .Y(n178) );
  OR2X2 U3 ( .A(n25), .B(n40), .Y(n1) );
  AND2X2 U4 ( .A(n137), .B(n185), .Y(n2) );
  OAI21X4 U5 ( .A0(A[11]), .A1(B[11]), .B0(n46), .Y(n186) );
  INVX2 U6 ( .A(n126), .Y(n10) );
  INVX4 U7 ( .A(n120), .Y(n111) );
  AOI21XL U8 ( .A0(n118), .A1(n119), .B0(n120), .Y(n113) );
  BUFX3 U9 ( .A(n80), .Y(n3) );
  NAND2X2 U10 ( .A(B[5]), .B(A[5]), .Y(n57) );
  NOR2BX1 U11 ( .AN(n57), .B(n81), .Y(n80) );
  OR2X4 U12 ( .A(A[12]), .B(B[12]), .Y(n112) );
  NAND2X1 U13 ( .A(n52), .B(n67), .Y(n71) );
  NAND2X4 U14 ( .A(n150), .B(n151), .Y(n17) );
  NAND4BX4 U15 ( .AN(n209), .B(n68), .C(n66), .D(n67), .Y(n43) );
  NOR2X1 U16 ( .A(A[7]), .B(B[7]), .Y(n209) );
  NAND3X1 U17 ( .A(n136), .B(n137), .C(n138), .Y(n135) );
  AND3X4 U18 ( .A(n137), .B(n138), .C(n136), .Y(n7) );
  NAND2BX2 U19 ( .AN(n174), .B(n173), .Y(n138) );
  XNOR2X1 U20 ( .A(B[16]), .B(A[16]), .Y(n24) );
  NOR2X2 U21 ( .A(n61), .B(n60), .Y(n204) );
  INVXL U22 ( .A(n40), .Y(n39) );
  CLKINVX3 U23 ( .A(n12), .Y(n31) );
  NAND3X1 U24 ( .A(n155), .B(n156), .C(n48), .Y(n152) );
  NAND3X1 U25 ( .A(A[12]), .B(B[12]), .C(n110), .Y(n160) );
  NOR2BX2 U26 ( .AN(n27), .B(n15), .Y(n90) );
  NAND2X1 U27 ( .A(B[1]), .B(A[1]), .Y(n63) );
  INVX1 U28 ( .A(n43), .Y(n123) );
  INVX1 U29 ( .A(n117), .Y(n115) );
  NOR2X2 U30 ( .A(n147), .B(n148), .Y(n145) );
  AND3X2 U31 ( .A(n55), .B(n56), .C(n57), .Y(n54) );
  NAND2X2 U32 ( .A(n172), .B(n9), .Y(n139) );
  NAND2X1 U33 ( .A(B[7]), .B(A[7]), .Y(n166) );
  CLKINVX3 U34 ( .A(n183), .Y(n9) );
  NAND2X2 U35 ( .A(n210), .B(n211), .Y(n199) );
  NOR2BX2 U36 ( .AN(n47), .B(n208), .Y(n210) );
  NAND3X2 U37 ( .A(n123), .B(n201), .C(n35), .Y(n200) );
  CLKINVX3 U38 ( .A(n208), .Y(n201) );
  NOR2X1 U39 ( .A(n183), .B(n184), .Y(n182) );
  INVX4 U40 ( .A(n66), .Y(n81) );
  CLKINVX3 U41 ( .A(n91), .Y(n61) );
  CLKBUFX8 U42 ( .A(n62), .Y(n27) );
  INVX4 U43 ( .A(n4), .Y(n15) );
  CLKBUFX8 U44 ( .A(n112), .Y(n14) );
  INVX1 U45 ( .A(n99), .Y(n98) );
  AND2X2 U46 ( .A(n136), .B(n133), .Y(n18) );
  NOR2BX1 U47 ( .AN(n31), .B(n32), .Y(n30) );
  NAND3X2 U48 ( .A(n4), .B(n69), .C(n207), .Y(n74) );
  AOI21X1 U49 ( .A0(A[4]), .A1(B[4]), .B0(n76), .Y(n75) );
  OR2X4 U50 ( .A(A[2]), .B(B[2]), .Y(n4) );
  INVX1 U51 ( .A(n48), .Y(n16) );
  AND2X2 U52 ( .A(n137), .B(n9), .Y(n5) );
  NOR2X1 U53 ( .A(A[14]), .B(B[14]), .Y(n147) );
  AND2X2 U54 ( .A(n102), .B(n104), .Y(n6) );
  AND3X2 U55 ( .A(n145), .B(n146), .C(n111), .Y(n8) );
  INVX1 U56 ( .A(n68), .Y(n84) );
  OAI2BB1X2 U57 ( .A0N(n34), .A1N(n35), .B0(n36), .Y(n29) );
  NOR2X1 U58 ( .A(n43), .B(n42), .Y(n34) );
  XOR2X1 U59 ( .A(n92), .B(n94), .Y(SUM[1]) );
  NOR2BX2 U60 ( .AN(n93), .B(n61), .Y(n94) );
  NAND2X1 U61 ( .A(B[4]), .B(A[4]), .Y(n56) );
  NAND3BX4 U62 ( .AN(n168), .B(n111), .C(n35), .Y(n179) );
  AND2X2 U63 ( .A(A[5]), .B(B[5]), .Y(n21) );
  NAND2XL U64 ( .A(n107), .B(n108), .Y(n106) );
  NAND3X1 U65 ( .A(A[13]), .B(B[13]), .C(n103), .Y(n131) );
  NOR2BX4 U66 ( .AN(n67), .B(n81), .Y(n181) );
  NAND3X2 U67 ( .A(n22), .B(n75), .C(n74), .Y(n73) );
  OR2X4 U68 ( .A(A[9]), .B(B[9]), .Y(n33) );
  INVX4 U69 ( .A(n173), .Y(n183) );
  NAND2X4 U70 ( .A(n8), .B(n10), .Y(n11) );
  NAND2X4 U71 ( .A(n11), .B(n127), .Y(n125) );
  OAI21X4 U72 ( .A0(A[9]), .A1(B[9]), .B0(n46), .Y(n208) );
  NOR2X2 U73 ( .A(n213), .B(n214), .Y(n23) );
  NAND3XL U74 ( .A(n52), .B(n143), .C(n144), .Y(n211) );
  NAND3XL U75 ( .A(n143), .B(n52), .C(n144), .Y(n157) );
  NAND3BXL U76 ( .AN(n141), .B(n142), .C(n143), .Y(n140) );
  INVX8 U77 ( .A(n13), .Y(n35) );
  NOR2X1 U78 ( .A(A[9]), .B(B[9]), .Y(n189) );
  INVX2 U79 ( .A(n46), .Y(n42) );
  NAND2X1 U80 ( .A(B[14]), .B(A[14]), .Y(n107) );
  NAND2X2 U81 ( .A(n14), .B(n110), .Y(n154) );
  NAND4X1 U82 ( .A(n14), .B(n103), .C(n110), .D(n133), .Y(n129) );
  AND2X2 U83 ( .A(B[9]), .B(A[9]), .Y(n12) );
  NOR2X4 U84 ( .A(n202), .B(n203), .Y(n13) );
  XNOR2X4 U85 ( .A(n175), .B(n176), .Y(SUM[12]) );
  OAI21X2 U86 ( .A0(n96), .A1(n97), .B0(n98), .Y(n95) );
  NOR2X1 U87 ( .A(n115), .B(n116), .Y(n114) );
  NAND3X2 U88 ( .A(n20), .B(n54), .C(n53), .Y(n51) );
  NAND2X2 U89 ( .A(B[6]), .B(A[6]), .Y(n52) );
  NOR2X1 U90 ( .A(A[6]), .B(B[6]), .Y(n215) );
  AND3X2 U91 ( .A(n14), .B(n110), .C(n133), .Y(n26) );
  NOR2X2 U92 ( .A(n134), .B(n135), .Y(n128) );
  OR2X4 U93 ( .A(A[11]), .B(B[11]), .Y(n133) );
  CLKINVX4 U94 ( .A(n196), .Y(n195) );
  NOR2X2 U95 ( .A(A[6]), .B(B[6]), .Y(n213) );
  OAI2BB1X4 U96 ( .A0N(n38), .A1N(n47), .B0(n48), .Y(n44) );
  OR2X4 U97 ( .A(A[1]), .B(B[1]), .Y(n91) );
  INVX4 U98 ( .A(n14), .Y(n148) );
  NAND2X2 U99 ( .A(B[11]), .B(A[11]), .Y(n136) );
  AOI31X2 U100 ( .A0(n56), .A1(n64), .A2(n57), .B0(n65), .Y(n50) );
  NAND4BX4 U101 ( .AN(n198), .B(n199), .C(n200), .D(n31), .Y(n197) );
  NOR2BX2 U102 ( .AN(n40), .B(n42), .Y(n45) );
  NAND4BX2 U103 ( .AN(n196), .B(n46), .C(n47), .D(n38), .Y(n193) );
  NAND2XL U104 ( .A(n103), .B(n107), .Y(n149) );
  NAND3X2 U105 ( .A(n107), .B(n132), .C(n131), .Y(n130) );
  NAND3BX4 U106 ( .AN(n180), .B(n68), .C(n181), .Y(n168) );
  NAND2X1 U107 ( .A(n66), .B(n67), .Y(n65) );
  NOR2X2 U108 ( .A(A[5]), .B(B[5]), .Y(n214) );
  NOR2BX1 U109 ( .AN(n14), .B(n120), .Y(n165) );
  NAND2XL U110 ( .A(B[1]), .B(A[1]), .Y(n93) );
  OAI21X2 U111 ( .A0(n88), .A1(n15), .B0(n27), .Y(n85) );
  INVX8 U112 ( .A(n69), .Y(n87) );
  NAND2X2 U113 ( .A(n68), .B(n69), .Y(n64) );
  NAND4BX4 U114 ( .AN(n177), .B(n178), .C(n136), .D(n179), .Y(n175) );
  NOR2X1 U115 ( .A(n154), .B(n120), .Y(n153) );
  AOI2BB1X4 U116 ( .A0N(n128), .A1N(n129), .B0(n130), .Y(n127) );
  NAND2BX2 U117 ( .AN(n159), .B(n160), .Y(n158) );
  NAND2X1 U118 ( .A(B[13]), .B(A[13]), .Y(n108) );
  OAI21X2 U119 ( .A0(n100), .A1(n101), .B0(n102), .Y(n99) );
  AOI21X2 U120 ( .A0(n31), .A1(n40), .B0(n196), .Y(n192) );
  NOR2BX2 U121 ( .AN(n78), .B(n87), .Y(n86) );
  XOR2X4 U122 ( .A(n85), .B(n86), .Y(SUM[3]) );
  NAND2X1 U123 ( .A(B[3]), .B(A[3]), .Y(n78) );
  XOR2X2 U124 ( .A(n35), .B(n83), .Y(SUM[4]) );
  NAND2X2 U125 ( .A(B[8]), .B(A[8]), .Y(n40) );
  NAND4BX2 U126 ( .AN(n43), .B(n46), .C(n195), .D(n35), .Y(n194) );
  NAND4BBX4 U127 ( .AN(n191), .BN(n192), .C(n193), .D(n194), .Y(n190) );
  AOI21X2 U128 ( .A0(n37), .A1(n38), .B0(n39), .Y(n36) );
  INVX2 U129 ( .A(n89), .Y(n88) );
  NAND2BX4 U130 ( .AN(n168), .B(n35), .Y(n48) );
  OAI2BB1X4 U131 ( .A0N(n68), .A1N(n35), .B0(n82), .Y(n79) );
  OR2X4 U132 ( .A(A[6]), .B(B[6]), .Y(n67) );
  NAND3X2 U133 ( .A(n166), .B(n167), .C(n48), .Y(n164) );
  NOR2X1 U134 ( .A(A[9]), .B(B[9]), .Y(n25) );
  NOR2X2 U135 ( .A(n40), .B(n25), .Y(n172) );
  NAND2X2 U136 ( .A(n164), .B(n165), .Y(n163) );
  NOR2XL U137 ( .A(B[10]), .B(A[10]), .Y(n188) );
  NAND2X2 U138 ( .A(B[10]), .B(A[10]), .Y(n137) );
  XNOR2X2 U139 ( .A(n95), .B(n24), .Y(SUM[16]) );
  NAND2X2 U140 ( .A(n152), .B(n153), .Y(n151) );
  NOR3BX2 U141 ( .AN(n38), .B(n41), .C(n120), .Y(n177) );
  AOI21X2 U142 ( .A0(n216), .A1(n40), .B0(n208), .Y(n198) );
  OR2X4 U143 ( .A(A[3]), .B(B[3]), .Y(n69) );
  XOR2X4 U144 ( .A(n125), .B(n6), .Y(SUM[15]) );
  OR2X4 U145 ( .A(A[5]), .B(B[5]), .Y(n66) );
  AOI21X2 U146 ( .A0(n47), .A1(n140), .B0(n16), .Y(n126) );
  XOR2X2 U147 ( .A(n89), .B(n90), .Y(SUM[2]) );
  XOR2X4 U148 ( .A(n44), .B(n45), .Y(SUM[8]) );
  INVX1 U149 ( .A(n137), .Y(n191) );
  OR2X4 U150 ( .A(A[10]), .B(B[10]), .Y(n173) );
  NAND2X4 U151 ( .A(n7), .B(n139), .Y(n117) );
  AOI21X2 U152 ( .A0(n26), .A1(n117), .B0(n158), .Y(n150) );
  AOI21X4 U153 ( .A0(n169), .A1(n117), .B0(n170), .Y(n162) );
  XOR2X4 U154 ( .A(n29), .B(n30), .Y(SUM[9]) );
  NAND3BX1 U155 ( .AN(n109), .B(n103), .C(n110), .Y(n132) );
  NOR2X2 U156 ( .A(n116), .B(n148), .Y(n169) );
  NOR2BX1 U157 ( .AN(n110), .B(n109), .Y(n105) );
  INVXL U158 ( .A(n171), .Y(n170) );
  INVXL U159 ( .A(n133), .Y(n116) );
  INVX1 U160 ( .A(n133), .Y(n184) );
  OAI2BB1X1 U161 ( .A0N(n91), .A1N(n92), .B0(n93), .Y(n89) );
  NAND2X2 U162 ( .A(n171), .B(n14), .Y(n176) );
  NAND2BXL U163 ( .AN(n76), .B(n74), .Y(n122) );
  NOR2X2 U164 ( .A(n41), .B(n42), .Y(n37) );
  NAND4X4 U165 ( .A(n143), .B(n166), .C(n144), .D(n52), .Y(n38) );
  NAND2BX4 U166 ( .AN(n27), .B(n69), .Y(n124) );
  XNOR2X4 U167 ( .A(n17), .B(n149), .Y(SUM[14]) );
  NAND2X4 U168 ( .A(n78), .B(n77), .Y(n203) );
  XOR2X4 U169 ( .A(n161), .B(n19), .Y(SUM[13]) );
  AND2X1 U170 ( .A(n110), .B(n108), .Y(n19) );
  OR2XL U171 ( .A(n15), .B(n63), .Y(n20) );
  INVXL U172 ( .A(n27), .Y(n58) );
  AND2X1 U173 ( .A(n66), .B(n68), .Y(n72) );
  OR2X4 U174 ( .A(B[8]), .B(A[8]), .Y(n46) );
  OR2X4 U175 ( .A(A[7]), .B(B[7]), .Y(n47) );
  NAND2BX4 U176 ( .AN(n215), .B(n21), .Y(n143) );
  AND2X1 U177 ( .A(n77), .B(n78), .Y(n22) );
  OR2XL U178 ( .A(A[13]), .B(B[13]), .Y(n146) );
  NAND2BX4 U179 ( .AN(n212), .B(n23), .Y(n144) );
  NOR3X1 U180 ( .A(n15), .B(n60), .C(n61), .Y(n59) );
  INVXL U181 ( .A(n33), .Y(n32) );
  INVX1 U182 ( .A(n124), .Y(n76) );
  INVX1 U183 ( .A(n139), .Y(n134) );
  INVX1 U184 ( .A(n63), .Y(n207) );
  NAND2X2 U185 ( .A(n74), .B(n124), .Y(n202) );
  NOR2X1 U186 ( .A(n58), .B(n59), .Y(n53) );
  NOR2BX2 U187 ( .AN(n82), .B(n84), .Y(n83) );
  XNOR2X4 U188 ( .A(n70), .B(n71), .Y(SUM[6]) );
  INVX1 U189 ( .A(n47), .Y(n41) );
  NOR2X1 U190 ( .A(n113), .B(n114), .Y(n96) );
  OAI21XL U191 ( .A0(n121), .A1(n122), .B0(n123), .Y(n118) );
  NAND2X1 U192 ( .A(n157), .B(n47), .Y(n155) );
  NAND2XL U193 ( .A(n77), .B(n78), .Y(n121) );
  NAND2X1 U194 ( .A(n157), .B(n47), .Y(n167) );
  NAND2XL U195 ( .A(n103), .B(n104), .Y(n101) );
  NOR2X1 U196 ( .A(n105), .B(n106), .Y(n100) );
  INVX1 U197 ( .A(n108), .Y(n159) );
  NOR2X2 U198 ( .A(n188), .B(n189), .Y(n187) );
  XNOR2X4 U199 ( .A(n49), .B(n28), .Y(SUM[7]) );
  OR2X2 U200 ( .A(A[15]), .B(B[15]), .Y(n104) );
  NAND2X1 U201 ( .A(B[15]), .B(A[15]), .Y(n102) );
  NAND2XL U202 ( .A(B[3]), .B(A[3]), .Y(n55) );
  INVX1 U203 ( .A(n60), .Y(n92) );
  NAND4BXL U204 ( .AN(n147), .B(n104), .C(n14), .D(n110), .Y(n97) );
  NAND2X1 U205 ( .A(B[0]), .B(A[0]), .Y(n60) );
  AND2X2 U206 ( .A(n60), .B(n206), .Y(SUM[0]) );
  OR2X2 U207 ( .A(A[0]), .B(B[0]), .Y(n206) );
  NAND2XL U208 ( .A(B[4]), .B(A[4]), .Y(n82) );
  NAND2XL U209 ( .A(B[4]), .B(A[4]), .Y(n212) );
  NAND2XL U210 ( .A(B[12]), .B(A[12]), .Y(n171) );
  NAND2XL U211 ( .A(B[12]), .B(A[12]), .Y(n109) );
  OAI2BB1X1 U212 ( .A0N(B[7]), .A1N(A[7]), .B0(n47), .Y(n28) );
  NAND2XL U213 ( .A(B[2]), .B(A[2]), .Y(n62) );
  NAND2XL U214 ( .A(n38), .B(n47), .Y(n119) );
  NAND2XL U215 ( .A(n144), .B(n52), .Y(n141) );
  NAND2XL U216 ( .A(B[9]), .B(A[9]), .Y(n185) );
  NAND2XL U217 ( .A(A[9]), .B(B[9]), .Y(n174) );
  NAND2XL U218 ( .A(B[7]), .B(A[7]), .Y(n156) );
  NAND2XL U219 ( .A(A[7]), .B(B[7]), .Y(n142) );
  NAND2XL U220 ( .A(B[7]), .B(A[7]), .Y(n216) );
  NOR2XL U221 ( .A(A[7]), .B(B[7]), .Y(n180) );
  OAI2BB1X4 U222 ( .A0N(n50), .A1N(n51), .B0(n52), .Y(n49) );
  OAI2BB1X4 U223 ( .A0N(n72), .A1N(n73), .B0(n57), .Y(n70) );
  XOR2X4 U224 ( .A(n79), .B(n3), .Y(SUM[5]) );
  OR2X4 U225 ( .A(A[14]), .B(B[14]), .Y(n103) );
  OR2X4 U226 ( .A(A[13]), .B(B[13]), .Y(n110) );
  NAND2X4 U227 ( .A(n162), .B(n163), .Y(n161) );
  NAND2BX4 U228 ( .AN(n186), .B(n187), .Y(n120) );
  XOR2X4 U229 ( .A(n190), .B(n18), .Y(SUM[11]) );
  NAND2X4 U230 ( .A(n173), .B(n33), .Y(n196) );
  XOR2X4 U231 ( .A(n197), .B(n5), .Y(SUM[10]) );
  NAND2X4 U232 ( .A(n204), .B(n205), .Y(n77) );
  NOR2X4 U233 ( .A(n87), .B(n15), .Y(n205) );
  OR2X4 U234 ( .A(A[4]), .B(B[4]), .Y(n68) );
endmodule


module butterfly_DW01_add_113 ( A, B, SUM );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184;

  NAND2X4 U2 ( .A(n61), .B(n62), .Y(n25) );
  NAND3X2 U3 ( .A(A[9]), .B(B[9]), .C(n138), .Y(n136) );
  NAND2X2 U4 ( .A(n139), .B(n140), .Y(n135) );
  NOR3BX4 U5 ( .AN(n161), .B(n163), .C(n175), .Y(n173) );
  INVX4 U6 ( .A(n108), .Y(n127) );
  NAND2X2 U7 ( .A(n61), .B(n62), .Y(n27) );
  NAND2X2 U8 ( .A(n128), .B(n129), .Y(n122) );
  NOR2X4 U9 ( .A(n72), .B(n31), .Y(n181) );
  CLKINVX8 U10 ( .A(n182), .Y(n72) );
  CLKINVX3 U11 ( .A(n53), .Y(n162) );
  CLKINVX2 U12 ( .A(n47), .Y(n145) );
  INVX1 U13 ( .A(n42), .Y(n129) );
  NAND2X4 U14 ( .A(n3), .B(n12), .Y(n13) );
  NAND2X1 U15 ( .A(B[5]), .B(A[5]), .Y(n57) );
  NOR2X4 U16 ( .A(n91), .B(n131), .Y(n121) );
  XOR2X2 U17 ( .A(n70), .B(n71), .Y(SUM[3]) );
  CLKINVX8 U18 ( .A(n66), .Y(n11) );
  OAI2BB1X4 U19 ( .A0N(n68), .A1N(n20), .B0(n175), .Y(n66) );
  NOR2X4 U20 ( .A(n79), .B(n31), .Y(n183) );
  NOR2X1 U21 ( .A(n104), .B(n105), .Y(n100) );
  INVX4 U22 ( .A(n109), .Y(n104) );
  NOR2X2 U23 ( .A(n81), .B(n82), .Y(n180) );
  NOR2X1 U24 ( .A(n178), .B(n179), .Y(n176) );
  NOR2X2 U25 ( .A(n7), .B(n143), .Y(n169) );
  INVX1 U26 ( .A(n146), .Y(n110) );
  CLKINVX3 U27 ( .A(n138), .Y(n144) );
  NAND2BX2 U28 ( .AN(n74), .B(n182), .Y(n62) );
  CLKINVX3 U29 ( .A(n77), .Y(n81) );
  NOR2BX2 U30 ( .AN(n53), .B(n52), .Y(n55) );
  CLKINVX3 U31 ( .A(n6), .Y(n7) );
  NAND4X2 U32 ( .A(n28), .B(n171), .C(n172), .D(n39), .Y(n170) );
  OR2X2 U33 ( .A(n176), .B(n177), .Y(n28) );
  BUFX4 U34 ( .A(n35), .Y(n19) );
  INVX2 U35 ( .A(n46), .Y(n130) );
  NOR2X1 U36 ( .A(n30), .B(n127), .Y(n124) );
  NAND2X2 U37 ( .A(n48), .B(n16), .Y(n17) );
  XOR2X1 U38 ( .A(n75), .B(n76), .Y(SUM[2]) );
  NAND2BX1 U39 ( .AN(n94), .B(n85), .Y(n83) );
  OAI21XL U40 ( .A0(n95), .A1(n96), .B0(n97), .Y(n94) );
  OAI21XL U41 ( .A0(n86), .A1(n87), .B0(n88), .Y(n85) );
  INVX8 U42 ( .A(n10), .Y(n15) );
  INVX4 U43 ( .A(n60), .Y(n20) );
  OR2X4 U44 ( .A(A[5]), .B(B[5]), .Y(n161) );
  NAND2X1 U45 ( .A(B[9]), .B(A[9]), .Y(n1) );
  NAND2X1 U46 ( .A(B[10]), .B(A[10]), .Y(n140) );
  AND2X4 U47 ( .A(n63), .B(n64), .Y(n2) );
  OAI2BB1X2 U48 ( .A0N(n68), .A1N(n20), .B0(n175), .Y(n3) );
  NAND2X1 U49 ( .A(B[4]), .B(A[4]), .Y(n175) );
  OAI2BB1X2 U50 ( .A0N(n121), .A1N(n122), .B0(n123), .Y(n114) );
  NAND2XL U51 ( .A(n40), .B(n41), .Y(n157) );
  NAND2XL U52 ( .A(n65), .B(n64), .Y(n179) );
  NAND2X2 U53 ( .A(n2), .B(n65), .Y(n26) );
  AOI2BB1X4 U54 ( .A0N(n37), .A1N(n36), .B0(n155), .Y(n151) );
  INVX1 U55 ( .A(n98), .Y(n116) );
  BUFX3 U56 ( .A(n69), .Y(n4) );
  NOR2BX2 U57 ( .AN(n103), .B(n104), .Y(n120) );
  NOR2X2 U58 ( .A(n144), .B(n30), .Y(n141) );
  NOR2X4 U59 ( .A(A[11]), .B(B[11]), .Y(n30) );
  NAND2X4 U60 ( .A(n65), .B(n64), .Y(n24) );
  NAND3BX4 U61 ( .AN(n39), .B(n19), .C(n138), .Y(n137) );
  OR2X4 U62 ( .A(A[1]), .B(B[1]), .Y(n77) );
  AOI21X2 U63 ( .A0(n160), .A1(n148), .B0(n162), .Y(n159) );
  NOR2XL U64 ( .A(n52), .B(n59), .Y(n22) );
  OAI21X1 U65 ( .A0(n73), .A1(n31), .B0(n74), .Y(n70) );
  NAND2BX2 U66 ( .AN(n164), .B(n53), .Y(n174) );
  NOR2BX1 U67 ( .AN(n64), .B(n72), .Y(n71) );
  NOR2BXL U68 ( .AN(n74), .B(n31), .Y(n76) );
  XNOR2X4 U69 ( .A(n168), .B(n5), .Y(SUM[10]) );
  NAND2XL U70 ( .A(n140), .B(n138), .Y(n5) );
  NAND3BX4 U71 ( .AN(n45), .B(n41), .C(n42), .Y(n38) );
  INVX2 U72 ( .A(n45), .Y(n6) );
  OR2X4 U73 ( .A(A[12]), .B(B[12]), .Y(n108) );
  INVX8 U74 ( .A(n54), .Y(n51) );
  NAND4XL U75 ( .A(n146), .B(n167), .C(n161), .D(n147), .Y(n177) );
  OR2X4 U76 ( .A(A[6]), .B(B[6]), .Y(n167) );
  OAI21X4 U77 ( .A0(n134), .A1(n91), .B0(n89), .Y(n132) );
  INVX2 U78 ( .A(n49), .Y(n16) );
  AOI21X2 U79 ( .A0(B[7]), .A1(A[7]), .B0(n50), .Y(n49) );
  NAND2X4 U80 ( .A(B[1]), .B(A[1]), .Y(n79) );
  NAND2X1 U81 ( .A(B[11]), .B(A[11]), .Y(n139) );
  NAND2X2 U82 ( .A(B[3]), .B(A[3]), .Y(n64) );
  AND2X2 U83 ( .A(A[5]), .B(B[5]), .Y(n33) );
  OR2X2 U84 ( .A(A[9]), .B(B[9]), .Y(n35) );
  OAI2BB1X4 U85 ( .A0N(n121), .A1N(n122), .B0(n123), .Y(n8) );
  OAI21X4 U86 ( .A0(n173), .A1(n174), .B0(n41), .Y(n171) );
  NOR2X4 U87 ( .A(A[6]), .B(B[6]), .Y(n163) );
  XOR2X4 U88 ( .A(n114), .B(n120), .Y(SUM[13]) );
  NAND2X2 U89 ( .A(B[8]), .B(A[8]), .Y(n39) );
  NAND4X2 U90 ( .A(n167), .B(n146), .C(n20), .D(n161), .Y(n46) );
  AOI21X4 U91 ( .A0(n130), .A1(n9), .B0(n145), .Y(n134) );
  NOR2BX4 U92 ( .AN(n57), .B(n59), .Y(n67) );
  AOI21X4 U93 ( .A0(n125), .A1(n124), .B0(n126), .Y(n123) );
  NAND2X4 U94 ( .A(n165), .B(n166), .Y(n37) );
  NAND2X4 U95 ( .A(n11), .B(n67), .Y(n14) );
  XOR2X4 U96 ( .A(n9), .B(n4), .Y(SUM[4]) );
  NAND2X2 U97 ( .A(n130), .B(n9), .Y(n128) );
  OAI21X4 U98 ( .A0(n52), .A1(n51), .B0(n53), .Y(n48) );
  XOR2X4 U99 ( .A(n112), .B(n111), .Y(SUM[15]) );
  NAND2BX4 U100 ( .AN(n30), .B(n125), .Y(n89) );
  AND2X2 U101 ( .A(n1), .B(n19), .Y(n23) );
  OAI211X2 U102 ( .A0(n37), .A1(n36), .B0(n38), .C0(n39), .Y(n34) );
  NAND2X2 U103 ( .A(n183), .B(n182), .Y(n61) );
  OAI21X4 U104 ( .A0(n26), .A1(n27), .B0(n58), .Y(n56) );
  NOR2X4 U105 ( .A(n59), .B(n60), .Y(n58) );
  INVX4 U106 ( .A(n67), .Y(n12) );
  AOI21X2 U107 ( .A0(n113), .A1(n8), .B0(n115), .Y(n112) );
  OR2X4 U108 ( .A(A[6]), .B(B[6]), .Y(n32) );
  NAND2X1 U109 ( .A(B[12]), .B(A[12]), .Y(n105) );
  INVX8 U110 ( .A(n36), .Y(n9) );
  CLKINVX8 U111 ( .A(n68), .Y(n36) );
  NAND2X1 U112 ( .A(n108), .B(n41), .Y(n131) );
  NAND2BX2 U113 ( .AN(n157), .B(n42), .Y(n156) );
  NOR2X2 U114 ( .A(n63), .B(n163), .Y(n160) );
  NOR2BX1 U115 ( .AN(n139), .B(n30), .Y(n150) );
  OAI21X4 U116 ( .A0(n51), .A1(n52), .B0(n53), .Y(n10) );
  NAND2X4 U117 ( .A(B[6]), .B(A[6]), .Y(n53) );
  NOR2BX2 U118 ( .AN(n79), .B(n81), .Y(n80) );
  NAND2X4 U119 ( .A(B[2]), .B(A[2]), .Y(n74) );
  OAI2BB1X4 U120 ( .A0N(n77), .A1N(n78), .B0(n79), .Y(n75) );
  OR2X4 U121 ( .A(A[3]), .B(B[3]), .Y(n182) );
  INVX12 U122 ( .A(n167), .Y(n52) );
  AOI21X4 U123 ( .A0(B[7]), .A1(A[7]), .B0(n164), .Y(n158) );
  NOR2BX1 U124 ( .AN(n63), .B(n60), .Y(n69) );
  XOR2X4 U125 ( .A(n132), .B(n133), .Y(SUM[12]) );
  NAND2X2 U126 ( .A(n156), .B(n39), .Y(n155) );
  INVX8 U127 ( .A(n148), .Y(n59) );
  INVX8 U128 ( .A(n19), .Y(n143) );
  XOR2X2 U129 ( .A(n78), .B(n80), .Y(SUM[1]) );
  NOR2X4 U130 ( .A(A[2]), .B(B[2]), .Y(n31) );
  OR2X4 U131 ( .A(A[8]), .B(B[8]), .Y(n40) );
  NOR2X4 U132 ( .A(n110), .B(n45), .Y(n165) );
  OAI21X2 U133 ( .A0(n36), .A1(n46), .B0(n47), .Y(n43) );
  NAND2X4 U134 ( .A(n42), .B(n41), .Y(n47) );
  AND2X4 U135 ( .A(n33), .B(n32), .Y(n164) );
  NAND3BX4 U136 ( .AN(n135), .B(n136), .C(n137), .Y(n125) );
  INVX8 U137 ( .A(n40), .Y(n45) );
  OR2X4 U138 ( .A(A[10]), .B(B[10]), .Y(n138) );
  OR2X4 U139 ( .A(A[14]), .B(B[14]), .Y(n98) );
  XOR2X4 U140 ( .A(n34), .B(n23), .Y(SUM[9]) );
  OR2X4 U141 ( .A(A[7]), .B(B[7]), .Y(n41) );
  INVX3 U142 ( .A(n41), .Y(n50) );
  XOR2X2 U143 ( .A(n54), .B(n55), .Y(SUM[6]) );
  XOR2X2 U144 ( .A(n43), .B(n44), .Y(SUM[8]) );
  NAND2X4 U145 ( .A(n13), .B(n14), .Y(SUM[5]) );
  NAND2X4 U146 ( .A(n15), .B(n49), .Y(n18) );
  NAND2X4 U147 ( .A(n17), .B(n18), .Y(SUM[7]) );
  NAND2X4 U148 ( .A(B[4]), .B(A[4]), .Y(n63) );
  NOR3BX2 U149 ( .AN(n167), .B(n60), .C(n59), .Y(n166) );
  OR2X4 U150 ( .A(A[7]), .B(B[7]), .Y(n146) );
  OR2X4 U151 ( .A(B[5]), .B(A[5]), .Y(n148) );
  NOR2BX2 U152 ( .AN(n105), .B(n127), .Y(n133) );
  INVX1 U153 ( .A(n105), .Y(n126) );
  NOR2BX1 U154 ( .AN(n39), .B(n45), .Y(n44) );
  INVXL U155 ( .A(n89), .Y(n87) );
  AND2X2 U156 ( .A(n21), .B(n22), .Y(n29) );
  NOR2XL U157 ( .A(n60), .B(n110), .Y(n21) );
  OR2X4 U158 ( .A(n24), .B(n25), .Y(n68) );
  NAND2X2 U159 ( .A(n97), .B(n99), .Y(n111) );
  OAI21XL U160 ( .A0(n116), .A1(n103), .B0(n102), .Y(n115) );
  INVX2 U161 ( .A(n75), .Y(n73) );
  NAND2XL U162 ( .A(n98), .B(n99), .Y(n96) );
  INVXL U163 ( .A(n140), .Y(n154) );
  NOR2XL U164 ( .A(n104), .B(n116), .Y(n113) );
  NAND2X1 U165 ( .A(n98), .B(n102), .Y(n117) );
  INVXL U166 ( .A(n103), .Y(n119) );
  NAND2XL U167 ( .A(n61), .B(n62), .Y(n178) );
  NAND2XL U168 ( .A(n138), .B(n19), .Y(n152) );
  AOI2BB1X2 U169 ( .A0N(n144), .A1N(n1), .B0(n154), .Y(n153) );
  OAI21XL U170 ( .A0(n92), .A1(n93), .B0(n29), .Y(n90) );
  NAND2XL U171 ( .A(n62), .B(n61), .Y(n93) );
  NOR2X1 U172 ( .A(n100), .B(n101), .Y(n95) );
  NAND2XL U173 ( .A(n102), .B(n103), .Y(n101) );
  NOR2X1 U174 ( .A(n106), .B(n107), .Y(n88) );
  NAND2XL U175 ( .A(n108), .B(n109), .Y(n107) );
  NAND2X1 U176 ( .A(n99), .B(n98), .Y(n106) );
  NAND2XL U177 ( .A(B[14]), .B(A[14]), .Y(n102) );
  OR2X2 U178 ( .A(A[15]), .B(B[15]), .Y(n99) );
  NAND2X1 U179 ( .A(B[15]), .B(A[15]), .Y(n97) );
  INVX1 U180 ( .A(n82), .Y(n78) );
  XOR2X1 U181 ( .A(B[16]), .B(A[16]), .Y(n84) );
  AND2X2 U182 ( .A(n82), .B(n184), .Y(SUM[0]) );
  OR2X2 U183 ( .A(A[0]), .B(B[0]), .Y(n184) );
  NAND2X1 U184 ( .A(B[0]), .B(A[0]), .Y(n82) );
  OR2X2 U185 ( .A(A[13]), .B(B[13]), .Y(n109) );
  NAND2X1 U186 ( .A(B[13]), .B(A[13]), .Y(n103) );
  AOI21XL U187 ( .A0(n90), .A1(n47), .B0(n91), .Y(n86) );
  NAND2XL U188 ( .A(n65), .B(n64), .Y(n92) );
  INVX8 U189 ( .A(n147), .Y(n60) );
  NAND2XL U190 ( .A(B[7]), .B(A[7]), .Y(n172) );
  NAND2X4 U191 ( .A(n56), .B(n57), .Y(n54) );
  XOR2X4 U192 ( .A(n83), .B(n84), .Y(SUM[16]) );
  XOR2X4 U193 ( .A(n117), .B(n118), .Y(SUM[14]) );
  AOI21X4 U194 ( .A0(n109), .A1(n8), .B0(n119), .Y(n118) );
  NAND2X4 U195 ( .A(n141), .B(n142), .Y(n91) );
  NOR2X4 U196 ( .A(n7), .B(n143), .Y(n142) );
  XOR2X4 U197 ( .A(n149), .B(n150), .Y(SUM[11]) );
  OAI21X4 U198 ( .A0(n151), .A1(n152), .B0(n153), .Y(n149) );
  NAND2X4 U199 ( .A(n158), .B(n159), .Y(n42) );
  OAI2BB1X4 U200 ( .A0N(n169), .A1N(n170), .B0(n1), .Y(n168) );
  OR2X4 U201 ( .A(B[4]), .B(A[4]), .Y(n147) );
  NAND2X4 U202 ( .A(n180), .B(n181), .Y(n65) );
endmodule


module butterfly_DW01_sub_95 ( A, B, DIFF );
  input [16:0] A;
  input [16:0] B;
  output [16:0] DIFF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201;

  NAND4X2 U3 ( .A(n122), .B(n108), .C(n63), .D(n21), .Y(n41) );
  INVX4 U4 ( .A(n169), .Y(n33) );
  NAND3X4 U5 ( .A(n169), .B(n167), .C(n38), .Y(n165) );
  NAND2X4 U6 ( .A(n53), .B(n4), .Y(n61) );
  NAND2BX4 U7 ( .AN(A[2]), .B(B[2]), .Y(n76) );
  NAND2X2 U8 ( .A(n78), .B(n79), .Y(n122) );
  NAND2X4 U9 ( .A(n38), .B(n47), .Y(n193) );
  OAI21X4 U10 ( .A0(n36), .A1(n37), .B0(n38), .Y(n31) );
  OR2X2 U11 ( .A(n131), .B(n114), .Y(n138) );
  OAI21X4 U12 ( .A0(A[7]), .A1(n39), .B0(n53), .Y(n197) );
  INVX3 U13 ( .A(B[7]), .Y(n39) );
  NOR2X4 U14 ( .A(n48), .B(n193), .Y(n192) );
  INVX2 U15 ( .A(A[7]), .Y(n30) );
  OAI21X1 U16 ( .A0(A[7]), .A1(n39), .B0(n40), .Y(n37) );
  AOI21X4 U17 ( .A0(n2), .A1(n42), .B0(n43), .Y(n36) );
  NAND2X2 U18 ( .A(n10), .B(n22), .Y(n170) );
  AOI21X4 U19 ( .A0(n54), .A1(n125), .B0(n126), .Y(n124) );
  OAI2BB1X4 U20 ( .A0N(n148), .A1N(n14), .B0(n127), .Y(n126) );
  NOR2X2 U21 ( .A(n135), .B(n105), .Y(n125) );
  OAI21X4 U22 ( .A0(n44), .A1(n45), .B0(n46), .Y(n43) );
  AOI21X2 U23 ( .A0(n53), .A1(n2), .B0(n71), .Y(n70) );
  NAND2X1 U24 ( .A(n53), .B(n29), .Y(n51) );
  INVX4 U25 ( .A(n53), .Y(n73) );
  NAND2XL U26 ( .A(n114), .B(n22), .Y(n157) );
  INVX8 U27 ( .A(n114), .Y(n148) );
  NAND2X2 U28 ( .A(n133), .B(n100), .Y(n132) );
  NAND4BX2 U29 ( .AN(n99), .B(n100), .C(n110), .D(n102), .Y(n91) );
  INVX8 U30 ( .A(n111), .Y(n99) );
  NOR2X4 U31 ( .A(A[11]), .B(n15), .Y(n161) );
  AOI21X2 U32 ( .A0(n148), .A1(n110), .B0(n149), .Y(n147) );
  NAND2X4 U33 ( .A(n15), .B(A[11]), .Y(n115) );
  NAND2XL U34 ( .A(n133), .B(n110), .Y(n145) );
  INVX4 U35 ( .A(n110), .Y(n153) );
  NAND2BX1 U36 ( .AN(B[2]), .B(A[2]), .Y(n201) );
  OAI21X2 U37 ( .A0(n142), .A1(n104), .B0(n103), .Y(n128) );
  BUFX8 U38 ( .A(n115), .Y(n22) );
  NAND2X2 U39 ( .A(n82), .B(n86), .Y(n200) );
  XOR2X2 U40 ( .A(n11), .B(n12), .Y(DIFF[2]) );
  INVXL U41 ( .A(n77), .Y(n11) );
  NAND2BX2 U42 ( .AN(B[1]), .B(A[1]), .Y(n82) );
  NAND2X1 U43 ( .A(n134), .B(n100), .Y(n135) );
  NOR2X1 U44 ( .A(n144), .B(n142), .Y(n143) );
  AOI21X2 U45 ( .A0(n33), .A1(n162), .B0(n176), .Y(n175) );
  CLKINVX3 U46 ( .A(n170), .Y(n17) );
  NAND2X1 U47 ( .A(n8), .B(n9), .Y(n10) );
  INVX1 U48 ( .A(n50), .Y(n44) );
  CLKBUFX8 U49 ( .A(n82), .Y(n28) );
  INVX1 U50 ( .A(n67), .Y(n71) );
  NOR3BX2 U51 ( .AN(n93), .B(n94), .C(n95), .Y(n92) );
  XOR2X1 U52 ( .A(n2), .B(n72), .Y(DIFF[4]) );
  NOR2X1 U53 ( .A(n71), .B(n73), .Y(n72) );
  CLKINVX3 U54 ( .A(n122), .Y(n65) );
  INVX4 U55 ( .A(n105), .Y(n140) );
  CLKINVX4 U56 ( .A(n41), .Y(n1) );
  INVX8 U57 ( .A(n1), .Y(n2) );
  AOI21X2 U58 ( .A0(n118), .A1(n106), .B0(n119), .Y(n116) );
  NOR2X2 U59 ( .A(n180), .B(n196), .Y(n195) );
  BUFX8 U60 ( .A(n52), .Y(n27) );
  NAND4BXL U61 ( .AN(n121), .B(n53), .C(n4), .D(n29), .Y(n109) );
  INVX1 U62 ( .A(n109), .Y(n106) );
  NAND2BX1 U63 ( .AN(n78), .B(n76), .Y(n12) );
  INVX8 U64 ( .A(n59), .Y(n3) );
  INVX8 U65 ( .A(n29), .Y(n59) );
  BUFX8 U66 ( .A(n49), .Y(n29) );
  NAND2X1 U67 ( .A(n29), .B(n27), .Y(n45) );
  NAND2BX2 U68 ( .AN(B[6]), .B(A[6]), .Y(n194) );
  INVX8 U69 ( .A(n180), .Y(n4) );
  INVX4 U70 ( .A(n52), .Y(n180) );
  INVX2 U71 ( .A(B[11]), .Y(n15) );
  AND3X4 U72 ( .A(n50), .B(n3), .C(n179), .Y(n5) );
  NOR2X4 U73 ( .A(n180), .B(n181), .Y(n179) );
  NOR2X2 U74 ( .A(n131), .B(n22), .Y(n141) );
  NAND2BX2 U75 ( .AN(A[6]), .B(B[6]), .Y(n49) );
  NAND3XL U76 ( .A(n117), .B(n47), .C(n6), .Y(n159) );
  NOR2BX2 U77 ( .AN(B[7]), .B(A[7]), .Y(n181) );
  NAND4BX2 U78 ( .AN(n105), .B(n106), .C(n107), .D(n64), .Y(n93) );
  CLKINVX3 U79 ( .A(n91), .Y(n107) );
  INVX2 U80 ( .A(n162), .Y(n186) );
  NAND3BX2 U81 ( .AN(n131), .B(n54), .C(n140), .Y(n139) );
  INVXL U82 ( .A(A[11]), .Y(n9) );
  NAND2BX4 U83 ( .AN(B[7]), .B(A[7]), .Y(n47) );
  NOR2BX2 U84 ( .AN(n154), .B(n5), .Y(n150) );
  AOI21X4 U85 ( .A0(n2), .A1(n189), .B0(n190), .Y(n187) );
  NAND2X4 U86 ( .A(n191), .B(n192), .Y(n190) );
  NOR2X2 U87 ( .A(n112), .B(n113), .Y(n90) );
  NAND2X2 U88 ( .A(n67), .B(n21), .Y(n66) );
  NAND2BX4 U89 ( .AN(B[4]), .B(A[4]), .Y(n67) );
  CLKINVX3 U90 ( .A(n5), .Y(n6) );
  NAND2BX4 U91 ( .AN(n17), .B(n18), .Y(n19) );
  NAND2XL U92 ( .A(n103), .B(n104), .Y(n101) );
  NAND2BX2 U93 ( .AN(B[13]), .B(A[13]), .Y(n103) );
  INVX4 U94 ( .A(n28), .Y(n85) );
  NAND2BXL U95 ( .AN(B[15]), .B(A[15]), .Y(n96) );
  NOR2BXL U96 ( .AN(B[7]), .B(A[7]), .Y(n121) );
  NAND2X4 U97 ( .A(n29), .B(n27), .Y(n178) );
  NAND2XL U98 ( .A(n120), .B(n47), .Y(n119) );
  NOR2BX4 U99 ( .AN(n47), .B(n48), .Y(n46) );
  NAND3BX4 U100 ( .AN(n7), .B(n199), .C(n200), .Y(n63) );
  NAND2X4 U101 ( .A(n79), .B(n76), .Y(n7) );
  NOR2X4 U102 ( .A(n178), .B(n197), .Y(n177) );
  NAND2BX4 U103 ( .AN(A[5]), .B(B[5]), .Y(n52) );
  NAND2BX4 U104 ( .AN(B[9]), .B(A[9]), .Y(n169) );
  NAND2X4 U105 ( .A(n62), .B(n67), .Y(n50) );
  AOI21XL U106 ( .A0(n116), .A1(n117), .B0(n105), .Y(n112) );
  NAND2BX4 U107 ( .AN(A[1]), .B(B[1]), .Y(n199) );
  INVX1 U108 ( .A(n183), .Y(n8) );
  INVXL U109 ( .A(B[11]), .Y(n183) );
  NAND2XL U110 ( .A(n62), .B(n27), .Y(n69) );
  NAND2XL U111 ( .A(n38), .B(n40), .Y(n23) );
  NAND2BX4 U112 ( .AN(A[3]), .B(B[3]), .Y(n79) );
  OR2X2 U113 ( .A(n58), .B(n59), .Y(n24) );
  INVX4 U114 ( .A(n131), .Y(n134) );
  INVXL U115 ( .A(n107), .Y(n13) );
  AND2X2 U116 ( .A(n134), .B(n100), .Y(n14) );
  NAND2BX4 U117 ( .AN(B[5]), .B(A[5]), .Y(n62) );
  NAND3X2 U118 ( .A(n50), .B(n3), .C(n195), .Y(n191) );
  NAND3X2 U119 ( .A(n167), .B(n168), .C(B[9]), .Y(n166) );
  INVX4 U120 ( .A(n167), .Y(n176) );
  NAND2BX4 U121 ( .AN(B[10]), .B(A[10]), .Y(n167) );
  NOR2X2 U122 ( .A(n51), .B(n180), .Y(n42) );
  INVX4 U123 ( .A(n201), .Y(n78) );
  INVX3 U124 ( .A(n22), .Y(n133) );
  NOR2BXL U125 ( .AN(B[7]), .B(A[7]), .Y(n196) );
  NOR2X2 U126 ( .A(n176), .B(n186), .Y(n185) );
  NOR2X2 U127 ( .A(n153), .B(n105), .Y(n152) );
  NAND2BX4 U128 ( .AN(A[9]), .B(B[9]), .Y(n35) );
  INVX3 U129 ( .A(A[9]), .Y(n168) );
  NOR2X4 U130 ( .A(n149), .B(n153), .Y(n156) );
  NOR4BX4 U131 ( .AN(n63), .B(n64), .C(n65), .D(n66), .Y(n60) );
  INVX1 U132 ( .A(n103), .Y(n144) );
  NOR2X2 U133 ( .A(n141), .B(n128), .Y(n137) );
  INVX4 U134 ( .A(n194), .Y(n58) );
  XOR2X4 U135 ( .A(n69), .B(n70), .Y(DIFF[5]) );
  NAND2X4 U136 ( .A(n2), .B(n177), .Y(n151) );
  NOR3BX1 U137 ( .AN(n2), .B(n163), .C(n164), .Y(n160) );
  NAND2X4 U138 ( .A(n17), .B(n171), .Y(n20) );
  OAI21X4 U139 ( .A0(n174), .A1(n38), .B0(n175), .Y(n173) );
  XOR2X4 U140 ( .A(n124), .B(n123), .Y(DIFF[15]) );
  AOI21X4 U141 ( .A0(n172), .A1(n54), .B0(n173), .Y(n16) );
  AOI21X2 U142 ( .A0(n54), .A1(n172), .B0(n173), .Y(n171) );
  NOR2X2 U143 ( .A(n33), .B(n34), .Y(n32) );
  NAND2XL U144 ( .A(n79), .B(n21), .Y(n74) );
  NAND4X2 U145 ( .A(n76), .B(n79), .C(n87), .D(n199), .Y(n108) );
  INVX4 U146 ( .A(n102), .Y(n142) );
  NOR2X4 U147 ( .A(n174), .B(n182), .Y(n172) );
  NAND2X4 U148 ( .A(n162), .B(n35), .Y(n174) );
  NAND2BX4 U149 ( .AN(A[13]), .B(B[13]), .Y(n102) );
  INVX8 U150 ( .A(n117), .Y(n48) );
  NAND3X1 U151 ( .A(n100), .B(n101), .C(n102), .Y(n97) );
  NOR2X4 U152 ( .A(n85), .B(n81), .Y(n84) );
  NAND4BX4 U153 ( .AN(n161), .B(n162), .C(n35), .D(n40), .Y(n105) );
  NOR2X2 U154 ( .A(n131), .B(n132), .Y(n129) );
  OAI21X2 U155 ( .A0(n90), .A1(n13), .B0(n92), .Y(n88) );
  NAND4BX4 U156 ( .AN(n161), .B(n165), .C(n166), .D(n162), .Y(n114) );
  NAND2BX4 U157 ( .AN(A[8]), .B(B[8]), .Y(n40) );
  XNOR2X4 U158 ( .A(n54), .B(n23), .Y(DIFF[8]) );
  NAND2BX4 U159 ( .AN(B[8]), .B(A[8]), .Y(n38) );
  XOR2X2 U160 ( .A(n74), .B(n75), .Y(DIFF[3]) );
  AOI21X2 U161 ( .A0(n76), .A1(n77), .B0(n78), .Y(n75) );
  OAI21X4 U162 ( .A0(n80), .A1(n81), .B0(n28), .Y(n77) );
  INVX4 U163 ( .A(n199), .Y(n81) );
  NAND2BX4 U164 ( .AN(B[14]), .B(A[14]), .Y(n98) );
  XOR2X4 U165 ( .A(n55), .B(n56), .Y(DIFF[7]) );
  CLKINVX3 U166 ( .A(n108), .Y(n64) );
  NAND2X4 U167 ( .A(n20), .B(n19), .Y(DIFF[11]) );
  INVX4 U168 ( .A(n16), .Y(n18) );
  NAND2BX4 U169 ( .AN(B[12]), .B(A[12]), .Y(n104) );
  BUFX8 U170 ( .A(n68), .Y(n21) );
  NAND2BX1 U171 ( .AN(B[3]), .B(A[3]), .Y(n68) );
  XOR2X4 U172 ( .A(n31), .B(n32), .Y(DIFF[9]) );
  NAND2BX4 U173 ( .AN(A[10]), .B(B[10]), .Y(n162) );
  NAND2BX4 U174 ( .AN(A[4]), .B(B[4]), .Y(n53) );
  XOR2X4 U175 ( .A(n26), .B(n136), .Y(DIFF[14]) );
  AND3X4 U176 ( .A(n137), .B(n138), .C(n139), .Y(n26) );
  NAND2XL U177 ( .A(n98), .B(n100), .Y(n136) );
  XNOR2X4 U178 ( .A(n57), .B(n24), .Y(DIFF[6]) );
  OAI21X2 U179 ( .A0(n159), .A1(n160), .B0(n140), .Y(n158) );
  XNOR2X4 U180 ( .A(n25), .B(n143), .Y(DIFF[13]) );
  AND3X4 U181 ( .A(n145), .B(n146), .C(n147), .Y(n25) );
  NAND2XL U182 ( .A(n29), .B(n27), .Y(n198) );
  NAND2BX4 U183 ( .AN(A[15]), .B(B[15]), .Y(n111) );
  INVX1 U184 ( .A(n35), .Y(n34) );
  INVX1 U185 ( .A(n40), .Y(n182) );
  NAND2X1 U186 ( .A(n35), .B(n40), .Y(n188) );
  OAI21XL U187 ( .A0(A[7]), .A1(n39), .B0(n47), .Y(n55) );
  INVX1 U188 ( .A(n98), .Y(n130) );
  NAND2X1 U189 ( .A(n96), .B(n111), .Y(n123) );
  NOR2X2 U190 ( .A(n197), .B(n198), .Y(n189) );
  OAI2BB1X2 U191 ( .A0N(n150), .A1N(n151), .B0(n152), .Y(n146) );
  INVX1 U192 ( .A(n96), .Y(n95) );
  AOI21X1 U193 ( .A0(n97), .A1(n98), .B0(n99), .Y(n94) );
  INVX1 U194 ( .A(n104), .Y(n149) );
  NAND2XL U195 ( .A(n3), .B(n4), .Y(n164) );
  INVX1 U196 ( .A(n83), .Y(n80) );
  NAND3XL U197 ( .A(n21), .B(n122), .C(n63), .Y(n118) );
  XOR2X2 U198 ( .A(n83), .B(n84), .Y(DIFF[1]) );
  XOR2X2 U199 ( .A(n88), .B(n89), .Y(DIFF[16]) );
  XNOR2X1 U200 ( .A(B[16]), .B(A[16]), .Y(n89) );
  NAND2X1 U201 ( .A(n86), .B(n87), .Y(DIFF[0]) );
  NAND2BX1 U202 ( .AN(n87), .B(n86), .Y(n83) );
  NAND2BX1 U203 ( .AN(B[0]), .B(A[0]), .Y(n86) );
  NAND2BX1 U204 ( .AN(A[0]), .B(B[0]), .Y(n87) );
  OAI21XL U205 ( .A0(A[7]), .A1(n39), .B0(n53), .Y(n163) );
  NOR2BX1 U206 ( .AN(n47), .B(n48), .Y(n154) );
  NAND2XL U207 ( .A(n114), .B(n22), .Y(n113) );
  AOI21X4 U208 ( .A0(n3), .A1(n57), .B0(n58), .Y(n56) );
  OAI21X4 U209 ( .A0(n60), .A1(n61), .B0(n62), .Y(n57) );
  AOI211X2 U210 ( .A0(n128), .A1(n100), .B0(n129), .C0(n130), .Y(n127) );
  NAND2BX4 U211 ( .AN(A[14]), .B(B[14]), .Y(n100) );
  NAND2X4 U212 ( .A(n110), .B(n102), .Y(n131) );
  XOR2X4 U213 ( .A(n155), .B(n156), .Y(DIFF[12]) );
  NAND2BX4 U214 ( .AN(A[12]), .B(B[12]), .Y(n110) );
  NAND2BX4 U215 ( .AN(n157), .B(n158), .Y(n155) );
  NAND4BX4 U216 ( .AN(n48), .B(n120), .C(n47), .D(n151), .Y(n54) );
  NAND3X4 U217 ( .A(n50), .B(n3), .C(n179), .Y(n120) );
  XOR2X4 U218 ( .A(n184), .B(n185), .Y(DIFF[10]) );
  OAI21X4 U219 ( .A0(n187), .A1(n188), .B0(n169), .Y(n184) );
  OAI2BB1X4 U220 ( .A0N(n30), .A1N(B[7]), .B0(n58), .Y(n117) );
endmodule


module butterfly_DW01_add_123 ( A, B, SUM );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146;

  NOR2BX1 U2 ( .AN(n126), .B(n133), .Y(n141) );
  INVX4 U3 ( .A(n125), .Y(n133) );
  NAND2X2 U4 ( .A(n22), .B(n20), .Y(n124) );
  CLKINVX8 U5 ( .A(n90), .Y(n122) );
  AOI21X4 U6 ( .A0(n17), .A1(n18), .B0(n19), .Y(n16) );
  BUFX8 U7 ( .A(n51), .Y(n1) );
  XNOR2X2 U8 ( .A(B[16]), .B(A[16]), .Y(n8) );
  INVX4 U9 ( .A(n18), .Y(n24) );
  NAND2X2 U10 ( .A(n42), .B(n43), .Y(n37) );
  NOR2BX2 U11 ( .AN(n27), .B(n28), .Y(n26) );
  INVX1 U12 ( .A(n107), .Y(n112) );
  NOR2X1 U13 ( .A(n80), .B(n81), .Y(n76) );
  NOR2BX2 U14 ( .AN(n36), .B(n47), .Y(n49) );
  INVX2 U15 ( .A(n35), .Y(n41) );
  INVX1 U16 ( .A(n20), .Y(n19) );
  NAND2BX2 U17 ( .AN(n126), .B(n12), .Y(n94) );
  OAI21X1 U18 ( .A0(n50), .A1(n1), .B0(n54), .Y(n129) );
  CLKINVX3 U19 ( .A(n137), .Y(n136) );
  OR2X2 U20 ( .A(A[6]), .B(B[6]), .Y(n34) );
  NOR2BX1 U21 ( .AN(n79), .B(n80), .Y(n116) );
  NOR2BX1 U22 ( .AN(n78), .B(n86), .Y(n111) );
  INVX1 U23 ( .A(n109), .Y(n14) );
  INVX1 U24 ( .A(n78), .Y(n108) );
  INVX1 U25 ( .A(n43), .Y(n47) );
  NAND2X1 U26 ( .A(n37), .B(n36), .Y(n40) );
  OR2X2 U27 ( .A(A[6]), .B(B[6]), .Y(n5) );
  NAND2X1 U28 ( .A(B[7]), .B(A[7]), .Y(n27) );
  AND2X2 U29 ( .A(n37), .B(n10), .Y(n30) );
  NAND2X2 U30 ( .A(B[8]), .B(A[8]), .Y(n20) );
  OR2X2 U31 ( .A(A[8]), .B(B[8]), .Y(n18) );
  NOR2X1 U32 ( .A(n80), .B(n87), .Y(n83) );
  OAI21XL U33 ( .A0(n71), .A1(n72), .B0(n73), .Y(n70) );
  INVX1 U34 ( .A(n57), .Y(n55) );
  XOR2X1 U35 ( .A(n60), .B(n62), .Y(SUM[1]) );
  NOR2X1 U36 ( .A(A[3]), .B(B[3]), .Y(n2) );
  NAND2X1 U37 ( .A(B[11]), .B(A[11]), .Y(n3) );
  NAND2X2 U38 ( .A(B[9]), .B(A[9]), .Y(n22) );
  NAND2X1 U39 ( .A(B[6]), .B(A[6]), .Y(n32) );
  NAND2XL U40 ( .A(n21), .B(n22), .Y(n15) );
  AND2X4 U41 ( .A(n99), .B(n27), .Y(n143) );
  INVX1 U42 ( .A(n27), .Y(n100) );
  OAI2BB1X4 U43 ( .A0N(n69), .A1N(n119), .B0(n120), .Y(n4) );
  OR2X4 U44 ( .A(A[11]), .B(B[11]), .Y(n12) );
  CLKINVX4 U45 ( .A(n98), .Y(n69) );
  INVX8 U46 ( .A(n33), .Y(n46) );
  NAND2X1 U47 ( .A(B[15]), .B(A[15]), .Y(n73) );
  OR2X2 U48 ( .A(B[15]), .B(A[15]), .Y(n75) );
  NAND2X2 U49 ( .A(n99), .B(n27), .Y(n138) );
  XOR2X2 U50 ( .A(n117), .B(n118), .Y(SUM[12]) );
  OAI2BB1X2 U51 ( .A0N(n117), .A1N(n14), .B0(n112), .Y(n110) );
  NAND2X4 U52 ( .A(B[5]), .B(A[5]), .Y(n35) );
  OR2X2 U53 ( .A(A[7]), .B(B[7]), .Y(n11) );
  NAND2X2 U54 ( .A(B[3]), .B(A[3]), .Y(n54) );
  NAND3BX4 U55 ( .AN(n138), .B(n127), .C(n95), .Y(n135) );
  XOR2X4 U56 ( .A(n102), .B(n103), .Y(SUM[15]) );
  AND2X2 U57 ( .A(n35), .B(n36), .Y(n10) );
  NOR2BX2 U58 ( .AN(n35), .B(n46), .Y(n45) );
  OR2X4 U59 ( .A(A[4]), .B(B[4]), .Y(n43) );
  NOR2BX1 U60 ( .AN(n61), .B(n63), .Y(n62) );
  XNOR2X4 U61 ( .A(n65), .B(n8), .Y(SUM[16]) );
  OAI21X2 U62 ( .A0(n66), .A1(n67), .B0(n68), .Y(n65) );
  NAND2X2 U63 ( .A(n21), .B(n18), .Y(n139) );
  NAND2X4 U64 ( .A(A[1]), .B(B[1]), .Y(n61) );
  OR2X2 U65 ( .A(A[14]), .B(B[14]), .Y(n74) );
  AND2X2 U66 ( .A(n3), .B(n12), .Y(n7) );
  AND3X4 U67 ( .A(n142), .B(n95), .C(n143), .Y(n6) );
  NAND2BXL U68 ( .AN(n82), .B(n101), .Y(n96) );
  NAND2X1 U69 ( .A(B[13]), .B(A[13]), .Y(n79) );
  NAND2BX4 U70 ( .AN(n82), .B(n129), .Y(n127) );
  NAND2X2 U71 ( .A(n113), .B(n114), .Y(n109) );
  INVX3 U72 ( .A(n113), .Y(n87) );
  OR2X1 U73 ( .A(A[12]), .B(B[12]), .Y(n113) );
  NAND3X2 U74 ( .A(A[6]), .B(B[6]), .C(n29), .Y(n95) );
  AOI21X4 U75 ( .A0(n134), .A1(n135), .B0(n136), .Y(n132) );
  OAI21X4 U76 ( .A0(n6), .A1(n139), .B0(n137), .Y(n140) );
  NOR2BX4 U77 ( .AN(n54), .B(n2), .Y(n53) );
  XOR2X2 U78 ( .A(n57), .B(n58), .Y(SUM[2]) );
  XOR2X4 U79 ( .A(n17), .B(n23), .Y(SUM[8]) );
  NAND2X2 U80 ( .A(B[14]), .B(A[14]), .Y(n78) );
  NOR2BX4 U81 ( .AN(n81), .B(n87), .Y(n118) );
  NAND2X2 U82 ( .A(B[10]), .B(A[10]), .Y(n126) );
  OAI21X4 U83 ( .A0(n104), .A1(n87), .B0(n81), .Y(n115) );
  OAI21X2 U84 ( .A0(n80), .A1(n81), .B0(n79), .Y(n107) );
  NAND2X2 U85 ( .A(B[12]), .B(A[12]), .Y(n81) );
  NAND2X1 U86 ( .A(n78), .B(n79), .Y(n77) );
  OAI21X2 U87 ( .A0(n55), .A1(n13), .B0(n56), .Y(n52) );
  NOR2BX2 U88 ( .AN(n56), .B(n13), .Y(n58) );
  NOR2X1 U89 ( .A(A[2]), .B(B[2]), .Y(n13) );
  XOR2X2 U90 ( .A(n42), .B(n49), .Y(SUM[4]) );
  INVX8 U91 ( .A(n114), .Y(n80) );
  OR2X4 U92 ( .A(A[13]), .B(B[13]), .Y(n114) );
  NAND3X4 U93 ( .A(n12), .B(n125), .C(n130), .Y(n98) );
  OR2X4 U94 ( .A(A[10]), .B(B[10]), .Y(n125) );
  AOI21X4 U95 ( .A0(B[2]), .A1(A[2]), .B0(n146), .Y(n50) );
  INVX4 U96 ( .A(n74), .Y(n86) );
  NAND2X4 U97 ( .A(B[0]), .B(A[0]), .Y(n64) );
  AOI21X2 U98 ( .A0(n40), .A1(n33), .B0(n41), .Y(n39) );
  NOR2XL U99 ( .A(n85), .B(n86), .Y(n84) );
  INVXL U100 ( .A(n94), .Y(n93) );
  INVX2 U101 ( .A(n139), .Y(n134) );
  NAND3BX2 U102 ( .AN(n138), .B(n127), .C(n128), .Y(n119) );
  XOR2X4 U103 ( .A(n131), .B(n7), .Y(SUM[11]) );
  OAI21X4 U104 ( .A0(n30), .A1(n31), .B0(n32), .Y(n25) );
  XOR2X4 U105 ( .A(n115), .B(n116), .Y(SUM[13]) );
  NOR2BX1 U106 ( .AN(n64), .B(n9), .Y(SUM[0]) );
  NOR2XL U107 ( .A(A[0]), .B(B[0]), .Y(n9) );
  OR2X2 U108 ( .A(n86), .B(n109), .Y(n105) );
  NAND2X1 U109 ( .A(n83), .B(n84), .Y(n67) );
  NOR2BX2 U110 ( .AN(n20), .B(n24), .Y(n23) );
  NAND2XL U111 ( .A(n5), .B(n32), .Y(n38) );
  INVXL U112 ( .A(n29), .Y(n28) );
  NOR2BX1 U113 ( .AN(n73), .B(n85), .Y(n103) );
  OAI21X2 U114 ( .A0(n104), .A1(n105), .B0(n106), .Y(n102) );
  AOI21X1 U115 ( .A0(n107), .A1(n74), .B0(n108), .Y(n106) );
  OAI2BB1X2 U116 ( .A0N(n22), .A1N(n20), .B0(n21), .Y(n137) );
  XOR2X2 U117 ( .A(n52), .B(n53), .Y(SUM[3]) );
  INVX1 U118 ( .A(n75), .Y(n85) );
  OAI2BB1X1 U119 ( .A0N(n59), .A1N(n60), .B0(n61), .Y(n57) );
  NOR2X1 U120 ( .A(n88), .B(n89), .Y(n66) );
  NAND2XL U121 ( .A(n90), .B(n91), .Y(n89) );
  AOI31X1 U122 ( .A0(n95), .A1(n96), .A2(n97), .B0(n98), .Y(n88) );
  NOR2X1 U123 ( .A(n92), .B(n93), .Y(n91) );
  NOR2X1 U124 ( .A(n76), .B(n77), .Y(n71) );
  NAND2X1 U125 ( .A(n74), .B(n75), .Y(n72) );
  INVX1 U126 ( .A(n64), .Y(n60) );
  NAND2XL U127 ( .A(n33), .B(n34), .Y(n31) );
  INVXL U128 ( .A(n3), .Y(n92) );
  OAI21XL U129 ( .A0(n50), .A1(n1), .B0(n54), .Y(n101) );
  NAND4X2 U130 ( .A(n11), .B(n43), .C(n33), .D(n34), .Y(n82) );
  NAND2XL U131 ( .A(B[2]), .B(A[2]), .Y(n56) );
  INVX1 U132 ( .A(n70), .Y(n68) );
  OAI22X2 U133 ( .A0(A[2]), .A1(B[2]), .B0(A[3]), .B1(B[3]), .Y(n51) );
  NAND3XL U134 ( .A(A[6]), .B(B[6]), .C(n29), .Y(n128) );
  INVX8 U135 ( .A(n21), .Y(n123) );
  INVX2 U136 ( .A(n42), .Y(n48) );
  NOR2X4 U137 ( .A(n24), .B(n123), .Y(n130) );
  NOR2BX1 U138 ( .AN(n99), .B(n100), .Y(n97) );
  INVX8 U139 ( .A(n4), .Y(n104) );
  XOR2X4 U140 ( .A(n16), .B(n15), .Y(SUM[9]) );
  XOR2X4 U141 ( .A(n25), .B(n26), .Y(SUM[7]) );
  XOR2X4 U142 ( .A(n38), .B(n39), .Y(SUM[6]) );
  XOR2X4 U143 ( .A(n44), .B(n45), .Y(SUM[5]) );
  OAI21X4 U144 ( .A0(n47), .A1(n48), .B0(n36), .Y(n44) );
  OAI21X4 U145 ( .A0(n50), .A1(n1), .B0(n54), .Y(n42) );
  XOR2X4 U146 ( .A(n110), .B(n111), .Y(SUM[14]) );
  OAI2BB1X4 U147 ( .A0N(n69), .A1N(n119), .B0(n120), .Y(n117) );
  NOR2X4 U148 ( .A(n121), .B(n122), .Y(n120) );
  NAND4BX4 U149 ( .AN(n123), .B(n124), .C(n12), .D(n125), .Y(n90) );
  NAND2X4 U150 ( .A(n94), .B(n3), .Y(n121) );
  OAI21X4 U151 ( .A0(n132), .A1(n133), .B0(n126), .Y(n131) );
  XOR2X4 U152 ( .A(n140), .B(n141), .Y(SUM[10]) );
  OR2X4 U153 ( .A(A[9]), .B(B[9]), .Y(n21) );
  NAND3X4 U154 ( .A(n142), .B(n95), .C(n143), .Y(n17) );
  NAND2BX4 U155 ( .AN(n144), .B(n145), .Y(n99) );
  AOI21X4 U156 ( .A0(n35), .A1(n36), .B0(n46), .Y(n145) );
  NAND2X4 U157 ( .A(B[4]), .B(A[4]), .Y(n36) );
  NAND2X4 U158 ( .A(n5), .B(n29), .Y(n144) );
  OR2X4 U159 ( .A(A[7]), .B(B[7]), .Y(n29) );
  NAND2BX4 U160 ( .AN(n82), .B(n129), .Y(n142) );
  OAI21X4 U161 ( .A0(n64), .A1(n63), .B0(n61), .Y(n146) );
  CLKINVX3 U162 ( .A(n59), .Y(n63) );
  OR2X4 U163 ( .A(B[1]), .B(A[1]), .Y(n59) );
  OR2X4 U164 ( .A(B[5]), .B(A[5]), .Y(n33) );
endmodule


module butterfly_DW01_sub_100 ( A, B, DIFF );
  input [16:0] A;
  input [16:0] B;
  output [16:0] DIFF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199;

  AOI21X2 U3 ( .A0(n155), .A1(n156), .B0(n157), .Y(n154) );
  OAI21X4 U4 ( .A0(n140), .A1(n118), .B0(n158), .Y(n157) );
  AOI2BB1X4 U5 ( .A0N(n42), .A1N(n41), .B0(n199), .Y(n197) );
  INVX3 U6 ( .A(n31), .Y(n30) );
  NAND2BX2 U7 ( .AN(B[13]), .B(A[13]), .Y(n132) );
  NOR2X4 U8 ( .A(n112), .B(n113), .Y(n111) );
  AOI21X4 U9 ( .A0(n114), .A1(n115), .B0(n97), .Y(n113) );
  OAI2BB1X4 U10 ( .A0N(n171), .A1N(A[9]), .B0(n172), .Y(n162) );
  CLKINVX1 U11 ( .A(B[9]), .Y(n171) );
  NAND2BX2 U12 ( .AN(B[8]), .B(A[8]), .Y(n172) );
  NAND2BX4 U13 ( .AN(B[8]), .B(A[8]), .Y(n139) );
  NOR2BX2 U14 ( .AN(n101), .B(n144), .Y(n164) );
  CLKINVX3 U15 ( .A(n44), .Y(n144) );
  NAND4X4 U16 ( .A(n14), .B(n13), .C(n39), .D(n6), .Y(n183) );
  BUFX20 U17 ( .A(n123), .Y(n1) );
  CLKINVX8 U18 ( .A(n4), .Y(n6) );
  XOR2X2 U19 ( .A(B[16]), .B(A[16]), .Y(n75) );
  NOR2X2 U20 ( .A(n193), .B(n192), .Y(n191) );
  OAI21X2 U21 ( .A0(n84), .A1(n85), .B0(n132), .Y(n131) );
  AND2X1 U22 ( .A(n39), .B(n50), .Y(n11) );
  NAND2X2 U23 ( .A(n122), .B(n1), .Y(n8) );
  INVX2 U24 ( .A(n24), .Y(n186) );
  NAND3X1 U25 ( .A(n163), .B(n100), .C(n164), .Y(n153) );
  NAND3X2 U26 ( .A(n190), .B(n58), .C(n191), .Y(n103) );
  NOR2X2 U27 ( .A(n194), .B(n16), .Y(n15) );
  OAI21X2 U28 ( .A0(n85), .A1(n119), .B0(n120), .Y(n112) );
  AOI21X2 U29 ( .A0(n87), .A1(n121), .B0(n88), .Y(n120) );
  INVX1 U30 ( .A(A[11]), .Y(n3) );
  AOI21X2 U31 ( .A0(n183), .A1(n188), .B0(n189), .Y(n187) );
  NAND3X2 U32 ( .A(n118), .B(n133), .C(n115), .Y(n105) );
  OAI21X1 U33 ( .A0(n65), .A1(n66), .B0(n67), .Y(n59) );
  NAND2X2 U34 ( .A(n37), .B(n49), .Y(n47) );
  INVX1 U35 ( .A(n27), .Y(n19) );
  AOI21X1 U36 ( .A0(n81), .A1(n82), .B0(n83), .Y(n80) );
  OAI21XL U37 ( .A0(n84), .A1(n85), .B0(n86), .Y(n82) );
  NOR2X2 U38 ( .A(n88), .B(n90), .Y(n125) );
  XOR2X2 U39 ( .A(n52), .B(n53), .Y(DIFF[5]) );
  XOR2X1 U40 ( .A(n68), .B(n69), .Y(DIFF[1]) );
  NOR2X1 U41 ( .A(n70), .B(n66), .Y(n69) );
  INVX1 U42 ( .A(n67), .Y(n70) );
  NOR2X1 U43 ( .A(n55), .B(n41), .Y(n54) );
  INVX1 U44 ( .A(n50), .Y(n55) );
  AOI21X2 U45 ( .A0(n36), .A1(n37), .B0(n38), .Y(n35) );
  INVX1 U46 ( .A(n7), .Y(n2) );
  NAND2X1 U47 ( .A(n39), .B(n7), .Y(n52) );
  BUFX3 U48 ( .A(n48), .Y(n7) );
  INVX4 U49 ( .A(n133), .Y(n116) );
  INVX1 U50 ( .A(n194), .Y(n60) );
  INVX1 U51 ( .A(n135), .Y(n160) );
  INVX1 U52 ( .A(A[9]), .Y(n138) );
  CLKINVXL U53 ( .A(n99), .Y(n91) );
  NAND2BXL U54 ( .AN(n97), .B(n96), .Y(n78) );
  INVX4 U55 ( .A(n170), .Y(n141) );
  NAND2X1 U56 ( .A(n122), .B(n121), .Y(n119) );
  NAND2BX2 U57 ( .AN(B[9]), .B(A[9]), .Y(n24) );
  NAND4X2 U58 ( .A(n71), .B(n73), .C(n61), .D(n58), .Y(n93) );
  NAND2BX1 U59 ( .AN(B[6]), .B(A[6]), .Y(n51) );
  NAND2BX2 U60 ( .AN(A[6]), .B(B[6]), .Y(n148) );
  NAND2BX1 U61 ( .AN(A[15]), .B(B[15]), .Y(n96) );
  NAND2X1 U62 ( .A(n39), .B(n40), .Y(n38) );
  NAND2X1 U63 ( .A(n39), .B(n50), .Y(n147) );
  NOR2BX1 U64 ( .AN(B[5]), .B(A[5]), .Y(n199) );
  NOR2BX2 U65 ( .AN(n136), .B(n161), .Y(n155) );
  NAND3X1 U66 ( .A(n100), .B(n44), .C(n101), .Y(n31) );
  OAI21X1 U67 ( .A0(B[9]), .A1(n138), .B0(n139), .Y(n137) );
  NAND2BX4 U68 ( .AN(A[10]), .B(B[10]), .Y(n135) );
  NAND2BX1 U69 ( .AN(B[14]), .B(A[14]), .Y(n126) );
  NOR2BX2 U70 ( .AN(n101), .B(n144), .Y(n175) );
  AOI21X4 U71 ( .A0(n116), .A1(n1), .B0(n159), .Y(n158) );
  AOI21X4 U72 ( .A0(n47), .A1(n39), .B0(n2), .Y(n46) );
  NOR2X2 U73 ( .A(n99), .B(n97), .Y(n109) );
  NOR2BX2 U74 ( .AN(n101), .B(n144), .Y(n143) );
  NAND2BX1 U75 ( .AN(B[3]), .B(A[3]), .Y(n62) );
  NOR2BX2 U76 ( .AN(B[3]), .B(A[3]), .Y(n193) );
  AND2X2 U77 ( .A(n43), .B(n148), .Y(n14) );
  NAND2X1 U78 ( .A(n43), .B(n1), .Y(n166) );
  CLKINVX4 U79 ( .A(n8), .Y(n9) );
  NAND2BX4 U80 ( .AN(B[4]), .B(A[4]), .Y(n49) );
  INVX8 U81 ( .A(n49), .Y(n41) );
  NAND3BX2 U82 ( .AN(n182), .B(n27), .C(n22), .Y(n180) );
  NOR2X4 U83 ( .A(n76), .B(n77), .Y(n74) );
  AOI21X2 U84 ( .A0(n94), .A1(n95), .B0(n78), .Y(n76) );
  INVX4 U85 ( .A(n96), .Y(n89) );
  NAND2BX2 U86 ( .AN(B[7]), .B(A[7]), .Y(n44) );
  NAND2XL U87 ( .A(n135), .B(n173), .Y(n184) );
  OAI21X1 U88 ( .A0(n182), .A1(n24), .B0(n173), .Y(n179) );
  INVX4 U89 ( .A(n118), .Y(n117) );
  NAND2BX4 U90 ( .AN(A[2]), .B(B[2]), .Y(n58) );
  NOR2BX2 U91 ( .AN(B[1]), .B(A[1]), .Y(n192) );
  NAND2BX4 U92 ( .AN(n182), .B(n21), .Y(n181) );
  NAND2XL U93 ( .A(n23), .B(n27), .Y(n189) );
  NAND2BX2 U94 ( .AN(A[6]), .B(B[6]), .Y(n40) );
  INVX2 U95 ( .A(n61), .Y(n16) );
  INVX3 U96 ( .A(n101), .Y(n195) );
  NAND2BX2 U97 ( .AN(A[1]), .B(B[1]), .Y(n71) );
  NAND2BX2 U98 ( .AN(B[10]), .B(A[10]), .Y(n173) );
  OR2X4 U99 ( .A(B[11]), .B(n3), .Y(n133) );
  XOR2X4 U100 ( .A(n45), .B(n46), .Y(DIFF[6]) );
  NOR2X4 U101 ( .A(n116), .B(n117), .Y(n114) );
  INVX4 U102 ( .A(n126), .Y(n88) );
  INVX4 U103 ( .A(n1), .Y(n140) );
  NAND2X2 U104 ( .A(n1), .B(n85), .Y(n167) );
  NOR3BX4 U105 ( .AN(n1), .B(n84), .C(n141), .Y(n129) );
  NAND2X2 U106 ( .A(n1), .B(n122), .Y(n149) );
  NAND3X2 U107 ( .A(n142), .B(n100), .C(n143), .Y(n110) );
  AOI21X4 U108 ( .A0(n130), .A1(n129), .B0(n131), .Y(n128) );
  OAI2BB1X4 U109 ( .A0N(n28), .A1N(n6), .B0(n30), .Y(n25) );
  NOR2X2 U110 ( .A(n149), .B(n99), .Y(n127) );
  NAND3X4 U111 ( .A(n100), .B(n44), .C(n101), .Y(n22) );
  NAND2XL U112 ( .A(n23), .B(n24), .Y(n17) );
  NOR2X2 U113 ( .A(n87), .B(n88), .Y(n86) );
  OAI21X2 U114 ( .A0(n78), .A1(n79), .B0(n80), .Y(n77) );
  INVX4 U115 ( .A(n22), .Y(n20) );
  OAI2BB1X4 U116 ( .A0N(n110), .A1N(n109), .B0(n111), .Y(n106) );
  OAI2BB1X4 U117 ( .A0N(n152), .A1N(n153), .B0(n154), .Y(n150) );
  NAND2BX2 U118 ( .AN(A[9]), .B(B[9]), .Y(n136) );
  NOR2BX1 U119 ( .AN(B[9]), .B(A[9]), .Y(n176) );
  NAND2XL U120 ( .A(n40), .B(n51), .Y(n45) );
  NAND2BX2 U121 ( .AN(A[9]), .B(B[9]), .Y(n23) );
  INVX1 U122 ( .A(n58), .Y(n64) );
  NAND2BX2 U123 ( .AN(B[2]), .B(A[2]), .Y(n194) );
  AOI21XL U124 ( .A0(n58), .A1(n59), .B0(n60), .Y(n57) );
  NAND3X2 U125 ( .A(n118), .B(n133), .C(n134), .Y(n130) );
  INVX4 U126 ( .A(n71), .Y(n66) );
  NAND2X4 U127 ( .A(n12), .B(n100), .Y(n196) );
  NAND2BX4 U128 ( .AN(A[5]), .B(B[5]), .Y(n39) );
  AND2X4 U129 ( .A(n50), .B(n27), .Y(n13) );
  XNOR2X4 U130 ( .A(n25), .B(n10), .Y(DIFF[8]) );
  AND2X4 U131 ( .A(n172), .B(n44), .Y(n12) );
  NAND2XL U132 ( .A(n148), .B(n43), .Y(n146) );
  NAND2XL U133 ( .A(n43), .B(n44), .Y(n32) );
  XOR2X2 U134 ( .A(n6), .B(n54), .Y(DIFF[4]) );
  NOR2X4 U135 ( .A(n195), .B(n196), .Y(n188) );
  OAI2BB1X4 U136 ( .A0N(n127), .A1N(n110), .B0(n128), .Y(n124) );
  NAND3X1 U137 ( .A(n135), .B(n136), .C(n137), .Y(n134) );
  INVX4 U138 ( .A(n121), .Y(n90) );
  NAND2X4 U139 ( .A(n9), .B(n121), .Y(n97) );
  NAND2BX4 U140 ( .AN(A[14]), .B(B[14]), .Y(n121) );
  NOR2X2 U141 ( .A(n116), .B(n141), .Y(n178) );
  NOR3X4 U142 ( .A(n140), .B(n160), .C(n141), .Y(n156) );
  NAND2BX2 U143 ( .AN(B[1]), .B(A[1]), .Y(n67) );
  AOI21X2 U144 ( .A0(n5), .A1(n50), .B0(n41), .Y(n53) );
  NAND2X4 U145 ( .A(n183), .B(n139), .Y(n21) );
  INVX2 U146 ( .A(n85), .Y(n159) );
  INVX8 U147 ( .A(n122), .Y(n84) );
  NAND2BX4 U148 ( .AN(A[13]), .B(B[13]), .Y(n122) );
  CLKINVX8 U149 ( .A(n29), .Y(n4) );
  INVX8 U150 ( .A(n4), .Y(n5) );
  NAND2XL U151 ( .A(n6), .B(n165), .Y(n163) );
  NAND2XL U152 ( .A(n6), .B(n145), .Y(n142) );
  NAND2BXL U153 ( .AN(n92), .B(n6), .Y(n174) );
  NAND2BX2 U154 ( .AN(B[5]), .B(A[5]), .Y(n48) );
  NAND2BX4 U155 ( .AN(A[7]), .B(B[7]), .Y(n43) );
  NAND4X2 U156 ( .A(n43), .B(n50), .C(n148), .D(n39), .Y(n92) );
  NAND3BX4 U157 ( .AN(n179), .B(n180), .C(n181), .Y(n177) );
  NAND2BX4 U158 ( .AN(A[3]), .B(B[3]), .Y(n61) );
  INVX4 U159 ( .A(n132), .Y(n87) );
  NAND4X2 U160 ( .A(n170), .B(n162), .C(n136), .D(n135), .Y(n115) );
  NAND2BX4 U161 ( .AN(A[11]), .B(B[11]), .Y(n170) );
  AND2X4 U162 ( .A(n43), .B(n40), .Y(n198) );
  XOR2X4 U163 ( .A(n124), .B(n125), .Y(DIFF[14]) );
  NAND2BX4 U164 ( .AN(A[8]), .B(B[8]), .Y(n27) );
  INVX4 U165 ( .A(n51), .Y(n34) );
  NAND4BX4 U166 ( .AN(n176), .B(n170), .C(n135), .D(n27), .Y(n99) );
  XOR2X4 U167 ( .A(n106), .B(n107), .Y(DIFF[15]) );
  XOR2X2 U168 ( .A(n56), .B(n57), .Y(DIFF[3]) );
  XOR2X4 U169 ( .A(n150), .B(n151), .Y(DIFF[13]) );
  NAND2X4 U170 ( .A(n34), .B(n43), .Y(n100) );
  NAND2BX4 U171 ( .AN(n173), .B(n170), .Y(n118) );
  NOR2X1 U172 ( .A(n60), .B(n64), .Y(n63) );
  NAND3BXL U173 ( .AN(n93), .B(n28), .C(n91), .Y(n79) );
  CLKINVX3 U174 ( .A(n92), .Y(n28) );
  INVX4 U175 ( .A(n48), .Y(n42) );
  INVXL U176 ( .A(n105), .Y(n94) );
  INVXL U177 ( .A(n162), .Y(n161) );
  NOR2X2 U178 ( .A(n166), .B(n99), .Y(n152) );
  NAND2BX4 U179 ( .AN(A[4]), .B(B[4]), .Y(n50) );
  OR2X2 U180 ( .A(n26), .B(n19), .Y(n10) );
  AND2X1 U181 ( .A(n11), .B(n148), .Y(n165) );
  NAND2BXL U182 ( .AN(B[15]), .B(A[15]), .Y(n108) );
  NOR2X1 U183 ( .A(n41), .B(n42), .Y(n36) );
  INVXL U184 ( .A(n139), .Y(n26) );
  NOR2X2 U185 ( .A(n146), .B(n147), .Y(n145) );
  XOR2X1 U186 ( .A(n59), .B(n63), .Y(DIFF[2]) );
  NAND2X1 U187 ( .A(n61), .B(n62), .Y(n56) );
  NOR2XL U188 ( .A(n89), .B(n90), .Y(n81) );
  OAI21XL U189 ( .A0(n98), .A1(n31), .B0(n91), .Y(n95) );
  INVX1 U190 ( .A(n68), .Y(n65) );
  AOI21XL U191 ( .A0(n102), .A1(n103), .B0(n92), .Y(n98) );
  INVXL U192 ( .A(n62), .Y(n104) );
  NAND2X2 U193 ( .A(n67), .B(n72), .Y(n190) );
  NAND2X1 U194 ( .A(n72), .B(n73), .Y(DIFF[0]) );
  NAND2BX1 U195 ( .AN(n73), .B(n72), .Y(n68) );
  NAND2BX1 U196 ( .AN(B[0]), .B(A[0]), .Y(n72) );
  NAND2BX1 U197 ( .AN(A[0]), .B(B[0]), .Y(n73) );
  NOR2X1 U198 ( .A(n104), .B(n15), .Y(n102) );
  XOR2X4 U199 ( .A(n18), .B(n17), .Y(DIFF[9]) );
  AOI2BB1X4 U200 ( .A0N(n19), .A1N(n20), .B0(n21), .Y(n18) );
  XOR2X4 U201 ( .A(n32), .B(n33), .Y(DIFF[7]) );
  NOR2X4 U202 ( .A(n34), .B(n35), .Y(n33) );
  NAND2X4 U203 ( .A(n5), .B(n50), .Y(n37) );
  XOR2X4 U204 ( .A(n74), .B(n75), .Y(DIFF[16]) );
  NOR2X4 U205 ( .A(n89), .B(n83), .Y(n107) );
  CLKINVX3 U206 ( .A(n108), .Y(n83) );
  NOR2X4 U207 ( .A(n87), .B(n84), .Y(n151) );
  XOR2X4 U208 ( .A(n168), .B(n167), .Y(DIFF[12]) );
  NOR2X4 U209 ( .A(n169), .B(n105), .Y(n168) );
  AOI31X2 U210 ( .A0(n174), .A1(n100), .A2(n175), .B0(n99), .Y(n169) );
  NAND2BX4 U211 ( .AN(B[12]), .B(A[12]), .Y(n85) );
  NAND2BX4 U212 ( .AN(A[12]), .B(B[12]), .Y(n123) );
  XOR2X4 U213 ( .A(n177), .B(n178), .Y(DIFF[11]) );
  NAND2X4 U214 ( .A(n135), .B(n23), .Y(n182) );
  XOR2X4 U215 ( .A(n185), .B(n184), .Y(DIFF[10]) );
  NOR2X4 U216 ( .A(n187), .B(n186), .Y(n185) );
  NAND4BX4 U217 ( .AN(n15), .B(n93), .C(n103), .D(n62), .Y(n29) );
  NAND2X4 U218 ( .A(n198), .B(n197), .Y(n101) );
endmodule


module butterfly_DW01_sub_98 ( A, B, DIFF );
  input [16:0] A;
  input [16:0] B;
  output [16:0] DIFF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175;

  OR2X2 U3 ( .A(n66), .B(n68), .Y(n16) );
  AND2X4 U4 ( .A(n55), .B(n56), .Y(n170) );
  INVX2 U5 ( .A(n99), .Y(n120) );
  BUFX8 U6 ( .A(n47), .Y(n12) );
  INVX1 U7 ( .A(n59), .Y(n9) );
  NAND2X2 U8 ( .A(n149), .B(n1), .Y(n147) );
  AND2X2 U9 ( .A(n32), .B(n3), .Y(n1) );
  BUFX16 U10 ( .A(n22), .Y(n2) );
  NAND3BX4 U11 ( .AN(B[9]), .B(A[9]), .C(n13), .Y(n138) );
  BUFX8 U12 ( .A(n78), .Y(n7) );
  AOI21X4 U13 ( .A0(n34), .A1(n123), .B0(n124), .Y(n122) );
  BUFX16 U14 ( .A(n67), .Y(n10) );
  INVX2 U15 ( .A(n71), .Y(n74) );
  NAND2X4 U16 ( .A(n161), .B(n3), .Y(n160) );
  CLKINVX8 U17 ( .A(n3), .Y(n141) );
  BUFX8 U18 ( .A(n26), .Y(n3) );
  XOR2X4 U19 ( .A(n121), .B(n122), .Y(DIFF[14]) );
  AOI21X2 U20 ( .A0(n90), .A1(n91), .B0(n127), .Y(n126) );
  INVX1 U21 ( .A(A[6]), .Y(n166) );
  CLKINVX3 U22 ( .A(n56), .Y(n108) );
  NOR2X1 U23 ( .A(n27), .B(n28), .Y(n24) );
  INVX1 U24 ( .A(n2), .Y(n5) );
  NAND2BX1 U25 ( .AN(B[8]), .B(A[8]), .Y(n26) );
  OR2X2 U26 ( .A(n98), .B(n120), .Y(n18) );
  OAI21X2 U27 ( .A0(n117), .A1(n98), .B0(n93), .Y(n116) );
  INVX1 U28 ( .A(n119), .Y(n129) );
  OAI21X2 U29 ( .A0(n69), .A1(n70), .B0(n71), .Y(n65) );
  INVX1 U30 ( .A(n54), .Y(n59) );
  NAND2X2 U31 ( .A(n12), .B(n2), .Y(n8) );
  NAND2BX2 U32 ( .AN(B[7]), .B(A[7]), .Y(n40) );
  AND2X2 U33 ( .A(n142), .B(n119), .Y(n17) );
  NAND2X1 U34 ( .A(n13), .B(n31), .Y(n146) );
  NAND2X1 U35 ( .A(n88), .B(n93), .Y(n121) );
  NOR2X1 U36 ( .A(n130), .B(n105), .Y(n123) );
  INVX1 U37 ( .A(n81), .Y(n97) );
  NAND3BX2 U38 ( .AN(n98), .B(n99), .C(n89), .Y(n81) );
  INVX4 U39 ( .A(n117), .Y(n90) );
  NAND2BX1 U40 ( .AN(n129), .B(n114), .Y(n102) );
  INVX2 U41 ( .A(n37), .Y(n42) );
  OR2X2 U42 ( .A(n156), .B(n157), .Y(n15) );
  INVX1 U43 ( .A(n143), .Y(n157) );
  NOR2X1 U44 ( .A(n127), .B(n128), .Y(n132) );
  NAND2XL U45 ( .A(n91), .B(n99), .Y(n130) );
  AOI21XL U46 ( .A0(n90), .A1(n91), .B0(n92), .Y(n85) );
  OR2X2 U47 ( .A(n30), .B(n28), .Y(n4) );
  NAND3X4 U48 ( .A(n31), .B(n13), .C(n141), .Y(n139) );
  NAND2X1 U49 ( .A(n55), .B(n56), .Y(n49) );
  NAND4BBX2 U50 ( .AN(n152), .BN(B[4]), .C(n153), .D(n154), .Y(n150) );
  NAND2BX2 U51 ( .AN(A[5]), .B(B[5]), .Y(n153) );
  NOR2X2 U52 ( .A(n90), .B(n120), .Y(n136) );
  CLKINVX4 U53 ( .A(n105), .Y(n96) );
  NAND2XL U54 ( .A(n88), .B(n89), .Y(n86) );
  NAND2X4 U55 ( .A(n10), .B(n77), .Y(n172) );
  NAND4BX4 U56 ( .AN(n76), .B(n75), .C(n64), .D(n10), .Y(n53) );
  NAND2BXL U57 ( .AN(B[15]), .B(A[15]), .Y(n87) );
  NOR2X4 U58 ( .A(n4), .B(n5), .Y(n6) );
  NOR2X4 U59 ( .A(n6), .B(n23), .Y(n21) );
  OAI2BB1X2 U60 ( .A0N(n24), .A1N(n25), .B0(n3), .Y(n23) );
  NAND2BX2 U61 ( .AN(B[14]), .B(A[14]), .Y(n93) );
  NAND2BX1 U62 ( .AN(A[6]), .B(B[6]), .Y(n37) );
  NAND2BX2 U63 ( .AN(A[6]), .B(B[6]), .Y(n154) );
  NAND2BX2 U64 ( .AN(B[4]), .B(A[4]), .Y(n54) );
  NAND2BX2 U65 ( .AN(B[2]), .B(A[2]), .Y(n171) );
  OAI21X2 U66 ( .A0(n80), .A1(n81), .B0(n82), .Y(n78) );
  INVX1 U67 ( .A(B[6]), .Y(n168) );
  INVX8 U68 ( .A(n30), .Y(n95) );
  NAND2BX4 U69 ( .AN(A[3]), .B(B[3]), .Y(n67) );
  NOR2X1 U70 ( .A(n74), .B(n70), .Y(n73) );
  CLKINVX4 U71 ( .A(n75), .Y(n70) );
  NOR2X4 U72 ( .A(n147), .B(n148), .Y(n145) );
  XNOR2X4 U73 ( .A(n34), .B(n14), .Y(DIFF[8]) );
  OAI21X4 U74 ( .A0(n145), .A1(n146), .B0(n143), .Y(n144) );
  NAND2BX2 U75 ( .AN(A[5]), .B(B[5]), .Y(n48) );
  NOR2BX2 U76 ( .AN(A[5]), .B(B[5]), .Y(n167) );
  NAND2BXL U77 ( .AN(B[5]), .B(A[5]), .Y(n46) );
  NAND2BX2 U78 ( .AN(A[7]), .B(B[7]), .Y(n29) );
  NAND2X4 U79 ( .A(n66), .B(n10), .Y(n56) );
  NAND2BX4 U80 ( .AN(A[8]), .B(B[8]), .Y(n33) );
  NAND4BX4 U81 ( .AN(n51), .B(n52), .C(n11), .D(n54), .Y(n50) );
  NOR2X4 U82 ( .A(n49), .B(n50), .Y(n44) );
  NAND3X1 U83 ( .A(n99), .B(n119), .C(n114), .Y(n133) );
  XOR2X4 U84 ( .A(n109), .B(n110), .Y(DIFF[15]) );
  AOI21X4 U85 ( .A0(n34), .A1(n111), .B0(n112), .Y(n110) );
  AOI21X2 U86 ( .A0(n64), .A1(n65), .B0(n66), .Y(n63) );
  NAND3X4 U87 ( .A(n64), .B(n74), .C(n10), .Y(n55) );
  OAI21X4 U88 ( .A0(n164), .A1(n165), .B0(n151), .Y(n163) );
  NAND2BX2 U89 ( .AN(B[10]), .B(A[10]), .Y(n143) );
  NAND2BX2 U90 ( .AN(A[10]), .B(B[10]), .Y(n140) );
  NAND2XL U91 ( .A(n33), .B(n3), .Y(n14) );
  OAI21X4 U92 ( .A0(n162), .A1(n163), .B0(n29), .Y(n161) );
  NAND2BX2 U93 ( .AN(B[1]), .B(A[1]), .Y(n71) );
  NOR2X4 U94 ( .A(n39), .B(n42), .Y(n41) );
  NAND2X2 U95 ( .A(n25), .B(n29), .Y(n104) );
  NOR3BX2 U96 ( .AN(n2), .B(n30), .C(n28), .Y(n148) );
  XOR2X2 U97 ( .A(n62), .B(n63), .Y(DIFF[3]) );
  NAND2BX4 U98 ( .AN(B[6]), .B(A[6]), .Y(n43) );
  OAI21X2 U99 ( .A0(n168), .A1(A[6]), .B0(A[4]), .Y(n165) );
  NAND2BX2 U100 ( .AN(B[11]), .B(A[11]), .Y(n142) );
  AOI21X4 U101 ( .A0(n37), .A1(n38), .B0(n39), .Y(n36) );
  XOR2X4 U102 ( .A(n38), .B(n41), .Y(DIFF[6]) );
  OAI2BB1X2 U103 ( .A0N(n34), .A1N(n96), .B0(n102), .Y(n135) );
  INVX4 U104 ( .A(n29), .Y(n27) );
  NAND2XL U105 ( .A(n31), .B(n32), .Y(n20) );
  NAND2BX2 U106 ( .AN(B[9]), .B(A[9]), .Y(n32) );
  OAI2BB1X4 U107 ( .A0N(n125), .A1N(n114), .B0(n126), .Y(n124) );
  NOR3X2 U108 ( .A(n120), .B(n128), .C(n129), .Y(n125) );
  AOI2BB1X2 U109 ( .A0N(n98), .A1N(n94), .B0(n116), .Y(n115) );
  NOR2X1 U110 ( .A(n118), .B(n98), .Y(n113) );
  NOR2X2 U111 ( .A(n18), .B(n105), .Y(n111) );
  XOR2X4 U112 ( .A(n20), .B(n21), .Y(DIFF[9]) );
  NAND2BX4 U113 ( .AN(A[14]), .B(B[14]), .Y(n88) );
  BUFX8 U114 ( .A(n53), .Y(n11) );
  INVX4 U115 ( .A(n94), .Y(n127) );
  NAND2X2 U116 ( .A(n93), .B(n94), .Y(n92) );
  NAND2BX2 U117 ( .AN(B[13]), .B(A[13]), .Y(n94) );
  NAND2BX2 U118 ( .AN(B[12]), .B(A[12]), .Y(n117) );
  NAND2BX2 U119 ( .AN(B[3]), .B(A[3]), .Y(n52) );
  XNOR2X2 U120 ( .A(n65), .B(n16), .Y(DIFF[2]) );
  NOR2X2 U121 ( .A(n83), .B(n84), .Y(n82) );
  XOR2X2 U122 ( .A(n72), .B(n73), .Y(DIFF[1]) );
  NAND2BX2 U123 ( .AN(A[4]), .B(B[4]), .Y(n47) );
  NAND2X1 U124 ( .A(n10), .B(n52), .Y(n62) );
  INVX2 U125 ( .A(n43), .Y(n39) );
  NAND2X1 U126 ( .A(n40), .B(n43), .Y(n162) );
  NAND2X2 U127 ( .A(n64), .B(n75), .Y(n173) );
  NAND2BX4 U128 ( .AN(A[1]), .B(B[1]), .Y(n75) );
  XOR2X2 U129 ( .A(n2), .B(n60), .Y(DIFF[4]) );
  AND4X2 U130 ( .A(n51), .B(n95), .C(n96), .D(n97), .Y(n83) );
  NOR2X4 U131 ( .A(n172), .B(n173), .Y(n51) );
  INVX4 U132 ( .A(n91), .Y(n128) );
  NAND2BX4 U133 ( .AN(A[13]), .B(B[13]), .Y(n91) );
  NAND3X2 U134 ( .A(n99), .B(n96), .C(n34), .Y(n134) );
  XNOR2X4 U135 ( .A(n155), .B(n15), .Y(DIFF[10]) );
  OAI21X4 U136 ( .A0(n158), .A1(n159), .B0(n32), .Y(n155) );
  OAI2BB1X4 U137 ( .A0N(n166), .A1N(B[6]), .B0(n167), .Y(n151) );
  NAND3X4 U138 ( .A(n19), .B(n150), .C(n151), .Y(n25) );
  OAI2BB1X2 U139 ( .A0N(n113), .A1N(n114), .B0(n115), .Y(n112) );
  INVX4 U140 ( .A(n171), .Y(n66) );
  NAND4BX4 U141 ( .AN(n174), .B(n175), .C(n12), .D(n48), .Y(n30) );
  AOI21X2 U142 ( .A0(n95), .A1(n2), .B0(n160), .Y(n158) );
  NAND2BX4 U143 ( .AN(A[2]), .B(B[2]), .Y(n64) );
  AND2X4 U144 ( .A(n8), .B(n9), .Y(n58) );
  XOR2X4 U145 ( .A(n57), .B(n58), .Y(DIFF[5]) );
  NAND3X2 U146 ( .A(n133), .B(n117), .C(n134), .Y(n131) );
  NAND2XL U147 ( .A(n29), .B(n40), .Y(n35) );
  AND2X2 U148 ( .A(n40), .B(n43), .Y(n19) );
  INVX8 U149 ( .A(n33), .Y(n28) );
  NAND2X1 U150 ( .A(n99), .B(n119), .Y(n118) );
  NAND2BX4 U151 ( .AN(A[11]), .B(B[11]), .Y(n119) );
  NAND2BX4 U152 ( .AN(A[9]), .B(B[9]), .Y(n31) );
  BUFX8 U153 ( .A(n140), .Y(n13) );
  NAND2X4 U154 ( .A(n91), .B(n88), .Y(n98) );
  NAND2XL U155 ( .A(n87), .B(n89), .Y(n109) );
  XOR2X4 U156 ( .A(n144), .B(n17), .Y(DIFF[11]) );
  OAI21X1 U157 ( .A0(n85), .A1(n86), .B0(n87), .Y(n84) );
  INVX1 U158 ( .A(n102), .Y(n101) );
  NAND2X1 U159 ( .A(n31), .B(n33), .Y(n159) );
  NAND2X2 U160 ( .A(n142), .B(n143), .Y(n137) );
  NOR2BX1 U161 ( .AN(B[7]), .B(A[7]), .Y(n174) );
  NAND2X2 U162 ( .A(n153), .B(n169), .Y(n164) );
  INVX1 U163 ( .A(n13), .Y(n156) );
  NOR2X2 U164 ( .A(n59), .B(n61), .Y(n60) );
  INVXL U165 ( .A(n12), .Y(n61) );
  NOR2X1 U166 ( .A(n100), .B(n101), .Y(n80) );
  AOI21XL U167 ( .A0(n103), .A1(n104), .B0(n105), .Y(n100) );
  INVX1 U168 ( .A(n64), .Y(n68) );
  NAND2XL U169 ( .A(n48), .B(n46), .Y(n57) );
  INVXL U170 ( .A(B[4]), .Y(n169) );
  INVX1 U171 ( .A(n72), .Y(n69) );
  OAI21XL U172 ( .A0(n106), .A1(n107), .B0(n95), .Y(n103) );
  NAND2XL U173 ( .A(n11), .B(n52), .Y(n106) );
  NAND2BXL U174 ( .AN(n108), .B(n55), .Y(n107) );
  XNOR2X1 U175 ( .A(B[16]), .B(A[16]), .Y(n79) );
  NAND2X1 U176 ( .A(n76), .B(n77), .Y(DIFF[0]) );
  NAND2BX1 U177 ( .AN(n77), .B(n76), .Y(n72) );
  NAND2BX1 U178 ( .AN(A[0]), .B(B[0]), .Y(n77) );
  NAND2BX1 U179 ( .AN(B[0]), .B(A[0]), .Y(n76) );
  INVXL U180 ( .A(A[4]), .Y(n152) );
  NAND3X1 U181 ( .A(n33), .B(n29), .C(n25), .Y(n149) );
  NAND2BX1 U182 ( .AN(A[6]), .B(B[6]), .Y(n175) );
  NAND2X2 U183 ( .A(n12), .B(n48), .Y(n45) );
  XOR2X4 U184 ( .A(n35), .B(n36), .Y(DIFF[7]) );
  OAI21X4 U185 ( .A0(n44), .A1(n45), .B0(n46), .Y(n38) );
  XOR2X4 U186 ( .A(n7), .B(n79), .Y(DIFF[16]) );
  NAND2BX4 U187 ( .AN(A[15]), .B(B[15]), .Y(n89) );
  XOR2X4 U188 ( .A(n131), .B(n132), .Y(DIFF[13]) );
  XOR2X4 U189 ( .A(n135), .B(n136), .Y(DIFF[12]) );
  NAND2BX4 U190 ( .AN(A[12]), .B(B[12]), .Y(n99) );
  NAND3BX4 U191 ( .AN(n137), .B(n138), .C(n139), .Y(n114) );
  NAND4BX4 U192 ( .AN(n28), .B(n31), .C(n119), .D(n13), .Y(n105) );
  OAI2BB1X4 U193 ( .A0N(n95), .A1N(n2), .B0(n104), .Y(n34) );
  NAND4BX4 U194 ( .AN(n51), .B(n170), .C(n11), .D(n52), .Y(n22) );
endmodule


module butterfly_DW01_add_140 ( A, B, SUM );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  wire   n180, n181, n182, n183, n184, n185, n186, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179;

  BUFX3 U2 ( .A(n56), .Y(n5) );
  NAND2X1 U3 ( .A(B[6]), .B(A[6]), .Y(n56) );
  NAND3BX2 U4 ( .AN(n94), .B(n3), .C(n92), .Y(n140) );
  NOR2X1 U5 ( .A(n94), .B(n119), .Y(n132) );
  NAND2X4 U6 ( .A(n11), .B(n48), .Y(n94) );
  NOR2X1 U7 ( .A(A[5]), .B(B[5]), .Y(n178) );
  INVX4 U8 ( .A(n41), .Y(n1) );
  CLKINVX3 U9 ( .A(n1), .Y(n2) );
  CLKINVX8 U10 ( .A(n1), .Y(n3) );
  INVX8 U11 ( .A(n60), .Y(n65) );
  INVX4 U12 ( .A(n119), .Y(n127) );
  BUFX20 U13 ( .A(n183), .Y(SUM[8]) );
  NAND3X2 U14 ( .A(n74), .B(n73), .C(n72), .Y(n112) );
  NOR2X4 U15 ( .A(A[5]), .B(B[5]), .Y(n4) );
  INVX20 U16 ( .A(n4), .Y(n59) );
  INVX8 U17 ( .A(n14), .Y(SUM[1]) );
  NAND2X2 U18 ( .A(B[2]), .B(A[2]), .Y(n80) );
  NAND4X1 U19 ( .A(n46), .B(n48), .C(n49), .D(n47), .Y(n160) );
  NAND2X4 U20 ( .A(n142), .B(n45), .Y(n125) );
  OR2X4 U21 ( .A(A[6]), .B(B[6]), .Y(n48) );
  NAND3X2 U22 ( .A(n133), .B(n131), .C(n130), .Y(n137) );
  INVX3 U23 ( .A(n72), .Y(n78) );
  NAND3X1 U24 ( .A(A[9]), .B(B[9]), .C(n145), .Y(n143) );
  CLKINVX4 U25 ( .A(n71), .Y(n69) );
  NAND2X4 U26 ( .A(B[3]), .B(A[3]), .Y(n71) );
  OAI2BB1X4 U27 ( .A0N(B[5]), .A1N(A[5]), .B0(n171), .Y(n47) );
  NAND2XL U28 ( .A(B[13]), .B(A[13]), .Y(n102) );
  OR2X4 U29 ( .A(A[13]), .B(B[13]), .Y(n126) );
  NAND3BX4 U30 ( .AN(n179), .B(B[6]), .C(A[6]), .Y(n45) );
  OR2X4 U31 ( .A(A[6]), .B(B[6]), .Y(n39) );
  NOR2BX4 U32 ( .AN(n5), .B(n62), .Y(n64) );
  NOR2X4 U33 ( .A(n61), .B(n62), .Y(n55) );
  INVX8 U34 ( .A(n58), .Y(n62) );
  BUFX8 U35 ( .A(n39), .Y(n6) );
  AND2X1 U36 ( .A(B[6]), .B(A[6]), .Y(n162) );
  OR2X4 U37 ( .A(A[6]), .B(B[6]), .Y(n58) );
  OAI21X4 U38 ( .A0(n100), .A1(n101), .B0(n102), .Y(n98) );
  INVX1 U39 ( .A(n120), .Y(n19) );
  INVX4 U40 ( .A(n54), .Y(n151) );
  NAND2BX1 U41 ( .AN(n129), .B(n130), .Y(n122) );
  NAND2X1 U42 ( .A(n127), .B(n131), .Y(n129) );
  NOR2BX1 U43 ( .AN(n118), .B(n107), .Y(n120) );
  NAND2BX1 U44 ( .AN(n163), .B(n42), .Y(n37) );
  INVX1 U45 ( .A(n131), .Y(n154) );
  NAND2X1 U46 ( .A(B[11]), .B(A[11]), .Y(n146) );
  NAND4BBX2 U47 ( .AN(n15), .BN(n52), .C(n36), .D(n45), .Y(n169) );
  NAND2X1 U48 ( .A(B[9]), .B(A[9]), .Y(n34) );
  INVX1 U49 ( .A(n133), .Y(n108) );
  INVX1 U50 ( .A(n15), .Y(n111) );
  NAND2X1 U51 ( .A(B[12]), .B(A[12]), .Y(n101) );
  INVX1 U52 ( .A(n126), .Y(n100) );
  OR2X2 U53 ( .A(A[14]), .B(B[14]), .Y(n97) );
  NOR2X1 U54 ( .A(A[15]), .B(B[15]), .Y(n25) );
  AOI22X2 U55 ( .A0(B[2]), .A1(A[2]), .B0(B[1]), .B1(A[1]), .Y(n174) );
  INVX4 U56 ( .A(n49), .Y(n163) );
  AND2X2 U57 ( .A(n102), .B(n126), .Y(n7) );
  AND2X2 U58 ( .A(n44), .B(n54), .Y(n8) );
  AND2X2 U59 ( .A(n36), .B(n49), .Y(n9) );
  AND2X2 U60 ( .A(n34), .B(n35), .Y(n10) );
  AND2X4 U61 ( .A(n150), .B(n70), .Y(n11) );
  NAND3BX1 U62 ( .AN(n128), .B(n3), .C(n132), .Y(n121) );
  NOR2X1 U63 ( .A(A[7]), .B(B[7]), .Y(n179) );
  XOR2X4 U64 ( .A(n12), .B(n9), .Y(n183) );
  NAND3X4 U65 ( .A(n50), .B(n51), .C(n45), .Y(n12) );
  AND3X4 U66 ( .A(n6), .B(n40), .C(n2), .Y(n13) );
  NAND2X2 U67 ( .A(n92), .B(n125), .Y(n141) );
  CLKINVX8 U68 ( .A(n128), .Y(n92) );
  XOR2X4 U69 ( .A(n87), .B(n86), .Y(n14) );
  NAND3X1 U70 ( .A(n49), .B(n54), .C(n162), .Y(n161) );
  NOR2X2 U71 ( .A(n164), .B(n165), .Y(n157) );
  NOR2BX2 U72 ( .AN(n61), .B(n4), .Y(n66) );
  NAND3X1 U73 ( .A(n46), .B(n47), .C(n48), .Y(n43) );
  OAI2BB1X4 U74 ( .A0N(n81), .A1N(n73), .B0(n80), .Y(n76) );
  NAND2X2 U75 ( .A(B[5]), .B(A[5]), .Y(n61) );
  NAND4BX4 U76 ( .AN(n135), .B(n138), .C(n136), .D(n137), .Y(n134) );
  INVX8 U77 ( .A(n164), .Y(n40) );
  AND3X4 U78 ( .A(n39), .B(n46), .C(n47), .Y(n15) );
  NAND3X2 U79 ( .A(n58), .B(n11), .C(n2), .Y(n51) );
  AND2X1 U80 ( .A(n171), .B(n70), .Y(n75) );
  OR2X4 U81 ( .A(A[4]), .B(B[4]), .Y(n16) );
  NAND2X4 U82 ( .A(n35), .B(n49), .Y(n148) );
  NAND3BX4 U83 ( .AN(n159), .B(n160), .C(n161), .Y(n158) );
  OAI211X2 U84 ( .A0(n163), .A1(n44), .B0(n36), .C0(n34), .Y(n159) );
  NAND3BX2 U85 ( .AN(n128), .B(n133), .C(n125), .Y(n136) );
  NAND2X2 U86 ( .A(B[4]), .B(A[4]), .Y(n171) );
  NAND2X4 U87 ( .A(n69), .B(n70), .Y(n68) );
  AOI21XL U88 ( .A0(n112), .A1(n71), .B0(n94), .Y(n109) );
  OAI2BB1X2 U89 ( .A0N(n115), .A1N(n116), .B0(n117), .Y(n113) );
  NAND3X2 U90 ( .A(n6), .B(n40), .C(n3), .Y(n38) );
  OAI21X4 U91 ( .A0(A[11]), .A1(B[11]), .B0(n145), .Y(n149) );
  NAND3X2 U92 ( .A(n60), .B(n58), .C(n59), .Y(n57) );
  NAND3X2 U93 ( .A(n43), .B(n44), .C(n45), .Y(n42) );
  XNOR2X4 U94 ( .A(n81), .B(n82), .Y(n21) );
  NAND2X4 U95 ( .A(B[8]), .B(A[8]), .Y(n36) );
  NAND4X2 U96 ( .A(n74), .B(n16), .C(n73), .D(n72), .Y(n67) );
  NAND2X2 U97 ( .A(B[10]), .B(A[10]), .Y(n147) );
  OAI21X4 U98 ( .A0(n155), .A1(n156), .B0(n147), .Y(n152) );
  INVX3 U99 ( .A(n73), .Y(n79) );
  INVX8 U100 ( .A(n18), .Y(SUM[14]) );
  NAND4BBX2 U101 ( .AN(n128), .BN(n94), .C(n3), .D(n133), .Y(n138) );
  XNOR2X4 U102 ( .A(n65), .B(n66), .Y(SUM[5]) );
  AOI21X2 U103 ( .A0(n124), .A1(n125), .B0(n98), .Y(n123) );
  NOR2BX2 U104 ( .AN(n127), .B(n128), .Y(n124) );
  AOI21X2 U105 ( .A0(n157), .A1(n3), .B0(n158), .Y(n155) );
  OAI21X1 U106 ( .A0(A[8]), .A1(B[8]), .B0(n70), .Y(n176) );
  NAND3X4 U107 ( .A(n140), .B(n103), .C(n141), .Y(n116) );
  BUFX20 U108 ( .A(n180), .Y(SUM[13]) );
  NAND3BX4 U109 ( .AN(n55), .B(n5), .C(n57), .Y(n53) );
  BUFX20 U110 ( .A(n186), .Y(SUM[4]) );
  AOI31X2 U111 ( .A0(n6), .A1(n46), .A2(n47), .B0(n52), .Y(n142) );
  OAI22X2 U112 ( .A0(A[5]), .A1(B[5]), .B0(A[7]), .B1(B[7]), .Y(n172) );
  NOR2X4 U113 ( .A(B[1]), .B(A[1]), .Y(n173) );
  OR2X4 U114 ( .A(A[4]), .B(B[4]), .Y(n70) );
  INVX4 U115 ( .A(n172), .Y(n46) );
  BUFX20 U116 ( .A(n181), .Y(SUM[11]) );
  BUFX20 U117 ( .A(n185), .Y(SUM[6]) );
  BUFX20 U118 ( .A(n184), .Y(SUM[7]) );
  BUFX20 U119 ( .A(n182), .Y(SUM[9]) );
  NAND2XL U120 ( .A(B[15]), .B(A[15]), .Y(n96) );
  INVX8 U121 ( .A(n21), .Y(SUM[2]) );
  XOR2X4 U122 ( .A(n134), .B(n7), .Y(n180) );
  AOI21XL U123 ( .A0(n98), .A1(n97), .B0(n99), .Y(n117) );
  INVXL U124 ( .A(n101), .Y(n135) );
  NOR2X2 U125 ( .A(n52), .B(n15), .Y(n50) );
  OAI21X4 U126 ( .A0(n65), .A1(n4), .B0(n61), .Y(n63) );
  INVX4 U127 ( .A(n44), .Y(n52) );
  NOR2BX1 U128 ( .AN(n35), .B(n163), .Y(n170) );
  NOR2XL U129 ( .A(n100), .B(n108), .Y(n105) );
  NAND2X2 U130 ( .A(n130), .B(n131), .Y(n103) );
  AND2X4 U131 ( .A(n146), .B(n147), .Y(n22) );
  OR2X4 U132 ( .A(B[1]), .B(A[1]), .Y(n83) );
  NAND2XL U133 ( .A(B[14]), .B(A[14]), .Y(n118) );
  INVX1 U134 ( .A(n6), .Y(n165) );
  XOR2X4 U135 ( .A(n166), .B(n167), .Y(n17) );
  INVX8 U136 ( .A(n17), .Y(SUM[10]) );
  NAND3BXL U137 ( .AN(n52), .B(n45), .C(n111), .Y(n110) );
  XNOR2X4 U138 ( .A(n20), .B(n19), .Y(n18) );
  AND3X4 U139 ( .A(n121), .B(n122), .C(n123), .Y(n20) );
  NAND2X2 U140 ( .A(B[7]), .B(A[7]), .Y(n44) );
  NOR2BX1 U141 ( .AN(n146), .B(n154), .Y(n153) );
  NAND3X4 U142 ( .A(n22), .B(n143), .C(n144), .Y(n130) );
  XOR2X4 U143 ( .A(n116), .B(n24), .Y(n23) );
  INVX8 U144 ( .A(n23), .Y(SUM[12]) );
  CLKINVX20 U145 ( .A(n139), .Y(n24) );
  NOR2BX1 U146 ( .AN(n96), .B(n25), .Y(n114) );
  NOR2XL U147 ( .A(n119), .B(n107), .Y(n115) );
  INVX1 U148 ( .A(n97), .Y(n107) );
  INVX1 U149 ( .A(n118), .Y(n99) );
  OAI21XL U150 ( .A0(n95), .A1(n25), .B0(n96), .Y(n91) );
  AOI21X1 U151 ( .A0(n97), .A1(n98), .B0(n99), .Y(n95) );
  NAND2XL U152 ( .A(n147), .B(n145), .Y(n167) );
  AOI21XL U153 ( .A0(n103), .A1(n104), .B0(n93), .Y(n90) );
  NAND2X1 U154 ( .A(n105), .B(n106), .Y(n93) );
  OAI21XL U155 ( .A0(n109), .A1(n110), .B0(n92), .Y(n104) );
  NOR2XL U156 ( .A(n25), .B(n107), .Y(n106) );
  NAND2XL U157 ( .A(n145), .B(n35), .Y(n156) );
  XOR2X2 U158 ( .A(n88), .B(n89), .Y(SUM[16]) );
  XNOR2X1 U159 ( .A(B[16]), .B(A[16]), .Y(n88) );
  NOR2X1 U160 ( .A(n90), .B(n91), .Y(n89) );
  OR2X2 U161 ( .A(A[11]), .B(B[11]), .Y(n131) );
  INVX1 U162 ( .A(n87), .Y(n84) );
  AND2X2 U163 ( .A(n87), .B(n175), .Y(SUM[0]) );
  OR2X2 U164 ( .A(A[0]), .B(B[0]), .Y(n175) );
  NAND2X1 U165 ( .A(B[0]), .B(A[0]), .Y(n87) );
  NAND2X4 U166 ( .A(n71), .B(n112), .Y(n41) );
  NOR2BX4 U167 ( .AN(n71), .B(n78), .Y(n77) );
  NAND2X2 U168 ( .A(A[1]), .B(B[1]), .Y(n85) );
  NAND3BX2 U169 ( .AN(n36), .B(n145), .C(n35), .Y(n144) );
  XOR2X4 U170 ( .A(n33), .B(n10), .Y(n182) );
  NAND3X4 U171 ( .A(n36), .B(n37), .C(n38), .Y(n33) );
  XOR2X4 U172 ( .A(n53), .B(n8), .Y(n184) );
  XOR2X4 U173 ( .A(n63), .B(n64), .Y(n185) );
  NAND3X4 U174 ( .A(n67), .B(n171), .C(n68), .Y(n60) );
  XOR2X4 U175 ( .A(n3), .B(n75), .Y(n186) );
  XOR2X4 U176 ( .A(n76), .B(n77), .Y(SUM[3]) );
  NOR2BX4 U177 ( .AN(n80), .B(n79), .Y(n82) );
  OAI2BB1X4 U178 ( .A0N(n83), .A1N(n84), .B0(n85), .Y(n81) );
  NOR2BX4 U179 ( .AN(n85), .B(n173), .Y(n86) );
  XOR2X4 U180 ( .A(n113), .B(n114), .Y(SUM[15]) );
  NAND2X4 U181 ( .A(n133), .B(n126), .Y(n119) );
  NOR2BX4 U182 ( .AN(n101), .B(n108), .Y(n139) );
  OR2X4 U183 ( .A(A[12]), .B(B[12]), .Y(n133) );
  OR2X4 U184 ( .A(n148), .B(n149), .Y(n128) );
  NOR2X4 U185 ( .A(n151), .B(n4), .Y(n150) );
  XOR2X4 U186 ( .A(n152), .B(n153), .Y(n181) );
  OR2X4 U187 ( .A(A[10]), .B(B[10]), .Y(n145) );
  NAND2X4 U188 ( .A(n34), .B(n168), .Y(n166) );
  OAI21X4 U189 ( .A0(n13), .A1(n169), .B0(n170), .Y(n168) );
  OR2X4 U190 ( .A(A[8]), .B(B[8]), .Y(n49) );
  OR2X4 U191 ( .A(A[9]), .B(B[9]), .Y(n35) );
  OR2X4 U192 ( .A(A[7]), .B(B[7]), .Y(n54) );
  OAI21X4 U193 ( .A0(n173), .A1(n87), .B0(n174), .Y(n74) );
  OR2X4 U194 ( .A(A[2]), .B(B[2]), .Y(n73) );
  OR2X4 U195 ( .A(A[3]), .B(B[3]), .Y(n72) );
  NAND2BX4 U196 ( .AN(n176), .B(n177), .Y(n164) );
  NOR2X4 U197 ( .A(n178), .B(n151), .Y(n177) );
endmodule


module butterfly_DW01_sub_112 ( A, B, DIFF );
  input [16:0] A;
  input [16:0] B;
  output [16:0] DIFF;
  wire   n253, n254, n255, n256, n257, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n24, n26,
         n27, n28, n29, n31, n32, n33, n34, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252;

  INVX4 U3 ( .A(n16), .Y(n210) );
  CLKINVX2 U4 ( .A(n74), .Y(n18) );
  NAND2X4 U5 ( .A(n73), .B(n74), .Y(n198) );
  OR2X2 U6 ( .A(n191), .B(n197), .Y(n32) );
  OAI21X4 U7 ( .A0(n235), .A1(n234), .B0(n236), .Y(n233) );
  NAND3BX4 U8 ( .AN(n78), .B(n68), .C(n49), .Y(n204) );
  OR2X4 U9 ( .A(n31), .B(n194), .Y(n205) );
  NOR2X2 U10 ( .A(n20), .B(n76), .Y(n72) );
  INVX1 U11 ( .A(n38), .Y(n27) );
  NAND2X2 U12 ( .A(n5), .B(n57), .Y(n93) );
  NOR2X2 U13 ( .A(n114), .B(n124), .Y(n8) );
  INVX4 U14 ( .A(n2), .Y(n114) );
  INVX8 U15 ( .A(n15), .Y(n124) );
  NOR2X4 U16 ( .A(n86), .B(n87), .Y(n81) );
  NAND3X2 U17 ( .A(n88), .B(n22), .C(n62), .Y(n86) );
  AND2X4 U18 ( .A(n57), .B(n88), .Y(n38) );
  NOR4X4 U19 ( .A(n176), .B(n177), .C(n178), .D(n179), .Y(n175) );
  BUFX12 U20 ( .A(n257), .Y(DIFF[1]) );
  BUFX8 U21 ( .A(n60), .Y(n24) );
  AOI21X2 U22 ( .A0(n189), .A1(n151), .B0(n190), .Y(n188) );
  CLKINVX3 U23 ( .A(n31), .Y(n161) );
  INVX1 U24 ( .A(n108), .Y(n9) );
  INVX1 U25 ( .A(n174), .Y(n171) );
  NOR2X1 U26 ( .A(n174), .B(n182), .Y(n176) );
  NOR2X1 U27 ( .A(n174), .B(n153), .Y(n178) );
  NOR2X2 U28 ( .A(n119), .B(n120), .Y(n115) );
  NOR2BX1 U29 ( .AN(n58), .B(n31), .Y(n225) );
  INVX1 U30 ( .A(n69), .Y(n66) );
  INVX1 U31 ( .A(n242), .Y(n111) );
  AOI21X1 U32 ( .A0(n195), .A1(n196), .B0(n197), .Y(n186) );
  INVX1 U33 ( .A(n143), .Y(n197) );
  INVX1 U34 ( .A(n168), .Y(n136) );
  OAI21XL U35 ( .A0(n142), .A1(n143), .B0(n144), .Y(n139) );
  NAND3X2 U36 ( .A(n50), .B(n215), .C(n69), .Y(n212) );
  AND2X2 U37 ( .A(n39), .B(n84), .Y(n83) );
  NAND2BX1 U38 ( .AN(n31), .B(n57), .Y(n82) );
  INVX8 U39 ( .A(n6), .Y(DIFF[6]) );
  XOR2X2 U40 ( .A(n89), .B(n90), .Y(n6) );
  NAND2X1 U41 ( .A(n84), .B(n91), .Y(n90) );
  XOR2X2 U42 ( .A(n128), .B(n129), .Y(DIFF[16]) );
  CLKINVX4 U43 ( .A(n71), .Y(n26) );
  BUFX16 U44 ( .A(n98), .Y(n2) );
  CLKINVX3 U45 ( .A(A[4]), .Y(n244) );
  AND2X2 U46 ( .A(n56), .B(n80), .Y(n3) );
  BUFX8 U47 ( .A(n63), .Y(n22) );
  CLKINVX3 U48 ( .A(n22), .Y(n101) );
  AND2X2 U49 ( .A(n49), .B(n50), .Y(n4) );
  AND2X2 U50 ( .A(n2), .B(n96), .Y(n5) );
  INVX8 U51 ( .A(n40), .Y(DIFF[11]) );
  NAND3BX2 U52 ( .AN(B[2]), .B(n11), .C(n2), .Y(n60) );
  NAND2BXL U53 ( .AN(A[8]), .B(B[8]), .Y(n200) );
  NOR2X4 U54 ( .A(n97), .B(n111), .Y(n110) );
  INVX2 U55 ( .A(n216), .Y(n7) );
  CLKINVX3 U56 ( .A(A[9]), .Y(n216) );
  NOR2X2 U57 ( .A(n191), .B(n158), .Y(n195) );
  NAND2BXL U58 ( .AN(n16), .B(n150), .Y(n132) );
  NAND2X4 U59 ( .A(n239), .B(n50), .Y(n238) );
  OAI22X4 U60 ( .A0(n229), .A1(n227), .B0(n227), .B1(n54), .Y(n219) );
  CLKINVX4 U61 ( .A(n55), .Y(n229) );
  OAI22X4 U62 ( .A0(n54), .A1(n240), .B0(n240), .B1(n69), .Y(n237) );
  NAND2XL U63 ( .A(n214), .B(n153), .Y(n218) );
  INVX2 U64 ( .A(n153), .Y(n189) );
  OR2X2 U65 ( .A(n31), .B(n85), .Y(n39) );
  NAND3X2 U66 ( .A(n151), .B(n49), .C(n68), .Y(n193) );
  NAND4BBX2 U67 ( .AN(n31), .BN(n240), .C(n57), .D(n56), .Y(n234) );
  NAND2BX2 U68 ( .AN(B[7]), .B(A[7]), .Y(n80) );
  NAND2X2 U69 ( .A(n62), .B(n22), .Y(n36) );
  INVX3 U70 ( .A(n85), .Y(n97) );
  INVX4 U71 ( .A(n56), .Y(n245) );
  INVX2 U72 ( .A(n152), .Y(n142) );
  INVX4 U73 ( .A(n10), .Y(n11) );
  NOR2X2 U74 ( .A(n174), .B(n154), .Y(n179) );
  NOR2X2 U75 ( .A(n101), .B(n208), .Y(n202) );
  NAND3X1 U76 ( .A(n225), .B(n226), .C(n71), .Y(n220) );
  NAND2BX2 U77 ( .AN(A[11]), .B(B[11]), .Y(n214) );
  NAND2X1 U78 ( .A(n24), .B(n61), .Y(n209) );
  NAND2BX1 U79 ( .AN(B[12]), .B(A[12]), .Y(n143) );
  NAND4X1 U80 ( .A(n161), .B(n56), .C(n57), .D(n58), .Y(n52) );
  NAND2BX4 U81 ( .AN(A[10]), .B(B[10]), .Y(n207) );
  NAND2BX2 U82 ( .AN(B[3]), .B(A[3]), .Y(n63) );
  NAND2XL U83 ( .A(n71), .B(n192), .Y(n187) );
  NAND3X2 U84 ( .A(n186), .B(n187), .C(n188), .Y(n183) );
  NAND4BX2 U85 ( .AN(n240), .B(n74), .C(n75), .D(n232), .Y(n239) );
  NAND3X2 U86 ( .A(n9), .B(n107), .C(n15), .Y(n103) );
  NAND4X2 U87 ( .A(n104), .B(n103), .C(n102), .D(n22), .Y(n100) );
  INVX3 U88 ( .A(B[1]), .Y(n250) );
  NAND4BX4 U89 ( .AN(n249), .B(n106), .C(n250), .D(n2), .Y(n61) );
  NAND2BXL U90 ( .AN(A[5]), .B(B[5]), .Y(n242) );
  NAND2BX2 U91 ( .AN(B[6]), .B(A[6]), .Y(n246) );
  INVX1 U92 ( .A(A[2]), .Y(n10) );
  OR2X4 U93 ( .A(n51), .B(n52), .Y(n12) );
  NAND2X4 U94 ( .A(n12), .B(n53), .Y(n48) );
  NAND2BX2 U95 ( .AN(A[1]), .B(B[1]), .Y(n118) );
  INVX4 U96 ( .A(n223), .Y(n211) );
  INVX4 U97 ( .A(B[4]), .Y(n199) );
  NAND2BX2 U98 ( .AN(A[6]), .B(B[6]), .Y(n243) );
  AOI21X4 U99 ( .A0(n95), .A1(n242), .B0(n97), .Y(n94) );
  NOR3BX1 U100 ( .AN(n59), .B(n247), .C(n248), .Y(n235) );
  INVX4 U101 ( .A(A[1]), .Y(n249) );
  NAND2X1 U102 ( .A(n57), .B(n56), .Y(n228) );
  OAI2BB1X2 U103 ( .A0N(n80), .A1N(n246), .B0(n56), .Y(n77) );
  INVX4 U104 ( .A(n88), .Y(n95) );
  CLKINVX3 U105 ( .A(n121), .Y(n119) );
  NOR3BX2 U106 ( .AN(n59), .B(n36), .C(n37), .Y(n51) );
  NOR4X1 U107 ( .A(n193), .B(n78), .C(n31), .D(n194), .Y(n192) );
  NAND2BX4 U108 ( .AN(A[8]), .B(B[8]), .Y(n68) );
  NAND2BX1 U109 ( .AN(A[8]), .B(B[8]), .Y(n231) );
  NAND3BX2 U110 ( .AN(n105), .B(n106), .C(n107), .Y(n104) );
  NOR2X4 U111 ( .A(n237), .B(n238), .Y(n236) );
  INVX2 U112 ( .A(n73), .Y(n17) );
  NAND2BX2 U113 ( .AN(B[2]), .B(A[2]), .Y(n117) );
  NAND3X1 U114 ( .A(n250), .B(n14), .C(n106), .Y(n102) );
  OAI21X4 U115 ( .A0(n174), .A1(n180), .B0(n181), .Y(n177) );
  NAND3X1 U116 ( .A(n215), .B(n13), .C(n216), .Y(n213) );
  NAND2BX4 U117 ( .AN(n13), .B(n7), .Y(n50) );
  NAND2X2 U118 ( .A(n71), .B(n27), .Y(n28) );
  BUFX8 U119 ( .A(B[9]), .Y(n13) );
  NAND2X2 U120 ( .A(n62), .B(n22), .Y(n247) );
  INVX2 U121 ( .A(n62), .Y(n208) );
  CLKINVX8 U122 ( .A(n249), .Y(n14) );
  NOR3X4 U123 ( .A(n17), .B(n18), .C(n19), .Y(n20) );
  NAND2BX2 U124 ( .AN(n199), .B(n85), .Y(n73) );
  NAND4X4 U125 ( .A(n75), .B(n231), .C(n232), .D(n74), .Y(n230) );
  NAND2X1 U126 ( .A(n118), .B(n106), .Y(n116) );
  OAI21X4 U127 ( .A0(n115), .A1(n116), .B0(n117), .Y(n112) );
  AOI21X2 U128 ( .A0(n171), .A1(n172), .B0(n173), .Y(n169) );
  NAND3X2 U129 ( .A(n61), .B(n24), .C(n16), .Y(n87) );
  NAND2X2 U130 ( .A(n223), .B(n49), .Y(n227) );
  NAND2BX2 U131 ( .AN(A[7]), .B(B[7]), .Y(n241) );
  NAND2BX1 U132 ( .AN(B[6]), .B(A[6]), .Y(n84) );
  NOR2X2 U133 ( .A(n142), .B(n185), .Y(n184) );
  OAI21X4 U134 ( .A0(n162), .A1(n198), .B0(n77), .Y(n196) );
  NAND2BX4 U135 ( .AN(B[4]), .B(A[4]), .Y(n88) );
  NOR2BX4 U136 ( .AN(n107), .B(n105), .Y(n251) );
  NOR2X1 U137 ( .A(n78), .B(n31), .Y(n70) );
  NAND2BX4 U138 ( .AN(A[2]), .B(B[2]), .Y(n15) );
  NAND2X4 U139 ( .A(n251), .B(n8), .Y(n16) );
  OAI2BB1X2 U140 ( .A0N(n70), .A1N(n71), .B0(n72), .Y(n64) );
  NAND2BX4 U141 ( .AN(B[8]), .B(A[8]), .Y(n69) );
  BUFX20 U142 ( .A(n33), .Y(DIFF[10]) );
  NAND2X4 U143 ( .A(n24), .B(n61), .Y(n248) );
  INVX8 U144 ( .A(n45), .Y(DIFF[2]) );
  NOR2X4 U145 ( .A(n209), .B(n210), .Y(n201) );
  OAI21X2 U146 ( .A0(n142), .A1(n143), .B0(n144), .Y(n173) );
  NAND2BX2 U147 ( .AN(n199), .B(n85), .Y(n232) );
  BUFX20 U148 ( .A(n256), .Y(DIFF[5]) );
  AOI2BB1X4 U149 ( .A0N(B[2]), .A1N(n99), .B0(n100), .Y(n92) );
  OAI2BB1X4 U150 ( .A0N(n57), .A1N(n71), .B0(n88), .Y(n109) );
  INVX8 U151 ( .A(n41), .Y(DIFF[14]) );
  NAND2BX4 U152 ( .AN(B[1]), .B(n14), .Y(n121) );
  NOR2X4 U153 ( .A(n114), .B(n124), .Y(n252) );
  NAND2BX4 U154 ( .AN(A[10]), .B(B[10]), .Y(n223) );
  INVX4 U155 ( .A(n75), .Y(n19) );
  CLKINVX8 U156 ( .A(n162), .Y(n75) );
  BUFX20 U157 ( .A(n253), .Y(DIFF[9]) );
  OR2X2 U158 ( .A(A[4]), .B(n199), .Y(n21) );
  NAND2X4 U159 ( .A(n21), .B(n56), .Y(n78) );
  NAND2X4 U160 ( .A(n151), .B(n152), .Y(n174) );
  BUFX20 U161 ( .A(n254), .Y(DIFF[8]) );
  XOR2X4 U162 ( .A(n233), .B(n34), .Y(n33) );
  NAND2X4 U163 ( .A(n26), .B(n38), .Y(n29) );
  NAND2X4 U164 ( .A(n28), .B(n29), .Y(DIFF[4]) );
  NAND2BX4 U165 ( .AN(B[10]), .B(A[10]), .Y(n215) );
  INVX1 U166 ( .A(n68), .Y(n67) );
  AND2X4 U167 ( .A(n107), .B(n121), .Y(n43) );
  NOR2X2 U168 ( .A(n191), .B(n154), .Y(n190) );
  NAND2BX1 U169 ( .AN(B[14]), .B(A[14]), .Y(n141) );
  NAND2X4 U170 ( .A(n96), .B(n91), .Y(n31) );
  NAND2X4 U171 ( .A(n58), .B(n49), .Y(n240) );
  INVX2 U172 ( .A(n77), .Y(n76) );
  NAND2BX1 U173 ( .AN(B[13]), .B(A[13]), .Y(n144) );
  NAND2BX1 U174 ( .AN(B[11]), .B(A[11]), .Y(n153) );
  NAND2X4 U175 ( .A(n145), .B(n196), .Y(n180) );
  XNOR2X4 U176 ( .A(n172), .B(n32), .Y(DIFF[12]) );
  NOR2XL U177 ( .A(n224), .B(n211), .Y(n34) );
  NAND2BX4 U178 ( .AN(A[5]), .B(B[5]), .Y(n96) );
  NAND2BX4 U179 ( .AN(A[6]), .B(B[6]), .Y(n91) );
  XNOR2X4 U180 ( .A(n122), .B(n123), .Y(n45) );
  NAND2X4 U181 ( .A(n44), .B(n180), .Y(n172) );
  XOR2X4 U182 ( .A(n42), .B(n175), .Y(n41) );
  AOI21XL U183 ( .A0(n222), .A1(n223), .B0(n224), .Y(n221) );
  NAND2XL U184 ( .A(n24), .B(n61), .Y(n37) );
  NAND2BX4 U185 ( .AN(A[12]), .B(B[12]), .Y(n151) );
  INVX2 U186 ( .A(A[11]), .Y(n206) );
  NAND2BX4 U187 ( .AN(A[14]), .B(B[14]), .Y(n138) );
  NAND2BXL U188 ( .AN(B[15]), .B(A[15]), .Y(n137) );
  NOR2X1 U189 ( .A(n66), .B(n67), .Y(n65) );
  NOR2X2 U190 ( .A(n227), .B(n228), .Y(n226) );
  INVXL U191 ( .A(n164), .Y(n155) );
  XOR2X4 U192 ( .A(n217), .B(n218), .Y(n40) );
  AND2X2 U193 ( .A(n141), .B(n138), .Y(n42) );
  XOR2X4 U194 ( .A(n120), .B(n43), .Y(n257) );
  AND3X4 U195 ( .A(n153), .B(n154), .C(n182), .Y(n44) );
  NOR2X1 U196 ( .A(n136), .B(n167), .Y(n166) );
  INVX1 U197 ( .A(n137), .Y(n167) );
  INVX1 U198 ( .A(n144), .Y(n185) );
  INVX1 U199 ( .A(n151), .Y(n191) );
  NAND4BXL U200 ( .AN(n136), .B(n138), .C(n151), .D(n152), .Y(n147) );
  INVX1 U201 ( .A(n215), .Y(n224) );
  NAND3BXL U202 ( .AN(n162), .B(n163), .C(n74), .Y(n156) );
  NAND2XL U203 ( .A(B[4]), .B(n85), .Y(n163) );
  OAI21XL U204 ( .A0(n148), .A1(n149), .B0(n150), .Y(n130) );
  INVX1 U205 ( .A(n147), .Y(n150) );
  NAND2XL U206 ( .A(n153), .B(n154), .Y(n149) );
  AOI31XL U207 ( .A0(n155), .A1(n156), .A2(n157), .B0(n158), .Y(n148) );
  AOI21X1 U208 ( .A0(n138), .A1(n139), .B0(n140), .Y(n135) );
  INVX1 U209 ( .A(n141), .Y(n140) );
  OAI21XL U210 ( .A0(n159), .A1(n160), .B0(n146), .Y(n157) );
  NAND2XL U211 ( .A(n24), .B(n61), .Y(n159) );
  INVXL U212 ( .A(n50), .Y(n222) );
  AOI2BB1X1 U213 ( .A0N(n132), .A1N(n133), .B0(n134), .Y(n131) );
  OAI21XL U214 ( .A0(n135), .A1(n136), .B0(n137), .Y(n134) );
  NAND2XL U215 ( .A(n145), .B(n146), .Y(n133) );
  INVX1 U216 ( .A(n138), .Y(n170) );
  INVX1 U217 ( .A(n120), .Y(n125) );
  XNOR2X1 U218 ( .A(B[16]), .B(A[16]), .Y(n129) );
  NAND2X1 U219 ( .A(n130), .B(n131), .Y(n128) );
  NAND2BX1 U220 ( .AN(A[15]), .B(B[15]), .Y(n168) );
  NAND2X1 U221 ( .A(n108), .B(n127), .Y(DIFF[0]) );
  NAND2BX1 U222 ( .AN(n127), .B(n108), .Y(n120) );
  INVX1 U223 ( .A(n127), .Y(n105) );
  NAND2BX1 U224 ( .AN(B[0]), .B(A[0]), .Y(n108) );
  NAND2BX1 U225 ( .AN(A[0]), .B(B[0]), .Y(n127) );
  BUFX20 U226 ( .A(n255), .Y(DIFF[7]) );
  INVXL U227 ( .A(n11), .Y(n99) );
  NAND2XL U228 ( .A(n62), .B(n22), .Y(n160) );
  OAI21X2 U229 ( .A0(n125), .A1(n126), .B0(n121), .Y(n122) );
  INVX2 U230 ( .A(n118), .Y(n126) );
  AND3X1 U231 ( .A(n161), .B(n56), .C(n57), .Y(n146) );
  NOR2BX4 U232 ( .AN(n117), .B(n124), .Y(n123) );
  XOR2X4 U233 ( .A(n48), .B(n4), .Y(n253) );
  NOR2BX4 U234 ( .AN(n54), .B(n55), .Y(n53) );
  XOR2X4 U235 ( .A(n64), .B(n65), .Y(n254) );
  XOR2X4 U236 ( .A(n79), .B(n3), .Y(n255) );
  OAI21X4 U237 ( .A0(n81), .A1(n82), .B0(n83), .Y(n79) );
  OAI21X4 U238 ( .A0(n92), .A1(n93), .B0(n94), .Y(n89) );
  XOR2X4 U239 ( .A(n109), .B(n110), .Y(n256) );
  XOR2X4 U240 ( .A(n112), .B(n113), .Y(DIFF[3]) );
  NOR2X4 U241 ( .A(n101), .B(n114), .Y(n113) );
  XOR2X4 U242 ( .A(n165), .B(n166), .Y(DIFF[15]) );
  OAI21X4 U243 ( .A0(n169), .A1(n170), .B0(n141), .Y(n165) );
  CLKINVX3 U244 ( .A(n173), .Y(n181) );
  XOR2X4 U245 ( .A(n183), .B(n184), .Y(DIFF[13]) );
  NAND2BX4 U246 ( .AN(A[13]), .B(B[13]), .Y(n152) );
  CLKINVX3 U247 ( .A(n158), .Y(n145) );
  NAND3BX4 U248 ( .AN(n194), .B(n200), .C(n49), .Y(n158) );
  OAI2BB1X4 U249 ( .A0N(n201), .A1N(n202), .B0(n203), .Y(n182) );
  NOR2X4 U250 ( .A(n204), .B(n205), .Y(n203) );
  OAI2BB1X4 U251 ( .A0N(n206), .A1N(B[11]), .B0(n207), .Y(n194) );
  NAND4BX4 U252 ( .AN(n211), .B(n212), .C(n213), .D(n214), .Y(n154) );
  NAND3BX4 U253 ( .AN(n219), .B(n220), .C(n221), .Y(n217) );
  NAND4BX4 U254 ( .AN(n248), .B(n59), .C(n62), .D(n22), .Y(n71) );
  NAND2X4 U255 ( .A(n230), .B(n69), .Y(n55) );
  NAND3X4 U256 ( .A(n241), .B(n96), .C(n243), .Y(n162) );
  NAND2X4 U257 ( .A(n85), .B(n244), .Y(n74) );
  NAND2BX4 U258 ( .AN(B[5]), .B(A[5]), .Y(n85) );
  NAND2X4 U259 ( .A(n164), .B(n68), .Y(n54) );
  OAI21X4 U260 ( .A0(n245), .A1(n246), .B0(n80), .Y(n164) );
  NAND4BX4 U261 ( .AN(n108), .B(n107), .C(n15), .D(n2), .Y(n62) );
  NAND2X4 U262 ( .A(n251), .B(n252), .Y(n59) );
  NAND2BX4 U263 ( .AN(A[2]), .B(B[2]), .Y(n106) );
  NAND2BX4 U264 ( .AN(A[3]), .B(B[3]), .Y(n98) );
  NAND2BX4 U265 ( .AN(A[1]), .B(B[1]), .Y(n107) );
  NAND2BX4 U266 ( .AN(A[7]), .B(B[7]), .Y(n56) );
  NAND2BX4 U267 ( .AN(A[4]), .B(B[4]), .Y(n57) );
  NAND2BX4 U268 ( .AN(A[9]), .B(B[9]), .Y(n49) );
  NAND2BX4 U269 ( .AN(A[8]), .B(B[8]), .Y(n58) );
endmodule


module butterfly_DW01_sub_114 ( A, B, DIFF );
  input [16:0] A;
  input [16:0] B;
  output [16:0] DIFF;
  wire   n204, n205, n206, n207, n208, n209, n210, n1, n2, n3, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n30, n31, n32, n33, n34, n35, n36, n37, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203;

  NAND4BX1 U3 ( .AN(n133), .B(n5), .C(n134), .D(n127), .Y(n120) );
  NAND2X4 U4 ( .A(n93), .B(n37), .Y(n92) );
  NAND3X4 U5 ( .A(n37), .B(n95), .C(n1), .Y(n90) );
  BUFX3 U6 ( .A(n74), .Y(n1) );
  NOR2BX2 U7 ( .AN(n2), .B(n86), .Y(n78) );
  CLKINVX3 U8 ( .A(n159), .Y(n119) );
  AOI21X4 U9 ( .A0(n194), .A1(n96), .B0(n195), .Y(n193) );
  OAI21X4 U10 ( .A0(n196), .A1(n188), .B0(n45), .Y(n195) );
  INVX2 U11 ( .A(B[7]), .Y(n198) );
  BUFX20 U12 ( .A(n208), .Y(DIFF[6]) );
  INVX4 U13 ( .A(n75), .Y(n94) );
  CLKINVX3 U14 ( .A(n158), .Y(n139) );
  OAI21X4 U15 ( .A0(n145), .A1(n153), .B0(n154), .Y(n152) );
  BUFX20 U16 ( .A(n50), .Y(n2) );
  OAI21X4 U17 ( .A0(n81), .A1(n82), .B0(n83), .Y(n65) );
  INVX4 U18 ( .A(n9), .Y(n81) );
  BUFX16 U19 ( .A(n55), .Y(n3) );
  NAND2X4 U20 ( .A(n75), .B(n76), .Y(n178) );
  INVX8 U21 ( .A(n101), .Y(n104) );
  XOR2X4 U22 ( .A(n111), .B(n112), .Y(DIFF[16]) );
  NAND4BX4 U23 ( .AN(n57), .B(n44), .C(n183), .D(n173), .Y(n159) );
  BUFX12 U24 ( .A(n204), .Y(DIFF[15]) );
  INVX1 U25 ( .A(n62), .Y(n60) );
  NAND2X4 U26 ( .A(n182), .B(n62), .Y(n53) );
  AND2X4 U27 ( .A(n46), .B(n62), .Y(n32) );
  NAND2BX4 U28 ( .AN(B[7]), .B(A[7]), .Y(n62) );
  NAND2BX4 U29 ( .AN(n104), .B(n102), .Y(n100) );
  NAND2XL U30 ( .A(n26), .B(n75), .Y(n79) );
  NOR2X2 U31 ( .A(n175), .B(n176), .Y(n168) );
  NOR2BX2 U32 ( .AN(B[9]), .B(A[9]), .Y(n175) );
  INVX3 U33 ( .A(n76), .Y(n93) );
  NAND2BX4 U34 ( .AN(B[3]), .B(n10), .Y(n76) );
  BUFX8 U35 ( .A(n128), .Y(n5) );
  CLKINVX3 U36 ( .A(n183), .Y(n172) );
  NAND2BX4 U37 ( .AN(A[11]), .B(B[11]), .Y(n183) );
  NOR2X1 U38 ( .A(n139), .B(n172), .Y(n184) );
  NOR2X1 U39 ( .A(n165), .B(n129), .Y(n166) );
  INVX1 U40 ( .A(n46), .Y(n56) );
  INVX1 U41 ( .A(n173), .Y(n171) );
  BUFX3 U42 ( .A(A[3]), .Y(n10) );
  CLKINVX3 U43 ( .A(n82), .Y(n89) );
  CLKINVX3 U44 ( .A(n189), .Y(n196) );
  AOI21X1 U45 ( .A0(n190), .A1(n173), .B0(n191), .Y(n185) );
  INVX1 U46 ( .A(n45), .Y(n190) );
  NOR2X1 U47 ( .A(n139), .B(n140), .Y(n167) );
  NAND2BX2 U48 ( .AN(B[8]), .B(A[8]), .Y(n46) );
  NAND2X2 U49 ( .A(n164), .B(n157), .Y(n163) );
  INVX1 U50 ( .A(n121), .Y(n133) );
  OR2X2 U51 ( .A(n18), .B(n19), .Y(n147) );
  NOR2X1 U52 ( .A(n156), .B(n157), .Y(n18) );
  NAND2BX1 U53 ( .AN(A[14]), .B(B[14]), .Y(n128) );
  INVX1 U54 ( .A(n120), .Y(n118) );
  INVX1 U55 ( .A(n142), .Y(n123) );
  INVX4 U56 ( .A(n153), .Y(n140) );
  INVX1 U57 ( .A(n67), .Y(n66) );
  INVX3 U58 ( .A(n68), .Y(n14) );
  NAND2XL U59 ( .A(n9), .B(n68), .Y(n86) );
  INVX8 U60 ( .A(n14), .Y(n13) );
  AND2X2 U61 ( .A(n64), .B(n67), .Y(n6) );
  NAND2BX2 U62 ( .AN(B[11]), .B(A[11]), .Y(n158) );
  OAI21X4 U63 ( .A0(n72), .A1(n73), .B0(n74), .Y(n84) );
  OR2X2 U64 ( .A(n56), .B(n57), .Y(n34) );
  XNOR2X4 U65 ( .A(n141), .B(n7), .Y(n204) );
  OR2X2 U66 ( .A(n133), .B(n123), .Y(n7) );
  BUFX3 U67 ( .A(A[1]), .Y(n8) );
  CLKINVX8 U68 ( .A(n107), .Y(n72) );
  NAND3X2 U69 ( .A(n85), .B(n99), .C(n107), .Y(n95) );
  CLKBUFX20 U70 ( .A(n207), .Y(DIFF[7]) );
  NAND2BX4 U71 ( .AN(A[5]), .B(B[5]), .Y(n9) );
  NAND2BX2 U72 ( .AN(A[5]), .B(B[5]), .Y(n69) );
  OAI21X1 U73 ( .A0(n72), .A1(n73), .B0(n74), .Y(n70) );
  NAND2BX4 U74 ( .AN(A[7]), .B(B[7]), .Y(n203) );
  NAND2BX4 U75 ( .AN(A[2]), .B(B[2]), .Y(n74) );
  NAND3BX2 U76 ( .AN(B[4]), .B(A[4]), .C(n69), .Y(n197) );
  OAI2BB1X4 U77 ( .A0N(n11), .A1N(n12), .B0(n63), .Y(n58) );
  NAND2X2 U78 ( .A(n27), .B(n28), .Y(n11) );
  AND4X1 U79 ( .A(n13), .B(n9), .C(n2), .D(n64), .Y(n12) );
  NAND2X4 U80 ( .A(n32), .B(n137), .Y(n189) );
  NAND2XL U81 ( .A(n44), .B(n45), .Y(n43) );
  NAND2BX2 U82 ( .AN(A[9]), .B(B[9]), .Y(n44) );
  NAND2BX4 U83 ( .AN(B[9]), .B(A[9]), .Y(n45) );
  AND2X4 U84 ( .A(n67), .B(n83), .Y(n36) );
  NAND3BX2 U85 ( .AN(n145), .B(n5), .C(n146), .Y(n144) );
  NAND2X4 U86 ( .A(n94), .B(n37), .Y(n91) );
  NAND4BBX2 U87 ( .AN(n49), .BN(n188), .C(n173), .D(n96), .Y(n187) );
  BUFX20 U88 ( .A(n205), .Y(DIFF[10]) );
  NOR2X1 U89 ( .A(n159), .B(n165), .Y(n162) );
  NAND4BX2 U90 ( .AN(n49), .B(n2), .C(n51), .D(n52), .Y(n48) );
  AOI21XL U91 ( .A0(n131), .A1(n132), .B0(n120), .Y(n113) );
  NAND3X2 U92 ( .A(n1), .B(n2), .C(n95), .Y(n138) );
  AND3X4 U93 ( .A(n76), .B(n84), .C(n71), .Y(n26) );
  AND2X2 U94 ( .A(n70), .B(n71), .Y(n28) );
  NAND2X4 U95 ( .A(n143), .B(n144), .Y(n141) );
  NAND2X1 U96 ( .A(n74), .B(n180), .Y(n179) );
  NOR2X4 U97 ( .A(n155), .B(n147), .Y(n154) );
  NAND2BX2 U98 ( .AN(B[4]), .B(A[4]), .Y(n82) );
  XOR2X4 U99 ( .A(n193), .B(n192), .Y(n205) );
  NOR2BX2 U100 ( .AN(n13), .B(n89), .Y(n97) );
  BUFX20 U101 ( .A(n209), .Y(DIFF[4]) );
  AOI21XL U102 ( .A0(n138), .A1(n76), .B0(n49), .Y(n135) );
  NAND2X2 U103 ( .A(n2), .B(n76), .Y(n98) );
  INVX20 U104 ( .A(n30), .Y(DIFF[5]) );
  AND2X2 U105 ( .A(n75), .B(n76), .Y(n27) );
  NOR2X4 U106 ( .A(n72), .B(n106), .Y(n25) );
  NAND2X4 U107 ( .A(n71), .B(n100), .Y(n24) );
  NOR2X4 U108 ( .A(n171), .B(n172), .Y(n170) );
  NAND3X1 U109 ( .A(n53), .B(n51), .C(n54), .Y(n47) );
  OAI21X4 U110 ( .A0(A[7]), .A1(n198), .B0(n64), .Y(n182) );
  BUFX20 U111 ( .A(n210), .Y(DIFF[2]) );
  BUFX20 U112 ( .A(n23), .Y(DIFF[3]) );
  NAND3BX4 U113 ( .AN(n49), .B(n52), .C(n2), .Y(n177) );
  INVX4 U114 ( .A(n203), .Y(n61) );
  BUFX20 U115 ( .A(n206), .Y(DIFF[9]) );
  NAND2BX4 U116 ( .AN(n182), .B(n181), .Y(n137) );
  NAND2X4 U117 ( .A(n36), .B(n197), .Y(n181) );
  AOI21X2 U118 ( .A0(n64), .A1(n65), .B0(n66), .Y(n63) );
  AND2X4 U119 ( .A(n68), .B(n2), .Y(n37) );
  NAND2X2 U120 ( .A(n134), .B(n127), .Y(n145) );
  NAND2BX4 U121 ( .AN(A[2]), .B(B[2]), .Y(n101) );
  NAND2BX4 U122 ( .AN(B[2]), .B(A[2]), .Y(n99) );
  XNOR2X4 U123 ( .A(n42), .B(n43), .Y(n206) );
  NAND3X2 U124 ( .A(n48), .B(n47), .C(n46), .Y(n42) );
  NAND2X4 U125 ( .A(n44), .B(n51), .Y(n188) );
  NAND2BX4 U126 ( .AN(B[2]), .B(A[2]), .Y(n71) );
  NAND3X4 U127 ( .A(n2), .B(n101), .C(n201), .Y(n75) );
  XOR2X4 U128 ( .A(n102), .B(n103), .Y(n210) );
  NAND2BX4 U129 ( .AN(B[1]), .B(n8), .Y(n107) );
  INVX4 U130 ( .A(n85), .Y(n73) );
  NAND2BX4 U131 ( .AN(n110), .B(n200), .Y(n85) );
  INVX1 U132 ( .A(n65), .Y(n80) );
  NAND2BX4 U133 ( .AN(B[13]), .B(A[13]), .Y(n130) );
  NAND2BX4 U134 ( .AN(B[12]), .B(A[12]), .Y(n157) );
  AOI21XL U135 ( .A0(n147), .A1(n5), .B0(n148), .Y(n143) );
  INVXL U136 ( .A(n130), .Y(n19) );
  NAND2BX4 U137 ( .AN(A[12]), .B(B[12]), .Y(n134) );
  NAND2BX4 U138 ( .AN(A[13]), .B(B[13]), .Y(n127) );
  INVX2 U139 ( .A(n25), .Y(n20) );
  NAND2BX4 U140 ( .AN(B[6]), .B(A[6]), .Y(n67) );
  NAND2BX4 U141 ( .AN(B[5]), .B(A[5]), .Y(n83) );
  OAI21X4 U142 ( .A0(n105), .A1(n106), .B0(n107), .Y(n102) );
  OAI2BB1X4 U143 ( .A0N(n78), .A1N(n79), .B0(n80), .Y(n77) );
  XOR2X4 U144 ( .A(n77), .B(n6), .Y(n208) );
  NOR2BX4 U145 ( .AN(n99), .B(n104), .Y(n103) );
  NAND2BX4 U146 ( .AN(n181), .B(n62), .Y(n54) );
  NAND2X1 U147 ( .A(n109), .B(n110), .Y(n108) );
  NAND2X4 U148 ( .A(n108), .B(n20), .Y(n21) );
  NAND2X2 U149 ( .A(n105), .B(n25), .Y(n22) );
  NAND2X4 U150 ( .A(n21), .B(n22), .Y(DIFF[1]) );
  XNOR2X4 U151 ( .A(n24), .B(n98), .Y(n23) );
  NAND2XL U152 ( .A(n126), .B(n5), .Y(n149) );
  AOI21X4 U153 ( .A0(n151), .A1(n3), .B0(n152), .Y(n150) );
  AOI21X4 U154 ( .A0(n162), .A1(n3), .B0(n163), .Y(n161) );
  NAND2BX4 U155 ( .AN(A[4]), .B(B[4]), .Y(n68) );
  NOR2X2 U156 ( .A(n145), .B(n158), .Y(n155) );
  NAND2BX4 U157 ( .AN(A[8]), .B(B[8]), .Y(n51) );
  NAND2XL U158 ( .A(n85), .B(n107), .Y(n180) );
  XNOR2X4 U159 ( .A(n35), .B(n184), .Y(DIFF[11]) );
  NAND2XL U160 ( .A(n127), .B(n5), .Y(n125) );
  XOR2X4 U161 ( .A(n87), .B(n31), .Y(n30) );
  OR2X2 U162 ( .A(n88), .B(n81), .Y(n31) );
  XOR2X4 U163 ( .A(n3), .B(n34), .Y(n33) );
  INVX8 U164 ( .A(n33), .Y(DIFF[8]) );
  INVX1 U165 ( .A(n51), .Y(n57) );
  NOR2XL U166 ( .A(n139), .B(n140), .Y(n131) );
  OAI21XL U167 ( .A0(n135), .A1(n136), .B0(n119), .Y(n132) );
  NAND2XL U168 ( .A(n137), .B(n62), .Y(n136) );
  INVXL U169 ( .A(n49), .Y(n117) );
  AND3X4 U170 ( .A(n185), .B(n186), .C(n187), .Y(n35) );
  NAND2X1 U171 ( .A(n127), .B(n130), .Y(n160) );
  NAND2XL U172 ( .A(n173), .B(n174), .Y(n192) );
  NOR2X1 U173 ( .A(n188), .B(n49), .Y(n194) );
  NOR2X1 U174 ( .A(n145), .B(n159), .Y(n151) );
  INVX1 U175 ( .A(n127), .Y(n156) );
  INVX1 U176 ( .A(n108), .Y(n105) );
  INVX1 U177 ( .A(n134), .Y(n165) );
  INVX1 U178 ( .A(n157), .Y(n129) );
  NAND2X1 U179 ( .A(n115), .B(n116), .Y(n114) );
  AOI21X1 U180 ( .A0(n121), .A1(n122), .B0(n123), .Y(n115) );
  OAI21XL U181 ( .A0(n124), .A1(n125), .B0(n126), .Y(n122) );
  NAND3BXL U182 ( .AN(n188), .B(n173), .C(n189), .Y(n186) );
  NOR2BXL U183 ( .AN(n130), .B(n129), .Y(n124) );
  INVX1 U184 ( .A(n83), .Y(n88) );
  NAND2BXL U185 ( .AN(B[8]), .B(A[8]), .Y(n176) );
  INVX1 U186 ( .A(n126), .Y(n148) );
  INVXL U187 ( .A(n174), .Y(n191) );
  XOR2X1 U188 ( .A(B[16]), .B(A[16]), .Y(n112) );
  NOR2X1 U189 ( .A(n113), .B(n114), .Y(n111) );
  NAND2BX1 U190 ( .AN(B[14]), .B(A[14]), .Y(n126) );
  NAND2BX1 U191 ( .AN(B[15]), .B(A[15]), .Y(n142) );
  NAND2BX1 U192 ( .AN(A[15]), .B(B[15]), .Y(n121) );
  NAND2X1 U193 ( .A(n110), .B(n202), .Y(DIFF[0]) );
  INVX1 U194 ( .A(n202), .Y(n109) );
  NAND2BX1 U195 ( .AN(B[0]), .B(A[0]), .Y(n110) );
  NAND2BX1 U196 ( .AN(A[0]), .B(B[0]), .Y(n202) );
  NAND4XL U197 ( .A(n94), .B(n117), .C(n118), .D(n119), .Y(n116) );
  INVX8 U198 ( .A(n200), .Y(n106) );
  XOR2X4 U199 ( .A(n58), .B(n59), .Y(n207) );
  NOR2X4 U200 ( .A(n60), .B(n61), .Y(n59) );
  NAND4BX4 U201 ( .AN(n89), .B(n91), .C(n90), .D(n92), .Y(n87) );
  XOR2X4 U202 ( .A(n96), .B(n97), .Y(n209) );
  XOR2X4 U203 ( .A(n149), .B(n150), .Y(DIFF[14]) );
  XOR2X4 U204 ( .A(n160), .B(n161), .Y(DIFF[13]) );
  OAI21X4 U205 ( .A0(n139), .A1(n140), .B0(n134), .Y(n164) );
  XOR2X4 U206 ( .A(n146), .B(n166), .Y(DIFF[12]) );
  OAI2BB1X4 U207 ( .A0N(n119), .A1N(n3), .B0(n167), .Y(n146) );
  OAI21X4 U208 ( .A0(n168), .A1(n169), .B0(n170), .Y(n153) );
  NAND2X4 U209 ( .A(n45), .B(n174), .Y(n169) );
  OAI2BB1X4 U210 ( .A0N(n53), .A1N(n54), .B0(n177), .Y(n55) );
  NAND3BX4 U211 ( .AN(n178), .B(n179), .C(n71), .Y(n52) );
  NAND2X4 U212 ( .A(n199), .B(n138), .Y(n96) );
  NOR2X4 U213 ( .A(n94), .B(n93), .Y(n199) );
  NOR2X4 U214 ( .A(n106), .B(n109), .Y(n201) );
  NAND2BX4 U215 ( .AN(A[1]), .B(B[1]), .Y(n200) );
  NAND2BX4 U216 ( .AN(A[3]), .B(B[3]), .Y(n50) );
  NAND4BX4 U217 ( .AN(n61), .B(n13), .C(n64), .D(n9), .Y(n49) );
  NAND2BX4 U218 ( .AN(A[6]), .B(B[6]), .Y(n64) );
  NAND2BX4 U219 ( .AN(B[10]), .B(A[10]), .Y(n174) );
  NAND2BX4 U220 ( .AN(A[10]), .B(B[10]), .Y(n173) );
endmodule


module butterfly_DW01_add_129 ( A, B, SUM );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  wire   n156, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155;

  AOI21X1 U2 ( .A0(n107), .A1(n63), .B0(n93), .Y(n103) );
  NAND2X2 U3 ( .A(n21), .B(n154), .Y(n107) );
  INVX4 U4 ( .A(n58), .Y(n56) );
  NOR2X2 U5 ( .A(n51), .B(n55), .Y(n152) );
  INVX4 U6 ( .A(n60), .Y(n55) );
  OAI211X1 U7 ( .A0(n75), .A1(n76), .B0(n73), .C0(n67), .Y(n154) );
  NAND2BX4 U8 ( .AN(n92), .B(n35), .Y(n96) );
  CLKBUFX3 U9 ( .A(n37), .Y(n1) );
  OAI21X4 U10 ( .A0(n7), .A1(n126), .B0(n90), .Y(n119) );
  BUFX16 U11 ( .A(n116), .Y(n25) );
  NOR2BX1 U12 ( .AN(n57), .B(n55), .Y(n59) );
  NOR2BX2 U13 ( .AN(n90), .B(n7), .Y(n128) );
  AOI21X1 U14 ( .A0(n31), .A1(n32), .B0(n33), .Y(n30) );
  NAND4X4 U15 ( .A(n22), .B(n23), .C(n111), .D(n112), .Y(n94) );
  NAND3X2 U16 ( .A(A[5]), .B(B[5]), .C(n49), .Y(n106) );
  BUFX16 U17 ( .A(n156), .Y(SUM[8]) );
  XOR2X4 U18 ( .A(n38), .B(n39), .Y(n156) );
  NAND2X1 U19 ( .A(n100), .B(n101), .Y(n98) );
  NOR2X4 U20 ( .A(n87), .B(n88), .Y(n82) );
  NAND2X2 U21 ( .A(n89), .B(n90), .Y(n88) );
  AOI21X1 U22 ( .A0(B[7]), .A1(A[7]), .B0(n41), .Y(n44) );
  INVX8 U23 ( .A(n99), .Y(n133) );
  OAI2BB1X4 U24 ( .A0N(n47), .A1N(n49), .B0(n46), .Y(n43) );
  CLKINVX3 U25 ( .A(n71), .Y(n75) );
  OAI21X4 U26 ( .A0(n55), .A1(n56), .B0(n57), .Y(n53) );
  NAND2X2 U27 ( .A(B[4]), .B(A[4]), .Y(n57) );
  NAND2X4 U28 ( .A(n17), .B(n18), .Y(SUM[10]) );
  NAND2X4 U29 ( .A(n15), .B(n16), .Y(n18) );
  OAI21X4 U30 ( .A0(n25), .A1(n129), .B0(n91), .Y(n127) );
  XNOR2X4 U31 ( .A(n127), .B(n5), .Y(SUM[13]) );
  NOR2X2 U32 ( .A(n110), .B(n94), .Y(n78) );
  NAND2X1 U33 ( .A(B[7]), .B(A[7]), .Y(n105) );
  INVX1 U34 ( .A(n133), .Y(n6) );
  NAND2X2 U35 ( .A(A[13]), .B(B[13]), .Y(n90) );
  AND2X2 U36 ( .A(n105), .B(n106), .Y(n20) );
  AND2X2 U37 ( .A(n70), .B(n155), .Y(n21) );
  OR2X2 U38 ( .A(A[4]), .B(B[4]), .Y(n60) );
  INVX1 U39 ( .A(n141), .Y(n15) );
  NAND2X2 U40 ( .A(B[2]), .B(A[2]), .Y(n67) );
  INVX1 U41 ( .A(n128), .Y(n5) );
  INVX1 U42 ( .A(n124), .Y(n26) );
  NAND2X1 U43 ( .A(n141), .B(n144), .Y(n17) );
  INVX1 U44 ( .A(n144), .Y(n16) );
  NAND2X1 U45 ( .A(n2), .B(n25), .Y(n12) );
  XOR2X2 U46 ( .A(n47), .B(n48), .Y(SUM[6]) );
  NOR2BX1 U47 ( .AN(n46), .B(n45), .Y(n48) );
  NOR2X4 U48 ( .A(n57), .B(n51), .Y(n150) );
  AND2X2 U49 ( .A(n112), .B(n91), .Y(n2) );
  NAND2X2 U50 ( .A(n63), .B(n107), .Y(n58) );
  NOR2BX4 U51 ( .AN(n35), .B(n92), .Y(n130) );
  INVX2 U52 ( .A(n36), .Y(n149) );
  INVXL U53 ( .A(n110), .Y(n3) );
  INVX3 U54 ( .A(n136), .Y(n110) );
  XNOR2X4 U55 ( .A(n77), .B(n4), .Y(SUM[16]) );
  XNOR2X4 U56 ( .A(B[16]), .B(A[16]), .Y(n4) );
  NAND2X2 U57 ( .A(B[9]), .B(A[9]), .Y(n37) );
  OR2X4 U58 ( .A(B[11]), .B(A[11]), .Y(n24) );
  INVX1 U59 ( .A(n25), .Y(n11) );
  OR2X2 U60 ( .A(n145), .B(n32), .Y(n9) );
  INVX1 U61 ( .A(n35), .Y(n41) );
  NAND2X4 U62 ( .A(n35), .B(n49), .Y(n153) );
  AOI21X4 U63 ( .A0(n147), .A1(n42), .B0(n148), .Y(n146) );
  INVX8 U64 ( .A(n108), .Y(n51) );
  NOR2X4 U65 ( .A(A[13]), .B(B[13]), .Y(n7) );
  NAND4X4 U66 ( .A(n20), .B(n46), .C(n109), .D(n32), .Y(n131) );
  NAND2X4 U67 ( .A(n138), .B(n36), .Y(n134) );
  OAI21X1 U68 ( .A0(n149), .A1(n29), .B0(n1), .Y(n148) );
  NOR2X2 U69 ( .A(n6), .B(n98), .Y(n97) );
  NAND2XL U70 ( .A(n3), .B(n101), .Y(n139) );
  NOR2BX2 U71 ( .AN(n89), .B(n121), .Y(n124) );
  NOR2X4 U72 ( .A(n153), .B(n56), .Y(n151) );
  NAND2X4 U73 ( .A(n37), .B(n29), .Y(n138) );
  NAND2X4 U74 ( .A(n150), .B(n49), .Y(n109) );
  NAND2X4 U75 ( .A(n112), .B(n111), .Y(n122) );
  NAND2X2 U76 ( .A(n85), .B(n86), .Y(n83) );
  INVX4 U77 ( .A(n86), .Y(n115) );
  OR2X4 U78 ( .A(A[15]), .B(B[15]), .Y(n86) );
  OR2X4 U79 ( .A(A[15]), .B(B[15]), .Y(n23) );
  NAND2XL U80 ( .A(n143), .B(n137), .Y(n144) );
  NAND2X4 U81 ( .A(n24), .B(n137), .Y(n135) );
  NAND2X1 U82 ( .A(B[11]), .B(A[11]), .Y(n101) );
  OR2X4 U83 ( .A(n121), .B(n122), .Y(n117) );
  NAND2X1 U84 ( .A(B[15]), .B(A[15]), .Y(n84) );
  NAND2X2 U85 ( .A(B[6]), .B(A[6]), .Y(n46) );
  INVX4 U86 ( .A(n81), .Y(n80) );
  OAI21X4 U87 ( .A0(n82), .A1(n83), .B0(n84), .Y(n81) );
  BUFX3 U88 ( .A(n44), .Y(n8) );
  AOI21X2 U89 ( .A0(n85), .A1(n119), .B0(n120), .Y(n118) );
  OAI21X2 U90 ( .A0(n95), .A1(n96), .B0(n97), .Y(n79) );
  NOR2BX2 U91 ( .AN(n35), .B(n145), .Y(n147) );
  NAND2X2 U92 ( .A(n36), .B(n34), .Y(n145) );
  NAND2X2 U93 ( .A(n10), .B(n11), .Y(n13) );
  OAI21X2 U94 ( .A0(n41), .A1(n31), .B0(n32), .Y(n38) );
  NOR2X2 U95 ( .A(n7), .B(n91), .Y(n87) );
  NAND2X4 U96 ( .A(n9), .B(n146), .Y(n141) );
  NAND2X4 U97 ( .A(n12), .B(n13), .Y(SUM[12]) );
  INVX1 U98 ( .A(n2), .Y(n10) );
  OAI21X4 U99 ( .A0(n50), .A1(n51), .B0(n52), .Y(n47) );
  INVX4 U100 ( .A(n53), .Y(n50) );
  OR2X4 U101 ( .A(A[8]), .B(B[8]), .Y(n34) );
  XOR2X4 U102 ( .A(n27), .B(n28), .Y(SUM[9]) );
  NOR2BX2 U103 ( .AN(n29), .B(n30), .Y(n28) );
  XOR2X4 U104 ( .A(n43), .B(n8), .Y(SUM[7]) );
  XOR2X2 U105 ( .A(n53), .B(n54), .Y(SUM[5]) );
  INVX1 U106 ( .A(n119), .Y(n125) );
  NAND2X2 U107 ( .A(B[12]), .B(A[12]), .Y(n91) );
  OAI21X4 U108 ( .A0(n25), .A1(n122), .B0(n125), .Y(n123) );
  NOR2BXL U109 ( .AN(n67), .B(n66), .Y(n69) );
  OAI21XL U110 ( .A0(n65), .A1(n66), .B0(n67), .Y(n61) );
  OR2X2 U111 ( .A(A[3]), .B(B[3]), .Y(n155) );
  NAND2XL U112 ( .A(B[3]), .B(A[3]), .Y(n63) );
  NOR2XL U113 ( .A(A[0]), .B(B[0]), .Y(n19) );
  INVX4 U114 ( .A(n42), .Y(n31) );
  INVXL U115 ( .A(n68), .Y(n65) );
  INVXL U116 ( .A(n89), .Y(n120) );
  INVXL U117 ( .A(n112), .Y(n129) );
  NAND2XL U118 ( .A(n105), .B(n106), .Y(n104) );
  NAND2XL U119 ( .A(n109), .B(n46), .Y(n102) );
  INVXL U120 ( .A(n76), .Y(n72) );
  OR2X4 U121 ( .A(A[2]), .B(B[2]), .Y(n70) );
  NOR2BX1 U122 ( .AN(n76), .B(n19), .Y(SUM[0]) );
  NOR2BX1 U123 ( .AN(n29), .B(n40), .Y(n39) );
  INVX1 U124 ( .A(n34), .Y(n40) );
  INVX1 U125 ( .A(n143), .Y(n142) );
  NOR3X1 U126 ( .A(n102), .B(n103), .C(n104), .Y(n95) );
  NAND4X2 U127 ( .A(n46), .B(n109), .C(n105), .D(n106), .Y(n42) );
  NOR2BXL U128 ( .AN(n52), .B(n51), .Y(n54) );
  XOR2X1 U129 ( .A(n58), .B(n59), .Y(SUM[4]) );
  XOR2X1 U130 ( .A(n61), .B(n62), .Y(SUM[3]) );
  NOR2BX1 U131 ( .AN(n63), .B(n64), .Y(n62) );
  INVX1 U132 ( .A(n155), .Y(n64) );
  XOR2X1 U133 ( .A(n68), .B(n69), .Y(SUM[2]) );
  INVXL U134 ( .A(n49), .Y(n45) );
  INVX1 U135 ( .A(n70), .Y(n66) );
  XOR2X1 U136 ( .A(n72), .B(n74), .Y(SUM[1]) );
  NOR2BXL U137 ( .AN(n73), .B(n75), .Y(n74) );
  NAND3XL U138 ( .A(n108), .B(n60), .C(n49), .Y(n93) );
  OAI2BB1X1 U139 ( .A0N(n71), .A1N(n72), .B0(n73), .Y(n68) );
  NAND2XL U140 ( .A(n34), .B(n35), .Y(n33) );
  OR2X2 U141 ( .A(A[14]), .B(B[14]), .Y(n22) );
  NAND2XL U142 ( .A(A[12]), .B(B[12]), .Y(n126) );
  NAND4X2 U143 ( .A(n136), .B(n137), .C(n36), .D(n34), .Y(n92) );
  NAND2X2 U144 ( .A(B[14]), .B(A[14]), .Y(n89) );
  NAND2X1 U145 ( .A(B[0]), .B(A[0]), .Y(n76) );
  NAND2X1 U146 ( .A(B[1]), .B(A[1]), .Y(n73) );
  NAND2XL U147 ( .A(B[5]), .B(A[5]), .Y(n52) );
  NAND2XL U148 ( .A(B[10]), .B(A[10]), .Y(n100) );
  NAND2XL U149 ( .A(B[10]), .B(A[10]), .Y(n143) );
  AOI21X4 U150 ( .A0(n137), .A1(n141), .B0(n142), .Y(n140) );
  NAND2XL U151 ( .A(n36), .B(n1), .Y(n27) );
  XNOR2X4 U152 ( .A(n123), .B(n26), .Y(SUM[14]) );
  OAI2BB1X4 U153 ( .A0N(n78), .A1N(n79), .B0(n80), .Y(n77) );
  XOR2X4 U154 ( .A(n113), .B(n114), .Y(SUM[15]) );
  NOR2BX4 U155 ( .AN(n84), .B(n115), .Y(n114) );
  OAI21X4 U156 ( .A0(n25), .A1(n117), .B0(n118), .Y(n113) );
  CLKINVX3 U157 ( .A(n85), .Y(n121) );
  OR2X4 U158 ( .A(A[14]), .B(B[14]), .Y(n85) );
  OR2X4 U159 ( .A(A[13]), .B(B[13]), .Y(n111) );
  AOI21X4 U160 ( .A0(n130), .A1(n131), .B0(n132), .Y(n116) );
  OAI211X2 U161 ( .A0(n110), .A1(n100), .B0(n133), .C0(n101), .Y(n132) );
  NOR2X4 U162 ( .A(n134), .B(n135), .Y(n99) );
  OR2X4 U163 ( .A(A[12]), .B(B[12]), .Y(n112) );
  XOR2X4 U164 ( .A(n139), .B(n140), .Y(SUM[11]) );
  OR2X4 U165 ( .A(A[11]), .B(B[11]), .Y(n136) );
  OR2X4 U166 ( .A(A[10]), .B(B[10]), .Y(n137) );
  NAND2X4 U167 ( .A(B[8]), .B(A[8]), .Y(n29) );
  NAND2X4 U168 ( .A(n151), .B(n152), .Y(n32) );
  OR2X4 U169 ( .A(A[5]), .B(B[5]), .Y(n108) );
  OR2X4 U170 ( .A(A[1]), .B(B[1]), .Y(n71) );
  OR2X4 U171 ( .A(A[6]), .B(B[6]), .Y(n49) );
  OR2X4 U172 ( .A(A[7]), .B(B[7]), .Y(n35) );
  OR2X4 U173 ( .A(A[9]), .B(B[9]), .Y(n36) );
endmodule


module butterfly_DW01_add_147 ( A, B, SUM );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  wire   n194, n195, n196, n197, n198, n199, n1, n2, n3, n4, n5, n6, n8, n9,
         n10, n11, n12, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193;

  BUFX16 U2 ( .A(n194), .Y(SUM[13]) );
  NOR2X1 U3 ( .A(n116), .B(n119), .Y(n149) );
  OAI2BB1X4 U4 ( .A0N(n49), .A1N(n4), .B0(n82), .Y(n78) );
  INVX3 U5 ( .A(n89), .Y(n87) );
  NAND2X2 U6 ( .A(n123), .B(n124), .Y(n150) );
  NAND2BX2 U7 ( .AN(n164), .B(n163), .Y(n123) );
  AOI2BB1X4 U8 ( .A0N(n70), .A1N(n71), .B0(n72), .Y(n66) );
  XOR2X4 U9 ( .A(n141), .B(n151), .Y(n195) );
  INVX8 U10 ( .A(n4), .Y(n5) );
  CLKINVX8 U11 ( .A(n81), .Y(n4) );
  NAND2XL U12 ( .A(B[4]), .B(A[4]), .Y(n77) );
  NAND4BX1 U13 ( .AN(n155), .B(n45), .C(n40), .D(n173), .Y(n178) );
  NAND2X2 U14 ( .A(n40), .B(n45), .Y(n174) );
  NOR2BX1 U15 ( .AN(n40), .B(n39), .Y(n57) );
  XOR2X4 U16 ( .A(n97), .B(n98), .Y(SUM[16]) );
  AND2X4 U17 ( .A(n68), .B(n69), .Y(n23) );
  NOR2BX4 U18 ( .AN(n69), .B(n86), .Y(n85) );
  CLKINVX2 U19 ( .A(n69), .Y(n10) );
  NAND2X4 U20 ( .A(B[3]), .B(n34), .Y(n69) );
  OAI21X1 U21 ( .A0(n116), .A1(n137), .B0(n110), .Y(n148) );
  INVX2 U22 ( .A(n142), .Y(n116) );
  NOR3X4 U23 ( .A(n41), .B(n42), .C(n43), .Y(n38) );
  NAND2X2 U24 ( .A(B[10]), .B(A[10]), .Y(n164) );
  OAI21X2 U25 ( .A0(n116), .A1(n146), .B0(n147), .Y(n144) );
  NAND2XL U26 ( .A(n124), .B(n163), .Y(n165) );
  CLKINVX3 U27 ( .A(n59), .Y(n19) );
  NOR2X1 U28 ( .A(n117), .B(n118), .Y(n99) );
  OAI21XL U29 ( .A0(n103), .A1(n27), .B0(n104), .Y(n102) );
  NOR2X1 U30 ( .A(n148), .B(n149), .Y(n147) );
  INVX1 U31 ( .A(n150), .Y(n137) );
  OR2X2 U32 ( .A(A[12]), .B(B[12]), .Y(n142) );
  NAND3BX1 U33 ( .AN(n39), .B(n37), .C(n168), .Y(n170) );
  NOR2BX2 U34 ( .AN(n172), .B(n127), .Y(n169) );
  OAI21XL U35 ( .A0(n160), .A1(n36), .B0(n164), .Y(n167) );
  INVX4 U36 ( .A(n91), .Y(n95) );
  CLKINVX3 U37 ( .A(n54), .Y(n81) );
  NOR3X2 U38 ( .A(n154), .B(n155), .C(n156), .Y(n153) );
  INVX1 U39 ( .A(n45), .Y(n156) );
  INVX1 U40 ( .A(n46), .Y(n64) );
  NOR2BX2 U41 ( .AN(n45), .B(n60), .Y(n59) );
  NAND2X2 U42 ( .A(B[8]), .B(A[8]), .Y(n40) );
  NAND2X1 U43 ( .A(B[9]), .B(A[9]), .Y(n36) );
  NAND2X2 U44 ( .A(n157), .B(n158), .Y(n112) );
  NOR2X2 U45 ( .A(n160), .B(n161), .Y(n157) );
  NAND2X1 U46 ( .A(B[14]), .B(A[14]), .Y(n108) );
  OR2X2 U47 ( .A(A[14]), .B(B[14]), .Y(n105) );
  NOR2X1 U48 ( .A(A[15]), .B(B[15]), .Y(n27) );
  INVX4 U49 ( .A(n187), .Y(n86) );
  CLKINVX3 U50 ( .A(n90), .Y(n17) );
  NOR2BX2 U51 ( .AN(n88), .B(n11), .Y(n90) );
  OAI21X1 U52 ( .A0(n99), .A1(n100), .B0(n101), .Y(n97) );
  OAI21X2 U53 ( .A0(n133), .A1(n134), .B0(n108), .Y(n131) );
  AOI21X1 U54 ( .A0(n6), .A1(n56), .B0(n136), .Y(n133) );
  NAND2X2 U55 ( .A(n46), .B(n82), .Y(n189) );
  AND2X4 U56 ( .A(n46), .B(n82), .Y(n18) );
  AND2X2 U57 ( .A(n36), .B(n37), .Y(n1) );
  INVX1 U58 ( .A(n112), .Y(n6) );
  AND2X2 U59 ( .A(n129), .B(n130), .Y(n2) );
  AND2X2 U60 ( .A(n164), .B(n168), .Y(n3) );
  NAND2X4 U61 ( .A(n6), .B(n56), .Y(n146) );
  INVX1 U62 ( .A(n52), .Y(n60) );
  INVX8 U63 ( .A(n9), .Y(SUM[1]) );
  INVX1 U64 ( .A(A[4]), .Y(n70) );
  XOR2X4 U65 ( .A(n75), .B(n8), .Y(SUM[6]) );
  AND2X1 U66 ( .A(n63), .B(n53), .Y(n8) );
  CLKINVX4 U67 ( .A(n152), .Y(n179) );
  INVX1 U68 ( .A(n55), .Y(n80) );
  NOR2X2 U69 ( .A(n18), .B(n48), .Y(n154) );
  OAI2BB1X2 U70 ( .A0N(n91), .A1N(n92), .B0(n93), .Y(n89) );
  NAND2X2 U71 ( .A(B[2]), .B(A[2]), .Y(n88) );
  XOR2X4 U72 ( .A(n96), .B(n94), .Y(n9) );
  NAND2X2 U73 ( .A(B[7]), .B(A[7]), .Y(n45) );
  INVX8 U74 ( .A(n21), .Y(SUM[11]) );
  NOR2BX4 U75 ( .AN(n68), .B(n10), .Y(n25) );
  BUFX3 U76 ( .A(B[2]), .Y(n12) );
  AND2X4 U77 ( .A(B[1]), .B(A[1]), .Y(n188) );
  BUFX2 U78 ( .A(A[3]), .Y(n34) );
  BUFX20 U79 ( .A(n196), .Y(SUM[9]) );
  AOI21X1 U80 ( .A0(n46), .A1(n47), .B0(n48), .Y(n42) );
  NOR2BX2 U81 ( .AN(n46), .B(n80), .Y(n79) );
  NAND2X2 U82 ( .A(n52), .B(n53), .Y(n182) );
  NOR2X4 U83 ( .A(A[6]), .B(B[6]), .Y(n192) );
  NAND2X2 U84 ( .A(n73), .B(n74), .Y(n72) );
  OAI21X4 U85 ( .A0(n38), .A1(n39), .B0(n40), .Y(n35) );
  INVX4 U86 ( .A(n44), .Y(n155) );
  AND2X4 U87 ( .A(n23), .B(n24), .Y(n76) );
  AND3X2 U88 ( .A(n74), .B(n77), .C(n73), .Y(n24) );
  NOR2X4 U89 ( .A(n191), .B(n192), .Y(n190) );
  NOR2X2 U90 ( .A(A[7]), .B(B[7]), .Y(n191) );
  NOR2X4 U91 ( .A(A[2]), .B(B[2]), .Y(n11) );
  XOR2X2 U92 ( .A(n49), .B(n83), .Y(n199) );
  NAND2X2 U93 ( .A(n54), .B(n55), .Y(n181) );
  BUFX16 U94 ( .A(n195), .Y(SUM[12]) );
  NAND2X4 U95 ( .A(n73), .B(n74), .Y(n183) );
  BUFX20 U96 ( .A(n198), .Y(SUM[5]) );
  NAND2X4 U97 ( .A(B[4]), .B(A[4]), .Y(n82) );
  NOR2X2 U98 ( .A(n155), .B(n174), .Y(n172) );
  NAND3X1 U99 ( .A(n137), .B(n138), .C(n119), .Y(n136) );
  NOR2X4 U100 ( .A(n39), .B(n159), .Y(n158) );
  INVX8 U101 ( .A(n171), .Y(n39) );
  NAND2X4 U102 ( .A(n54), .B(n55), .Y(n67) );
  BUFX20 U103 ( .A(n197), .Y(SUM[7]) );
  AOI21X2 U104 ( .A0(n169), .A1(n152), .B0(n170), .Y(n166) );
  NAND2X4 U105 ( .A(n49), .B(n180), .Y(n152) );
  NAND2XL U106 ( .A(B[15]), .B(A[15]), .Y(n104) );
  NOR2BX4 U107 ( .AN(n82), .B(n5), .Y(n83) );
  NAND2X2 U108 ( .A(B[1]), .B(A[1]), .Y(n93) );
  NOR2BXL U109 ( .AN(n110), .B(n116), .Y(n151) );
  INVX3 U110 ( .A(n168), .Y(n160) );
  NAND2X1 U111 ( .A(B[13]), .B(A[13]), .Y(n111) );
  XNOR2X4 U112 ( .A(n56), .B(n57), .Y(n20) );
  INVXL U113 ( .A(n53), .Y(n62) );
  NOR3BX4 U114 ( .AN(n49), .B(n50), .C(n51), .Y(n41) );
  XOR2X4 U115 ( .A(n78), .B(n79), .Y(n198) );
  INVXL U116 ( .A(n123), .Y(n122) );
  OR2X4 U117 ( .A(A[8]), .B(B[8]), .Y(n171) );
  OR2X4 U118 ( .A(n166), .B(n167), .Y(n22) );
  AND2X1 U119 ( .A(n142), .B(n143), .Y(n26) );
  XOR2X4 U120 ( .A(n139), .B(n140), .Y(SUM[14]) );
  INVXL U121 ( .A(n124), .Y(n121) );
  NAND2X2 U122 ( .A(B[12]), .B(A[12]), .Y(n110) );
  NOR2X1 U123 ( .A(n60), .B(n62), .Y(n130) );
  NOR2XL U124 ( .A(n80), .B(n5), .Y(n129) );
  NAND2XL U125 ( .A(n44), .B(n45), .Y(n43) );
  XNOR2X4 U126 ( .A(n175), .B(n3), .Y(n14) );
  INVX8 U127 ( .A(n14), .Y(SUM[10]) );
  XNOR2X4 U128 ( .A(n84), .B(n85), .Y(n15) );
  INVX8 U129 ( .A(n15), .Y(SUM[3]) );
  XOR2X2 U130 ( .A(n89), .B(n17), .Y(n16) );
  INVX8 U131 ( .A(n16), .Y(SUM[2]) );
  XNOR2X4 U132 ( .A(n58), .B(n19), .Y(n197) );
  INVX8 U133 ( .A(n20), .Y(SUM[8]) );
  NAND2XL U134 ( .A(n119), .B(n120), .Y(n118) );
  AOI31XL U135 ( .A0(n44), .A1(n125), .A2(n126), .B0(n112), .Y(n117) );
  NOR2X1 U136 ( .A(n121), .B(n122), .Y(n120) );
  NOR2BXL U137 ( .AN(n45), .B(n127), .Y(n126) );
  NAND2XL U138 ( .A(n52), .B(n53), .Y(n51) );
  NAND2XL U139 ( .A(n54), .B(n55), .Y(n50) );
  NAND2XL U140 ( .A(n37), .B(n171), .Y(n177) );
  XOR2X4 U141 ( .A(n165), .B(n22), .Y(n21) );
  NOR2BX1 U142 ( .AN(n111), .B(n109), .Y(n145) );
  INVX1 U143 ( .A(B[4]), .Y(n71) );
  NOR2BX1 U144 ( .AN(n104), .B(n27), .Y(n132) );
  OAI21XL U145 ( .A0(n26), .A1(n135), .B0(n105), .Y(n134) );
  OAI21XL U146 ( .A0(n109), .A1(n110), .B0(n111), .Y(n106) );
  INVX1 U147 ( .A(n105), .Y(n115) );
  OAI21XL U148 ( .A0(n128), .A1(n183), .B0(n2), .Y(n125) );
  NAND2XL U149 ( .A(n68), .B(n69), .Y(n128) );
  NAND2XL U150 ( .A(B[4]), .B(A[4]), .Y(n47) );
  NAND2X1 U151 ( .A(n113), .B(n114), .Y(n100) );
  NOR2XL U152 ( .A(n27), .B(n115), .Y(n114) );
  NOR2XL U153 ( .A(n109), .B(n116), .Y(n113) );
  INVX1 U154 ( .A(n102), .Y(n101) );
  AOI21X1 U155 ( .A0(n105), .A1(n106), .B0(n107), .Y(n103) );
  INVX1 U156 ( .A(n108), .Y(n107) );
  XOR2X1 U157 ( .A(B[16]), .B(A[16]), .Y(n98) );
  NAND2X1 U158 ( .A(B[11]), .B(A[11]), .Y(n124) );
  INVX1 U159 ( .A(n96), .Y(n92) );
  AND2X2 U160 ( .A(n96), .B(n193), .Y(SUM[0]) );
  OR2X2 U161 ( .A(A[0]), .B(B[0]), .Y(n193) );
  NAND2X1 U162 ( .A(B[0]), .B(A[0]), .Y(n96) );
  NAND3BX4 U163 ( .AN(n183), .B(n68), .C(n69), .Y(n49) );
  BUFX16 U164 ( .A(n199), .Y(SUM[4]) );
  OAI21X4 U165 ( .A0(n87), .A1(n11), .B0(n88), .Y(n84) );
  NOR3X2 U166 ( .A(n159), .B(n160), .C(n161), .Y(n162) );
  NAND3X4 U167 ( .A(A[2]), .B(n12), .C(n187), .Y(n73) );
  NAND3X4 U168 ( .A(n186), .B(n187), .C(n188), .Y(n74) );
  XOR2X4 U169 ( .A(n35), .B(n1), .Y(n196) );
  OAI21X4 U170 ( .A0(n61), .A1(n62), .B0(n63), .Y(n58) );
  NOR2X4 U171 ( .A(n65), .B(n64), .Y(n61) );
  AOI21X4 U172 ( .A0(n25), .A1(n66), .B0(n67), .Y(n65) );
  OAI21X4 U173 ( .A0(n76), .A1(n67), .B0(n46), .Y(n75) );
  NOR2BX4 U174 ( .AN(n93), .B(n95), .Y(n94) );
  XOR2X4 U175 ( .A(n131), .B(n132), .Y(SUM[15]) );
  NOR2BX4 U176 ( .AN(n108), .B(n115), .Y(n140) );
  OAI2BB1X4 U177 ( .A0N(n26), .A1N(n141), .B0(n138), .Y(n139) );
  CLKINVX3 U178 ( .A(n135), .Y(n138) );
  OAI21X4 U179 ( .A0(n109), .A1(n110), .B0(n111), .Y(n135) );
  XOR2X4 U180 ( .A(n144), .B(n145), .Y(n194) );
  CLKINVX3 U181 ( .A(n143), .Y(n109) );
  OR2X4 U182 ( .A(A[13]), .B(B[13]), .Y(n143) );
  NAND3BX4 U183 ( .AN(n150), .B(n146), .C(n119), .Y(n141) );
  NAND2X4 U184 ( .A(n152), .B(n153), .Y(n56) );
  OAI2BB1X4 U185 ( .A0N(n36), .A1N(n40), .B0(n162), .Y(n119) );
  CLKINVX3 U186 ( .A(n163), .Y(n161) );
  CLKINVX3 U187 ( .A(n37), .Y(n159) );
  CLKINVX3 U188 ( .A(n173), .Y(n127) );
  OR2X4 U189 ( .A(A[11]), .B(B[11]), .Y(n163) );
  OR2X4 U190 ( .A(A[10]), .B(B[10]), .Y(n168) );
  OAI21X4 U191 ( .A0(n176), .A1(n177), .B0(n36), .Y(n175) );
  OR2X4 U192 ( .A(A[9]), .B(B[9]), .Y(n37) );
  NOR2X4 U193 ( .A(n178), .B(n179), .Y(n176) );
  NOR2X4 U194 ( .A(n181), .B(n182), .Y(n180) );
  OR2X4 U195 ( .A(A[6]), .B(B[6]), .Y(n53) );
  OR2X4 U196 ( .A(A[5]), .B(B[5]), .Y(n55) );
  OR2X4 U197 ( .A(A[4]), .B(B[4]), .Y(n54) );
  NAND2X4 U198 ( .A(n185), .B(n184), .Y(n68) );
  NOR2X4 U199 ( .A(n86), .B(n11), .Y(n185) );
  NOR2X4 U200 ( .A(n95), .B(n96), .Y(n184) );
  OR2X4 U201 ( .A(B[1]), .B(A[1]), .Y(n91) );
  OR2X4 U202 ( .A(A[2]), .B(B[2]), .Y(n186) );
  OR2X4 U203 ( .A(A[3]), .B(B[3]), .Y(n187) );
  NAND2BX4 U204 ( .AN(n48), .B(n189), .Y(n173) );
  NAND2X4 U205 ( .A(B[5]), .B(A[5]), .Y(n46) );
  OAI21X4 U206 ( .A0(A[5]), .A1(B[5]), .B0(n190), .Y(n48) );
  NAND2BX4 U207 ( .AN(n63), .B(n52), .Y(n44) );
  OR2X4 U208 ( .A(A[7]), .B(B[7]), .Y(n52) );
  NAND2X4 U209 ( .A(B[6]), .B(A[6]), .Y(n63) );
endmodule


module butterfly_DW01_add_145 ( A, B, SUM );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184;

  NAND2XL U2 ( .A(B[13]), .B(A[13]), .Y(n114) );
  NAND3X1 U3 ( .A(n119), .B(n120), .C(n121), .Y(n116) );
  OAI21X4 U4 ( .A0(n23), .A1(n24), .B0(n107), .Y(n91) );
  NAND2X4 U5 ( .A(B[8]), .B(A[8]), .Y(n141) );
  NAND4X2 U6 ( .A(n26), .B(n142), .C(n143), .D(n35), .Y(n103) );
  NOR2BX1 U7 ( .AN(n50), .B(n3), .Y(n54) );
  AND2X4 U8 ( .A(n93), .B(n154), .Y(n25) );
  NAND2X1 U9 ( .A(n144), .B(n45), .Y(n168) );
  AND2X4 U10 ( .A(n144), .B(n45), .Y(n15) );
  CLKINVX3 U11 ( .A(n139), .Y(n172) );
  NAND2X1 U12 ( .A(B[10]), .B(A[10]), .Y(n119) );
  INVX3 U13 ( .A(n39), .Y(n36) );
  OAI2BB1X4 U14 ( .A0N(n48), .A1N(n49), .B0(n50), .Y(n46) );
  NAND4BX4 U15 ( .AN(n14), .B(n21), .C(n56), .D(n95), .Y(n5) );
  NAND2X4 U16 ( .A(n96), .B(n39), .Y(n14) );
  NOR2X2 U17 ( .A(A[3]), .B(B[3]), .Y(n28) );
  NOR2X4 U18 ( .A(A[2]), .B(B[2]), .Y(n27) );
  OAI21X2 U19 ( .A0(n182), .A1(n69), .B0(n183), .Y(n180) );
  NAND3X2 U20 ( .A(n5), .B(n141), .C(n176), .Y(n175) );
  INVX1 U21 ( .A(n3), .Y(n154) );
  INVX1 U22 ( .A(n4), .Y(n96) );
  NAND2X2 U23 ( .A(n147), .B(n148), .Y(n145) );
  NOR2X2 U24 ( .A(n129), .B(n149), .Y(n147) );
  OAI2BB1X2 U25 ( .A0N(n15), .A1N(n16), .B0(n170), .Y(n176) );
  AND3X2 U26 ( .A(n139), .B(n7), .C(n153), .Y(n24) );
  NAND2X1 U27 ( .A(n116), .B(n117), .Y(n97) );
  NOR2X1 U28 ( .A(n118), .B(n104), .Y(n117) );
  NAND4BX1 U29 ( .AN(n100), .B(n101), .C(n102), .D(n103), .Y(n99) );
  INVX1 U30 ( .A(n104), .Y(n102) );
  NOR2X2 U31 ( .A(n105), .B(n106), .Y(n101) );
  NAND2X2 U32 ( .A(B[5]), .B(A[5]), .Y(n50) );
  NOR2X1 U33 ( .A(n3), .B(n4), .Y(n48) );
  NAND3X1 U34 ( .A(n51), .B(n52), .C(n6), .Y(n49) );
  OAI2BB1X1 U35 ( .A0N(n51), .A1N(n52), .B0(n19), .Y(n92) );
  OAI21XL U36 ( .A0(n74), .A1(n75), .B0(n76), .Y(n73) );
  AND2X4 U37 ( .A(B[4]), .B(A[4]), .Y(n1) );
  AND2X2 U38 ( .A(B[2]), .B(A[2]), .Y(n2) );
  NOR2X4 U39 ( .A(A[5]), .B(B[5]), .Y(n3) );
  AND2X4 U40 ( .A(n38), .B(n141), .Y(n165) );
  INVX1 U41 ( .A(n108), .Y(n42) );
  OR2X2 U42 ( .A(A[6]), .B(B[6]), .Y(n20) );
  OR2X2 U43 ( .A(A[7]), .B(B[7]), .Y(n108) );
  NOR2XL U44 ( .A(A[7]), .B(B[7]), .Y(n13) );
  NOR2BX2 U45 ( .AN(n164), .B(n172), .Y(n174) );
  NAND2X1 U46 ( .A(n119), .B(n120), .Y(n23) );
  AND2X2 U47 ( .A(n119), .B(n120), .Y(n138) );
  AND2X2 U48 ( .A(n93), .B(n154), .Y(n21) );
  AOI21XL U49 ( .A0(n92), .A1(n34), .B0(n85), .Y(n89) );
  NAND3X2 U50 ( .A(n166), .B(n165), .C(n167), .Y(n163) );
  NAND4BX2 U51 ( .AN(n126), .B(n127), .C(n128), .D(n103), .Y(n124) );
  AOI21X4 U52 ( .A0(n130), .A1(n131), .B0(n132), .Y(n123) );
  CLKINVX3 U53 ( .A(n177), .Y(n170) );
  NOR2X1 U54 ( .A(A[1]), .B(B[1]), .Y(n182) );
  NOR2X4 U55 ( .A(B[4]), .B(A[4]), .Y(n4) );
  NAND2X2 U56 ( .A(B[3]), .B(A[3]), .Y(n51) );
  OAI22X1 U57 ( .A0(A[8]), .A1(B[8]), .B0(A[7]), .B1(B[7]), .Y(n177) );
  INVX1 U58 ( .A(n77), .Y(n115) );
  NAND2X2 U59 ( .A(B[12]), .B(A[12]), .Y(n84) );
  OR2X4 U60 ( .A(A[12]), .B(B[12]), .Y(n109) );
  OAI21X2 U61 ( .A0(n60), .A1(n27), .B0(n61), .Y(n58) );
  NAND3X2 U62 ( .A(n119), .B(n120), .C(n121), .Y(n130) );
  NOR2BX2 U63 ( .AN(n61), .B(n27), .Y(n63) );
  NOR2X4 U64 ( .A(n28), .B(n27), .Y(n181) );
  INVX4 U65 ( .A(n93), .Y(n44) );
  NAND2BX2 U66 ( .AN(n50), .B(n93), .Y(n171) );
  NAND2X2 U67 ( .A(n34), .B(n35), .Y(n40) );
  NOR2X4 U68 ( .A(n145), .B(n146), .Y(n135) );
  NOR2BX4 U69 ( .AN(n66), .B(n68), .Y(n67) );
  OR2X2 U70 ( .A(A[15]), .B(B[15]), .Y(n78) );
  NAND2X2 U71 ( .A(B[9]), .B(A[9]), .Y(n38) );
  NOR2X1 U72 ( .A(n42), .B(n36), .Y(n148) );
  OAI2BB1X2 U73 ( .A0N(B[9]), .A1N(A[9]), .B0(n141), .Y(n140) );
  NAND3X1 U74 ( .A(n110), .B(n107), .C(n109), .Y(n126) );
  NAND2X4 U75 ( .A(n109), .B(n107), .Y(n118) );
  NOR2BX2 U76 ( .AN(n112), .B(n118), .Y(n131) );
  NAND2XL U77 ( .A(B[2]), .B(A[2]), .Y(n61) );
  OR2X4 U78 ( .A(A[14]), .B(B[14]), .Y(n77) );
  NAND2X2 U79 ( .A(n112), .B(n77), .Y(n104) );
  OR2X2 U80 ( .A(A[9]), .B(B[9]), .Y(n37) );
  NAND2X1 U81 ( .A(n107), .B(n7), .Y(n106) );
  OAI21X2 U82 ( .A0(n168), .A1(n169), .B0(n170), .Y(n167) );
  OR2X1 U83 ( .A(A[1]), .B(B[1]), .Y(n64) );
  OAI2BB1X4 U84 ( .A0N(n7), .A1N(n175), .B0(n38), .Y(n173) );
  NAND2X1 U85 ( .A(n7), .B(n38), .Y(n30) );
  NOR2BX4 U86 ( .AN(n120), .B(n149), .Y(n161) );
  INVX4 U87 ( .A(n56), .Y(n55) );
  OR2X2 U88 ( .A(A[10]), .B(B[10]), .Y(n110) );
  XOR2X2 U89 ( .A(n62), .B(n63), .Y(SUM[2]) );
  NAND4BX4 U90 ( .AN(n14), .B(n21), .C(n56), .D(n95), .Y(n166) );
  OR2X4 U91 ( .A(A[6]), .B(B[6]), .Y(n93) );
  XOR2X4 U92 ( .A(n70), .B(n71), .Y(SUM[16]) );
  NAND4BX4 U93 ( .AN(n13), .B(n25), .C(n96), .D(n56), .Y(n35) );
  XOR2X4 U94 ( .A(n58), .B(n59), .Y(SUM[3]) );
  OAI2BB1X1 U95 ( .A0N(B[7]), .A1N(A[7]), .B0(n171), .Y(n169) );
  AOI21X2 U96 ( .A0(n138), .A1(n121), .B0(n118), .Y(n137) );
  OR2X4 U97 ( .A(A[10]), .B(B[10]), .Y(n139) );
  OR2X4 U98 ( .A(A[8]), .B(B[8]), .Y(n39) );
  NAND2X1 U99 ( .A(n77), .B(n78), .Y(n75) );
  INVX4 U100 ( .A(n112), .Y(n83) );
  OR2X4 U101 ( .A(A[13]), .B(B[13]), .Y(n112) );
  INVX8 U102 ( .A(n107), .Y(n149) );
  OR2X4 U103 ( .A(A[11]), .B(B[11]), .Y(n107) );
  NOR2X4 U104 ( .A(n3), .B(n6), .Y(n179) );
  INVX8 U105 ( .A(n1), .Y(n6) );
  XOR2X4 U106 ( .A(n56), .B(n57), .Y(SUM[4]) );
  NOR2X2 U107 ( .A(n36), .B(n129), .Y(n158) );
  INVX8 U108 ( .A(n7), .Y(n129) );
  BUFX8 U109 ( .A(n37), .Y(n7) );
  NAND2X2 U110 ( .A(n141), .B(n39), .Y(n10) );
  NOR2BX2 U111 ( .AN(n6), .B(n4), .Y(n57) );
  AND2X2 U112 ( .A(n171), .B(n178), .Y(n16) );
  XOR2X4 U113 ( .A(n133), .B(n134), .Y(SUM[13]) );
  OAI2BB1X4 U114 ( .A0N(n135), .A1N(n103), .B0(n136), .Y(n133) );
  INVX1 U115 ( .A(n82), .Y(n132) );
  NOR2BX2 U116 ( .AN(n45), .B(n44), .Y(n47) );
  AND2X2 U117 ( .A(n8), .B(n9), .Y(n19) );
  NOR2X1 U118 ( .A(n4), .B(n94), .Y(n8) );
  NOR2XL U119 ( .A(n44), .B(n3), .Y(n9) );
  XNOR2X4 U120 ( .A(n40), .B(n10), .Y(SUM[8]) );
  NOR2XL U121 ( .A(n83), .B(n88), .Y(n86) );
  XNOR2X4 U122 ( .A(n22), .B(n11), .Y(SUM[15]) );
  AND2X2 U123 ( .A(n76), .B(n78), .Y(n11) );
  INVX4 U124 ( .A(n46), .Y(n43) );
  AND2X1 U125 ( .A(n81), .B(n77), .Y(n12) );
  OAI2BB1X2 U126 ( .A0N(n17), .A1N(n18), .B0(n72), .Y(n70) );
  OR2X2 U127 ( .A(n89), .B(n90), .Y(n17) );
  AND2X2 U128 ( .A(n86), .B(n87), .Y(n18) );
  NOR2BX2 U129 ( .AN(n84), .B(n137), .Y(n136) );
  AND2X1 U130 ( .A(n78), .B(n77), .Y(n87) );
  OAI2BB1X2 U131 ( .A0N(n64), .A1N(n65), .B0(n66), .Y(n62) );
  NAND2XL U132 ( .A(B[15]), .B(A[15]), .Y(n76) );
  NOR2BX1 U133 ( .AN(n82), .B(n83), .Y(n134) );
  NAND2XL U134 ( .A(n39), .B(n108), .Y(n105) );
  INVX1 U135 ( .A(n95), .Y(n94) );
  INVX1 U136 ( .A(n91), .Y(n90) );
  NAND2X1 U137 ( .A(n109), .B(n110), .Y(n100) );
  XNOR2X4 U138 ( .A(n41), .B(n29), .Y(SUM[7]) );
  AND3X4 U139 ( .A(n97), .B(n98), .C(n99), .Y(n22) );
  AOI21X2 U140 ( .A0(n111), .A1(n112), .B0(n113), .Y(n98) );
  INVX1 U141 ( .A(n81), .Y(n113) );
  AOI21X1 U142 ( .A0(n84), .A1(n114), .B0(n115), .Y(n111) );
  OAI2BB1X1 U143 ( .A0N(B[7]), .A1N(A[7]), .B0(n108), .Y(n29) );
  AND2X1 U144 ( .A(n144), .B(n45), .Y(n26) );
  NOR2BX1 U145 ( .AN(n51), .B(n28), .Y(n59) );
  INVX1 U146 ( .A(n62), .Y(n60) );
  NAND2X1 U147 ( .A(B[13]), .B(A[13]), .Y(n82) );
  NOR2XL U148 ( .A(n42), .B(n36), .Y(n127) );
  INVX1 U149 ( .A(n109), .Y(n88) );
  INVX1 U150 ( .A(n73), .Y(n72) );
  NOR2X1 U151 ( .A(n79), .B(n80), .Y(n74) );
  NAND2XL U152 ( .A(n81), .B(n82), .Y(n80) );
  NAND2X1 U153 ( .A(n110), .B(n109), .Y(n146) );
  XOR2X2 U154 ( .A(n65), .B(n67), .Y(SUM[1]) );
  NAND2XL U155 ( .A(B[14]), .B(A[14]), .Y(n81) );
  XOR2X1 U156 ( .A(B[16]), .B(A[16]), .Y(n71) );
  INVX1 U157 ( .A(n69), .Y(n65) );
  AND2X2 U158 ( .A(n69), .B(n184), .Y(SUM[0]) );
  OR2X2 U159 ( .A(A[0]), .B(B[0]), .Y(n184) );
  NAND2X1 U160 ( .A(B[0]), .B(A[0]), .Y(n69) );
  NAND2X4 U161 ( .A(n51), .B(n52), .Y(n56) );
  CLKINVX3 U162 ( .A(n141), .Y(n32) );
  OAI2BB1X1 U163 ( .A0N(B[9]), .A1N(A[9]), .B0(n141), .Y(n153) );
  NAND2XL U164 ( .A(B[10]), .B(A[10]), .Y(n164) );
  NAND2X2 U165 ( .A(B[6]), .B(A[6]), .Y(n45) );
  INVX2 U166 ( .A(n64), .Y(n68) );
  NOR2XL U167 ( .A(n83), .B(n84), .Y(n79) );
  NOR2BX2 U168 ( .AN(n84), .B(n88), .Y(n151) );
  NAND2BX1 U169 ( .AN(n84), .B(n112), .Y(n125) );
  NOR2X2 U170 ( .A(n129), .B(n172), .Y(n162) );
  NAND2X2 U171 ( .A(B[11]), .B(A[11]), .Y(n120) );
  NOR2X2 U172 ( .A(n129), .B(n83), .Y(n128) );
  NAND2XL U173 ( .A(B[7]), .B(A[7]), .Y(n156) );
  OR2X2 U174 ( .A(A[7]), .B(B[7]), .Y(n95) );
  NAND2XL U175 ( .A(B[7]), .B(A[7]), .Y(n178) );
  NAND2XL U176 ( .A(B[7]), .B(A[7]), .Y(n142) );
  NAND2XL U177 ( .A(B[1]), .B(A[1]), .Y(n66) );
  NAND2XL U178 ( .A(B[1]), .B(A[1]), .Y(n183) );
  XOR2X4 U179 ( .A(n30), .B(n31), .Y(SUM[9]) );
  NOR2X4 U180 ( .A(n32), .B(n33), .Y(n31) );
  AOI21X4 U181 ( .A0(n34), .A1(n35), .B0(n36), .Y(n33) );
  OAI21X4 U182 ( .A0(n43), .A1(n44), .B0(n45), .Y(n41) );
  XOR2X4 U183 ( .A(n46), .B(n47), .Y(SUM[6]) );
  XOR2X4 U184 ( .A(n53), .B(n54), .Y(SUM[5]) );
  OAI21X4 U185 ( .A0(n55), .A1(n4), .B0(n6), .Y(n53) );
  XOR2X4 U186 ( .A(n122), .B(n12), .Y(SUM[14]) );
  NAND3X4 U187 ( .A(n123), .B(n124), .C(n125), .Y(n122) );
  NAND3X4 U188 ( .A(n139), .B(n7), .C(n140), .Y(n121) );
  XOR2X4 U189 ( .A(n150), .B(n151), .Y(SUM[12]) );
  OAI2BB1X4 U190 ( .A0N(n152), .A1N(n40), .B0(n91), .Y(n150) );
  NAND2X4 U191 ( .A(n155), .B(n108), .Y(n34) );
  NAND4X2 U192 ( .A(n143), .B(n156), .C(n45), .D(n144), .Y(n155) );
  NAND2BX4 U193 ( .AN(n50), .B(n93), .Y(n143) );
  CLKINVX3 U194 ( .A(n85), .Y(n152) );
  NAND2X4 U195 ( .A(n157), .B(n158), .Y(n85) );
  NOR2X4 U196 ( .A(n149), .B(n159), .Y(n157) );
  CLKINVX3 U197 ( .A(n110), .Y(n159) );
  XOR2X4 U198 ( .A(n160), .B(n161), .Y(SUM[11]) );
  OAI2BB1X4 U199 ( .A0N(n162), .A1N(n163), .B0(n164), .Y(n160) );
  XOR2X4 U200 ( .A(n173), .B(n174), .Y(SUM[10]) );
  NAND2X4 U201 ( .A(n179), .B(n20), .Y(n144) );
  OAI21X4 U202 ( .A0(n2), .A1(n180), .B0(n181), .Y(n52) );
endmodule


module butterfly_DW01_sub_120 ( A, B, DIFF );
  input [16:0] A;
  input [16:0] B;
  output [16:0] DIFF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190;

  INVX1 U3 ( .A(n28), .Y(n1) );
  INVX2 U4 ( .A(n64), .Y(n59) );
  INVX2 U5 ( .A(n31), .Y(n184) );
  OAI2BB1X2 U6 ( .A0N(n25), .A1N(n10), .B0(n162), .Y(n158) );
  OR2X1 U7 ( .A(n45), .B(n15), .Y(n18) );
  NAND2BX2 U8 ( .AN(n182), .B(n183), .Y(n180) );
  AOI21X1 U9 ( .A0(n94), .A1(n118), .B0(n96), .Y(n117) );
  XNOR2X4 U10 ( .A(n20), .B(n52), .Y(DIFF[5]) );
  INVX2 U11 ( .A(n71), .Y(n66) );
  NAND3X1 U12 ( .A(n169), .B(n100), .C(n130), .Y(n132) );
  NAND3X2 U13 ( .A(n137), .B(n26), .C(n31), .Y(n121) );
  XNOR2X2 U14 ( .A(n12), .B(n17), .Y(DIFF[4]) );
  NAND2X2 U15 ( .A(n38), .B(n3), .Y(n4) );
  NAND2X2 U16 ( .A(n2), .B(n39), .Y(n5) );
  NAND2X4 U17 ( .A(n4), .B(n5), .Y(DIFF[7]) );
  CLKINVX4 U18 ( .A(n38), .Y(n2) );
  INVX1 U19 ( .A(n39), .Y(n3) );
  OAI2BB1X4 U20 ( .A0N(n42), .A1N(n43), .B0(n44), .Y(n38) );
  NOR2X2 U21 ( .A(n40), .B(n41), .Y(n39) );
  AOI21X4 U22 ( .A0(n134), .A1(n110), .B0(n135), .Y(n133) );
  NAND2BX4 U23 ( .AN(A[13]), .B(B[13]), .Y(n130) );
  OAI21X4 U24 ( .A0(A[13]), .A1(n123), .B0(n99), .Y(n120) );
  INVXL U25 ( .A(B[13]), .Y(n123) );
  NAND2X2 U26 ( .A(n42), .B(n49), .Y(n155) );
  INVX8 U27 ( .A(n15), .Y(n42) );
  INVX3 U28 ( .A(n174), .Y(n41) );
  NAND2BX2 U29 ( .AN(A[7]), .B(B[7]), .Y(n174) );
  AOI21X2 U30 ( .A0(n116), .A1(n130), .B0(n92), .Y(n129) );
  CLKINVX3 U31 ( .A(n101), .Y(n95) );
  NAND2BX1 U32 ( .AN(A[5]), .B(B[5]), .Y(n173) );
  NAND2X1 U33 ( .A(n104), .B(n44), .Y(n182) );
  NAND2BX1 U34 ( .AN(A[1]), .B(B[1]), .Y(n71) );
  NAND2X2 U35 ( .A(n13), .B(n6), .Y(n14) );
  AOI21X2 U36 ( .A0(n115), .A1(n116), .B0(n117), .Y(n114) );
  INVX1 U37 ( .A(n110), .Y(n7) );
  NAND2BX2 U38 ( .AN(B[11]), .B(A[11]), .Y(n149) );
  NAND2BX2 U39 ( .AN(B[1]), .B(A[1]), .Y(n67) );
  AND2X2 U40 ( .A(n16), .B(B[6]), .Y(n15) );
  NAND2X1 U41 ( .A(n99), .B(n94), .Y(n124) );
  NOR2X1 U42 ( .A(n132), .B(n121), .Y(n126) );
  INVX1 U43 ( .A(n83), .Y(n82) );
  AOI21X1 U44 ( .A0(n85), .A1(n86), .B0(n87), .Y(n78) );
  OAI21XL U45 ( .A0(n89), .A1(n90), .B0(n91), .Y(n86) );
  NOR2X2 U46 ( .A(n28), .B(n29), .Y(n27) );
  NAND2BX2 U47 ( .AN(A[0]), .B(B[0]), .Y(n73) );
  INVX1 U48 ( .A(n50), .Y(n53) );
  AOI21X2 U49 ( .A0(n50), .A1(n36), .B0(n51), .Y(n52) );
  INVX2 U50 ( .A(n104), .Y(n40) );
  NAND3X1 U51 ( .A(n143), .B(n147), .C(n169), .Y(n6) );
  CLKINVX3 U52 ( .A(n103), .Y(n153) );
  NAND4BXL U53 ( .AN(n29), .B(n31), .C(n169), .D(n137), .Y(n157) );
  XOR2X4 U54 ( .A(n74), .B(n75), .Y(DIFF[16]) );
  AOI2BB1X4 U55 ( .A0N(n7), .A1N(n8), .B0(n111), .Y(n109) );
  OR3X2 U56 ( .A(n121), .B(n122), .C(n120), .Y(n8) );
  NAND2BX2 U57 ( .AN(B[8]), .B(A[8]), .Y(n37) );
  NAND2BX2 U58 ( .AN(A[9]), .B(B[9]), .Y(n143) );
  INVX1 U59 ( .A(n143), .Y(n142) );
  AOI21X1 U60 ( .A0(n141), .A1(B[10]), .B0(n142), .Y(n138) );
  AND2X1 U61 ( .A(n49), .B(n48), .Y(n20) );
  INVX4 U62 ( .A(n30), .Y(n28) );
  NAND2X1 U63 ( .A(n169), .B(n100), .Y(n122) );
  NAND2BX4 U64 ( .AN(B[4]), .B(A[4]), .Y(n54) );
  NAND3BX4 U65 ( .AN(n187), .B(n188), .C(n189), .Y(n106) );
  AND2X4 U66 ( .A(B[7]), .B(n9), .Y(n172) );
  CLKINVX20 U67 ( .A(A[7]), .Y(n9) );
  INVX2 U68 ( .A(B[12]), .Y(n136) );
  OAI21X4 U69 ( .A0(n11), .A1(n128), .B0(n129), .Y(n127) );
  NAND2X1 U70 ( .A(n32), .B(n37), .Y(n139) );
  INVX2 U71 ( .A(n90), .Y(n116) );
  OAI21X4 U72 ( .A0(n11), .A1(n113), .B0(n114), .Y(n111) );
  NAND2BX2 U73 ( .AN(A[12]), .B(B[12]), .Y(n100) );
  INVX1 U74 ( .A(n99), .Y(n96) );
  NAND2X2 U75 ( .A(n130), .B(n119), .Y(n128) );
  NAND2BX2 U76 ( .AN(B[14]), .B(A[14]), .Y(n94) );
  NAND2BX2 U77 ( .AN(B[6]), .B(A[6]), .Y(n44) );
  NAND2BX1 U78 ( .AN(n73), .B(n72), .Y(n68) );
  OAI21X4 U79 ( .A0(n65), .A1(n66), .B0(n67), .Y(n58) );
  CLKINVX3 U80 ( .A(n68), .Y(n65) );
  NAND2BX2 U81 ( .AN(B[0]), .B(A[0]), .Y(n72) );
  NAND3X2 U82 ( .A(n67), .B(n72), .C(n64), .Y(n188) );
  NAND2X1 U83 ( .A(n104), .B(n105), .Y(n152) );
  NAND2BX4 U84 ( .AN(A[14]), .B(B[14]), .Y(n99) );
  AOI21X2 U85 ( .A0(n57), .A1(n58), .B0(n59), .Y(n56) );
  AOI21X2 U86 ( .A0(n35), .A1(n12), .B0(n30), .Y(n34) );
  NAND2X2 U87 ( .A(n57), .B(n60), .Y(n187) );
  NOR2X4 U88 ( .A(n51), .B(n36), .Y(n46) );
  OAI21X4 U89 ( .A0(n161), .A1(n177), .B0(n178), .Y(n175) );
  INVX4 U90 ( .A(n25), .Y(n161) );
  AOI21X2 U91 ( .A0(n179), .A1(n180), .B0(n181), .Y(n178) );
  NAND2X2 U92 ( .A(n78), .B(n79), .Y(n77) );
  NAND4X1 U93 ( .A(n80), .B(n35), .C(n81), .D(n82), .Y(n79) );
  AOI21X4 U94 ( .A0(n25), .A1(n26), .B0(n27), .Y(n24) );
  NOR3X2 U95 ( .A(n184), .B(n41), .C(n29), .Y(n179) );
  CLKINVX2 U96 ( .A(n140), .Y(n13) );
  XNOR2X4 U97 ( .A(n19), .B(n133), .Y(DIFF[13]) );
  NAND2BX2 U98 ( .AN(A[15]), .B(B[15]), .Y(n101) );
  NAND2BX1 U99 ( .AN(B[15]), .B(A[15]), .Y(n88) );
  XOR2X4 U100 ( .A(n23), .B(n24), .Y(DIFF[9]) );
  AND3X1 U101 ( .A(n31), .B(n26), .C(n169), .Y(n10) );
  NAND2BX4 U102 ( .AN(A[10]), .B(B[10]), .Y(n169) );
  NAND4BX2 U103 ( .AN(n95), .B(n99), .C(n100), .D(n130), .Y(n83) );
  INVX2 U104 ( .A(n94), .Y(n93) );
  NOR2X2 U105 ( .A(n92), .B(n93), .Y(n91) );
  NOR2X4 U106 ( .A(n163), .B(n164), .Y(n162) );
  AOI21XL U107 ( .A0(n97), .A1(n98), .B0(n83), .Y(n76) );
  OAI21X2 U108 ( .A0(n112), .A1(n131), .B0(n90), .Y(n135) );
  NAND4BX2 U109 ( .AN(n107), .B(n50), .C(n49), .D(n42), .Y(n84) );
  NOR2BX2 U110 ( .AN(B[7]), .B(A[7]), .Y(n107) );
  BUFX8 U111 ( .A(n112), .Y(n11) );
  NAND2X4 U112 ( .A(n45), .B(n174), .Y(n103) );
  NAND3X2 U113 ( .A(n31), .B(n26), .C(n169), .Y(n168) );
  INVX4 U114 ( .A(n169), .Y(n165) );
  INVX3 U115 ( .A(n84), .Y(n35) );
  AOI21X4 U116 ( .A0(n139), .A1(n138), .B0(n140), .Y(n112) );
  INVX4 U117 ( .A(n54), .Y(n51) );
  NOR2BX4 U118 ( .AN(n173), .B(n172), .Y(n171) );
  BUFX8 U119 ( .A(n36), .Y(n12) );
  NAND2BX4 U120 ( .AN(B[3]), .B(A[3]), .Y(n61) );
  OAI2BB1X4 U121 ( .A0N(n12), .A1N(n185), .B0(n37), .Y(n25) );
  AOI21X2 U122 ( .A0(n167), .A1(n105), .B0(n168), .Y(n163) );
  NOR2X2 U123 ( .A(n40), .B(n153), .Y(n167) );
  AND2X4 U124 ( .A(n21), .B(n22), .Y(n80) );
  NAND2X2 U125 ( .A(n115), .B(n119), .Y(n113) );
  INVX2 U126 ( .A(n131), .Y(n119) );
  OAI2BB1X4 U127 ( .A0N(n12), .A1N(n150), .B0(n151), .Y(n110) );
  INVX4 U128 ( .A(n120), .Y(n115) );
  OAI21X4 U129 ( .A0(n46), .A1(n47), .B0(n48), .Y(n43) );
  NAND2BX4 U130 ( .AN(B[5]), .B(A[5]), .Y(n48) );
  CLKINVX1 U131 ( .A(n130), .Y(n89) );
  XOR2X4 U132 ( .A(n108), .B(n109), .Y(DIFF[15]) );
  OAI2BB1X4 U133 ( .A0N(n148), .A1N(A[10]), .B0(n149), .Y(n140) );
  NAND2BX4 U134 ( .AN(B[7]), .B(A[7]), .Y(n104) );
  INVX4 U135 ( .A(n67), .Y(n70) );
  AND2X2 U136 ( .A(n130), .B(n118), .Y(n19) );
  INVX4 U137 ( .A(n118), .Y(n92) );
  NAND2BX2 U138 ( .AN(B[13]), .B(A[13]), .Y(n118) );
  NAND2BX4 U139 ( .AN(B[2]), .B(A[2]), .Y(n64) );
  OAI21XL U140 ( .A0(A[7]), .A1(n156), .B0(n50), .Y(n186) );
  INVX4 U141 ( .A(B[7]), .Y(n156) );
  NAND2BX4 U142 ( .AN(A[4]), .B(B[4]), .Y(n50) );
  NAND2BX4 U143 ( .AN(A[3]), .B(B[3]), .Y(n60) );
  NAND2BX4 U144 ( .AN(B[9]), .B(A[9]), .Y(n32) );
  NAND2BX4 U145 ( .AN(A[11]), .B(B[11]), .Y(n137) );
  NAND3X4 U146 ( .A(n103), .B(n104), .C(n105), .Y(n30) );
  NAND2X2 U147 ( .A(n14), .B(n137), .Y(n97) );
  INVX4 U148 ( .A(n97), .Y(n146) );
  OAI21X1 U149 ( .A0(A[7]), .A1(n156), .B0(n50), .Y(n154) );
  NAND2X1 U150 ( .A(n49), .B(n50), .Y(n47) );
  INVX4 U151 ( .A(n44), .Y(n45) );
  INVXL U152 ( .A(A[6]), .Y(n16) );
  XOR2X2 U153 ( .A(n58), .B(n62), .Y(DIFF[2]) );
  NOR2X1 U154 ( .A(n59), .B(n63), .Y(n62) );
  NOR2X2 U155 ( .A(n70), .B(n66), .Y(n69) );
  OR2X2 U156 ( .A(n51), .B(n53), .Y(n17) );
  AND2X2 U157 ( .A(n57), .B(n60), .Y(n22) );
  NAND2X2 U158 ( .A(n48), .B(n54), .Y(n170) );
  XNOR2X2 U159 ( .A(n43), .B(n18), .Y(DIFF[6]) );
  INVX4 U160 ( .A(n26), .Y(n29) );
  NOR2X2 U161 ( .A(n152), .B(n153), .Y(n151) );
  INVXL U162 ( .A(A[10]), .Y(n141) );
  OAI21X2 U163 ( .A0(A[12]), .A1(n136), .B0(n137), .Y(n131) );
  NOR2X2 U164 ( .A(n76), .B(n77), .Y(n74) );
  NAND3BX4 U165 ( .AN(n80), .B(n61), .C(n106), .Y(n36) );
  NAND2XL U166 ( .A(n73), .B(n72), .Y(DIFF[0]) );
  NOR2X2 U167 ( .A(n121), .B(n122), .Y(n134) );
  NOR2X1 U168 ( .A(n95), .B(n96), .Y(n85) );
  NAND2X1 U169 ( .A(n32), .B(n37), .Y(n147) );
  NAND2XL U170 ( .A(n31), .B(n26), .Y(n177) );
  NAND2BX2 U171 ( .AN(n190), .B(n64), .Y(n189) );
  NAND2XL U172 ( .A(n100), .B(n90), .Y(n144) );
  NAND2X1 U173 ( .A(n88), .B(n101), .Y(n108) );
  INVXL U174 ( .A(n137), .Y(n160) );
  NAND2XL U175 ( .A(n31), .B(n32), .Y(n23) );
  INVX1 U176 ( .A(n32), .Y(n181) );
  OAI21X2 U177 ( .A0(n165), .A1(n32), .B0(n166), .Y(n164) );
  AOI21XL U178 ( .A0(n106), .A1(n61), .B0(n84), .Y(n102) );
  INVXL U179 ( .A(n57), .Y(n63) );
  AND2X2 U180 ( .A(n73), .B(n71), .Y(n21) );
  XOR2X2 U181 ( .A(n33), .B(n34), .Y(DIFF[8]) );
  NAND2XL U182 ( .A(n26), .B(n37), .Y(n33) );
  XOR2X2 U183 ( .A(n55), .B(n56), .Y(DIFF[3]) );
  NAND2X1 U184 ( .A(n60), .B(n61), .Y(n55) );
  XOR2X2 U185 ( .A(n68), .B(n69), .Y(DIFF[1]) );
  NAND3XL U186 ( .A(n170), .B(n173), .C(n42), .Y(n183) );
  INVX1 U187 ( .A(n88), .Y(n87) );
  NOR2X2 U188 ( .A(n186), .B(n155), .Y(n185) );
  NOR2X1 U189 ( .A(n154), .B(n155), .Y(n150) );
  XOR2X1 U190 ( .A(B[16]), .B(A[16]), .Y(n75) );
  NAND2BX2 U191 ( .AN(A[5]), .B(B[5]), .Y(n49) );
  NAND2BX1 U192 ( .AN(B[10]), .B(A[10]), .Y(n166) );
  INVXL U193 ( .A(B[10]), .Y(n148) );
  OAI21XL U194 ( .A0(n102), .A1(n1), .B0(n81), .Y(n98) );
  NAND2BX2 U195 ( .AN(B[12]), .B(A[12]), .Y(n90) );
  NAND2BXL U196 ( .AN(A[1]), .B(B[1]), .Y(n190) );
  XOR2X4 U197 ( .A(n124), .B(n125), .Y(DIFF[14]) );
  AOI21X4 U198 ( .A0(n110), .A1(n126), .B0(n127), .Y(n125) );
  XOR2X4 U199 ( .A(n144), .B(n145), .Y(DIFF[12]) );
  AOI21X4 U200 ( .A0(n81), .A1(n110), .B0(n146), .Y(n145) );
  CLKINVX3 U201 ( .A(n157), .Y(n81) );
  XOR2X4 U202 ( .A(n158), .B(n159), .Y(DIFF[11]) );
  NOR2BX4 U203 ( .AN(n149), .B(n160), .Y(n159) );
  NAND3X4 U204 ( .A(n170), .B(n42), .C(n171), .Y(n105) );
  XOR2X4 U205 ( .A(n175), .B(n176), .Y(DIFF[10]) );
  NOR2BX4 U206 ( .AN(n166), .B(n165), .Y(n176) );
  NAND2BX4 U207 ( .AN(A[8]), .B(B[8]), .Y(n26) );
  NAND2BX4 U208 ( .AN(A[9]), .B(B[9]), .Y(n31) );
  NAND2BX4 U209 ( .AN(A[2]), .B(B[2]), .Y(n57) );
endmodule


module butterfly ( calc_in, rotation, calc_out );
  input [135:0] calc_in;
  input [2:0] rotation;
  output [135:0] calc_out;
  wire   n109, n110, n111, n112, N9, N42, N43, n7, n9, N306, N305, N304, N303,
         N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292,
         N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281,
         N280, N279, N278, N277, N276, N275, N274, N273, N238, N237, N236,
         N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225,
         N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214,
         N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203,
         N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192,
         N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181,
         N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N136,
         N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125,
         N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114,
         N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103,
         N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330,
         N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319,
         N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308,
         N307, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263,
         N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252,
         N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241,
         N240, N239, N170, N169, N168, N167, N166, N165, N164, N163, N162,
         N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151,
         N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140,
         N139, N138, N137, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90,
         N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76,
         N75, N74, N73, N72, N71, N70, N69, N102, N101, N100, n8, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n54, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84;
  wire   [16:0] temp_2_1_real;
  wire   [16:0] temp_2_2_real;
  wire   [16:0] temp_2_1_imag;
  wire   [16:0] temp_2_2_imag;
  wire   [16:0] temp_3_1_real;
  wire   [16:0] temp_3_2_real;
  wire   [16:0] temp_3_1_imag;
  wire   [16:0] temp_3_2_imag;
  wire   [16:0] temp_4_1_real;
  wire   [16:0] temp_4_2_real;
  wire   [16:0] temp_4_1_imag;
  wire   [16:0] temp_4_2_imag;
  wire   [16:0] temp_1_real;
  wire   [16:0] temp_1_imag;
  wire   [16:0] temp_2_real;
  wire   [16:0] temp_2_imag;
  wire   [16:0] temp_3_real;
  wire   [16:0] temp_3_imag;

  multi16_0 multiBRR ( .in_17bit({n79, calc_in[66:51]}), .in_8bit({1'b0, n72, 
        n7, 1'b1, n13, n63, n72, n76}), .out(temp_2_1_real) );
  multi16_11 multiBII ( .in_17bit(calc_in[50:34]), .in_8bit({n66, n68, n65, 
        1'b0, n70, n78, n61, n67}), .out(temp_2_2_real) );
  multi16_10 multiBRI ( .in_17bit({n79, calc_in[66:51]}), .in_8bit({n66, n68, 
        n65, 1'b0, n70, n78, n61, n67}), .out(temp_2_1_imag) );
  multi16_9 multiBIR ( .in_17bit(calc_in[50:34]), .in_8bit({1'b0, n72, n7, 
        1'b1, n14, n63, n72, n77}), .out(temp_2_2_imag) );
  multi16_8 multiCRR ( .in_17bit({n80, calc_in[100:85]}), .in_8bit({n73, n63, 
        n77, n63, n63, n75, n7, N42}), .out(temp_3_1_real) );
  multi16_7 multiCII ( .in_17bit(calc_in[84:68]), .in_8bit({n58, 1'b0, n70, 
        1'b0, 1'b0, n70, n70, n65}), .out(temp_3_2_real) );
  multi16_6 multiCRI ( .in_17bit({n80, calc_in[100:85]}), .in_8bit({n66, 1'b0, 
        n70, 1'b0, 1'b0, n70, n70, n65}), .out(temp_3_1_imag) );
  multi16_5 multiCIR ( .in_17bit(calc_in[84:68]), .in_8bit({n73, n63, n77, n63, 
        n63, n76, n7, N42}), .out(temp_3_2_imag) );
  multi16_4 multiDRR ( .in_17bit({n81, calc_in[134:119]}), .in_8bit({n9, N42, 
        n72, n63, n76, n14, n69, n63}), .out(temp_4_1_real) );
  multi16_3 multiDII ( .in_17bit(calc_in[118:102]), .in_8bit({n78, 1'b0, n64, 
        n74, n67, n65, n78, n73}), .out(temp_4_2_real) );
  multi16_2 multiDRI ( .in_17bit({n81, calc_in[134:119]}), .in_8bit({n78, 1'b0, 
        n64, n74, n67, n65, n78, n73}), .out(temp_4_1_imag) );
  multi16_1 multiDIR ( .in_17bit(calc_in[118:102]), .in_8bit({n9, N42, n72, 
        n63, n75, n13, n69, n63}), .out(temp_4_2_imag) );
  butterfly_DW01_sub_14 sub_0_root_sub_0_root_sub_300_2 ( .A({N306, N305, N304, 
        N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, 
        N291, N290}), .B({N289, N288, N287, N286, N285, N284, N283, N282, N281, 
        N280, N279, N278, N277, N276, N275, N274, N273}), .DIFF(
        calc_out[67:51]) );
  butterfly_DW01_add_21 add_0_root_add_0_root_add_292_3 ( .A({N102, N101, N100, 
        N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86}), 
        .B({N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, 
        N72, N71, N70, N69}), .SUM({calc_out[33:31], n112, calc_out[29:17]})
         );
  butterfly_DW01_sub_36 sub_2_root_sub_0_root_sub_299_2 ( .A(calc_in[16:0]), 
        .B({temp_3_real[16:15], n10, n15, n48, n51, temp_3_real[10:2], n21, 
        temp_3_real[0]}), .DIFF({N272, N271, N270, N269, N268, N267, N266, 
        N265, N264, N263, N262, N261, N260, N259, N258, N257, N256}) );
  butterfly_DW01_add_43 add_2_root_sub_0_root_sub_300_2 ( .A(calc_in[33:17]), 
        .B({temp_1_imag[16:6], n47, temp_1_imag[4], n57, temp_1_imag[2:0]}), 
        .SUM({N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, 
        N295, N294, N293, N292, N291, N290}) );
  butterfly_DW01_sub_38 sub_1_root_sub_0_root_sub_299_2 ( .A({temp_1_real[16], 
        n27, temp_1_real[14:12], n42, n50, n16, n45, temp_1_real[7:4], n26, 
        n38, n18, temp_1_real[0]}), .B({temp_2_imag[16:15], n28, 
        temp_2_imag[13:7], n29, temp_2_imag[5:0]}), .DIFF({N255, N254, N253, 
        N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, 
        N240, N239}) );
  butterfly_DW01_add_52 add_0_root_sub_0_root_add_301 ( .A({N340, N339, N338, 
        N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, 
        N325, N324}), .B({N323, N322, N321, N320, N319, N318, N317, N316, N315, 
        N314, N313, N312, N311, N310, N309, N308, N307}), .SUM(calc_out[50:34]) );
  butterfly_DW01_add_64 add_0_root_sub_0_root_sub_296_2 ( .A({N204, N203, N202, 
        N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, 
        N189, N188}), .B({N187, N186, N185, N184, N183, N182, N181, N180, N179, 
        N178, N177, N176, N175, N174, N173, N172, N171}), .SUM(calc_out[84:68]) );
  butterfly_DW01_add_69 add_2_root_add_0_root_add_292_3 ( .A(calc_in[33:17]), 
        .B({temp_2_real[16:14], n19, n37, temp_2_real[11:5], n24, n34, 
        temp_2_real[2:0]}), .SUM({N102, N101, N100, N99, N98, N97, N96, N95, 
        N94, N93, N92, N91, N90, N89, N88, N87, N86}) );
  butterfly_DW01_sub_68 sub_2_root_sub_0_root_add_301 ( .A(calc_in[16:0]), .B(
        {temp_1_real[16], n27, temp_1_real[14:12], n42, n50, n16, 
        temp_1_real[8:4], n26, n38, n18, temp_1_real[0]}), .DIFF({N340, N339, 
        N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, 
        N326, N325, N324}) );
  butterfly_DW01_add_94 add_1_root_sub_0_root_sub_300_2 ( .A({
        temp_3_imag[16:11], n20, temp_3_imag[9:8], n71, temp_3_imag[6], n49, 
        n22, n44, n36, temp_3_imag[1:0]}), .B({temp_2_real[16:14], n19, n37, 
        temp_2_real[11:5], n24, n34, temp_2_real[2:0]}), .SUM({N289, N288, 
        N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, 
        N275, N274, N273}) );
  butterfly_DW01_sub_69 sub_0_root_sub_0_root_sub_295_2 ( .A({N170, N169, N168, 
        N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, 
        N155, N154}), .B({N153, N152, N151, N150, N149, n46, N147, N146, N145, 
        N144, N143, N142, N141, N140, N139, N138, N137}), .DIFF({
        calc_out[101:93], n111, calc_out[91:85]}) );
  butterfly_DW01_sub_82 sub_2_root_sub_0_root_sub_296_2 ( .A(calc_in[16:0]), 
        .B({temp_1_imag[16:6], n47, temp_1_imag[4], n57, temp_1_imag[2:0]}), 
        .DIFF({N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, 
        N194, N193, N192, N191, N190, N189, N188}) );
  butterfly_DW01_add_88 add_0_root_add_0_root_add_293_3 ( .A({N136, N135, N134, 
        N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, n41, 
        N121, N120}), .B({N119, N118, N117, N116, N115, N114, N113, N112, N111, 
        N110, N109, N108, N107, N106, N105, N104, N103}), .SUM(calc_out[16:0])
         );
  butterfly_DW01_add_103 add_2_root_sub_0_root_sub_295_2 ( .A(calc_in[33:17]), 
        .B({temp_2_real[16:14], n19, n37, temp_2_real[11:5], n24, n34, 
        temp_2_real[2:0]}), .SUM({N170, N169, N168, N167, N166, N165, N164, 
        N163, N162, N161, N160, N159, N158, N157, N156, N155, N154}) );
  butterfly_DW01_sub_79 sub_275 ( .A(temp_2_1_real), .B({temp_2_2_real[16:2], 
        n39, temp_2_2_real[0]}), .DIFF(temp_1_real) );
  butterfly_DW01_add_114 add_282 ( .A(temp_4_1_imag), .B({temp_4_2_imag[16:2], 
        n40, temp_4_2_imag[0]}), .SUM(temp_3_imag) );
  butterfly_DW01_add_108 add_0_root_sub_0_root_sub_299_2 ( .A({N272, N271, 
        N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, 
        N258, N257, N256}), .B({N255, N254, N253, N252, N251, N250, N249, N248, 
        N247, N246, N245, N244, N243, N242, N241, N240, N239}), .SUM({
        calc_out[118:114], n110, calc_out[112:102]}) );
  butterfly_DW01_add_112 add_1_root_sub_0_root_sub_295_2 ( .A({temp_1_real[16], 
        n27, temp_1_real[14:12], n42, n50, n16, n45, temp_1_real[7:4], n26, 
        n38, n18, temp_1_real[0]}), .B({temp_3_real[16:15], n10, n31, n48, n51, 
        temp_3_real[10:2], n21, temp_3_real[0]}), .SUM({N153, N152, N151, N150, 
        N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, 
        N137}) );
  butterfly_DW01_add_113 add_1_root_add_0_root_add_292_3 ( .A({temp_1_real[16], 
        n27, temp_1_real[14:12], n42, n50, n16, n45, temp_1_real[7:3], n38, 
        n18, temp_1_real[0]}), .B({temp_3_real[16:15], n10, n31, n48, n51, 
        temp_3_real[10:2], n21, temp_3_real[0]}), .SUM({N85, N84, N83, N82, 
        N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69}) );
  butterfly_DW01_sub_95 sub_1_root_sub_0_root_add_298 ( .A({temp_3_imag[16:11], 
        n20, temp_3_imag[9:8], n71, temp_3_imag[6], n49, n22, n44, 
        temp_3_imag[2:0]}), .B({temp_2_real[16:14], n19, n37, 
        temp_2_real[11:5], n24, n34, temp_2_real[2:0]}), .DIFF({N221, N220, 
        N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, 
        N207, N206, N205}) );
  butterfly_DW01_add_123 add_2_root_add_0_root_add_293_3 ( .A(calc_in[16:0]), 
        .B({temp_2_imag[16:15], n28, temp_2_imag[13:7], n29, temp_2_imag[5:0]}), .SUM({N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, 
        N124, N123, N122, N121, N120}) );
  butterfly_DW01_sub_100 sub_1_root_sub_0_root_sub_296_2 ( .A({
        temp_2_imag[16:15], n28, temp_2_imag[13:7], n29, temp_2_imag[5:0]}), 
        .B({n8, temp_3_imag[15:11], n20, temp_3_imag[9:8], n71, temp_3_imag[6], 
        n49, n22, n44, n36, temp_3_imag[1:0]}), .DIFF({N187, N186, N185, N184, 
        N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, 
        N171}) );
  butterfly_DW01_sub_98 sub_1_root_sub_0_root_add_301 ( .A({temp_3_real[16:15], 
        n10, n15, n48, n51, temp_3_real[10:2], n21, temp_3_real[0]}), .B({
        temp_2_imag[16:15], n28, temp_2_imag[13:7], n29, temp_2_imag[5:0]}), 
        .DIFF({N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, 
        N313, N312, N311, N310, N309, N308, N307}) );
  butterfly_DW01_add_140 add_276 ( .A(temp_2_1_imag), .B({temp_2_2_imag[16:9], 
        n43, temp_2_2_imag[7:0]}), .SUM(temp_1_imag) );
  butterfly_DW01_sub_112 sub_278 ( .A(temp_3_1_real), .B(temp_3_2_real), 
        .DIFF(temp_2_real) );
  butterfly_DW01_sub_114 sub_281 ( .A({temp_4_1_real[16:3], n35, 
        temp_4_1_real[1:0]}), .B(temp_4_2_real), .DIFF(temp_3_real) );
  butterfly_DW01_add_129 add_0_root_sub_0_root_add_298 ( .A({N238, N237, N236, 
        N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, 
        N223, N222}), .B({N221, N220, N219, N218, N217, N216, N215, N214, N213, 
        N212, N211, N210, n25, N208, N207, N206, N205}), .SUM({
        calc_out[135:132], n109, calc_out[130:119]}) );
  butterfly_DW01_add_147 add_279 ( .A(temp_3_1_imag), .B(temp_3_2_imag), .SUM(
        temp_2_imag) );
  butterfly_DW01_add_145 add_1_root_add_0_root_add_293_3 ( .A({
        temp_1_imag[16:6], n47, temp_1_imag[4], n57, temp_1_imag[2:0]}), .B({
        temp_3_imag[16:11], n20, temp_3_imag[9:8], n71, temp_3_imag[6], n49, 
        n22, n44, n36, temp_3_imag[1:0]}), .SUM({N119, N118, N117, N116, N115, 
        N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103}) );
  butterfly_DW01_sub_120 sub_2_root_sub_0_root_add_298 ( .A(calc_in[33:17]), 
        .B({temp_1_imag[16:6], n47, temp_1_imag[4], n57, temp_1_imag[2:0]}), 
        .DIFF({N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, 
        N228, N227, N226, N225, N224, N223, N222}) );
  BUFX3 U9 ( .A(temp_3_imag[16]), .Y(n8) );
  BUFX12 U10 ( .A(temp_3_real[13]), .Y(n15) );
  BUFX20 U11 ( .A(temp_3_imag[2]), .Y(n36) );
  BUFX16 U12 ( .A(n112), .Y(calc_out[30]) );
  INVX8 U13 ( .A(n30), .Y(n31) );
  BUFX16 U14 ( .A(calc_in[101]), .Y(n80) );
  NAND2X4 U15 ( .A(n62), .B(rotation[2]), .Y(n83) );
  BUFX8 U16 ( .A(N209), .Y(n25) );
  BUFX16 U17 ( .A(temp_4_1_real[2]), .Y(n35) );
  CLKINVX3 U18 ( .A(n83), .Y(n9) );
  BUFX16 U19 ( .A(n58), .Y(n66) );
  CLKINVX1 U20 ( .A(n58), .Y(N42) );
  INVX20 U21 ( .A(N43), .Y(n73) );
  BUFX12 U22 ( .A(rotation[0]), .Y(n56) );
  BUFX12 U23 ( .A(rotation[1]), .Y(n62) );
  BUFX12 U24 ( .A(temp_2_2_real[1]), .Y(n39) );
  CLKINVX3 U25 ( .A(temp_3_real[13]), .Y(n30) );
  BUFX12 U26 ( .A(N148), .Y(n46) );
  BUFX12 U27 ( .A(temp_3_real[14]), .Y(n10) );
  AND2X1 U28 ( .A(n56), .B(rotation[2]), .Y(n11) );
  BUFX16 U29 ( .A(calc_in[135]), .Y(n81) );
  NAND2X2 U30 ( .A(n60), .B(rotation[2]), .Y(N9) );
  OR2XL U31 ( .A(n13), .B(n62), .Y(n12) );
  INVXL U32 ( .A(N43), .Y(n74) );
  INVXL U33 ( .A(n11), .Y(n13) );
  INVXL U34 ( .A(n11), .Y(n14) );
  BUFX20 U35 ( .A(temp_1_real[2]), .Y(n38) );
  BUFX20 U36 ( .A(temp_3_imag[3]), .Y(n44) );
  BUFX20 U37 ( .A(temp_1_imag[3]), .Y(n57) );
  BUFX20 U38 ( .A(temp_2_imag[14]), .Y(n28) );
  BUFX20 U39 ( .A(temp_1_imag[5]), .Y(n47) );
  BUFX20 U40 ( .A(temp_2_real[13]), .Y(n19) );
  BUFX20 U41 ( .A(temp_1_real[9]), .Y(n16) );
  BUFX16 U42 ( .A(temp_1_real[8]), .Y(n45) );
  INVX4 U43 ( .A(temp_1_real[1]), .Y(n17) );
  INVX8 U44 ( .A(n17), .Y(n18) );
  BUFX20 U45 ( .A(temp_3_real[12]), .Y(n48) );
  BUFX20 U46 ( .A(temp_2_real[4]), .Y(n24) );
  INVX2 U47 ( .A(rotation[2]), .Y(n59) );
  BUFX20 U48 ( .A(temp_3_imag[10]), .Y(n20) );
  BUFX12 U49 ( .A(temp_3_real[1]), .Y(n21) );
  BUFX20 U50 ( .A(temp_2_real[12]), .Y(n37) );
  BUFX20 U51 ( .A(temp_3_imag[5]), .Y(n49) );
  BUFX20 U52 ( .A(temp_1_real[11]), .Y(n42) );
  BUFX20 U53 ( .A(temp_3_imag[4]), .Y(n22) );
  BUFX12 U54 ( .A(temp_2_2_imag[8]), .Y(n43) );
  BUFX20 U55 ( .A(temp_1_real[10]), .Y(n50) );
  BUFX20 U56 ( .A(temp_1_real[3]), .Y(n26) );
  BUFX12 U57 ( .A(temp_1_real[15]), .Y(n27) );
  BUFX20 U58 ( .A(temp_2_imag[6]), .Y(n29) );
  CLKINVX8 U59 ( .A(n111), .Y(n32) );
  INVX8 U60 ( .A(n32), .Y(calc_out[92]) );
  BUFX12 U61 ( .A(temp_2_real[3]), .Y(n34) );
  BUFX8 U62 ( .A(temp_4_2_imag[1]), .Y(n40) );
  BUFX8 U63 ( .A(N122), .Y(n41) );
  BUFX20 U64 ( .A(temp_3_real[11]), .Y(n51) );
  CLKINVX8 U65 ( .A(n110), .Y(n52) );
  INVX8 U66 ( .A(n52), .Y(calc_out[113]) );
  CLKINVX8 U67 ( .A(n109), .Y(n54) );
  INVX8 U68 ( .A(n54), .Y(calc_out[131]) );
  BUFX20 U69 ( .A(calc_in[67]), .Y(n79) );
  AOI2BB1X4 U70 ( .A0N(n56), .A1N(n62), .B0(n59), .Y(n58) );
  NAND2BX4 U71 ( .AN(n83), .B(n56), .Y(N43) );
  INVX8 U72 ( .A(N9), .Y(n78) );
  XOR2X4 U73 ( .A(n56), .B(n62), .Y(n60) );
  INVXL U74 ( .A(n74), .Y(n72) );
  INVX1 U75 ( .A(n68), .Y(n69) );
  CLKBUFXL U76 ( .A(n66), .Y(n61) );
  INVX1 U77 ( .A(n12), .Y(n68) );
  CLKINVX3 U78 ( .A(n64), .Y(n63) );
  INVXL U79 ( .A(n83), .Y(n64) );
  INVX1 U80 ( .A(n12), .Y(n67) );
  INVX1 U81 ( .A(n78), .Y(n75) );
  INVX1 U82 ( .A(n78), .Y(n76) );
  INVX1 U83 ( .A(n78), .Y(n77) );
  BUFX3 U84 ( .A(n11), .Y(n70) );
  BUFX3 U85 ( .A(n84), .Y(n65) );
  INVX1 U86 ( .A(n7), .Y(n84) );
  NAND2X2 U87 ( .A(n64), .B(n82), .Y(n7) );
  INVXL U88 ( .A(n56), .Y(n82) );
  BUFX20 U89 ( .A(temp_3_imag[7]), .Y(n71) );
endmodule


module reg1 ( clk, rst_n, data_in_2, reg_datain_flag, data_out_2 );
  input [135:0] data_in_2;
  output [135:0] data_out_2;
  input clk, rst_n, reg_datain_flag;
  wire   reg_flag_mux, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62,
         N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76,
         N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90,
         N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, N124, N125,
         N126, N127, N128, N129, N130, N131, N132, N133, N134, N135, N136,
         N137, N138, N139, N140, N141, N142, N143, N144, N145, N146, N147,
         N148, N149, N150, N151, N152, N153, N154, N155, N156, N157, N158,
         N159, N160, N161, N162, N163, N164, N165, N166, N167, N168, N169,
         N170, N171, N172, N173, N174, N175, N176, N177, N178, N179, N180,
         N181, N182, N183, N184, N185, N186, N187, n150, n151, n152, n153,
         n165, n167, n168, n169, n170, n184, n185, n186, n195, n201, n203,
         n204, n286, n287, n288, n289, n301, n303, n304, n305, n306, n320,
         n321, n322, n331, n337, n339, n340, n422, n423, n424, n425, n437,
         n439, n440, n441, n442, n456, n457, n458, n467, n473, n475, n476,
         n524, n525, n526, n535, n541, n543, n544, n558, n559, n560, n561,
         n573, n575, n576, n577, n578, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n961, n962, n963, n964, n965, n966, n968, n969, n971,
         n973, n974, n975, n976, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
         n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
         n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
         n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
         n1116, n2, n6, n7, n30, n58, n59, n78, n114, n115, n603, n604, n605,
         n606, n607, n608, n609, n610, n612, n614, n616, n618, n620, n622,
         n624, n626, n628, n630, n632, n634, n636, n638, n640, n642, n644,
         n646, n648, n650, n652, n654, n656, n658, n660, n662, n664, n666,
         n668, n670, n672, n674, n676, n678, n680, n682, n684, n958, n960,
         n970, n977, n1118, n1120, n1122, n1124, n1126, n1128, n1130, n1132,
         n1134, n1136, n1138, n1140, n1142, n1144, n1146, n1148, n1150, n1152,
         n1154, n1156, n1158, n1160, n1162, n1164, n1166, n1168, n1170, n1172,
         n1174, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
         n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
         n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
         n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
         n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
         n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
         n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
         n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
         n1327, n1328, n1329;
  wire   [1:0] counter1;
  wire   [33:0] R0;
  wire   [33:0] R1;
  wire   [33:0] R4;
  wire   [33:0] R5;
  wire   [33:0] R8;
  wire   [33:0] R9;
  wire   [33:0] R12;
  wire   [33:0] R13;
  wire   [1:0] counter2;

  CLKINVX4 U302 ( .A(rst_n), .Y(n961) );
  EDFFXL R10_reg_31_ ( .D(data_in_2[99]), .E(n1258), .CK(clk), .QN(n722) );
  EDFFXL R14_reg_31_ ( .D(data_in_2[99]), .E(n1283), .CK(clk), .QN(n756) );
  EDFFXL R2_reg_31_ ( .D(data_in_2[99]), .E(n115), .CK(clk), .QN(n824) );
  EDFFXL R6_reg_31_ ( .D(data_in_2[99]), .E(n1292), .CK(clk), .QN(n892) );
  EDFFXL R13_reg_13_ ( .D(data_in_2[47]), .E(n1286), .CK(clk), .Q(R13[13]) );
  EDFFXL R9_reg_13_ ( .D(data_in_2[47]), .E(n1254), .CK(clk), .Q(R9[13]) );
  EDFFXL R1_reg_13_ ( .D(data_in_2[47]), .E(n1266), .CK(clk), .Q(R1[13]) );
  EDFFXL R5_reg_13_ ( .D(data_in_2[47]), .E(n1291), .CK(clk), .Q(R5[13]) );
  EDFFXL R4_reg_16_ ( .D(data_in_2[16]), .E(n1289), .CK(clk), .Q(R4[16]) );
  EDFFXL R0_reg_16_ ( .D(data_in_2[16]), .E(n1264), .CK(clk), .Q(R0[16]) );
  EDFFXL R12_reg_16_ ( .D(data_in_2[16]), .E(n1284), .CK(clk), .Q(R12[16]) );
  EDFFXL R8_reg_16_ ( .D(data_in_2[16]), .E(n1262), .CK(clk), .Q(R8[16]) );
  DFFXL R14_reg_14_ ( .D(n1236), .CK(clk), .Q(n457), .QN(n773) );
  DFFXL R10_reg_14_ ( .D(n1235), .CK(clk), .Q(n525), .QN(n739) );
  DFFXL R6_reg_14_ ( .D(n1234), .CK(clk), .Q(n185), .QN(n909) );
  DFFXL R2_reg_14_ ( .D(n1233), .CK(clk), .Q(n321), .QN(n841) );
  MX2X1 R15_reg_28__U3 ( .A(n437), .B(data_in_2[130]), .S0(n1280), .Y(n1232)
         );
  DFFXL R15_reg_28_ ( .D(n1232), .CK(clk), .Q(n437), .QN(n793) );
  MX2X1 R11_reg_28__U3 ( .A(n573), .B(data_in_2[130]), .S0(n1261), .Y(n1231)
         );
  DFFXL R11_reg_28_ ( .D(n1231), .CK(clk), .Q(n573), .QN(n691) );
  MX2X1 R7_reg_28__U3 ( .A(n165), .B(data_in_2[130]), .S0(n1294), .Y(n1230) );
  DFFXL R7_reg_28_ ( .D(n1230), .CK(clk), .Q(n165), .QN(n929) );
  MX2X1 R3_reg_28__U3 ( .A(n301), .B(data_in_2[130]), .S0(n1267), .Y(n1229) );
  DFFXL R3_reg_28_ ( .D(n1229), .CK(clk), .Q(n301), .QN(n861) );
  MX2X1 R15_reg_31__U3 ( .A(n440), .B(data_in_2[133]), .S0(n1280), .Y(n1228)
         );
  DFFXL R15_reg_31_ ( .D(n1228), .CK(clk), .Q(n440), .QN(n790) );
  MX2X1 R11_reg_31__U3 ( .A(n576), .B(data_in_2[133]), .S0(n1261), .Y(n1227)
         );
  DFFXL R11_reg_31_ ( .D(n1227), .CK(clk), .Q(n576), .QN(n688) );
  MX2X1 R7_reg_31__U3 ( .A(n168), .B(data_in_2[133]), .S0(n1294), .Y(n1226) );
  DFFXL R7_reg_31_ ( .D(n1226), .CK(clk), .Q(n168), .QN(n926) );
  MX2X1 R3_reg_31__U3 ( .A(n304), .B(data_in_2[133]), .S0(n1267), .Y(n1225) );
  DFFXL R3_reg_31_ ( .D(n1225), .CK(clk), .Q(n304), .QN(n858) );
  MX2X1 R14_reg_15__U3 ( .A(n458), .B(data_in_2[83]), .S0(n1282), .Y(n1224) );
  DFFXL R14_reg_15_ ( .D(n1224), .CK(clk), .Q(n458), .QN(n772) );
  MX2X1 R10_reg_15__U3 ( .A(n526), .B(data_in_2[83]), .S0(n1257), .Y(n1223) );
  DFFXL R10_reg_15_ ( .D(n1223), .CK(clk), .Q(n526), .QN(n738) );
  MX2X1 R6_reg_15__U3 ( .A(n186), .B(data_in_2[83]), .S0(n1293), .Y(n1222) );
  DFFXL R6_reg_15_ ( .D(n1222), .CK(clk), .Q(n186), .QN(n908) );
  MX2X1 R2_reg_15__U3 ( .A(n322), .B(data_in_2[83]), .S0(n1267), .Y(n1221) );
  DFFXL R2_reg_15_ ( .D(n1221), .CK(clk), .Q(n322), .QN(n840) );
  MX2X1 R14_reg_16__U3 ( .A(n1250), .B(data_in_2[84]), .S0(n1282), .Y(n1220)
         );
  DFFXL R14_reg_16_ ( .D(n1220), .CK(clk), .Q(n1250), .QN(n771) );
  MX2X1 R10_reg_16__U3 ( .A(n1249), .B(data_in_2[84]), .S0(n1257), .Y(n1219)
         );
  DFFXL R10_reg_16_ ( .D(n1219), .CK(clk), .Q(n1249), .QN(n737) );
  MX2X1 R6_reg_16__U3 ( .A(n1252), .B(data_in_2[84]), .S0(n1293), .Y(n1218) );
  DFFXL R6_reg_16_ ( .D(n1218), .CK(clk), .Q(n1252), .QN(n907) );
  MX2X1 R2_reg_16__U3 ( .A(n1251), .B(data_in_2[84]), .S0(n115), .Y(n1217) );
  DFFXL R2_reg_16_ ( .D(n1217), .CK(clk), .Q(n1251), .QN(n839) );
  DFFXL R15_reg_32_ ( .D(n1216), .CK(clk), .Q(n441), .QN(n789) );
  MX2X1 R11_reg_32__U3 ( .A(n577), .B(data_in_2[134]), .S0(n1261), .Y(n1215)
         );
  DFFXL R11_reg_32_ ( .D(n1215), .CK(clk), .Q(n577), .QN(n687) );
  MX2X1 R7_reg_32__U3 ( .A(n169), .B(data_in_2[134]), .S0(n1293), .Y(n1214) );
  DFFXL R7_reg_32_ ( .D(n1214), .CK(clk), .Q(n169), .QN(n925) );
  MX2X1 R3_reg_32__U3 ( .A(n305), .B(data_in_2[134]), .S0(n1267), .Y(n1213) );
  DFFXL R3_reg_32_ ( .D(n1213), .CK(clk), .Q(n305), .QN(n857) );
  DFFXL R15_reg_30_ ( .D(n1212), .CK(clk), .Q(n439), .QN(n791) );
  DFFXL R11_reg_30_ ( .D(n1211), .CK(clk), .Q(n575), .QN(n689) );
  DFFXL R7_reg_30_ ( .D(n1210), .CK(clk), .Q(n167), .QN(n927) );
  DFFXL R3_reg_30_ ( .D(n1209), .CK(clk), .Q(n303), .QN(n859) );
  MX2X1 R15_reg_16__U3 ( .A(n425), .B(data_in_2[118]), .S0(n1279), .Y(n1208)
         );
  DFFXL R15_reg_16_ ( .D(n1208), .CK(clk), .Q(n425), .QN(n805) );
  MX2X1 R11_reg_16__U3 ( .A(n561), .B(data_in_2[118]), .S0(n1260), .Y(n1207)
         );
  DFFXL R11_reg_16_ ( .D(n1207), .CK(clk), .Q(n561), .QN(n703) );
  MX2X1 R7_reg_16__U3 ( .A(n153), .B(data_in_2[118]), .S0(n1294), .Y(n1206) );
  DFFXL R7_reg_16_ ( .D(n1206), .CK(clk), .Q(n153), .QN(n941) );
  MX2X1 R3_reg_16__U3 ( .A(n289), .B(data_in_2[118]), .S0(n1268), .Y(n1205) );
  DFFXL R3_reg_16_ ( .D(n1205), .CK(clk), .Q(n289), .QN(n873) );
  MX2X1 R15_reg_13__U3 ( .A(n422), .B(data_in_2[115]), .S0(n1279), .Y(n1204)
         );
  DFFXL R15_reg_13_ ( .D(n1204), .CK(clk), .Q(n422), .QN(n808) );
  MX2X1 R11_reg_13__U3 ( .A(n558), .B(data_in_2[115]), .S0(n1259), .Y(n1203)
         );
  DFFXL R11_reg_13_ ( .D(n1203), .CK(clk), .Q(n558), .QN(n706) );
  MX2X1 R7_reg_13__U3 ( .A(n150), .B(data_in_2[115]), .S0(n1294), .Y(n1202) );
  DFFXL R7_reg_13_ ( .D(n1202), .CK(clk), .Q(n150), .QN(n944) );
  MX2X1 R3_reg_13__U3 ( .A(n286), .B(data_in_2[115]), .S0(n1268), .Y(n1201) );
  DFFXL R3_reg_13_ ( .D(n1201), .CK(clk), .Q(n286), .QN(n876) );
  MX2X1 R14_reg_24__U3 ( .A(n467), .B(data_in_2[92]), .S0(n1282), .Y(n1200) );
  DFFXL R14_reg_24_ ( .D(n1200), .CK(clk), .Q(n467), .QN(n763) );
  MX2X1 R10_reg_24__U3 ( .A(n535), .B(data_in_2[92]), .S0(n1257), .Y(n1199) );
  DFFXL R10_reg_24_ ( .D(n1199), .CK(clk), .Q(n535), .QN(n729) );
  MX2X1 R6_reg_24__U3 ( .A(n195), .B(data_in_2[92]), .S0(n1292), .Y(n1198) );
  DFFXL R6_reg_24_ ( .D(n1198), .CK(clk), .Q(n195), .QN(n899) );
  MX2X1 R2_reg_24__U3 ( .A(n331), .B(data_in_2[92]), .S0(n1266), .Y(n1197) );
  DFFXL R2_reg_24_ ( .D(n1197), .CK(clk), .Q(n331), .QN(n831) );
  MX2X1 R14_reg_32__U3 ( .A(n475), .B(data_in_2[100]), .S0(n1283), .Y(n1196)
         );
  DFFXL R14_reg_32_ ( .D(n1196), .CK(clk), .Q(n475), .QN(n755) );
  MX2X1 R10_reg_32__U3 ( .A(n543), .B(data_in_2[100]), .S0(n1258), .Y(n1195)
         );
  DFFXL R10_reg_32_ ( .D(n1195), .CK(clk), .Q(n543), .QN(n721) );
  MX2X1 R6_reg_32__U3 ( .A(n203), .B(data_in_2[100]), .S0(n1292), .Y(n1194) );
  DFFXL R6_reg_32_ ( .D(n1194), .CK(clk), .Q(n203), .QN(n891) );
  MX2X1 R2_reg_32__U3 ( .A(n339), .B(data_in_2[100]), .S0(n115), .Y(n1193) );
  DFFXL R2_reg_32_ ( .D(n1193), .CK(clk), .Q(n339), .QN(n823) );
  MX2X1 R14_reg_30__U3 ( .A(n473), .B(data_in_2[98]), .S0(n1283), .Y(n1192) );
  DFFXL R14_reg_30_ ( .D(n1192), .CK(clk), .Q(n473), .QN(n757) );
  MX2X1 R10_reg_30__U3 ( .A(n541), .B(data_in_2[98]), .S0(n1258), .Y(n1191) );
  DFFXL R10_reg_30_ ( .D(n1191), .CK(clk), .Q(n541), .QN(n723) );
  MX2X1 R6_reg_30__U3 ( .A(n201), .B(data_in_2[98]), .S0(n1292), .Y(n1190) );
  DFFXL R6_reg_30_ ( .D(n1190), .CK(clk), .Q(n201), .QN(n893) );
  MX2X1 R2_reg_30__U3 ( .A(n337), .B(data_in_2[98]), .S0(n1267), .Y(n1189) );
  DFFXL R2_reg_30_ ( .D(n1189), .CK(clk), .Q(n337), .QN(n825) );
  MX2X1 R15_reg_33__U3 ( .A(n442), .B(data_in_2[135]), .S0(n1280), .Y(n1188)
         );
  DFFXL R15_reg_33_ ( .D(n1188), .CK(clk), .Q(n442), .QN(n788) );
  MX2X1 R11_reg_33__U3 ( .A(n578), .B(data_in_2[135]), .S0(n1261), .Y(n1187)
         );
  DFFXL R11_reg_33_ ( .D(n1187), .CK(clk), .Q(n578), .QN(n686) );
  MX2X1 R7_reg_33__U3 ( .A(n170), .B(data_in_2[135]), .S0(n1293), .Y(n1186) );
  DFFXL R7_reg_33_ ( .D(n1186), .CK(clk), .Q(n170), .QN(n924) );
  MX2X1 R3_reg_33__U3 ( .A(n306), .B(data_in_2[135]), .S0(n1267), .Y(n1185) );
  DFFXL R3_reg_33_ ( .D(n1185), .CK(clk), .Q(n306), .QN(n856) );
  MX2X1 R14_reg_13__U3 ( .A(n456), .B(data_in_2[81]), .S0(n1281), .Y(n1184) );
  DFFXL R14_reg_13_ ( .D(n1184), .CK(clk), .Q(n456), .QN(n774) );
  MX2X1 R10_reg_13__U3 ( .A(n524), .B(data_in_2[81]), .S0(n1256), .Y(n1183) );
  DFFXL R10_reg_13_ ( .D(n1183), .CK(clk), .Q(n524), .QN(n740) );
  MX2X1 R6_reg_13__U3 ( .A(n184), .B(data_in_2[81]), .S0(n1293), .Y(n1182) );
  DFFXL R6_reg_13_ ( .D(n1182), .CK(clk), .Q(n184), .QN(n910) );
  MX2X1 R2_reg_13__U3 ( .A(n320), .B(data_in_2[81]), .S0(n1267), .Y(n1181) );
  DFFXL R2_reg_13_ ( .D(n1181), .CK(clk), .Q(n320), .QN(n842) );
  MX2X1 R14_reg_33__U3 ( .A(n476), .B(data_in_2[101]), .S0(n1283), .Y(n1180)
         );
  DFFXL R14_reg_33_ ( .D(n1180), .CK(clk), .Q(n476), .QN(n754) );
  MX2X1 R10_reg_33__U3 ( .A(n544), .B(data_in_2[101]), .S0(n1258), .Y(n1179)
         );
  DFFXL R10_reg_33_ ( .D(n1179), .CK(clk), .Q(n544), .QN(n720) );
  DFFXL R6_reg_33_ ( .D(n1178), .CK(clk), .Q(n204), .QN(n890) );
  MX2X1 R2_reg_33__U3 ( .A(n340), .B(data_in_2[101]), .S0(n1268), .Y(n1177) );
  DFFXL R2_reg_33_ ( .D(n1177), .CK(clk), .Q(n340), .QN(n822) );
  DFFXL R12_reg_33_ ( .D(n1176), .CK(clk), .Q(R12[33]) );
  DFFXL R8_reg_33_ ( .D(n1174), .CK(clk), .Q(R8[33]) );
  DFFXL R4_reg_33_ ( .D(n1172), .CK(clk), .Q(R4[33]) );
  DFFXL R0_reg_33_ ( .D(n1170), .CK(clk), .Q(R0[33]) );
  MX2X1 R12_reg_14__U3 ( .A(R12[14]), .B(data_in_2[14]), .S0(n1284), .Y(n1168)
         );
  DFFXL R12_reg_14_ ( .D(n1168), .CK(clk), .Q(R12[14]) );
  MX2X1 R8_reg_14__U3 ( .A(R8[14]), .B(data_in_2[14]), .S0(n1262), .Y(n1166)
         );
  DFFXL R8_reg_14_ ( .D(n1166), .CK(clk), .Q(R8[14]) );
  MX2X1 R4_reg_14__U3 ( .A(R4[14]), .B(data_in_2[14]), .S0(n1289), .Y(n1164)
         );
  DFFXL R4_reg_14_ ( .D(n1164), .CK(clk), .Q(R4[14]) );
  MX2X1 R0_reg_14__U3 ( .A(R0[14]), .B(data_in_2[14]), .S0(n1264), .Y(n1162)
         );
  DFFXL R0_reg_14_ ( .D(n1162), .CK(clk), .Q(R0[14]) );
  DFFXL R12_reg_13_ ( .D(n1160), .CK(clk), .Q(R12[13]) );
  DFFXL R8_reg_13_ ( .D(n1158), .CK(clk), .Q(R8[13]) );
  DFFXL R4_reg_13_ ( .D(n1156), .CK(clk), .Q(R4[13]) );
  DFFXL R0_reg_13_ ( .D(n1154), .CK(clk), .Q(R0[13]) );
  MX2X1 R12_reg_11__U3 ( .A(R12[11]), .B(data_in_2[11]), .S0(n1284), .Y(n1152)
         );
  DFFXL R12_reg_11_ ( .D(n1152), .CK(clk), .Q(R12[11]) );
  MX2X1 R8_reg_11__U3 ( .A(R8[11]), .B(data_in_2[11]), .S0(n1262), .Y(n1150)
         );
  DFFXL R8_reg_11_ ( .D(n1150), .CK(clk), .Q(R8[11]) );
  MX2X1 R4_reg_11__U3 ( .A(R4[11]), .B(data_in_2[11]), .S0(n1290), .Y(n1148)
         );
  DFFXL R4_reg_11_ ( .D(n1148), .CK(clk), .Q(R4[11]) );
  MX2X1 R0_reg_11__U3 ( .A(R0[11]), .B(data_in_2[11]), .S0(n1265), .Y(n1146)
         );
  DFFXL R0_reg_11_ ( .D(n1146), .CK(clk), .Q(R0[11]) );
  MX2X1 R12_reg_30__U3 ( .A(R12[30]), .B(data_in_2[30]), .S0(n1285), .Y(n1144)
         );
  DFFXL R12_reg_30_ ( .D(n1144), .CK(clk), .Q(R12[30]) );
  MX2X1 R8_reg_30__U3 ( .A(R8[30]), .B(data_in_2[30]), .S0(n114), .Y(n1142) );
  DFFXL R8_reg_30_ ( .D(n1142), .CK(clk), .Q(R8[30]) );
  MX2X1 R4_reg_30__U3 ( .A(R4[30]), .B(data_in_2[30]), .S0(n1289), .Y(n1140)
         );
  DFFXL R4_reg_30_ ( .D(n1140), .CK(clk), .Q(R4[30]) );
  MX2X1 R0_reg_30__U3 ( .A(R0[30]), .B(data_in_2[30]), .S0(n1264), .Y(n1138)
         );
  DFFXL R0_reg_30_ ( .D(n1138), .CK(clk), .Q(R0[30]) );
  MX2X1 R13_reg_28__U3 ( .A(R13[28]), .B(data_in_2[62]), .S0(n1287), .Y(n1136)
         );
  DFFXL R13_reg_28_ ( .D(n1136), .CK(clk), .Q(R13[28]) );
  MX2X1 R9_reg_28__U3 ( .A(R9[28]), .B(data_in_2[62]), .S0(n1255), .Y(n1134)
         );
  DFFXL R9_reg_28_ ( .D(n1134), .CK(clk), .Q(R9[28]) );
  MX2X1 R5_reg_28__U3 ( .A(R5[28]), .B(data_in_2[62]), .S0(n1290), .Y(n1132)
         );
  DFFXL R5_reg_28_ ( .D(n1132), .CK(clk), .Q(R5[28]) );
  MX2X1 R1_reg_28__U3 ( .A(R1[28]), .B(data_in_2[62]), .S0(n1265), .Y(n1130)
         );
  DFFXL R1_reg_28_ ( .D(n1130), .CK(clk), .Q(R1[28]) );
  DFFXL R12_reg_15_ ( .D(n1128), .CK(clk), .Q(R12[15]) );
  DFFXL R8_reg_15_ ( .D(n1126), .CK(clk), .Q(R8[15]) );
  DFFXL R4_reg_15_ ( .D(n1124), .CK(clk), .Q(R4[15]) );
  DFFXL R0_reg_15_ ( .D(n1122), .CK(clk), .Q(R0[15]) );
  MX2X1 R13_reg_16__U3 ( .A(R13[16]), .B(data_in_2[50]), .S0(n1286), .Y(n1120)
         );
  DFFXL R13_reg_16_ ( .D(n1120), .CK(clk), .Q(R13[16]) );
  MX2X1 R9_reg_16__U3 ( .A(R9[16]), .B(data_in_2[50]), .S0(n1254), .Y(n1118)
         );
  DFFXL R9_reg_16_ ( .D(n1118), .CK(clk), .Q(R9[16]) );
  MX2X1 R5_reg_16__U3 ( .A(R5[16]), .B(data_in_2[50]), .S0(n1291), .Y(n977) );
  DFFXL R5_reg_16_ ( .D(n977), .CK(clk), .Q(R5[16]) );
  MX2X1 R1_reg_16__U3 ( .A(R1[16]), .B(data_in_2[50]), .S0(n1266), .Y(n970) );
  DFFXL R1_reg_16_ ( .D(n970), .CK(clk), .Q(R1[16]) );
  DFFXL R12_reg_31_ ( .D(n960), .CK(clk), .Q(R12[31]) );
  DFFXL R8_reg_31_ ( .D(n958), .CK(clk), .Q(R8[31]) );
  DFFXL R4_reg_31_ ( .D(n684), .CK(clk), .Q(R4[31]) );
  DFFXL R0_reg_31_ ( .D(n682), .CK(clk), .Q(R0[31]) );
  DFFXL R12_reg_32_ ( .D(n680), .CK(clk), .Q(R12[32]) );
  DFFXL R8_reg_32_ ( .D(n678), .CK(clk), .Q(R8[32]) );
  DFFXL R4_reg_32_ ( .D(n676), .CK(clk), .Q(R4[32]) );
  DFFXL R0_reg_32_ ( .D(n674), .CK(clk), .Q(R0[32]) );
  MX2X1 R13_reg_31__U3 ( .A(R13[31]), .B(data_in_2[65]), .S0(n1287), .Y(n672)
         );
  DFFXL R13_reg_31_ ( .D(n672), .CK(clk), .Q(R13[31]) );
  MX2X1 R9_reg_31__U3 ( .A(R9[31]), .B(data_in_2[65]), .S0(n1255), .Y(n670) );
  DFFXL R9_reg_31_ ( .D(n670), .CK(clk), .Q(R9[31]) );
  MX2X1 R5_reg_31__U3 ( .A(R5[31]), .B(data_in_2[65]), .S0(n1290), .Y(n668) );
  DFFXL R5_reg_31_ ( .D(n668), .CK(clk), .Q(R5[31]) );
  MX2X1 R1_reg_31__U3 ( .A(R1[31]), .B(data_in_2[65]), .S0(n1265), .Y(n666) );
  DFFXL R1_reg_31_ ( .D(n666), .CK(clk), .Q(R1[31]) );
  MX2X1 R13_reg_15__U3 ( .A(R13[15]), .B(data_in_2[49]), .S0(n1286), .Y(n664)
         );
  DFFXL R13_reg_15_ ( .D(n664), .CK(clk), .Q(R13[15]) );
  DFFXL R13_reg_14_ ( .D(n662), .CK(clk), .Q(R13[14]) );
  MX2X1 R9_reg_15__U3 ( .A(R9[15]), .B(data_in_2[49]), .S0(n1254), .Y(n660) );
  DFFXL R9_reg_15_ ( .D(n660), .CK(clk), .Q(R9[15]) );
  MX2X1 R9_reg_14__U3 ( .A(R9[14]), .B(data_in_2[48]), .S0(n1254), .Y(n658) );
  DFFXL R9_reg_14_ ( .D(n658), .CK(clk), .Q(R9[14]) );
  MX2X1 R5_reg_15__U3 ( .A(R5[15]), .B(data_in_2[49]), .S0(n1291), .Y(n656) );
  DFFXL R5_reg_15_ ( .D(n656), .CK(clk), .Q(R5[15]) );
  MX2X1 R5_reg_14__U3 ( .A(R5[14]), .B(data_in_2[48]), .S0(n1291), .Y(n654) );
  DFFXL R5_reg_14_ ( .D(n654), .CK(clk), .Q(R5[14]) );
  MX2X1 R1_reg_15__U3 ( .A(R1[15]), .B(data_in_2[49]), .S0(n1266), .Y(n652) );
  DFFXL R1_reg_15_ ( .D(n652), .CK(clk), .Q(R1[15]) );
  MX2X1 R1_reg_14__U3 ( .A(R1[14]), .B(data_in_2[48]), .S0(n1266), .Y(n650) );
  DFFXL R1_reg_14_ ( .D(n650), .CK(clk), .Q(R1[14]) );
  DFFXL R13_reg_32_ ( .D(n648), .CK(clk), .Q(R13[32]) );
  MX2X1 R9_reg_32__U3 ( .A(R9[32]), .B(data_in_2[66]), .S0(n1255), .Y(n646) );
  DFFXL R9_reg_32_ ( .D(n646), .CK(clk), .Q(R9[32]) );
  MX2X1 R5_reg_32__U3 ( .A(R5[32]), .B(data_in_2[66]), .S0(n1290), .Y(n644) );
  DFFXL R5_reg_32_ ( .D(n644), .CK(clk), .Q(R5[32]) );
  MX2X1 R1_reg_32__U3 ( .A(R1[32]), .B(data_in_2[66]), .S0(n1265), .Y(n642) );
  DFFXL R1_reg_32_ ( .D(n642), .CK(clk), .Q(R1[32]) );
  MX2X1 R13_reg_12__U3 ( .A(R13[12]), .B(data_in_2[46]), .S0(n1286), .Y(n640)
         );
  DFFXL R13_reg_12_ ( .D(n640), .CK(clk), .Q(R13[12]) );
  MX2X1 R9_reg_12__U3 ( .A(R9[12]), .B(data_in_2[46]), .S0(n1254), .Y(n638) );
  DFFXL R9_reg_12_ ( .D(n638), .CK(clk), .Q(R9[12]) );
  MX2X1 R1_reg_12__U3 ( .A(R1[12]), .B(data_in_2[46]), .S0(n1266), .Y(n636) );
  DFFXL R1_reg_12_ ( .D(n636), .CK(clk), .Q(R1[12]) );
  MX2X1 R13_reg_9__U3 ( .A(R13[9]), .B(data_in_2[43]), .S0(n1286), .Y(n634) );
  DFFXL R13_reg_9_ ( .D(n634), .CK(clk), .Q(R13[9]) );
  MX2X1 R9_reg_9__U3 ( .A(R9[9]), .B(data_in_2[43]), .S0(n1253), .Y(n632) );
  DFFXL R9_reg_9_ ( .D(n632), .CK(clk), .Q(R9[9]) );
  MX2X1 R5_reg_9__U3 ( .A(R5[9]), .B(data_in_2[43]), .S0(n1291), .Y(n630) );
  DFFXL R5_reg_9_ ( .D(n630), .CK(clk), .Q(R5[9]) );
  MX2X1 R1_reg_9__U3 ( .A(R1[9]), .B(data_in_2[43]), .S0(n1266), .Y(n628) );
  DFFXL R1_reg_9_ ( .D(n628), .CK(clk), .Q(R1[9]) );
  MX2X1 R13_reg_11__U3 ( .A(R13[11]), .B(data_in_2[45]), .S0(n1286), .Y(n626)
         );
  DFFXL R13_reg_11_ ( .D(n626), .CK(clk), .Q(R13[11]) );
  MX2X1 R9_reg_11__U3 ( .A(R9[11]), .B(data_in_2[45]), .S0(n1253), .Y(n624) );
  DFFXL R9_reg_11_ ( .D(n624), .CK(clk), .Q(R9[11]) );
  MX2X1 R5_reg_11__U3 ( .A(R5[11]), .B(data_in_2[45]), .S0(n1291), .Y(n622) );
  DFFXL R5_reg_11_ ( .D(n622), .CK(clk), .Q(R5[11]) );
  MX2X1 R1_reg_11__U3 ( .A(R1[11]), .B(data_in_2[45]), .S0(n1266), .Y(n620) );
  DFFXL R1_reg_11_ ( .D(n620), .CK(clk), .Q(R1[11]) );
  MX2X1 R13_reg_33__U3 ( .A(R13[33]), .B(data_in_2[67]), .S0(n1278), .Y(n618)
         );
  DFFXL R13_reg_33_ ( .D(n618), .CK(clk), .Q(R13[33]) );
  DFFXL R9_reg_33_ ( .D(n616), .CK(clk), .Q(R9[33]) );
  MX2X1 R5_reg_33__U3 ( .A(R5[33]), .B(data_in_2[67]), .S0(n1290), .Y(n614) );
  DFFXL R5_reg_33_ ( .D(n614), .CK(clk), .Q(R5[33]) );
  MX2X1 R1_reg_33__U3 ( .A(R1[33]), .B(data_in_2[67]), .S0(n1265), .Y(n612) );
  DFFXL R1_reg_33_ ( .D(n612), .CK(clk), .Q(R1[33]) );
  MX2X1 R15_reg_15__U3 ( .A(n424), .B(data_in_2[117]), .S0(n1279), .Y(n610) );
  DFFXL R15_reg_15_ ( .D(n610), .CK(clk), .Q(n424), .QN(n806) );
  MX2X1 R15_reg_14__U3 ( .A(n423), .B(data_in_2[116]), .S0(n1279), .Y(n609) );
  DFFXL R15_reg_14_ ( .D(n609), .CK(clk), .Q(n423), .QN(n807) );
  MX2X1 R11_reg_15__U3 ( .A(n560), .B(data_in_2[117]), .S0(n1259), .Y(n608) );
  DFFXL R11_reg_15_ ( .D(n608), .CK(clk), .Q(n560), .QN(n704) );
  MX2X1 R11_reg_14__U3 ( .A(n559), .B(data_in_2[116]), .S0(n1259), .Y(n607) );
  DFFXL R11_reg_14_ ( .D(n607), .CK(clk), .Q(n559), .QN(n705) );
  MX2X1 R7_reg_15__U3 ( .A(n152), .B(data_in_2[117]), .S0(n1294), .Y(n606) );
  DFFXL R7_reg_15_ ( .D(n606), .CK(clk), .Q(n152), .QN(n942) );
  MX2X1 R7_reg_14__U3 ( .A(n151), .B(data_in_2[116]), .S0(n1294), .Y(n605) );
  DFFXL R7_reg_14_ ( .D(n605), .CK(clk), .Q(n151), .QN(n943) );
  MX2X1 R3_reg_15__U3 ( .A(n288), .B(data_in_2[117]), .S0(n1268), .Y(n604) );
  DFFXL R3_reg_15_ ( .D(n604), .CK(clk), .Q(n288), .QN(n874) );
  MX2X1 R3_reg_14__U3 ( .A(n287), .B(data_in_2[116]), .S0(n1268), .Y(n603) );
  DFFXL R3_reg_14_ ( .D(n603), .CK(clk), .Q(n287), .QN(n875) );
  EDFFX1 data_out_2_reg_134_ ( .D(N186), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[134]) );
  EDFFX1 data_out_2_reg_133_ ( .D(N185), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[133]) );
  EDFFX1 data_out_2_reg_132_ ( .D(N184), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[132]) );
  EDFFX1 data_out_2_reg_131_ ( .D(N183), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[131]) );
  EDFFX1 data_out_2_reg_130_ ( .D(N182), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[130]) );
  EDFFX1 data_out_2_reg_129_ ( .D(N181), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[129]) );
  EDFFX1 data_out_2_reg_128_ ( .D(N180), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[128]) );
  EDFFX1 data_out_2_reg_127_ ( .D(N179), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[127]) );
  EDFFX1 data_out_2_reg_126_ ( .D(N178), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[126]) );
  EDFFX1 data_out_2_reg_125_ ( .D(N177), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[125]) );
  EDFFX1 data_out_2_reg_124_ ( .D(N176), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[124]) );
  EDFFX1 data_out_2_reg_123_ ( .D(N175), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[123]) );
  EDFFX1 data_out_2_reg_122_ ( .D(N174), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[122]) );
  EDFFX1 data_out_2_reg_121_ ( .D(N173), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[121]) );
  EDFFX1 data_out_2_reg_120_ ( .D(N172), .E(n1323), .CK(clk), .Q(
        data_out_2[120]) );
  EDFFX1 data_out_2_reg_117_ ( .D(N169), .E(n1322), .CK(clk), .Q(
        data_out_2[117]) );
  EDFFX1 data_out_2_reg_116_ ( .D(N168), .E(n1323), .CK(clk), .Q(
        data_out_2[116]) );
  EDFFX1 data_out_2_reg_115_ ( .D(N167), .E(n1321), .CK(clk), .Q(
        data_out_2[115]) );
  EDFFX1 data_out_2_reg_114_ ( .D(N166), .E(n1321), .CK(clk), .Q(
        data_out_2[114]) );
  EDFFX1 data_out_2_reg_113_ ( .D(N165), .E(n1322), .CK(clk), .Q(
        data_out_2[113]) );
  EDFFX1 data_out_2_reg_112_ ( .D(N164), .E(n1323), .CK(clk), .Q(
        data_out_2[112]) );
  EDFFX1 data_out_2_reg_111_ ( .D(N163), .E(n1323), .CK(clk), .Q(
        data_out_2[111]) );
  EDFFX1 data_out_2_reg_110_ ( .D(N162), .E(n1321), .CK(clk), .Q(
        data_out_2[110]) );
  EDFFX1 data_out_2_reg_109_ ( .D(N161), .E(n1322), .CK(clk), .Q(
        data_out_2[109]) );
  EDFFX1 data_out_2_reg_108_ ( .D(N160), .E(n1323), .CK(clk), .Q(
        data_out_2[108]) );
  EDFFX1 data_out_2_reg_107_ ( .D(N159), .E(n1322), .CK(clk), .Q(
        data_out_2[107]) );
  EDFFX1 data_out_2_reg_106_ ( .D(N158), .E(n1321), .CK(clk), .Q(
        data_out_2[106]) );
  EDFFX1 data_out_2_reg_105_ ( .D(N157), .E(n1322), .CK(clk), .Q(
        data_out_2[105]) );
  EDFFX1 data_out_2_reg_104_ ( .D(N156), .E(n1323), .CK(clk), .Q(
        data_out_2[104]) );
  EDFFX1 data_out_2_reg_103_ ( .D(N155), .E(n1321), .CK(clk), .Q(
        data_out_2[103]) );
  EDFFX1 data_out_2_reg_100_ ( .D(N152), .E(n1321), .CK(clk), .Q(
        data_out_2[100]) );
  EDFFX1 data_out_2_reg_99_ ( .D(N151), .E(n1322), .CK(clk), .Q(data_out_2[99]) );
  EDFFX1 data_out_2_reg_98_ ( .D(N150), .E(n1322), .CK(clk), .Q(data_out_2[98]) );
  EDFFX1 data_out_2_reg_97_ ( .D(N149), .E(n1321), .CK(clk), .Q(data_out_2[97]) );
  EDFFX1 data_out_2_reg_96_ ( .D(N148), .E(n1323), .CK(clk), .Q(data_out_2[96]) );
  EDFFX1 data_out_2_reg_95_ ( .D(N147), .E(n1322), .CK(clk), .Q(data_out_2[95]) );
  EDFFX1 data_out_2_reg_94_ ( .D(N146), .E(n1321), .CK(clk), .Q(data_out_2[94]) );
  EDFFX1 data_out_2_reg_93_ ( .D(N145), .E(n1323), .CK(clk), .Q(data_out_2[93]) );
  EDFFX1 data_out_2_reg_92_ ( .D(N144), .E(n1322), .CK(clk), .Q(data_out_2[92]) );
  EDFFX1 data_out_2_reg_91_ ( .D(N143), .E(n1321), .CK(clk), .Q(data_out_2[91]) );
  EDFFX1 data_out_2_reg_90_ ( .D(N142), .E(n1323), .CK(clk), .Q(data_out_2[90]) );
  EDFFX1 data_out_2_reg_89_ ( .D(N141), .E(n1322), .CK(clk), .Q(data_out_2[89]) );
  EDFFX1 data_out_2_reg_88_ ( .D(N140), .E(n1323), .CK(clk), .Q(data_out_2[88]) );
  EDFFX1 data_out_2_reg_87_ ( .D(N139), .E(n1321), .CK(clk), .Q(data_out_2[87]) );
  EDFFX1 data_out_2_reg_86_ ( .D(N138), .E(n1322), .CK(clk), .Q(data_out_2[86]) );
  EDFFX1 data_out_2_reg_83_ ( .D(N135), .E(n1323), .CK(clk), .Q(data_out_2[83]) );
  EDFFX1 data_out_2_reg_82_ ( .D(N134), .E(n1321), .CK(clk), .Q(data_out_2[82]) );
  EDFFX1 data_out_2_reg_81_ ( .D(N133), .E(n1322), .CK(clk), .Q(data_out_2[81]) );
  EDFFX1 data_out_2_reg_80_ ( .D(N132), .E(n1323), .CK(clk), .Q(data_out_2[80]) );
  EDFFX1 data_out_2_reg_79_ ( .D(N131), .E(n1321), .CK(clk), .Q(data_out_2[79]) );
  EDFFX1 data_out_2_reg_78_ ( .D(N130), .E(n1321), .CK(clk), .Q(data_out_2[78]) );
  EDFFX1 data_out_2_reg_77_ ( .D(N129), .E(n1321), .CK(clk), .Q(data_out_2[77]) );
  EDFFX1 data_out_2_reg_76_ ( .D(N128), .E(n1321), .CK(clk), .Q(data_out_2[76]) );
  EDFFX1 data_out_2_reg_75_ ( .D(N127), .E(n1321), .CK(clk), .Q(data_out_2[75]) );
  EDFFX1 data_out_2_reg_74_ ( .D(N126), .E(n1321), .CK(clk), .Q(data_out_2[74]) );
  EDFFX1 data_out_2_reg_73_ ( .D(N125), .E(n1321), .CK(clk), .Q(data_out_2[73]) );
  EDFFX1 data_out_2_reg_72_ ( .D(N124), .E(n1321), .CK(clk), .Q(data_out_2[72]) );
  EDFFX1 data_out_2_reg_71_ ( .D(N123), .E(n1321), .CK(clk), .Q(data_out_2[71]) );
  EDFFX1 data_out_2_reg_70_ ( .D(N122), .E(n1321), .CK(clk), .Q(data_out_2[70]) );
  EDFFX1 data_out_2_reg_69_ ( .D(N121), .E(n1321), .CK(clk), .Q(data_out_2[69]) );
  EDFFX1 data_out_2_reg_66_ ( .D(N118), .E(n1321), .CK(clk), .Q(data_out_2[66]) );
  EDFFX1 data_out_2_reg_65_ ( .D(N117), .E(n1321), .CK(clk), .Q(data_out_2[65]) );
  EDFFX1 data_out_2_reg_64_ ( .D(N116), .E(n1321), .CK(clk), .Q(data_out_2[64]) );
  EDFFX1 data_out_2_reg_63_ ( .D(N115), .E(n1321), .CK(clk), .Q(data_out_2[63]) );
  EDFFX1 data_out_2_reg_62_ ( .D(N114), .E(n1321), .CK(clk), .Q(data_out_2[62]) );
  EDFFX1 data_out_2_reg_61_ ( .D(N113), .E(n1321), .CK(clk), .Q(data_out_2[61]) );
  EDFFX1 data_out_2_reg_60_ ( .D(N112), .E(n1321), .CK(clk), .Q(data_out_2[60]) );
  EDFFX1 data_out_2_reg_59_ ( .D(N111), .E(n1322), .CK(clk), .Q(data_out_2[59]) );
  EDFFX1 data_out_2_reg_58_ ( .D(N110), .E(n1322), .CK(clk), .Q(data_out_2[58]) );
  EDFFX1 data_out_2_reg_57_ ( .D(N109), .E(n1322), .CK(clk), .Q(data_out_2[57]) );
  EDFFX1 data_out_2_reg_56_ ( .D(N108), .E(n1322), .CK(clk), .Q(data_out_2[56]) );
  EDFFX1 data_out_2_reg_55_ ( .D(N107), .E(n1322), .CK(clk), .Q(data_out_2[55]) );
  EDFFX1 data_out_2_reg_54_ ( .D(N106), .E(n1322), .CK(clk), .Q(data_out_2[54]) );
  EDFFX1 data_out_2_reg_53_ ( .D(N105), .E(n1322), .CK(clk), .Q(data_out_2[53]) );
  EDFFX1 data_out_2_reg_52_ ( .D(N104), .E(n1322), .CK(clk), .Q(data_out_2[52]) );
  EDFFX1 data_out_2_reg_49_ ( .D(N101), .E(n1322), .CK(clk), .Q(data_out_2[49]) );
  EDFFX1 data_out_2_reg_48_ ( .D(N100), .E(n1322), .CK(clk), .Q(data_out_2[48]) );
  EDFFX1 data_out_2_reg_47_ ( .D(N99), .E(n1322), .CK(clk), .Q(data_out_2[47])
         );
  EDFFX1 data_out_2_reg_46_ ( .D(N98), .E(n1322), .CK(clk), .Q(data_out_2[46])
         );
  EDFFX1 data_out_2_reg_45_ ( .D(N97), .E(n1322), .CK(clk), .Q(data_out_2[45])
         );
  EDFFX1 data_out_2_reg_44_ ( .D(N96), .E(n1322), .CK(clk), .Q(data_out_2[44])
         );
  EDFFX1 data_out_2_reg_43_ ( .D(N95), .E(n1322), .CK(clk), .Q(data_out_2[43])
         );
  EDFFX1 data_out_2_reg_42_ ( .D(N94), .E(n1322), .CK(clk), .Q(data_out_2[42])
         );
  EDFFX1 data_out_2_reg_41_ ( .D(N93), .E(n1322), .CK(clk), .Q(data_out_2[41])
         );
  EDFFX1 data_out_2_reg_40_ ( .D(N92), .E(n1322), .CK(clk), .Q(data_out_2[40])
         );
  EDFFX1 data_out_2_reg_39_ ( .D(N91), .E(n1323), .CK(clk), .Q(data_out_2[39])
         );
  EDFFX1 data_out_2_reg_38_ ( .D(N90), .E(n1322), .CK(clk), .Q(data_out_2[38])
         );
  EDFFX1 data_out_2_reg_37_ ( .D(N89), .E(n1323), .CK(clk), .Q(data_out_2[37])
         );
  EDFFX1 data_out_2_reg_36_ ( .D(N88), .E(n1321), .CK(clk), .Q(data_out_2[36])
         );
  EDFFX1 data_out_2_reg_35_ ( .D(N87), .E(n1323), .CK(clk), .Q(data_out_2[35])
         );
  EDFFX1 data_out_2_reg_119_ ( .D(N171), .E(n1322), .CK(clk), .Q(
        data_out_2[119]) );
  EDFFX1 data_out_2_reg_102_ ( .D(N154), .E(n1321), .CK(clk), .Q(
        data_out_2[102]) );
  EDFFX1 data_out_2_reg_85_ ( .D(N137), .E(n1322), .CK(clk), .Q(data_out_2[85]) );
  EDFFX1 data_out_2_reg_68_ ( .D(N120), .E(n1321), .CK(clk), .Q(data_out_2[68]) );
  EDFFX1 data_out_2_reg_51_ ( .D(N103), .E(n1322), .CK(clk), .Q(data_out_2[51]) );
  EDFFX1 data_out_2_reg_34_ ( .D(N86), .E(n1323), .CK(clk), .Q(data_out_2[34])
         );
  EDFFX1 R10_reg_23_ ( .D(data_in_2[91]), .E(n1257), .CK(clk), .QN(n730) );
  EDFFX1 R10_reg_22_ ( .D(n78), .E(n1257), .CK(clk), .QN(n731) );
  EDFFX1 R10_reg_21_ ( .D(data_in_2[89]), .E(n1257), .CK(clk), .QN(n732) );
  EDFFX1 R10_reg_20_ ( .D(data_in_2[88]), .E(n1257), .CK(clk), .QN(n733) );
  EDFFX1 R10_reg_19_ ( .D(data_in_2[87]), .E(n1257), .CK(clk), .QN(n734) );
  EDFFX1 R10_reg_18_ ( .D(data_in_2[86]), .E(n1257), .CK(clk), .QN(n735) );
  EDFFX1 R10_reg_17_ ( .D(data_in_2[85]), .E(n1257), .CK(clk), .QN(n736) );
  EDFFX1 R10_reg_8_ ( .D(data_in_2[76]), .E(n1256), .CK(clk), .QN(n745) );
  EDFFX1 R10_reg_6_ ( .D(data_in_2[74]), .E(n1256), .CK(clk), .QN(n747) );
  EDFFXL R10_reg_4_ ( .D(data_in_2[72]), .E(n1256), .CK(clk), .QN(n749) );
  EDFFX1 R10_reg_3_ ( .D(data_in_2[71]), .E(n1256), .CK(clk), .QN(n750) );
  EDFFX1 R10_reg_2_ ( .D(data_in_2[70]), .E(n1256), .CK(clk), .QN(n751) );
  EDFFX1 R10_reg_1_ ( .D(data_in_2[69]), .E(n1255), .CK(clk), .QN(n752) );
  EDFFX1 R10_reg_0_ ( .D(data_in_2[68]), .E(n1255), .CK(clk), .QN(n753) );
  EDFFX1 R14_reg_23_ ( .D(data_in_2[91]), .E(n1282), .CK(clk), .QN(n764) );
  EDFFX1 R14_reg_22_ ( .D(n78), .E(n1282), .CK(clk), .QN(n765) );
  EDFFX1 R14_reg_21_ ( .D(data_in_2[89]), .E(n1282), .CK(clk), .QN(n766) );
  EDFFX1 R14_reg_20_ ( .D(data_in_2[88]), .E(n1282), .CK(clk), .QN(n767) );
  EDFFX1 R14_reg_19_ ( .D(data_in_2[87]), .E(n1282), .CK(clk), .QN(n768) );
  EDFFX1 R14_reg_18_ ( .D(data_in_2[86]), .E(n1282), .CK(clk), .QN(n769) );
  EDFFX1 R14_reg_17_ ( .D(data_in_2[85]), .E(n1282), .CK(clk), .QN(n770) );
  EDFFX1 R14_reg_8_ ( .D(data_in_2[76]), .E(n1281), .CK(clk), .QN(n779) );
  EDFFX1 R14_reg_6_ ( .D(data_in_2[74]), .E(n1281), .CK(clk), .QN(n781) );
  EDFFXL R14_reg_4_ ( .D(data_in_2[72]), .E(n1281), .CK(clk), .QN(n783) );
  EDFFX1 R14_reg_3_ ( .D(data_in_2[71]), .E(n1281), .CK(clk), .QN(n784) );
  EDFFX1 R14_reg_2_ ( .D(data_in_2[70]), .E(n1281), .CK(clk), .QN(n785) );
  EDFFX1 R14_reg_1_ ( .D(data_in_2[69]), .E(n1280), .CK(clk), .QN(n786) );
  EDFFX1 R14_reg_0_ ( .D(data_in_2[68]), .E(n1280), .CK(clk), .QN(n787) );
  EDFFX1 R2_reg_23_ ( .D(data_in_2[91]), .E(n1265), .CK(clk), .QN(n832) );
  EDFFX1 R2_reg_22_ ( .D(data_in_2[90]), .E(n1268), .CK(clk), .QN(n833) );
  EDFFX1 R2_reg_21_ ( .D(data_in_2[89]), .E(n1267), .CK(clk), .QN(n834) );
  EDFFX1 R2_reg_20_ ( .D(data_in_2[88]), .E(n1266), .CK(clk), .QN(n835) );
  EDFFX1 R2_reg_19_ ( .D(data_in_2[87]), .E(n1265), .CK(clk), .QN(n836) );
  EDFFX1 R2_reg_18_ ( .D(data_in_2[86]), .E(n1268), .CK(clk), .QN(n837) );
  EDFFX1 R2_reg_17_ ( .D(data_in_2[85]), .E(n1267), .CK(clk), .QN(n838) );
  EDFFX1 R2_reg_8_ ( .D(data_in_2[76]), .E(n1267), .CK(clk), .QN(n847) );
  EDFFX1 R2_reg_6_ ( .D(data_in_2[74]), .E(n1267), .CK(clk), .QN(n849) );
  EDFFXL R2_reg_4_ ( .D(data_in_2[72]), .E(n1267), .CK(clk), .QN(n851) );
  EDFFX1 R2_reg_3_ ( .D(data_in_2[71]), .E(n1267), .CK(clk), .QN(n852) );
  EDFFX1 R2_reg_2_ ( .D(data_in_2[70]), .E(n1267), .CK(clk), .QN(n853) );
  EDFFX1 R2_reg_1_ ( .D(data_in_2[69]), .E(n1267), .CK(clk), .QN(n854) );
  EDFFX1 R2_reg_0_ ( .D(data_in_2[68]), .E(n1267), .CK(clk), .QN(n855) );
  EDFFXL R6_reg_29_ ( .D(data_in_2[97]), .E(n1292), .CK(clk), .QN(n894) );
  EDFFXL R6_reg_28_ ( .D(data_in_2[96]), .E(n1292), .CK(clk), .QN(n895) );
  EDFFXL R6_reg_27_ ( .D(data_in_2[95]), .E(n1292), .CK(clk), .QN(n896) );
  EDFFXL R6_reg_26_ ( .D(data_in_2[94]), .E(n1292), .CK(clk), .QN(n897) );
  EDFFXL R6_reg_25_ ( .D(data_in_2[93]), .E(n1292), .CK(clk), .QN(n898) );
  EDFFX1 R6_reg_20_ ( .D(data_in_2[88]), .E(n1292), .CK(clk), .QN(n903) );
  EDFFX1 R6_reg_19_ ( .D(data_in_2[87]), .E(n1292), .CK(clk), .QN(n904) );
  EDFFX1 R6_reg_18_ ( .D(data_in_2[86]), .E(n1293), .CK(clk), .QN(n905) );
  EDFFX1 R6_reg_17_ ( .D(data_in_2[85]), .E(n1293), .CK(clk), .QN(n906) );
  EDFFXL R6_reg_12_ ( .D(data_in_2[80]), .E(n1293), .CK(clk), .QN(n911) );
  EDFFXL R6_reg_11_ ( .D(data_in_2[79]), .E(n1293), .CK(clk), .QN(n912) );
  EDFFXL R6_reg_10_ ( .D(data_in_2[78]), .E(n1293), .CK(clk), .QN(n913) );
  EDFFXL R6_reg_9_ ( .D(data_in_2[77]), .E(n1293), .CK(clk), .QN(n914) );
  EDFFXL R6_reg_7_ ( .D(data_in_2[75]), .E(n1293), .CK(clk), .QN(n916) );
  EDFFXL R6_reg_4_ ( .D(data_in_2[72]), .E(n1293), .CK(clk), .QN(n919) );
  EDFFX1 R6_reg_3_ ( .D(data_in_2[71]), .E(n1293), .CK(clk), .QN(n920) );
  EDFFX1 R6_reg_2_ ( .D(data_in_2[70]), .E(n1293), .CK(clk), .QN(n921) );
  EDFFX1 R6_reg_1_ ( .D(data_in_2[69]), .E(n1293), .CK(clk), .QN(n922) );
  EDFFX1 R6_reg_0_ ( .D(data_in_2[68]), .E(n1293), .CK(clk), .QN(n923) );
  EDFFX1 R11_reg_25_ ( .D(data_in_2[127]), .E(n1260), .CK(clk), .QN(n694) );
  EDFFX1 R11_reg_24_ ( .D(data_in_2[126]), .E(n1260), .CK(clk), .QN(n695) );
  EDFFX1 R11_reg_23_ ( .D(data_in_2[125]), .E(n1260), .CK(clk), .QN(n696) );
  EDFFX1 R11_reg_22_ ( .D(data_in_2[124]), .E(n1260), .CK(clk), .QN(n697) );
  EDFFXL R11_reg_21_ ( .D(n2), .E(n1260), .CK(clk), .QN(n698) );
  EDFFX1 R11_reg_20_ ( .D(data_in_2[122]), .E(n1260), .CK(clk), .QN(n699) );
  EDFFX1 R11_reg_19_ ( .D(data_in_2[121]), .E(n1260), .CK(clk), .QN(n700) );
  EDFFX1 R11_reg_18_ ( .D(data_in_2[120]), .E(n1260), .CK(clk), .QN(n701) );
  EDFFX1 R11_reg_17_ ( .D(data_in_2[119]), .E(n1260), .CK(clk), .QN(n702) );
  EDFFX1 R11_reg_9_ ( .D(data_in_2[111]), .E(n1259), .CK(clk), .QN(n710) );
  EDFFX1 R11_reg_8_ ( .D(data_in_2[110]), .E(n1259), .CK(clk), .QN(n711) );
  EDFFX1 R11_reg_4_ ( .D(data_in_2[106]), .E(n1259), .CK(clk), .QN(n715) );
  EDFFX1 R11_reg_3_ ( .D(data_in_2[105]), .E(n1258), .CK(clk), .QN(n716) );
  EDFFX1 R11_reg_2_ ( .D(data_in_2[104]), .E(n1258), .CK(clk), .QN(n717) );
  EDFFX1 R11_reg_1_ ( .D(data_in_2[103]), .E(n1258), .CK(clk), .QN(n718) );
  EDFFX1 R11_reg_0_ ( .D(data_in_2[102]), .E(n1258), .CK(clk), .QN(n719) );
  EDFFX1 R15_reg_25_ ( .D(data_in_2[127]), .E(n1280), .CK(clk), .QN(n796) );
  EDFFX1 R15_reg_24_ ( .D(data_in_2[126]), .E(n1280), .CK(clk), .QN(n797) );
  EDFFX1 R15_reg_23_ ( .D(data_in_2[125]), .E(n1279), .CK(clk), .QN(n798) );
  EDFFX1 R15_reg_22_ ( .D(data_in_2[124]), .E(n1279), .CK(clk), .QN(n799) );
  EDFFXL R15_reg_21_ ( .D(n2), .E(n1279), .CK(clk), .QN(n800) );
  EDFFX1 R15_reg_20_ ( .D(data_in_2[122]), .E(n1279), .CK(clk), .QN(n801) );
  EDFFX1 R15_reg_19_ ( .D(data_in_2[121]), .E(n1279), .CK(clk), .QN(n802) );
  EDFFX1 R15_reg_18_ ( .D(data_in_2[120]), .E(n1279), .CK(clk), .QN(n803) );
  EDFFX1 R15_reg_17_ ( .D(data_in_2[119]), .E(n1279), .CK(clk), .QN(n804) );
  EDFFX1 R15_reg_9_ ( .D(data_in_2[111]), .E(n1278), .CK(clk), .QN(n812) );
  EDFFX1 R15_reg_8_ ( .D(data_in_2[110]), .E(n1278), .CK(clk), .QN(n813) );
  EDFFX1 R15_reg_4_ ( .D(data_in_2[106]), .E(n1278), .CK(clk), .QN(n817) );
  EDFFX1 R15_reg_3_ ( .D(data_in_2[105]), .E(n1278), .CK(clk), .QN(n818) );
  EDFFX1 R15_reg_2_ ( .D(data_in_2[104]), .E(n1278), .CK(clk), .QN(n819) );
  EDFFX1 R15_reg_1_ ( .D(data_in_2[103]), .E(n1278), .CK(clk), .QN(n820) );
  EDFFX1 R15_reg_0_ ( .D(data_in_2[102]), .E(n1278), .CK(clk), .QN(n821) );
  EDFFX1 R3_reg_25_ ( .D(data_in_2[127]), .E(n1268), .CK(clk), .QN(n864) );
  EDFFX1 R3_reg_24_ ( .D(data_in_2[126]), .E(n1268), .CK(clk), .QN(n865) );
  EDFFX1 R3_reg_23_ ( .D(data_in_2[125]), .E(n1268), .CK(clk), .QN(n866) );
  EDFFX1 R3_reg_22_ ( .D(data_in_2[124]), .E(n1268), .CK(clk), .QN(n867) );
  EDFFXL R3_reg_21_ ( .D(n2), .E(n1268), .CK(clk), .QN(n868) );
  EDFFX1 R3_reg_20_ ( .D(data_in_2[122]), .E(n1268), .CK(clk), .QN(n869) );
  EDFFX1 R3_reg_19_ ( .D(data_in_2[121]), .E(n1268), .CK(clk), .QN(n870) );
  EDFFX1 R3_reg_18_ ( .D(data_in_2[120]), .E(n1268), .CK(clk), .QN(n871) );
  EDFFX1 R3_reg_17_ ( .D(data_in_2[119]), .E(n1268), .CK(clk), .QN(n872) );
  EDFFX1 R3_reg_9_ ( .D(data_in_2[111]), .E(n1268), .CK(clk), .QN(n880) );
  EDFFX1 R3_reg_8_ ( .D(data_in_2[110]), .E(n1268), .CK(clk), .QN(n881) );
  EDFFX1 R3_reg_4_ ( .D(data_in_2[106]), .E(n1265), .CK(clk), .QN(n885) );
  EDFFX1 R3_reg_3_ ( .D(data_in_2[105]), .E(n1266), .CK(clk), .QN(n886) );
  EDFFX1 R3_reg_2_ ( .D(data_in_2[104]), .E(n1268), .CK(clk), .QN(n887) );
  EDFFX1 R3_reg_1_ ( .D(data_in_2[103]), .E(n1267), .CK(clk), .QN(n888) );
  EDFFX1 R3_reg_0_ ( .D(data_in_2[102]), .E(n1268), .CK(clk), .QN(n889) );
  EDFFXL R7_reg_29_ ( .D(data_in_2[131]), .E(n1294), .CK(clk), .QN(n928) );
  EDFFXL R7_reg_26_ ( .D(data_in_2[128]), .E(n1294), .CK(clk), .QN(n931) );
  EDFFXL R7_reg_21_ ( .D(n2), .E(n1294), .CK(clk), .QN(n936) );
  EDFFX1 R7_reg_20_ ( .D(data_in_2[122]), .E(n1294), .CK(clk), .QN(n937) );
  EDFFX1 R7_reg_19_ ( .D(data_in_2[121]), .E(n1294), .CK(clk), .QN(n938) );
  EDFFX1 R7_reg_18_ ( .D(data_in_2[120]), .E(n1294), .CK(clk), .QN(n939) );
  EDFFX1 R7_reg_17_ ( .D(data_in_2[119]), .E(n1294), .CK(clk), .QN(n940) );
  EDFFXL R7_reg_12_ ( .D(data_in_2[114]), .E(n1294), .CK(clk), .QN(n945) );
  EDFFXL R7_reg_11_ ( .D(data_in_2[113]), .E(n1294), .CK(clk), .QN(n946) );
  EDFFXL R7_reg_10_ ( .D(data_in_2[112]), .E(n1292), .CK(clk), .QN(n947) );
  EDFFXL R7_reg_7_ ( .D(data_in_2[109]), .E(n1294), .CK(clk), .QN(n950) );
  EDFFXL R7_reg_6_ ( .D(data_in_2[108]), .E(n1292), .CK(clk), .QN(n951) );
  EDFFXL R7_reg_4_ ( .D(data_in_2[106]), .E(n1293), .CK(clk), .QN(n953) );
  EDFFX1 R7_reg_3_ ( .D(data_in_2[105]), .E(n1294), .CK(clk), .QN(n954) );
  EDFFX1 R7_reg_2_ ( .D(data_in_2[104]), .E(n1293), .CK(clk), .QN(n955) );
  EDFFX1 R7_reg_1_ ( .D(data_in_2[103]), .E(n1292), .CK(clk), .QN(n956) );
  EDFFX1 R7_reg_0_ ( .D(data_in_2[102]), .E(n1294), .CK(clk), .QN(n957) );
  EDFFX1 R8_reg_27_ ( .D(data_in_2[27]), .E(n114), .CK(clk), .Q(R8[27]) );
  EDFFXL R8_reg_25_ ( .D(data_in_2[25]), .E(n114), .CK(clk), .Q(R8[25]) );
  EDFFX1 R8_reg_23_ ( .D(data_in_2[23]), .E(n114), .CK(clk), .Q(R8[23]) );
  EDFFX1 R8_reg_21_ ( .D(data_in_2[21]), .E(n114), .CK(clk), .Q(R8[21]) );
  EDFFX1 R8_reg_19_ ( .D(data_in_2[19]), .E(n114), .CK(clk), .Q(R8[19]) );
  EDFFX1 R8_reg_18_ ( .D(data_in_2[18]), .E(n114), .CK(clk), .Q(R8[18]) );
  EDFFX1 R8_reg_17_ ( .D(data_in_2[17]), .E(n1262), .CK(clk), .Q(R8[17]) );
  EDFFX1 R8_reg_9_ ( .D(data_in_2[9]), .E(n1262), .CK(clk), .Q(R8[9]) );
  EDFFX1 R8_reg_7_ ( .D(data_in_2[7]), .E(n1262), .CK(clk), .Q(R8[7]) );
  EDFFX1 R8_reg_6_ ( .D(data_in_2[6]), .E(n1262), .CK(clk), .Q(R8[6]) );
  EDFFX1 R8_reg_5_ ( .D(data_in_2[5]), .E(n1261), .CK(clk), .Q(R8[5]) );
  EDFFX1 R8_reg_4_ ( .D(data_in_2[4]), .E(n1261), .CK(clk), .Q(R8[4]) );
  EDFFX1 R8_reg_3_ ( .D(data_in_2[3]), .E(n1261), .CK(clk), .Q(R8[3]) );
  EDFFX1 R8_reg_2_ ( .D(data_in_2[2]), .E(n1261), .CK(clk), .Q(R8[2]) );
  EDFFX1 R8_reg_1_ ( .D(data_in_2[1]), .E(n1261), .CK(clk), .Q(R8[1]) );
  EDFFX1 R8_reg_0_ ( .D(data_in_2[0]), .E(n1261), .CK(clk), .Q(R8[0]) );
  EDFFX1 R12_reg_27_ ( .D(data_in_2[27]), .E(n1281), .CK(clk), .Q(R12[27]) );
  EDFFXL R12_reg_25_ ( .D(data_in_2[25]), .E(n1286), .CK(clk), .Q(R12[25]) );
  EDFFX1 R12_reg_23_ ( .D(data_in_2[23]), .E(n1279), .CK(clk), .Q(R12[23]) );
  EDFFX1 R12_reg_21_ ( .D(data_in_2[21]), .E(n1278), .CK(clk), .Q(R12[21]) );
  EDFFX1 R12_reg_19_ ( .D(data_in_2[19]), .E(n1280), .CK(clk), .Q(R12[19]) );
  EDFFX1 R12_reg_18_ ( .D(data_in_2[18]), .E(n1285), .CK(clk), .Q(R12[18]) );
  EDFFX1 R12_reg_17_ ( .D(data_in_2[17]), .E(n1285), .CK(clk), .Q(R12[17]) );
  EDFFX1 R12_reg_9_ ( .D(data_in_2[9]), .E(n1284), .CK(clk), .Q(R12[9]) );
  EDFFX1 R12_reg_7_ ( .D(data_in_2[7]), .E(n1284), .CK(clk), .Q(R12[7]) );
  EDFFX1 R12_reg_6_ ( .D(data_in_2[6]), .E(n1284), .CK(clk), .Q(R12[6]) );
  EDFFX1 R12_reg_5_ ( .D(data_in_2[5]), .E(n1284), .CK(clk), .Q(R12[5]) );
  EDFFX1 R12_reg_4_ ( .D(data_in_2[4]), .E(n1284), .CK(clk), .Q(R12[4]) );
  EDFFX1 R12_reg_3_ ( .D(data_in_2[3]), .E(n1283), .CK(clk), .Q(R12[3]) );
  EDFFX1 R12_reg_2_ ( .D(data_in_2[2]), .E(n1283), .CK(clk), .Q(R12[2]) );
  EDFFX1 R12_reg_1_ ( .D(data_in_2[1]), .E(n1283), .CK(clk), .Q(R12[1]) );
  EDFFX1 R12_reg_0_ ( .D(data_in_2[0]), .E(n1283), .CK(clk), .Q(R12[0]) );
  EDFFX1 R0_reg_27_ ( .D(data_in_2[27]), .E(n1264), .CK(clk), .Q(R0[27]) );
  EDFFXL R0_reg_25_ ( .D(data_in_2[25]), .E(n1264), .CK(clk), .Q(R0[25]) );
  EDFFX1 R0_reg_23_ ( .D(data_in_2[23]), .E(n1264), .CK(clk), .Q(R0[23]) );
  EDFFX1 R0_reg_21_ ( .D(data_in_2[21]), .E(n1264), .CK(clk), .Q(R0[21]) );
  EDFFX1 R0_reg_19_ ( .D(data_in_2[19]), .E(n1264), .CK(clk), .Q(R0[19]) );
  EDFFX1 R0_reg_18_ ( .D(data_in_2[18]), .E(n1264), .CK(clk), .Q(R0[18]) );
  EDFFX1 R0_reg_17_ ( .D(data_in_2[17]), .E(n1264), .CK(clk), .Q(R0[17]) );
  EDFFX1 R0_reg_9_ ( .D(data_in_2[9]), .E(n1265), .CK(clk), .Q(R0[9]) );
  EDFFX1 R0_reg_7_ ( .D(data_in_2[7]), .E(n1265), .CK(clk), .Q(R0[7]) );
  EDFFX1 R0_reg_6_ ( .D(data_in_2[6]), .E(n1265), .CK(clk), .Q(R0[6]) );
  EDFFX1 R0_reg_5_ ( .D(data_in_2[5]), .E(n1265), .CK(clk), .Q(R0[5]) );
  EDFFX1 R0_reg_4_ ( .D(data_in_2[4]), .E(n1265), .CK(clk), .Q(R0[4]) );
  EDFFX1 R0_reg_3_ ( .D(data_in_2[3]), .E(n1265), .CK(clk), .Q(R0[3]) );
  EDFFX1 R0_reg_2_ ( .D(data_in_2[2]), .E(n1265), .CK(clk), .Q(R0[2]) );
  EDFFX1 R0_reg_1_ ( .D(data_in_2[1]), .E(n1265), .CK(clk), .Q(R0[1]) );
  EDFFX1 R0_reg_0_ ( .D(data_in_2[0]), .E(n1265), .CK(clk), .Q(R0[0]) );
  EDFFXL R4_reg_29_ ( .D(data_in_2[29]), .E(n1289), .CK(clk), .Q(R4[29]) );
  EDFFXL R4_reg_28_ ( .D(data_in_2[28]), .E(n1289), .CK(clk), .Q(R4[28]) );
  EDFFXL R4_reg_27_ ( .D(n30), .E(n1289), .CK(clk), .Q(R4[27]) );
  EDFFXL R4_reg_26_ ( .D(data_in_2[26]), .E(n1289), .CK(clk), .Q(R4[26]) );
  EDFFXL R4_reg_25_ ( .D(data_in_2[25]), .E(n1289), .CK(clk), .Q(R4[25]) );
  EDFFXL R4_reg_24_ ( .D(data_in_2[24]), .E(n1289), .CK(clk), .Q(R4[24]) );
  EDFFXL R4_reg_23_ ( .D(data_in_2[23]), .E(n1289), .CK(clk), .Q(R4[23]) );
  EDFFXL R4_reg_22_ ( .D(n59), .E(n1289), .CK(clk), .Q(R4[22]) );
  EDFFXL R4_reg_21_ ( .D(data_in_2[21]), .E(n1289), .CK(clk), .Q(R4[21]) );
  EDFFX1 R4_reg_19_ ( .D(data_in_2[19]), .E(n1289), .CK(clk), .Q(R4[19]) );
  EDFFX1 R4_reg_18_ ( .D(data_in_2[18]), .E(n1289), .CK(clk), .Q(R4[18]) );
  EDFFX1 R4_reg_17_ ( .D(data_in_2[17]), .E(n1289), .CK(clk), .Q(R4[17]) );
  EDFFXL R4_reg_12_ ( .D(data_in_2[12]), .E(n1290), .CK(clk), .Q(R4[12]) );
  EDFFXL R4_reg_10_ ( .D(data_in_2[10]), .E(n1290), .CK(clk), .Q(R4[10]) );
  EDFFXL R4_reg_9_ ( .D(data_in_2[9]), .E(n1290), .CK(clk), .Q(R4[9]) );
  EDFFXL R4_reg_8_ ( .D(data_in_2[8]), .E(n1290), .CK(clk), .Q(R4[8]) );
  EDFFXL R4_reg_7_ ( .D(data_in_2[7]), .E(n1290), .CK(clk), .Q(R4[7]) );
  EDFFXL R4_reg_6_ ( .D(data_in_2[6]), .E(n1290), .CK(clk), .Q(R4[6]) );
  EDFFXL R4_reg_5_ ( .D(data_in_2[5]), .E(n1290), .CK(clk), .Q(R4[5]) );
  EDFFXL R4_reg_4_ ( .D(data_in_2[4]), .E(n1290), .CK(clk), .Q(R4[4]) );
  EDFFX1 R4_reg_3_ ( .D(data_in_2[3]), .E(n1290), .CK(clk), .Q(R4[3]) );
  EDFFX1 R4_reg_2_ ( .D(data_in_2[2]), .E(n1290), .CK(clk), .Q(R4[2]) );
  EDFFX1 R4_reg_1_ ( .D(data_in_2[1]), .E(n1290), .CK(clk), .Q(R4[1]) );
  EDFFX1 R4_reg_0_ ( .D(data_in_2[0]), .E(n1290), .CK(clk), .Q(R4[0]) );
  EDFFXL R13_reg_30_ ( .D(data_in_2[64]), .E(n1281), .CK(clk), .Q(R13[30]) );
  EDFFXL R13_reg_29_ ( .D(data_in_2[63]), .E(n1287), .CK(clk), .Q(R13[29]) );
  EDFFXL R13_reg_27_ ( .D(data_in_2[61]), .E(n1287), .CK(clk), .Q(R13[27]) );
  EDFFXL R13_reg_26_ ( .D(data_in_2[60]), .E(n1287), .CK(clk), .Q(R13[26]) );
  EDFFXL R13_reg_25_ ( .D(data_in_2[59]), .E(n1287), .CK(clk), .Q(R13[25]) );
  EDFFXL R13_reg_24_ ( .D(data_in_2[58]), .E(n1287), .CK(clk), .Q(R13[24]) );
  EDFFXL R13_reg_23_ ( .D(data_in_2[57]), .E(n1287), .CK(clk), .Q(R13[23]) );
  EDFFXL R13_reg_22_ ( .D(data_in_2[56]), .E(n1287), .CK(clk), .Q(R13[22]) );
  EDFFXL R13_reg_21_ ( .D(data_in_2[55]), .E(n1287), .CK(clk), .Q(R13[21]) );
  EDFFX1 R13_reg_20_ ( .D(data_in_2[54]), .E(n1287), .CK(clk), .Q(R13[20]) );
  EDFFX1 R13_reg_19_ ( .D(data_in_2[53]), .E(n1287), .CK(clk), .Q(R13[19]) );
  EDFFX1 R13_reg_18_ ( .D(data_in_2[52]), .E(n1287), .CK(clk), .Q(R13[18]) );
  EDFFX1 R13_reg_17_ ( .D(data_in_2[51]), .E(n1286), .CK(clk), .Q(R13[17]) );
  EDFFXL R13_reg_10_ ( .D(data_in_2[44]), .E(n1286), .CK(clk), .Q(R13[10]) );
  EDFFXL R13_reg_8_ ( .D(data_in_2[42]), .E(n1286), .CK(clk), .Q(R13[8]) );
  EDFFXL R13_reg_7_ ( .D(data_in_2[41]), .E(n1286), .CK(clk), .Q(R13[7]) );
  EDFFXL R13_reg_6_ ( .D(data_in_2[40]), .E(n1286), .CK(clk), .Q(R13[6]) );
  EDFFXL R13_reg_5_ ( .D(data_in_2[39]), .E(n1285), .CK(clk), .Q(R13[5]) );
  EDFFXL R13_reg_4_ ( .D(data_in_2[38]), .E(n1285), .CK(clk), .Q(R13[4]) );
  EDFFX1 R13_reg_3_ ( .D(data_in_2[37]), .E(n1285), .CK(clk), .Q(R13[3]) );
  EDFFX1 R13_reg_2_ ( .D(data_in_2[36]), .E(n1285), .CK(clk), .Q(R13[2]) );
  EDFFX1 R13_reg_1_ ( .D(data_in_2[35]), .E(n1285), .CK(clk), .Q(R13[1]) );
  EDFFX1 R13_reg_0_ ( .D(data_in_2[34]), .E(n1285), .CK(clk), .Q(R13[0]) );
  EDFFXL R9_reg_30_ ( .D(data_in_2[64]), .E(n1255), .CK(clk), .Q(R9[30]) );
  EDFFXL R9_reg_29_ ( .D(data_in_2[63]), .E(n1255), .CK(clk), .Q(R9[29]) );
  EDFFXL R9_reg_27_ ( .D(data_in_2[61]), .E(n1255), .CK(clk), .Q(R9[27]) );
  EDFFXL R9_reg_26_ ( .D(data_in_2[60]), .E(n1255), .CK(clk), .Q(R9[26]) );
  EDFFXL R9_reg_25_ ( .D(data_in_2[59]), .E(n1255), .CK(clk), .Q(R9[25]) );
  EDFFXL R9_reg_24_ ( .D(data_in_2[58]), .E(n1255), .CK(clk), .Q(R9[24]) );
  EDFFXL R9_reg_23_ ( .D(data_in_2[57]), .E(n1254), .CK(clk), .Q(R9[23]) );
  EDFFXL R9_reg_22_ ( .D(data_in_2[56]), .E(n1254), .CK(clk), .Q(R9[22]) );
  EDFFXL R9_reg_21_ ( .D(data_in_2[55]), .E(n1254), .CK(clk), .Q(R9[21]) );
  EDFFX1 R9_reg_20_ ( .D(data_in_2[54]), .E(n1254), .CK(clk), .Q(R9[20]) );
  EDFFX1 R9_reg_19_ ( .D(data_in_2[53]), .E(n1254), .CK(clk), .Q(R9[19]) );
  EDFFX1 R9_reg_18_ ( .D(data_in_2[52]), .E(n1254), .CK(clk), .Q(R9[18]) );
  EDFFX1 R9_reg_17_ ( .D(data_in_2[51]), .E(n1254), .CK(clk), .Q(R9[17]) );
  EDFFXL R9_reg_10_ ( .D(data_in_2[44]), .E(n1253), .CK(clk), .Q(R9[10]) );
  EDFFXL R9_reg_8_ ( .D(data_in_2[42]), .E(n1253), .CK(clk), .Q(R9[8]) );
  EDFFXL R9_reg_7_ ( .D(data_in_2[41]), .E(n1253), .CK(clk), .Q(R9[7]) );
  EDFFXL R9_reg_6_ ( .D(data_in_2[40]), .E(n1253), .CK(clk), .Q(R9[6]) );
  EDFFXL R9_reg_5_ ( .D(data_in_2[39]), .E(n1253), .CK(clk), .Q(R9[5]) );
  EDFFXL R9_reg_4_ ( .D(data_in_2[38]), .E(n1253), .CK(clk), .Q(R9[4]) );
  EDFFX1 R9_reg_3_ ( .D(data_in_2[37]), .E(n1253), .CK(clk), .Q(R9[3]) );
  EDFFX1 R9_reg_2_ ( .D(data_in_2[36]), .E(n1253), .CK(clk), .Q(R9[2]) );
  EDFFX1 R9_reg_1_ ( .D(data_in_2[35]), .E(n1253), .CK(clk), .Q(R9[1]) );
  EDFFX1 R9_reg_0_ ( .D(data_in_2[34]), .E(n1253), .CK(clk), .Q(R9[0]) );
  EDFFXL R1_reg_30_ ( .D(data_in_2[64]), .E(n1265), .CK(clk), .Q(R1[30]) );
  EDFFXL R1_reg_29_ ( .D(data_in_2[63]), .E(n1265), .CK(clk), .Q(R1[29]) );
  EDFFXL R1_reg_27_ ( .D(data_in_2[61]), .E(n1265), .CK(clk), .Q(R1[27]) );
  EDFFXL R1_reg_26_ ( .D(data_in_2[60]), .E(n1265), .CK(clk), .Q(R1[26]) );
  EDFFXL R1_reg_25_ ( .D(data_in_2[59]), .E(n1266), .CK(clk), .Q(R1[25]) );
  EDFFXL R1_reg_24_ ( .D(data_in_2[58]), .E(n1266), .CK(clk), .Q(R1[24]) );
  EDFFXL R1_reg_23_ ( .D(data_in_2[57]), .E(n1266), .CK(clk), .Q(R1[23]) );
  EDFFXL R1_reg_22_ ( .D(data_in_2[56]), .E(n1266), .CK(clk), .Q(R1[22]) );
  EDFFXL R1_reg_21_ ( .D(data_in_2[55]), .E(n1266), .CK(clk), .Q(R1[21]) );
  EDFFX1 R1_reg_20_ ( .D(data_in_2[54]), .E(n1266), .CK(clk), .Q(R1[20]) );
  EDFFX1 R1_reg_19_ ( .D(data_in_2[53]), .E(n1266), .CK(clk), .Q(R1[19]) );
  EDFFX1 R1_reg_18_ ( .D(data_in_2[52]), .E(n1266), .CK(clk), .Q(R1[18]) );
  EDFFX1 R1_reg_17_ ( .D(data_in_2[51]), .E(n1266), .CK(clk), .Q(R1[17]) );
  EDFFXL R1_reg_10_ ( .D(data_in_2[44]), .E(n1266), .CK(clk), .Q(R1[10]) );
  EDFFXL R1_reg_8_ ( .D(data_in_2[42]), .E(n1266), .CK(clk), .Q(R1[8]) );
  EDFFXL R1_reg_7_ ( .D(data_in_2[41]), .E(n1266), .CK(clk), .Q(R1[7]) );
  EDFFXL R1_reg_6_ ( .D(data_in_2[40]), .E(n1266), .CK(clk), .Q(R1[6]) );
  EDFFXL R1_reg_5_ ( .D(data_in_2[39]), .E(n1266), .CK(clk), .Q(R1[5]) );
  EDFFXL R1_reg_4_ ( .D(data_in_2[38]), .E(n1266), .CK(clk), .Q(R1[4]) );
  EDFFX1 R1_reg_3_ ( .D(data_in_2[37]), .E(n1267), .CK(clk), .Q(R1[3]) );
  EDFFX1 R1_reg_2_ ( .D(data_in_2[36]), .E(n1266), .CK(clk), .Q(R1[2]) );
  EDFFX1 R1_reg_1_ ( .D(data_in_2[35]), .E(n1265), .CK(clk), .Q(R1[1]) );
  EDFFX1 R1_reg_0_ ( .D(data_in_2[34]), .E(n1268), .CK(clk), .Q(R1[0]) );
  EDFFXL R5_reg_30_ ( .D(data_in_2[64]), .E(n1290), .CK(clk), .Q(R5[30]) );
  EDFFXL R5_reg_29_ ( .D(data_in_2[63]), .E(n1290), .CK(clk), .Q(R5[29]) );
  EDFFXL R5_reg_27_ ( .D(data_in_2[61]), .E(n1290), .CK(clk), .Q(R5[27]) );
  EDFFXL R5_reg_26_ ( .D(data_in_2[60]), .E(n1291), .CK(clk), .Q(R5[26]) );
  EDFFXL R5_reg_25_ ( .D(data_in_2[59]), .E(n1291), .CK(clk), .Q(R5[25]) );
  EDFFXL R5_reg_24_ ( .D(data_in_2[58]), .E(n1291), .CK(clk), .Q(R5[24]) );
  EDFFXL R5_reg_23_ ( .D(data_in_2[57]), .E(n1291), .CK(clk), .Q(R5[23]) );
  EDFFXL R5_reg_22_ ( .D(data_in_2[56]), .E(n1291), .CK(clk), .Q(R5[22]) );
  EDFFXL R5_reg_21_ ( .D(data_in_2[55]), .E(n1291), .CK(clk), .Q(R5[21]) );
  EDFFX1 R5_reg_20_ ( .D(data_in_2[54]), .E(n1291), .CK(clk), .Q(R5[20]) );
  EDFFX1 R5_reg_19_ ( .D(data_in_2[53]), .E(n1291), .CK(clk), .Q(R5[19]) );
  EDFFX1 R5_reg_18_ ( .D(data_in_2[52]), .E(n1291), .CK(clk), .Q(R5[18]) );
  EDFFX1 R5_reg_17_ ( .D(data_in_2[51]), .E(n1291), .CK(clk), .Q(R5[17]) );
  EDFFXL R5_reg_10_ ( .D(data_in_2[44]), .E(n1291), .CK(clk), .Q(R5[10]) );
  EDFFXL R5_reg_8_ ( .D(data_in_2[42]), .E(n1291), .CK(clk), .Q(R5[8]) );
  EDFFXL R5_reg_7_ ( .D(data_in_2[41]), .E(n1291), .CK(clk), .Q(R5[7]) );
  EDFFXL R5_reg_6_ ( .D(data_in_2[40]), .E(n1291), .CK(clk), .Q(R5[6]) );
  EDFFXL R5_reg_5_ ( .D(data_in_2[39]), .E(n1292), .CK(clk), .Q(R5[5]) );
  EDFFXL R5_reg_4_ ( .D(data_in_2[38]), .E(n1292), .CK(clk), .Q(R5[4]) );
  EDFFX1 R5_reg_3_ ( .D(data_in_2[37]), .E(n1292), .CK(clk), .Q(R5[3]) );
  EDFFX1 R5_reg_2_ ( .D(data_in_2[36]), .E(n1292), .CK(clk), .Q(R5[2]) );
  EDFFX1 R5_reg_1_ ( .D(data_in_2[35]), .E(n1292), .CK(clk), .Q(R5[1]) );
  EDFFX1 R5_reg_0_ ( .D(data_in_2[34]), .E(n1292), .CK(clk), .Q(R5[0]) );
  DFFHQX1 counter1_reg_1_ ( .D(n1115), .CK(clk), .Q(counter1[1]) );
  DFFHQX1 reg_flag_mux_reg ( .D(n1325), .CK(clk), .Q(reg_flag_mux) );
  DFFHQX1 counter2_reg_0_ ( .D(n1114), .CK(clk), .Q(counter2[0]) );
  DFFHQX1 counter2_reg_1_ ( .D(n1113), .CK(clk), .Q(counter2[1]) );
  EDFFX1 data_out_2_reg_16_ ( .D(N68), .E(n1323), .CK(clk), .Q(data_out_2[16])
         );
  EDFFX1 data_out_2_reg_33_ ( .D(N85), .E(n1322), .CK(clk), .Q(data_out_2[33])
         );
  EDFFX1 data_out_2_reg_32_ ( .D(N84), .E(n1322), .CK(clk), .Q(data_out_2[32])
         );
  EDFFX1 data_out_2_reg_31_ ( .D(N83), .E(n1321), .CK(clk), .Q(data_out_2[31])
         );
  EDFFX1 data_out_2_reg_15_ ( .D(N67), .E(n1323), .CK(clk), .Q(data_out_2[15])
         );
  EDFFX1 data_out_2_reg_14_ ( .D(N66), .E(n1323), .CK(clk), .Q(data_out_2[14])
         );
  EDFFX1 data_out_2_reg_13_ ( .D(N65), .E(n1323), .CK(clk), .Q(data_out_2[13])
         );
  EDFFX1 data_out_2_reg_24_ ( .D(N76), .E(n1321), .CK(clk), .Q(data_out_2[24])
         );
  EDFFX1 data_out_2_reg_22_ ( .D(N74), .E(n1323), .CK(clk), .Q(data_out_2[22])
         );
  EDFFX1 data_out_2_reg_7_ ( .D(N59), .E(n1323), .CK(clk), .Q(data_out_2[7])
         );
  EDFFX1 data_out_2_reg_30_ ( .D(N82), .E(n1322), .CK(clk), .Q(data_out_2[30])
         );
  EDFFX1 data_out_2_reg_29_ ( .D(N81), .E(n1321), .CK(clk), .Q(data_out_2[29])
         );
  EDFFX1 data_out_2_reg_28_ ( .D(N80), .E(n1321), .CK(clk), .Q(data_out_2[28])
         );
  EDFFX1 data_out_2_reg_27_ ( .D(N79), .E(n1322), .CK(clk), .Q(data_out_2[27])
         );
  EDFFX1 data_out_2_reg_26_ ( .D(N78), .E(n1323), .CK(clk), .Q(data_out_2[26])
         );
  EDFFX1 data_out_2_reg_25_ ( .D(N77), .E(n1322), .CK(clk), .Q(data_out_2[25])
         );
  EDFFX1 data_out_2_reg_23_ ( .D(N75), .E(n1321), .CK(clk), .Q(data_out_2[23])
         );
  EDFFX1 data_out_2_reg_21_ ( .D(N73), .E(n1321), .CK(clk), .Q(data_out_2[21])
         );
  EDFFX1 data_out_2_reg_20_ ( .D(N72), .E(n1323), .CK(clk), .Q(data_out_2[20])
         );
  EDFFX1 data_out_2_reg_17_ ( .D(N69), .E(n1323), .CK(clk), .Q(data_out_2[17])
         );
  EDFFX1 data_out_2_reg_12_ ( .D(N64), .E(n1323), .CK(clk), .Q(data_out_2[12])
         );
  EDFFX1 data_out_2_reg_11_ ( .D(N63), .E(n1323), .CK(clk), .Q(data_out_2[11])
         );
  EDFFX1 data_out_2_reg_10_ ( .D(N62), .E(n1323), .CK(clk), .Q(data_out_2[10])
         );
  EDFFX1 data_out_2_reg_9_ ( .D(N61), .E(n1323), .CK(clk), .Q(data_out_2[9])
         );
  EDFFX1 data_out_2_reg_8_ ( .D(N60), .E(n1323), .CK(clk), .Q(data_out_2[8])
         );
  EDFFX1 data_out_2_reg_6_ ( .D(N58), .E(n1323), .CK(clk), .Q(data_out_2[6])
         );
  EDFFX1 data_out_2_reg_5_ ( .D(N57), .E(n1323), .CK(clk), .Q(data_out_2[5])
         );
  EDFFX1 data_out_2_reg_4_ ( .D(N56), .E(n1323), .CK(clk), .Q(data_out_2[4])
         );
  EDFFX1 data_out_2_reg_19_ ( .D(N71), .E(n1323), .CK(clk), .Q(data_out_2[19])
         );
  EDFFX1 data_out_2_reg_18_ ( .D(N70), .E(n1323), .CK(clk), .Q(data_out_2[18])
         );
  EDFFX1 data_out_2_reg_3_ ( .D(N55), .E(n1323), .CK(clk), .Q(data_out_2[3])
         );
  EDFFX1 data_out_2_reg_2_ ( .D(N54), .E(n1323), .CK(clk), .Q(data_out_2[2])
         );
  EDFFX1 data_out_2_reg_1_ ( .D(N53), .E(n1323), .CK(clk), .Q(data_out_2[1])
         );
  EDFFX1 data_out_2_reg_0_ ( .D(N52), .E(n1322), .CK(clk), .Q(data_out_2[0])
         );
  EDFFX1 data_out_2_reg_118_ ( .D(N170), .E(n1321), .CK(clk), .Q(
        data_out_2[118]) );
  EDFFX1 data_out_2_reg_135_ ( .D(N187), .E(n1323), .CK(clk), .Q(
        data_out_2[135]) );
  EDFFX1 data_out_2_reg_50_ ( .D(N102), .E(n1322), .CK(clk), .Q(data_out_2[50]) );
  EDFFXL R8_reg_24_ ( .D(data_in_2[24]), .E(n114), .CK(clk), .Q(R8[24]) );
  EDFFXL R0_reg_24_ ( .D(data_in_2[24]), .E(n1264), .CK(clk), .Q(R0[24]) );
  EDFFXL R12_reg_24_ ( .D(data_in_2[24]), .E(n1280), .CK(clk), .Q(R12[24]) );
  EDFFXL R8_reg_20_ ( .D(data_in_2[20]), .E(n114), .CK(clk), .Q(R8[20]) );
  EDFFXL R12_reg_20_ ( .D(data_in_2[20]), .E(n1282), .CK(clk), .Q(R12[20]) );
  EDFFXL R0_reg_20_ ( .D(data_in_2[20]), .E(n1264), .CK(clk), .Q(R0[20]) );
  EDFFXL R4_reg_20_ ( .D(data_in_2[20]), .E(n1289), .CK(clk), .Q(R4[20]) );
  EDFFXL R11_reg_11_ ( .D(data_in_2[113]), .E(n1259), .CK(clk), .QN(n708) );
  EDFFXL R3_reg_11_ ( .D(data_in_2[113]), .E(n1268), .CK(clk), .QN(n878) );
  EDFFXL R15_reg_11_ ( .D(data_in_2[113]), .E(n1278), .CK(clk), .QN(n810) );
  EDFFXL R3_reg_29_ ( .D(data_in_2[131]), .E(n1267), .CK(clk), .QN(n860) );
  EDFFXL R15_reg_29_ ( .D(data_in_2[131]), .E(n1280), .CK(clk), .QN(n792) );
  EDFFXL R11_reg_29_ ( .D(data_in_2[131]), .E(n1261), .CK(clk), .QN(n690) );
  EDFFXL R3_reg_10_ ( .D(data_in_2[112]), .E(n1268), .CK(clk), .QN(n879) );
  EDFFXL R15_reg_10_ ( .D(data_in_2[112]), .E(n1278), .CK(clk), .QN(n811) );
  EDFFXL R11_reg_10_ ( .D(data_in_2[112]), .E(n1259), .CK(clk), .QN(n709) );
  EDFFXL R10_reg_12_ ( .D(data_in_2[80]), .E(n1256), .CK(clk), .QN(n741) );
  EDFFXL R14_reg_12_ ( .D(data_in_2[80]), .E(n1281), .CK(clk), .QN(n775) );
  EDFFXL R2_reg_12_ ( .D(data_in_2[80]), .E(n1267), .CK(clk), .QN(n843) );
  EDFFXL R10_reg_28_ ( .D(data_in_2[96]), .E(n1258), .CK(clk), .QN(n725) );
  EDFFXL R14_reg_28_ ( .D(data_in_2[96]), .E(n1283), .CK(clk), .QN(n759) );
  EDFFXL R2_reg_28_ ( .D(data_in_2[96]), .E(n115), .CK(clk), .QN(n827) );
  EDFFXL R11_reg_12_ ( .D(data_in_2[114]), .E(n1259), .CK(clk), .QN(n707) );
  EDFFXL R15_reg_12_ ( .D(data_in_2[114]), .E(n1279), .CK(clk), .QN(n809) );
  EDFFXL R3_reg_12_ ( .D(data_in_2[114]), .E(n1268), .CK(clk), .QN(n877) );
  EDFFXL R11_reg_7_ ( .D(data_in_2[109]), .E(n1259), .CK(clk), .QN(n712) );
  EDFFXL R15_reg_7_ ( .D(data_in_2[109]), .E(n1278), .CK(clk), .QN(n814) );
  EDFFXL R3_reg_7_ ( .D(data_in_2[109]), .E(n1268), .CK(clk), .QN(n882) );
  EDFFXL R10_reg_27_ ( .D(data_in_2[95]), .E(n1258), .CK(clk), .QN(n726) );
  EDFFXL R14_reg_27_ ( .D(data_in_2[95]), .E(n1283), .CK(clk), .QN(n760) );
  EDFFXL R2_reg_27_ ( .D(data_in_2[95]), .E(n115), .CK(clk), .QN(n828) );
  EDFFXL R10_reg_7_ ( .D(data_in_2[75]), .E(n1256), .CK(clk), .QN(n746) );
  EDFFXL R14_reg_7_ ( .D(data_in_2[75]), .E(n1281), .CK(clk), .QN(n780) );
  EDFFXL R2_reg_7_ ( .D(data_in_2[75]), .E(n1267), .CK(clk), .QN(n848) );
  EDFFX1 R7_reg_24_ ( .D(data_in_2[126]), .E(n1294), .CK(clk), .QN(n933) );
  EDFFXL R11_reg_26_ ( .D(data_in_2[128]), .E(n1260), .CK(clk), .QN(n693) );
  EDFFXL R15_reg_26_ ( .D(data_in_2[128]), .E(n1280), .CK(clk), .QN(n795) );
  EDFFXL R3_reg_26_ ( .D(data_in_2[128]), .E(n1268), .CK(clk), .QN(n863) );
  EDFFXL R8_reg_10_ ( .D(data_in_2[10]), .E(n1262), .CK(clk), .Q(R8[10]) );
  EDFFXL R12_reg_10_ ( .D(data_in_2[10]), .E(n1284), .CK(clk), .Q(R12[10]) );
  EDFFXL R0_reg_10_ ( .D(data_in_2[10]), .E(n1265), .CK(clk), .Q(R0[10]) );
  EDFFXL R10_reg_29_ ( .D(data_in_2[97]), .E(n1258), .CK(clk), .QN(n724) );
  EDFFXL R14_reg_29_ ( .D(data_in_2[97]), .E(n1283), .CK(clk), .QN(n758) );
  EDFFXL R2_reg_29_ ( .D(data_in_2[97]), .E(n115), .CK(clk), .QN(n826) );
  EDFFXL R10_reg_10_ ( .D(data_in_2[78]), .E(n1256), .CK(clk), .QN(n743) );
  EDFFXL R14_reg_10_ ( .D(data_in_2[78]), .E(n1281), .CK(clk), .QN(n777) );
  EDFFXL R2_reg_10_ ( .D(data_in_2[78]), .E(n1267), .CK(clk), .QN(n845) );
  EDFFXL R8_reg_22_ ( .D(n59), .E(n114), .CK(clk), .Q(R8[22]) );
  EDFFXL R12_reg_22_ ( .D(n59), .E(n1285), .CK(clk), .Q(R12[22]) );
  EDFFXL R0_reg_22_ ( .D(n59), .E(n1264), .CK(clk), .Q(R0[22]) );
  EDFFXL R10_reg_25_ ( .D(data_in_2[93]), .E(n1257), .CK(clk), .QN(n728) );
  EDFFXL R14_reg_25_ ( .D(data_in_2[93]), .E(n1282), .CK(clk), .QN(n762) );
  EDFFXL R2_reg_25_ ( .D(data_in_2[93]), .E(n115), .CK(clk), .QN(n830) );
  EDFFXL R10_reg_26_ ( .D(data_in_2[94]), .E(n1258), .CK(clk), .QN(n727) );
  EDFFXL R14_reg_26_ ( .D(data_in_2[94]), .E(n1283), .CK(clk), .QN(n761) );
  EDFFXL R2_reg_26_ ( .D(data_in_2[94]), .E(n115), .CK(clk), .QN(n829) );
  EDFFXL R10_reg_11_ ( .D(data_in_2[79]), .E(n1256), .CK(clk), .QN(n742) );
  EDFFXL R14_reg_11_ ( .D(data_in_2[79]), .E(n1281), .CK(clk), .QN(n776) );
  EDFFXL R2_reg_11_ ( .D(data_in_2[79]), .E(n1267), .CK(clk), .QN(n844) );
  EDFFXL R11_reg_6_ ( .D(data_in_2[108]), .E(n1259), .CK(clk), .QN(n713) );
  EDFFXL R15_reg_6_ ( .D(data_in_2[108]), .E(n1278), .CK(clk), .QN(n815) );
  EDFFXL R3_reg_6_ ( .D(data_in_2[108]), .E(n1268), .CK(clk), .QN(n883) );
  EDFFXL R8_reg_8_ ( .D(data_in_2[8]), .E(n1262), .CK(clk), .Q(R8[8]) );
  EDFFXL R12_reg_8_ ( .D(data_in_2[8]), .E(n1284), .CK(clk), .Q(R12[8]) );
  EDFFXL R0_reg_8_ ( .D(data_in_2[8]), .E(n1265), .CK(clk), .Q(R0[8]) );
  EDFFXL R8_reg_12_ ( .D(data_in_2[12]), .E(n1262), .CK(clk), .Q(R8[12]) );
  EDFFXL R12_reg_12_ ( .D(data_in_2[12]), .E(n1284), .CK(clk), .Q(R12[12]) );
  EDFFXL R0_reg_12_ ( .D(data_in_2[12]), .E(n1265), .CK(clk), .Q(R0[12]) );
  EDFFXL R8_reg_26_ ( .D(data_in_2[26]), .E(n114), .CK(clk), .Q(R8[26]) );
  EDFFXL R12_reg_26_ ( .D(data_in_2[26]), .E(n1283), .CK(clk), .Q(R12[26]) );
  EDFFXL R0_reg_26_ ( .D(data_in_2[26]), .E(n1264), .CK(clk), .Q(R0[26]) );
  EDFFXL R10_reg_9_ ( .D(data_in_2[77]), .E(n1256), .CK(clk), .QN(n744) );
  EDFFXL R14_reg_9_ ( .D(data_in_2[77]), .E(n1281), .CK(clk), .QN(n778) );
  EDFFXL R2_reg_9_ ( .D(data_in_2[77]), .E(n1267), .CK(clk), .QN(n846) );
  EDFFXL R8_reg_28_ ( .D(data_in_2[28]), .E(n114), .CK(clk), .Q(R8[28]) );
  EDFFXL R12_reg_28_ ( .D(data_in_2[28]), .E(n1285), .CK(clk), .Q(R12[28]) );
  EDFFXL R0_reg_28_ ( .D(data_in_2[28]), .E(n1264), .CK(clk), .Q(R0[28]) );
  EDFFXL R8_reg_29_ ( .D(data_in_2[29]), .E(n114), .CK(clk), .Q(R8[29]) );
  EDFFXL R12_reg_29_ ( .D(data_in_2[29]), .E(n1285), .CK(clk), .Q(R12[29]) );
  EDFFXL R0_reg_29_ ( .D(data_in_2[29]), .E(n1264), .CK(clk), .Q(R0[29]) );
  DFFXL counter1_reg_0_ ( .D(n1116), .CK(clk), .Q(counter1[0]), .QN(n1326) );
  EDFFXL R7_reg_23_ ( .D(data_in_2[125]), .E(n969), .CK(clk), .QN(n934) );
  EDFFXL R7_reg_22_ ( .D(data_in_2[124]), .E(n969), .CK(clk), .QN(n935) );
  EDFFXL R14_reg_5_ ( .D(data_in_2[73]), .E(n971), .CK(clk), .QN(n782) );
  EDFFXL R10_reg_5_ ( .D(data_in_2[73]), .E(n114), .CK(clk), .QN(n748) );
  EDFFXL R6_reg_5_ ( .D(data_in_2[73]), .E(n969), .CK(clk), .QN(n918) );
  EDFFXL R2_reg_5_ ( .D(data_in_2[73]), .E(n115), .CK(clk), .QN(n850) );
  EDFFXL R6_reg_23_ ( .D(data_in_2[91]), .E(n969), .CK(clk), .QN(n900) );
  EDFFXL R6_reg_6_ ( .D(data_in_2[74]), .E(n969), .CK(clk), .QN(n917) );
  EDFFXL R6_reg_8_ ( .D(data_in_2[76]), .E(n969), .CK(clk), .QN(n915) );
  EDFFXL R7_reg_25_ ( .D(data_in_2[127]), .E(n969), .CK(clk), .QN(n932) );
  EDFFXL R7_reg_9_ ( .D(data_in_2[111]), .E(n969), .CK(clk), .QN(n948) );
  EDFFXL R7_reg_8_ ( .D(data_in_2[110]), .E(n969), .CK(clk), .QN(n949) );
  EDFFXL R6_reg_22_ ( .D(data_in_2[90]), .E(n969), .CK(clk), .QN(n901) );
  EDFFXL R15_reg_5_ ( .D(data_in_2[107]), .E(n971), .CK(clk), .QN(n816) );
  EDFFXL R11_reg_5_ ( .D(data_in_2[107]), .E(n114), .CK(clk), .QN(n714) );
  EDFFXL R7_reg_5_ ( .D(data_in_2[107]), .E(n969), .CK(clk), .QN(n952) );
  EDFFXL R3_reg_5_ ( .D(data_in_2[107]), .E(n115), .CK(clk), .QN(n884) );
  EDFFXL R15_reg_27_ ( .D(data_in_2[129]), .E(n971), .CK(clk), .QN(n794) );
  EDFFXL R11_reg_27_ ( .D(data_in_2[129]), .E(n114), .CK(clk), .QN(n692) );
  EDFFXL R7_reg_27_ ( .D(data_in_2[129]), .E(n969), .CK(clk), .QN(n930) );
  EDFFXL R3_reg_27_ ( .D(data_in_2[129]), .E(n115), .CK(clk), .QN(n862) );
  EDFFXL R5_reg_12_ ( .D(data_in_2[46]), .E(n1291), .CK(clk), .Q(R5[12]) );
  EDFFX1 data_out_2_reg_101_ ( .D(N153), .E(n1323), .CK(clk), .Q(
        data_out_2[101]) );
  EDFFX2 data_out_2_reg_84_ ( .D(N136), .E(n1321), .CK(clk), .Q(data_out_2[84]) );
  EDFFX1 data_out_2_reg_67_ ( .D(N119), .E(n1321), .CK(clk), .Q(data_out_2[67]) );
  EDFFX1 R6_reg_21_ ( .D(data_in_2[89]), .E(n969), .CK(clk), .QN(n902) );
  MX2X1 U3 ( .A(data_in_2[48]), .B(R13[14]), .S0(n1288), .Y(n662) );
  BUFX3 U4 ( .A(data_in_2[123]), .Y(n2) );
  INVX1 U5 ( .A(n58), .Y(n59) );
  INVX1 U6 ( .A(data_in_2[22]), .Y(n58) );
  BUFX4 U7 ( .A(data_in_2[90]), .Y(n78) );
  MX2X1 U8 ( .A(n303), .B(data_in_2[132]), .S0(n1267), .Y(n1209) );
  MX2X1 U9 ( .A(n167), .B(data_in_2[132]), .S0(n1294), .Y(n1210) );
  MX2X1 U10 ( .A(n575), .B(data_in_2[132]), .S0(n1261), .Y(n1211) );
  MX2X1 U11 ( .A(n439), .B(data_in_2[132]), .S0(n1280), .Y(n1212) );
  OR2X2 U12 ( .A(counter2[0]), .B(counter2[1]), .Y(n6) );
  OR2X2 U13 ( .A(n1328), .B(counter2[1]), .Y(n7) );
  NOR2X2 U14 ( .A(n973), .B(n1327), .Y(n969) );
  BUFX1 U15 ( .A(data_in_2[27]), .Y(n30) );
  MX2X1 U16 ( .A(R13[32]), .B(data_in_2[66]), .S0(n1287), .Y(n648) );
  MX2X1 U17 ( .A(n441), .B(data_in_2[134]), .S0(n1280), .Y(n1216) );
  MX2X1 U18 ( .A(n204), .B(data_in_2[101]), .S0(n1292), .Y(n1178) );
  MX2X2 U19 ( .A(R4[31]), .B(data_in_2[31]), .S0(n1289), .Y(n684) );
  MX2X2 U20 ( .A(R0[31]), .B(data_in_2[31]), .S0(n1264), .Y(n682) );
  MX2X2 U21 ( .A(R8[31]), .B(data_in_2[31]), .S0(n1256), .Y(n958) );
  MX2X2 U22 ( .A(data_in_2[31]), .B(R12[31]), .S0(n1288), .Y(n960) );
  MX2X2 U23 ( .A(R0[13]), .B(data_in_2[13]), .S0(n1265), .Y(n1154) );
  MX2X2 U24 ( .A(R4[13]), .B(data_in_2[13]), .S0(n1290), .Y(n1156) );
  MX2X2 U25 ( .A(n185), .B(data_in_2[82]), .S0(n1293), .Y(n1234) );
  MX2X2 U26 ( .A(n321), .B(data_in_2[82]), .S0(n1267), .Y(n1233) );
  MX2X2 U27 ( .A(n525), .B(data_in_2[82]), .S0(n1257), .Y(n1235) );
  MX2X2 U28 ( .A(n457), .B(data_in_2[82]), .S0(n1282), .Y(n1236) );
  MX2X2 U29 ( .A(R4[33]), .B(data_in_2[33]), .S0(n1289), .Y(n1172) );
  MX2X2 U30 ( .A(R0[33]), .B(data_in_2[33]), .S0(n1264), .Y(n1170) );
  MX2X2 U31 ( .A(R8[33]), .B(data_in_2[33]), .S0(n1259), .Y(n1174) );
  MX2X2 U32 ( .A(data_in_2[33]), .B(R12[33]), .S0(n1288), .Y(n1176) );
  MX2X2 U33 ( .A(R8[13]), .B(data_in_2[13]), .S0(n1262), .Y(n1158) );
  MX2X2 U34 ( .A(R12[13]), .B(data_in_2[13]), .S0(n1284), .Y(n1160) );
  MX2X2 U35 ( .A(R8[15]), .B(data_in_2[15]), .S0(n1262), .Y(n1126) );
  MX2X2 U36 ( .A(R12[15]), .B(data_in_2[15]), .S0(n1284), .Y(n1128) );
  MX2X2 U37 ( .A(R4[15]), .B(data_in_2[15]), .S0(n1289), .Y(n1124) );
  MX2X2 U38 ( .A(R0[15]), .B(data_in_2[15]), .S0(n1264), .Y(n1122) );
  MX2X2 U39 ( .A(R12[32]), .B(data_in_2[32]), .S0(n1285), .Y(n680) );
  MX2X2 U40 ( .A(R4[32]), .B(data_in_2[32]), .S0(n1289), .Y(n676) );
  MX2X2 U41 ( .A(R0[32]), .B(data_in_2[32]), .S0(n1264), .Y(n674) );
  MX2X2 U42 ( .A(R8[32]), .B(data_in_2[32]), .S0(n1260), .Y(n678) );
  MX2X1 U43 ( .A(R9[33]), .B(data_in_2[67]), .S0(n1255), .Y(n616) );
  CLKINVX3 U44 ( .A(n1295), .Y(n1293) );
  CLKINVX3 U45 ( .A(n1295), .Y(n1290) );
  CLKINVX3 U46 ( .A(n1295), .Y(n1294) );
  CLKINVX3 U47 ( .A(n1295), .Y(n1292) );
  CLKINVX3 U48 ( .A(n1295), .Y(n1291) );
  CLKINVX3 U49 ( .A(n1295), .Y(n1289) );
  INVX1 U50 ( .A(n1288), .Y(n1278) );
  INVX1 U51 ( .A(n1288), .Y(n1281) );
  INVX1 U52 ( .A(n1288), .Y(n1287) );
  INVX1 U53 ( .A(n1288), .Y(n1279) );
  INVX1 U54 ( .A(n1288), .Y(n1282) );
  INVX1 U55 ( .A(n1288), .Y(n1284) );
  INVX1 U56 ( .A(n1288), .Y(n1285) );
  INVX1 U57 ( .A(n1288), .Y(n1280) );
  INVX1 U58 ( .A(n1288), .Y(n1283) );
  INVX1 U59 ( .A(n1288), .Y(n1286) );
  INVX1 U60 ( .A(n969), .Y(n1295) );
  INVX1 U61 ( .A(n7), .Y(n1312) );
  INVX1 U62 ( .A(n7), .Y(n1306) );
  INVX1 U63 ( .A(n7), .Y(n1307) );
  INVX1 U64 ( .A(n7), .Y(n1309) );
  INVX1 U65 ( .A(n7), .Y(n1310) );
  INVX1 U66 ( .A(n7), .Y(n1311) );
  CLKINVX3 U67 ( .A(n1269), .Y(n1268) );
  CLKINVX3 U68 ( .A(n1269), .Y(n1265) );
  CLKINVX3 U69 ( .A(n1269), .Y(n1267) );
  CLKINVX3 U70 ( .A(n1269), .Y(n1266) );
  INVX1 U71 ( .A(n7), .Y(n1305) );
  INVX1 U72 ( .A(n7), .Y(n1308) );
  INVX1 U73 ( .A(n6), .Y(n1276) );
  INVX1 U74 ( .A(n6), .Y(n1277) );
  INVX1 U75 ( .A(n6), .Y(n1270) );
  INVX1 U76 ( .A(n6), .Y(n1273) );
  INVX1 U77 ( .A(n6), .Y(n1274) );
  INVX1 U78 ( .A(n6), .Y(n1275) );
  INVX1 U79 ( .A(n6), .Y(n1271) );
  INVX1 U80 ( .A(n6), .Y(n1272) );
  INVX1 U81 ( .A(n1320), .Y(n1314) );
  INVX1 U82 ( .A(n1320), .Y(n1313) );
  INVX1 U83 ( .A(n1320), .Y(n1319) );
  INVX1 U84 ( .A(n1320), .Y(n1318) );
  INVX1 U85 ( .A(n1320), .Y(n1317) );
  INVX1 U86 ( .A(n1320), .Y(n1316) );
  INVX1 U87 ( .A(n1320), .Y(n1315) );
  INVX1 U88 ( .A(n1303), .Y(n1300) );
  INVX1 U89 ( .A(n1303), .Y(n1301) );
  INVX1 U90 ( .A(n1303), .Y(n1302) );
  INVX1 U91 ( .A(n1303), .Y(n1296) );
  INVX1 U92 ( .A(n1303), .Y(n1297) );
  INVX1 U93 ( .A(n1303), .Y(n1298) );
  INVX1 U94 ( .A(n1303), .Y(n1299) );
  INVX1 U95 ( .A(n1263), .Y(n1256) );
  INVX1 U96 ( .A(n1263), .Y(n1260) );
  INVX1 U97 ( .A(n1263), .Y(n1253) );
  INVX1 U98 ( .A(n1263), .Y(n1259) );
  INVX1 U99 ( .A(n1263), .Y(n1255) );
  INVX1 U100 ( .A(n1263), .Y(n1257) );
  INVX1 U101 ( .A(n1263), .Y(n1261) );
  INVX1 U102 ( .A(n1263), .Y(n1258) );
  INVX1 U103 ( .A(n1263), .Y(n1254) );
  INVX1 U104 ( .A(n1263), .Y(n1262) );
  INVX1 U105 ( .A(n966), .Y(n1329) );
  INVX1 U106 ( .A(n971), .Y(n1288) );
  NOR2X1 U107 ( .A(n1327), .B(n1326), .Y(n964) );
  INVX1 U108 ( .A(n7), .Y(n1304) );
  CLKINVX3 U109 ( .A(n1269), .Y(n1264) );
  INVX1 U110 ( .A(n115), .Y(n1269) );
  CLKINVX3 U111 ( .A(n1324), .Y(n1322) );
  CLKINVX3 U112 ( .A(n1324), .Y(n1321) );
  CLKINVX3 U113 ( .A(n1324), .Y(n1323) );
  INVX1 U114 ( .A(n968), .Y(n1303) );
  INVX1 U115 ( .A(n114), .Y(n1263) );
  INVX1 U116 ( .A(n963), .Y(n1320) );
  OAI32X1 U117 ( .A0(n961), .A1(counter2[0]), .A2(n966), .B0(n1328), .B1(n1329), .Y(n1114) );
  NOR2X1 U118 ( .A(n961), .B(reg_flag_mux), .Y(n966) );
  OAI22X1 U119 ( .A0(n1326), .A1(n974), .B0(n961), .B1(n973), .Y(n1116) );
  NAND2BX1 U120 ( .AN(reg_datain_flag), .B(rst_n), .Y(n974) );
  OAI21XL U121 ( .A0(n1327), .A1(n974), .B0(n975), .Y(n1115) );
  OAI21XL U122 ( .A0(n1264), .A1(n1289), .B0(rst_n), .Y(n975) );
  OAI2BB2X1 U123 ( .B0(n965), .B1(n961), .A0N(counter2[1]), .A1N(n966), .Y(
        n1113) );
  AOI21X1 U124 ( .A0(n1308), .A1(n1329), .B0(n1303), .Y(n965) );
  INVX1 U125 ( .A(n962), .Y(n1325) );
  AOI32X1 U126 ( .A0(reg_flag_mux), .A1(n1319), .A2(rst_n), .B0(n964), .B1(
        rst_n), .Y(n962) );
  NOR2X1 U127 ( .A(n973), .B(counter1[1]), .Y(n971) );
  NAND2X1 U128 ( .A(reg_datain_flag), .B(n1326), .Y(n973) );
  OAI221XL U129 ( .A0(n876), .A1(n1314), .B0(n842), .B1(n1300), .C0(n1011), 
        .Y(N65) );
  OAI221XL U130 ( .A0(n944), .A1(n1316), .B0(n910), .B1(n1297), .C0(n976), .Y(
        N99) );
  OAI221XL U131 ( .A0(n706), .A1(n1317), .B0(n740), .B1(n1298), .C0(n1079), 
        .Y(N133) );
  OAI221XL U132 ( .A0(n808), .A1(n1316), .B0(n774), .B1(n1301), .C0(n1045), 
        .Y(N167) );
  NAND2X1 U133 ( .A(counter2[1]), .B(n1328), .Y(n968) );
  NAND2X1 U134 ( .A(counter2[1]), .B(counter2[0]), .Y(n963) );
  OAI221XL U135 ( .A0(n858), .A1(n1313), .B0(n824), .B1(n1301), .C0(n993), .Y(
        N83) );
  AOI22X1 U136 ( .A0(R1[31]), .A1(n1312), .B0(n1276), .B1(R0[31]), .Y(n993) );
  OAI221XL U137 ( .A0(n926), .A1(n1319), .B0(n892), .B1(n1297), .C0(n1095), 
        .Y(N117) );
  AOI22X1 U138 ( .A0(R5[31]), .A1(n1312), .B0(n1270), .B1(R4[31]), .Y(n1095)
         );
  OAI221XL U139 ( .A0(n688), .A1(n1316), .B0(n722), .B1(n1297), .C0(n1061), 
        .Y(N151) );
  AOI22X1 U140 ( .A0(R9[31]), .A1(n1306), .B0(n1273), .B1(R8[31]), .Y(n1061)
         );
  OAI221XL U141 ( .A0(n790), .A1(n1315), .B0(n756), .B1(n1299), .C0(n1027), 
        .Y(N185) );
  AOI22X1 U142 ( .A0(R13[31]), .A1(n1309), .B0(n1275), .B1(R12[31]), .Y(n1027)
         );
  OAI221XL U143 ( .A0(n875), .A1(n1314), .B0(n841), .B1(n1300), .C0(n1010), 
        .Y(N66) );
  AOI22X1 U144 ( .A0(R1[14]), .A1(n1310), .B0(n1271), .B1(R0[14]), .Y(n1010)
         );
  OAI221XL U145 ( .A0(n874), .A1(n1314), .B0(n840), .B1(n1300), .C0(n1009), 
        .Y(N67) );
  AOI22X1 U146 ( .A0(R1[15]), .A1(n1310), .B0(n1276), .B1(R0[15]), .Y(n1009)
         );
  OAI221XL U147 ( .A0(n873), .A1(n1314), .B0(n839), .B1(n1300), .C0(n1008), 
        .Y(N68) );
  OAI221XL U148 ( .A0(n865), .A1(n1313), .B0(n831), .B1(n1301), .C0(n1000), 
        .Y(N76) );
  AOI22X1 U149 ( .A0(R1[24]), .A1(n1311), .B0(n1276), .B1(R0[24]), .Y(n1000)
         );
  OAI221XL U150 ( .A0(n859), .A1(n1313), .B0(n825), .B1(n1301), .C0(n994), .Y(
        N82) );
  AOI22X1 U151 ( .A0(R1[30]), .A1(n1312), .B0(n1276), .B1(R0[30]), .Y(n994) );
  OAI221XL U152 ( .A0(n857), .A1(n1313), .B0(n823), .B1(n1302), .C0(n992), .Y(
        N84) );
  AOI22X1 U153 ( .A0(R1[32]), .A1(n1312), .B0(n1277), .B1(R0[32]), .Y(n992) );
  OAI221XL U154 ( .A0(n856), .A1(n1313), .B0(n822), .B1(n1302), .C0(n991), .Y(
        N85) );
  AOI22X1 U155 ( .A0(R1[33]), .A1(n1312), .B0(n1277), .B1(R0[33]), .Y(n991) );
  OAI221XL U156 ( .A0(n943), .A1(n1319), .B0(n909), .B1(n1296), .C0(n1112), 
        .Y(N100) );
  AOI22X1 U157 ( .A0(R5[14]), .A1(n1304), .B0(n1272), .B1(R4[14]), .Y(n1112)
         );
  OAI221XL U158 ( .A0(n942), .A1(n1319), .B0(n908), .B1(n1296), .C0(n1111), 
        .Y(N101) );
  AOI22X1 U159 ( .A0(R5[15]), .A1(n1304), .B0(n1270), .B1(R4[15]), .Y(n1111)
         );
  OAI221XL U160 ( .A0(n941), .A1(n1319), .B0(n907), .B1(n1296), .C0(n1110), 
        .Y(N102) );
  OAI221XL U161 ( .A0(n933), .A1(n1319), .B0(n899), .B1(n1296), .C0(n1102), 
        .Y(N110) );
  AOI22X1 U162 ( .A0(R5[24]), .A1(n1304), .B0(n1273), .B1(R4[24]), .Y(n1102)
         );
  OAI221XL U163 ( .A0(n927), .A1(n1319), .B0(n893), .B1(n1297), .C0(n1096), 
        .Y(N116) );
  AOI22X1 U164 ( .A0(R5[30]), .A1(n1304), .B0(n1270), .B1(R4[30]), .Y(n1096)
         );
  OAI221XL U165 ( .A0(n925), .A1(n1319), .B0(n891), .B1(n1297), .C0(n1094), 
        .Y(N118) );
  AOI22X1 U166 ( .A0(R5[32]), .A1(n1312), .B0(n1270), .B1(R4[32]), .Y(n1094)
         );
  OAI221XL U167 ( .A0(n924), .A1(n1319), .B0(n890), .B1(n1297), .C0(n1093), 
        .Y(N119) );
  AOI22X1 U168 ( .A0(R5[33]), .A1(n1304), .B0(n1270), .B1(R4[33]), .Y(n1093)
         );
  OAI221XL U169 ( .A0(n705), .A1(n1317), .B0(n739), .B1(n1298), .C0(n1078), 
        .Y(N134) );
  AOI22X1 U170 ( .A0(R9[14]), .A1(n1305), .B0(n1271), .B1(R8[14]), .Y(n1078)
         );
  OAI221XL U171 ( .A0(n704), .A1(n1317), .B0(n738), .B1(n1298), .C0(n1077), 
        .Y(N135) );
  AOI22X1 U172 ( .A0(R9[15]), .A1(n1305), .B0(n1271), .B1(R8[15]), .Y(n1077)
         );
  OAI221XL U173 ( .A0(n703), .A1(n1317), .B0(n737), .B1(n968), .C0(n1076), .Y(
        N136) );
  OAI221XL U174 ( .A0(n695), .A1(n1317), .B0(n729), .B1(n1302), .C0(n1068), 
        .Y(N144) );
  AOI22X1 U175 ( .A0(R9[24]), .A1(n1306), .B0(n1272), .B1(R8[24]), .Y(n1068)
         );
  OAI221XL U176 ( .A0(n689), .A1(n1316), .B0(n723), .B1(n1301), .C0(n1062), 
        .Y(N150) );
  AOI22X1 U177 ( .A0(R9[30]), .A1(n1306), .B0(n1273), .B1(R8[30]), .Y(n1062)
         );
  OAI221XL U178 ( .A0(n687), .A1(n1316), .B0(n721), .B1(n1299), .C0(n1060), 
        .Y(N152) );
  AOI22X1 U179 ( .A0(R9[32]), .A1(n1307), .B0(n1273), .B1(R8[32]), .Y(n1060)
         );
  OAI221XL U180 ( .A0(n686), .A1(n1316), .B0(n720), .B1(n968), .C0(n1059), .Y(
        N153) );
  AOI22X1 U181 ( .A0(R9[33]), .A1(n1307), .B0(n1273), .B1(R8[33]), .Y(n1059)
         );
  OAI221XL U182 ( .A0(n807), .A1(n1317), .B0(n773), .B1(n1300), .C0(n1044), 
        .Y(N168) );
  AOI22X1 U183 ( .A0(R13[14]), .A1(n1308), .B0(n1270), .B1(R12[14]), .Y(n1044)
         );
  OAI221XL U184 ( .A0(n806), .A1(n1313), .B0(n772), .B1(n1299), .C0(n1043), 
        .Y(N169) );
  AOI22X1 U185 ( .A0(R13[15]), .A1(n1308), .B0(n1274), .B1(R12[15]), .Y(n1043)
         );
  OAI221XL U186 ( .A0(n805), .A1(n1314), .B0(n771), .B1(n1302), .C0(n1042), 
        .Y(N170) );
  OAI221XL U187 ( .A0(n797), .A1(n1316), .B0(n763), .B1(n1297), .C0(n1034), 
        .Y(N178) );
  AOI22X1 U188 ( .A0(R13[24]), .A1(n1309), .B0(n1274), .B1(R12[24]), .Y(n1034)
         );
  OAI221XL U189 ( .A0(n791), .A1(n1317), .B0(n757), .B1(n1299), .C0(n1028), 
        .Y(N184) );
  AOI22X1 U190 ( .A0(R13[30]), .A1(n1309), .B0(n1275), .B1(R12[30]), .Y(n1028)
         );
  OAI221XL U191 ( .A0(n789), .A1(n1315), .B0(n755), .B1(n1299), .C0(n1026), 
        .Y(N186) );
  AOI22X1 U192 ( .A0(R13[32]), .A1(n1309), .B0(n1275), .B1(R12[32]), .Y(n1026)
         );
  OAI221XL U193 ( .A0(n788), .A1(n1315), .B0(n754), .B1(n1299), .C0(n1025), 
        .Y(N187) );
  AOI22X1 U194 ( .A0(R13[33]), .A1(n1309), .B0(n1275), .B1(R12[33]), .Y(n1025)
         );
  OAI221XL U195 ( .A0(n889), .A1(n1315), .B0(n855), .B1(n1299), .C0(n1024), 
        .Y(N52) );
  AOI22X1 U196 ( .A0(R1[0]), .A1(n1309), .B0(n1275), .B1(R0[0]), .Y(n1024) );
  OAI221XL U197 ( .A0(n888), .A1(n1315), .B0(n854), .B1(n1299), .C0(n1023), 
        .Y(N53) );
  AOI22X1 U198 ( .A0(R1[1]), .A1(n1309), .B0(n1275), .B1(R0[1]), .Y(n1023) );
  OAI221XL U199 ( .A0(n887), .A1(n1315), .B0(n853), .B1(n1299), .C0(n1022), 
        .Y(N54) );
  AOI22X1 U200 ( .A0(R1[2]), .A1(n1309), .B0(n1275), .B1(R0[2]), .Y(n1022) );
  OAI221XL U201 ( .A0(n886), .A1(n1315), .B0(n852), .B1(n1299), .C0(n1021), 
        .Y(N55) );
  AOI22X1 U202 ( .A0(R1[3]), .A1(n1310), .B0(n1275), .B1(R0[3]), .Y(n1021) );
  OAI221XL U203 ( .A0(n885), .A1(n1315), .B0(n851), .B1(n1299), .C0(n1020), 
        .Y(N56) );
  AOI22X1 U204 ( .A0(R1[4]), .A1(n1310), .B0(n1275), .B1(R0[4]), .Y(n1020) );
  OAI221XL U205 ( .A0(n884), .A1(n1315), .B0(n850), .B1(n1299), .C0(n1019), 
        .Y(N57) );
  AOI22X1 U206 ( .A0(R1[5]), .A1(n1310), .B0(n1275), .B1(R0[5]), .Y(n1019) );
  OAI221XL U207 ( .A0(n883), .A1(n1315), .B0(n849), .B1(n1299), .C0(n1018), 
        .Y(N58) );
  AOI22X1 U208 ( .A0(R1[6]), .A1(n1310), .B0(n1275), .B1(R0[6]), .Y(n1018) );
  OAI221XL U209 ( .A0(n882), .A1(n1315), .B0(n848), .B1(n1299), .C0(n1017), 
        .Y(N59) );
  AOI22X1 U210 ( .A0(R1[7]), .A1(n1310), .B0(n1275), .B1(R0[7]), .Y(n1017) );
  OAI221XL U211 ( .A0(n881), .A1(n1315), .B0(n847), .B1(n1300), .C0(n1016), 
        .Y(N60) );
  AOI22X1 U212 ( .A0(R1[8]), .A1(n1310), .B0(n1274), .B1(R0[8]), .Y(n1016) );
  OAI221XL U213 ( .A0(n880), .A1(n1315), .B0(n846), .B1(n1300), .C0(n1015), 
        .Y(N61) );
  AOI22X1 U214 ( .A0(R1[9]), .A1(n1310), .B0(n1271), .B1(R0[9]), .Y(n1015) );
  OAI221XL U215 ( .A0(n879), .A1(n1314), .B0(n845), .B1(n1300), .C0(n1014), 
        .Y(N62) );
  AOI22X1 U216 ( .A0(R1[10]), .A1(n1310), .B0(n1276), .B1(R0[10]), .Y(n1014)
         );
  OAI221XL U217 ( .A0(n878), .A1(n1314), .B0(n844), .B1(n1300), .C0(n1013), 
        .Y(N63) );
  AOI22X1 U218 ( .A0(R1[11]), .A1(n1310), .B0(n1272), .B1(R0[11]), .Y(n1013)
         );
  OAI221XL U219 ( .A0(n877), .A1(n1314), .B0(n843), .B1(n1300), .C0(n1012), 
        .Y(N64) );
  AOI22X1 U220 ( .A0(R1[12]), .A1(n1310), .B0(n1272), .B1(R0[12]), .Y(n1012)
         );
  OAI221XL U221 ( .A0(n872), .A1(n1314), .B0(n838), .B1(n1300), .C0(n1007), 
        .Y(N69) );
  AOI22X1 U222 ( .A0(R1[17]), .A1(n1311), .B0(n1270), .B1(R0[17]), .Y(n1007)
         );
  OAI221XL U223 ( .A0(n871), .A1(n1314), .B0(n837), .B1(n1300), .C0(n1006), 
        .Y(N70) );
  AOI22X1 U224 ( .A0(R1[18]), .A1(n1311), .B0(n1273), .B1(R0[18]), .Y(n1006)
         );
  OAI221XL U225 ( .A0(n870), .A1(n1314), .B0(n836), .B1(n1300), .C0(n1005), 
        .Y(N71) );
  AOI22X1 U226 ( .A0(R1[19]), .A1(n1311), .B0(n1277), .B1(R0[19]), .Y(n1005)
         );
  OAI221XL U227 ( .A0(n869), .A1(n1314), .B0(n835), .B1(n1301), .C0(n1004), 
        .Y(N72) );
  AOI22X1 U228 ( .A0(R1[20]), .A1(n1311), .B0(n1276), .B1(R0[20]), .Y(n1004)
         );
  OAI221XL U229 ( .A0(n868), .A1(n1314), .B0(n834), .B1(n1301), .C0(n1003), 
        .Y(N73) );
  AOI22X1 U230 ( .A0(R1[21]), .A1(n1311), .B0(n1276), .B1(R0[21]), .Y(n1003)
         );
  OAI221XL U231 ( .A0(n867), .A1(n1314), .B0(n833), .B1(n1301), .C0(n1002), 
        .Y(N74) );
  AOI22X1 U232 ( .A0(R1[22]), .A1(n1311), .B0(n1276), .B1(R0[22]), .Y(n1002)
         );
  OAI221XL U233 ( .A0(n866), .A1(n1313), .B0(n832), .B1(n1301), .C0(n1001), 
        .Y(N75) );
  AOI22X1 U234 ( .A0(R1[23]), .A1(n1311), .B0(n1276), .B1(R0[23]), .Y(n1001)
         );
  OAI221XL U235 ( .A0(n864), .A1(n1313), .B0(n830), .B1(n1301), .C0(n999), .Y(
        N77) );
  AOI22X1 U236 ( .A0(R1[25]), .A1(n1311), .B0(n1276), .B1(R0[25]), .Y(n999) );
  OAI221XL U237 ( .A0(n863), .A1(n1313), .B0(n829), .B1(n1301), .C0(n998), .Y(
        N78) );
  AOI22X1 U238 ( .A0(R1[26]), .A1(n1311), .B0(n1276), .B1(R0[26]), .Y(n998) );
  OAI221XL U239 ( .A0(n862), .A1(n1313), .B0(n828), .B1(n1301), .C0(n997), .Y(
        N79) );
  AOI22X1 U240 ( .A0(R1[27]), .A1(n1311), .B0(n1276), .B1(R0[27]), .Y(n997) );
  OAI221XL U241 ( .A0(n861), .A1(n1313), .B0(n827), .B1(n1301), .C0(n996), .Y(
        N80) );
  AOI22X1 U242 ( .A0(R1[28]), .A1(n1311), .B0(n1276), .B1(R0[28]), .Y(n996) );
  OAI221XL U243 ( .A0(n860), .A1(n1313), .B0(n826), .B1(n1301), .C0(n995), .Y(
        N81) );
  AOI22X1 U244 ( .A0(R1[29]), .A1(n1312), .B0(n1276), .B1(R0[29]), .Y(n995) );
  OAI221XL U245 ( .A0(n957), .A1(n1313), .B0(n923), .B1(n1302), .C0(n990), .Y(
        N86) );
  AOI22X1 U246 ( .A0(R5[0]), .A1(n1312), .B0(n1277), .B1(R4[0]), .Y(n990) );
  OAI221XL U247 ( .A0(n956), .A1(n1313), .B0(n922), .B1(n1302), .C0(n989), .Y(
        N87) );
  AOI22X1 U248 ( .A0(R5[1]), .A1(n1312), .B0(n1277), .B1(R4[1]), .Y(n989) );
  OAI221XL U249 ( .A0(n955), .A1(n1313), .B0(n921), .B1(n1302), .C0(n988), .Y(
        N88) );
  AOI22X1 U250 ( .A0(R5[2]), .A1(n1312), .B0(n1277), .B1(R4[2]), .Y(n988) );
  OAI221XL U251 ( .A0(n954), .A1(n1315), .B0(n920), .B1(n1302), .C0(n987), .Y(
        N89) );
  AOI22X1 U252 ( .A0(R5[3]), .A1(n1312), .B0(n1277), .B1(R4[3]), .Y(n987) );
  OAI221XL U253 ( .A0(n953), .A1(n1314), .B0(n919), .B1(n1302), .C0(n986), .Y(
        N90) );
  AOI22X1 U254 ( .A0(R5[4]), .A1(n1312), .B0(n1277), .B1(R4[4]), .Y(n986) );
  OAI221XL U255 ( .A0(n952), .A1(n1318), .B0(n918), .B1(n1302), .C0(n985), .Y(
        N91) );
  AOI22X1 U256 ( .A0(R5[5]), .A1(n1312), .B0(n1277), .B1(R4[5]), .Y(n985) );
  OAI221XL U257 ( .A0(n951), .A1(n963), .B0(n917), .B1(n1302), .C0(n984), .Y(
        N92) );
  AOI22X1 U258 ( .A0(R5[6]), .A1(n1312), .B0(n1277), .B1(R4[6]), .Y(n984) );
  OAI221XL U259 ( .A0(n950), .A1(n963), .B0(n916), .B1(n1302), .C0(n983), .Y(
        N93) );
  AOI22X1 U260 ( .A0(R5[7]), .A1(n1312), .B0(n1277), .B1(R4[7]), .Y(n983) );
  OAI221XL U261 ( .A0(n949), .A1(n963), .B0(n915), .B1(n1302), .C0(n982), .Y(
        N94) );
  AOI22X1 U262 ( .A0(R5[8]), .A1(n1305), .B0(n1277), .B1(R4[8]), .Y(n982) );
  OAI221XL U263 ( .A0(n948), .A1(n963), .B0(n914), .B1(n1302), .C0(n981), .Y(
        N95) );
  AOI22X1 U264 ( .A0(R5[9]), .A1(n1307), .B0(n1277), .B1(R4[9]), .Y(n981) );
  OAI221XL U265 ( .A0(n947), .A1(n963), .B0(n913), .B1(n1301), .C0(n980), .Y(
        N96) );
  AOI22X1 U266 ( .A0(R5[10]), .A1(n1311), .B0(n1277), .B1(R4[10]), .Y(n980) );
  OAI221XL U267 ( .A0(n946), .A1(n963), .B0(n912), .B1(n1297), .C0(n979), .Y(
        N97) );
  AOI22X1 U268 ( .A0(R5[11]), .A1(n1310), .B0(n1277), .B1(R4[11]), .Y(n979) );
  OAI221XL U269 ( .A0(n945), .A1(n963), .B0(n911), .B1(n1301), .C0(n978), .Y(
        N98) );
  AOI22X1 U270 ( .A0(R5[12]), .A1(n1306), .B0(n1276), .B1(R4[12]), .Y(n978) );
  OAI221XL U271 ( .A0(n940), .A1(n1317), .B0(n906), .B1(n1296), .C0(n1109), 
        .Y(N103) );
  AOI22X1 U272 ( .A0(R5[17]), .A1(n1304), .B0(n1274), .B1(R4[17]), .Y(n1109)
         );
  OAI221XL U273 ( .A0(n939), .A1(n963), .B0(n905), .B1(n1296), .C0(n1108), .Y(
        N104) );
  AOI22X1 U274 ( .A0(R5[18]), .A1(n1304), .B0(n1272), .B1(R4[18]), .Y(n1108)
         );
  OAI221XL U275 ( .A0(n938), .A1(n963), .B0(n904), .B1(n1296), .C0(n1107), .Y(
        N105) );
  AOI22X1 U276 ( .A0(R5[19]), .A1(n1304), .B0(n1273), .B1(R4[19]), .Y(n1107)
         );
  OAI221XL U277 ( .A0(n937), .A1(n963), .B0(n903), .B1(n1296), .C0(n1106), .Y(
        N106) );
  AOI22X1 U278 ( .A0(R5[20]), .A1(n1304), .B0(n1275), .B1(R4[20]), .Y(n1106)
         );
  OAI221XL U279 ( .A0(n936), .A1(n1319), .B0(n902), .B1(n1296), .C0(n1105), 
        .Y(N107) );
  AOI22X1 U280 ( .A0(R5[21]), .A1(n1304), .B0(n1275), .B1(R4[21]), .Y(n1105)
         );
  OAI221XL U281 ( .A0(n935), .A1(n1319), .B0(n901), .B1(n1296), .C0(n1104), 
        .Y(N108) );
  AOI22X1 U282 ( .A0(R5[22]), .A1(n1304), .B0(n1271), .B1(R4[22]), .Y(n1104)
         );
  OAI221XL U283 ( .A0(n934), .A1(n1319), .B0(n900), .B1(n1296), .C0(n1103), 
        .Y(N109) );
  AOI22X1 U284 ( .A0(R5[23]), .A1(n1304), .B0(n1270), .B1(R4[23]), .Y(n1103)
         );
  OAI221XL U285 ( .A0(n932), .A1(n1319), .B0(n898), .B1(n1296), .C0(n1101), 
        .Y(N111) );
  AOI22X1 U286 ( .A0(R5[25]), .A1(n1304), .B0(n1270), .B1(R4[25]), .Y(n1101)
         );
  OAI221XL U287 ( .A0(n931), .A1(n1319), .B0(n897), .B1(n1297), .C0(n1100), 
        .Y(N112) );
  AOI22X1 U288 ( .A0(R5[26]), .A1(n1304), .B0(n1270), .B1(R4[26]), .Y(n1100)
         );
  OAI221XL U289 ( .A0(n930), .A1(n1319), .B0(n896), .B1(n1297), .C0(n1099), 
        .Y(N113) );
  AOI22X1 U290 ( .A0(R5[27]), .A1(n1304), .B0(n1270), .B1(R4[27]), .Y(n1099)
         );
  OAI221XL U291 ( .A0(n929), .A1(n1319), .B0(n895), .B1(n1297), .C0(n1098), 
        .Y(N114) );
  AOI22X1 U292 ( .A0(R5[28]), .A1(n1308), .B0(n1270), .B1(R4[28]), .Y(n1098)
         );
  OAI221XL U293 ( .A0(n928), .A1(n1319), .B0(n894), .B1(n1297), .C0(n1097), 
        .Y(N115) );
  AOI22X1 U294 ( .A0(R5[29]), .A1(n1305), .B0(n1270), .B1(R4[29]), .Y(n1097)
         );
  OAI221XL U295 ( .A0(n719), .A1(n1318), .B0(n753), .B1(n1297), .C0(n1092), 
        .Y(N120) );
  AOI22X1 U296 ( .A0(R9[0]), .A1(n1307), .B0(n1270), .B1(R8[0]), .Y(n1092) );
  OAI221XL U297 ( .A0(n718), .A1(n1318), .B0(n752), .B1(n1297), .C0(n1091), 
        .Y(N121) );
  AOI22X1 U298 ( .A0(R9[1]), .A1(n1311), .B0(n1270), .B1(R8[1]), .Y(n1091) );
  OAI221XL U299 ( .A0(n717), .A1(n1318), .B0(n751), .B1(n1297), .C0(n1090), 
        .Y(N122) );
  AOI22X1 U300 ( .A0(R9[2]), .A1(n1310), .B0(n1270), .B1(R8[2]), .Y(n1090) );
  OAI221XL U301 ( .A0(n716), .A1(n1318), .B0(n750), .B1(n1297), .C0(n1089), 
        .Y(N123) );
  AOI22X1 U303 ( .A0(R9[3]), .A1(n1309), .B0(n1270), .B1(R8[3]), .Y(n1089) );
  OAI221XL U304 ( .A0(n715), .A1(n1318), .B0(n749), .B1(n1298), .C0(n1088), 
        .Y(N124) );
  AOI22X1 U305 ( .A0(R9[4]), .A1(n1306), .B0(n1271), .B1(R8[4]), .Y(n1088) );
  OAI221XL U306 ( .A0(n714), .A1(n1318), .B0(n748), .B1(n1298), .C0(n1087), 
        .Y(N125) );
  AOI22X1 U307 ( .A0(R9[5]), .A1(n1312), .B0(n1271), .B1(R8[5]), .Y(n1087) );
  OAI221XL U308 ( .A0(n713), .A1(n1318), .B0(n747), .B1(n1298), .C0(n1086), 
        .Y(N126) );
  AOI22X1 U309 ( .A0(R9[6]), .A1(n1305), .B0(n1271), .B1(R8[6]), .Y(n1086) );
  OAI221XL U310 ( .A0(n712), .A1(n1318), .B0(n746), .B1(n1298), .C0(n1085), 
        .Y(N127) );
  AOI22X1 U311 ( .A0(R9[7]), .A1(n1305), .B0(n1271), .B1(R8[7]), .Y(n1085) );
  OAI221XL U312 ( .A0(n711), .A1(n1318), .B0(n745), .B1(n1298), .C0(n1084), 
        .Y(N128) );
  AOI22X1 U313 ( .A0(R9[8]), .A1(n1305), .B0(n1271), .B1(R8[8]), .Y(n1084) );
  OAI221XL U314 ( .A0(n710), .A1(n1318), .B0(n744), .B1(n1298), .C0(n1083), 
        .Y(N129) );
  AOI22X1 U315 ( .A0(R9[9]), .A1(n1305), .B0(n1271), .B1(R8[9]), .Y(n1083) );
  OAI221XL U316 ( .A0(n709), .A1(n1318), .B0(n743), .B1(n1298), .C0(n1082), 
        .Y(N130) );
  AOI22X1 U317 ( .A0(R9[10]), .A1(n1305), .B0(n1271), .B1(R8[10]), .Y(n1082)
         );
  OAI221XL U318 ( .A0(n708), .A1(n1318), .B0(n742), .B1(n1298), .C0(n1081), 
        .Y(N131) );
  AOI22X1 U319 ( .A0(R9[11]), .A1(n1305), .B0(n1271), .B1(R8[11]), .Y(n1081)
         );
  OAI221XL U320 ( .A0(n707), .A1(n1318), .B0(n741), .B1(n1298), .C0(n1080), 
        .Y(N132) );
  AOI22X1 U321 ( .A0(R9[12]), .A1(n1305), .B0(n1271), .B1(R8[12]), .Y(n1080)
         );
  OAI221XL U322 ( .A0(n702), .A1(n1317), .B0(n736), .B1(n1298), .C0(n1075), 
        .Y(N137) );
  AOI22X1 U323 ( .A0(R9[17]), .A1(n1305), .B0(n1272), .B1(R8[17]), .Y(n1075)
         );
  OAI221XL U324 ( .A0(n701), .A1(n1317), .B0(n735), .B1(n1296), .C0(n1074), 
        .Y(N138) );
  AOI22X1 U325 ( .A0(R9[18]), .A1(n1305), .B0(n1272), .B1(R8[18]), .Y(n1074)
         );
  OAI221XL U326 ( .A0(n700), .A1(n1317), .B0(n734), .B1(n968), .C0(n1073), .Y(
        N139) );
  AOI22X1 U327 ( .A0(R9[19]), .A1(n1306), .B0(n1272), .B1(R8[19]), .Y(n1073)
         );
  OAI221XL U328 ( .A0(n699), .A1(n1317), .B0(n733), .B1(n968), .C0(n1072), .Y(
        N140) );
  AOI22X1 U329 ( .A0(R9[20]), .A1(n1306), .B0(n1272), .B1(R8[20]), .Y(n1072)
         );
  OAI221XL U330 ( .A0(n698), .A1(n1317), .B0(n732), .B1(n968), .C0(n1071), .Y(
        N141) );
  AOI22X1 U331 ( .A0(R9[21]), .A1(n1306), .B0(n1272), .B1(R8[21]), .Y(n1071)
         );
  OAI221XL U332 ( .A0(n697), .A1(n1317), .B0(n731), .B1(n968), .C0(n1070), .Y(
        N142) );
  AOI22X1 U333 ( .A0(R9[22]), .A1(n1306), .B0(n1272), .B1(R8[22]), .Y(n1070)
         );
  OAI221XL U334 ( .A0(n696), .A1(n1317), .B0(n730), .B1(n968), .C0(n1069), .Y(
        N143) );
  AOI22X1 U335 ( .A0(R9[23]), .A1(n1306), .B0(n1272), .B1(R8[23]), .Y(n1069)
         );
  OAI221XL U336 ( .A0(n694), .A1(n1317), .B0(n728), .B1(n968), .C0(n1067), .Y(
        N145) );
  AOI22X1 U337 ( .A0(R9[25]), .A1(n1306), .B0(n1272), .B1(R8[25]), .Y(n1067)
         );
  OAI221XL U338 ( .A0(n693), .A1(n1316), .B0(n727), .B1(n968), .C0(n1066), .Y(
        N146) );
  AOI22X1 U339 ( .A0(R9[26]), .A1(n1306), .B0(n1272), .B1(R8[26]), .Y(n1066)
         );
  OAI221XL U340 ( .A0(n692), .A1(n1316), .B0(n726), .B1(n968), .C0(n1065), .Y(
        N147) );
  AOI22X1 U341 ( .A0(R9[27]), .A1(n1306), .B0(n1272), .B1(R8[27]), .Y(n1065)
         );
  OAI221XL U342 ( .A0(n691), .A1(n1316), .B0(n725), .B1(n1297), .C0(n1064), 
        .Y(N148) );
  AOI22X1 U343 ( .A0(R9[28]), .A1(n1306), .B0(n1273), .B1(R8[28]), .Y(n1064)
         );
  OAI221XL U344 ( .A0(n690), .A1(n1316), .B0(n724), .B1(n1301), .C0(n1063), 
        .Y(N149) );
  AOI22X1 U345 ( .A0(R9[29]), .A1(n1306), .B0(n1273), .B1(R8[29]), .Y(n1063)
         );
  OAI221XL U346 ( .A0(n821), .A1(n1316), .B0(n787), .B1(n1300), .C0(n1058), 
        .Y(N154) );
  AOI22X1 U347 ( .A0(R13[0]), .A1(n1307), .B0(n1273), .B1(R12[0]), .Y(n1058)
         );
  OAI221XL U348 ( .A0(n820), .A1(n1316), .B0(n786), .B1(n1300), .C0(n1057), 
        .Y(N155) );
  AOI22X1 U349 ( .A0(R13[1]), .A1(n1307), .B0(n1273), .B1(R12[1]), .Y(n1057)
         );
  OAI221XL U350 ( .A0(n819), .A1(n1316), .B0(n785), .B1(n1299), .C0(n1056), 
        .Y(N156) );
  AOI22X1 U351 ( .A0(R13[2]), .A1(n1307), .B0(n1273), .B1(R12[2]), .Y(n1056)
         );
  OAI221XL U352 ( .A0(n818), .A1(n1316), .B0(n784), .B1(n1298), .C0(n1055), 
        .Y(N157) );
  AOI22X1 U353 ( .A0(R13[3]), .A1(n1307), .B0(n1273), .B1(R12[3]), .Y(n1055)
         );
  OAI221XL U354 ( .A0(n817), .A1(n1316), .B0(n783), .B1(n1302), .C0(n1054), 
        .Y(N158) );
  AOI22X1 U355 ( .A0(R13[4]), .A1(n1307), .B0(n1273), .B1(R12[4]), .Y(n1054)
         );
  OAI221XL U356 ( .A0(n816), .A1(n1318), .B0(n782), .B1(n1296), .C0(n1053), 
        .Y(N159) );
  AOI22X1 U357 ( .A0(R13[5]), .A1(n1307), .B0(n1273), .B1(R12[5]), .Y(n1053)
         );
  OAI221XL U358 ( .A0(n815), .A1(n1315), .B0(n781), .B1(n1298), .C0(n1052), 
        .Y(N160) );
  AOI22X1 U359 ( .A0(R13[6]), .A1(n1307), .B0(n1273), .B1(R12[6]), .Y(n1052)
         );
  OAI221XL U360 ( .A0(n814), .A1(n1319), .B0(n780), .B1(n1296), .C0(n1051), 
        .Y(N161) );
  AOI22X1 U361 ( .A0(R13[7]), .A1(n1307), .B0(n1276), .B1(R12[7]), .Y(n1051)
         );
  OAI221XL U362 ( .A0(n813), .A1(n1316), .B0(n779), .B1(n968), .C0(n1050), .Y(
        N162) );
  AOI22X1 U363 ( .A0(R13[8]), .A1(n1307), .B0(n1277), .B1(R12[8]), .Y(n1050)
         );
  OAI221XL U364 ( .A0(n812), .A1(n1317), .B0(n778), .B1(n968), .C0(n1049), .Y(
        N163) );
  AOI22X1 U365 ( .A0(R13[9]), .A1(n1307), .B0(n1275), .B1(R12[9]), .Y(n1049)
         );
  OAI221XL U366 ( .A0(n811), .A1(n1313), .B0(n777), .B1(n968), .C0(n1048), .Y(
        N164) );
  AOI22X1 U367 ( .A0(R13[10]), .A1(n1307), .B0(n1276), .B1(R12[10]), .Y(n1048)
         );
  OAI221XL U368 ( .A0(n810), .A1(n1314), .B0(n776), .B1(n968), .C0(n1047), .Y(
        N165) );
  AOI22X1 U369 ( .A0(R13[11]), .A1(n1308), .B0(n1272), .B1(R12[11]), .Y(n1047)
         );
  OAI221XL U370 ( .A0(n809), .A1(n1318), .B0(n775), .B1(n968), .C0(n1046), .Y(
        N166) );
  AOI22X1 U371 ( .A0(R13[12]), .A1(n1308), .B0(n1273), .B1(R12[12]), .Y(n1046)
         );
  OAI221XL U372 ( .A0(n804), .A1(n1315), .B0(n770), .B1(n968), .C0(n1041), .Y(
        N171) );
  AOI22X1 U373 ( .A0(R13[17]), .A1(n1308), .B0(n1277), .B1(R12[17]), .Y(n1041)
         );
  OAI221XL U374 ( .A0(n803), .A1(n1313), .B0(n769), .B1(n1300), .C0(n1040), 
        .Y(N172) );
  AOI22X1 U375 ( .A0(R13[18]), .A1(n1308), .B0(n1274), .B1(R12[18]), .Y(n1040)
         );
  OAI221XL U376 ( .A0(n802), .A1(n1315), .B0(n768), .B1(n1299), .C0(n1039), 
        .Y(N173) );
  AOI22X1 U377 ( .A0(R13[19]), .A1(n1308), .B0(n1274), .B1(R12[19]), .Y(n1039)
         );
  OAI221XL U378 ( .A0(n801), .A1(n1314), .B0(n767), .B1(n1298), .C0(n1038), 
        .Y(N174) );
  AOI22X1 U379 ( .A0(R13[20]), .A1(n1308), .B0(n1274), .B1(R12[20]), .Y(n1038)
         );
  OAI221XL U380 ( .A0(n800), .A1(n1318), .B0(n766), .B1(n1302), .C0(n1037), 
        .Y(N175) );
  AOI22X1 U381 ( .A0(R13[21]), .A1(n1308), .B0(n1274), .B1(R12[21]), .Y(n1037)
         );
  OAI221XL U382 ( .A0(n799), .A1(n963), .B0(n765), .B1(n1296), .C0(n1036), .Y(
        N176) );
  AOI22X1 U383 ( .A0(R13[22]), .A1(n1308), .B0(n1274), .B1(R12[22]), .Y(n1036)
         );
  OAI221XL U384 ( .A0(n798), .A1(n963), .B0(n764), .B1(n968), .C0(n1035), .Y(
        N177) );
  AOI22X1 U385 ( .A0(R13[23]), .A1(n1308), .B0(n1274), .B1(R12[23]), .Y(n1035)
         );
  OAI221XL U386 ( .A0(n796), .A1(n963), .B0(n762), .B1(n1300), .C0(n1033), .Y(
        N179) );
  AOI22X1 U387 ( .A0(R13[25]), .A1(n1309), .B0(n1274), .B1(R12[25]), .Y(n1033)
         );
  OAI221XL U388 ( .A0(n795), .A1(n963), .B0(n761), .B1(n1299), .C0(n1032), .Y(
        N180) );
  AOI22X1 U389 ( .A0(R13[26]), .A1(n1309), .B0(n1274), .B1(R12[26]), .Y(n1032)
         );
  OAI221XL U390 ( .A0(n794), .A1(n963), .B0(n760), .B1(n1298), .C0(n1031), .Y(
        N181) );
  AOI22X1 U391 ( .A0(R13[27]), .A1(n1309), .B0(n1274), .B1(R12[27]), .Y(n1031)
         );
  OAI221XL U392 ( .A0(n793), .A1(n963), .B0(n759), .B1(n1302), .C0(n1030), .Y(
        N182) );
  AOI22X1 U393 ( .A0(R13[28]), .A1(n1309), .B0(n1274), .B1(R12[28]), .Y(n1030)
         );
  OAI221XL U394 ( .A0(n792), .A1(n963), .B0(n758), .B1(n1296), .C0(n1029), .Y(
        N183) );
  AOI22X1 U395 ( .A0(R13[29]), .A1(n1309), .B0(n1274), .B1(R12[29]), .Y(n1029)
         );
  AND2X2 U396 ( .A(reg_datain_flag), .B(n964), .Y(n114) );
  INVX1 U397 ( .A(counter1[1]), .Y(n1327) );
  INVX1 U398 ( .A(counter2[0]), .Y(n1328) );
  AND3X2 U399 ( .A(counter1[0]), .B(n1327), .C(reg_datain_flag), .Y(n115) );
  INVX1 U400 ( .A(reg_flag_mux), .Y(n1324) );
  AOI22X1 U401 ( .A0(R9[13]), .A1(n1305), .B0(n1271), .B1(R8[13]), .Y(n1079)
         );
  AOI22X1 U402 ( .A0(R13[13]), .A1(n1308), .B0(n1275), .B1(R12[13]), .Y(n1045)
         );
  AOI22X1 U403 ( .A0(R1[13]), .A1(n1310), .B0(n1275), .B1(R0[13]), .Y(n1011)
         );
  AOI22X1 U404 ( .A0(R5[13]), .A1(n1309), .B0(n1271), .B1(R4[13]), .Y(n976) );
  AOI22X1 U405 ( .A0(R9[16]), .A1(n1305), .B0(n1272), .B1(R8[16]), .Y(n1076)
         );
  AOI22X1 U406 ( .A0(R13[16]), .A1(n1308), .B0(n1271), .B1(R12[16]), .Y(n1042)
         );
  AOI22X1 U407 ( .A0(R1[16]), .A1(n1311), .B0(n1274), .B1(R0[16]), .Y(n1008)
         );
  AOI22X1 U408 ( .A0(R5[16]), .A1(n1304), .B0(n1274), .B1(R4[16]), .Y(n1110)
         );
endmodule


module p_s ( clk, rst_n, data_in_3, p_s_flag_in, data_out_3 );
  input [135:0] data_in_3;
  output [33:0] data_out_3;
  input clk, rst_n, p_s_flag_in;
  wire   N26, N50, N52, N119, N120, N121, N122, N123, N124, N125, N126, N127,
         N128, N129, N130, N131, N132, N133, N134, N135, N136, N137, N138,
         N139, N140, N141, N142, N143, N144, N145, N146, N147, N148, N149,
         N150, N151, N152, n85, n86, n87, n96, n102, n104, n105, n115, n117,
         n118, n120, n121, n122, n134, n137, n138, n139, n221, n222, n223,
         n232, n238, n240, n241, n251, n253, n254, n256, n257, n258, n270,
         n273, n274, n275, n357, n358, n359, n368, n374, n375, n376, n377,
         n387, n389, n390, n391, n392, n393, n394, n406, n409, n410, n411,
         n425, n426, n427, n436, n442, n443, n444, n445, n523, n525, n527,
         n528, n529, n530, n542, n545, n546, n547, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n861, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n882, n883, n884,
         n886, n887, n888, n889, n892, n894, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
         n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
         n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
         n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
         n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
         n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
         n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
         n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
         n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
         n1160, n1161, n1162, n1163, n1164, n8, n9, n10, n19, n20, n21, n22,
         n23, n24, n25, n26, n71, n81, n82, n83, n98, n151, n152, n153, n511,
         n513, n515, n517, n519, n521, n524, n531, n533, n535, n537, n539,
         n541, n544, n549, n551, n553, n555, n557, n559, n561, n563, n565,
         n567, n569, n571, n573, n575, n577, n579, n581, n857, n859, n862,
         n864, n866, n881, n890, n893, n1165, n1167, n1169, n1171, n1173,
         n1175, n1177, n1179, n1181, n1183, n1185, n1187, n1189, n1191, n1193,
         n1195, n1197, n1199, n1201, n1203, n1205, n1207, n1209, n1211, n1213,
         n1215, n1217, n1219, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
         n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
         n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
         n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1305,
         n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
         n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
         n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
         n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
         n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
         n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
         n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
         n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
         n1386, n1387, n1388, n1389, n1390, n1391;
  wire   [1:0] counter_1;
  wire   [33:0] R0;
  wire   [33:0] R12;
  wire   [33:0] R1;
  wire   [33:0] R13;
  wire   [33:0] R2;
  wire   [33:0] R14;
  wire   [33:0] R3;
  wire   [33:0] R15;
  wire   [3:0] counter_2;

  AND2X2 U321 ( .A(n1157), .B(n869), .Y(n886) );
  AND2X2 U324 ( .A(counter_2[3]), .B(n861), .Y(n1157) );
  AND2X2 U326 ( .A(counter_2[3]), .B(counter_2[0]), .Y(n1158) );
  EDFFXL R8_reg_31_ ( .D(data_in_3[99]), .E(n1357), .CK(clk), .QN(n757) );
  EDFFXL R9_reg_31_ ( .D(data_in_3[99]), .E(n1368), .CK(clk), .QN(n825) );
  EDFFXL R4_reg_13_ ( .D(data_in_3[47]), .E(n1358), .CK(clk), .QN(n741) );
  EDFFXL R5_reg_13_ ( .D(data_in_3[47]), .E(n1369), .CK(clk), .QN(n809) );
  EDFFXL R1_reg_16_ ( .D(data_in_3[16]), .E(n1372), .CK(clk), .Q(R1[16]) );
  EDFFXL R0_reg_16_ ( .D(data_in_3[16]), .E(n1361), .CK(clk), .Q(R0[16]) );
  EDFFXL R3_reg_16_ ( .D(data_in_3[16]), .E(n1346), .CK(clk), .Q(R3[16]) );
  EDFFXL R2_reg_16_ ( .D(data_in_3[16]), .E(n1374), .CK(clk), .Q(R2[16]) );
  DFFXL R11_reg_14_ ( .D(n1296), .CK(clk), .Q(n358), .QN(n706) );
  DFFXL R10_reg_14_ ( .D(n1295), .CK(clk), .Q(n426), .QN(n638) );
  DFFXL R9_reg_14_ ( .D(n1294), .CK(clk), .Q(n86), .QN(n842) );
  DFFXL R8_reg_14_ ( .D(n1293), .CK(clk), .Q(n222), .QN(n774) );
  MX2X1 R11_reg_15__U3 ( .A(n359), .B(data_in_3[83]), .S0(n1343), .Y(n1292) );
  DFFXL R11_reg_15_ ( .D(n1292), .CK(clk), .Q(n359), .QN(n705) );
  MX2X1 R10_reg_15__U3 ( .A(n427), .B(data_in_3[83]), .S0(n1379), .Y(n1291) );
  DFFXL R10_reg_15_ ( .D(n1291), .CK(clk), .Q(n427), .QN(n637) );
  MX2X1 R9_reg_15__U3 ( .A(n87), .B(data_in_3[83]), .S0(n1367), .Y(n1290) );
  DFFXL R9_reg_15_ ( .D(n1290), .CK(clk), .Q(n87), .QN(n841) );
  MX2X1 R8_reg_15__U3 ( .A(n223), .B(data_in_3[83]), .S0(n1356), .Y(n1289) );
  DFFXL R8_reg_15_ ( .D(n1289), .CK(clk), .Q(n223), .QN(n773) );
  MX2X1 R11_reg_16__U3 ( .A(n1306), .B(data_in_3[84]), .S0(n1343), .Y(n1288)
         );
  DFFXL R11_reg_16_ ( .D(n1288), .CK(clk), .Q(n1306), .QN(n704) );
  MX2X1 R10_reg_16__U3 ( .A(n1305), .B(data_in_3[84]), .S0(n1379), .Y(n1287)
         );
  DFFXL R10_reg_16_ ( .D(n1287), .CK(clk), .Q(n1305), .QN(n636) );
  MX2X1 R9_reg_16__U3 ( .A(n1308), .B(data_in_3[84]), .S0(n1367), .Y(n1286) );
  DFFXL R9_reg_16_ ( .D(n1286), .CK(clk), .Q(n1308), .QN(n840) );
  MX2X1 R8_reg_16__U3 ( .A(n1307), .B(data_in_3[84]), .S0(n1356), .Y(n1285) );
  DFFXL R8_reg_16_ ( .D(n1285), .CK(clk), .Q(n1307), .QN(n772) );
  MX2X1 R7_reg_28__U3 ( .A(n542), .B(data_in_3[62]), .S0(n1341), .Y(n1284) );
  DFFXL R7_reg_28_ ( .D(n1284), .CK(clk), .Q(n542), .QN(n590) );
  MX2X1 R6_reg_28__U3 ( .A(n406), .B(data_in_3[62]), .S0(n1377), .Y(n1283) );
  DFFXL R6_reg_28_ ( .D(n1283), .CK(clk), .Q(n406), .QN(n658) );
  MX2X1 R5_reg_28__U3 ( .A(n134), .B(data_in_3[62]), .S0(n1371), .Y(n1282) );
  DFFXL R5_reg_28_ ( .D(n1282), .CK(clk), .Q(n134), .QN(n794) );
  MX2X1 R4_reg_28__U3 ( .A(n270), .B(data_in_3[62]), .S0(n1360), .Y(n1281) );
  DFFXL R4_reg_28_ ( .D(n1281), .CK(clk), .Q(n270), .QN(n726) );
  DFFXL R7_reg_16_ ( .D(n1280), .CK(clk), .Q(n530), .QN(n602) );
  MX2X1 R6_reg_16__U3 ( .A(n394), .B(data_in_3[50]), .S0(n1376), .Y(n1279) );
  DFFXL R6_reg_16_ ( .D(n1279), .CK(clk), .Q(n394), .QN(n670) );
  MX2X1 R5_reg_16__U3 ( .A(n122), .B(data_in_3[50]), .S0(n1370), .Y(n1278) );
  DFFXL R5_reg_16_ ( .D(n1278), .CK(clk), .Q(n122), .QN(n806) );
  MX2X1 R4_reg_16__U3 ( .A(n258), .B(data_in_3[50]), .S0(n1359), .Y(n1277) );
  DFFXL R4_reg_16_ ( .D(n1277), .CK(clk), .Q(n258), .QN(n738) );
  MX2X1 R11_reg_24__U3 ( .A(n368), .B(data_in_3[92]), .S0(n1343), .Y(n1276) );
  DFFXL R11_reg_24_ ( .D(n1276), .CK(clk), .Q(n368), .QN(n696) );
  MX2X1 R10_reg_24__U3 ( .A(n436), .B(data_in_3[92]), .S0(n1379), .Y(n1275) );
  DFFXL R10_reg_24_ ( .D(n1275), .CK(clk), .Q(n436), .QN(n628) );
  MX2X1 R9_reg_24__U3 ( .A(n96), .B(data_in_3[92]), .S0(n1367), .Y(n1274) );
  DFFXL R9_reg_24_ ( .D(n1274), .CK(clk), .Q(n96), .QN(n832) );
  MX2X1 R8_reg_24__U3 ( .A(n232), .B(data_in_3[92]), .S0(n1356), .Y(n1273) );
  DFFXL R8_reg_24_ ( .D(n1273), .CK(clk), .Q(n232), .QN(n764) );
  MX2X1 R7_reg_31__U3 ( .A(n545), .B(data_in_3[65]), .S0(n1348), .Y(n1272) );
  DFFXL R7_reg_31_ ( .D(n1272), .CK(clk), .Q(n545), .QN(n587) );
  MX2X1 R6_reg_31__U3 ( .A(n409), .B(data_in_3[65]), .S0(n1377), .Y(n1271) );
  DFFXL R6_reg_31_ ( .D(n1271), .CK(clk), .Q(n409), .QN(n655) );
  DFFXL R5_reg_31_ ( .D(n1270), .CK(clk), .Q(n137), .QN(n791) );
  DFFXL R4_reg_31_ ( .D(n1269), .CK(clk), .Q(n273), .QN(n723) );
  DFFXL R11_reg_32_ ( .D(n1268), .CK(clk), .Q(n376), .QN(n688) );
  DFFXL R10_reg_32_ ( .D(n1267), .CK(clk), .Q(n444), .QN(n620) );
  DFFXL R9_reg_32_ ( .D(n1266), .CK(clk), .Q(n104), .QN(n824) );
  MX2X1 R8_reg_32__U3 ( .A(n240), .B(data_in_3[100]), .S0(n1357), .Y(n1265) );
  DFFXL R8_reg_32_ ( .D(n1265), .CK(clk), .Q(n240), .QN(n756) );
  DFFXL R11_reg_30_ ( .D(n1264), .CK(clk), .Q(n374), .QN(n690) );
  DFFXL R10_reg_30_ ( .D(n1263), .CK(clk), .Q(n442), .QN(n622) );
  MX2X1 R9_reg_30__U3 ( .A(n102), .B(data_in_3[98]), .S0(n1368), .Y(n1262) );
  DFFXL R9_reg_30_ ( .D(n1262), .CK(clk), .Q(n102), .QN(n826) );
  MX2X1 R8_reg_30__U3 ( .A(n238), .B(data_in_3[98]), .S0(n1357), .Y(n1261) );
  DFFXL R8_reg_30_ ( .D(n1261), .CK(clk), .Q(n238), .QN(n758) );
  DFFXL R11_reg_31_ ( .D(n1260), .CK(clk), .Q(n375), .QN(n689) );
  DFFXL R10_reg_31_ ( .D(n1259), .CK(clk), .Q(n443), .QN(n621) );
  MX2X1 R7_reg_15__U3 ( .A(n529), .B(data_in_3[49]), .S0(n1348), .Y(n1258) );
  DFFXL R7_reg_15_ ( .D(n1258), .CK(clk), .Q(n529), .QN(n603) );
  DFFXL R7_reg_14_ ( .D(n1257), .CK(clk), .Q(n528), .QN(n604) );
  MX2X1 R6_reg_15__U3 ( .A(n393), .B(data_in_3[49]), .S0(n1376), .Y(n1256) );
  DFFXL R6_reg_15_ ( .D(n1256), .CK(clk), .Q(n393), .QN(n671) );
  DFFXL R6_reg_14_ ( .D(n1255), .CK(clk), .Q(n392), .QN(n672) );
  MX2X1 R5_reg_15__U3 ( .A(n121), .B(data_in_3[49]), .S0(n1369), .Y(n1254) );
  DFFXL R5_reg_15_ ( .D(n1254), .CK(clk), .Q(n121), .QN(n807) );
  DFFXL R5_reg_14_ ( .D(n1253), .CK(clk), .Q(n120), .QN(n808) );
  DFFXL R4_reg_15_ ( .D(n1252), .CK(clk), .Q(n257), .QN(n739) );
  DFFXL R4_reg_14_ ( .D(n1251), .CK(clk), .Q(n256), .QN(n740) );
  MX2X1 R7_reg_32__U3 ( .A(n546), .B(data_in_3[66]), .S0(n1344), .Y(n1250) );
  DFFXL R7_reg_32_ ( .D(n1250), .CK(clk), .Q(n546), .QN(n586) );
  MX2X1 R6_reg_32__U3 ( .A(n410), .B(data_in_3[66]), .S0(n1377), .Y(n1249) );
  DFFXL R6_reg_32_ ( .D(n1249), .CK(clk), .Q(n410), .QN(n654) );
  MX2X1 R5_reg_32__U3 ( .A(n138), .B(data_in_3[66]), .S0(n1371), .Y(n1248) );
  DFFXL R5_reg_32_ ( .D(n1248), .CK(clk), .Q(n138), .QN(n790) );
  MX2X1 R4_reg_32__U3 ( .A(n274), .B(data_in_3[66]), .S0(n1360), .Y(n1247) );
  DFFXL R4_reg_32_ ( .D(n1247), .CK(clk), .Q(n274), .QN(n722) );
  MX2X1 R6_reg_12__U3 ( .A(n390), .B(data_in_3[46]), .S0(n1376), .Y(n1246) );
  DFFXL R6_reg_12_ ( .D(n1246), .CK(clk), .Q(n390), .QN(n674) );
  MX2X1 R5_reg_12__U3 ( .A(n118), .B(data_in_3[46]), .S0(n1369), .Y(n1245) );
  DFFXL R5_reg_12_ ( .D(n1245), .CK(clk), .Q(n118), .QN(n810) );
  MX2X1 R4_reg_12__U3 ( .A(n254), .B(data_in_3[46]), .S0(n1358), .Y(n1244) );
  DFFXL R4_reg_12_ ( .D(n1244), .CK(clk), .Q(n254), .QN(n742) );
  MX2X1 R7_reg_9__U3 ( .A(n523), .B(data_in_3[43]), .S0(n1348), .Y(n1243) );
  DFFXL R7_reg_9_ ( .D(n1243), .CK(clk), .Q(n523), .QN(n609) );
  MX2X1 R6_reg_9__U3 ( .A(n387), .B(data_in_3[43]), .S0(n1375), .Y(n1242) );
  DFFXL R6_reg_9_ ( .D(n1242), .CK(clk), .Q(n387), .QN(n677) );
  MX2X1 R5_reg_9__U3 ( .A(n115), .B(data_in_3[43]), .S0(n1369), .Y(n1241) );
  DFFXL R5_reg_9_ ( .D(n1241), .CK(clk), .Q(n115), .QN(n813) );
  MX2X1 R4_reg_9__U3 ( .A(n251), .B(data_in_3[43]), .S0(n1358), .Y(n1240) );
  DFFXL R4_reg_9_ ( .D(n1240), .CK(clk), .Q(n251), .QN(n745) );
  DFFXL R7_reg_13_ ( .D(n1239), .CK(clk), .Q(n527), .QN(n605) );
  DFFXL R6_reg_13_ ( .D(n1238), .CK(clk), .Q(n391), .QN(n673) );
  DFFXL R11_reg_13_ ( .D(n1237), .CK(clk), .Q(n357), .QN(n707) );
  MX2X1 R10_reg_13__U3 ( .A(n425), .B(data_in_3[81]), .S0(n1378), .Y(n1236) );
  DFFXL R10_reg_13_ ( .D(n1236), .CK(clk), .Q(n425), .QN(n639) );
  MX2X1 R9_reg_13__U3 ( .A(n85), .B(data_in_3[81]), .S0(n1366), .Y(n1235) );
  DFFXL R9_reg_13_ ( .D(n1235), .CK(clk), .Q(n85), .QN(n843) );
  MX2X1 R8_reg_13__U3 ( .A(n221), .B(data_in_3[81]), .S0(n1355), .Y(n1234) );
  DFFXL R8_reg_13_ ( .D(n1234), .CK(clk), .Q(n221), .QN(n775) );
  DFFXL R11_reg_33_ ( .D(n1233), .CK(clk), .Q(n377), .QN(n687) );
  MX2X1 R10_reg_33__U3 ( .A(n445), .B(data_in_3[101]), .S0(n1380), .Y(n1232)
         );
  DFFXL R10_reg_33_ ( .D(n1232), .CK(clk), .Q(n445), .QN(n619) );
  MX2X1 R9_reg_33__U3 ( .A(n105), .B(data_in_3[101]), .S0(n1368), .Y(n1231) );
  DFFXL R9_reg_33_ ( .D(n1231), .CK(clk), .Q(n105), .QN(n823) );
  MX2X1 R8_reg_33__U3 ( .A(n241), .B(data_in_3[101]), .S0(n1357), .Y(n1230) );
  DFFXL R8_reg_33_ ( .D(n1230), .CK(clk), .Q(n241), .QN(n755) );
  MX2X1 R7_reg_11__U3 ( .A(n525), .B(data_in_3[45]), .S0(n1348), .Y(n1229) );
  DFFXL R7_reg_11_ ( .D(n1229), .CK(clk), .Q(n525), .QN(n607) );
  MX2X1 R6_reg_11__U3 ( .A(n389), .B(data_in_3[45]), .S0(n1375), .Y(n1228) );
  DFFXL R6_reg_11_ ( .D(n1228), .CK(clk), .Q(n389), .QN(n675) );
  MX2X1 R5_reg_11__U3 ( .A(n117), .B(data_in_3[45]), .S0(n1369), .Y(n1227) );
  DFFXL R5_reg_11_ ( .D(n1227), .CK(clk), .Q(n117), .QN(n811) );
  DFFXL R4_reg_11_ ( .D(n1226), .CK(clk), .Q(n253), .QN(n743) );
  MX2X1 R7_reg_33__U3 ( .A(n547), .B(data_in_3[67]), .S0(n1346), .Y(n1225) );
  DFFXL R7_reg_33_ ( .D(n1225), .CK(clk), .Q(n547), .QN(n585) );
  DFFXL R6_reg_33_ ( .D(n1224), .CK(clk), .Q(n411), .QN(n653) );
  DFFXL R5_reg_33_ ( .D(n1223), .CK(clk), .Q(n139), .QN(n789) );
  DFFXL R4_reg_33_ ( .D(n1222), .CK(clk), .Q(n275), .QN(n721) );
  DFFXL R3_reg_33_ ( .D(n1221), .CK(clk), .Q(R3[33]) );
  DFFXL R2_reg_33_ ( .D(n1219), .CK(clk), .Q(R2[33]) );
  DFFXL R1_reg_33_ ( .D(n1217), .CK(clk), .Q(R1[33]) );
  DFFXL R0_reg_33_ ( .D(n1215), .CK(clk), .Q(R0[33]) );
  MX2X1 R15_reg_28__U3 ( .A(R15[28]), .B(data_in_3[130]), .S0(n1342), .Y(n1213) );
  DFFXL R15_reg_28_ ( .D(n1213), .CK(clk), .Q(R15[28]) );
  MX2X1 R14_reg_28__U3 ( .A(R14[28]), .B(data_in_3[130]), .S0(n1381), .Y(n1211) );
  DFFXL R14_reg_28_ ( .D(n1211), .CK(clk), .Q(R14[28]) );
  MX2X1 R13_reg_28__U3 ( .A(R13[28]), .B(data_in_3[130]), .S0(n1365), .Y(n1209) );
  DFFXL R13_reg_28_ ( .D(n1209), .CK(clk), .Q(R13[28]) );
  MX2X1 R12_reg_28__U3 ( .A(R12[28]), .B(data_in_3[130]), .S0(n1354), .Y(n1207) );
  DFFXL R12_reg_28_ ( .D(n1207), .CK(clk), .Q(R12[28]) );
  MX2X1 R3_reg_14__U3 ( .A(R3[14]), .B(data_in_3[14]), .S0(n1345), .Y(n1205)
         );
  DFFXL R3_reg_14_ ( .D(n1205), .CK(clk), .Q(R3[14]) );
  MX2X1 R2_reg_14__U3 ( .A(R2[14]), .B(data_in_3[14]), .S0(n1376), .Y(n1203)
         );
  DFFXL R2_reg_14_ ( .D(n1203), .CK(clk), .Q(R2[14]) );
  DFFXL R1_reg_14_ ( .D(n1201), .CK(clk), .Q(R1[14]) );
  MX2X1 R0_reg_14__U3 ( .A(R0[14]), .B(data_in_3[14]), .S0(n1361), .Y(n1199)
         );
  DFFXL R0_reg_14_ ( .D(n1199), .CK(clk), .Q(R0[14]) );
  DFFXL R3_reg_13_ ( .D(n1197), .CK(clk), .Q(R3[13]) );
  DFFXL R2_reg_13_ ( .D(n1195), .CK(clk), .Q(R2[13]) );
  DFFXL R1_reg_13_ ( .D(n1193), .CK(clk), .Q(R1[13]) );
  DFFXL R0_reg_13_ ( .D(n1191), .CK(clk), .Q(R0[13]) );
  MX2X1 R15_reg_31__U3 ( .A(R15[31]), .B(data_in_3[133]), .S0(n1342), .Y(n1189) );
  DFFXL R15_reg_31_ ( .D(n1189), .CK(clk), .Q(R15[31]) );
  MX2X1 R14_reg_31__U3 ( .A(R14[31]), .B(data_in_3[133]), .S0(n1383), .Y(n1187) );
  DFFXL R14_reg_31_ ( .D(n1187), .CK(clk), .Q(R14[31]) );
  MX2X1 R13_reg_31__U3 ( .A(R13[31]), .B(data_in_3[133]), .S0(n1365), .Y(n1185) );
  DFFXL R13_reg_31_ ( .D(n1185), .CK(clk), .Q(R13[31]) );
  DFFXL R12_reg_31_ ( .D(n1183), .CK(clk), .Q(R12[31]) );
  MX2X1 R3_reg_11__U3 ( .A(R3[11]), .B(data_in_3[11]), .S0(n1345), .Y(n1181)
         );
  DFFXL R3_reg_11_ ( .D(n1181), .CK(clk), .Q(R3[11]) );
  MX2X1 R2_reg_11__U3 ( .A(R2[11]), .B(data_in_3[11]), .S0(n1382), .Y(n1179)
         );
  DFFXL R2_reg_11_ ( .D(n1179), .CK(clk), .Q(R2[11]) );
  MX2X1 R1_reg_11__U3 ( .A(R1[11]), .B(data_in_3[11]), .S0(n1372), .Y(n1177)
         );
  DFFXL R1_reg_11_ ( .D(n1177), .CK(clk), .Q(R1[11]) );
  MX2X1 R0_reg_11__U3 ( .A(R0[11]), .B(data_in_3[11]), .S0(n1361), .Y(n1175)
         );
  DFFXL R0_reg_11_ ( .D(n1175), .CK(clk), .Q(R0[11]) );
  DFFXL R3_reg_30_ ( .D(n1173), .CK(clk), .Q(R3[30]) );
  MX2X1 R2_reg_30__U3 ( .A(R2[30]), .B(data_in_3[30]), .S0(n1383), .Y(n1171)
         );
  DFFXL R2_reg_30_ ( .D(n1171), .CK(clk), .Q(R2[30]) );
  MX2X1 R1_reg_30__U3 ( .A(R1[30]), .B(data_in_3[30]), .S0(n1366), .Y(n1169)
         );
  DFFXL R1_reg_30_ ( .D(n1169), .CK(clk), .Q(R1[30]) );
  MX2X1 R0_reg_30__U3 ( .A(R0[30]), .B(data_in_3[30]), .S0(n1355), .Y(n1167)
         );
  DFFXL R0_reg_30_ ( .D(n1167), .CK(clk), .Q(R0[30]) );
  MX2X1 R15_reg_32__U3 ( .A(R15[32]), .B(data_in_3[134]), .S0(n1342), .Y(n1165) );
  DFFXL R15_reg_32_ ( .D(n1165), .CK(clk), .Q(R15[32]) );
  DFFXL R14_reg_32_ ( .D(n893), .CK(clk), .Q(R14[32]) );
  MX2X1 R13_reg_32__U3 ( .A(R13[32]), .B(data_in_3[134]), .S0(n1365), .Y(n890)
         );
  DFFXL R13_reg_32_ ( .D(n890), .CK(clk), .Q(R13[32]) );
  DFFXL R12_reg_32_ ( .D(n881), .CK(clk), .Q(R12[32]) );
  DFFXL R15_reg_30_ ( .D(n866), .CK(clk), .Q(R15[30]) );
  DFFXL R14_reg_30_ ( .D(n864), .CK(clk), .Q(R14[30]) );
  DFFXL R13_reg_30_ ( .D(n862), .CK(clk), .Q(R13[30]) );
  DFFXL R12_reg_30_ ( .D(n859), .CK(clk), .Q(R12[30]) );
  DFFXL R3_reg_15_ ( .D(n857), .CK(clk), .Q(R3[15]) );
  DFFXL R2_reg_15_ ( .D(n581), .CK(clk), .Q(R2[15]) );
  DFFXL R1_reg_15_ ( .D(n579), .CK(clk), .Q(R1[15]) );
  DFFXL R0_reg_15_ ( .D(n577), .CK(clk), .Q(R0[15]) );
  DFFXL R3_reg_31_ ( .D(n575), .CK(clk), .Q(R3[31]) );
  DFFXL R2_reg_31_ ( .D(n573), .CK(clk), .Q(R2[31]) );
  DFFXL R1_reg_31_ ( .D(n571), .CK(clk), .Q(R1[31]) );
  DFFXL R0_reg_31_ ( .D(n569), .CK(clk), .Q(R0[31]) );
  DFFXL R3_reg_32_ ( .D(n567), .CK(clk), .Q(R3[32]) );
  DFFXL R2_reg_32_ ( .D(n565), .CK(clk), .Q(R2[32]) );
  DFFXL R1_reg_32_ ( .D(n563), .CK(clk), .Q(R1[32]) );
  DFFXL R0_reg_32_ ( .D(n561), .CK(clk), .Q(R0[32]) );
  MX2X1 R15_reg_16__U3 ( .A(R15[16]), .B(data_in_3[118]), .S0(n1341), .Y(n559)
         );
  DFFXL R15_reg_16_ ( .D(n559), .CK(clk), .Q(R15[16]) );
  MX2X1 R14_reg_16__U3 ( .A(R14[16]), .B(data_in_3[118]), .S0(n1382), .Y(n557)
         );
  DFFXL R14_reg_16_ ( .D(n557), .CK(clk), .Q(R14[16]) );
  MX2X1 R13_reg_16__U3 ( .A(R13[16]), .B(data_in_3[118]), .S0(n1364), .Y(n555)
         );
  DFFXL R13_reg_16_ ( .D(n555), .CK(clk), .Q(R13[16]) );
  MX2X1 R12_reg_16__U3 ( .A(R12[16]), .B(data_in_3[118]), .S0(n1353), .Y(n553)
         );
  DFFXL R12_reg_16_ ( .D(n553), .CK(clk), .Q(R12[16]) );
  MX2X1 R15_reg_13__U3 ( .A(R15[13]), .B(data_in_3[115]), .S0(n1341), .Y(n551)
         );
  DFFXL R15_reg_13_ ( .D(n551), .CK(clk), .Q(R15[13]) );
  DFFXL R14_reg_13_ ( .D(n549), .CK(clk), .Q(R14[13]) );
  MX2X1 R13_reg_13__U3 ( .A(R13[13]), .B(data_in_3[115]), .S0(n1364), .Y(n544)
         );
  DFFXL R13_reg_13_ ( .D(n544), .CK(clk), .Q(R13[13]) );
  DFFXL R12_reg_13_ ( .D(n541), .CK(clk), .Q(R12[13]) );
  DFFXL R15_reg_33_ ( .D(n539), .CK(clk), .Q(R15[33]) );
  MX2X1 R14_reg_33__U3 ( .A(R14[33]), .B(data_in_3[135]), .S0(n1379), .Y(n537)
         );
  DFFXL R14_reg_33_ ( .D(n537), .CK(clk), .Q(R14[33]) );
  MX2X1 R13_reg_33__U3 ( .A(R13[33]), .B(data_in_3[135]), .S0(n1365), .Y(n535)
         );
  DFFXL R13_reg_33_ ( .D(n535), .CK(clk), .Q(R13[33]) );
  MX2X1 R12_reg_33__U3 ( .A(R12[33]), .B(data_in_3[135]), .S0(n1354), .Y(n533)
         );
  DFFXL R12_reg_33_ ( .D(n533), .CK(clk), .Q(R12[33]) );
  MX2X1 R15_reg_15__U3 ( .A(R15[15]), .B(data_in_3[117]), .S0(n1341), .Y(n531)
         );
  DFFXL R15_reg_15_ ( .D(n531), .CK(clk), .Q(R15[15]) );
  MX2X1 R15_reg_14__U3 ( .A(R15[14]), .B(data_in_3[116]), .S0(n1341), .Y(n524)
         );
  DFFXL R15_reg_14_ ( .D(n524), .CK(clk), .Q(R15[14]) );
  DFFXL R14_reg_15_ ( .D(n521), .CK(clk), .Q(R14[15]) );
  DFFXL R14_reg_14_ ( .D(n519), .CK(clk), .Q(R14[14]) );
  MX2X1 R13_reg_15__U3 ( .A(R13[15]), .B(data_in_3[117]), .S0(n1364), .Y(n517)
         );
  DFFXL R13_reg_15_ ( .D(n517), .CK(clk), .Q(R13[15]) );
  MX2X1 R13_reg_14__U3 ( .A(R13[14]), .B(data_in_3[116]), .S0(n1364), .Y(n515)
         );
  DFFXL R13_reg_14_ ( .D(n515), .CK(clk), .Q(R13[14]) );
  DFFXL R12_reg_15_ ( .D(n513), .CK(clk), .Q(R12[15]) );
  MX2X1 R12_reg_14__U3 ( .A(R12[14]), .B(data_in_3[116]), .S0(n1353), .Y(n511)
         );
  DFFXL R12_reg_14_ ( .D(n511), .CK(clk), .Q(R12[14]) );
  EDFFX1 R7_reg_23_ ( .D(data_in_3[57]), .E(n1348), .CK(clk), .QN(n595) );
  EDFFX1 R7_reg_22_ ( .D(data_in_3[56]), .E(n19), .CK(clk), .QN(n596) );
  EDFFXL R7_reg_21_ ( .D(data_in_3[55]), .E(n19), .CK(clk), .QN(n597) );
  EDFFX1 R7_reg_20_ ( .D(data_in_3[54]), .E(n19), .CK(clk), .QN(n598) );
  EDFFX1 R7_reg_19_ ( .D(data_in_3[53]), .E(n1347), .CK(clk), .QN(n599) );
  EDFFX1 R7_reg_18_ ( .D(data_in_3[52]), .E(n1343), .CK(clk), .QN(n600) );
  EDFFX1 R7_reg_17_ ( .D(data_in_3[51]), .E(n1348), .CK(clk), .QN(n601) );
  EDFFX1 R7_reg_10_ ( .D(data_in_3[44]), .E(n1348), .CK(clk), .QN(n608) );
  EDFFX1 R7_reg_7_ ( .D(data_in_3[41]), .E(n1348), .CK(clk), .QN(n611) );
  EDFFX1 R7_reg_3_ ( .D(data_in_3[37]), .E(n1347), .CK(clk), .QN(n615) );
  EDFFX1 R7_reg_2_ ( .D(data_in_3[36]), .E(n1347), .CK(clk), .QN(n616) );
  EDFFX1 R7_reg_1_ ( .D(data_in_3[35]), .E(n1347), .CK(clk), .QN(n617) );
  EDFFX1 R7_reg_0_ ( .D(data_in_3[34]), .E(n1347), .CK(clk), .QN(n618) );
  EDFFX1 R6_reg_23_ ( .D(data_in_3[57]), .E(n1376), .CK(clk), .QN(n663) );
  EDFFX1 R6_reg_22_ ( .D(data_in_3[56]), .E(n1376), .CK(clk), .QN(n664) );
  EDFFXL R6_reg_21_ ( .D(data_in_3[55]), .E(n1376), .CK(clk), .QN(n665) );
  EDFFX1 R6_reg_20_ ( .D(data_in_3[54]), .E(n1376), .CK(clk), .QN(n666) );
  EDFFX1 R6_reg_19_ ( .D(data_in_3[53]), .E(n1376), .CK(clk), .QN(n667) );
  EDFFX1 R6_reg_18_ ( .D(data_in_3[52]), .E(n1376), .CK(clk), .QN(n668) );
  EDFFX1 R6_reg_17_ ( .D(data_in_3[51]), .E(n1376), .CK(clk), .QN(n669) );
  EDFFX1 R6_reg_10_ ( .D(data_in_3[44]), .E(n1375), .CK(clk), .QN(n676) );
  EDFFX1 R6_reg_7_ ( .D(data_in_3[41]), .E(n1375), .CK(clk), .QN(n679) );
  EDFFX1 R6_reg_3_ ( .D(data_in_3[37]), .E(n1375), .CK(clk), .QN(n683) );
  EDFFX1 R6_reg_2_ ( .D(data_in_3[36]), .E(n1375), .CK(clk), .QN(n684) );
  EDFFX1 R6_reg_1_ ( .D(data_in_3[35]), .E(n1375), .CK(clk), .QN(n685) );
  EDFFX1 R6_reg_0_ ( .D(data_in_3[34]), .E(n1375), .CK(clk), .QN(n686) );
  EDFFX1 R4_reg_23_ ( .D(data_in_3[57]), .E(n1359), .CK(clk), .QN(n731) );
  EDFFX1 R4_reg_22_ ( .D(data_in_3[56]), .E(n1359), .CK(clk), .QN(n732) );
  EDFFXL R4_reg_21_ ( .D(data_in_3[55]), .E(n1359), .CK(clk), .QN(n733) );
  EDFFX1 R4_reg_20_ ( .D(data_in_3[54]), .E(n1359), .CK(clk), .QN(n734) );
  EDFFX1 R4_reg_19_ ( .D(data_in_3[53]), .E(n1359), .CK(clk), .QN(n735) );
  EDFFX1 R4_reg_18_ ( .D(data_in_3[52]), .E(n1359), .CK(clk), .QN(n736) );
  EDFFX1 R4_reg_17_ ( .D(data_in_3[51]), .E(n1359), .CK(clk), .QN(n737) );
  EDFFX1 R4_reg_10_ ( .D(data_in_3[44]), .E(n1358), .CK(clk), .QN(n744) );
  EDFFX1 R4_reg_7_ ( .D(data_in_3[41]), .E(n1358), .CK(clk), .QN(n747) );
  EDFFX1 R4_reg_3_ ( .D(data_in_3[37]), .E(n1357), .CK(clk), .QN(n751) );
  EDFFX1 R4_reg_2_ ( .D(data_in_3[36]), .E(n1357), .CK(clk), .QN(n752) );
  EDFFX1 R4_reg_1_ ( .D(data_in_3[35]), .E(n1357), .CK(clk), .QN(n753) );
  EDFFX1 R4_reg_0_ ( .D(data_in_3[34]), .E(n1357), .CK(clk), .QN(n754) );
  EDFFXL R5_reg_30_ ( .D(data_in_3[64]), .E(n1371), .CK(clk), .QN(n792) );
  EDFFXL R5_reg_29_ ( .D(data_in_3[63]), .E(n1371), .CK(clk), .QN(n793) );
  EDFFXL R5_reg_25_ ( .D(data_in_3[59]), .E(n1370), .CK(clk), .QN(n797) );
  EDFFXL R5_reg_24_ ( .D(data_in_3[58]), .E(n1370), .CK(clk), .QN(n798) );
  EDFFXL R5_reg_21_ ( .D(data_in_3[55]), .E(n1370), .CK(clk), .QN(n801) );
  EDFFX1 R5_reg_20_ ( .D(data_in_3[54]), .E(n1370), .CK(clk), .QN(n802) );
  EDFFX1 R5_reg_19_ ( .D(data_in_3[53]), .E(n1370), .CK(clk), .QN(n803) );
  EDFFX1 R5_reg_18_ ( .D(data_in_3[52]), .E(n1370), .CK(clk), .QN(n804) );
  EDFFX1 R5_reg_17_ ( .D(data_in_3[51]), .E(n1370), .CK(clk), .QN(n805) );
  EDFFXL R5_reg_8_ ( .D(data_in_3[42]), .E(n1369), .CK(clk), .QN(n814) );
  EDFFXL R5_reg_5_ ( .D(n83), .E(n1369), .CK(clk), .QN(n817) );
  EDFFXL R5_reg_4_ ( .D(data_in_3[38]), .E(n1369), .CK(clk), .QN(n818) );
  EDFFX1 R5_reg_3_ ( .D(data_in_3[37]), .E(n1368), .CK(clk), .QN(n819) );
  EDFFX1 R5_reg_2_ ( .D(data_in_3[36]), .E(n1368), .CK(clk), .QN(n820) );
  EDFFX1 R5_reg_1_ ( .D(data_in_3[35]), .E(n1368), .CK(clk), .QN(n821) );
  EDFFX1 R5_reg_0_ ( .D(data_in_3[34]), .E(n1368), .CK(clk), .QN(n822) );
  EDFFXL R10_reg_29_ ( .D(data_in_3[97]), .E(n1380), .CK(clk), .QN(n623) );
  EDFFXL R10_reg_28_ ( .D(data_in_3[96]), .E(n1380), .CK(clk), .QN(n624) );
  EDFFXL R10_reg_27_ ( .D(data_in_3[95]), .E(n1380), .CK(clk), .QN(n625) );
  EDFFXL R10_reg_26_ ( .D(data_in_3[94]), .E(n1380), .CK(clk), .QN(n626) );
  EDFFXL R10_reg_25_ ( .D(data_in_3[93]), .E(n1379), .CK(clk), .QN(n627) );
  EDFFX1 R10_reg_20_ ( .D(data_in_3[88]), .E(n1379), .CK(clk), .QN(n632) );
  EDFFX1 R10_reg_19_ ( .D(data_in_3[87]), .E(n1379), .CK(clk), .QN(n633) );
  EDFFX1 R10_reg_18_ ( .D(data_in_3[86]), .E(n1379), .CK(clk), .QN(n634) );
  EDFFX1 R10_reg_17_ ( .D(data_in_3[85]), .E(n1379), .CK(clk), .QN(n635) );
  EDFFXL R10_reg_12_ ( .D(data_in_3[80]), .E(n1378), .CK(clk), .QN(n640) );
  EDFFXL R10_reg_11_ ( .D(data_in_3[79]), .E(n1378), .CK(clk), .QN(n641) );
  EDFFXL R10_reg_10_ ( .D(data_in_3[78]), .E(n1378), .CK(clk), .QN(n642) );
  EDFFXL R10_reg_9_ ( .D(data_in_3[77]), .E(n1378), .CK(clk), .QN(n643) );
  EDFFXL R10_reg_7_ ( .D(data_in_3[75]), .E(n1378), .CK(clk), .QN(n645) );
  EDFFXL R10_reg_4_ ( .D(data_in_3[72]), .E(n1378), .CK(clk), .QN(n648) );
  EDFFX1 R10_reg_3_ ( .D(data_in_3[71]), .E(n1378), .CK(clk), .QN(n649) );
  EDFFX1 R10_reg_2_ ( .D(data_in_3[70]), .E(n1378), .CK(clk), .QN(n650) );
  EDFFX1 R10_reg_1_ ( .D(data_in_3[69]), .E(n1377), .CK(clk), .QN(n651) );
  EDFFX1 R10_reg_0_ ( .D(data_in_3[68]), .E(n1377), .CK(clk), .QN(n652) );
  EDFFXL R11_reg_29_ ( .D(data_in_3[97]), .E(n1344), .CK(clk), .QN(n691) );
  EDFFXL R11_reg_28_ ( .D(data_in_3[96]), .E(n1344), .CK(clk), .QN(n692) );
  EDFFXL R11_reg_27_ ( .D(data_in_3[95]), .E(n1344), .CK(clk), .QN(n693) );
  EDFFXL R11_reg_26_ ( .D(data_in_3[94]), .E(n1344), .CK(clk), .QN(n694) );
  EDFFXL R11_reg_25_ ( .D(data_in_3[93]), .E(n1343), .CK(clk), .QN(n695) );
  EDFFX1 R11_reg_20_ ( .D(data_in_3[88]), .E(n1343), .CK(clk), .QN(n700) );
  EDFFX1 R11_reg_19_ ( .D(data_in_3[87]), .E(n1343), .CK(clk), .QN(n701) );
  EDFFX1 R11_reg_18_ ( .D(data_in_3[86]), .E(n1343), .CK(clk), .QN(n702) );
  EDFFX1 R11_reg_17_ ( .D(data_in_3[85]), .E(n1343), .CK(clk), .QN(n703) );
  EDFFXL R11_reg_12_ ( .D(data_in_3[80]), .E(n1347), .CK(clk), .QN(n708) );
  EDFFXL R11_reg_11_ ( .D(data_in_3[79]), .E(n1343), .CK(clk), .QN(n709) );
  EDFFXL R11_reg_10_ ( .D(data_in_3[78]), .E(n1346), .CK(clk), .QN(n710) );
  EDFFXL R11_reg_9_ ( .D(data_in_3[77]), .E(n1342), .CK(clk), .QN(n711) );
  EDFFXL R11_reg_7_ ( .D(data_in_3[75]), .E(n1347), .CK(clk), .QN(n713) );
  EDFFXL R11_reg_4_ ( .D(data_in_3[72]), .E(n1347), .CK(clk), .QN(n716) );
  EDFFX1 R11_reg_3_ ( .D(data_in_3[71]), .E(n1347), .CK(clk), .QN(n717) );
  EDFFX1 R11_reg_2_ ( .D(data_in_3[70]), .E(n1347), .CK(clk), .QN(n718) );
  EDFFX1 R11_reg_1_ ( .D(data_in_3[69]), .E(n1342), .CK(clk), .QN(n719) );
  EDFFX1 R11_reg_0_ ( .D(data_in_3[68]), .E(n1342), .CK(clk), .QN(n720) );
  EDFFXL R8_reg_29_ ( .D(data_in_3[97]), .E(n1357), .CK(clk), .QN(n759) );
  EDFFXL R8_reg_28_ ( .D(data_in_3[96]), .E(n1357), .CK(clk), .QN(n760) );
  EDFFXL R8_reg_27_ ( .D(data_in_3[95]), .E(n1357), .CK(clk), .QN(n761) );
  EDFFXL R8_reg_26_ ( .D(data_in_3[94]), .E(n1357), .CK(clk), .QN(n762) );
  EDFFXL R8_reg_25_ ( .D(data_in_3[93]), .E(n1356), .CK(clk), .QN(n763) );
  EDFFX1 R8_reg_20_ ( .D(data_in_3[88]), .E(n1356), .CK(clk), .QN(n768) );
  EDFFX1 R8_reg_19_ ( .D(data_in_3[87]), .E(n1356), .CK(clk), .QN(n769) );
  EDFFX1 R8_reg_18_ ( .D(data_in_3[86]), .E(n1356), .CK(clk), .QN(n770) );
  EDFFX1 R8_reg_17_ ( .D(data_in_3[85]), .E(n1356), .CK(clk), .QN(n771) );
  EDFFXL R8_reg_12_ ( .D(data_in_3[80]), .E(n1355), .CK(clk), .QN(n776) );
  EDFFXL R8_reg_11_ ( .D(data_in_3[79]), .E(n1355), .CK(clk), .QN(n777) );
  EDFFXL R8_reg_10_ ( .D(data_in_3[78]), .E(n1355), .CK(clk), .QN(n778) );
  EDFFXL R8_reg_9_ ( .D(data_in_3[77]), .E(n1355), .CK(clk), .QN(n779) );
  EDFFXL R8_reg_7_ ( .D(data_in_3[75]), .E(n1355), .CK(clk), .QN(n781) );
  EDFFXL R8_reg_4_ ( .D(data_in_3[72]), .E(n1355), .CK(clk), .QN(n784) );
  EDFFX1 R8_reg_3_ ( .D(data_in_3[71]), .E(n1355), .CK(clk), .QN(n785) );
  EDFFX1 R8_reg_2_ ( .D(data_in_3[70]), .E(n1355), .CK(clk), .QN(n786) );
  EDFFX1 R8_reg_1_ ( .D(data_in_3[69]), .E(n1354), .CK(clk), .QN(n787) );
  EDFFX1 R8_reg_0_ ( .D(data_in_3[68]), .E(n1354), .CK(clk), .QN(n788) );
  EDFFXL R9_reg_29_ ( .D(data_in_3[97]), .E(n1368), .CK(clk), .QN(n827) );
  EDFFXL R9_reg_28_ ( .D(data_in_3[96]), .E(n1368), .CK(clk), .QN(n828) );
  EDFFXL R9_reg_27_ ( .D(data_in_3[95]), .E(n1368), .CK(clk), .QN(n829) );
  EDFFXL R9_reg_26_ ( .D(data_in_3[94]), .E(n1368), .CK(clk), .QN(n830) );
  EDFFXL R9_reg_25_ ( .D(data_in_3[93]), .E(n1367), .CK(clk), .QN(n831) );
  EDFFX1 R9_reg_20_ ( .D(data_in_3[88]), .E(n1367), .CK(clk), .QN(n836) );
  EDFFX1 R9_reg_19_ ( .D(data_in_3[87]), .E(n1367), .CK(clk), .QN(n837) );
  EDFFX1 R9_reg_18_ ( .D(data_in_3[86]), .E(n1367), .CK(clk), .QN(n838) );
  EDFFX1 R9_reg_17_ ( .D(data_in_3[85]), .E(n1367), .CK(clk), .QN(n839) );
  EDFFXL R9_reg_12_ ( .D(data_in_3[80]), .E(n1366), .CK(clk), .QN(n844) );
  EDFFXL R9_reg_11_ ( .D(data_in_3[79]), .E(n1366), .CK(clk), .QN(n845) );
  EDFFXL R9_reg_10_ ( .D(data_in_3[78]), .E(n1366), .CK(clk), .QN(n846) );
  EDFFXL R9_reg_9_ ( .D(data_in_3[77]), .E(n1366), .CK(clk), .QN(n847) );
  EDFFXL R9_reg_7_ ( .D(data_in_3[75]), .E(n1366), .CK(clk), .QN(n849) );
  EDFFXL R9_reg_4_ ( .D(data_in_3[72]), .E(n1366), .CK(clk), .QN(n852) );
  EDFFX1 R9_reg_3_ ( .D(data_in_3[71]), .E(n1366), .CK(clk), .QN(n853) );
  EDFFX1 R9_reg_2_ ( .D(data_in_3[70]), .E(n1366), .CK(clk), .QN(n854) );
  EDFFX1 R9_reg_1_ ( .D(data_in_3[69]), .E(n1365), .CK(clk), .QN(n855) );
  EDFFX1 R9_reg_0_ ( .D(data_in_3[68]), .E(n1365), .CK(clk), .QN(n856) );
  EDFFXL R15_reg_29_ ( .D(data_in_3[131]), .E(n1342), .CK(clk), .Q(R15[29]) );
  EDFFXL R15_reg_27_ ( .D(data_in_3[129]), .E(n1342), .CK(clk), .Q(R15[27]) );
  EDFFXL R15_reg_26_ ( .D(data_in_3[128]), .E(n1342), .CK(clk), .Q(R15[26]) );
  EDFFXL R15_reg_25_ ( .D(data_in_3[127]), .E(n1342), .CK(clk), .Q(R15[25]) );
  EDFFXL R15_reg_23_ ( .D(data_in_3[125]), .E(n1341), .CK(clk), .Q(R15[23]) );
  EDFFXL R15_reg_22_ ( .D(data_in_3[124]), .E(n1341), .CK(clk), .Q(R15[22]) );
  EDFFX1 R15_reg_20_ ( .D(data_in_3[122]), .E(n1341), .CK(clk), .Q(R15[20]) );
  EDFFX1 R15_reg_19_ ( .D(data_in_3[121]), .E(n1341), .CK(clk), .Q(R15[19]) );
  EDFFX1 R15_reg_18_ ( .D(data_in_3[120]), .E(n1341), .CK(clk), .Q(R15[18]) );
  EDFFX1 R15_reg_17_ ( .D(data_in_3[119]), .E(n1341), .CK(clk), .Q(R15[17]) );
  EDFFXL R15_reg_12_ ( .D(data_in_3[114]), .E(n1341), .CK(clk), .Q(R15[12]) );
  EDFFXL R15_reg_11_ ( .D(data_in_3[113]), .E(n1342), .CK(clk), .Q(R15[11]) );
  EDFFXL R15_reg_10_ ( .D(data_in_3[112]), .E(n1343), .CK(clk), .Q(R15[10]) );
  EDFFXL R15_reg_9_ ( .D(data_in_3[111]), .E(n1341), .CK(clk), .Q(R15[9]) );
  EDFFXL R15_reg_8_ ( .D(data_in_3[110]), .E(n1344), .CK(clk), .Q(R15[8]) );
  EDFFXL R15_reg_7_ ( .D(data_in_3[109]), .E(n1346), .CK(clk), .Q(R15[7]) );
  EDFFXL R15_reg_6_ ( .D(data_in_3[108]), .E(n1348), .CK(clk), .Q(R15[6]) );
  EDFFXL R15_reg_4_ ( .D(data_in_3[106]), .E(n1345), .CK(clk), .Q(R15[4]) );
  EDFFX1 R15_reg_3_ ( .D(data_in_3[105]), .E(n1346), .CK(clk), .Q(R15[3]) );
  EDFFX1 R15_reg_2_ ( .D(data_in_3[104]), .E(n1345), .CK(clk), .Q(R15[2]) );
  EDFFX1 R15_reg_1_ ( .D(data_in_3[103]), .E(n1346), .CK(clk), .Q(R15[1]) );
  EDFFX1 R15_reg_0_ ( .D(data_in_3[102]), .E(n1345), .CK(clk), .Q(R15[0]) );
  EDFFXL R12_reg_29_ ( .D(data_in_3[131]), .E(n1354), .CK(clk), .Q(R12[29]) );
  EDFFXL R12_reg_27_ ( .D(data_in_3[129]), .E(n1354), .CK(clk), .Q(R12[27]) );
  EDFFXL R12_reg_26_ ( .D(data_in_3[128]), .E(n1354), .CK(clk), .Q(R12[26]) );
  EDFFXL R12_reg_25_ ( .D(data_in_3[127]), .E(n1354), .CK(clk), .Q(R12[25]) );
  EDFFXL R12_reg_23_ ( .D(data_in_3[125]), .E(n1353), .CK(clk), .Q(R12[23]) );
  EDFFXL R12_reg_22_ ( .D(data_in_3[124]), .E(n1353), .CK(clk), .Q(R12[22]) );
  EDFFX1 R12_reg_20_ ( .D(data_in_3[122]), .E(n1353), .CK(clk), .Q(R12[20]) );
  EDFFX1 R12_reg_19_ ( .D(data_in_3[121]), .E(n1353), .CK(clk), .Q(R12[19]) );
  EDFFX1 R12_reg_18_ ( .D(data_in_3[120]), .E(n1353), .CK(clk), .Q(R12[18]) );
  EDFFX1 R12_reg_17_ ( .D(data_in_3[119]), .E(n1353), .CK(clk), .Q(R12[17]) );
  EDFFXL R12_reg_12_ ( .D(data_in_3[114]), .E(n1353), .CK(clk), .Q(R12[12]) );
  EDFFXL R12_reg_11_ ( .D(data_in_3[113]), .E(n1354), .CK(clk), .Q(R12[11]) );
  EDFFXL R12_reg_10_ ( .D(data_in_3[112]), .E(n1355), .CK(clk), .Q(R12[10]) );
  EDFFXL R12_reg_9_ ( .D(data_in_3[111]), .E(n1355), .CK(clk), .Q(R12[9]) );
  EDFFXL R12_reg_8_ ( .D(data_in_3[110]), .E(n1355), .CK(clk), .Q(R12[8]) );
  EDFFXL R12_reg_7_ ( .D(data_in_3[109]), .E(n1360), .CK(clk), .Q(R12[7]) );
  EDFFXL R12_reg_6_ ( .D(data_in_3[108]), .E(n1353), .CK(clk), .Q(R12[6]) );
  EDFFXL R12_reg_4_ ( .D(data_in_3[106]), .E(n1361), .CK(clk), .Q(R12[4]) );
  EDFFX1 R12_reg_3_ ( .D(data_in_3[105]), .E(n1353), .CK(clk), .Q(R12[3]) );
  EDFFX1 R12_reg_2_ ( .D(data_in_3[104]), .E(n1361), .CK(clk), .Q(R12[2]) );
  EDFFX1 R12_reg_1_ ( .D(data_in_3[103]), .E(n1360), .CK(clk), .Q(R12[1]) );
  EDFFX1 R12_reg_0_ ( .D(data_in_3[102]), .E(n1353), .CK(clk), .Q(R12[0]) );
  EDFFXL R3_reg_29_ ( .D(data_in_3[29]), .E(n1347), .CK(clk), .Q(R3[29]) );
  EDFFXL R3_reg_28_ ( .D(data_in_3[28]), .E(n1347), .CK(clk), .Q(R3[28]) );
  EDFFXL R3_reg_26_ ( .D(data_in_3[26]), .E(n1346), .CK(clk), .Q(R3[26]) );
  EDFFXL R3_reg_25_ ( .D(data_in_3[25]), .E(n1346), .CK(clk), .Q(R3[25]) );
  EDFFXL R3_reg_24_ ( .D(data_in_3[24]), .E(n1346), .CK(clk), .Q(R3[24]) );
  EDFFXL R3_reg_23_ ( .D(data_in_3[23]), .E(n1346), .CK(clk), .Q(R3[23]) );
  EDFFXL R3_reg_22_ ( .D(data_in_3[22]), .E(n1346), .CK(clk), .Q(R3[22]) );
  EDFFXL R3_reg_21_ ( .D(data_in_3[21]), .E(n1346), .CK(clk), .Q(R3[21]) );
  EDFFX1 R3_reg_19_ ( .D(data_in_3[19]), .E(n1346), .CK(clk), .Q(R3[19]) );
  EDFFX1 R3_reg_18_ ( .D(data_in_3[18]), .E(n1346), .CK(clk), .Q(R3[18]) );
  EDFFX1 R3_reg_17_ ( .D(data_in_3[17]), .E(n1346), .CK(clk), .Q(R3[17]) );
  EDFFXL R3_reg_12_ ( .D(data_in_3[12]), .E(n1345), .CK(clk), .Q(R3[12]) );
  EDFFXL R3_reg_10_ ( .D(data_in_3[10]), .E(n1345), .CK(clk), .Q(R3[10]) );
  EDFFXL R3_reg_9_ ( .D(data_in_3[9]), .E(n1345), .CK(clk), .Q(R3[9]) );
  EDFFXL R3_reg_8_ ( .D(data_in_3[8]), .E(n1345), .CK(clk), .Q(R3[8]) );
  EDFFXL R3_reg_7_ ( .D(data_in_3[7]), .E(n1345), .CK(clk), .Q(R3[7]) );
  EDFFXL R3_reg_6_ ( .D(data_in_3[6]), .E(n1345), .CK(clk), .Q(R3[6]) );
  EDFFXL R3_reg_5_ ( .D(data_in_3[5]), .E(n1345), .CK(clk), .Q(R3[5]) );
  EDFFXL R3_reg_4_ ( .D(data_in_3[4]), .E(n1345), .CK(clk), .Q(R3[4]) );
  EDFFX1 R3_reg_3_ ( .D(data_in_3[3]), .E(n1344), .CK(clk), .Q(R3[3]) );
  EDFFX1 R3_reg_2_ ( .D(data_in_3[2]), .E(n1344), .CK(clk), .Q(R3[2]) );
  EDFFX1 R3_reg_1_ ( .D(data_in_3[1]), .E(n1344), .CK(clk), .Q(R3[1]) );
  EDFFX1 R3_reg_0_ ( .D(data_in_3[0]), .E(n1344), .CK(clk), .Q(R3[0]) );
  EDFFXL R0_reg_29_ ( .D(data_in_3[29]), .E(n1357), .CK(clk), .Q(R0[29]) );
  EDFFXL R0_reg_28_ ( .D(data_in_3[28]), .E(n1356), .CK(clk), .Q(R0[28]) );
  EDFFXL R0_reg_26_ ( .D(data_in_3[26]), .E(n1358), .CK(clk), .Q(R0[26]) );
  EDFFXL R0_reg_25_ ( .D(data_in_3[25]), .E(n1354), .CK(clk), .Q(R0[25]) );
  EDFFXL R0_reg_24_ ( .D(data_in_3[24]), .E(n1356), .CK(clk), .Q(R0[24]) );
  EDFFXL R0_reg_23_ ( .D(data_in_3[23]), .E(n1356), .CK(clk), .Q(R0[23]) );
  EDFFXL R0_reg_22_ ( .D(data_in_3[22]), .E(n1359), .CK(clk), .Q(R0[22]) );
  EDFFXL R0_reg_21_ ( .D(data_in_3[21]), .E(n1354), .CK(clk), .Q(R0[21]) );
  EDFFX1 R0_reg_19_ ( .D(data_in_3[19]), .E(n1355), .CK(clk), .Q(R0[19]) );
  EDFFX1 R0_reg_18_ ( .D(data_in_3[18]), .E(n1354), .CK(clk), .Q(R0[18]) );
  EDFFX1 R0_reg_17_ ( .D(data_in_3[17]), .E(n1361), .CK(clk), .Q(R0[17]) );
  EDFFXL R0_reg_12_ ( .D(data_in_3[12]), .E(n1361), .CK(clk), .Q(R0[12]) );
  EDFFXL R0_reg_10_ ( .D(data_in_3[10]), .E(n1361), .CK(clk), .Q(R0[10]) );
  EDFFXL R0_reg_9_ ( .D(data_in_3[9]), .E(n1361), .CK(clk), .Q(R0[9]) );
  EDFFXL R0_reg_8_ ( .D(data_in_3[8]), .E(n1361), .CK(clk), .Q(R0[8]) );
  EDFFXL R0_reg_7_ ( .D(data_in_3[7]), .E(n1361), .CK(clk), .Q(R0[7]) );
  EDFFXL R0_reg_6_ ( .D(data_in_3[6]), .E(n1361), .CK(clk), .Q(R0[6]) );
  EDFFXL R0_reg_5_ ( .D(data_in_3[5]), .E(n1360), .CK(clk), .Q(R0[5]) );
  EDFFXL R0_reg_4_ ( .D(data_in_3[4]), .E(n1360), .CK(clk), .Q(R0[4]) );
  EDFFX1 R0_reg_3_ ( .D(data_in_3[3]), .E(n1360), .CK(clk), .Q(R0[3]) );
  EDFFX1 R0_reg_2_ ( .D(data_in_3[2]), .E(n1360), .CK(clk), .Q(R0[2]) );
  EDFFX1 R0_reg_1_ ( .D(data_in_3[1]), .E(n1360), .CK(clk), .Q(R0[1]) );
  EDFFX1 R0_reg_0_ ( .D(data_in_3[0]), .E(n1360), .CK(clk), .Q(R0[0]) );
  EDFFXL R1_reg_29_ ( .D(data_in_3[29]), .E(n1371), .CK(clk), .Q(R1[29]) );
  EDFFXL R1_reg_28_ ( .D(data_in_3[28]), .E(n1368), .CK(clk), .Q(R1[28]) );
  EDFFXL R1_reg_26_ ( .D(data_in_3[26]), .E(n1365), .CK(clk), .Q(R1[26]) );
  EDFFXL R1_reg_25_ ( .D(data_in_3[25]), .E(n1367), .CK(clk), .Q(R1[25]) );
  EDFFXL R1_reg_24_ ( .D(data_in_3[24]), .E(n1367), .CK(clk), .Q(R1[24]) );
  EDFFXL R1_reg_23_ ( .D(data_in_3[23]), .E(n1371), .CK(clk), .Q(R1[23]) );
  EDFFXL R1_reg_22_ ( .D(data_in_3[22]), .E(n1367), .CK(clk), .Q(R1[22]) );
  EDFFXL R1_reg_21_ ( .D(data_in_3[21]), .E(n1368), .CK(clk), .Q(R1[21]) );
  EDFFX1 R1_reg_19_ ( .D(data_in_3[19]), .E(n1365), .CK(clk), .Q(R1[19]) );
  EDFFX1 R1_reg_18_ ( .D(data_in_3[18]), .E(n1364), .CK(clk), .Q(R1[18]) );
  EDFFX1 R1_reg_17_ ( .D(data_in_3[17]), .E(n1372), .CK(clk), .Q(R1[17]) );
  EDFFXL R1_reg_12_ ( .D(data_in_3[12]), .E(n1372), .CK(clk), .Q(R1[12]) );
  EDFFXL R1_reg_10_ ( .D(data_in_3[10]), .E(n1372), .CK(clk), .Q(R1[10]) );
  EDFFXL R1_reg_9_ ( .D(data_in_3[9]), .E(n1372), .CK(clk), .Q(R1[9]) );
  EDFFXL R1_reg_8_ ( .D(data_in_3[8]), .E(n1372), .CK(clk), .Q(R1[8]) );
  EDFFXL R1_reg_7_ ( .D(data_in_3[7]), .E(n1372), .CK(clk), .Q(R1[7]) );
  EDFFXL R1_reg_6_ ( .D(data_in_3[6]), .E(n1372), .CK(clk), .Q(R1[6]) );
  EDFFXL R1_reg_5_ ( .D(data_in_3[5]), .E(n1371), .CK(clk), .Q(R1[5]) );
  EDFFXL R1_reg_4_ ( .D(data_in_3[4]), .E(n1371), .CK(clk), .Q(R1[4]) );
  EDFFX1 R1_reg_3_ ( .D(data_in_3[3]), .E(n1371), .CK(clk), .Q(R1[3]) );
  EDFFX1 R1_reg_2_ ( .D(data_in_3[2]), .E(n1371), .CK(clk), .Q(R1[2]) );
  EDFFX1 R1_reg_1_ ( .D(data_in_3[1]), .E(n1371), .CK(clk), .Q(R1[1]) );
  EDFFX1 R1_reg_0_ ( .D(data_in_3[0]), .E(n1371), .CK(clk), .Q(R1[0]) );
  EDFFXL R14_reg_29_ ( .D(data_in_3[131]), .E(n1381), .CK(clk), .Q(R14[29]) );
  EDFFXL R14_reg_27_ ( .D(data_in_3[129]), .E(n1382), .CK(clk), .Q(R14[27]) );
  EDFFXL R14_reg_26_ ( .D(data_in_3[128]), .E(n1382), .CK(clk), .Q(R14[26]) );
  EDFFXL R14_reg_25_ ( .D(data_in_3[127]), .E(n1382), .CK(clk), .Q(R14[25]) );
  EDFFXL R14_reg_23_ ( .D(data_in_3[125]), .E(n1382), .CK(clk), .Q(R14[23]) );
  EDFFXL R14_reg_22_ ( .D(data_in_3[124]), .E(n1382), .CK(clk), .Q(R14[22]) );
  EDFFX1 R14_reg_20_ ( .D(data_in_3[122]), .E(n1382), .CK(clk), .Q(R14[20]) );
  EDFFX1 R14_reg_19_ ( .D(data_in_3[121]), .E(n1382), .CK(clk), .Q(R14[19]) );
  EDFFX1 R14_reg_18_ ( .D(data_in_3[120]), .E(n1382), .CK(clk), .Q(R14[18]) );
  EDFFX1 R14_reg_17_ ( .D(data_in_3[119]), .E(n1382), .CK(clk), .Q(R14[17]) );
  EDFFXL R14_reg_12_ ( .D(data_in_3[114]), .E(n1381), .CK(clk), .Q(R14[12]) );
  EDFFXL R14_reg_11_ ( .D(data_in_3[113]), .E(n1381), .CK(clk), .Q(R14[11]) );
  EDFFXL R14_reg_10_ ( .D(data_in_3[112]), .E(n1381), .CK(clk), .Q(R14[10]) );
  EDFFXL R14_reg_9_ ( .D(data_in_3[111]), .E(n1381), .CK(clk), .Q(R14[9]) );
  EDFFXL R14_reg_8_ ( .D(data_in_3[110]), .E(n1381), .CK(clk), .Q(R14[8]) );
  EDFFXL R14_reg_7_ ( .D(data_in_3[109]), .E(n1381), .CK(clk), .Q(R14[7]) );
  EDFFXL R14_reg_6_ ( .D(data_in_3[108]), .E(n1381), .CK(clk), .Q(R14[6]) );
  EDFFXL R14_reg_4_ ( .D(data_in_3[106]), .E(n1381), .CK(clk), .Q(R14[4]) );
  EDFFX1 R14_reg_3_ ( .D(data_in_3[105]), .E(n1380), .CK(clk), .Q(R14[3]) );
  EDFFX1 R14_reg_2_ ( .D(data_in_3[104]), .E(n1380), .CK(clk), .Q(R14[2]) );
  EDFFX1 R14_reg_1_ ( .D(data_in_3[103]), .E(n1380), .CK(clk), .Q(R14[1]) );
  EDFFX1 R14_reg_0_ ( .D(data_in_3[102]), .E(n1380), .CK(clk), .Q(R14[0]) );
  EDFFXL R13_reg_29_ ( .D(data_in_3[131]), .E(n1365), .CK(clk), .Q(R13[29]) );
  EDFFXL R13_reg_27_ ( .D(data_in_3[129]), .E(n1365), .CK(clk), .Q(R13[27]) );
  EDFFXL R13_reg_26_ ( .D(data_in_3[128]), .E(n1365), .CK(clk), .Q(R13[26]) );
  EDFFXL R13_reg_25_ ( .D(data_in_3[127]), .E(n1365), .CK(clk), .Q(R13[25]) );
  EDFFXL R13_reg_23_ ( .D(data_in_3[125]), .E(n1364), .CK(clk), .Q(R13[23]) );
  EDFFXL R13_reg_22_ ( .D(data_in_3[124]), .E(n1364), .CK(clk), .Q(R13[22]) );
  EDFFXL R13_reg_21_ ( .D(data_in_3[123]), .E(n1364), .CK(clk), .Q(R13[21]) );
  EDFFX1 R13_reg_20_ ( .D(data_in_3[122]), .E(n1364), .CK(clk), .Q(R13[20]) );
  EDFFX1 R13_reg_19_ ( .D(data_in_3[121]), .E(n1364), .CK(clk), .Q(R13[19]) );
  EDFFX1 R13_reg_18_ ( .D(data_in_3[120]), .E(n1364), .CK(clk), .Q(R13[18]) );
  EDFFX1 R13_reg_17_ ( .D(data_in_3[119]), .E(n1364), .CK(clk), .Q(R13[17]) );
  EDFFXL R13_reg_12_ ( .D(data_in_3[114]), .E(n1364), .CK(clk), .Q(R13[12]) );
  EDFFXL R13_reg_11_ ( .D(data_in_3[113]), .E(n1371), .CK(clk), .Q(R13[11]) );
  EDFFXL R13_reg_10_ ( .D(data_in_3[112]), .E(n1364), .CK(clk), .Q(R13[10]) );
  EDFFXL R13_reg_9_ ( .D(data_in_3[111]), .E(n1368), .CK(clk), .Q(R13[9]) );
  EDFFXL R13_reg_8_ ( .D(data_in_3[110]), .E(n1370), .CK(clk), .Q(R13[8]) );
  EDFFXL R13_reg_7_ ( .D(data_in_3[109]), .E(n1366), .CK(clk), .Q(R13[7]) );
  EDFFXL R13_reg_6_ ( .D(data_in_3[108]), .E(n1372), .CK(clk), .Q(R13[6]) );
  EDFFXL R13_reg_4_ ( .D(data_in_3[106]), .E(n1369), .CK(clk), .Q(R13[4]) );
  EDFFX1 R13_reg_3_ ( .D(data_in_3[105]), .E(n1366), .CK(clk), .Q(R13[3]) );
  EDFFX1 R13_reg_2_ ( .D(data_in_3[104]), .E(n1372), .CK(clk), .Q(R13[2]) );
  EDFFX1 R13_reg_1_ ( .D(data_in_3[103]), .E(n1370), .CK(clk), .Q(R13[1]) );
  EDFFX1 R13_reg_0_ ( .D(data_in_3[102]), .E(n1366), .CK(clk), .Q(R13[0]) );
  EDFFXL R2_reg_29_ ( .D(data_in_3[29]), .E(n1383), .CK(clk), .Q(R2[29]) );
  EDFFXL R2_reg_28_ ( .D(data_in_3[28]), .E(n1377), .CK(clk), .Q(R2[28]) );
  EDFFXL R2_reg_26_ ( .D(data_in_3[26]), .E(n1375), .CK(clk), .Q(R2[26]) );
  EDFFXL R2_reg_25_ ( .D(data_in_3[25]), .E(n1383), .CK(clk), .Q(R2[25]) );
  EDFFXL R2_reg_24_ ( .D(data_in_3[24]), .E(n1383), .CK(clk), .Q(R2[24]) );
  EDFFXL R2_reg_23_ ( .D(data_in_3[23]), .E(n1383), .CK(clk), .Q(R2[23]) );
  EDFFXL R2_reg_22_ ( .D(data_in_3[22]), .E(n1383), .CK(clk), .Q(R2[22]) );
  EDFFXL R2_reg_21_ ( .D(data_in_3[21]), .E(n1383), .CK(clk), .Q(R2[21]) );
  EDFFX1 R2_reg_19_ ( .D(data_in_3[19]), .E(n1383), .CK(clk), .Q(R2[19]) );
  EDFFX1 R2_reg_18_ ( .D(data_in_3[18]), .E(n1383), .CK(clk), .Q(R2[18]) );
  EDFFX1 R2_reg_17_ ( .D(data_in_3[17]), .E(n1381), .CK(clk), .Q(R2[17]) );
  EDFFXL R2_reg_12_ ( .D(data_in_3[12]), .E(n1380), .CK(clk), .Q(R2[12]) );
  EDFFXL R2_reg_10_ ( .D(data_in_3[10]), .E(n1378), .CK(clk), .Q(R2[10]) );
  EDFFXL R2_reg_9_ ( .D(data_in_3[9]), .E(n1377), .CK(clk), .Q(R2[9]) );
  EDFFXL R2_reg_8_ ( .D(data_in_3[8]), .E(n1381), .CK(clk), .Q(R2[8]) );
  EDFFXL R2_reg_7_ ( .D(data_in_3[7]), .E(n1375), .CK(clk), .Q(R2[7]) );
  EDFFXL R2_reg_6_ ( .D(data_in_3[6]), .E(n1376), .CK(clk), .Q(R2[6]) );
  EDFFXL R2_reg_5_ ( .D(data_in_3[5]), .E(n1382), .CK(clk), .Q(R2[5]) );
  EDFFXL R2_reg_4_ ( .D(data_in_3[4]), .E(n1380), .CK(clk), .Q(R2[4]) );
  EDFFX1 R2_reg_3_ ( .D(data_in_3[3]), .E(n1378), .CK(clk), .Q(R2[3]) );
  EDFFX1 R2_reg_2_ ( .D(data_in_3[2]), .E(n1382), .CK(clk), .Q(R2[2]) );
  EDFFX1 R2_reg_1_ ( .D(data_in_3[1]), .E(n1377), .CK(clk), .Q(R2[1]) );
  EDFFX1 R2_reg_0_ ( .D(data_in_3[0]), .E(n1375), .CK(clk), .Q(R2[0]) );
  JKFFRXL counter_1_reg_0_ ( .J(1'b1), .K(1'b1), .CK(clk), .RN(rst_n), .Q(
        counter_1[0]), .QN(n584) );
  JKFFRXL counter_2_reg_0_ ( .J(1'b1), .K(1'b1), .CK(clk), .RN(rst_n), .Q(
        counter_2[0]), .QN(n861) );
  DFFRHQX1 counter_2_reg_1_ ( .D(N50), .CK(clk), .RN(rst_n), .Q(counter_2[1])
         );
  DFFRHQX1 counter_1_reg_1_ ( .D(N26), .CK(clk), .RN(rst_n), .Q(counter_1[1])
         );
  DFFRHQX1 counter_2_reg_2_ ( .D(n1388), .CK(clk), .RN(rst_n), .Q(counter_2[2]) );
  DFFRHQX1 counter_2_reg_3_ ( .D(N52), .CK(clk), .RN(rst_n), .Q(counter_2[3])
         );
  EDFFX1 data_out_3_reg_33_ ( .D(N152), .E(n1386), .CK(clk), .Q(data_out_3[33]) );
  EDFFX1 data_out_3_reg_32_ ( .D(N151), .E(n1386), .CK(clk), .Q(data_out_3[32]) );
  EDFFX1 data_out_3_reg_31_ ( .D(N150), .E(n1386), .CK(clk), .Q(data_out_3[31]) );
  EDFFX1 data_out_3_reg_30_ ( .D(N149), .E(n1386), .CK(clk), .Q(data_out_3[30]) );
  EDFFX1 data_out_3_reg_29_ ( .D(N148), .E(n1386), .CK(clk), .Q(data_out_3[29]) );
  EDFFX1 data_out_3_reg_28_ ( .D(N147), .E(n1386), .CK(clk), .Q(data_out_3[28]) );
  EDFFX1 data_out_3_reg_27_ ( .D(N146), .E(n1386), .CK(clk), .Q(data_out_3[27]) );
  EDFFX1 data_out_3_reg_26_ ( .D(N145), .E(n1386), .CK(clk), .Q(data_out_3[26]) );
  EDFFX1 data_out_3_reg_25_ ( .D(N144), .E(n1386), .CK(clk), .Q(data_out_3[25]) );
  EDFFX1 data_out_3_reg_24_ ( .D(N143), .E(n1386), .CK(clk), .Q(data_out_3[24]) );
  EDFFX1 data_out_3_reg_23_ ( .D(N142), .E(n1386), .CK(clk), .Q(data_out_3[23]) );
  EDFFX1 data_out_3_reg_22_ ( .D(N141), .E(n1386), .CK(clk), .Q(data_out_3[22]) );
  EDFFX1 data_out_3_reg_21_ ( .D(N140), .E(n1386), .CK(clk), .Q(data_out_3[21]) );
  EDFFX1 data_out_3_reg_20_ ( .D(N139), .E(n1386), .CK(clk), .Q(data_out_3[20]) );
  EDFFX1 data_out_3_reg_19_ ( .D(N138), .E(n1386), .CK(clk), .Q(data_out_3[19]) );
  EDFFX1 data_out_3_reg_18_ ( .D(N137), .E(n1386), .CK(clk), .Q(data_out_3[18]) );
  EDFFX1 data_out_3_reg_17_ ( .D(N136), .E(n1386), .CK(clk), .Q(data_out_3[17]) );
  EDFFX1 data_out_3_reg_16_ ( .D(N135), .E(n1386), .CK(clk), .Q(data_out_3[16]) );
  EDFFX1 data_out_3_reg_15_ ( .D(N134), .E(n1386), .CK(clk), .Q(data_out_3[15]) );
  EDFFX1 data_out_3_reg_14_ ( .D(N133), .E(n1386), .CK(clk), .Q(data_out_3[14]) );
  EDFFX1 data_out_3_reg_13_ ( .D(N132), .E(n1386), .CK(clk), .Q(data_out_3[13]) );
  EDFFX1 data_out_3_reg_12_ ( .D(N131), .E(n1386), .CK(clk), .Q(data_out_3[12]) );
  EDFFX1 data_out_3_reg_11_ ( .D(N130), .E(n1386), .CK(clk), .Q(data_out_3[11]) );
  EDFFX1 data_out_3_reg_10_ ( .D(N129), .E(n1386), .CK(clk), .Q(data_out_3[10]) );
  EDFFX1 data_out_3_reg_9_ ( .D(N128), .E(n1386), .CK(clk), .Q(data_out_3[9])
         );
  EDFFX1 data_out_3_reg_8_ ( .D(N127), .E(n1386), .CK(clk), .Q(data_out_3[8])
         );
  EDFFX1 data_out_3_reg_7_ ( .D(N126), .E(n1386), .CK(clk), .Q(data_out_3[7])
         );
  EDFFX1 data_out_3_reg_6_ ( .D(N125), .E(n1386), .CK(clk), .Q(data_out_3[6])
         );
  EDFFX1 data_out_3_reg_5_ ( .D(N124), .E(n1386), .CK(clk), .Q(data_out_3[5])
         );
  EDFFX1 data_out_3_reg_4_ ( .D(N123), .E(n1386), .CK(clk), .Q(data_out_3[4])
         );
  EDFFX1 data_out_3_reg_3_ ( .D(N122), .E(n1386), .CK(clk), .Q(data_out_3[3])
         );
  EDFFX1 data_out_3_reg_2_ ( .D(N121), .E(n1386), .CK(clk), .Q(data_out_3[2])
         );
  EDFFX1 data_out_3_reg_1_ ( .D(N120), .E(n1386), .CK(clk), .Q(data_out_3[1])
         );
  EDFFX1 data_out_3_reg_0_ ( .D(N119), .E(n1386), .CK(clk), .Q(data_out_3[0])
         );
  EDFFXL R2_reg_20_ ( .D(data_in_3[20]), .E(n1383), .CK(clk), .Q(R2[20]) );
  EDFFXL R3_reg_20_ ( .D(data_in_3[20]), .E(n1346), .CK(clk), .Q(R3[20]) );
  EDFFXL R0_reg_20_ ( .D(data_in_3[20]), .E(n1355), .CK(clk), .Q(R0[20]) );
  EDFFXL R1_reg_20_ ( .D(data_in_3[20]), .E(n1367), .CK(clk), .Q(R1[20]) );
  EDFFXL R4_reg_8_ ( .D(data_in_3[42]), .E(n1358), .CK(clk), .QN(n746) );
  EDFFXL R7_reg_29_ ( .D(data_in_3[63]), .E(n19), .CK(clk), .QN(n589) );
  EDFFXL R6_reg_29_ ( .D(data_in_3[63]), .E(n1377), .CK(clk), .QN(n657) );
  EDFFXL R4_reg_29_ ( .D(data_in_3[63]), .E(n1360), .CK(clk), .QN(n725) );
  EDFFXL R7_reg_30_ ( .D(data_in_3[64]), .E(n19), .CK(clk), .QN(n588) );
  EDFFXL R6_reg_30_ ( .D(data_in_3[64]), .E(n1377), .CK(clk), .QN(n656) );
  EDFFXL R4_reg_30_ ( .D(data_in_3[64]), .E(n1360), .CK(clk), .QN(n724) );
  EDFFX1 R13_reg_24_ ( .D(data_in_3[126]), .E(n1365), .CK(clk), .Q(R13[24]) );
  EDFFX1 R14_reg_24_ ( .D(data_in_3[126]), .E(n1382), .CK(clk), .Q(R14[24]) );
  EDFFX1 R12_reg_24_ ( .D(data_in_3[126]), .E(n1354), .CK(clk), .Q(R12[24]) );
  EDFFX1 R15_reg_24_ ( .D(data_in_3[126]), .E(n1342), .CK(clk), .Q(R15[24]) );
  EDFFXL R4_reg_5_ ( .D(n83), .E(n1358), .CK(clk), .QN(n749) );
  EDFFXL R6_reg_5_ ( .D(n83), .E(n1375), .CK(clk), .QN(n681) );
  EDFFXL R7_reg_5_ ( .D(n83), .E(n1347), .CK(clk), .QN(n613) );
  EDFFXL R4_reg_25_ ( .D(data_in_3[59]), .E(n1359), .CK(clk), .QN(n729) );
  EDFFXL R6_reg_25_ ( .D(data_in_3[59]), .E(n1377), .CK(clk), .QN(n661) );
  EDFFXL R7_reg_25_ ( .D(data_in_3[59]), .E(n1348), .CK(clk), .QN(n593) );
  EDFFXL R7_reg_4_ ( .D(data_in_3[38]), .E(n1347), .CK(clk), .QN(n614) );
  EDFFXL R6_reg_4_ ( .D(data_in_3[38]), .E(n1375), .CK(clk), .QN(n682) );
  EDFFXL R4_reg_4_ ( .D(data_in_3[38]), .E(n1358), .CK(clk), .QN(n750) );
  EDFFXL R7_reg_24_ ( .D(data_in_3[58]), .E(n19), .CK(clk), .QN(n594) );
  EDFFXL R6_reg_24_ ( .D(data_in_3[58]), .E(n1377), .CK(clk), .QN(n662) );
  EDFFXL R4_reg_24_ ( .D(data_in_3[58]), .E(n1359), .CK(clk), .QN(n730) );
  EDFFXL R11_reg_22_ ( .D(data_in_3[90]), .E(n19), .CK(clk), .QN(n698) );
  EDFFXL R10_reg_22_ ( .D(data_in_3[90]), .E(n1374), .CK(clk), .QN(n630) );
  EDFFXL R9_reg_22_ ( .D(data_in_3[90]), .E(n1372), .CK(clk), .QN(n834) );
  EDFFXL R8_reg_22_ ( .D(data_in_3[90]), .E(n1352), .CK(clk), .QN(n766) );
  EDFFXL R11_reg_5_ ( .D(data_in_3[73]), .E(n19), .CK(clk), .QN(n715) );
  EDFFXL R10_reg_5_ ( .D(data_in_3[73]), .E(n1374), .CK(clk), .QN(n647) );
  EDFFXL R9_reg_5_ ( .D(data_in_3[73]), .E(n1370), .CK(clk), .QN(n851) );
  EDFFXL R8_reg_5_ ( .D(data_in_3[73]), .E(n1352), .CK(clk), .QN(n783) );
  EDFFXL R11_reg_23_ ( .D(data_in_3[91]), .E(n19), .CK(clk), .QN(n697) );
  EDFFXL R10_reg_23_ ( .D(data_in_3[91]), .E(n1374), .CK(clk), .QN(n629) );
  EDFFXL R9_reg_23_ ( .D(data_in_3[91]), .E(n1366), .CK(clk), .QN(n833) );
  EDFFXL R8_reg_23_ ( .D(data_in_3[91]), .E(n1352), .CK(clk), .QN(n765) );
  EDFFXL R6_reg_26_ ( .D(data_in_3[60]), .E(n1374), .CK(clk), .QN(n660) );
  EDFFXL R5_reg_26_ ( .D(data_in_3[60]), .E(n1366), .CK(clk), .QN(n796) );
  EDFFXL R4_reg_26_ ( .D(data_in_3[60]), .E(n1361), .CK(clk), .QN(n728) );
  EDFFXL R11_reg_6_ ( .D(data_in_3[74]), .E(n19), .CK(clk), .QN(n714) );
  EDFFXL R10_reg_6_ ( .D(data_in_3[74]), .E(n1374), .CK(clk), .QN(n646) );
  EDFFXL R9_reg_6_ ( .D(data_in_3[74]), .E(n1369), .CK(clk), .QN(n850) );
  EDFFXL R8_reg_6_ ( .D(data_in_3[74]), .E(n1352), .CK(clk), .QN(n782) );
  EDFFXL R5_reg_23_ ( .D(data_in_3[57]), .E(n1370), .CK(clk), .QN(n799) );
  EDFFXL R11_reg_8_ ( .D(data_in_3[76]), .E(n19), .CK(clk), .QN(n712) );
  EDFFXL R10_reg_8_ ( .D(data_in_3[76]), .E(n1374), .CK(clk), .QN(n644) );
  EDFFXL R9_reg_8_ ( .D(data_in_3[76]), .E(n1369), .CK(clk), .QN(n848) );
  EDFFXL R8_reg_8_ ( .D(data_in_3[76]), .E(n1352), .CK(clk), .QN(n780) );
  EDFFXL R5_reg_7_ ( .D(data_in_3[41]), .E(n1367), .CK(clk), .QN(n815) );
  EDFFXL R5_reg_10_ ( .D(data_in_3[44]), .E(n1369), .CK(clk), .QN(n812) );
  EDFFXL R7_reg_27_ ( .D(data_in_3[61]), .E(n1341), .CK(clk), .QN(n591) );
  EDFFXL R6_reg_27_ ( .D(data_in_3[61]), .E(n1374), .CK(clk), .QN(n659) );
  EDFFXL R5_reg_27_ ( .D(data_in_3[61]), .E(n1366), .CK(clk), .QN(n795) );
  EDFFXL R4_reg_27_ ( .D(data_in_3[61]), .E(n1360), .CK(clk), .QN(n727) );
  EDFFXL R5_reg_22_ ( .D(data_in_3[56]), .E(n1370), .CK(clk), .QN(n800) );
  EDFFXL R7_reg_6_ ( .D(data_in_3[40]), .E(n1343), .CK(clk), .QN(n612) );
  EDFFXL R6_reg_6_ ( .D(data_in_3[40]), .E(n1374), .CK(clk), .QN(n680) );
  EDFFXL R5_reg_6_ ( .D(data_in_3[40]), .E(n1370), .CK(clk), .QN(n816) );
  EDFFXL R4_reg_6_ ( .D(data_in_3[40]), .E(n1353), .CK(clk), .QN(n748) );
  EDFFXL R7_reg_26_ ( .D(data_in_3[60]), .E(n1343), .CK(clk), .QN(n592) );
  EDFFXL R7_reg_8_ ( .D(data_in_3[42]), .E(n1343), .CK(clk), .QN(n610) );
  EDFFXL R6_reg_8_ ( .D(data_in_3[42]), .E(n1374), .CK(clk), .QN(n678) );
  EDFFXL R7_reg_12_ ( .D(data_in_3[46]), .E(n1348), .CK(clk), .QN(n606) );
  JKFFRX2 p_s_flag_out_reg ( .J(n1391), .K(1'b0), .CK(clk), .RN(rst_n), .Q(
        n1386) );
  EDFFX1 R2_reg_27_ ( .D(data_in_3[27]), .E(n1383), .CK(clk), .Q(R2[27]) );
  EDFFX1 R1_reg_27_ ( .D(data_in_3[27]), .E(n1364), .CK(clk), .Q(R1[27]) );
  EDFFX1 R0_reg_27_ ( .D(data_in_3[27]), .E(n1359), .CK(clk), .Q(R0[27]) );
  EDFFX1 R3_reg_27_ ( .D(data_in_3[27]), .E(n1346), .CK(clk), .Q(R3[27]) );
  EDFFX1 R13_reg_5_ ( .D(data_in_3[107]), .E(n1370), .CK(clk), .Q(R13[5]) );
  EDFFX1 R14_reg_5_ ( .D(data_in_3[107]), .E(n1381), .CK(clk), .Q(R14[5]) );
  EDFFX1 R12_reg_5_ ( .D(data_in_3[107]), .E(n1360), .CK(clk), .Q(R12[5]) );
  EDFFX1 R15_reg_5_ ( .D(data_in_3[107]), .E(n19), .CK(clk), .Q(R15[5]) );
  EDFFX1 R8_reg_21_ ( .D(data_in_3[89]), .E(n1352), .CK(clk), .QN(n767) );
  EDFFX1 R9_reg_21_ ( .D(data_in_3[89]), .E(n1369), .CK(clk), .QN(n835) );
  EDFFX1 R10_reg_21_ ( .D(data_in_3[89]), .E(n1374), .CK(clk), .QN(n631) );
  EDFFX1 R11_reg_21_ ( .D(data_in_3[89]), .E(n19), .CK(clk), .QN(n699) );
  EDFFX1 R14_reg_21_ ( .D(data_in_3[123]), .E(n1382), .CK(clk), .Q(R14[21]) );
  EDFFX1 R12_reg_21_ ( .D(data_in_3[123]), .E(n1353), .CK(clk), .Q(R12[21]) );
  EDFFX1 R15_reg_21_ ( .D(data_in_3[123]), .E(n1341), .CK(clk), .Q(R15[21]) );
  MX2X1 U3 ( .A(data_in_3[48]), .B(n256), .S0(n1362), .Y(n1251) );
  MX2X1 U6 ( .A(data_in_3[48]), .B(n528), .S0(n1349), .Y(n1257) );
  MX2X1 U7 ( .A(data_in_3[100]), .B(n444), .S0(n1385), .Y(n1267) );
  MX2X1 U8 ( .A(data_in_3[100]), .B(n104), .S0(n1373), .Y(n1266) );
  MX2X2 U9 ( .A(R12[30]), .B(data_in_3[132]), .S0(n1354), .Y(n859) );
  MX2X2 U10 ( .A(data_in_3[33]), .B(R2[33]), .S0(n153), .Y(n1219) );
  MX2X2 U11 ( .A(n392), .B(data_in_3[48]), .S0(n1376), .Y(n1255) );
  MX2X1 U12 ( .A(data_in_3[65]), .B(n137), .S0(n1373), .Y(n1270) );
  MX2X2 U13 ( .A(R14[13]), .B(data_in_3[115]), .S0(n1381), .Y(n549) );
  MX2X2 U14 ( .A(n273), .B(data_in_3[65]), .S0(n1360), .Y(n1269) );
  MX2X2 U15 ( .A(R12[15]), .B(data_in_3[117]), .S0(n1353), .Y(n513) );
  MX2X2 U16 ( .A(R12[13]), .B(data_in_3[115]), .S0(n1353), .Y(n541) );
  NAND2X2 U17 ( .A(n120), .B(n8), .Y(n9) );
  NAND2X1 U18 ( .A(data_in_3[48]), .B(n1369), .Y(n10) );
  NAND2X2 U19 ( .A(n9), .B(n10), .Y(n1253) );
  INVX1 U20 ( .A(n1369), .Y(n8) );
  INVX20 U21 ( .A(n151), .Y(n1369) );
  MX2X1 U22 ( .A(R15[33]), .B(data_in_3[135]), .S0(n1342), .Y(n539) );
  MX2X1 U23 ( .A(R13[30]), .B(data_in_3[132]), .S0(n1365), .Y(n862) );
  MX2X1 U24 ( .A(R14[30]), .B(data_in_3[132]), .S0(n1379), .Y(n864) );
  MX2X1 U25 ( .A(R15[30]), .B(data_in_3[132]), .S0(n1342), .Y(n866) );
  MX2X1 U26 ( .A(R12[31]), .B(data_in_3[133]), .S0(n1354), .Y(n1183) );
  MX2X1 U27 ( .A(R1[14]), .B(data_in_3[14]), .S0(n1372), .Y(n1201) );
  MX2X1 U28 ( .A(n253), .B(data_in_3[45]), .S0(n1358), .Y(n1226) );
  MX2X1 U29 ( .A(n357), .B(data_in_3[81]), .S0(n1347), .Y(n1237) );
  INVX1 U30 ( .A(n1376), .Y(n71) );
  MX2X2 U31 ( .A(n443), .B(data_in_3[99]), .S0(n1380), .Y(n1259) );
  INVX1 U32 ( .A(n1344), .Y(n98) );
  MX2X1 U33 ( .A(data_in_3[98]), .B(n442), .S0(n1385), .Y(n1263) );
  MX2X1 U34 ( .A(n374), .B(data_in_3[98]), .S0(n1344), .Y(n1264) );
  NOR3X2 U35 ( .A(counter_1[1]), .B(p_s_flag_in), .C(n584), .Y(n19) );
  INVX1 U36 ( .A(n1348), .Y(n81) );
  AND2X2 U37 ( .A(n1162), .B(n872), .Y(n20) );
  NAND2X1 U38 ( .A(n1158), .B(n871), .Y(n21) );
  NAND2X1 U39 ( .A(n1158), .B(n869), .Y(n22) );
  NAND2X1 U40 ( .A(n871), .B(n1163), .Y(n23) );
  NAND2X1 U41 ( .A(n1157), .B(n871), .Y(n24) );
  NAND2X1 U42 ( .A(n1162), .B(n871), .Y(n25) );
  NAND2X1 U43 ( .A(n1162), .B(n869), .Y(n26) );
  MX2X1 U45 ( .A(data_in_3[49]), .B(n257), .S0(n1362), .Y(n1252) );
  MX2X1 U46 ( .A(R14[15]), .B(data_in_3[117]), .S0(n1381), .Y(n521) );
  MX2X1 U47 ( .A(n411), .B(data_in_3[67]), .S0(n1377), .Y(n1224) );
  MX2X1 U48 ( .A(data_in_3[100]), .B(n376), .S0(n1351), .Y(n1268) );
  MX2X1 U49 ( .A(data_in_3[30]), .B(R3[30]), .S0(n1350), .Y(n1173) );
  MX2X1 U50 ( .A(data_in_3[116]), .B(R14[14]), .S0(n1384), .Y(n519) );
  MX2X1 U51 ( .A(n377), .B(data_in_3[101]), .S0(n1344), .Y(n1233) );
  MX2X2 U52 ( .A(data_in_3[31]), .B(R3[31]), .S0(n81), .Y(n575) );
  MX2X1 U53 ( .A(data_in_3[134]), .B(R12[32]), .S0(n1363), .Y(n881) );
  MX2X1 U54 ( .A(R14[32]), .B(data_in_3[134]), .S0(n1378), .Y(n893) );
  MX2X2 U55 ( .A(R0[31]), .B(data_in_3[31]), .S0(n1356), .Y(n569) );
  MX2X2 U56 ( .A(R1[31]), .B(data_in_3[31]), .S0(n1367), .Y(n571) );
  MX2X2 U57 ( .A(R2[31]), .B(data_in_3[31]), .S0(n1383), .Y(n573) );
  MX2X2 U58 ( .A(data_in_3[47]), .B(n391), .S0(n71), .Y(n1238) );
  MX2X2 U59 ( .A(n222), .B(data_in_3[82]), .S0(n1356), .Y(n1293) );
  MX2X2 U60 ( .A(n426), .B(data_in_3[82]), .S0(n1379), .Y(n1295) );
  MX2X2 U61 ( .A(n358), .B(data_in_3[82]), .S0(n1343), .Y(n1296) );
  MX2X2 U62 ( .A(n86), .B(data_in_3[82]), .S0(n1367), .Y(n1294) );
  MX2X2 U63 ( .A(R0[33]), .B(data_in_3[33]), .S0(n1358), .Y(n1215) );
  MX2X2 U64 ( .A(R1[33]), .B(data_in_3[33]), .S0(n1369), .Y(n1217) );
  MX2X2 U65 ( .A(data_in_3[33]), .B(R3[33]), .S0(n1349), .Y(n1221) );
  MX2X2 U66 ( .A(R1[13]), .B(data_in_3[13]), .S0(n1372), .Y(n1193) );
  MX2X2 U67 ( .A(R3[13]), .B(data_in_3[13]), .S0(n1345), .Y(n1197) );
  MX2X2 U68 ( .A(R0[13]), .B(data_in_3[13]), .S0(n1361), .Y(n1191) );
  MX2X2 U69 ( .A(R2[13]), .B(data_in_3[13]), .S0(n1378), .Y(n1195) );
  MX2X2 U70 ( .A(R0[15]), .B(data_in_3[15]), .S0(n1361), .Y(n577) );
  MX2X2 U71 ( .A(R1[15]), .B(data_in_3[15]), .S0(n1372), .Y(n579) );
  MX2X2 U72 ( .A(R3[32]), .B(data_in_3[32]), .S0(n1347), .Y(n567) );
  MX2X2 U73 ( .A(R0[32]), .B(data_in_3[32]), .S0(n1359), .Y(n561) );
  MX2X2 U74 ( .A(R1[32]), .B(data_in_3[32]), .S0(n1370), .Y(n563) );
  MX2X2 U75 ( .A(R2[32]), .B(data_in_3[32]), .S0(n1383), .Y(n565) );
  INVX4 U76 ( .A(n82), .Y(n83) );
  INVX4 U77 ( .A(data_in_3[39]), .Y(n82) );
  MX2X2 U78 ( .A(R2[15]), .B(data_in_3[15]), .S0(n1379), .Y(n581) );
  MX2X1 U79 ( .A(data_in_3[50]), .B(n530), .S0(n1349), .Y(n1280) );
  MX2X2 U80 ( .A(data_in_3[47]), .B(n527), .S0(n81), .Y(n1239) );
  MX2X2 U81 ( .A(data_in_3[99]), .B(n375), .S0(n98), .Y(n1260) );
  MX2X1 U82 ( .A(n275), .B(data_in_3[67]), .S0(n1360), .Y(n1222) );
  MX2X1 U83 ( .A(n139), .B(data_in_3[67]), .S0(n1371), .Y(n1223) );
  MX2X2 U84 ( .A(R3[15]), .B(data_in_3[15]), .S0(n1345), .Y(n857) );
  INVX1 U85 ( .A(n867), .Y(n1309) );
  INVX1 U86 ( .A(n867), .Y(n1310) );
  INVX1 U87 ( .A(n22), .Y(n1328) );
  INVX1 U88 ( .A(n24), .Y(n1334) );
  INVX1 U89 ( .A(n25), .Y(n1318) );
  INVX1 U90 ( .A(n26), .Y(n1312) );
  INVX1 U91 ( .A(n21), .Y(n1336) );
  INVX1 U92 ( .A(n23), .Y(n1320) );
  INVX1 U93 ( .A(n1326), .Y(n1325) );
  INVX1 U94 ( .A(n1340), .Y(n1339) );
  INVX1 U95 ( .A(n1332), .Y(n1331) );
  INVX1 U96 ( .A(n1324), .Y(n1323) );
  INVX1 U97 ( .A(n1316), .Y(n1315) );
  INVX1 U98 ( .A(n20), .Y(n1314) );
  INVX1 U99 ( .A(n1338), .Y(n1337) );
  INVX1 U100 ( .A(n1330), .Y(n1329) );
  INVX1 U101 ( .A(n1322), .Y(n1321) );
  INVX1 U102 ( .A(n151), .Y(n1366) );
  INVX1 U103 ( .A(n151), .Y(n1370) );
  INVX1 U104 ( .A(n1363), .Y(n1355) );
  INVX1 U105 ( .A(n1362), .Y(n1359) );
  INVX1 U106 ( .A(n1385), .Y(n1378) );
  INVX1 U107 ( .A(n1384), .Y(n1382) );
  INVX1 U108 ( .A(n1385), .Y(n1375) );
  INVX1 U109 ( .A(n1384), .Y(n1381) );
  INVX1 U110 ( .A(n1373), .Y(n1364) );
  INVX1 U111 ( .A(n151), .Y(n1367) );
  INVX1 U112 ( .A(n1373), .Y(n1371) );
  INVX1 U113 ( .A(n152), .Y(n1353) );
  INVX1 U114 ( .A(n1362), .Y(n1356) );
  INVX1 U115 ( .A(n152), .Y(n1360) );
  INVX1 U116 ( .A(n1351), .Y(n1341) );
  INVX1 U117 ( .A(n1351), .Y(n1343) );
  INVX1 U118 ( .A(n1385), .Y(n1377) );
  INVX1 U119 ( .A(n1385), .Y(n1379) );
  INVX1 U120 ( .A(n1385), .Y(n1380) );
  INVX1 U121 ( .A(n1351), .Y(n1344) );
  INVX1 U122 ( .A(n1350), .Y(n1345) );
  INVX1 U123 ( .A(n1349), .Y(n1347) );
  INVX1 U124 ( .A(n1373), .Y(n1365) );
  INVX1 U125 ( .A(n1363), .Y(n1354) );
  INVX1 U126 ( .A(n1351), .Y(n1342) );
  INVX1 U127 ( .A(n1384), .Y(n1376) );
  INVX1 U128 ( .A(n1350), .Y(n1346) );
  INVX1 U129 ( .A(n1349), .Y(n1348) );
  INVX1 U130 ( .A(n1373), .Y(n1368) );
  INVX1 U131 ( .A(n1362), .Y(n1357) );
  INVX1 U132 ( .A(n151), .Y(n1372) );
  INVX1 U133 ( .A(n152), .Y(n1361) );
  INVX1 U134 ( .A(n1362), .Y(n1358) );
  INVX1 U135 ( .A(n153), .Y(n1383) );
  INVX1 U136 ( .A(n21), .Y(n1335) );
  INVX1 U137 ( .A(n22), .Y(n1327) );
  INVX1 U138 ( .A(n23), .Y(n1319) );
  INVX1 U139 ( .A(n24), .Y(n1333) );
  INVX1 U140 ( .A(n26), .Y(n1311) );
  INVX1 U141 ( .A(n887), .Y(n1324) );
  INVX1 U142 ( .A(n892), .Y(n1316) );
  INVX1 U143 ( .A(n20), .Y(n1313) );
  INVX1 U144 ( .A(n1367), .Y(n1373) );
  INVX1 U145 ( .A(n1352), .Y(n1363) );
  INVX1 U146 ( .A(n1352), .Y(n1362) );
  INVX1 U147 ( .A(n1374), .Y(n1385) );
  INVX1 U148 ( .A(n1374), .Y(n1384) );
  INVX1 U149 ( .A(n19), .Y(n1351) );
  INVX1 U150 ( .A(n19), .Y(n1350) );
  INVX1 U151 ( .A(n19), .Y(n1349) );
  INVX1 U152 ( .A(n882), .Y(n1332) );
  INVX1 U153 ( .A(n883), .Y(n1330) );
  INVX1 U154 ( .A(n877), .Y(n1340) );
  INVX1 U155 ( .A(n878), .Y(n1338) );
  INVX1 U156 ( .A(n886), .Y(n1326) );
  INVX1 U157 ( .A(n888), .Y(n1322) );
  INVX1 U158 ( .A(n25), .Y(n1317) );
  NOR2X1 U159 ( .A(n1390), .B(n1389), .Y(n869) );
  NAND2X1 U160 ( .A(n1163), .B(n869), .Y(n867) );
  NAND2X1 U161 ( .A(n1159), .B(n1158), .Y(n877) );
  NAND2X1 U162 ( .A(n872), .B(n1158), .Y(n882) );
  NAND2X1 U163 ( .A(n1159), .B(n1157), .Y(n878) );
  NAND2X1 U164 ( .A(n872), .B(n1157), .Y(n883) );
  NAND2X1 U165 ( .A(n872), .B(n1163), .Y(n892) );
  NAND2X1 U166 ( .A(n1159), .B(n1163), .Y(n887) );
  NAND2X1 U167 ( .A(n1162), .B(n1159), .Y(n888) );
  INVX1 U168 ( .A(n152), .Y(n1352) );
  INVX1 U169 ( .A(n153), .Y(n1374) );
  NOR2X1 U170 ( .A(n1390), .B(counter_2[1]), .Y(n872) );
  NOR2X1 U171 ( .A(counter_2[2]), .B(counter_2[1]), .Y(n1159) );
  NOR2X1 U172 ( .A(n861), .B(counter_2[3]), .Y(n1163) );
  OAI221XL U173 ( .A0(n843), .A1(n1339), .B0(n809), .B1(n878), .C0(n1052), .Y(
        n1051) );
  OAI221XL U174 ( .A0(n847), .A1(n1339), .B0(n813), .B1(n1337), .C0(n1084), 
        .Y(n1083) );
  AOI22X1 U175 ( .A0(n1335), .A1(R2[9]), .B0(n1333), .B1(R13[9]), .Y(n1084) );
  OAI221XL U176 ( .A0(n845), .A1(n1339), .B0(n811), .B1(n878), .C0(n1068), .Y(
        n1067) );
  AOI22X1 U177 ( .A0(n1335), .A1(R2[11]), .B0(n1333), .B1(R13[11]), .Y(n1068)
         );
  OAI221XL U178 ( .A0(n844), .A1(n1339), .B0(n810), .B1(n878), .C0(n1060), .Y(
        n1059) );
  AOI22X1 U179 ( .A0(n1335), .A1(R2[12]), .B0(n1334), .B1(R13[12]), .Y(n1060)
         );
  OAI221XL U180 ( .A0(n842), .A1(n1339), .B0(n808), .B1(n878), .C0(n1044), .Y(
        n1043) );
  AOI22X1 U181 ( .A0(n1336), .A1(R2[14]), .B0(n1334), .B1(R13[14]), .Y(n1044)
         );
  OAI221XL U182 ( .A0(n841), .A1(n1339), .B0(n807), .B1(n878), .C0(n1036), .Y(
        n1035) );
  AOI22X1 U183 ( .A0(n1335), .A1(R2[15]), .B0(n1334), .B1(R13[15]), .Y(n1036)
         );
  OAI221XL U184 ( .A0(n840), .A1(n1339), .B0(n806), .B1(n878), .C0(n1028), .Y(
        n1027) );
  OAI221XL U185 ( .A0(n828), .A1(n877), .B0(n794), .B1(n1337), .C0(n932), .Y(
        n931) );
  AOI22X1 U186 ( .A0(n1336), .A1(R2[28]), .B0(n1334), .B1(R13[28]), .Y(n932)
         );
  OAI221XL U187 ( .A0(n825), .A1(n877), .B0(n791), .B1(n1337), .C0(n908), .Y(
        n907) );
  AOI22X1 U188 ( .A0(n1336), .A1(R2[31]), .B0(n1333), .B1(R13[31]), .Y(n908)
         );
  OAI221XL U189 ( .A0(n824), .A1(n877), .B0(n790), .B1(n878), .C0(n900), .Y(
        n899) );
  AOI22X1 U190 ( .A0(n1336), .A1(R2[32]), .B0(n1334), .B1(R13[32]), .Y(n900)
         );
  OAI221XL U191 ( .A0(n823), .A1(n877), .B0(n789), .B1(n1337), .C0(n879), .Y(
        n876) );
  AOI22X1 U192 ( .A0(n1336), .A1(R2[33]), .B0(n1333), .B1(R13[33]), .Y(n879)
         );
  OAI221XL U193 ( .A0(n856), .A1(n877), .B0(n822), .B1(n1337), .C0(n1156), .Y(
        n1155) );
  AOI22X1 U194 ( .A0(n1335), .A1(R2[0]), .B0(n1333), .B1(R13[0]), .Y(n1156) );
  OAI221XL U195 ( .A0(n855), .A1(n1339), .B0(n821), .B1(n1337), .C0(n1148), 
        .Y(n1147) );
  AOI22X1 U196 ( .A0(n1335), .A1(R2[1]), .B0(n1333), .B1(R13[1]), .Y(n1148) );
  OAI221XL U197 ( .A0(n854), .A1(n877), .B0(n820), .B1(n1337), .C0(n1140), .Y(
        n1139) );
  AOI22X1 U198 ( .A0(n1335), .A1(R2[2]), .B0(n1333), .B1(R13[2]), .Y(n1140) );
  OAI221XL U199 ( .A0(n853), .A1(n877), .B0(n819), .B1(n1337), .C0(n1132), .Y(
        n1131) );
  AOI22X1 U200 ( .A0(n1335), .A1(R2[3]), .B0(n1333), .B1(R13[3]), .Y(n1132) );
  OAI221XL U201 ( .A0(n852), .A1(n877), .B0(n818), .B1(n1337), .C0(n1124), .Y(
        n1123) );
  AOI22X1 U202 ( .A0(n1335), .A1(R2[4]), .B0(n1333), .B1(R13[4]), .Y(n1124) );
  OAI221XL U203 ( .A0(n851), .A1(n877), .B0(n817), .B1(n1337), .C0(n1116), .Y(
        n1115) );
  AOI22X1 U204 ( .A0(n1335), .A1(R2[5]), .B0(n1333), .B1(R13[5]), .Y(n1116) );
  OAI221XL U205 ( .A0(n850), .A1(n877), .B0(n816), .B1(n1337), .C0(n1108), .Y(
        n1107) );
  AOI22X1 U206 ( .A0(n1335), .A1(R2[6]), .B0(n1333), .B1(R13[6]), .Y(n1108) );
  OAI221XL U207 ( .A0(n849), .A1(n877), .B0(n815), .B1(n1337), .C0(n1100), .Y(
        n1099) );
  AOI22X1 U208 ( .A0(n1335), .A1(R2[7]), .B0(n1333), .B1(R13[7]), .Y(n1100) );
  OAI221XL U209 ( .A0(n848), .A1(n1339), .B0(n814), .B1(n1337), .C0(n1092), 
        .Y(n1091) );
  AOI22X1 U210 ( .A0(n1335), .A1(R2[8]), .B0(n1333), .B1(R13[8]), .Y(n1092) );
  OAI221XL U211 ( .A0(n846), .A1(n1339), .B0(n812), .B1(n878), .C0(n1076), .Y(
        n1075) );
  AOI22X1 U212 ( .A0(n1335), .A1(R2[10]), .B0(n1333), .B1(R13[10]), .Y(n1076)
         );
  OAI221XL U213 ( .A0(n839), .A1(n1339), .B0(n805), .B1(n1337), .C0(n1020), 
        .Y(n1019) );
  AOI22X1 U214 ( .A0(n1336), .A1(R2[17]), .B0(n1334), .B1(R13[17]), .Y(n1020)
         );
  OAI221XL U215 ( .A0(n838), .A1(n1339), .B0(n804), .B1(n1337), .C0(n1012), 
        .Y(n1011) );
  AOI22X1 U216 ( .A0(n1335), .A1(R2[18]), .B0(n1334), .B1(R13[18]), .Y(n1012)
         );
  OAI221XL U217 ( .A0(n837), .A1(n1339), .B0(n803), .B1(n1337), .C0(n1004), 
        .Y(n1003) );
  AOI22X1 U218 ( .A0(n1336), .A1(R2[19]), .B0(n1334), .B1(R13[19]), .Y(n1004)
         );
  OAI221XL U219 ( .A0(n836), .A1(n1339), .B0(n802), .B1(n1337), .C0(n996), .Y(
        n995) );
  AOI22X1 U220 ( .A0(n1335), .A1(R2[20]), .B0(n1334), .B1(R13[20]), .Y(n996)
         );
  OAI221XL U221 ( .A0(n835), .A1(n877), .B0(n801), .B1(n878), .C0(n988), .Y(
        n987) );
  AOI22X1 U222 ( .A0(n1336), .A1(R2[21]), .B0(n1334), .B1(R13[21]), .Y(n988)
         );
  OAI221XL U223 ( .A0(n834), .A1(n877), .B0(n800), .B1(n878), .C0(n980), .Y(
        n979) );
  AOI22X1 U224 ( .A0(n1336), .A1(R2[22]), .B0(n1334), .B1(R13[22]), .Y(n980)
         );
  OAI221XL U225 ( .A0(n833), .A1(n877), .B0(n799), .B1(n878), .C0(n972), .Y(
        n971) );
  AOI22X1 U226 ( .A0(n1336), .A1(R2[23]), .B0(n1334), .B1(R13[23]), .Y(n972)
         );
  OAI221XL U227 ( .A0(n832), .A1(n877), .B0(n798), .B1(n878), .C0(n964), .Y(
        n963) );
  AOI22X1 U228 ( .A0(n1336), .A1(R2[24]), .B0(n1334), .B1(R13[24]), .Y(n964)
         );
  OAI221XL U229 ( .A0(n831), .A1(n877), .B0(n797), .B1(n878), .C0(n956), .Y(
        n955) );
  AOI22X1 U230 ( .A0(n1336), .A1(R2[25]), .B0(n1333), .B1(R13[25]), .Y(n956)
         );
  OAI221XL U231 ( .A0(n830), .A1(n877), .B0(n796), .B1(n878), .C0(n948), .Y(
        n947) );
  AOI22X1 U232 ( .A0(n1336), .A1(R2[26]), .B0(n1334), .B1(R13[26]), .Y(n948)
         );
  OAI221XL U233 ( .A0(n829), .A1(n1339), .B0(n795), .B1(n878), .C0(n940), .Y(
        n939) );
  AOI22X1 U234 ( .A0(n1336), .A1(R2[27]), .B0(n1333), .B1(R13[27]), .Y(n940)
         );
  OAI221XL U235 ( .A0(n827), .A1(n1339), .B0(n793), .B1(n878), .C0(n924), .Y(
        n923) );
  AOI22X1 U236 ( .A0(n1336), .A1(R2[29]), .B0(n1334), .B1(R13[29]), .Y(n924)
         );
  OAI221XL U237 ( .A0(n826), .A1(n1339), .B0(n792), .B1(n878), .C0(n916), .Y(
        n915) );
  AOI22X1 U238 ( .A0(n1336), .A1(R2[30]), .B0(n1333), .B1(R13[30]), .Y(n916)
         );
  NOR2X1 U239 ( .A(counter_2[3]), .B(counter_2[0]), .Y(n1162) );
  NOR2X1 U240 ( .A(n1389), .B(counter_2[2]), .Y(n871) );
  INVX1 U241 ( .A(counter_2[1]), .Y(n1389) );
  OR3XL U242 ( .A(n584), .B(p_s_flag_in), .C(n1387), .Y(n151) );
  OR3XL U243 ( .A(counter_1[0]), .B(p_s_flag_in), .C(n1387), .Y(n152) );
  OR3XL U244 ( .A(counter_1[1]), .B(p_s_flag_in), .C(counter_1[0]), .Y(n153)
         );
  INVX1 U245 ( .A(counter_1[1]), .Y(n1387) );
  AOI22X1 U246 ( .A0(n1327), .A1(R3[11]), .B0(n1325), .B1(R14[11]), .Y(n1069)
         );
  AOI22X1 U247 ( .A0(n1319), .A1(R0[11]), .B0(n1317), .B1(R15[11]), .Y(n1070)
         );
  AOI22X1 U248 ( .A0(n1309), .A1(R1[11]), .B0(n1311), .B1(R12[11]), .Y(n1071)
         );
  AOI22X1 U249 ( .A0(n1328), .A1(R3[14]), .B0(n886), .B1(R14[14]), .Y(n1045)
         );
  AOI22X1 U250 ( .A0(n1320), .A1(R0[14]), .B0(n1318), .B1(R15[14]), .Y(n1046)
         );
  AOI22X1 U251 ( .A0(n1309), .A1(R1[14]), .B0(n1312), .B1(R12[14]), .Y(n1047)
         );
  AOI22X1 U252 ( .A0(n1328), .A1(R3[15]), .B0(n886), .B1(R14[15]), .Y(n1037)
         );
  AOI22X1 U253 ( .A0(n1320), .A1(R0[15]), .B0(n1318), .B1(R15[15]), .Y(n1038)
         );
  AOI22X1 U254 ( .A0(n1309), .A1(R1[15]), .B0(n1312), .B1(R12[15]), .Y(n1039)
         );
  AOI22X1 U255 ( .A0(n1328), .A1(R3[30]), .B0(n1325), .B1(R14[30]), .Y(n917)
         );
  AOI22X1 U256 ( .A0(n1320), .A1(R0[30]), .B0(n1317), .B1(R15[30]), .Y(n918)
         );
  AOI22X1 U257 ( .A0(n1310), .A1(R1[30]), .B0(n1311), .B1(R12[30]), .Y(n919)
         );
  AOI22X1 U258 ( .A0(n1327), .A1(R3[31]), .B0(n1325), .B1(R14[31]), .Y(n909)
         );
  AOI22X1 U259 ( .A0(n1320), .A1(R0[31]), .B0(n1318), .B1(R15[31]), .Y(n910)
         );
  AOI22X1 U260 ( .A0(n1310), .A1(R1[31]), .B0(n1312), .B1(R12[31]), .Y(n911)
         );
  AOI22X1 U261 ( .A0(n1328), .A1(R3[32]), .B0(n1325), .B1(R14[32]), .Y(n901)
         );
  AOI22X1 U262 ( .A0(n1320), .A1(R0[32]), .B0(n1318), .B1(R15[32]), .Y(n902)
         );
  AOI22X1 U263 ( .A0(n1310), .A1(R1[32]), .B0(n1312), .B1(R12[32]), .Y(n903)
         );
  AOI22X1 U264 ( .A0(n1327), .A1(R3[33]), .B0(n1325), .B1(R14[33]), .Y(n884)
         );
  AOI22X1 U265 ( .A0(n1320), .A1(R0[33]), .B0(n1317), .B1(R15[33]), .Y(n889)
         );
  AOI22X1 U266 ( .A0(n1309), .A1(R1[33]), .B0(n1311), .B1(R12[33]), .Y(n894)
         );
  AOI22X1 U267 ( .A0(n1328), .A1(R3[28]), .B0(n1325), .B1(R14[28]), .Y(n933)
         );
  AOI22X1 U268 ( .A0(n1320), .A1(R0[28]), .B0(n1317), .B1(R15[28]), .Y(n934)
         );
  AOI22X1 U269 ( .A0(n1310), .A1(R1[28]), .B0(n1312), .B1(R12[28]), .Y(n935)
         );
  INVX1 U270 ( .A(counter_2[2]), .Y(n1390) );
  AOI22X1 U271 ( .A0(n1327), .A1(R3[0]), .B0(n886), .B1(R14[0]), .Y(n1160) );
  AOI22X1 U272 ( .A0(n1319), .A1(R0[0]), .B0(n1317), .B1(R15[0]), .Y(n1161) );
  AOI22X1 U273 ( .A0(n1310), .A1(R1[0]), .B0(n1311), .B1(R12[0]), .Y(n1164) );
  AOI22X1 U274 ( .A0(n1327), .A1(R3[1]), .B0(n886), .B1(R14[1]), .Y(n1149) );
  AOI22X1 U275 ( .A0(n1319), .A1(R0[1]), .B0(n1317), .B1(R15[1]), .Y(n1150) );
  AOI22X1 U276 ( .A0(n1310), .A1(R1[1]), .B0(n1311), .B1(R12[1]), .Y(n1151) );
  AOI22X1 U277 ( .A0(n1327), .A1(R3[2]), .B0(n886), .B1(R14[2]), .Y(n1141) );
  AOI22X1 U278 ( .A0(n1319), .A1(R0[2]), .B0(n1317), .B1(R15[2]), .Y(n1142) );
  AOI22X1 U279 ( .A0(n1310), .A1(R1[2]), .B0(n1311), .B1(R12[2]), .Y(n1143) );
  AOI22X1 U280 ( .A0(n1327), .A1(R3[3]), .B0(n886), .B1(R14[3]), .Y(n1133) );
  AOI22X1 U281 ( .A0(n1319), .A1(R0[3]), .B0(n1317), .B1(R15[3]), .Y(n1134) );
  AOI22X1 U282 ( .A0(n1310), .A1(R1[3]), .B0(n1311), .B1(R12[3]), .Y(n1135) );
  AOI22X1 U283 ( .A0(n1327), .A1(R3[4]), .B0(n886), .B1(R14[4]), .Y(n1125) );
  AOI22X1 U284 ( .A0(n1319), .A1(R0[4]), .B0(n1317), .B1(R15[4]), .Y(n1126) );
  AOI22X1 U285 ( .A0(n1310), .A1(R1[4]), .B0(n1311), .B1(R12[4]), .Y(n1127) );
  AOI22X1 U286 ( .A0(n1327), .A1(R3[5]), .B0(n886), .B1(R14[5]), .Y(n1117) );
  AOI22X1 U287 ( .A0(n1319), .A1(R0[5]), .B0(n1317), .B1(R15[5]), .Y(n1118) );
  AOI22X1 U288 ( .A0(n1310), .A1(R1[5]), .B0(n1311), .B1(R12[5]), .Y(n1119) );
  AOI22X1 U289 ( .A0(n1327), .A1(R3[6]), .B0(n886), .B1(R14[6]), .Y(n1109) );
  AOI22X1 U290 ( .A0(n1319), .A1(R0[6]), .B0(n1317), .B1(R15[6]), .Y(n1110) );
  AOI22X1 U291 ( .A0(n1310), .A1(R1[6]), .B0(n1311), .B1(R12[6]), .Y(n1111) );
  AOI22X1 U292 ( .A0(n1327), .A1(R3[7]), .B0(n886), .B1(R14[7]), .Y(n1101) );
  AOI22X1 U293 ( .A0(n1319), .A1(R0[7]), .B0(n1317), .B1(R15[7]), .Y(n1102) );
  AOI22X1 U294 ( .A0(n1310), .A1(R1[7]), .B0(n1311), .B1(R12[7]), .Y(n1103) );
  AOI22X1 U295 ( .A0(n1327), .A1(R3[8]), .B0(n1325), .B1(R14[8]), .Y(n1093) );
  AOI22X1 U296 ( .A0(n1319), .A1(R0[8]), .B0(n1317), .B1(R15[8]), .Y(n1094) );
  AOI22X1 U297 ( .A0(n1310), .A1(R1[8]), .B0(n1311), .B1(R12[8]), .Y(n1095) );
  AOI22X1 U298 ( .A0(n1327), .A1(R3[9]), .B0(n886), .B1(R14[9]), .Y(n1085) );
  AOI22X1 U299 ( .A0(n1319), .A1(R0[9]), .B0(n1317), .B1(R15[9]), .Y(n1086) );
  AOI22X1 U300 ( .A0(n1310), .A1(R1[9]), .B0(n1311), .B1(R12[9]), .Y(n1087) );
  AOI22X1 U301 ( .A0(n1327), .A1(R3[10]), .B0(n886), .B1(R14[10]), .Y(n1077)
         );
  AOI22X1 U302 ( .A0(n1319), .A1(R0[10]), .B0(n1317), .B1(R15[10]), .Y(n1078)
         );
  AOI22X1 U303 ( .A0(n1309), .A1(R1[10]), .B0(n1311), .B1(R12[10]), .Y(n1079)
         );
  AOI22X1 U304 ( .A0(n1328), .A1(R3[12]), .B0(n886), .B1(R14[12]), .Y(n1061)
         );
  AOI22X1 U305 ( .A0(n1319), .A1(R0[12]), .B0(n1318), .B1(R15[12]), .Y(n1062)
         );
  AOI22X1 U306 ( .A0(n1309), .A1(R1[12]), .B0(n1312), .B1(R12[12]), .Y(n1063)
         );
  AOI22X1 U307 ( .A0(n1328), .A1(R3[17]), .B0(n886), .B1(R14[17]), .Y(n1021)
         );
  AOI22X1 U308 ( .A0(n1320), .A1(R0[17]), .B0(n1318), .B1(R15[17]), .Y(n1022)
         );
  AOI22X1 U309 ( .A0(n1309), .A1(R1[17]), .B0(n1312), .B1(R12[17]), .Y(n1023)
         );
  AOI22X1 U310 ( .A0(n1328), .A1(R3[18]), .B0(n886), .B1(R14[18]), .Y(n1013)
         );
  AOI22X1 U311 ( .A0(n1319), .A1(R0[18]), .B0(n1318), .B1(R15[18]), .Y(n1014)
         );
  AOI22X1 U312 ( .A0(n1309), .A1(R1[18]), .B0(n1312), .B1(R12[18]), .Y(n1015)
         );
  AOI22X1 U313 ( .A0(n1328), .A1(R3[19]), .B0(n886), .B1(R14[19]), .Y(n1005)
         );
  AOI22X1 U314 ( .A0(n1320), .A1(R0[19]), .B0(n1318), .B1(R15[19]), .Y(n1006)
         );
  AOI22X1 U315 ( .A0(n1309), .A1(R1[19]), .B0(n1312), .B1(R12[19]), .Y(n1007)
         );
  AOI22X1 U316 ( .A0(n1328), .A1(R3[20]), .B0(n886), .B1(R14[20]), .Y(n997) );
  AOI22X1 U317 ( .A0(n1319), .A1(R0[20]), .B0(n1318), .B1(R15[20]), .Y(n998)
         );
  AOI22X1 U318 ( .A0(n1309), .A1(R1[20]), .B0(n1312), .B1(R12[20]), .Y(n999)
         );
  AOI22X1 U319 ( .A0(n1328), .A1(R3[21]), .B0(n886), .B1(R14[21]), .Y(n989) );
  AOI22X1 U320 ( .A0(n1320), .A1(R0[21]), .B0(n1318), .B1(R15[21]), .Y(n990)
         );
  AOI22X1 U322 ( .A0(n1309), .A1(R1[21]), .B0(n1312), .B1(R12[21]), .Y(n991)
         );
  AOI22X1 U323 ( .A0(n1328), .A1(R3[22]), .B0(n886), .B1(R14[22]), .Y(n981) );
  AOI22X1 U325 ( .A0(n1319), .A1(R0[22]), .B0(n1318), .B1(R15[22]), .Y(n982)
         );
  AOI22X1 U327 ( .A0(n1309), .A1(R1[22]), .B0(n1312), .B1(R12[22]), .Y(n983)
         );
  AOI22X1 U328 ( .A0(n1328), .A1(R3[23]), .B0(n886), .B1(R14[23]), .Y(n973) );
  AOI22X1 U329 ( .A0(n1320), .A1(R0[23]), .B0(n1318), .B1(R15[23]), .Y(n974)
         );
  AOI22X1 U330 ( .A0(n1310), .A1(R1[23]), .B0(n1312), .B1(R12[23]), .Y(n975)
         );
  AOI22X1 U331 ( .A0(n1327), .A1(R3[24]), .B0(n1325), .B1(R14[24]), .Y(n965)
         );
  AOI22X1 U332 ( .A0(n1320), .A1(R0[24]), .B0(n1318), .B1(R15[24]), .Y(n966)
         );
  AOI22X1 U333 ( .A0(n1309), .A1(R1[24]), .B0(n1311), .B1(R12[24]), .Y(n967)
         );
  AOI22X1 U334 ( .A0(n1328), .A1(R3[25]), .B0(n1325), .B1(R14[25]), .Y(n957)
         );
  AOI22X1 U335 ( .A0(n1320), .A1(R0[25]), .B0(n1317), .B1(R15[25]), .Y(n958)
         );
  AOI22X1 U336 ( .A0(n1310), .A1(R1[25]), .B0(n1312), .B1(R12[25]), .Y(n959)
         );
  AOI22X1 U337 ( .A0(n1327), .A1(R3[26]), .B0(n1325), .B1(R14[26]), .Y(n949)
         );
  AOI22X1 U338 ( .A0(n1320), .A1(R0[26]), .B0(n1318), .B1(R15[26]), .Y(n950)
         );
  AOI22X1 U339 ( .A0(n1309), .A1(R1[26]), .B0(n1311), .B1(R12[26]), .Y(n951)
         );
  AOI22X1 U340 ( .A0(n1328), .A1(R3[27]), .B0(n1325), .B1(R14[27]), .Y(n941)
         );
  AOI22X1 U341 ( .A0(n1320), .A1(R0[27]), .B0(n1317), .B1(R15[27]), .Y(n942)
         );
  AOI22X1 U342 ( .A0(n1310), .A1(R1[27]), .B0(n1312), .B1(R12[27]), .Y(n943)
         );
  AOI22X1 U343 ( .A0(n1327), .A1(R3[29]), .B0(n1325), .B1(R14[29]), .Y(n925)
         );
  AOI22X1 U344 ( .A0(n1320), .A1(R0[29]), .B0(n1318), .B1(R15[29]), .Y(n926)
         );
  AOI22X1 U345 ( .A0(n1309), .A1(R1[29]), .B0(n1311), .B1(R12[29]), .Y(n927)
         );
  OR4X2 U346 ( .A(n1048), .B(n1049), .C(n1050), .D(n1051), .Y(N132) );
  OAI221XL U347 ( .A0(n775), .A1(n1315), .B0(n741), .B1(n1314), .C0(n1055), 
        .Y(n1048) );
  OAI221XL U348 ( .A0(n707), .A1(n1323), .B0(n605), .B1(n888), .C0(n1054), .Y(
        n1049) );
  OAI221XL U349 ( .A0(n639), .A1(n1331), .B0(n673), .B1(n883), .C0(n1053), .Y(
        n1050) );
  OR4X2 U350 ( .A(n1024), .B(n1025), .C(n1026), .D(n1027), .Y(N135) );
  OAI221XL U351 ( .A0(n772), .A1(n1315), .B0(n738), .B1(n1314), .C0(n1031), 
        .Y(n1024) );
  OAI221XL U352 ( .A0(n704), .A1(n1323), .B0(n602), .B1(n888), .C0(n1030), .Y(
        n1025) );
  OAI221XL U353 ( .A0(n636), .A1(n1331), .B0(n670), .B1(n883), .C0(n1029), .Y(
        n1026) );
  OR4X2 U354 ( .A(n1064), .B(n1065), .C(n1066), .D(n1067), .Y(N130) );
  OAI221XL U355 ( .A0(n777), .A1(n1315), .B0(n743), .B1(n1314), .C0(n1071), 
        .Y(n1064) );
  OAI221XL U356 ( .A0(n709), .A1(n1323), .B0(n607), .B1(n888), .C0(n1070), .Y(
        n1065) );
  OAI221XL U357 ( .A0(n641), .A1(n1331), .B0(n675), .B1(n883), .C0(n1069), .Y(
        n1066) );
  OR4X2 U358 ( .A(n1040), .B(n1041), .C(n1042), .D(n1043), .Y(N133) );
  OAI221XL U359 ( .A0(n774), .A1(n1315), .B0(n740), .B1(n1314), .C0(n1047), 
        .Y(n1040) );
  OAI221XL U360 ( .A0(n706), .A1(n1323), .B0(n604), .B1(n888), .C0(n1046), .Y(
        n1041) );
  OAI221XL U361 ( .A0(n638), .A1(n1331), .B0(n672), .B1(n883), .C0(n1045), .Y(
        n1042) );
  OR4X2 U362 ( .A(n1032), .B(n1033), .C(n1034), .D(n1035), .Y(N134) );
  OAI221XL U363 ( .A0(n773), .A1(n1315), .B0(n739), .B1(n1314), .C0(n1039), 
        .Y(n1032) );
  OAI221XL U364 ( .A0(n705), .A1(n1323), .B0(n603), .B1(n888), .C0(n1038), .Y(
        n1033) );
  OAI221XL U365 ( .A0(n637), .A1(n1331), .B0(n671), .B1(n883), .C0(n1037), .Y(
        n1034) );
  OR4X2 U366 ( .A(n912), .B(n913), .C(n914), .D(n915), .Y(N149) );
  OAI221XL U367 ( .A0(n758), .A1(n892), .B0(n724), .B1(n1313), .C0(n919), .Y(
        n912) );
  OAI221XL U368 ( .A0(n690), .A1(n887), .B0(n588), .B1(n1321), .C0(n918), .Y(
        n913) );
  OAI221XL U369 ( .A0(n622), .A1(n882), .B0(n656), .B1(n1329), .C0(n917), .Y(
        n914) );
  OR4X2 U370 ( .A(n904), .B(n905), .C(n906), .D(n907), .Y(N150) );
  OAI221XL U371 ( .A0(n757), .A1(n1315), .B0(n723), .B1(n1313), .C0(n911), .Y(
        n904) );
  OAI221XL U372 ( .A0(n689), .A1(n1323), .B0(n587), .B1(n1321), .C0(n910), .Y(
        n905) );
  OAI221XL U373 ( .A0(n621), .A1(n882), .B0(n655), .B1(n1329), .C0(n909), .Y(
        n906) );
  OR4X2 U374 ( .A(n896), .B(n897), .C(n898), .D(n899), .Y(N151) );
  OAI221XL U375 ( .A0(n756), .A1(n892), .B0(n722), .B1(n1313), .C0(n903), .Y(
        n896) );
  OAI221XL U376 ( .A0(n688), .A1(n887), .B0(n586), .B1(n888), .C0(n902), .Y(
        n897) );
  OAI221XL U377 ( .A0(n620), .A1(n882), .B0(n654), .B1(n1329), .C0(n901), .Y(
        n898) );
  OR4X2 U378 ( .A(n873), .B(n874), .C(n875), .D(n876), .Y(N152) );
  OAI221XL U379 ( .A0(n755), .A1(n1315), .B0(n721), .B1(n1313), .C0(n894), .Y(
        n873) );
  OAI221XL U380 ( .A0(n687), .A1(n1323), .B0(n585), .B1(n1321), .C0(n889), .Y(
        n874) );
  OAI221XL U381 ( .A0(n619), .A1(n882), .B0(n653), .B1(n1329), .C0(n884), .Y(
        n875) );
  OR4X2 U382 ( .A(n928), .B(n929), .C(n930), .D(n931), .Y(N147) );
  OAI221XL U383 ( .A0(n760), .A1(n892), .B0(n726), .B1(n1313), .C0(n935), .Y(
        n928) );
  OAI221XL U384 ( .A0(n692), .A1(n887), .B0(n590), .B1(n888), .C0(n934), .Y(
        n929) );
  OAI221XL U385 ( .A0(n624), .A1(n882), .B0(n658), .B1(n883), .C0(n933), .Y(
        n930) );
  OR4X2 U386 ( .A(n1152), .B(n1153), .C(n1154), .D(n1155), .Y(N119) );
  OAI221XL U387 ( .A0(n788), .A1(n892), .B0(n754), .B1(n1314), .C0(n1164), .Y(
        n1152) );
  OAI221XL U388 ( .A0(n720), .A1(n887), .B0(n618), .B1(n1321), .C0(n1161), .Y(
        n1153) );
  OAI221XL U389 ( .A0(n652), .A1(n882), .B0(n686), .B1(n1329), .C0(n1160), .Y(
        n1154) );
  OR4X2 U390 ( .A(n1144), .B(n1145), .C(n1146), .D(n1147), .Y(N120) );
  OAI221XL U391 ( .A0(n787), .A1(n1315), .B0(n753), .B1(n1313), .C0(n1151), 
        .Y(n1144) );
  OAI221XL U392 ( .A0(n719), .A1(n1323), .B0(n617), .B1(n1321), .C0(n1150), 
        .Y(n1145) );
  OAI221XL U393 ( .A0(n651), .A1(n1331), .B0(n685), .B1(n1329), .C0(n1149), 
        .Y(n1146) );
  OR4X2 U394 ( .A(n1136), .B(n1137), .C(n1138), .D(n1139), .Y(N121) );
  OAI221XL U395 ( .A0(n786), .A1(n892), .B0(n752), .B1(n1314), .C0(n1143), .Y(
        n1136) );
  OAI221XL U396 ( .A0(n718), .A1(n887), .B0(n616), .B1(n1321), .C0(n1142), .Y(
        n1137) );
  OAI221XL U397 ( .A0(n650), .A1(n882), .B0(n684), .B1(n1329), .C0(n1141), .Y(
        n1138) );
  OR4X2 U398 ( .A(n1128), .B(n1129), .C(n1130), .D(n1131), .Y(N122) );
  OAI221XL U399 ( .A0(n785), .A1(n892), .B0(n751), .B1(n1313), .C0(n1135), .Y(
        n1128) );
  OAI221XL U400 ( .A0(n717), .A1(n887), .B0(n615), .B1(n1321), .C0(n1134), .Y(
        n1129) );
  OAI221XL U401 ( .A0(n649), .A1(n882), .B0(n683), .B1(n1329), .C0(n1133), .Y(
        n1130) );
  OR4X2 U402 ( .A(n1120), .B(n1121), .C(n1122), .D(n1123), .Y(N123) );
  OAI221XL U403 ( .A0(n784), .A1(n892), .B0(n750), .B1(n1314), .C0(n1127), .Y(
        n1120) );
  OAI221XL U404 ( .A0(n716), .A1(n887), .B0(n614), .B1(n1321), .C0(n1126), .Y(
        n1121) );
  OAI221XL U405 ( .A0(n648), .A1(n882), .B0(n682), .B1(n1329), .C0(n1125), .Y(
        n1122) );
  OR4X2 U406 ( .A(n1112), .B(n1113), .C(n1114), .D(n1115), .Y(N124) );
  OAI221XL U407 ( .A0(n783), .A1(n892), .B0(n749), .B1(n1313), .C0(n1119), .Y(
        n1112) );
  OAI221XL U408 ( .A0(n715), .A1(n887), .B0(n613), .B1(n1321), .C0(n1118), .Y(
        n1113) );
  OAI221XL U409 ( .A0(n647), .A1(n882), .B0(n681), .B1(n1329), .C0(n1117), .Y(
        n1114) );
  OR4X2 U410 ( .A(n1104), .B(n1105), .C(n1106), .D(n1107), .Y(N125) );
  OAI221XL U411 ( .A0(n782), .A1(n892), .B0(n748), .B1(n1314), .C0(n1111), .Y(
        n1104) );
  OAI221XL U412 ( .A0(n714), .A1(n887), .B0(n612), .B1(n1321), .C0(n1110), .Y(
        n1105) );
  OAI221XL U413 ( .A0(n646), .A1(n882), .B0(n680), .B1(n1329), .C0(n1109), .Y(
        n1106) );
  OR4X2 U414 ( .A(n1096), .B(n1097), .C(n1098), .D(n1099), .Y(N126) );
  OAI221XL U415 ( .A0(n781), .A1(n892), .B0(n747), .B1(n1313), .C0(n1103), .Y(
        n1096) );
  OAI221XL U416 ( .A0(n713), .A1(n887), .B0(n611), .B1(n1321), .C0(n1102), .Y(
        n1097) );
  OAI221XL U417 ( .A0(n645), .A1(n882), .B0(n679), .B1(n1329), .C0(n1101), .Y(
        n1098) );
  OR4X2 U418 ( .A(n1088), .B(n1089), .C(n1090), .D(n1091), .Y(N127) );
  OAI221XL U419 ( .A0(n780), .A1(n1315), .B0(n746), .B1(n1314), .C0(n1095), 
        .Y(n1088) );
  OAI221XL U420 ( .A0(n712), .A1(n1323), .B0(n610), .B1(n1321), .C0(n1094), 
        .Y(n1089) );
  OAI221XL U421 ( .A0(n644), .A1(n1331), .B0(n678), .B1(n1329), .C0(n1093), 
        .Y(n1090) );
  OR4X2 U422 ( .A(n1080), .B(n1081), .C(n1082), .D(n1083), .Y(N128) );
  OAI221XL U423 ( .A0(n779), .A1(n1315), .B0(n745), .B1(n1313), .C0(n1087), 
        .Y(n1080) );
  OAI221XL U424 ( .A0(n711), .A1(n1323), .B0(n609), .B1(n1321), .C0(n1086), 
        .Y(n1081) );
  OAI221XL U425 ( .A0(n643), .A1(n1331), .B0(n677), .B1(n1329), .C0(n1085), 
        .Y(n1082) );
  OR4X2 U426 ( .A(n1072), .B(n1073), .C(n1074), .D(n1075), .Y(N129) );
  OAI221XL U427 ( .A0(n778), .A1(n1315), .B0(n744), .B1(n1314), .C0(n1079), 
        .Y(n1072) );
  OAI221XL U428 ( .A0(n710), .A1(n1323), .B0(n608), .B1(n888), .C0(n1078), .Y(
        n1073) );
  OAI221XL U429 ( .A0(n642), .A1(n1331), .B0(n676), .B1(n883), .C0(n1077), .Y(
        n1074) );
  OR4X2 U430 ( .A(n1056), .B(n1057), .C(n1058), .D(n1059), .Y(N131) );
  OAI221XL U431 ( .A0(n776), .A1(n1315), .B0(n742), .B1(n1314), .C0(n1063), 
        .Y(n1056) );
  OAI221XL U432 ( .A0(n708), .A1(n1323), .B0(n606), .B1(n888), .C0(n1062), .Y(
        n1057) );
  OAI221XL U433 ( .A0(n640), .A1(n1331), .B0(n674), .B1(n883), .C0(n1061), .Y(
        n1058) );
  OR4X2 U434 ( .A(n1016), .B(n1017), .C(n1018), .D(n1019), .Y(N136) );
  OAI221XL U435 ( .A0(n771), .A1(n1315), .B0(n737), .B1(n1314), .C0(n1023), 
        .Y(n1016) );
  OAI221XL U436 ( .A0(n703), .A1(n1323), .B0(n601), .B1(n888), .C0(n1022), .Y(
        n1017) );
  OAI221XL U437 ( .A0(n635), .A1(n1331), .B0(n669), .B1(n883), .C0(n1021), .Y(
        n1018) );
  OR4X2 U438 ( .A(n1008), .B(n1009), .C(n1010), .D(n1011), .Y(N137) );
  OAI221XL U439 ( .A0(n770), .A1(n1315), .B0(n736), .B1(n1314), .C0(n1015), 
        .Y(n1008) );
  OAI221XL U440 ( .A0(n702), .A1(n1323), .B0(n600), .B1(n1321), .C0(n1014), 
        .Y(n1009) );
  OAI221XL U441 ( .A0(n634), .A1(n1331), .B0(n668), .B1(n883), .C0(n1013), .Y(
        n1010) );
  OR4X2 U442 ( .A(n1000), .B(n1001), .C(n1002), .D(n1003), .Y(N138) );
  OAI221XL U443 ( .A0(n769), .A1(n1315), .B0(n735), .B1(n1314), .C0(n1007), 
        .Y(n1000) );
  OAI221XL U444 ( .A0(n701), .A1(n1323), .B0(n599), .B1(n1321), .C0(n1006), 
        .Y(n1001) );
  OAI221XL U445 ( .A0(n633), .A1(n1331), .B0(n667), .B1(n1329), .C0(n1005), 
        .Y(n1002) );
  OR4X2 U446 ( .A(n992), .B(n993), .C(n994), .D(n995), .Y(N139) );
  OAI221XL U447 ( .A0(n768), .A1(n1315), .B0(n734), .B1(n1314), .C0(n999), .Y(
        n992) );
  OAI221XL U448 ( .A0(n700), .A1(n1323), .B0(n598), .B1(n1321), .C0(n998), .Y(
        n993) );
  OAI221XL U449 ( .A0(n632), .A1(n1331), .B0(n666), .B1(n1329), .C0(n997), .Y(
        n994) );
  OR4X2 U450 ( .A(n984), .B(n985), .C(n986), .D(n987), .Y(N140) );
  OAI221XL U451 ( .A0(n767), .A1(n1315), .B0(n733), .B1(n1314), .C0(n991), .Y(
        n984) );
  OAI221XL U452 ( .A0(n699), .A1(n1323), .B0(n597), .B1(n1321), .C0(n990), .Y(
        n985) );
  OAI221XL U453 ( .A0(n631), .A1(n882), .B0(n665), .B1(n883), .C0(n989), .Y(
        n986) );
  OR4X2 U454 ( .A(n976), .B(n977), .C(n978), .D(n979), .Y(N141) );
  OAI221XL U455 ( .A0(n766), .A1(n892), .B0(n732), .B1(n1313), .C0(n983), .Y(
        n976) );
  OAI221XL U456 ( .A0(n698), .A1(n887), .B0(n596), .B1(n888), .C0(n982), .Y(
        n977) );
  OAI221XL U457 ( .A0(n630), .A1(n882), .B0(n664), .B1(n1329), .C0(n981), .Y(
        n978) );
  OR4X2 U458 ( .A(n968), .B(n969), .C(n970), .D(n971), .Y(N142) );
  OAI221XL U459 ( .A0(n765), .A1(n892), .B0(n731), .B1(n1313), .C0(n975), .Y(
        n968) );
  OAI221XL U460 ( .A0(n697), .A1(n887), .B0(n595), .B1(n888), .C0(n974), .Y(
        n969) );
  OAI221XL U461 ( .A0(n629), .A1(n882), .B0(n663), .B1(n883), .C0(n973), .Y(
        n970) );
  OR4X2 U462 ( .A(n960), .B(n961), .C(n962), .D(n963), .Y(N143) );
  OAI221XL U463 ( .A0(n764), .A1(n892), .B0(n730), .B1(n1313), .C0(n967), .Y(
        n960) );
  OAI221XL U464 ( .A0(n696), .A1(n887), .B0(n594), .B1(n888), .C0(n966), .Y(
        n961) );
  OAI221XL U465 ( .A0(n628), .A1(n882), .B0(n662), .B1(n883), .C0(n965), .Y(
        n962) );
  OR4X2 U466 ( .A(n952), .B(n953), .C(n954), .D(n955), .Y(N144) );
  OAI221XL U467 ( .A0(n763), .A1(n892), .B0(n729), .B1(n1313), .C0(n959), .Y(
        n952) );
  OAI221XL U468 ( .A0(n695), .A1(n887), .B0(n593), .B1(n888), .C0(n958), .Y(
        n953) );
  OAI221XL U469 ( .A0(n627), .A1(n882), .B0(n661), .B1(n883), .C0(n957), .Y(
        n954) );
  OR4X2 U470 ( .A(n944), .B(n945), .C(n946), .D(n947), .Y(N145) );
  OAI221XL U471 ( .A0(n762), .A1(n892), .B0(n728), .B1(n1313), .C0(n951), .Y(
        n944) );
  OAI221XL U472 ( .A0(n694), .A1(n887), .B0(n592), .B1(n888), .C0(n950), .Y(
        n945) );
  OAI221XL U473 ( .A0(n626), .A1(n1331), .B0(n660), .B1(n883), .C0(n949), .Y(
        n946) );
  OR4X2 U474 ( .A(n936), .B(n937), .C(n938), .D(n939), .Y(N146) );
  OAI221XL U475 ( .A0(n761), .A1(n892), .B0(n727), .B1(n1313), .C0(n943), .Y(
        n936) );
  OAI221XL U476 ( .A0(n693), .A1(n887), .B0(n591), .B1(n888), .C0(n942), .Y(
        n937) );
  OAI221XL U477 ( .A0(n625), .A1(n1331), .B0(n659), .B1(n883), .C0(n941), .Y(
        n938) );
  OR4X2 U478 ( .A(n920), .B(n921), .C(n922), .D(n923), .Y(N148) );
  OAI221XL U479 ( .A0(n759), .A1(n892), .B0(n725), .B1(n1313), .C0(n927), .Y(
        n920) );
  OAI221XL U480 ( .A0(n691), .A1(n887), .B0(n589), .B1(n888), .C0(n926), .Y(
        n921) );
  OAI221XL U481 ( .A0(n623), .A1(n1331), .B0(n657), .B1(n883), .C0(n925), .Y(
        n922) );
  INVX1 U482 ( .A(n870), .Y(n1388) );
  AOI221X1 U483 ( .A0(counter_2[0]), .A1(n871), .B0(n861), .B1(counter_2[2]), 
        .C0(n872), .Y(n870) );
  NAND2X1 U484 ( .A(n867), .B(n868), .Y(N52) );
  OAI2BB1X1 U485 ( .A0N(n869), .A1N(counter_2[0]), .B0(counter_2[3]), .Y(n868)
         );
  INVX1 U486 ( .A(p_s_flag_in), .Y(n1391) );
  XNOR2X1 U487 ( .A(n1389), .B(counter_2[0]), .Y(N50) );
  XNOR2X1 U488 ( .A(n1387), .B(counter_1[0]), .Y(N26) );
  AOI22X1 U489 ( .A0(n1336), .A1(R2[13]), .B0(n1334), .B1(R13[13]), .Y(n1052)
         );
  AOI22X1 U490 ( .A0(n1328), .A1(R3[13]), .B0(n886), .B1(R14[13]), .Y(n1053)
         );
  AOI22X1 U491 ( .A0(n1319), .A1(R0[13]), .B0(n1318), .B1(R15[13]), .Y(n1054)
         );
  AOI22X1 U492 ( .A0(n1309), .A1(R1[13]), .B0(n1312), .B1(R12[13]), .Y(n1055)
         );
  AOI22X1 U493 ( .A0(n1335), .A1(R2[16]), .B0(n1334), .B1(R13[16]), .Y(n1028)
         );
  AOI22X1 U494 ( .A0(n1328), .A1(R3[16]), .B0(n886), .B1(R14[16]), .Y(n1029)
         );
  AOI22X1 U495 ( .A0(n1320), .A1(R0[16]), .B0(n1318), .B1(R15[16]), .Y(n1030)
         );
  AOI22X1 U496 ( .A0(n1309), .A1(R1[16]), .B0(n1312), .B1(R12[16]), .Y(n1031)
         );
endmodule


module fft ( clk, rst_n, data_in, data_out );
  input [33:0] data_in;
  output [33:0] data_out;
  input clk, rst_n;
  wire   s_p_flag, mux_flag, demux_flag, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37;
  wire   [2:0] rotation;
  wire   [135:0] data_1;
  wire   [135:0] data_2;
  wire   [135:0] data_4;
  wire   [135:0] data_3;

  ctrl ctrl0 ( .clk(clk), .rst_n(rst_n), .s_p_flag_in(s_p_flag), .mux_flag(
        mux_flag), .rotation(rotation), .demux_flag(demux_flag) );
  s_p s_p0 ( .clk(clk), .rst_n(rst_n), .data_in_1(data_in), .data_out_1(data_1), .s_p_flag_out(s_p_flag) );
  mux mux0 ( .mux_flag(mux_flag), .clk(clk), .rst_n(rst_n), .data_in_1(data_2), 
        .data_in_2(data_1), .data_out(data_3), .data_in_3_33_(n10), 
        .data_in_3_32_(n21), .data_in_3_31_(n2), .data_in_3_30_(data_4[30]), 
        .data_in_3_29_(data_4[29]), .data_in_3_28_(data_4[28]), 
        .data_in_3_27_(data_4[27]), .data_in_3_26_(data_4[26]), 
        .data_in_3_25_(data_4[25]), .data_in_3_24_(data_4[24]), 
        .data_in_3_23_(data_4[23]), .data_in_3_22_(data_4[22]), 
        .data_in_3_21_(data_4[21]), .data_in_3_20_(data_4[20]), 
        .data_in_3_19_(data_4[19]), .data_in_3_18_(data_4[18]), 
        .data_in_3_17_(data_4[17]), .data_in_3_16_(n23), .data_in_3_15_(
        data_4[15]), .data_in_3_14_(n27), .data_in_3_13_(n1), .data_in_3_12_(
        data_4[12]), .data_in_3_11_(n6), .data_in_3_10_(data_4[10]), 
        .data_in_3_9_(data_4[9]), .data_in_3_8_(data_4[8]), .data_in_3_7_(
        data_4[7]), .data_in_3_6_(data_4[6]), .data_in_3_5_(n36), 
        .data_in_3_4_(data_4[4]), .data_in_3_3_(data_4[3]), .data_in_3_2_(
        data_4[2]), .data_in_3_1_(data_4[1]), .data_in_3_0_(data_4[0]) );
  butterfly butterfly0 ( .calc_in(data_3), .rotation({n37, rotation[1:0]}), 
        .calc_out(data_4) );
  reg1 reg10 ( .clk(clk), .rst_n(rst_n), .data_in_2({n30, n17, n20, n19, 
        data_4[131], n13, data_4[129:119], n12, n9, data_4[116], n7, 
        data_4[114:102], n33, n31, n11, n15, data_4[97:85], n28, n25, n26, n16, 
        data_4[80:68], n32, n24, n5, n4, data_4[63], n29, data_4[61:51], n22, 
        n18, n14, data_4[47:46], n34, data_4[44:15], n8, data_4[13:12], n3, 
        data_4[10:6], n36, data_4[4:0]}), .reg_datain_flag(demux_flag), 
        .data_out_2(data_2) );
  p_s p_s0 ( .clk(clk), .rst_n(rst_n), .data_in_3({n30, n17, n20, n19, 
        data_4[131], n13, data_4[129:119], n12, n9, data_4[116], n7, 
        data_4[114:102], n33, n31, n11, n15, data_4[97:85], n28, n25, n26, n16, 
        data_4[80:68], n32, n24, n5, n4, data_4[63], n29, data_4[61:51], n22, 
        n18, n14, data_4[47:46], n34, data_4[44:15], n8, data_4[13:12], n3, 
        data_4[10:6], n36, data_4[4:0]}), .p_s_flag_in(demux_flag), 
        .data_out_3(data_out) );
  BUFX20 U1 ( .A(data_4[101]), .Y(n33) );
  BUFX20 U2 ( .A(data_4[132]), .Y(n19) );
  BUFX20 U3 ( .A(data_4[66]), .Y(n24) );
  BUFX20 U4 ( .A(data_4[118]), .Y(n12) );
  BUFX16 U5 ( .A(data_4[65]), .Y(n5) );
  BUFX20 U6 ( .A(data_4[67]), .Y(n32) );
  BUFX16 U7 ( .A(data_4[50]), .Y(n22) );
  BUFX20 U8 ( .A(data_4[117]), .Y(n9) );
  BUFX20 U9 ( .A(data_4[84]), .Y(n28) );
  BUFX16 U10 ( .A(data_4[115]), .Y(n7) );
  DLY1X1 U11 ( .A(data_4[16]), .Y(n23) );
  INVX8 U12 ( .A(n35), .Y(n36) );
  BUFX12 U13 ( .A(rotation[2]), .Y(n37) );
  BUFX12 U14 ( .A(data_4[62]), .Y(n29) );
  BUFX16 U15 ( .A(data_4[135]), .Y(n30) );
  BUFX16 U16 ( .A(data_4[98]), .Y(n15) );
  BUFX16 U17 ( .A(data_4[100]), .Y(n31) );
  BUFX16 U18 ( .A(data_4[134]), .Y(n17) );
  BUFX16 U19 ( .A(data_4[83]), .Y(n25) );
  BUFX12 U20 ( .A(data_4[133]), .Y(n20) );
  BUFX16 U21 ( .A(data_4[14]), .Y(n8) );
  BUFX3 U22 ( .A(n3), .Y(n6) );
  CLKINVX3 U23 ( .A(data_4[5]), .Y(n35) );
  CLKBUFX3 U24 ( .A(data_4[31]), .Y(n2) );
  BUFX3 U25 ( .A(data_4[32]), .Y(n21) );
  BUFX3 U26 ( .A(data_4[33]), .Y(n10) );
  BUFX3 U27 ( .A(n8), .Y(n27) );
  BUFX3 U28 ( .A(data_4[13]), .Y(n1) );
  BUFX16 U29 ( .A(data_4[11]), .Y(n3) );
  BUFX20 U30 ( .A(data_4[81]), .Y(n16) );
  BUFX20 U31 ( .A(data_4[82]), .Y(n26) );
  BUFX16 U32 ( .A(data_4[130]), .Y(n13) );
  BUFX16 U33 ( .A(data_4[49]), .Y(n18) );
  BUFX16 U34 ( .A(data_4[45]), .Y(n34) );
  BUFX16 U35 ( .A(data_4[48]), .Y(n14) );
  BUFX8 U36 ( .A(data_4[64]), .Y(n4) );
  BUFX12 U37 ( .A(data_4[99]), .Y(n11) );
endmodule


module fft_chip ( clk, rst_n, data_in, data_out );
  input [33:0] data_in;
  output [33:0] data_out;
  input clk, rst_n;
  wire   net_clk, net_rst_n;
  wire   [33:0] net_data_in;
  wire   [33:0] net_data_out;

  PIW PIW_clk ( .PAD(clk), .C(net_clk) );
  PIW PIW_rst_n ( .PAD(rst_n), .C(net_rst_n) );
  PIW PIW_data_in0 ( .PAD(data_in[0]), .C(net_data_in[0]) );
  PIW PIW_data_in1 ( .PAD(data_in[1]), .C(net_data_in[1]) );
  PIW PIW_data_in2 ( .PAD(data_in[2]), .C(net_data_in[2]) );
  PIW PIW_data_in3 ( .PAD(data_in[3]), .C(net_data_in[3]) );
  PIW PIW_data_in4 ( .PAD(data_in[4]), .C(net_data_in[4]) );
  PIW PIW_data_in5 ( .PAD(data_in[5]), .C(net_data_in[5]) );
  PIW PIW_data_in6 ( .PAD(data_in[6]), .C(net_data_in[6]) );
  PIW PIW_data_in7 ( .PAD(data_in[7]), .C(net_data_in[7]) );
  PIW PIW_data_in8 ( .PAD(data_in[8]), .C(net_data_in[8]) );
  PIW PIW_data_in9 ( .PAD(data_in[9]), .C(net_data_in[9]) );
  PIW PIW_data_in10 ( .PAD(data_in[10]), .C(net_data_in[10]) );
  PIW PIW_data_in11 ( .PAD(data_in[11]), .C(net_data_in[11]) );
  PIW PIW_data_in12 ( .PAD(data_in[12]), .C(net_data_in[12]) );
  PIW PIW_data_in13 ( .PAD(data_in[13]), .C(net_data_in[13]) );
  PIW PIW_data_in14 ( .PAD(data_in[14]), .C(net_data_in[14]) );
  PIW PIW_data_in15 ( .PAD(data_in[15]), .C(net_data_in[15]) );
  PIW PIW_data_in16 ( .PAD(data_in[16]), .C(net_data_in[16]) );
  PIW PIW_data_in17 ( .PAD(data_in[17]), .C(net_data_in[17]) );
  PIW PIW_data_in18 ( .PAD(data_in[18]), .C(net_data_in[18]) );
  PIW PIW_data_in19 ( .PAD(data_in[19]), .C(net_data_in[19]) );
  PIW PIW_data_in20 ( .PAD(data_in[20]), .C(net_data_in[20]) );
  PIW PIW_data_in21 ( .PAD(data_in[21]), .C(net_data_in[21]) );
  PIW PIW_data_in22 ( .PAD(data_in[22]), .C(net_data_in[22]) );
  PIW PIW_data_in23 ( .PAD(data_in[23]), .C(net_data_in[23]) );
  PIW PIW_data_in24 ( .PAD(data_in[24]), .C(net_data_in[24]) );
  PIW PIW_data_in25 ( .PAD(data_in[25]), .C(net_data_in[25]) );
  PIW PIW_data_in26 ( .PAD(data_in[26]), .C(net_data_in[26]) );
  PIW PIW_data_in27 ( .PAD(data_in[27]), .C(net_data_in[27]) );
  PIW PIW_data_in28 ( .PAD(data_in[28]), .C(net_data_in[28]) );
  PIW PIW_data_in29 ( .PAD(data_in[29]), .C(net_data_in[29]) );
  PIW PIW_data_in30 ( .PAD(data_in[30]), .C(net_data_in[30]) );
  PIW PIW_data_in31 ( .PAD(data_in[31]), .C(net_data_in[31]) );
  PIW PIW_data_in32 ( .PAD(data_in[32]), .C(net_data_in[32]) );
  PIW PIW_data_in33 ( .PAD(data_in[33]), .C(net_data_in[33]) );
  PO8W PO8W_data_out0 ( .I(net_data_out[0]), .PAD(data_out[0]) );
  PO8W PO8W_data_out1 ( .I(net_data_out[1]), .PAD(data_out[1]) );
  PO8W PO8W_data_out2 ( .I(net_data_out[2]), .PAD(data_out[2]) );
  PO8W PO8W_data_out3 ( .I(net_data_out[3]), .PAD(data_out[3]) );
  PO8W PO8W_data_out4 ( .I(net_data_out[4]), .PAD(data_out[4]) );
  PO8W PO8W_data_out5 ( .I(net_data_out[5]), .PAD(data_out[5]) );
  PO8W PO8W_data_out6 ( .I(net_data_out[6]), .PAD(data_out[6]) );
  PO8W PO8W_data_out7 ( .I(net_data_out[7]), .PAD(data_out[7]) );
  PO8W PO8W_data_out8 ( .I(net_data_out[8]), .PAD(data_out[8]) );
  PO8W PO8W_data_out9 ( .I(net_data_out[9]), .PAD(data_out[9]) );
  PO8W PO8W_data_out10 ( .I(net_data_out[10]), .PAD(data_out[10]) );
  PO8W PO8W_data_out11 ( .I(net_data_out[11]), .PAD(data_out[11]) );
  PO8W PO8W_data_out12 ( .I(net_data_out[12]), .PAD(data_out[12]) );
  PO8W PO8W_data_out13 ( .I(net_data_out[13]), .PAD(data_out[13]) );
  PO8W PO8W_data_out14 ( .I(net_data_out[14]), .PAD(data_out[14]) );
  PO8W PO8W_data_out15 ( .I(net_data_out[15]), .PAD(data_out[15]) );
  PO8W PO8W_data_out16 ( .I(net_data_out[16]), .PAD(data_out[16]) );
  PO8W PO8W_data_out17 ( .I(net_data_out[17]), .PAD(data_out[17]) );
  PO8W PO8W_data_out18 ( .I(net_data_out[18]), .PAD(data_out[18]) );
  PO8W PO8W_data_out19 ( .I(net_data_out[19]), .PAD(data_out[19]) );
  PO8W PO8W_data_out20 ( .I(net_data_out[20]), .PAD(data_out[20]) );
  PO8W PO8W_data_out21 ( .I(net_data_out[21]), .PAD(data_out[21]) );
  PO8W PO8W_data_out22 ( .I(net_data_out[22]), .PAD(data_out[22]) );
  PO8W PO8W_data_out23 ( .I(net_data_out[23]), .PAD(data_out[23]) );
  PO8W PO8W_data_out24 ( .I(net_data_out[24]), .PAD(data_out[24]) );
  PO8W PO8W_data_out25 ( .I(net_data_out[25]), .PAD(data_out[25]) );
  PO8W PO8W_data_out26 ( .I(net_data_out[26]), .PAD(data_out[26]) );
  PO8W PO8W_data_out27 ( .I(net_data_out[27]), .PAD(data_out[27]) );
  PO8W PO8W_data_out28 ( .I(net_data_out[28]), .PAD(data_out[28]) );
  PO8W PO8W_data_out29 ( .I(net_data_out[29]), .PAD(data_out[29]) );
  PO8W PO8W_data_out30 ( .I(net_data_out[30]), .PAD(data_out[30]) );
  PO8W PO8W_data_out31 ( .I(net_data_out[31]), .PAD(data_out[31]) );
  PO8W PO8W_data_out32 ( .I(net_data_out[32]), .PAD(data_out[32]) );
  PO8W PO8W_data_out33 ( .I(net_data_out[33]), .PAD(data_out[33]) );
  fft inst_fft ( .clk(net_clk), .rst_n(net_rst_n), .data_in(net_data_in), 
        .data_out(net_data_out) );
endmodule

