//**********************************************************
// Author: @VenciFreeman, copyright 2020
// e-mail: vencifreeman16@sjtu.edu.cn
// School: Shanghai Jiao Tong University
//
// File Name: butterfly
//
// Type: Combinational
//
// Purpose: <Specific Function Description>
// 
//
// Details:
//
//
// Release History:
// - Version 1.0 20/03/30: Create;
//
// Notes:
//
//**********************************************************

module mult(a_in, b_in, c_out)

  input a_in[16:0];
  input b_in[7:0];

  output c_out[16:0];

endmodule