
module ctrl ( clk, rst_n, s_p_flag_in, mux_flag, rotation, demux_flag );
  output [2:0] rotation;
  input clk, rst_n, s_p_flag_in;
  output mux_flag, demux_flag;
  wire   n7, n8, n9, N17, N18, N19, n3, n1, n6;
  wire   [2:0] core_tick;

  DFFRHQX4 mux_flag_reg ( .D(core_tick[2]), .CK(clk), .RN(rst_n), .Q(mux_flag)
         );
  DFFRHQX4 rotation_reg_2_ ( .D(core_tick[2]), .CK(clk), .RN(rst_n), .Q(n7) );
  DFFRHQX4 rotation_reg_1_ ( .D(core_tick[1]), .CK(clk), .RN(rst_n), .Q(n8) );
  DFFRHQX4 rotation_reg_0_ ( .D(core_tick[0]), .CK(clk), .RN(rst_n), .Q(n9) );
  DFFRHQX1 core_tick_reg_2_ ( .D(N19), .CK(clk), .RN(rst_n), .Q(core_tick[2])
         );
  DFFRHQX1 core_tick_reg_1_ ( .D(N18), .CK(clk), .RN(rst_n), .Q(core_tick[1])
         );
  DFFRHQX1 core_tick_reg_0_ ( .D(N17), .CK(clk), .RN(rst_n), .Q(core_tick[0])
         );
  DFFRHQX1 demux_flag_reg ( .D(n6), .CK(clk), .RN(rst_n), .Q(demux_flag) );
  BUFX16 U3 ( .A(n9), .Y(rotation[0]) );
  BUFX20 U4 ( .A(n7), .Y(rotation[2]) );
  BUFX16 U5 ( .A(n8), .Y(rotation[1]) );
  INVX1 U6 ( .A(core_tick[2]), .Y(n6) );
  AOI2BB1X1 U7 ( .A0N(n1), .A1N(core_tick[1]), .B0(core_tick[0]), .Y(N17) );
  OR2X2 U8 ( .A(s_p_flag_in), .B(core_tick[2]), .Y(n1) );
  XOR2X1 U9 ( .A(core_tick[1]), .B(core_tick[0]), .Y(N18) );
  XOR2X1 U10 ( .A(n6), .B(n3), .Y(N19) );
  NAND2X1 U11 ( .A(core_tick[1]), .B(core_tick[0]), .Y(n3) );
endmodule


module s_p ( clk, rst_n, data_in_1, data_out_1, s_p_flag_out );
  input [33:0] data_in_1;
  output [135:0] data_out_1;
  input clk, rst_n;
  output s_p_flag_out;
  wire   N13, N14, N15, N230, n550, n551, n552, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045;
  wire   [3:0] counter;
  wire   [33:0] R15;
  wire   [33:0] R11;
  wire   [33:0] R7;
  wire   [33:0] R3;
  wire   [33:0] R12;
  wire   [33:0] R8;
  wire   [33:0] R4;
  wire   [33:0] R0;
  wire   [33:0] R13;
  wire   [33:0] R9;
  wire   [33:0] R5;
  wire   [33:0] R1;
  wire   [33:0] R14;
  wire   [33:0] R10;
  wire   [33:0] R6;
  wire   [33:0] R2;

  DFFHQX4 data_out_1_reg_67_ ( .D(n900), .CK(clk), .Q(data_out_1[67]) );
  DFFHQX4 data_out_1_reg_64_ ( .D(n903), .CK(clk), .Q(data_out_1[64]) );
  DFFHQX4 data_out_1_reg_63_ ( .D(n904), .CK(clk), .Q(data_out_1[63]) );
  DFFHQX4 data_out_1_reg_62_ ( .D(n905), .CK(clk), .Q(data_out_1[62]) );
  DFFHQX4 data_out_1_reg_61_ ( .D(n906), .CK(clk), .Q(data_out_1[61]) );
  DFFHQX4 data_out_1_reg_60_ ( .D(n907), .CK(clk), .Q(data_out_1[60]) );
  DFFHQX4 data_out_1_reg_59_ ( .D(n908), .CK(clk), .Q(data_out_1[59]) );
  DFFHQX4 data_out_1_reg_58_ ( .D(n909), .CK(clk), .Q(data_out_1[58]) );
  DFFHQX4 data_out_1_reg_56_ ( .D(n911), .CK(clk), .Q(data_out_1[56]) );
  DFFHQX4 data_out_1_reg_55_ ( .D(n912), .CK(clk), .Q(data_out_1[55]) );
  DFFHQX4 data_out_1_reg_51_ ( .D(n916), .CK(clk), .Q(data_out_1[51]) );
  DFFHQX4 data_out_1_reg_50_ ( .D(n917), .CK(clk), .Q(data_out_1[50]) );
  DFFHQX4 data_out_1_reg_101_ ( .D(n866), .CK(clk), .Q(data_out_1[101]) );
  DFFHQX4 data_out_1_reg_94_ ( .D(n873), .CK(clk), .Q(data_out_1[94]) );
  DFFHQX4 data_out_1_reg_85_ ( .D(n882), .CK(clk), .Q(data_out_1[85]) );
  DFFHQX4 data_out_1_reg_84_ ( .D(n883), .CK(clk), .Q(data_out_1[84]) );
  DFFHQX4 data_out_1_reg_73_ ( .D(n894), .CK(clk), .Q(data_out_1[73]) );
  DFFHQX4 data_out_1_reg_71_ ( .D(n896), .CK(clk), .Q(data_out_1[71]) );
  DFFHQX4 data_out_1_reg_69_ ( .D(n898), .CK(clk), .Q(data_out_1[69]) );
  DFFHQX4 data_out_1_reg_68_ ( .D(n899), .CK(clk), .Q(data_out_1[68]) );
  DFFHQX4 data_out_1_reg_130_ ( .D(n837), .CK(clk), .Q(data_out_1[130]) );
  DFFHQX4 data_out_1_reg_129_ ( .D(n838), .CK(clk), .Q(data_out_1[129]) );
  DFFHQX4 data_out_1_reg_128_ ( .D(n839), .CK(clk), .Q(data_out_1[128]) );
  DFFHQX4 data_out_1_reg_127_ ( .D(n840), .CK(clk), .Q(data_out_1[127]) );
  DFFHQX4 data_out_1_reg_126_ ( .D(n841), .CK(clk), .Q(data_out_1[126]) );
  DFFHQX4 data_out_1_reg_125_ ( .D(n842), .CK(clk), .Q(data_out_1[125]) );
  DFFHQX4 data_out_1_reg_124_ ( .D(n843), .CK(clk), .Q(data_out_1[124]) );
  DFFHQX4 data_out_1_reg_123_ ( .D(n844), .CK(clk), .Q(data_out_1[123]) );
  DFFHQX4 data_out_1_reg_122_ ( .D(n845), .CK(clk), .Q(data_out_1[122]) );
  DFFHQX4 data_out_1_reg_120_ ( .D(n847), .CK(clk), .Q(data_out_1[120]) );
  DFFHQX4 data_out_1_reg_119_ ( .D(n848), .CK(clk), .Q(data_out_1[119]) );
  DFFHQX4 data_out_1_reg_118_ ( .D(n849), .CK(clk), .Q(data_out_1[118]) );
  DFFHQX4 data_out_1_reg_114_ ( .D(n853), .CK(clk), .Q(data_out_1[114]) );
  DFFHQX4 data_out_1_reg_113_ ( .D(n854), .CK(clk), .Q(data_out_1[113]) );
  DFFHQX4 data_out_1_reg_112_ ( .D(n855), .CK(clk), .Q(data_out_1[112]) );
  DFFHQX4 data_out_1_reg_111_ ( .D(n856), .CK(clk), .Q(data_out_1[111]) );
  DFFHQX4 data_out_1_reg_110_ ( .D(n857), .CK(clk), .Q(data_out_1[110]) );
  DFFHQX4 data_out_1_reg_109_ ( .D(n858), .CK(clk), .Q(data_out_1[109]) );
  DFFHQX4 data_out_1_reg_108_ ( .D(n859), .CK(clk), .Q(data_out_1[108]) );
  DFFHQX4 data_out_1_reg_107_ ( .D(n860), .CK(clk), .Q(data_out_1[107]) );
  DFFHQX4 data_out_1_reg_106_ ( .D(n861), .CK(clk), .Q(data_out_1[106]) );
  DFFHQX4 data_out_1_reg_105_ ( .D(n862), .CK(clk), .Q(data_out_1[105]) );
  DFFHQX4 data_out_1_reg_102_ ( .D(n865), .CK(clk), .Q(data_out_1[102]) );
  EDFFX1 R13_reg_33_ ( .D(data_in_1[33]), .E(n969), .CK(clk), .Q(R13[33]) );
  EDFFX1 R13_reg_32_ ( .D(data_in_1[32]), .E(n1011), .CK(clk), .Q(R13[32]) );
  EDFFX1 R13_reg_31_ ( .D(data_in_1[31]), .E(n1010), .CK(clk), .Q(R13[31]) );
  EDFFX1 R13_reg_30_ ( .D(data_in_1[30]), .E(n969), .CK(clk), .Q(R13[30]) );
  EDFFX1 R13_reg_29_ ( .D(data_in_1[29]), .E(n1011), .CK(clk), .Q(R13[29]) );
  EDFFX1 R13_reg_28_ ( .D(data_in_1[28]), .E(n1010), .CK(clk), .Q(R13[28]) );
  EDFFX1 R13_reg_27_ ( .D(data_in_1[27]), .E(n969), .CK(clk), .Q(R13[27]) );
  EDFFX1 R13_reg_26_ ( .D(data_in_1[26]), .E(n1011), .CK(clk), .Q(R13[26]) );
  EDFFX1 R13_reg_25_ ( .D(data_in_1[25]), .E(n969), .CK(clk), .Q(R13[25]) );
  EDFFX1 R13_reg_24_ ( .D(data_in_1[24]), .E(n1010), .CK(clk), .Q(R13[24]) );
  EDFFX1 R13_reg_23_ ( .D(data_in_1[23]), .E(n1011), .CK(clk), .Q(R13[23]) );
  EDFFX1 R13_reg_22_ ( .D(data_in_1[22]), .E(n1009), .CK(clk), .Q(R13[22]) );
  EDFFX1 R13_reg_21_ ( .D(data_in_1[21]), .E(n1010), .CK(clk), .Q(R13[21]) );
  EDFFX1 R13_reg_20_ ( .D(data_in_1[20]), .E(n1011), .CK(clk), .Q(R13[20]) );
  EDFFX1 R13_reg_19_ ( .D(data_in_1[19]), .E(n969), .CK(clk), .Q(R13[19]) );
  EDFFX1 R13_reg_18_ ( .D(data_in_1[18]), .E(n1010), .CK(clk), .Q(R13[18]) );
  EDFFX1 R13_reg_17_ ( .D(data_in_1[17]), .E(n1010), .CK(clk), .Q(R13[17]) );
  EDFFX1 R13_reg_16_ ( .D(data_in_1[16]), .E(n1009), .CK(clk), .Q(R13[16]) );
  EDFFX1 R13_reg_15_ ( .D(data_in_1[15]), .E(n969), .CK(clk), .Q(R13[15]) );
  EDFFX1 R13_reg_14_ ( .D(data_in_1[14]), .E(n1011), .CK(clk), .Q(R13[14]) );
  EDFFX1 R13_reg_13_ ( .D(data_in_1[13]), .E(n969), .CK(clk), .Q(R13[13]) );
  EDFFX1 R13_reg_12_ ( .D(data_in_1[12]), .E(n1010), .CK(clk), .Q(R13[12]) );
  EDFFX1 R13_reg_11_ ( .D(data_in_1[11]), .E(n1011), .CK(clk), .Q(R13[11]) );
  EDFFX1 R13_reg_10_ ( .D(data_in_1[10]), .E(n1009), .CK(clk), .Q(R13[10]) );
  EDFFX1 R13_reg_9_ ( .D(data_in_1[9]), .E(n1011), .CK(clk), .Q(R13[9]) );
  EDFFX1 R13_reg_8_ ( .D(data_in_1[8]), .E(n1009), .CK(clk), .Q(R13[8]) );
  EDFFX1 R13_reg_7_ ( .D(data_in_1[7]), .E(n1009), .CK(clk), .Q(R13[7]) );
  EDFFX1 R13_reg_6_ ( .D(data_in_1[6]), .E(n1009), .CK(clk), .Q(R13[6]) );
  EDFFX1 R13_reg_5_ ( .D(data_in_1[5]), .E(n1010), .CK(clk), .Q(R13[5]) );
  EDFFX1 R13_reg_4_ ( .D(data_in_1[4]), .E(n1009), .CK(clk), .Q(R13[4]) );
  EDFFX1 R13_reg_3_ ( .D(data_in_1[3]), .E(n1009), .CK(clk), .Q(R13[3]) );
  EDFFX1 R13_reg_2_ ( .D(data_in_1[2]), .E(n1010), .CK(clk), .Q(R13[2]) );
  EDFFX1 R13_reg_1_ ( .D(data_in_1[1]), .E(n969), .CK(clk), .Q(R13[1]) );
  EDFFX1 R13_reg_0_ ( .D(data_in_1[0]), .E(n1009), .CK(clk), .Q(R13[0]) );
  EDFFX1 R1_reg_33_ ( .D(data_in_1[33]), .E(n979), .CK(clk), .Q(R1[33]) );
  EDFFX1 R1_reg_32_ ( .D(data_in_1[32]), .E(n979), .CK(clk), .Q(R1[32]) );
  EDFFX1 R1_reg_31_ ( .D(data_in_1[31]), .E(n979), .CK(clk), .Q(R1[31]) );
  EDFFX1 R1_reg_30_ ( .D(data_in_1[30]), .E(n979), .CK(clk), .Q(R1[30]) );
  EDFFX1 R1_reg_29_ ( .D(data_in_1[29]), .E(n979), .CK(clk), .Q(R1[29]) );
  EDFFX1 R1_reg_28_ ( .D(data_in_1[28]), .E(n979), .CK(clk), .Q(R1[28]) );
  EDFFX1 R1_reg_27_ ( .D(data_in_1[27]), .E(n979), .CK(clk), .Q(R1[27]) );
  EDFFX1 R1_reg_26_ ( .D(data_in_1[26]), .E(n979), .CK(clk), .Q(R1[26]) );
  EDFFX1 R1_reg_25_ ( .D(data_in_1[25]), .E(n979), .CK(clk), .Q(R1[25]) );
  EDFFX1 R1_reg_24_ ( .D(data_in_1[24]), .E(n979), .CK(clk), .Q(R1[24]) );
  EDFFX1 R1_reg_23_ ( .D(data_in_1[23]), .E(n979), .CK(clk), .Q(R1[23]) );
  EDFFX1 R1_reg_22_ ( .D(data_in_1[22]), .E(n979), .CK(clk), .Q(R1[22]) );
  EDFFX1 R1_reg_21_ ( .D(data_in_1[21]), .E(n980), .CK(clk), .Q(R1[21]) );
  EDFFX1 R1_reg_20_ ( .D(data_in_1[20]), .E(n980), .CK(clk), .Q(R1[20]) );
  EDFFX1 R1_reg_19_ ( .D(data_in_1[19]), .E(n980), .CK(clk), .Q(R1[19]) );
  EDFFX1 R1_reg_18_ ( .D(data_in_1[18]), .E(n980), .CK(clk), .Q(R1[18]) );
  EDFFX1 R1_reg_17_ ( .D(data_in_1[17]), .E(n980), .CK(clk), .Q(R1[17]) );
  EDFFX1 R1_reg_16_ ( .D(data_in_1[16]), .E(n980), .CK(clk), .Q(R1[16]) );
  EDFFX1 R1_reg_15_ ( .D(data_in_1[15]), .E(n980), .CK(clk), .Q(R1[15]) );
  EDFFX1 R1_reg_14_ ( .D(data_in_1[14]), .E(n980), .CK(clk), .Q(R1[14]) );
  EDFFX1 R1_reg_13_ ( .D(data_in_1[13]), .E(n980), .CK(clk), .Q(R1[13]) );
  EDFFX1 R1_reg_12_ ( .D(data_in_1[12]), .E(n980), .CK(clk), .Q(R1[12]) );
  EDFFX1 R1_reg_11_ ( .D(data_in_1[11]), .E(n980), .CK(clk), .Q(R1[11]) );
  EDFFX1 R1_reg_10_ ( .D(data_in_1[10]), .E(n980), .CK(clk), .Q(R1[10]) );
  EDFFX1 R1_reg_9_ ( .D(data_in_1[9]), .E(n979), .CK(clk), .Q(R1[9]) );
  EDFFX1 R1_reg_8_ ( .D(data_in_1[8]), .E(n980), .CK(clk), .Q(R1[8]) );
  EDFFX1 R1_reg_7_ ( .D(data_in_1[7]), .E(n979), .CK(clk), .Q(R1[7]) );
  EDFFX1 R1_reg_6_ ( .D(data_in_1[6]), .E(n980), .CK(clk), .Q(R1[6]) );
  EDFFX1 R1_reg_5_ ( .D(data_in_1[5]), .E(n979), .CK(clk), .Q(R1[5]) );
  EDFFX1 R1_reg_4_ ( .D(data_in_1[4]), .E(n980), .CK(clk), .Q(R1[4]) );
  EDFFX1 R1_reg_3_ ( .D(data_in_1[3]), .E(n979), .CK(clk), .Q(R1[3]) );
  EDFFX1 R1_reg_2_ ( .D(data_in_1[2]), .E(n980), .CK(clk), .Q(R1[2]) );
  EDFFX1 R1_reg_1_ ( .D(data_in_1[1]), .E(n979), .CK(clk), .Q(R1[1]) );
  EDFFX1 R1_reg_0_ ( .D(data_in_1[0]), .E(n980), .CK(clk), .Q(R1[0]) );
  EDFFX1 R5_reg_33_ ( .D(data_in_1[33]), .E(n987), .CK(clk), .Q(R5[33]) );
  EDFFX1 R5_reg_32_ ( .D(data_in_1[32]), .E(n987), .CK(clk), .Q(R5[32]) );
  EDFFX1 R5_reg_31_ ( .D(data_in_1[31]), .E(n987), .CK(clk), .Q(R5[31]) );
  EDFFX1 R5_reg_30_ ( .D(data_in_1[30]), .E(n987), .CK(clk), .Q(R5[30]) );
  EDFFX1 R5_reg_29_ ( .D(data_in_1[29]), .E(n987), .CK(clk), .Q(R5[29]) );
  EDFFX1 R5_reg_28_ ( .D(data_in_1[28]), .E(n987), .CK(clk), .Q(R5[28]) );
  EDFFX1 R5_reg_27_ ( .D(data_in_1[27]), .E(n987), .CK(clk), .Q(R5[27]) );
  EDFFX1 R5_reg_26_ ( .D(data_in_1[26]), .E(n987), .CK(clk), .Q(R5[26]) );
  EDFFX1 R5_reg_25_ ( .D(data_in_1[25]), .E(n987), .CK(clk), .Q(R5[25]) );
  EDFFX1 R5_reg_24_ ( .D(data_in_1[24]), .E(n987), .CK(clk), .Q(R5[24]) );
  EDFFX1 R5_reg_23_ ( .D(data_in_1[23]), .E(n987), .CK(clk), .Q(R5[23]) );
  EDFFX1 R5_reg_22_ ( .D(data_in_1[22]), .E(n987), .CK(clk), .Q(R5[22]) );
  EDFFX1 R5_reg_21_ ( .D(data_in_1[21]), .E(n988), .CK(clk), .Q(R5[21]) );
  EDFFX1 R5_reg_20_ ( .D(data_in_1[20]), .E(n988), .CK(clk), .Q(R5[20]) );
  EDFFX1 R5_reg_19_ ( .D(data_in_1[19]), .E(n988), .CK(clk), .Q(R5[19]) );
  EDFFX1 R5_reg_18_ ( .D(data_in_1[18]), .E(n988), .CK(clk), .Q(R5[18]) );
  EDFFX1 R5_reg_17_ ( .D(data_in_1[17]), .E(n988), .CK(clk), .Q(R5[17]) );
  EDFFX1 R5_reg_16_ ( .D(data_in_1[16]), .E(n988), .CK(clk), .Q(R5[16]) );
  EDFFX1 R5_reg_15_ ( .D(data_in_1[15]), .E(n988), .CK(clk), .Q(R5[15]) );
  EDFFX1 R5_reg_14_ ( .D(data_in_1[14]), .E(n988), .CK(clk), .Q(R5[14]) );
  EDFFX1 R5_reg_13_ ( .D(data_in_1[13]), .E(n988), .CK(clk), .Q(R5[13]) );
  EDFFX1 R5_reg_12_ ( .D(data_in_1[12]), .E(n988), .CK(clk), .Q(R5[12]) );
  EDFFX1 R5_reg_11_ ( .D(data_in_1[11]), .E(n988), .CK(clk), .Q(R5[11]) );
  EDFFX1 R5_reg_10_ ( .D(data_in_1[10]), .E(n988), .CK(clk), .Q(R5[10]) );
  EDFFX1 R5_reg_9_ ( .D(data_in_1[9]), .E(n987), .CK(clk), .Q(R5[9]) );
  EDFFX1 R5_reg_8_ ( .D(data_in_1[8]), .E(n988), .CK(clk), .Q(R5[8]) );
  EDFFX1 R5_reg_7_ ( .D(data_in_1[7]), .E(n987), .CK(clk), .Q(R5[7]) );
  EDFFX1 R5_reg_6_ ( .D(data_in_1[6]), .E(n988), .CK(clk), .Q(R5[6]) );
  EDFFX1 R5_reg_5_ ( .D(data_in_1[5]), .E(n987), .CK(clk), .Q(R5[5]) );
  EDFFX1 R5_reg_4_ ( .D(data_in_1[4]), .E(n988), .CK(clk), .Q(R5[4]) );
  EDFFX1 R5_reg_3_ ( .D(data_in_1[3]), .E(n987), .CK(clk), .Q(R5[3]) );
  EDFFX1 R5_reg_2_ ( .D(data_in_1[2]), .E(n988), .CK(clk), .Q(R5[2]) );
  EDFFX1 R5_reg_1_ ( .D(data_in_1[1]), .E(n987), .CK(clk), .Q(R5[1]) );
  EDFFX1 R5_reg_0_ ( .D(data_in_1[0]), .E(n988), .CK(clk), .Q(R5[0]) );
  EDFFX1 R9_reg_33_ ( .D(data_in_1[33]), .E(n973), .CK(clk), .Q(R9[33]) );
  EDFFX1 R9_reg_32_ ( .D(data_in_1[32]), .E(n973), .CK(clk), .Q(R9[32]) );
  EDFFX1 R9_reg_31_ ( .D(data_in_1[31]), .E(n973), .CK(clk), .Q(R9[31]) );
  EDFFX1 R9_reg_30_ ( .D(data_in_1[30]), .E(n973), .CK(clk), .Q(R9[30]) );
  EDFFX1 R9_reg_29_ ( .D(data_in_1[29]), .E(n973), .CK(clk), .Q(R9[29]) );
  EDFFX1 R9_reg_28_ ( .D(data_in_1[28]), .E(n973), .CK(clk), .Q(R9[28]) );
  EDFFX1 R9_reg_27_ ( .D(data_in_1[27]), .E(n973), .CK(clk), .Q(R9[27]) );
  EDFFX1 R9_reg_26_ ( .D(data_in_1[26]), .E(n973), .CK(clk), .Q(R9[26]) );
  EDFFX1 R9_reg_25_ ( .D(data_in_1[25]), .E(n997), .CK(clk), .Q(R9[25]) );
  EDFFX1 R9_reg_24_ ( .D(data_in_1[24]), .E(n996), .CK(clk), .Q(R9[24]) );
  EDFFX1 R9_reg_23_ ( .D(data_in_1[23]), .E(n997), .CK(clk), .Q(R9[23]) );
  EDFFX1 R9_reg_22_ ( .D(data_in_1[22]), .E(n997), .CK(clk), .Q(R9[22]) );
  EDFFX1 R9_reg_21_ ( .D(data_in_1[21]), .E(n996), .CK(clk), .Q(R9[21]) );
  EDFFX1 R9_reg_20_ ( .D(data_in_1[20]), .E(n996), .CK(clk), .Q(R9[20]) );
  EDFFX1 R9_reg_19_ ( .D(data_in_1[19]), .E(n996), .CK(clk), .Q(R9[19]) );
  EDFFX1 R9_reg_18_ ( .D(data_in_1[18]), .E(n996), .CK(clk), .Q(R9[18]) );
  EDFFX1 R9_reg_17_ ( .D(data_in_1[17]), .E(n996), .CK(clk), .Q(R9[17]) );
  EDFFX1 R9_reg_16_ ( .D(data_in_1[16]), .E(n996), .CK(clk), .Q(R9[16]) );
  EDFFX1 R9_reg_15_ ( .D(data_in_1[15]), .E(n996), .CK(clk), .Q(R9[15]) );
  EDFFX1 R9_reg_14_ ( .D(data_in_1[14]), .E(n996), .CK(clk), .Q(R9[14]) );
  EDFFX1 R9_reg_13_ ( .D(data_in_1[13]), .E(n996), .CK(clk), .Q(R9[13]) );
  EDFFX1 R9_reg_12_ ( .D(data_in_1[12]), .E(n996), .CK(clk), .Q(R9[12]) );
  EDFFX1 R9_reg_11_ ( .D(data_in_1[11]), .E(n996), .CK(clk), .Q(R9[11]) );
  EDFFX1 R9_reg_10_ ( .D(data_in_1[10]), .E(n996), .CK(clk), .Q(R9[10]) );
  EDFFX1 R9_reg_9_ ( .D(data_in_1[9]), .E(n997), .CK(clk), .Q(R9[9]) );
  EDFFX1 R9_reg_8_ ( .D(data_in_1[8]), .E(n997), .CK(clk), .Q(R9[8]) );
  EDFFX1 R9_reg_7_ ( .D(data_in_1[7]), .E(n997), .CK(clk), .Q(R9[7]) );
  EDFFX1 R9_reg_6_ ( .D(data_in_1[6]), .E(n997), .CK(clk), .Q(R9[6]) );
  EDFFX1 R9_reg_5_ ( .D(data_in_1[5]), .E(n997), .CK(clk), .Q(R9[5]) );
  EDFFX1 R9_reg_4_ ( .D(data_in_1[4]), .E(n997), .CK(clk), .Q(R9[4]) );
  EDFFX1 R9_reg_3_ ( .D(data_in_1[3]), .E(n997), .CK(clk), .Q(R9[3]) );
  EDFFX1 R9_reg_2_ ( .D(data_in_1[2]), .E(n997), .CK(clk), .Q(R9[2]) );
  EDFFX1 R9_reg_1_ ( .D(data_in_1[1]), .E(n997), .CK(clk), .Q(R9[1]) );
  EDFFX1 R9_reg_0_ ( .D(data_in_1[0]), .E(n997), .CK(clk), .Q(R9[0]) );
  EDFFX1 R14_reg_33_ ( .D(data_in_1[33]), .E(n1016), .CK(clk), .Q(R14[33]) );
  EDFFX1 R14_reg_32_ ( .D(data_in_1[32]), .E(n1016), .CK(clk), .Q(R14[32]) );
  EDFFX1 R14_reg_31_ ( .D(data_in_1[31]), .E(n1016), .CK(clk), .Q(R14[31]) );
  EDFFX1 R14_reg_30_ ( .D(data_in_1[30]), .E(n1016), .CK(clk), .Q(R14[30]) );
  EDFFX1 R14_reg_29_ ( .D(data_in_1[29]), .E(n1016), .CK(clk), .Q(R14[29]) );
  EDFFX1 R14_reg_28_ ( .D(data_in_1[28]), .E(n1016), .CK(clk), .Q(R14[28]) );
  EDFFX1 R14_reg_27_ ( .D(data_in_1[27]), .E(n1016), .CK(clk), .Q(R14[27]) );
  EDFFX1 R14_reg_26_ ( .D(data_in_1[26]), .E(n1016), .CK(clk), .Q(R14[26]) );
  EDFFX1 R14_reg_25_ ( .D(data_in_1[25]), .E(n1015), .CK(clk), .Q(R14[25]) );
  EDFFX1 R14_reg_24_ ( .D(data_in_1[24]), .E(n968), .CK(clk), .Q(R14[24]) );
  EDFFX1 R14_reg_23_ ( .D(data_in_1[23]), .E(n1013), .CK(clk), .Q(R14[23]) );
  EDFFX1 R14_reg_22_ ( .D(data_in_1[22]), .E(n1016), .CK(clk), .Q(R14[22]) );
  EDFFX1 R14_reg_21_ ( .D(data_in_1[21]), .E(n1015), .CK(clk), .Q(R14[21]) );
  EDFFX1 R14_reg_20_ ( .D(data_in_1[20]), .E(n968), .CK(clk), .Q(R14[20]) );
  EDFFX1 R14_reg_19_ ( .D(data_in_1[19]), .E(n1016), .CK(clk), .Q(R14[19]) );
  EDFFX1 R14_reg_18_ ( .D(data_in_1[18]), .E(n1016), .CK(clk), .Q(R14[18]) );
  EDFFX1 R14_reg_17_ ( .D(data_in_1[17]), .E(n968), .CK(clk), .Q(R14[17]) );
  EDFFX1 R14_reg_16_ ( .D(data_in_1[16]), .E(n1015), .CK(clk), .Q(R14[16]) );
  EDFFX1 R14_reg_15_ ( .D(data_in_1[15]), .E(n1016), .CK(clk), .Q(R14[15]) );
  EDFFX1 R14_reg_14_ ( .D(data_in_1[14]), .E(n1016), .CK(clk), .Q(R14[14]) );
  EDFFX1 R14_reg_13_ ( .D(data_in_1[13]), .E(n968), .CK(clk), .Q(R14[13]) );
  EDFFX1 R14_reg_12_ ( .D(data_in_1[12]), .E(n1015), .CK(clk), .Q(R14[12]) );
  EDFFX1 R14_reg_11_ ( .D(data_in_1[11]), .E(n1016), .CK(clk), .Q(R14[11]) );
  EDFFX1 R14_reg_10_ ( .D(data_in_1[10]), .E(n1015), .CK(clk), .Q(R14[10]) );
  EDFFX1 R14_reg_9_ ( .D(data_in_1[9]), .E(n968), .CK(clk), .Q(R14[9]) );
  EDFFX1 R14_reg_8_ ( .D(data_in_1[8]), .E(n1015), .CK(clk), .Q(R14[8]) );
  EDFFX1 R14_reg_7_ ( .D(data_in_1[7]), .E(n1016), .CK(clk), .Q(R14[7]) );
  EDFFX1 R14_reg_6_ ( .D(data_in_1[6]), .E(n1013), .CK(clk), .Q(R14[6]) );
  EDFFX1 R14_reg_5_ ( .D(data_in_1[5]), .E(n968), .CK(clk), .Q(R14[5]) );
  EDFFX1 R14_reg_4_ ( .D(data_in_1[4]), .E(n1015), .CK(clk), .Q(R14[4]) );
  EDFFX1 R14_reg_3_ ( .D(data_in_1[3]), .E(n1014), .CK(clk), .Q(R14[3]) );
  EDFFX1 R14_reg_2_ ( .D(data_in_1[2]), .E(n1016), .CK(clk), .Q(R14[2]) );
  EDFFX1 R14_reg_1_ ( .D(data_in_1[1]), .E(n1014), .CK(clk), .Q(R14[1]) );
  EDFFX1 R14_reg_0_ ( .D(data_in_1[0]), .E(n1014), .CK(clk), .Q(R14[0]) );
  EDFFX1 R2_reg_33_ ( .D(data_in_1[33]), .E(n981), .CK(clk), .Q(R2[33]) );
  EDFFX1 R2_reg_32_ ( .D(data_in_1[32]), .E(n981), .CK(clk), .Q(R2[32]) );
  EDFFX1 R2_reg_31_ ( .D(data_in_1[31]), .E(n981), .CK(clk), .Q(R2[31]) );
  EDFFX1 R2_reg_30_ ( .D(data_in_1[30]), .E(n981), .CK(clk), .Q(R2[30]) );
  EDFFX1 R2_reg_29_ ( .D(data_in_1[29]), .E(n981), .CK(clk), .Q(R2[29]) );
  EDFFX1 R2_reg_28_ ( .D(data_in_1[28]), .E(n981), .CK(clk), .Q(R2[28]) );
  EDFFX1 R2_reg_27_ ( .D(data_in_1[27]), .E(n981), .CK(clk), .Q(R2[27]) );
  EDFFX1 R2_reg_26_ ( .D(data_in_1[26]), .E(n981), .CK(clk), .Q(R2[26]) );
  EDFFX1 R2_reg_25_ ( .D(data_in_1[25]), .E(n981), .CK(clk), .Q(R2[25]) );
  EDFFX1 R2_reg_24_ ( .D(data_in_1[24]), .E(n981), .CK(clk), .Q(R2[24]) );
  EDFFX1 R2_reg_23_ ( .D(data_in_1[23]), .E(n981), .CK(clk), .Q(R2[23]) );
  EDFFX1 R2_reg_22_ ( .D(data_in_1[22]), .E(n981), .CK(clk), .Q(R2[22]) );
  EDFFX1 R2_reg_21_ ( .D(data_in_1[21]), .E(n982), .CK(clk), .Q(R2[21]) );
  EDFFX1 R2_reg_20_ ( .D(data_in_1[20]), .E(n982), .CK(clk), .Q(R2[20]) );
  EDFFX1 R2_reg_19_ ( .D(data_in_1[19]), .E(n982), .CK(clk), .Q(R2[19]) );
  EDFFX1 R2_reg_18_ ( .D(data_in_1[18]), .E(n982), .CK(clk), .Q(R2[18]) );
  EDFFX1 R2_reg_17_ ( .D(data_in_1[17]), .E(n982), .CK(clk), .Q(R2[17]) );
  EDFFX1 R2_reg_16_ ( .D(data_in_1[16]), .E(n982), .CK(clk), .Q(R2[16]) );
  EDFFX1 R2_reg_15_ ( .D(data_in_1[15]), .E(n982), .CK(clk), .Q(R2[15]) );
  EDFFX1 R2_reg_14_ ( .D(data_in_1[14]), .E(n982), .CK(clk), .Q(R2[14]) );
  EDFFX1 R2_reg_13_ ( .D(data_in_1[13]), .E(n982), .CK(clk), .Q(R2[13]) );
  EDFFX1 R2_reg_12_ ( .D(data_in_1[12]), .E(n982), .CK(clk), .Q(R2[12]) );
  EDFFX1 R2_reg_11_ ( .D(data_in_1[11]), .E(n982), .CK(clk), .Q(R2[11]) );
  EDFFX1 R2_reg_10_ ( .D(data_in_1[10]), .E(n982), .CK(clk), .Q(R2[10]) );
  EDFFX1 R2_reg_9_ ( .D(data_in_1[9]), .E(n981), .CK(clk), .Q(R2[9]) );
  EDFFX1 R2_reg_8_ ( .D(data_in_1[8]), .E(n982), .CK(clk), .Q(R2[8]) );
  EDFFX1 R2_reg_7_ ( .D(data_in_1[7]), .E(n981), .CK(clk), .Q(R2[7]) );
  EDFFX1 R2_reg_6_ ( .D(data_in_1[6]), .E(n982), .CK(clk), .Q(R2[6]) );
  EDFFX1 R2_reg_5_ ( .D(data_in_1[5]), .E(n981), .CK(clk), .Q(R2[5]) );
  EDFFX1 R2_reg_4_ ( .D(data_in_1[4]), .E(n982), .CK(clk), .Q(R2[4]) );
  EDFFX1 R2_reg_3_ ( .D(data_in_1[3]), .E(n981), .CK(clk), .Q(R2[3]) );
  EDFFX1 R2_reg_2_ ( .D(data_in_1[2]), .E(n982), .CK(clk), .Q(R2[2]) );
  EDFFX1 R2_reg_1_ ( .D(data_in_1[1]), .E(n981), .CK(clk), .Q(R2[1]) );
  EDFFX1 R2_reg_0_ ( .D(data_in_1[0]), .E(n982), .CK(clk), .Q(R2[0]) );
  EDFFX1 R6_reg_33_ ( .D(data_in_1[33]), .E(n989), .CK(clk), .Q(R6[33]) );
  EDFFX1 R6_reg_32_ ( .D(data_in_1[32]), .E(n989), .CK(clk), .Q(R6[32]) );
  EDFFX1 R6_reg_31_ ( .D(data_in_1[31]), .E(n989), .CK(clk), .Q(R6[31]) );
  EDFFX1 R6_reg_30_ ( .D(data_in_1[30]), .E(n989), .CK(clk), .Q(R6[30]) );
  EDFFX1 R6_reg_29_ ( .D(data_in_1[29]), .E(n989), .CK(clk), .Q(R6[29]) );
  EDFFX1 R6_reg_28_ ( .D(data_in_1[28]), .E(n989), .CK(clk), .Q(R6[28]) );
  EDFFX1 R6_reg_27_ ( .D(data_in_1[27]), .E(n989), .CK(clk), .Q(R6[27]) );
  EDFFX1 R6_reg_26_ ( .D(data_in_1[26]), .E(n989), .CK(clk), .Q(R6[26]) );
  EDFFX1 R6_reg_25_ ( .D(data_in_1[25]), .E(n989), .CK(clk), .Q(R6[25]) );
  EDFFX1 R6_reg_24_ ( .D(data_in_1[24]), .E(n989), .CK(clk), .Q(R6[24]) );
  EDFFX1 R6_reg_23_ ( .D(data_in_1[23]), .E(n989), .CK(clk), .Q(R6[23]) );
  EDFFX1 R6_reg_22_ ( .D(data_in_1[22]), .E(n989), .CK(clk), .Q(R6[22]) );
  EDFFX1 R6_reg_21_ ( .D(data_in_1[21]), .E(n990), .CK(clk), .Q(R6[21]) );
  EDFFX1 R6_reg_20_ ( .D(data_in_1[20]), .E(n990), .CK(clk), .Q(R6[20]) );
  EDFFX1 R6_reg_19_ ( .D(data_in_1[19]), .E(n990), .CK(clk), .Q(R6[19]) );
  EDFFX1 R6_reg_18_ ( .D(data_in_1[18]), .E(n990), .CK(clk), .Q(R6[18]) );
  EDFFX1 R6_reg_17_ ( .D(data_in_1[17]), .E(n990), .CK(clk), .Q(R6[17]) );
  EDFFX1 R6_reg_16_ ( .D(data_in_1[16]), .E(n990), .CK(clk), .Q(R6[16]) );
  EDFFX1 R6_reg_15_ ( .D(data_in_1[15]), .E(n990), .CK(clk), .Q(R6[15]) );
  EDFFX1 R6_reg_14_ ( .D(data_in_1[14]), .E(n990), .CK(clk), .Q(R6[14]) );
  EDFFX1 R6_reg_13_ ( .D(data_in_1[13]), .E(n990), .CK(clk), .Q(R6[13]) );
  EDFFX1 R6_reg_12_ ( .D(data_in_1[12]), .E(n990), .CK(clk), .Q(R6[12]) );
  EDFFX1 R6_reg_11_ ( .D(data_in_1[11]), .E(n990), .CK(clk), .Q(R6[11]) );
  EDFFX1 R6_reg_10_ ( .D(data_in_1[10]), .E(n990), .CK(clk), .Q(R6[10]) );
  EDFFX1 R6_reg_9_ ( .D(data_in_1[9]), .E(n989), .CK(clk), .Q(R6[9]) );
  EDFFX1 R6_reg_8_ ( .D(data_in_1[8]), .E(n990), .CK(clk), .Q(R6[8]) );
  EDFFX1 R6_reg_7_ ( .D(data_in_1[7]), .E(n989), .CK(clk), .Q(R6[7]) );
  EDFFX1 R6_reg_6_ ( .D(data_in_1[6]), .E(n990), .CK(clk), .Q(R6[6]) );
  EDFFX1 R6_reg_5_ ( .D(data_in_1[5]), .E(n989), .CK(clk), .Q(R6[5]) );
  EDFFX1 R6_reg_4_ ( .D(data_in_1[4]), .E(n990), .CK(clk), .Q(R6[4]) );
  EDFFX1 R6_reg_3_ ( .D(data_in_1[3]), .E(n989), .CK(clk), .Q(R6[3]) );
  EDFFX1 R6_reg_2_ ( .D(data_in_1[2]), .E(n990), .CK(clk), .Q(R6[2]) );
  EDFFX1 R6_reg_1_ ( .D(data_in_1[1]), .E(n989), .CK(clk), .Q(R6[1]) );
  EDFFX1 R6_reg_0_ ( .D(data_in_1[0]), .E(n990), .CK(clk), .Q(R6[0]) );
  EDFFX1 R10_reg_33_ ( .D(data_in_1[33]), .E(n972), .CK(clk), .Q(R10[33]) );
  EDFFX1 R10_reg_32_ ( .D(data_in_1[32]), .E(n972), .CK(clk), .Q(R10[32]) );
  EDFFX1 R10_reg_31_ ( .D(data_in_1[31]), .E(n972), .CK(clk), .Q(R10[31]) );
  EDFFX1 R10_reg_30_ ( .D(data_in_1[30]), .E(n972), .CK(clk), .Q(R10[30]) );
  EDFFX1 R10_reg_29_ ( .D(data_in_1[29]), .E(n972), .CK(clk), .Q(R10[29]) );
  EDFFX1 R10_reg_28_ ( .D(data_in_1[28]), .E(n972), .CK(clk), .Q(R10[28]) );
  EDFFX1 R10_reg_27_ ( .D(data_in_1[27]), .E(n972), .CK(clk), .Q(R10[27]) );
  EDFFX1 R10_reg_26_ ( .D(data_in_1[26]), .E(n972), .CK(clk), .Q(R10[26]) );
  EDFFX1 R10_reg_25_ ( .D(data_in_1[25]), .E(n1000), .CK(clk), .Q(R10[25]) );
  EDFFX1 R10_reg_24_ ( .D(data_in_1[24]), .E(n999), .CK(clk), .Q(R10[24]) );
  EDFFX1 R10_reg_23_ ( .D(data_in_1[23]), .E(n1000), .CK(clk), .Q(R10[23]) );
  EDFFX1 R10_reg_22_ ( .D(data_in_1[22]), .E(n1000), .CK(clk), .Q(R10[22]) );
  EDFFX1 R10_reg_21_ ( .D(data_in_1[21]), .E(n999), .CK(clk), .Q(R10[21]) );
  EDFFX1 R10_reg_20_ ( .D(data_in_1[20]), .E(n999), .CK(clk), .Q(R10[20]) );
  EDFFX1 R10_reg_19_ ( .D(data_in_1[19]), .E(n999), .CK(clk), .Q(R10[19]) );
  EDFFX1 R10_reg_18_ ( .D(data_in_1[18]), .E(n999), .CK(clk), .Q(R10[18]) );
  EDFFX1 R10_reg_17_ ( .D(data_in_1[17]), .E(n999), .CK(clk), .Q(R10[17]) );
  EDFFX1 R10_reg_16_ ( .D(data_in_1[16]), .E(n999), .CK(clk), .Q(R10[16]) );
  EDFFX1 R10_reg_15_ ( .D(data_in_1[15]), .E(n999), .CK(clk), .Q(R10[15]) );
  EDFFX1 R10_reg_14_ ( .D(data_in_1[14]), .E(n999), .CK(clk), .Q(R10[14]) );
  EDFFX1 R10_reg_13_ ( .D(data_in_1[13]), .E(n999), .CK(clk), .Q(R10[13]) );
  EDFFX1 R10_reg_12_ ( .D(data_in_1[12]), .E(n999), .CK(clk), .Q(R10[12]) );
  EDFFX1 R10_reg_11_ ( .D(data_in_1[11]), .E(n999), .CK(clk), .Q(R10[11]) );
  EDFFX1 R10_reg_10_ ( .D(data_in_1[10]), .E(n999), .CK(clk), .Q(R10[10]) );
  EDFFX1 R10_reg_9_ ( .D(data_in_1[9]), .E(n1000), .CK(clk), .Q(R10[9]) );
  EDFFX1 R10_reg_8_ ( .D(data_in_1[8]), .E(n1000), .CK(clk), .Q(R10[8]) );
  EDFFX1 R10_reg_7_ ( .D(data_in_1[7]), .E(n1000), .CK(clk), .Q(R10[7]) );
  EDFFX1 R10_reg_6_ ( .D(data_in_1[6]), .E(n1000), .CK(clk), .Q(R10[6]) );
  EDFFX1 R10_reg_5_ ( .D(data_in_1[5]), .E(n1000), .CK(clk), .Q(R10[5]) );
  EDFFX1 R10_reg_4_ ( .D(data_in_1[4]), .E(n1000), .CK(clk), .Q(R10[4]) );
  EDFFX1 R10_reg_3_ ( .D(data_in_1[3]), .E(n1000), .CK(clk), .Q(R10[3]) );
  EDFFX1 R10_reg_2_ ( .D(data_in_1[2]), .E(n1000), .CK(clk), .Q(R10[2]) );
  EDFFX1 R10_reg_1_ ( .D(data_in_1[1]), .E(n1000), .CK(clk), .Q(R10[1]) );
  EDFFX1 R10_reg_0_ ( .D(data_in_1[0]), .E(n1000), .CK(clk), .Q(R10[0]) );
  EDFFX1 R0_reg_33_ ( .D(data_in_1[33]), .E(n1042), .CK(clk), .Q(R0[33]) );
  EDFFX1 R0_reg_32_ ( .D(data_in_1[32]), .E(n1042), .CK(clk), .Q(R0[32]) );
  EDFFX1 R0_reg_31_ ( .D(data_in_1[31]), .E(n1042), .CK(clk), .Q(R0[31]) );
  EDFFX1 R0_reg_30_ ( .D(data_in_1[30]), .E(n1042), .CK(clk), .Q(R0[30]) );
  EDFFX1 R0_reg_29_ ( .D(data_in_1[29]), .E(n1042), .CK(clk), .Q(R0[29]) );
  EDFFX1 R0_reg_28_ ( .D(data_in_1[28]), .E(n1042), .CK(clk), .Q(R0[28]) );
  EDFFX1 R0_reg_27_ ( .D(data_in_1[27]), .E(n1042), .CK(clk), .Q(R0[27]) );
  EDFFX1 R0_reg_26_ ( .D(data_in_1[26]), .E(n1042), .CK(clk), .Q(R0[26]) );
  EDFFX1 R0_reg_25_ ( .D(data_in_1[25]), .E(n1042), .CK(clk), .Q(R0[25]) );
  EDFFX1 R0_reg_24_ ( .D(data_in_1[24]), .E(n1042), .CK(clk), .Q(R0[24]) );
  EDFFX1 R0_reg_23_ ( .D(data_in_1[23]), .E(n1041), .CK(clk), .Q(R0[23]) );
  EDFFX1 R0_reg_22_ ( .D(data_in_1[22]), .E(n1040), .CK(clk), .Q(R0[22]) );
  EDFFX1 R0_reg_21_ ( .D(data_in_1[21]), .E(n1035), .CK(clk), .Q(R0[21]) );
  EDFFX1 R0_reg_20_ ( .D(data_in_1[20]), .E(n1034), .CK(clk), .Q(R0[20]) );
  EDFFX1 R0_reg_19_ ( .D(data_in_1[19]), .E(n1039), .CK(clk), .Q(R0[19]) );
  EDFFX1 R0_reg_18_ ( .D(data_in_1[18]), .E(n1037), .CK(clk), .Q(R0[18]) );
  EDFFX1 R0_reg_17_ ( .D(data_in_1[17]), .E(n1038), .CK(clk), .Q(R0[17]) );
  EDFFX1 R0_reg_16_ ( .D(data_in_1[16]), .E(n1036), .CK(clk), .Q(R0[16]) );
  EDFFX1 R0_reg_15_ ( .D(data_in_1[15]), .E(n1034), .CK(clk), .Q(R0[15]) );
  EDFFX1 R0_reg_14_ ( .D(data_in_1[14]), .E(n1041), .CK(clk), .Q(R0[14]) );
  EDFFX1 R0_reg_13_ ( .D(data_in_1[13]), .E(n1040), .CK(clk), .Q(R0[13]) );
  EDFFX1 R0_reg_12_ ( .D(data_in_1[12]), .E(n1035), .CK(clk), .Q(R0[12]) );
  EDFFX1 R0_reg_11_ ( .D(data_in_1[11]), .E(n1034), .CK(clk), .Q(R0[11]) );
  EDFFX1 R0_reg_10_ ( .D(data_in_1[10]), .E(n1039), .CK(clk), .Q(R0[10]) );
  EDFFX1 R0_reg_9_ ( .D(data_in_1[9]), .E(n1037), .CK(clk), .Q(R0[9]) );
  EDFFX1 R0_reg_8_ ( .D(data_in_1[8]), .E(n1038), .CK(clk), .Q(R0[8]) );
  EDFFX1 R0_reg_7_ ( .D(data_in_1[7]), .E(n1036), .CK(clk), .Q(R0[7]) );
  EDFFX1 R0_reg_6_ ( .D(data_in_1[6]), .E(n1040), .CK(clk), .Q(R0[6]) );
  EDFFX1 R0_reg_5_ ( .D(data_in_1[5]), .E(n1035), .CK(clk), .Q(R0[5]) );
  EDFFX1 R0_reg_4_ ( .D(data_in_1[4]), .E(n1034), .CK(clk), .Q(R0[4]) );
  EDFFX1 R0_reg_3_ ( .D(data_in_1[3]), .E(n1039), .CK(clk), .Q(R0[3]) );
  EDFFX1 R0_reg_2_ ( .D(data_in_1[2]), .E(n1037), .CK(clk), .Q(R0[2]) );
  EDFFX1 R0_reg_1_ ( .D(data_in_1[1]), .E(n1038), .CK(clk), .Q(R0[1]) );
  EDFFX1 R0_reg_0_ ( .D(data_in_1[0]), .E(n1036), .CK(clk), .Q(R0[0]) );
  EDFFX1 R4_reg_33_ ( .D(data_in_1[33]), .E(n985), .CK(clk), .Q(R4[33]) );
  EDFFX1 R4_reg_32_ ( .D(data_in_1[32]), .E(n985), .CK(clk), .Q(R4[32]) );
  EDFFX1 R4_reg_31_ ( .D(data_in_1[31]), .E(n985), .CK(clk), .Q(R4[31]) );
  EDFFX1 R4_reg_30_ ( .D(data_in_1[30]), .E(n985), .CK(clk), .Q(R4[30]) );
  EDFFX1 R4_reg_29_ ( .D(data_in_1[29]), .E(n985), .CK(clk), .Q(R4[29]) );
  EDFFX1 R4_reg_28_ ( .D(data_in_1[28]), .E(n985), .CK(clk), .Q(R4[28]) );
  EDFFX1 R4_reg_27_ ( .D(data_in_1[27]), .E(n985), .CK(clk), .Q(R4[27]) );
  EDFFX1 R4_reg_26_ ( .D(data_in_1[26]), .E(n985), .CK(clk), .Q(R4[26]) );
  EDFFX1 R4_reg_25_ ( .D(data_in_1[25]), .E(n985), .CK(clk), .Q(R4[25]) );
  EDFFX1 R4_reg_24_ ( .D(data_in_1[24]), .E(n985), .CK(clk), .Q(R4[24]) );
  EDFFX1 R4_reg_23_ ( .D(data_in_1[23]), .E(n985), .CK(clk), .Q(R4[23]) );
  EDFFX1 R4_reg_22_ ( .D(data_in_1[22]), .E(n985), .CK(clk), .Q(R4[22]) );
  EDFFX1 R4_reg_21_ ( .D(data_in_1[21]), .E(n986), .CK(clk), .Q(R4[21]) );
  EDFFX1 R4_reg_20_ ( .D(data_in_1[20]), .E(n986), .CK(clk), .Q(R4[20]) );
  EDFFX1 R4_reg_19_ ( .D(data_in_1[19]), .E(n986), .CK(clk), .Q(R4[19]) );
  EDFFX1 R4_reg_18_ ( .D(data_in_1[18]), .E(n986), .CK(clk), .Q(R4[18]) );
  EDFFX1 R4_reg_17_ ( .D(data_in_1[17]), .E(n986), .CK(clk), .Q(R4[17]) );
  EDFFX1 R4_reg_16_ ( .D(data_in_1[16]), .E(n986), .CK(clk), .Q(R4[16]) );
  EDFFX1 R4_reg_15_ ( .D(data_in_1[15]), .E(n986), .CK(clk), .Q(R4[15]) );
  EDFFX1 R4_reg_14_ ( .D(data_in_1[14]), .E(n986), .CK(clk), .Q(R4[14]) );
  EDFFX1 R4_reg_13_ ( .D(data_in_1[13]), .E(n986), .CK(clk), .Q(R4[13]) );
  EDFFX1 R4_reg_12_ ( .D(data_in_1[12]), .E(n986), .CK(clk), .Q(R4[12]) );
  EDFFX1 R4_reg_11_ ( .D(data_in_1[11]), .E(n986), .CK(clk), .Q(R4[11]) );
  EDFFX1 R4_reg_10_ ( .D(data_in_1[10]), .E(n986), .CK(clk), .Q(R4[10]) );
  EDFFX1 R4_reg_9_ ( .D(data_in_1[9]), .E(n985), .CK(clk), .Q(R4[9]) );
  EDFFX1 R4_reg_8_ ( .D(data_in_1[8]), .E(n986), .CK(clk), .Q(R4[8]) );
  EDFFX1 R4_reg_7_ ( .D(data_in_1[7]), .E(n985), .CK(clk), .Q(R4[7]) );
  EDFFX1 R4_reg_6_ ( .D(data_in_1[6]), .E(n986), .CK(clk), .Q(R4[6]) );
  EDFFX1 R4_reg_5_ ( .D(data_in_1[5]), .E(n985), .CK(clk), .Q(R4[5]) );
  EDFFX1 R4_reg_4_ ( .D(data_in_1[4]), .E(n986), .CK(clk), .Q(R4[4]) );
  EDFFX1 R4_reg_3_ ( .D(data_in_1[3]), .E(n985), .CK(clk), .Q(R4[3]) );
  EDFFX1 R4_reg_2_ ( .D(data_in_1[2]), .E(n986), .CK(clk), .Q(R4[2]) );
  EDFFX1 R4_reg_1_ ( .D(data_in_1[1]), .E(n985), .CK(clk), .Q(R4[1]) );
  EDFFX1 R4_reg_0_ ( .D(data_in_1[0]), .E(n986), .CK(clk), .Q(R4[0]) );
  EDFFX1 R8_reg_33_ ( .D(data_in_1[33]), .E(n974), .CK(clk), .Q(R8[33]) );
  EDFFX1 R8_reg_32_ ( .D(data_in_1[32]), .E(n974), .CK(clk), .Q(R8[32]) );
  EDFFX1 R8_reg_31_ ( .D(data_in_1[31]), .E(n974), .CK(clk), .Q(R8[31]) );
  EDFFX1 R8_reg_30_ ( .D(data_in_1[30]), .E(n974), .CK(clk), .Q(R8[30]) );
  EDFFX1 R8_reg_29_ ( .D(data_in_1[29]), .E(n974), .CK(clk), .Q(R8[29]) );
  EDFFX1 R8_reg_28_ ( .D(data_in_1[28]), .E(n974), .CK(clk), .Q(R8[28]) );
  EDFFX1 R8_reg_27_ ( .D(data_in_1[27]), .E(n974), .CK(clk), .Q(R8[27]) );
  EDFFX1 R8_reg_26_ ( .D(data_in_1[26]), .E(n974), .CK(clk), .Q(R8[26]) );
  EDFFX1 R8_reg_25_ ( .D(data_in_1[25]), .E(n994), .CK(clk), .Q(R8[25]) );
  EDFFX1 R8_reg_24_ ( .D(data_in_1[24]), .E(n993), .CK(clk), .Q(R8[24]) );
  EDFFX1 R8_reg_23_ ( .D(data_in_1[23]), .E(n994), .CK(clk), .Q(R8[23]) );
  EDFFX1 R8_reg_22_ ( .D(data_in_1[22]), .E(n994), .CK(clk), .Q(R8[22]) );
  EDFFX1 R8_reg_21_ ( .D(data_in_1[21]), .E(n993), .CK(clk), .Q(R8[21]) );
  EDFFX1 R8_reg_20_ ( .D(data_in_1[20]), .E(n993), .CK(clk), .Q(R8[20]) );
  EDFFX1 R8_reg_19_ ( .D(data_in_1[19]), .E(n993), .CK(clk), .Q(R8[19]) );
  EDFFX1 R8_reg_18_ ( .D(data_in_1[18]), .E(n993), .CK(clk), .Q(R8[18]) );
  EDFFX1 R8_reg_17_ ( .D(data_in_1[17]), .E(n993), .CK(clk), .Q(R8[17]) );
  EDFFX1 R8_reg_16_ ( .D(data_in_1[16]), .E(n993), .CK(clk), .Q(R8[16]) );
  EDFFX1 R8_reg_15_ ( .D(data_in_1[15]), .E(n993), .CK(clk), .Q(R8[15]) );
  EDFFX1 R8_reg_14_ ( .D(data_in_1[14]), .E(n993), .CK(clk), .Q(R8[14]) );
  EDFFX1 R8_reg_13_ ( .D(data_in_1[13]), .E(n993), .CK(clk), .Q(R8[13]) );
  EDFFX1 R8_reg_12_ ( .D(data_in_1[12]), .E(n993), .CK(clk), .Q(R8[12]) );
  EDFFX1 R8_reg_11_ ( .D(data_in_1[11]), .E(n993), .CK(clk), .Q(R8[11]) );
  EDFFX1 R8_reg_10_ ( .D(data_in_1[10]), .E(n993), .CK(clk), .Q(R8[10]) );
  EDFFX1 R8_reg_9_ ( .D(data_in_1[9]), .E(n994), .CK(clk), .Q(R8[9]) );
  EDFFX1 R8_reg_8_ ( .D(data_in_1[8]), .E(n994), .CK(clk), .Q(R8[8]) );
  EDFFX1 R8_reg_7_ ( .D(data_in_1[7]), .E(n994), .CK(clk), .Q(R8[7]) );
  EDFFX1 R8_reg_6_ ( .D(data_in_1[6]), .E(n994), .CK(clk), .Q(R8[6]) );
  EDFFX1 R8_reg_5_ ( .D(data_in_1[5]), .E(n994), .CK(clk), .Q(R8[5]) );
  EDFFX1 R8_reg_4_ ( .D(data_in_1[4]), .E(n994), .CK(clk), .Q(R8[4]) );
  EDFFX1 R8_reg_3_ ( .D(data_in_1[3]), .E(n994), .CK(clk), .Q(R8[3]) );
  EDFFX1 R8_reg_2_ ( .D(data_in_1[2]), .E(n994), .CK(clk), .Q(R8[2]) );
  EDFFX1 R8_reg_1_ ( .D(data_in_1[1]), .E(n994), .CK(clk), .Q(R8[1]) );
  EDFFX1 R8_reg_0_ ( .D(data_in_1[0]), .E(n994), .CK(clk), .Q(R8[0]) );
  EDFFX1 R12_reg_33_ ( .D(data_in_1[33]), .E(n1006), .CK(clk), .Q(R12[33]) );
  EDFFX1 R12_reg_32_ ( .D(data_in_1[32]), .E(n1006), .CK(clk), .Q(R12[32]) );
  EDFFX1 R12_reg_31_ ( .D(data_in_1[31]), .E(n1006), .CK(clk), .Q(R12[31]) );
  EDFFX1 R12_reg_30_ ( .D(data_in_1[30]), .E(n1006), .CK(clk), .Q(R12[30]) );
  EDFFX1 R12_reg_29_ ( .D(data_in_1[29]), .E(n1006), .CK(clk), .Q(R12[29]) );
  EDFFX1 R12_reg_28_ ( .D(data_in_1[28]), .E(n1006), .CK(clk), .Q(R12[28]) );
  EDFFX1 R12_reg_27_ ( .D(data_in_1[27]), .E(n1006), .CK(clk), .Q(R12[27]) );
  EDFFX1 R12_reg_26_ ( .D(data_in_1[26]), .E(n1006), .CK(clk), .Q(R12[26]) );
  EDFFX1 R12_reg_25_ ( .D(data_in_1[25]), .E(n1006), .CK(clk), .Q(R12[25]) );
  EDFFX1 R12_reg_24_ ( .D(data_in_1[24]), .E(n1006), .CK(clk), .Q(R12[24]) );
  EDFFX1 R12_reg_23_ ( .D(data_in_1[23]), .E(n1005), .CK(clk), .Q(R12[23]) );
  EDFFX1 R12_reg_22_ ( .D(data_in_1[22]), .E(n1005), .CK(clk), .Q(R12[22]) );
  EDFFX1 R12_reg_21_ ( .D(data_in_1[21]), .E(n1005), .CK(clk), .Q(R12[21]) );
  EDFFX1 R12_reg_20_ ( .D(data_in_1[20]), .E(n1005), .CK(clk), .Q(R12[20]) );
  EDFFX1 R12_reg_19_ ( .D(data_in_1[19]), .E(n1005), .CK(clk), .Q(R12[19]) );
  EDFFX1 R12_reg_18_ ( .D(data_in_1[18]), .E(n1005), .CK(clk), .Q(R12[18]) );
  EDFFX1 R12_reg_17_ ( .D(data_in_1[17]), .E(n1005), .CK(clk), .Q(R12[17]) );
  EDFFX1 R12_reg_16_ ( .D(data_in_1[16]), .E(n1005), .CK(clk), .Q(R12[16]) );
  EDFFX1 R12_reg_15_ ( .D(data_in_1[15]), .E(n1005), .CK(clk), .Q(R12[15]) );
  EDFFX1 R12_reg_14_ ( .D(data_in_1[14]), .E(n1005), .CK(clk), .Q(R12[14]) );
  EDFFX1 R12_reg_13_ ( .D(data_in_1[13]), .E(n1005), .CK(clk), .Q(R12[13]) );
  EDFFX1 R12_reg_12_ ( .D(data_in_1[12]), .E(n1005), .CK(clk), .Q(R12[12]) );
  EDFFX1 R12_reg_11_ ( .D(data_in_1[11]), .E(n970), .CK(clk), .Q(R12[11]) );
  EDFFX1 R12_reg_10_ ( .D(data_in_1[10]), .E(n970), .CK(clk), .Q(R12[10]) );
  EDFFX1 R12_reg_9_ ( .D(data_in_1[9]), .E(n970), .CK(clk), .Q(R12[9]) );
  EDFFX1 R12_reg_8_ ( .D(data_in_1[8]), .E(n970), .CK(clk), .Q(R12[8]) );
  EDFFX1 R12_reg_7_ ( .D(data_in_1[7]), .E(n970), .CK(clk), .Q(R12[7]) );
  EDFFX1 R12_reg_6_ ( .D(data_in_1[6]), .E(n970), .CK(clk), .Q(R12[6]) );
  EDFFX1 R12_reg_5_ ( .D(data_in_1[5]), .E(n970), .CK(clk), .Q(R12[5]) );
  EDFFX1 R12_reg_4_ ( .D(data_in_1[4]), .E(n1005), .CK(clk), .Q(R12[4]) );
  EDFFX1 R12_reg_3_ ( .D(data_in_1[3]), .E(n1006), .CK(clk), .Q(R12[3]) );
  EDFFX1 R12_reg_2_ ( .D(data_in_1[2]), .E(n1005), .CK(clk), .Q(R12[2]) );
  EDFFX1 R12_reg_1_ ( .D(data_in_1[1]), .E(n1006), .CK(clk), .Q(R12[1]) );
  EDFFX1 R12_reg_0_ ( .D(data_in_1[0]), .E(n1006), .CK(clk), .Q(R12[0]) );
  EDFFX1 R15_reg_33_ ( .D(data_in_1[33]), .E(n1031), .CK(clk), .Q(R15[33]) );
  EDFFX1 R15_reg_32_ ( .D(data_in_1[32]), .E(n1031), .CK(clk), .Q(R15[32]) );
  EDFFX1 R15_reg_31_ ( .D(data_in_1[31]), .E(n1031), .CK(clk), .Q(R15[31]) );
  EDFFX1 R15_reg_30_ ( .D(data_in_1[30]), .E(n1031), .CK(clk), .Q(R15[30]) );
  EDFFX1 R15_reg_29_ ( .D(data_in_1[29]), .E(n1031), .CK(clk), .Q(R15[29]) );
  EDFFX1 R15_reg_28_ ( .D(data_in_1[28]), .E(n1031), .CK(clk), .Q(R15[28]) );
  EDFFX1 R15_reg_27_ ( .D(data_in_1[27]), .E(n1031), .CK(clk), .Q(R15[27]) );
  EDFFX1 R15_reg_26_ ( .D(data_in_1[26]), .E(n1031), .CK(clk), .Q(R15[26]) );
  EDFFX1 R15_reg_25_ ( .D(data_in_1[25]), .E(n1031), .CK(clk), .Q(R15[25]) );
  EDFFX1 R15_reg_24_ ( .D(data_in_1[24]), .E(n1031), .CK(clk), .Q(R15[24]) );
  EDFFX1 R15_reg_23_ ( .D(data_in_1[23]), .E(n1031), .CK(clk), .Q(R15[23]) );
  EDFFX1 R15_reg_22_ ( .D(data_in_1[22]), .E(n1031), .CK(clk), .Q(R15[22]) );
  EDFFX1 R15_reg_21_ ( .D(data_in_1[21]), .E(n1031), .CK(clk), .Q(R15[21]) );
  EDFFX1 R15_reg_20_ ( .D(data_in_1[20]), .E(n1031), .CK(clk), .Q(R15[20]) );
  EDFFX1 R15_reg_19_ ( .D(data_in_1[19]), .E(n1031), .CK(clk), .Q(R15[19]) );
  EDFFX1 R15_reg_18_ ( .D(data_in_1[18]), .E(n1031), .CK(clk), .Q(R15[18]) );
  EDFFX1 R15_reg_17_ ( .D(data_in_1[17]), .E(n1031), .CK(clk), .Q(R15[17]) );
  EDFFX1 R15_reg_16_ ( .D(data_in_1[16]), .E(n1031), .CK(clk), .Q(R15[16]) );
  EDFFX1 R15_reg_15_ ( .D(data_in_1[15]), .E(n1031), .CK(clk), .Q(R15[15]) );
  EDFFX1 R15_reg_14_ ( .D(data_in_1[14]), .E(n1031), .CK(clk), .Q(R15[14]) );
  EDFFX1 R15_reg_13_ ( .D(data_in_1[13]), .E(n1031), .CK(clk), .Q(R15[13]) );
  EDFFX1 R15_reg_12_ ( .D(data_in_1[12]), .E(n1031), .CK(clk), .Q(R15[12]) );
  EDFFX1 R15_reg_11_ ( .D(data_in_1[11]), .E(n1031), .CK(clk), .Q(R15[11]) );
  EDFFX1 R15_reg_10_ ( .D(data_in_1[10]), .E(n1031), .CK(clk), .Q(R15[10]) );
  EDFFX1 R15_reg_9_ ( .D(data_in_1[9]), .E(n1031), .CK(clk), .Q(R15[9]) );
  EDFFX1 R15_reg_8_ ( .D(data_in_1[8]), .E(n1031), .CK(clk), .Q(R15[8]) );
  EDFFX1 R15_reg_7_ ( .D(data_in_1[7]), .E(n1031), .CK(clk), .Q(R15[7]) );
  EDFFX1 R15_reg_6_ ( .D(data_in_1[6]), .E(n1031), .CK(clk), .Q(R15[6]) );
  EDFFX1 R15_reg_5_ ( .D(data_in_1[5]), .E(n1031), .CK(clk), .Q(R15[5]) );
  EDFFX1 R15_reg_4_ ( .D(data_in_1[4]), .E(n1031), .CK(clk), .Q(R15[4]) );
  EDFFX1 R15_reg_3_ ( .D(data_in_1[3]), .E(n1031), .CK(clk), .Q(R15[3]) );
  EDFFX1 R15_reg_2_ ( .D(data_in_1[2]), .E(n1031), .CK(clk), .Q(R15[2]) );
  EDFFX1 R15_reg_1_ ( .D(data_in_1[1]), .E(n1031), .CK(clk), .Q(R15[1]) );
  EDFFX1 R15_reg_0_ ( .D(data_in_1[0]), .E(n1031), .CK(clk), .Q(R15[0]) );
  EDFFX1 R3_reg_33_ ( .D(data_in_1[33]), .E(n983), .CK(clk), .Q(R3[33]) );
  EDFFX1 R3_reg_32_ ( .D(data_in_1[32]), .E(n983), .CK(clk), .Q(R3[32]) );
  EDFFX1 R3_reg_31_ ( .D(data_in_1[31]), .E(n983), .CK(clk), .Q(R3[31]) );
  EDFFX1 R3_reg_30_ ( .D(data_in_1[30]), .E(n983), .CK(clk), .Q(R3[30]) );
  EDFFX1 R3_reg_29_ ( .D(data_in_1[29]), .E(n983), .CK(clk), .Q(R3[29]) );
  EDFFX1 R3_reg_28_ ( .D(data_in_1[28]), .E(n983), .CK(clk), .Q(R3[28]) );
  EDFFX1 R3_reg_27_ ( .D(data_in_1[27]), .E(n983), .CK(clk), .Q(R3[27]) );
  EDFFX1 R3_reg_26_ ( .D(data_in_1[26]), .E(n983), .CK(clk), .Q(R3[26]) );
  EDFFX1 R3_reg_25_ ( .D(data_in_1[25]), .E(n983), .CK(clk), .Q(R3[25]) );
  EDFFX1 R3_reg_24_ ( .D(data_in_1[24]), .E(n983), .CK(clk), .Q(R3[24]) );
  EDFFX1 R3_reg_23_ ( .D(data_in_1[23]), .E(n983), .CK(clk), .Q(R3[23]) );
  EDFFX1 R3_reg_22_ ( .D(data_in_1[22]), .E(n983), .CK(clk), .Q(R3[22]) );
  EDFFX1 R3_reg_21_ ( .D(data_in_1[21]), .E(n984), .CK(clk), .Q(R3[21]) );
  EDFFX1 R3_reg_20_ ( .D(data_in_1[20]), .E(n984), .CK(clk), .Q(R3[20]) );
  EDFFX1 R3_reg_19_ ( .D(data_in_1[19]), .E(n984), .CK(clk), .Q(R3[19]) );
  EDFFX1 R3_reg_18_ ( .D(data_in_1[18]), .E(n984), .CK(clk), .Q(R3[18]) );
  EDFFX1 R3_reg_17_ ( .D(data_in_1[17]), .E(n984), .CK(clk), .Q(R3[17]) );
  EDFFX1 R3_reg_16_ ( .D(data_in_1[16]), .E(n984), .CK(clk), .Q(R3[16]) );
  EDFFX1 R3_reg_15_ ( .D(data_in_1[15]), .E(n984), .CK(clk), .Q(R3[15]) );
  EDFFX1 R3_reg_14_ ( .D(data_in_1[14]), .E(n984), .CK(clk), .Q(R3[14]) );
  EDFFX1 R3_reg_13_ ( .D(data_in_1[13]), .E(n984), .CK(clk), .Q(R3[13]) );
  EDFFX1 R3_reg_12_ ( .D(data_in_1[12]), .E(n984), .CK(clk), .Q(R3[12]) );
  EDFFX1 R3_reg_11_ ( .D(data_in_1[11]), .E(n984), .CK(clk), .Q(R3[11]) );
  EDFFX1 R3_reg_10_ ( .D(data_in_1[10]), .E(n984), .CK(clk), .Q(R3[10]) );
  EDFFX1 R3_reg_9_ ( .D(data_in_1[9]), .E(n983), .CK(clk), .Q(R3[9]) );
  EDFFX1 R3_reg_8_ ( .D(data_in_1[8]), .E(n984), .CK(clk), .Q(R3[8]) );
  EDFFX1 R3_reg_7_ ( .D(data_in_1[7]), .E(n983), .CK(clk), .Q(R3[7]) );
  EDFFX1 R3_reg_6_ ( .D(data_in_1[6]), .E(n984), .CK(clk), .Q(R3[6]) );
  EDFFX1 R3_reg_5_ ( .D(data_in_1[5]), .E(n983), .CK(clk), .Q(R3[5]) );
  EDFFX1 R3_reg_4_ ( .D(data_in_1[4]), .E(n984), .CK(clk), .Q(R3[4]) );
  EDFFX1 R3_reg_3_ ( .D(data_in_1[3]), .E(n983), .CK(clk), .Q(R3[3]) );
  EDFFX1 R3_reg_2_ ( .D(data_in_1[2]), .E(n984), .CK(clk), .Q(R3[2]) );
  EDFFX1 R3_reg_1_ ( .D(data_in_1[1]), .E(n983), .CK(clk), .Q(R3[1]) );
  EDFFX1 R3_reg_0_ ( .D(data_in_1[0]), .E(n984), .CK(clk), .Q(R3[0]) );
  EDFFX1 R7_reg_33_ ( .D(data_in_1[33]), .E(n991), .CK(clk), .Q(R7[33]) );
  EDFFX1 R7_reg_32_ ( .D(data_in_1[32]), .E(n992), .CK(clk), .Q(R7[32]) );
  EDFFX1 R7_reg_31_ ( .D(data_in_1[31]), .E(n991), .CK(clk), .Q(R7[31]) );
  EDFFX1 R7_reg_30_ ( .D(data_in_1[30]), .E(n992), .CK(clk), .Q(R7[30]) );
  EDFFX1 R7_reg_29_ ( .D(data_in_1[29]), .E(n991), .CK(clk), .Q(R7[29]) );
  EDFFX1 R7_reg_28_ ( .D(data_in_1[28]), .E(n992), .CK(clk), .Q(R7[28]) );
  EDFFX1 R7_reg_27_ ( .D(data_in_1[27]), .E(n991), .CK(clk), .Q(R7[27]) );
  EDFFX1 R7_reg_26_ ( .D(data_in_1[26]), .E(n992), .CK(clk), .Q(R7[26]) );
  EDFFX1 R7_reg_25_ ( .D(data_in_1[25]), .E(n991), .CK(clk), .Q(R7[25]) );
  EDFFX1 R7_reg_24_ ( .D(data_in_1[24]), .E(n992), .CK(clk), .Q(R7[24]) );
  EDFFX1 R7_reg_23_ ( .D(data_in_1[23]), .E(n992), .CK(clk), .Q(R7[23]) );
  EDFFX1 R7_reg_22_ ( .D(data_in_1[22]), .E(n992), .CK(clk), .Q(R7[22]) );
  EDFFX1 R7_reg_21_ ( .D(data_in_1[21]), .E(n992), .CK(clk), .Q(R7[21]) );
  EDFFX1 R7_reg_20_ ( .D(data_in_1[20]), .E(n992), .CK(clk), .Q(R7[20]) );
  EDFFX1 R7_reg_19_ ( .D(data_in_1[19]), .E(n992), .CK(clk), .Q(R7[19]) );
  EDFFX1 R7_reg_18_ ( .D(data_in_1[18]), .E(n992), .CK(clk), .Q(R7[18]) );
  EDFFX1 R7_reg_17_ ( .D(data_in_1[17]), .E(n992), .CK(clk), .Q(R7[17]) );
  EDFFX1 R7_reg_16_ ( .D(data_in_1[16]), .E(n992), .CK(clk), .Q(R7[16]) );
  EDFFX1 R7_reg_15_ ( .D(data_in_1[15]), .E(n992), .CK(clk), .Q(R7[15]) );
  EDFFX1 R7_reg_14_ ( .D(data_in_1[14]), .E(n992), .CK(clk), .Q(R7[14]) );
  EDFFX1 R7_reg_13_ ( .D(data_in_1[13]), .E(n992), .CK(clk), .Q(R7[13]) );
  EDFFX1 R7_reg_12_ ( .D(data_in_1[12]), .E(n992), .CK(clk), .Q(R7[12]) );
  EDFFX1 R7_reg_11_ ( .D(data_in_1[11]), .E(n991), .CK(clk), .Q(R7[11]) );
  EDFFX1 R7_reg_10_ ( .D(data_in_1[10]), .E(n991), .CK(clk), .Q(R7[10]) );
  EDFFX1 R7_reg_9_ ( .D(data_in_1[9]), .E(n991), .CK(clk), .Q(R7[9]) );
  EDFFX1 R7_reg_8_ ( .D(data_in_1[8]), .E(n991), .CK(clk), .Q(R7[8]) );
  EDFFX1 R7_reg_7_ ( .D(data_in_1[7]), .E(n991), .CK(clk), .Q(R7[7]) );
  EDFFX1 R7_reg_6_ ( .D(data_in_1[6]), .E(n991), .CK(clk), .Q(R7[6]) );
  EDFFX1 R7_reg_5_ ( .D(data_in_1[5]), .E(n991), .CK(clk), .Q(R7[5]) );
  EDFFX1 R7_reg_4_ ( .D(data_in_1[4]), .E(n991), .CK(clk), .Q(R7[4]) );
  EDFFX1 R7_reg_3_ ( .D(data_in_1[3]), .E(n991), .CK(clk), .Q(R7[3]) );
  EDFFX1 R7_reg_2_ ( .D(data_in_1[2]), .E(n991), .CK(clk), .Q(R7[2]) );
  EDFFX1 R7_reg_1_ ( .D(data_in_1[1]), .E(n991), .CK(clk), .Q(R7[1]) );
  EDFFX1 R7_reg_0_ ( .D(data_in_1[0]), .E(n991), .CK(clk), .Q(R7[0]) );
  EDFFX1 R11_reg_33_ ( .D(data_in_1[33]), .E(n971), .CK(clk), .Q(R11[33]) );
  EDFFX1 R11_reg_32_ ( .D(data_in_1[32]), .E(n971), .CK(clk), .Q(R11[32]) );
  EDFFX1 R11_reg_31_ ( .D(data_in_1[31]), .E(n971), .CK(clk), .Q(R11[31]) );
  EDFFX1 R11_reg_30_ ( .D(data_in_1[30]), .E(n971), .CK(clk), .Q(R11[30]) );
  EDFFX1 R11_reg_29_ ( .D(data_in_1[29]), .E(n971), .CK(clk), .Q(R11[29]) );
  EDFFX1 R11_reg_28_ ( .D(data_in_1[28]), .E(n971), .CK(clk), .Q(R11[28]) );
  EDFFX1 R11_reg_27_ ( .D(data_in_1[27]), .E(n971), .CK(clk), .Q(R11[27]) );
  EDFFX1 R11_reg_26_ ( .D(data_in_1[26]), .E(n971), .CK(clk), .Q(R11[26]) );
  EDFFX1 R11_reg_25_ ( .D(data_in_1[25]), .E(n1003), .CK(clk), .Q(R11[25]) );
  EDFFX1 R11_reg_24_ ( .D(data_in_1[24]), .E(n1002), .CK(clk), .Q(R11[24]) );
  EDFFX1 R11_reg_23_ ( .D(data_in_1[23]), .E(n1003), .CK(clk), .Q(R11[23]) );
  EDFFX1 R11_reg_22_ ( .D(data_in_1[22]), .E(n1003), .CK(clk), .Q(R11[22]) );
  EDFFX1 R11_reg_21_ ( .D(data_in_1[21]), .E(n1002), .CK(clk), .Q(R11[21]) );
  EDFFX1 R11_reg_20_ ( .D(data_in_1[20]), .E(n1002), .CK(clk), .Q(R11[20]) );
  EDFFX1 R11_reg_19_ ( .D(data_in_1[19]), .E(n1002), .CK(clk), .Q(R11[19]) );
  EDFFX1 R11_reg_18_ ( .D(data_in_1[18]), .E(n1002), .CK(clk), .Q(R11[18]) );
  EDFFX1 R11_reg_17_ ( .D(data_in_1[17]), .E(n1002), .CK(clk), .Q(R11[17]) );
  EDFFX1 R11_reg_16_ ( .D(data_in_1[16]), .E(n1002), .CK(clk), .Q(R11[16]) );
  EDFFX1 R11_reg_15_ ( .D(data_in_1[15]), .E(n1002), .CK(clk), .Q(R11[15]) );
  EDFFX1 R11_reg_14_ ( .D(data_in_1[14]), .E(n1002), .CK(clk), .Q(R11[14]) );
  EDFFX1 R11_reg_13_ ( .D(data_in_1[13]), .E(n1002), .CK(clk), .Q(R11[13]) );
  EDFFX1 R11_reg_12_ ( .D(data_in_1[12]), .E(n1002), .CK(clk), .Q(R11[12]) );
  EDFFX1 R11_reg_11_ ( .D(data_in_1[11]), .E(n1002), .CK(clk), .Q(R11[11]) );
  EDFFX1 R11_reg_10_ ( .D(data_in_1[10]), .E(n1002), .CK(clk), .Q(R11[10]) );
  EDFFX1 R11_reg_9_ ( .D(data_in_1[9]), .E(n1003), .CK(clk), .Q(R11[9]) );
  EDFFX1 R11_reg_8_ ( .D(data_in_1[8]), .E(n1003), .CK(clk), .Q(R11[8]) );
  EDFFX1 R11_reg_7_ ( .D(data_in_1[7]), .E(n1003), .CK(clk), .Q(R11[7]) );
  EDFFX1 R11_reg_6_ ( .D(data_in_1[6]), .E(n1003), .CK(clk), .Q(R11[6]) );
  EDFFX1 R11_reg_5_ ( .D(data_in_1[5]), .E(n1003), .CK(clk), .Q(R11[5]) );
  EDFFX1 R11_reg_4_ ( .D(data_in_1[4]), .E(n1003), .CK(clk), .Q(R11[4]) );
  EDFFX1 R11_reg_3_ ( .D(data_in_1[3]), .E(n1003), .CK(clk), .Q(R11[3]) );
  EDFFX1 R11_reg_2_ ( .D(data_in_1[2]), .E(n1003), .CK(clk), .Q(R11[2]) );
  EDFFX1 R11_reg_1_ ( .D(data_in_1[1]), .E(n1003), .CK(clk), .Q(R11[1]) );
  EDFFX1 R11_reg_0_ ( .D(data_in_1[0]), .E(n1003), .CK(clk), .Q(R11[0]) );
  DFFRHQX1 s_p_flag_out_reg ( .D(n1006), .CK(clk), .RN(rst_n), .Q(s_p_flag_out) );
  DFFHQX1 data_out_1_reg_33_ ( .D(n934), .CK(clk), .Q(data_out_1[33]) );
  DFFHQX1 data_out_1_reg_16_ ( .D(n951), .CK(clk), .Q(data_out_1[16]) );
  JKFFRXL counter_reg_0_ ( .J(1'b1), .K(1'b1), .CK(clk), .RN(rst_n), .Q(
        counter[0]), .QN(n550) );
  DFFHQX1 data_out_1_reg_32_ ( .D(n935), .CK(clk), .Q(data_out_1[32]) );
  DFFHQX1 data_out_1_reg_31_ ( .D(n936), .CK(clk), .Q(data_out_1[31]) );
  DFFHQX1 data_out_1_reg_30_ ( .D(n937), .CK(clk), .Q(data_out_1[30]) );
  DFFHQX1 data_out_1_reg_28_ ( .D(n939), .CK(clk), .Q(data_out_1[28]) );
  DFFHQX1 data_out_1_reg_15_ ( .D(n952), .CK(clk), .Q(data_out_1[15]) );
  DFFHQX1 data_out_1_reg_14_ ( .D(n953), .CK(clk), .Q(data_out_1[14]) );
  DFFHQX1 data_out_1_reg_13_ ( .D(n954), .CK(clk), .Q(data_out_1[13]) );
  DFFHQX1 data_out_1_reg_11_ ( .D(n956), .CK(clk), .Q(data_out_1[11]) );
  DFFRHQX1 counter_reg_3_ ( .D(N15), .CK(clk), .RN(rst_n), .Q(counter[3]) );
  DFFRHQX1 counter_reg_1_ ( .D(N13), .CK(clk), .RN(rst_n), .Q(counter[1]) );
  DFFRHQX1 counter_reg_2_ ( .D(N14), .CK(clk), .RN(rst_n), .Q(counter[2]) );
  DFFHQX1 data_out_1_reg_27_ ( .D(n940), .CK(clk), .Q(data_out_1[27]) );
  DFFHQX1 data_out_1_reg_26_ ( .D(n941), .CK(clk), .Q(data_out_1[26]) );
  DFFHQX1 data_out_1_reg_25_ ( .D(n942), .CK(clk), .Q(data_out_1[25]) );
  DFFHQX1 data_out_1_reg_10_ ( .D(n957), .CK(clk), .Q(data_out_1[10]) );
  DFFHQX1 data_out_1_reg_9_ ( .D(n958), .CK(clk), .Q(data_out_1[9]) );
  DFFHQX1 data_out_1_reg_8_ ( .D(n959), .CK(clk), .Q(data_out_1[8]) );
  DFFHQX1 data_out_1_reg_29_ ( .D(n938), .CK(clk), .Q(data_out_1[29]) );
  DFFHQX1 data_out_1_reg_12_ ( .D(n955), .CK(clk), .Q(data_out_1[12]) );
  DFFHQX1 data_out_1_reg_24_ ( .D(n943), .CK(clk), .Q(data_out_1[24]) );
  DFFHQX1 data_out_1_reg_23_ ( .D(n944), .CK(clk), .Q(data_out_1[23]) );
  DFFHQX1 data_out_1_reg_22_ ( .D(n945), .CK(clk), .Q(data_out_1[22]) );
  DFFHQX1 data_out_1_reg_21_ ( .D(n946), .CK(clk), .Q(data_out_1[21]) );
  DFFHQX1 data_out_1_reg_20_ ( .D(n947), .CK(clk), .Q(data_out_1[20]) );
  DFFHQX1 data_out_1_reg_19_ ( .D(n948), .CK(clk), .Q(data_out_1[19]) );
  DFFHQX1 data_out_1_reg_18_ ( .D(n949), .CK(clk), .Q(data_out_1[18]) );
  DFFHQX1 data_out_1_reg_17_ ( .D(n950), .CK(clk), .Q(data_out_1[17]) );
  DFFHQX1 data_out_1_reg_7_ ( .D(n960), .CK(clk), .Q(data_out_1[7]) );
  DFFHQX1 data_out_1_reg_6_ ( .D(n961), .CK(clk), .Q(data_out_1[6]) );
  DFFHQX1 data_out_1_reg_5_ ( .D(n962), .CK(clk), .Q(data_out_1[5]) );
  DFFHQX1 data_out_1_reg_4_ ( .D(n963), .CK(clk), .Q(data_out_1[4]) );
  DFFHQX1 data_out_1_reg_3_ ( .D(n964), .CK(clk), .Q(data_out_1[3]) );
  DFFHQX1 data_out_1_reg_2_ ( .D(n965), .CK(clk), .Q(data_out_1[2]) );
  DFFHQX1 data_out_1_reg_0_ ( .D(n967), .CK(clk), .Q(data_out_1[0]) );
  DFFHQX1 data_out_1_reg_1_ ( .D(n966), .CK(clk), .Q(data_out_1[1]) );
  DFFHQX1 data_out_1_reg_49_ ( .D(n918), .CK(clk), .Q(data_out_1[49]) );
  DFFHQX1 data_out_1_reg_48_ ( .D(n919), .CK(clk), .Q(data_out_1[48]) );
  DFFHQX1 data_out_1_reg_100_ ( .D(n867), .CK(clk), .Q(data_out_1[100]) );
  DFFHQX1 data_out_1_reg_99_ ( .D(n868), .CK(clk), .Q(data_out_1[99]) );
  DFFHQX1 data_out_1_reg_83_ ( .D(n884), .CK(clk), .Q(data_out_1[83]) );
  DFFHQX1 data_out_1_reg_82_ ( .D(n885), .CK(clk), .Q(data_out_1[82]) );
  DFFHQX1 data_out_1_reg_134_ ( .D(n833), .CK(clk), .Q(data_out_1[134]) );
  DFFHQX1 data_out_1_reg_133_ ( .D(n834), .CK(clk), .Q(data_out_1[133]) );
  DFFHQX1 data_out_1_reg_117_ ( .D(n850), .CK(clk), .Q(data_out_1[117]) );
  DFFHQX1 data_out_1_reg_116_ ( .D(n851), .CK(clk), .Q(data_out_1[116]) );
  DFFHQX1 data_out_1_reg_81_ ( .D(n886), .CK(clk), .Q(data_out_1[81]) );
  DFFHQX1 data_out_1_reg_80_ ( .D(n887), .CK(clk), .Q(data_out_1[80]) );
  DFFHQX1 data_out_1_reg_79_ ( .D(n888), .CK(clk), .Q(data_out_1[79]) );
  DFFHQX1 data_out_1_reg_97_ ( .D(n870), .CK(clk), .Q(data_out_1[97]) );
  DFFHQX1 data_out_1_reg_98_ ( .D(n869), .CK(clk), .Q(data_out_1[98]) );
  DFFHQX1 data_out_1_reg_115_ ( .D(n852), .CK(clk), .Q(data_out_1[115]) );
  DFFHQX1 data_out_1_reg_46_ ( .D(n921), .CK(clk), .Q(data_out_1[46]) );
  DFFHQX1 data_out_1_reg_78_ ( .D(n889), .CK(clk), .Q(data_out_1[78]) );
  DFFHQX1 data_out_1_reg_77_ ( .D(n890), .CK(clk), .Q(data_out_1[77]) );
  DFFHQX1 data_out_1_reg_76_ ( .D(n891), .CK(clk), .Q(data_out_1[76]) );
  DFFHQX1 data_out_1_reg_75_ ( .D(n892), .CK(clk), .Q(data_out_1[75]) );
  DFFHQX1 data_out_1_reg_74_ ( .D(n893), .CK(clk), .Q(data_out_1[74]) );
  DFFHQX1 data_out_1_reg_72_ ( .D(n895), .CK(clk), .Q(data_out_1[72]) );
  DFFHQX1 data_out_1_reg_54_ ( .D(n913), .CK(clk), .Q(data_out_1[54]) );
  DFFHQX1 data_out_1_reg_36_ ( .D(n931), .CK(clk), .Q(data_out_1[36]) );
  DFFHQX1 data_out_1_reg_87_ ( .D(n880), .CK(clk), .Q(data_out_1[87]) );
  DFFHQX1 data_out_1_reg_70_ ( .D(n897), .CK(clk), .Q(data_out_1[70]) );
  DFFHQX1 data_out_1_reg_135_ ( .D(n832), .CK(clk), .Q(data_out_1[135]) );
  DFFHQX1 data_out_1_reg_53_ ( .D(n914), .CK(clk), .Q(data_out_1[53]) );
  DFFHQX1 data_out_1_reg_121_ ( .D(n846), .CK(clk), .Q(data_out_1[121]) );
  DFFHQX1 data_out_1_reg_86_ ( .D(n881), .CK(clk), .Q(data_out_1[86]) );
  DFFHQX1 data_out_1_reg_35_ ( .D(n932), .CK(clk), .Q(data_out_1[35]) );
  DFFHQX1 data_out_1_reg_104_ ( .D(n863), .CK(clk), .Q(data_out_1[104]) );
  DFFHQX1 data_out_1_reg_103_ ( .D(n864), .CK(clk), .Q(data_out_1[103]) );
  DFFHQX1 data_out_1_reg_34_ ( .D(n933), .CK(clk), .Q(data_out_1[34]) );
  DFFHQX4 data_out_1_reg_96_ ( .D(n871), .CK(clk), .Q(data_out_1[96]) );
  DFFHQX4 data_out_1_reg_95_ ( .D(n872), .CK(clk), .Q(data_out_1[95]) );
  DFFHQX4 data_out_1_reg_93_ ( .D(n874), .CK(clk), .Q(data_out_1[93]) );
  DFFHQX4 data_out_1_reg_92_ ( .D(n875), .CK(clk), .Q(data_out_1[92]) );
  DFFHQX4 data_out_1_reg_90_ ( .D(n877), .CK(clk), .Q(data_out_1[90]) );
  DFFHQX4 data_out_1_reg_88_ ( .D(n879), .CK(clk), .Q(data_out_1[88]) );
  DFFHQX4 data_out_1_reg_52_ ( .D(n915), .CK(clk), .Q(data_out_1[52]) );
  DFFHQX4 data_out_1_reg_89_ ( .D(n878), .CK(clk), .Q(data_out_1[89]) );
  DFFHQXL data_out_1_reg_132_ ( .D(n835), .CK(clk), .Q(data_out_1[132]) );
  DFFHQXL data_out_1_reg_66_ ( .D(n901), .CK(clk), .Q(data_out_1[66]) );
  DFFHQXL data_out_1_reg_47_ ( .D(n920), .CK(clk), .Q(data_out_1[47]) );
  DFFHQXL data_out_1_reg_131_ ( .D(n836), .CK(clk), .Q(data_out_1[131]) );
  DFFHQXL data_out_1_reg_45_ ( .D(n922), .CK(clk), .Q(data_out_1[45]) );
  DFFHQXL data_out_1_reg_44_ ( .D(n923), .CK(clk), .Q(data_out_1[44]) );
  DFFHQXL data_out_1_reg_43_ ( .D(n924), .CK(clk), .Q(data_out_1[43]) );
  DFFHQXL data_out_1_reg_42_ ( .D(n925), .CK(clk), .Q(data_out_1[42]) );
  DFFHQXL data_out_1_reg_41_ ( .D(n926), .CK(clk), .Q(data_out_1[41]) );
  DFFHQXL data_out_1_reg_40_ ( .D(n927), .CK(clk), .Q(data_out_1[40]) );
  DFFHQXL data_out_1_reg_57_ ( .D(n910), .CK(clk), .Q(data_out_1[57]) );
  DFFHQXL data_out_1_reg_91_ ( .D(n876), .CK(clk), .Q(data_out_1[91]) );
  DFFHQXL data_out_1_reg_39_ ( .D(n928), .CK(clk), .Q(data_out_1[39]) );
  DFFHQXL data_out_1_reg_38_ ( .D(n929), .CK(clk), .Q(data_out_1[38]) );
  DFFHQXL data_out_1_reg_37_ ( .D(n930), .CK(clk), .Q(data_out_1[37]) );
  DFFHQX1 data_out_1_reg_65_ ( .D(n902), .CK(clk), .Q(data_out_1[65]) );
  OR2X2 U4 ( .A(n830), .B(n828), .Y(n1) );
  OR2X2 U5 ( .A(n829), .B(n826), .Y(n2) );
  OR2X2 U6 ( .A(n826), .B(n830), .Y(n3) );
  OR2X2 U7 ( .A(n824), .B(n829), .Y(n4) );
  OR2X2 U8 ( .A(n824), .B(n830), .Y(n5) );
  OR2X2 U9 ( .A(n825), .B(n829), .Y(n6) );
  OR2X2 U10 ( .A(n825), .B(n830), .Y(n7) );
  OR2X2 U11 ( .A(n828), .B(n829), .Y(n8) );
  AOI22XL U12 ( .A0(R3[0]), .A1(n1042), .B0(data_out_1[0]), .B1(n1018), .Y(
        n822) );
  AOI22XL U13 ( .A0(R3[1]), .A1(n1042), .B0(data_out_1[1]), .B1(n1018), .Y(
        n820) );
  AOI22XL U14 ( .A0(R3[2]), .A1(n1042), .B0(data_out_1[2]), .B1(n1018), .Y(
        n818) );
  AOI22XL U15 ( .A0(R3[3]), .A1(n1042), .B0(data_out_1[3]), .B1(n1018), .Y(
        n816) );
  AOI22XL U16 ( .A0(R15[14]), .A1(n1034), .B0(data_out_1[116]), .B1(n1027), 
        .Y(n590) );
  AOI22XL U17 ( .A0(R15[15]), .A1(n1034), .B0(data_out_1[117]), .B1(n1027), 
        .Y(n588) );
  AOI22XL U18 ( .A0(R11[13]), .A1(n1037), .B0(data_out_1[81]), .B1(n1023), .Y(
        n660) );
  AOI22XL U19 ( .A0(R11[14]), .A1(n1037), .B0(data_out_1[82]), .B1(n1023), .Y(
        n658) );
  AOI22XL U20 ( .A0(R11[15]), .A1(n1037), .B0(data_out_1[83]), .B1(n1023), .Y(
        n656) );
  AOI22XL U21 ( .A0(R11[30]), .A1(n1035), .B0(data_out_1[98]), .B1(n1027), .Y(
        n626) );
  AOI22XL U22 ( .A0(R11[31]), .A1(n1035), .B0(data_out_1[99]), .B1(n1027), .Y(
        n624) );
  AOI22XL U23 ( .A0(R11[32]), .A1(n1035), .B0(data_out_1[100]), .B1(n1027), 
        .Y(n622) );
  AOI22XL U24 ( .A0(R7[13]), .A1(n1039), .B0(data_out_1[47]), .B1(n1021), .Y(
        n728) );
  AOI22XL U25 ( .A0(R7[14]), .A1(n1039), .B0(data_out_1[48]), .B1(n1022), .Y(
        n726) );
  AOI22XL U26 ( .A0(R7[15]), .A1(n1039), .B0(data_out_1[49]), .B1(n1022), .Y(
        n724) );
  AOI22XL U27 ( .A0(R3[17]), .A1(n1041), .B0(data_out_1[17]), .B1(n1019), .Y(
        n788) );
  AOI22XL U28 ( .A0(R3[18]), .A1(n1041), .B0(data_out_1[18]), .B1(n1019), .Y(
        n786) );
  AOI22XL U29 ( .A0(R3[19]), .A1(n1041), .B0(data_out_1[19]), .B1(n1019), .Y(
        n784) );
  AOI22XL U30 ( .A0(R3[20]), .A1(n1041), .B0(data_out_1[20]), .B1(n1019), .Y(
        n782) );
  AOI22XL U31 ( .A0(R15[31]), .A1(n1033), .B0(data_out_1[133]), .B1(n1023), 
        .Y(n556) );
  AOI22XL U32 ( .A0(R15[32]), .A1(n1033), .B0(data_out_1[134]), .B1(n1027), 
        .Y(n554) );
  INVX1 U33 ( .A(n1026), .Y(n1025) );
  INVX1 U34 ( .A(n1026), .Y(n1023) );
  INVX1 U35 ( .A(n1026), .Y(n1024) );
  INVX1 U36 ( .A(n9), .Y(n1021) );
  INVX1 U37 ( .A(n9), .Y(n1022) );
  INVX1 U38 ( .A(n9), .Y(n1018) );
  INVX1 U39 ( .A(n9), .Y(n1019) );
  INVX1 U40 ( .A(n9), .Y(n1020) );
  INVX1 U41 ( .A(n1027), .Y(n1026) );
  INVX1 U42 ( .A(n9), .Y(n1027) );
  CLKINVX3 U43 ( .A(n1032), .Y(n1028) );
  CLKINVX3 U44 ( .A(n1017), .Y(n1013) );
  CLKINVX3 U45 ( .A(n1012), .Y(n1008) );
  OR4X2 U46 ( .A(n1013), .B(n1008), .C(n1028), .D(n1033), .Y(n9) );
  CLKINVX3 U47 ( .A(n1012), .Y(n1010) );
  CLKINVX3 U48 ( .A(n1012), .Y(n1009) );
  CLKINVX3 U49 ( .A(n1012), .Y(n1011) );
  CLKINVX3 U50 ( .A(n1032), .Y(n1031) );
  INVX1 U51 ( .A(n1), .Y(n1034) );
  INVX1 U52 ( .A(n1), .Y(n1037) );
  INVX1 U53 ( .A(n1), .Y(n1036) );
  INVX1 U54 ( .A(n1), .Y(n1035) );
  INVX1 U55 ( .A(n1), .Y(n1039) );
  INVX1 U56 ( .A(n1), .Y(n1038) );
  INVX1 U57 ( .A(n1), .Y(n1041) );
  INVX1 U58 ( .A(n1), .Y(n1040) );
  CLKINVX3 U59 ( .A(n1032), .Y(n1029) );
  CLKINVX3 U60 ( .A(n1032), .Y(n1030) );
  INVX1 U61 ( .A(n1), .Y(n1042) );
  CLKINVX3 U62 ( .A(n1017), .Y(n1014) );
  CLKINVX3 U63 ( .A(n1017), .Y(n1015) );
  CLKINVX3 U64 ( .A(n1017), .Y(n1016) );
  INVX1 U65 ( .A(n1007), .Y(n1005) );
  INVX1 U66 ( .A(n1004), .Y(n1002) );
  INVX1 U67 ( .A(n1001), .Y(n999) );
  INVX1 U68 ( .A(n998), .Y(n996) );
  INVX1 U69 ( .A(n995), .Y(n993) );
  INVX1 U70 ( .A(n2), .Y(n991) );
  INVX1 U71 ( .A(n2), .Y(n992) );
  INVX1 U72 ( .A(n4), .Y(n990) );
  INVX1 U73 ( .A(n6), .Y(n988) );
  INVX1 U74 ( .A(n8), .Y(n986) );
  INVX1 U75 ( .A(n3), .Y(n984) );
  INVX1 U76 ( .A(n5), .Y(n982) );
  INVX1 U77 ( .A(n7), .Y(n980) );
  INVX1 U78 ( .A(n1007), .Y(n1006) );
  INVX1 U79 ( .A(n1004), .Y(n1003) );
  INVX1 U80 ( .A(n1001), .Y(n1000) );
  INVX1 U81 ( .A(n998), .Y(n997) );
  INVX1 U82 ( .A(n995), .Y(n994) );
  INVX1 U83 ( .A(n1), .Y(n1033) );
  INVX1 U84 ( .A(N230), .Y(n1032) );
  INVX1 U85 ( .A(n969), .Y(n1012) );
  INVX1 U86 ( .A(n968), .Y(n1017) );
  INVX1 U87 ( .A(n4), .Y(n989) );
  INVX1 U88 ( .A(n6), .Y(n987) );
  INVX1 U89 ( .A(n8), .Y(n985) );
  INVX1 U90 ( .A(n3), .Y(n983) );
  INVX1 U91 ( .A(n5), .Y(n981) );
  INVX1 U92 ( .A(n7), .Y(n979) );
  INVX1 U93 ( .A(n970), .Y(n1007) );
  INVX1 U94 ( .A(n971), .Y(n1004) );
  INVX1 U95 ( .A(n972), .Y(n1001) );
  INVX1 U96 ( .A(n973), .Y(n998) );
  INVX1 U97 ( .A(n974), .Y(n995) );
  NOR3X1 U98 ( .A(n1045), .B(n1044), .C(n825), .Y(n969) );
  NOR3X1 U99 ( .A(n1045), .B(n1044), .C(n824), .Y(n968) );
  NOR3X1 U100 ( .A(n1044), .B(n826), .C(n1045), .Y(N230) );
  NAND2X1 U101 ( .A(n1044), .B(n1045), .Y(n830) );
  NOR3X1 U102 ( .A(n1045), .B(n1044), .C(n828), .Y(n970) );
  OAI211X1 U103 ( .A0(n831), .A1(n1045), .B0(n827), .C0(n2), .Y(N15) );
  NOR2X1 U104 ( .A(n826), .B(n827), .Y(n971) );
  NOR2X1 U105 ( .A(n824), .B(n827), .Y(n972) );
  NOR2X1 U106 ( .A(n825), .B(n827), .Y(n973) );
  NOR2X1 U107 ( .A(n828), .B(n827), .Y(n974) );
  NAND2X1 U108 ( .A(n824), .B(n825), .Y(N13) );
  INVX1 U109 ( .A(counter[2]), .Y(n1044) );
  INVX1 U110 ( .A(counter[3]), .Y(n1045) );
  NAND2X1 U111 ( .A(counter[0]), .B(n1043), .Y(n825) );
  NAND2X1 U112 ( .A(counter[1]), .B(counter[0]), .Y(n826) );
  NAND2X1 U113 ( .A(counter[1]), .B(n550), .Y(n824) );
  NAND2X1 U114 ( .A(n550), .B(n1043), .Y(n828) );
  INVX1 U115 ( .A(counter[1]), .Y(n1043) );
  NAND2X1 U116 ( .A(n618), .B(n619), .Y(n865) );
  AOI222X1 U117 ( .A0(R12[0]), .A1(n1009), .B0(R14[0]), .B1(n1030), .C0(R13[0]), .C1(n1014), .Y(n619) );
  AOI22XL U118 ( .A0(R15[0]), .A1(n1035), .B0(data_out_1[102]), .B1(n1021), 
        .Y(n618) );
  NAND2X1 U119 ( .A(n616), .B(n617), .Y(n864) );
  AOI222X1 U120 ( .A0(R12[1]), .A1(n1009), .B0(R14[1]), .B1(n1030), .C0(R13[1]), .C1(n1014), .Y(n617) );
  AOI22XL U121 ( .A0(R15[1]), .A1(n1035), .B0(data_out_1[103]), .B1(n1027), 
        .Y(n616) );
  NAND2X1 U122 ( .A(n614), .B(n615), .Y(n863) );
  AOI222X1 U123 ( .A0(R12[2]), .A1(n1010), .B0(R14[2]), .B1(n1029), .C0(R13[2]), .C1(n1014), .Y(n615) );
  AOI22XL U124 ( .A0(R15[2]), .A1(n1035), .B0(data_out_1[104]), .B1(n1027), 
        .Y(n614) );
  NAND2X1 U125 ( .A(n612), .B(n613), .Y(n862) );
  AOI222X1 U126 ( .A0(R12[3]), .A1(n1009), .B0(R14[3]), .B1(n1031), .C0(R13[3]), .C1(n1014), .Y(n613) );
  AOI22XL U127 ( .A0(R15[3]), .A1(n1035), .B0(data_out_1[105]), .B1(n1024), 
        .Y(n612) );
  NAND2X1 U128 ( .A(n610), .B(n611), .Y(n861) );
  AOI222X1 U129 ( .A0(R12[4]), .A1(n1011), .B0(R14[4]), .B1(n1028), .C0(R13[4]), .C1(n1014), .Y(n611) );
  AOI22XL U130 ( .A0(R15[4]), .A1(n1035), .B0(data_out_1[106]), .B1(n1021), 
        .Y(n610) );
  NAND2X1 U131 ( .A(n608), .B(n609), .Y(n860) );
  AOI222X1 U132 ( .A0(R12[5]), .A1(n1009), .B0(R14[5]), .B1(n1030), .C0(R13[5]), .C1(n1014), .Y(n609) );
  AOI22XL U133 ( .A0(R15[5]), .A1(n1035), .B0(data_out_1[107]), .B1(n1025), 
        .Y(n608) );
  NAND2X1 U134 ( .A(n606), .B(n607), .Y(n859) );
  AOI222X1 U135 ( .A0(R12[6]), .A1(n1011), .B0(R14[6]), .B1(n1030), .C0(R13[6]), .C1(n1014), .Y(n607) );
  AOI22XL U136 ( .A0(R15[6]), .A1(n1035), .B0(data_out_1[108]), .B1(n1027), 
        .Y(n606) );
  NAND2X1 U137 ( .A(n604), .B(n605), .Y(n858) );
  AOI222X1 U138 ( .A0(R12[7]), .A1(n1010), .B0(R14[7]), .B1(n1029), .C0(R13[7]), .C1(n1014), .Y(n605) );
  AOI22XL U139 ( .A0(R15[7]), .A1(n1035), .B0(data_out_1[109]), .B1(n1027), 
        .Y(n604) );
  NAND2X1 U140 ( .A(n602), .B(n603), .Y(n857) );
  AOI222X1 U141 ( .A0(R12[8]), .A1(n1010), .B0(R14[8]), .B1(n1031), .C0(R13[8]), .C1(n1014), .Y(n603) );
  AOI22XL U142 ( .A0(R15[8]), .A1(n1034), .B0(data_out_1[110]), .B1(n1027), 
        .Y(n602) );
  NAND2X1 U143 ( .A(n600), .B(n601), .Y(n856) );
  AOI222X1 U144 ( .A0(R12[9]), .A1(n1010), .B0(R14[9]), .B1(n1030), .C0(R13[9]), .C1(n1014), .Y(n601) );
  AOI22XL U145 ( .A0(R15[9]), .A1(n1034), .B0(data_out_1[111]), .B1(n1027), 
        .Y(n600) );
  NAND2X1 U146 ( .A(n598), .B(n599), .Y(n855) );
  AOI222X1 U147 ( .A0(R12[10]), .A1(n1009), .B0(R14[10]), .B1(n1029), .C0(
        R13[10]), .C1(n1014), .Y(n599) );
  AOI22XL U148 ( .A0(R15[10]), .A1(n1034), .B0(data_out_1[112]), .B1(n1027), 
        .Y(n598) );
  NAND2X1 U149 ( .A(n596), .B(n597), .Y(n854) );
  AOI222X1 U150 ( .A0(R12[11]), .A1(n1011), .B0(R14[11]), .B1(n1030), .C0(
        R13[11]), .C1(n1014), .Y(n597) );
  AOI22XL U151 ( .A0(R15[11]), .A1(n1034), .B0(data_out_1[113]), .B1(n1027), 
        .Y(n596) );
  NAND2X1 U152 ( .A(n594), .B(n595), .Y(n853) );
  AOI222X1 U153 ( .A0(R12[12]), .A1(n1010), .B0(R14[12]), .B1(n1029), .C0(
        R13[12]), .C1(n1014), .Y(n595) );
  AOI22XL U154 ( .A0(R15[12]), .A1(n1034), .B0(data_out_1[114]), .B1(n1022), 
        .Y(n594) );
  NAND2X1 U155 ( .A(n592), .B(n593), .Y(n852) );
  AOI222X1 U156 ( .A0(R12[13]), .A1(n1009), .B0(R14[13]), .B1(n1030), .C0(
        R13[13]), .C1(n1014), .Y(n593) );
  AOI22XL U157 ( .A0(R15[13]), .A1(n1034), .B0(data_out_1[115]), .B1(n1027), 
        .Y(n592) );
  NAND2X1 U158 ( .A(n590), .B(n591), .Y(n851) );
  AOI222X1 U159 ( .A0(R12[14]), .A1(n1009), .B0(R14[14]), .B1(n1030), .C0(
        R13[14]), .C1(n1014), .Y(n591) );
  NAND2X1 U160 ( .A(n588), .B(n589), .Y(n850) );
  AOI222X1 U161 ( .A0(R12[15]), .A1(n1009), .B0(R14[15]), .B1(n1030), .C0(
        R13[15]), .C1(n1014), .Y(n589) );
  NAND2X1 U162 ( .A(n586), .B(n587), .Y(n849) );
  AOI222X1 U163 ( .A0(R12[16]), .A1(n1009), .B0(R14[16]), .B1(n1028), .C0(
        R13[16]), .C1(n1013), .Y(n587) );
  AOI22XL U164 ( .A0(R15[16]), .A1(n1034), .B0(data_out_1[118]), .B1(n1025), 
        .Y(n586) );
  NAND2X1 U165 ( .A(n584), .B(n585), .Y(n848) );
  AOI222X1 U166 ( .A0(R12[17]), .A1(n1008), .B0(R14[17]), .B1(n1028), .C0(
        R13[17]), .C1(n1013), .Y(n585) );
  AOI22XL U167 ( .A0(R15[17]), .A1(n1034), .B0(data_out_1[119]), .B1(n1024), 
        .Y(n584) );
  NAND2X1 U168 ( .A(n582), .B(n583), .Y(n847) );
  AOI222X1 U169 ( .A0(R12[18]), .A1(n1008), .B0(R14[18]), .B1(n1028), .C0(
        R13[18]), .C1(n1013), .Y(n583) );
  AOI22XL U170 ( .A0(R15[18]), .A1(n1034), .B0(data_out_1[120]), .B1(n1025), 
        .Y(n582) );
  NAND2X1 U171 ( .A(n580), .B(n581), .Y(n846) );
  AOI222X1 U172 ( .A0(R12[19]), .A1(n1008), .B0(R14[19]), .B1(n1028), .C0(
        R13[19]), .C1(n1013), .Y(n581) );
  AOI22XL U173 ( .A0(R15[19]), .A1(n1034), .B0(data_out_1[121]), .B1(n1025), 
        .Y(n580) );
  NAND2X1 U174 ( .A(n578), .B(n579), .Y(n845) );
  AOI222X1 U175 ( .A0(R12[20]), .A1(n1008), .B0(R14[20]), .B1(n1028), .C0(
        R13[20]), .C1(n1013), .Y(n579) );
  AOI22XL U176 ( .A0(R15[20]), .A1(n1034), .B0(data_out_1[122]), .B1(n1025), 
        .Y(n578) );
  NAND2X1 U177 ( .A(n576), .B(n577), .Y(n844) );
  AOI222X1 U178 ( .A0(R12[21]), .A1(n1008), .B0(R14[21]), .B1(n1028), .C0(
        R13[21]), .C1(n1013), .Y(n577) );
  AOI22XL U179 ( .A0(R15[21]), .A1(n1033), .B0(data_out_1[123]), .B1(n1025), 
        .Y(n576) );
  NAND2X1 U180 ( .A(n574), .B(n575), .Y(n843) );
  AOI222X1 U181 ( .A0(R12[22]), .A1(n1008), .B0(R14[22]), .B1(n1028), .C0(
        R13[22]), .C1(n1013), .Y(n575) );
  AOI22XL U182 ( .A0(R15[22]), .A1(n1033), .B0(data_out_1[124]), .B1(n1025), 
        .Y(n574) );
  NAND2X1 U183 ( .A(n572), .B(n573), .Y(n842) );
  AOI222X1 U184 ( .A0(R12[23]), .A1(n1008), .B0(R14[23]), .B1(n1028), .C0(
        R13[23]), .C1(n1013), .Y(n573) );
  AOI22XL U185 ( .A0(R15[23]), .A1(n1033), .B0(data_out_1[125]), .B1(n1025), 
        .Y(n572) );
  NAND2X1 U186 ( .A(n570), .B(n571), .Y(n841) );
  AOI222X1 U187 ( .A0(R12[24]), .A1(n1008), .B0(R14[24]), .B1(n1028), .C0(
        R13[24]), .C1(n1013), .Y(n571) );
  AOI22XL U188 ( .A0(R15[24]), .A1(n1033), .B0(data_out_1[126]), .B1(n1025), 
        .Y(n570) );
  NAND2X1 U189 ( .A(n568), .B(n569), .Y(n840) );
  AOI222X1 U190 ( .A0(R12[25]), .A1(n1008), .B0(R14[25]), .B1(n1028), .C0(
        R13[25]), .C1(n1013), .Y(n569) );
  AOI22XL U191 ( .A0(R15[25]), .A1(n1033), .B0(data_out_1[127]), .B1(n1025), 
        .Y(n568) );
  NAND2X1 U192 ( .A(n566), .B(n567), .Y(n839) );
  AOI222X1 U193 ( .A0(R12[26]), .A1(n1008), .B0(R14[26]), .B1(n1028), .C0(
        R13[26]), .C1(n1013), .Y(n567) );
  AOI22XL U194 ( .A0(R15[26]), .A1(n1033), .B0(data_out_1[128]), .B1(n1025), 
        .Y(n566) );
  NAND2X1 U195 ( .A(n564), .B(n565), .Y(n838) );
  AOI222X1 U196 ( .A0(R12[27]), .A1(n1008), .B0(R14[27]), .B1(n1028), .C0(
        R13[27]), .C1(n1013), .Y(n565) );
  AOI22XL U197 ( .A0(R15[27]), .A1(n1033), .B0(data_out_1[129]), .B1(n1025), 
        .Y(n564) );
  NAND2X1 U198 ( .A(n562), .B(n563), .Y(n837) );
  AOI222X1 U199 ( .A0(R12[28]), .A1(n1008), .B0(R14[28]), .B1(n1028), .C0(
        R13[28]), .C1(n1013), .Y(n563) );
  AOI22XL U200 ( .A0(R15[28]), .A1(n1033), .B0(data_out_1[130]), .B1(n1025), 
        .Y(n562) );
  NAND2X1 U201 ( .A(n560), .B(n561), .Y(n836) );
  AOI222X1 U202 ( .A0(R12[29]), .A1(n1008), .B0(R14[29]), .B1(n1028), .C0(
        R13[29]), .C1(n1013), .Y(n561) );
  AOI22XL U203 ( .A0(R15[29]), .A1(n1033), .B0(data_out_1[131]), .B1(n1025), 
        .Y(n560) );
  NAND2X1 U204 ( .A(n686), .B(n687), .Y(n899) );
  AOI222X1 U205 ( .A0(R8[0]), .A1(n1009), .B0(R10[0]), .B1(n1029), .C0(R9[0]), 
        .C1(n1015), .Y(n687) );
  AOI22XL U206 ( .A0(R11[0]), .A1(n1038), .B0(data_out_1[68]), .B1(n1022), .Y(
        n686) );
  NAND2X1 U207 ( .A(n684), .B(n685), .Y(n898) );
  AOI222X1 U208 ( .A0(R8[1]), .A1(n1009), .B0(R10[1]), .B1(n1031), .C0(R9[1]), 
        .C1(n1016), .Y(n685) );
  AOI22XL U209 ( .A0(R11[1]), .A1(n1038), .B0(data_out_1[69]), .B1(n1021), .Y(
        n684) );
  NAND2X1 U210 ( .A(n682), .B(n683), .Y(n897) );
  AOI222X1 U211 ( .A0(R8[2]), .A1(n1009), .B0(R10[2]), .B1(n1030), .C0(R9[2]), 
        .C1(n1015), .Y(n683) );
  AOI22XL U212 ( .A0(R11[2]), .A1(n1038), .B0(data_out_1[70]), .B1(n1021), .Y(
        n682) );
  NAND2X1 U213 ( .A(n680), .B(n681), .Y(n896) );
  AOI222X1 U214 ( .A0(R8[3]), .A1(n1009), .B0(R10[3]), .B1(n1030), .C0(R9[3]), 
        .C1(n1014), .Y(n681) );
  AOI22XL U215 ( .A0(R11[3]), .A1(n1037), .B0(data_out_1[71]), .B1(n1023), .Y(
        n680) );
  NAND2X1 U216 ( .A(n678), .B(n679), .Y(n895) );
  AOI222X1 U217 ( .A0(R8[4]), .A1(n1009), .B0(R10[4]), .B1(n1030), .C0(R9[4]), 
        .C1(n1014), .Y(n679) );
  AOI22XL U218 ( .A0(R11[4]), .A1(n1037), .B0(data_out_1[72]), .B1(n1023), .Y(
        n678) );
  NAND2X1 U219 ( .A(n676), .B(n677), .Y(n894) );
  AOI222X1 U220 ( .A0(R8[5]), .A1(n1009), .B0(R10[5]), .B1(n1029), .C0(R9[5]), 
        .C1(n1015), .Y(n677) );
  AOI22XL U221 ( .A0(R11[5]), .A1(n1037), .B0(data_out_1[73]), .B1(n1023), .Y(
        n676) );
  NAND2X1 U222 ( .A(n674), .B(n675), .Y(n893) );
  AOI222X1 U223 ( .A0(R8[6]), .A1(n1009), .B0(R10[6]), .B1(n1029), .C0(R9[6]), 
        .C1(n1015), .Y(n675) );
  AOI22XL U224 ( .A0(R11[6]), .A1(n1037), .B0(data_out_1[74]), .B1(n1023), .Y(
        n674) );
  NAND2X1 U225 ( .A(n672), .B(n673), .Y(n892) );
  AOI222X1 U226 ( .A0(R8[7]), .A1(n1009), .B0(R10[7]), .B1(n1030), .C0(R9[7]), 
        .C1(n1016), .Y(n673) );
  AOI22XL U227 ( .A0(R11[7]), .A1(n1037), .B0(data_out_1[75]), .B1(n1023), .Y(
        n672) );
  NAND2X1 U228 ( .A(n670), .B(n671), .Y(n891) );
  AOI222X1 U229 ( .A0(R8[8]), .A1(n1009), .B0(R10[8]), .B1(n1029), .C0(R9[8]), 
        .C1(n1014), .Y(n671) );
  AOI22XL U230 ( .A0(R11[8]), .A1(n1037), .B0(data_out_1[76]), .B1(n1023), .Y(
        n670) );
  NAND2X1 U231 ( .A(n668), .B(n669), .Y(n890) );
  AOI222X1 U232 ( .A0(R8[9]), .A1(n1009), .B0(R10[9]), .B1(n1029), .C0(R9[9]), 
        .C1(n1015), .Y(n669) );
  AOI22XL U233 ( .A0(R11[9]), .A1(n1037), .B0(data_out_1[77]), .B1(n1023), .Y(
        n668) );
  NAND2X1 U234 ( .A(n666), .B(n667), .Y(n889) );
  AOI222X1 U235 ( .A0(R8[10]), .A1(n1009), .B0(R10[10]), .B1(n1030), .C0(
        R9[10]), .C1(n1016), .Y(n667) );
  AOI22XL U236 ( .A0(R11[10]), .A1(n1037), .B0(data_out_1[78]), .B1(n1023), 
        .Y(n666) );
  NAND2X1 U237 ( .A(n664), .B(n665), .Y(n888) );
  AOI222X1 U238 ( .A0(R8[11]), .A1(n1009), .B0(R10[11]), .B1(n1031), .C0(
        R9[11]), .C1(n1014), .Y(n665) );
  AOI22XL U239 ( .A0(R11[11]), .A1(n1037), .B0(data_out_1[79]), .B1(n1023), 
        .Y(n664) );
  NAND2X1 U240 ( .A(n662), .B(n663), .Y(n887) );
  AOI222X1 U241 ( .A0(R8[12]), .A1(n1009), .B0(R10[12]), .B1(n1029), .C0(
        R9[12]), .C1(n1015), .Y(n663) );
  AOI22XL U242 ( .A0(R11[12]), .A1(n1037), .B0(data_out_1[80]), .B1(n1023), 
        .Y(n662) );
  NAND2X1 U243 ( .A(n660), .B(n661), .Y(n886) );
  AOI222X1 U244 ( .A0(R8[13]), .A1(n1009), .B0(R10[13]), .B1(n1031), .C0(
        R9[13]), .C1(n1016), .Y(n661) );
  NAND2X1 U245 ( .A(n658), .B(n659), .Y(n885) );
  AOI222X1 U246 ( .A0(R8[14]), .A1(n1009), .B0(R10[14]), .B1(n1029), .C0(
        R9[14]), .C1(n1016), .Y(n659) );
  NAND2X1 U247 ( .A(n656), .B(n657), .Y(n884) );
  AOI222X1 U248 ( .A0(R8[15]), .A1(n1010), .B0(R10[15]), .B1(n1029), .C0(
        R9[15]), .C1(n1015), .Y(n657) );
  NAND2X1 U249 ( .A(n654), .B(n655), .Y(n883) );
  AOI222X1 U250 ( .A0(R8[16]), .A1(n1009), .B0(R10[16]), .B1(n1029), .C0(
        R9[16]), .C1(n1016), .Y(n655) );
  AOI22XL U251 ( .A0(R11[16]), .A1(n1036), .B0(data_out_1[84]), .B1(n1024), 
        .Y(n654) );
  NAND2X1 U252 ( .A(n652), .B(n653), .Y(n882) );
  AOI222X1 U253 ( .A0(R8[17]), .A1(n1009), .B0(R10[17]), .B1(n1029), .C0(
        R9[17]), .C1(n1015), .Y(n653) );
  AOI22XL U254 ( .A0(R11[17]), .A1(n1036), .B0(data_out_1[85]), .B1(n1024), 
        .Y(n652) );
  NAND2X1 U255 ( .A(n650), .B(n651), .Y(n881) );
  AOI222X1 U256 ( .A0(R8[18]), .A1(n1011), .B0(R10[18]), .B1(n1029), .C0(
        R9[18]), .C1(n1014), .Y(n651) );
  AOI22XL U257 ( .A0(R11[18]), .A1(n1036), .B0(data_out_1[86]), .B1(n1024), 
        .Y(n650) );
  NAND2X1 U258 ( .A(n648), .B(n649), .Y(n880) );
  AOI222X1 U259 ( .A0(R8[19]), .A1(n1009), .B0(R10[19]), .B1(n1029), .C0(
        R9[19]), .C1(n1016), .Y(n649) );
  AOI22XL U260 ( .A0(R11[19]), .A1(n1036), .B0(data_out_1[87]), .B1(n1024), 
        .Y(n648) );
  NAND2X1 U261 ( .A(n646), .B(n647), .Y(n879) );
  AOI222X1 U262 ( .A0(R8[20]), .A1(n1011), .B0(R10[20]), .B1(n1029), .C0(
        R9[20]), .C1(n1016), .Y(n647) );
  AOI22XL U263 ( .A0(R11[20]), .A1(n1036), .B0(data_out_1[88]), .B1(n1024), 
        .Y(n646) );
  NAND2X1 U264 ( .A(n644), .B(n645), .Y(n878) );
  AOI222X1 U265 ( .A0(R8[21]), .A1(n1010), .B0(R10[21]), .B1(n1029), .C0(
        R9[21]), .C1(n1016), .Y(n645) );
  AOI22XL U266 ( .A0(R11[21]), .A1(n1036), .B0(data_out_1[89]), .B1(n1024), 
        .Y(n644) );
  NAND2X1 U267 ( .A(n642), .B(n643), .Y(n877) );
  AOI222X1 U268 ( .A0(R8[22]), .A1(n1010), .B0(R10[22]), .B1(n1029), .C0(
        R9[22]), .C1(n1015), .Y(n643) );
  AOI22XL U269 ( .A0(R11[22]), .A1(n1036), .B0(data_out_1[90]), .B1(n1024), 
        .Y(n642) );
  NAND2X1 U270 ( .A(n640), .B(n641), .Y(n876) );
  AOI222X1 U271 ( .A0(R8[23]), .A1(n1011), .B0(R10[23]), .B1(n1029), .C0(
        R9[23]), .C1(n1015), .Y(n641) );
  AOI22XL U272 ( .A0(R11[23]), .A1(n1036), .B0(data_out_1[91]), .B1(n1024), 
        .Y(n640) );
  NAND2X1 U273 ( .A(n638), .B(n639), .Y(n875) );
  AOI222X1 U274 ( .A0(R8[24]), .A1(n1009), .B0(R10[24]), .B1(n1029), .C0(
        R9[24]), .C1(n1014), .Y(n639) );
  AOI22XL U275 ( .A0(R11[24]), .A1(n1036), .B0(data_out_1[92]), .B1(n1024), 
        .Y(n638) );
  NAND2X1 U276 ( .A(n636), .B(n637), .Y(n874) );
  AOI222X1 U277 ( .A0(R8[25]), .A1(n1011), .B0(R10[25]), .B1(n1029), .C0(
        R9[25]), .C1(n1016), .Y(n637) );
  AOI22XL U278 ( .A0(R11[25]), .A1(n1036), .B0(data_out_1[93]), .B1(n1024), 
        .Y(n636) );
  NAND2X1 U279 ( .A(n634), .B(n635), .Y(n873) );
  AOI222X1 U280 ( .A0(R8[26]), .A1(n1010), .B0(R10[26]), .B1(n1029), .C0(
        R9[26]), .C1(n1015), .Y(n635) );
  AOI22XL U281 ( .A0(R11[26]), .A1(n1036), .B0(data_out_1[94]), .B1(n1024), 
        .Y(n634) );
  NAND2X1 U282 ( .A(n632), .B(n633), .Y(n872) );
  AOI222X1 U283 ( .A0(R8[27]), .A1(n1011), .B0(R10[27]), .B1(n1029), .C0(
        R9[27]), .C1(n1014), .Y(n633) );
  AOI22XL U284 ( .A0(R11[27]), .A1(n1036), .B0(data_out_1[95]), .B1(n1024), 
        .Y(n632) );
  NAND2X1 U285 ( .A(n630), .B(n631), .Y(n871) );
  AOI222X1 U286 ( .A0(R8[28]), .A1(n1009), .B0(R10[28]), .B1(n1029), .C0(
        R9[28]), .C1(n1016), .Y(n631) );
  AOI22XL U287 ( .A0(R11[28]), .A1(n1036), .B0(data_out_1[96]), .B1(n1019), 
        .Y(n630) );
  NAND2X1 U288 ( .A(n628), .B(n629), .Y(n870) );
  AOI222X1 U289 ( .A0(R8[29]), .A1(n1011), .B0(R10[29]), .B1(n1029), .C0(
        R9[29]), .C1(n1015), .Y(n629) );
  AOI22XL U290 ( .A0(R11[29]), .A1(n1035), .B0(data_out_1[97]), .B1(n1022), 
        .Y(n628) );
  NAND2X1 U291 ( .A(n626), .B(n627), .Y(n869) );
  AOI222X1 U292 ( .A0(R8[30]), .A1(n1010), .B0(R10[30]), .B1(n1029), .C0(
        R9[30]), .C1(n1015), .Y(n627) );
  NAND2X1 U293 ( .A(n624), .B(n625), .Y(n868) );
  AOI222X1 U294 ( .A0(R8[31]), .A1(n1011), .B0(R10[31]), .B1(n1029), .C0(
        R9[31]), .C1(n1016), .Y(n625) );
  NAND2X1 U295 ( .A(n622), .B(n623), .Y(n867) );
  AOI222X1 U296 ( .A0(R8[32]), .A1(n1011), .B0(R10[32]), .B1(n1031), .C0(
        R9[32]), .C1(n1014), .Y(n623) );
  NAND2X1 U297 ( .A(n620), .B(n621), .Y(n866) );
  AOI222X1 U298 ( .A0(R8[33]), .A1(n1011), .B0(R10[33]), .B1(n1029), .C0(
        R9[33]), .C1(n1014), .Y(n621) );
  AOI22XL U299 ( .A0(R11[33]), .A1(n1035), .B0(data_out_1[101]), .B1(n1018), 
        .Y(n620) );
  NAND2X1 U300 ( .A(n754), .B(n755), .Y(n933) );
  AOI222X1 U301 ( .A0(R4[0]), .A1(n1011), .B0(R6[0]), .B1(n1029), .C0(R5[0]), 
        .C1(n1015), .Y(n755) );
  AOI22XL U302 ( .A0(R7[0]), .A1(n1040), .B0(data_out_1[34]), .B1(n1020), .Y(
        n754) );
  NAND2X1 U303 ( .A(n752), .B(n753), .Y(n932) );
  AOI222X1 U304 ( .A0(R4[1]), .A1(n1009), .B0(R6[1]), .B1(n1029), .C0(R5[1]), 
        .C1(n1015), .Y(n753) );
  AOI22XL U305 ( .A0(R7[1]), .A1(n1040), .B0(data_out_1[35]), .B1(n1020), .Y(
        n752) );
  NAND2X1 U306 ( .A(n750), .B(n751), .Y(n931) );
  AOI222X1 U307 ( .A0(R4[2]), .A1(n1010), .B0(R6[2]), .B1(n1029), .C0(R5[2]), 
        .C1(n1015), .Y(n751) );
  AOI22XL U308 ( .A0(R7[2]), .A1(n1040), .B0(data_out_1[36]), .B1(n1021), .Y(
        n750) );
  NAND2X1 U309 ( .A(n748), .B(n749), .Y(n930) );
  AOI222X1 U310 ( .A0(R4[3]), .A1(n1010), .B0(R6[3]), .B1(n1029), .C0(R5[3]), 
        .C1(n1015), .Y(n749) );
  AOI22XL U311 ( .A0(R7[3]), .A1(n1040), .B0(data_out_1[37]), .B1(n1021), .Y(
        n748) );
  NAND2X1 U312 ( .A(n746), .B(n747), .Y(n929) );
  AOI222X1 U313 ( .A0(R4[4]), .A1(n1011), .B0(R6[4]), .B1(N230), .C0(R5[4]), 
        .C1(n1015), .Y(n747) );
  AOI22XL U314 ( .A0(R7[4]), .A1(n1040), .B0(data_out_1[38]), .B1(n1021), .Y(
        n746) );
  NAND2X1 U315 ( .A(n744), .B(n745), .Y(n928) );
  AOI222X1 U316 ( .A0(R4[5]), .A1(n1009), .B0(R6[5]), .B1(n1030), .C0(R5[5]), 
        .C1(n1015), .Y(n745) );
  AOI22XL U317 ( .A0(R7[5]), .A1(n1040), .B0(data_out_1[39]), .B1(n1021), .Y(
        n744) );
  NAND2X1 U318 ( .A(n742), .B(n743), .Y(n927) );
  AOI222X1 U319 ( .A0(R4[6]), .A1(n1010), .B0(R6[6]), .B1(N230), .C0(R5[6]), 
        .C1(n1015), .Y(n743) );
  AOI22XL U320 ( .A0(R7[6]), .A1(n1040), .B0(data_out_1[40]), .B1(n1021), .Y(
        n742) );
  NAND2X1 U321 ( .A(n740), .B(n741), .Y(n926) );
  AOI222X1 U322 ( .A0(R4[7]), .A1(n1011), .B0(R6[7]), .B1(n1029), .C0(R5[7]), 
        .C1(n1015), .Y(n741) );
  AOI22XL U323 ( .A0(R7[7]), .A1(n1040), .B0(data_out_1[41]), .B1(n1021), .Y(
        n740) );
  NAND2X1 U324 ( .A(n738), .B(n739), .Y(n925) );
  AOI222X1 U325 ( .A0(R4[8]), .A1(n1009), .B0(R6[8]), .B1(n1029), .C0(R5[8]), 
        .C1(n1015), .Y(n739) );
  AOI22XL U326 ( .A0(R7[8]), .A1(n1040), .B0(data_out_1[42]), .B1(n1021), .Y(
        n738) );
  NAND2X1 U327 ( .A(n736), .B(n737), .Y(n924) );
  AOI222X1 U328 ( .A0(R4[9]), .A1(n1010), .B0(R6[9]), .B1(n1030), .C0(R5[9]), 
        .C1(n1015), .Y(n737) );
  AOI22XL U329 ( .A0(R7[9]), .A1(n1040), .B0(data_out_1[43]), .B1(n1021), .Y(
        n736) );
  NAND2X1 U330 ( .A(n734), .B(n735), .Y(n923) );
  AOI222X1 U331 ( .A0(R4[10]), .A1(n1008), .B0(R6[10]), .B1(N230), .C0(R5[10]), 
        .C1(n1015), .Y(n735) );
  AOI22XL U332 ( .A0(R7[10]), .A1(n1040), .B0(data_out_1[44]), .B1(n1021), .Y(
        n734) );
  NAND2X1 U333 ( .A(n732), .B(n733), .Y(n922) );
  AOI222X1 U334 ( .A0(R4[11]), .A1(n1008), .B0(R6[11]), .B1(n1029), .C0(R5[11]), .C1(n1015), .Y(n733) );
  AOI22XL U335 ( .A0(R7[11]), .A1(n1040), .B0(data_out_1[45]), .B1(n1021), .Y(
        n732) );
  NAND2X1 U336 ( .A(n730), .B(n731), .Y(n921) );
  AOI222X1 U337 ( .A0(R4[12]), .A1(n1011), .B0(R6[12]), .B1(n1030), .C0(R5[12]), .C1(n1015), .Y(n731) );
  AOI22XL U338 ( .A0(R7[12]), .A1(n1039), .B0(data_out_1[46]), .B1(n1021), .Y(
        n730) );
  NAND2X1 U339 ( .A(n728), .B(n729), .Y(n920) );
  AOI222X1 U340 ( .A0(R4[13]), .A1(n1009), .B0(R6[13]), .B1(N230), .C0(R5[13]), 
        .C1(n1014), .Y(n729) );
  NAND2X1 U341 ( .A(n726), .B(n727), .Y(n919) );
  AOI222X1 U342 ( .A0(R4[14]), .A1(n1010), .B0(R6[14]), .B1(n1030), .C0(R5[14]), .C1(n1014), .Y(n727) );
  NAND2X1 U343 ( .A(n724), .B(n725), .Y(n918) );
  AOI222X1 U344 ( .A0(R4[15]), .A1(n1010), .B0(R6[15]), .B1(n1029), .C0(R5[15]), .C1(n1014), .Y(n725) );
  NAND2X1 U345 ( .A(n722), .B(n723), .Y(n917) );
  AOI222X1 U346 ( .A0(R4[16]), .A1(n1010), .B0(R6[16]), .B1(n1031), .C0(R5[16]), .C1(n1014), .Y(n723) );
  AOI22XL U347 ( .A0(R7[16]), .A1(n1039), .B0(data_out_1[50]), .B1(n1022), .Y(
        n722) );
  NAND2X1 U348 ( .A(n720), .B(n721), .Y(n916) );
  AOI222X1 U349 ( .A0(R4[17]), .A1(n1010), .B0(R6[17]), .B1(n1030), .C0(R5[17]), .C1(n1014), .Y(n721) );
  AOI22XL U350 ( .A0(R7[17]), .A1(n1039), .B0(data_out_1[51]), .B1(n1022), .Y(
        n720) );
  NAND2X1 U351 ( .A(n718), .B(n719), .Y(n915) );
  AOI222X1 U352 ( .A0(R4[18]), .A1(n1010), .B0(R6[18]), .B1(n1029), .C0(R5[18]), .C1(n1014), .Y(n719) );
  AOI22XL U353 ( .A0(R7[18]), .A1(n1039), .B0(data_out_1[52]), .B1(n1022), .Y(
        n718) );
  NAND2X1 U354 ( .A(n716), .B(n717), .Y(n914) );
  AOI222X1 U355 ( .A0(R4[19]), .A1(n1010), .B0(R6[19]), .B1(n1031), .C0(R5[19]), .C1(n1014), .Y(n717) );
  AOI22XL U356 ( .A0(R7[19]), .A1(n1039), .B0(data_out_1[53]), .B1(n1022), .Y(
        n716) );
  NAND2X1 U357 ( .A(n714), .B(n715), .Y(n913) );
  AOI222X1 U358 ( .A0(R4[20]), .A1(n1010), .B0(R6[20]), .B1(n1030), .C0(R5[20]), .C1(n1014), .Y(n715) );
  AOI22XL U359 ( .A0(R7[20]), .A1(n1039), .B0(data_out_1[54]), .B1(n1022), .Y(
        n714) );
  NAND2X1 U360 ( .A(n712), .B(n713), .Y(n912) );
  AOI222X1 U361 ( .A0(R4[21]), .A1(n1010), .B0(R6[21]), .B1(n1031), .C0(R5[21]), .C1(n1014), .Y(n713) );
  AOI22XL U362 ( .A0(R7[21]), .A1(n1039), .B0(data_out_1[55]), .B1(n1022), .Y(
        n712) );
  NAND2X1 U363 ( .A(n710), .B(n711), .Y(n911) );
  AOI222X1 U364 ( .A0(R4[22]), .A1(n1010), .B0(R6[22]), .B1(n1030), .C0(R5[22]), .C1(n1014), .Y(n711) );
  AOI22XL U365 ( .A0(R7[22]), .A1(n1039), .B0(data_out_1[56]), .B1(n1022), .Y(
        n710) );
  NAND2X1 U366 ( .A(n708), .B(n709), .Y(n910) );
  AOI222X1 U367 ( .A0(R4[23]), .A1(n1010), .B0(R6[23]), .B1(n1028), .C0(R5[23]), .C1(n1015), .Y(n709) );
  AOI22XL U368 ( .A0(R7[23]), .A1(n1039), .B0(data_out_1[57]), .B1(n1022), .Y(
        n708) );
  NAND2X1 U369 ( .A(n706), .B(n707), .Y(n909) );
  AOI222X1 U370 ( .A0(R4[24]), .A1(n1010), .B0(R6[24]), .B1(n1029), .C0(R5[24]), .C1(n1014), .Y(n707) );
  AOI22XL U371 ( .A0(R7[24]), .A1(n1038), .B0(data_out_1[58]), .B1(n1022), .Y(
        n706) );
  NAND2X1 U372 ( .A(n704), .B(n705), .Y(n908) );
  AOI222X1 U373 ( .A0(R4[25]), .A1(n1010), .B0(R6[25]), .B1(n1031), .C0(R5[25]), .C1(n1014), .Y(n705) );
  AOI22XL U374 ( .A0(R7[25]), .A1(n1038), .B0(data_out_1[59]), .B1(n1022), .Y(
        n704) );
  NAND2X1 U375 ( .A(n702), .B(n703), .Y(n907) );
  AOI222X1 U376 ( .A0(R4[26]), .A1(n1010), .B0(R6[26]), .B1(n1030), .C0(R5[26]), .C1(n1014), .Y(n703) );
  AOI22XL U377 ( .A0(R7[26]), .A1(n1038), .B0(data_out_1[60]), .B1(n1022), .Y(
        n702) );
  NAND2X1 U378 ( .A(n700), .B(n701), .Y(n906) );
  AOI222X1 U379 ( .A0(R4[27]), .A1(n1010), .B0(R6[27]), .B1(n1029), .C0(R5[27]), .C1(n1014), .Y(n701) );
  AOI22XL U380 ( .A0(R7[27]), .A1(n1038), .B0(data_out_1[61]), .B1(n1019), .Y(
        n700) );
  NAND2X1 U381 ( .A(n698), .B(n699), .Y(n905) );
  AOI222X1 U382 ( .A0(R4[28]), .A1(n1010), .B0(R6[28]), .B1(n1031), .C0(R5[28]), .C1(n1014), .Y(n699) );
  AOI22XL U383 ( .A0(R7[28]), .A1(n1038), .B0(data_out_1[62]), .B1(n1021), .Y(
        n698) );
  NAND2X1 U384 ( .A(n696), .B(n697), .Y(n904) );
  AOI222X1 U385 ( .A0(R4[29]), .A1(n1010), .B0(R6[29]), .B1(n1030), .C0(R5[29]), .C1(n1014), .Y(n697) );
  AOI22XL U386 ( .A0(R7[29]), .A1(n1038), .B0(data_out_1[63]), .B1(n1018), .Y(
        n696) );
  NAND2X1 U387 ( .A(n694), .B(n695), .Y(n903) );
  AOI222X1 U388 ( .A0(R4[30]), .A1(n1010), .B0(R6[30]), .B1(n1030), .C0(R5[30]), .C1(n1016), .Y(n695) );
  AOI22XL U389 ( .A0(R7[30]), .A1(n1038), .B0(data_out_1[64]), .B1(n1023), .Y(
        n694) );
  NAND2X1 U390 ( .A(n692), .B(n693), .Y(n902) );
  AOI222X1 U391 ( .A0(R4[31]), .A1(n1009), .B0(R6[31]), .B1(n1029), .C0(R5[31]), .C1(n1014), .Y(n693) );
  AOI22XL U392 ( .A0(R7[31]), .A1(n1038), .B0(data_out_1[65]), .B1(n1022), .Y(
        n692) );
  NAND2X1 U393 ( .A(n690), .B(n691), .Y(n901) );
  AOI222X1 U394 ( .A0(R4[32]), .A1(n1009), .B0(R6[32]), .B1(n1031), .C0(R5[32]), .C1(n1016), .Y(n691) );
  AOI22XL U395 ( .A0(R7[32]), .A1(n1038), .B0(data_out_1[66]), .B1(n1025), .Y(
        n690) );
  NAND2X1 U396 ( .A(n688), .B(n689), .Y(n900) );
  AOI222X1 U397 ( .A0(R4[33]), .A1(n1009), .B0(R6[33]), .B1(n1031), .C0(R5[33]), .C1(n1015), .Y(n689) );
  AOI22XL U398 ( .A0(R7[33]), .A1(n1038), .B0(data_out_1[67]), .B1(n1020), .Y(
        n688) );
  NAND2X1 U399 ( .A(n822), .B(n823), .Y(n967) );
  AOI222X1 U400 ( .A0(R0[0]), .A1(n1009), .B0(R2[0]), .B1(n1030), .C0(R1[0]), 
        .C1(n1016), .Y(n823) );
  NAND2X1 U401 ( .A(n820), .B(n821), .Y(n966) );
  AOI222X1 U402 ( .A0(R0[1]), .A1(n1011), .B0(R2[1]), .B1(n1029), .C0(R1[1]), 
        .C1(n1016), .Y(n821) );
  NAND2X1 U403 ( .A(n818), .B(n819), .Y(n965) );
  AOI222X1 U404 ( .A0(R0[2]), .A1(n1010), .B0(R2[2]), .B1(n1031), .C0(R1[2]), 
        .C1(n1016), .Y(n819) );
  NAND2X1 U405 ( .A(n816), .B(n817), .Y(n964) );
  AOI222X1 U406 ( .A0(R0[3]), .A1(n1010), .B0(R2[3]), .B1(n1030), .C0(R1[3]), 
        .C1(n1016), .Y(n817) );
  NAND2X1 U407 ( .A(n814), .B(n815), .Y(n963) );
  AOI222X1 U408 ( .A0(R0[4]), .A1(n1011), .B0(R2[4]), .B1(n1029), .C0(R1[4]), 
        .C1(n1016), .Y(n815) );
  AOI22X1 U409 ( .A0(R3[4]), .A1(n1042), .B0(data_out_1[4]), .B1(n1018), .Y(
        n814) );
  NAND2X1 U410 ( .A(n812), .B(n813), .Y(n962) );
  AOI222X1 U411 ( .A0(R0[5]), .A1(n1010), .B0(R2[5]), .B1(n1029), .C0(R1[5]), 
        .C1(n1016), .Y(n813) );
  AOI22X1 U412 ( .A0(R3[5]), .A1(n1042), .B0(data_out_1[5]), .B1(n1018), .Y(
        n812) );
  NAND2X1 U413 ( .A(n810), .B(n811), .Y(n961) );
  AOI222X1 U414 ( .A0(R0[6]), .A1(n1009), .B0(R2[6]), .B1(n1030), .C0(R1[6]), 
        .C1(n1016), .Y(n811) );
  AOI22X1 U415 ( .A0(R3[6]), .A1(n1042), .B0(data_out_1[6]), .B1(n1018), .Y(
        n810) );
  NAND2X1 U416 ( .A(n808), .B(n809), .Y(n960) );
  AOI222X1 U417 ( .A0(R0[7]), .A1(n1010), .B0(R2[7]), .B1(n1029), .C0(R1[7]), 
        .C1(n1016), .Y(n809) );
  AOI22X1 U418 ( .A0(R3[7]), .A1(n1041), .B0(data_out_1[7]), .B1(n1018), .Y(
        n808) );
  NAND2X1 U419 ( .A(n806), .B(n807), .Y(n959) );
  AOI222X1 U420 ( .A0(R0[8]), .A1(n1011), .B0(R2[8]), .B1(n1030), .C0(R1[8]), 
        .C1(n1016), .Y(n807) );
  AOI22X1 U421 ( .A0(R3[8]), .A1(n1041), .B0(data_out_1[8]), .B1(n1018), .Y(
        n806) );
  NAND2X1 U422 ( .A(n804), .B(n805), .Y(n958) );
  AOI222X1 U423 ( .A0(R0[9]), .A1(n1010), .B0(R2[9]), .B1(n1029), .C0(R1[9]), 
        .C1(n1016), .Y(n805) );
  AOI22X1 U424 ( .A0(R3[9]), .A1(n1041), .B0(data_out_1[9]), .B1(n1018), .Y(
        n804) );
  NAND2X1 U425 ( .A(n802), .B(n803), .Y(n957) );
  AOI222X1 U426 ( .A0(R0[10]), .A1(n1010), .B0(R2[10]), .B1(n1030), .C0(R1[10]), .C1(n1016), .Y(n803) );
  AOI22X1 U427 ( .A0(R3[10]), .A1(n1041), .B0(data_out_1[10]), .B1(n1018), .Y(
        n802) );
  NAND2X1 U428 ( .A(n800), .B(n801), .Y(n956) );
  AOI222X1 U429 ( .A0(R0[11]), .A1(n1011), .B0(R2[11]), .B1(n1030), .C0(R1[11]), .C1(n1015), .Y(n801) );
  AOI22X1 U430 ( .A0(R3[11]), .A1(n1041), .B0(data_out_1[11]), .B1(n1018), .Y(
        n800) );
  NAND2X1 U431 ( .A(n798), .B(n799), .Y(n955) );
  AOI222X1 U432 ( .A0(R0[12]), .A1(n1011), .B0(R2[12]), .B1(n1030), .C0(R1[12]), .C1(n1016), .Y(n799) );
  AOI22X1 U433 ( .A0(R3[12]), .A1(n1041), .B0(data_out_1[12]), .B1(n1019), .Y(
        n798) );
  NAND2X1 U434 ( .A(n796), .B(n797), .Y(n954) );
  AOI222X1 U435 ( .A0(R0[13]), .A1(n1011), .B0(R2[13]), .B1(n1030), .C0(R1[13]), .C1(n1015), .Y(n797) );
  AOI22X1 U436 ( .A0(R3[13]), .A1(n1041), .B0(data_out_1[13]), .B1(n1019), .Y(
        n796) );
  NAND2X1 U437 ( .A(n794), .B(n795), .Y(n953) );
  AOI222X1 U438 ( .A0(R0[14]), .A1(n1011), .B0(R2[14]), .B1(n1030), .C0(R1[14]), .C1(n1016), .Y(n795) );
  AOI22X1 U439 ( .A0(R3[14]), .A1(n1041), .B0(data_out_1[14]), .B1(n1019), .Y(
        n794) );
  NAND2X1 U440 ( .A(n792), .B(n793), .Y(n952) );
  AOI222X1 U441 ( .A0(R0[15]), .A1(n1011), .B0(R2[15]), .B1(n1030), .C0(R1[15]), .C1(n1014), .Y(n793) );
  AOI22X1 U442 ( .A0(R3[15]), .A1(n1041), .B0(data_out_1[15]), .B1(n1019), .Y(
        n792) );
  NAND2X1 U443 ( .A(n790), .B(n791), .Y(n951) );
  AOI222X1 U444 ( .A0(R0[16]), .A1(n1011), .B0(R2[16]), .B1(n1030), .C0(R1[16]), .C1(n1016), .Y(n791) );
  AOI22X1 U445 ( .A0(R3[16]), .A1(n1041), .B0(data_out_1[16]), .B1(n1019), .Y(
        n790) );
  NAND2X1 U446 ( .A(n788), .B(n789), .Y(n950) );
  AOI222X1 U447 ( .A0(R0[17]), .A1(n1011), .B0(R2[17]), .B1(n1030), .C0(R1[17]), .C1(n1016), .Y(n789) );
  NAND2X1 U448 ( .A(n786), .B(n787), .Y(n949) );
  AOI222X1 U449 ( .A0(R0[18]), .A1(n1011), .B0(R2[18]), .B1(n1030), .C0(R1[18]), .C1(n1015), .Y(n787) );
  NAND2X1 U450 ( .A(n784), .B(n785), .Y(n948) );
  AOI222X1 U451 ( .A0(R0[19]), .A1(n1011), .B0(R2[19]), .B1(n1030), .C0(R1[19]), .C1(n1014), .Y(n785) );
  NAND2X1 U452 ( .A(n782), .B(n783), .Y(n947) );
  AOI222X1 U453 ( .A0(R0[20]), .A1(n1011), .B0(R2[20]), .B1(n1030), .C0(R1[20]), .C1(n1015), .Y(n783) );
  NAND2X1 U454 ( .A(n780), .B(n781), .Y(n946) );
  AOI222X1 U455 ( .A0(R0[21]), .A1(n1011), .B0(R2[21]), .B1(n1030), .C0(R1[21]), .C1(n1015), .Y(n781) );
  AOI22X1 U456 ( .A0(R3[21]), .A1(n1038), .B0(data_out_1[21]), .B1(n1019), .Y(
        n780) );
  NAND2X1 U457 ( .A(n778), .B(n779), .Y(n945) );
  AOI222X1 U458 ( .A0(R0[22]), .A1(n1011), .B0(R2[22]), .B1(n1030), .C0(R1[22]), .C1(n1015), .Y(n779) );
  AOI22X1 U459 ( .A0(R3[22]), .A1(n1034), .B0(data_out_1[22]), .B1(n1019), .Y(
        n778) );
  NAND2X1 U460 ( .A(n776), .B(n777), .Y(n944) );
  AOI222X1 U461 ( .A0(R0[23]), .A1(n1011), .B0(R2[23]), .B1(n1030), .C0(R1[23]), .C1(n1015), .Y(n777) );
  AOI22X1 U462 ( .A0(R3[23]), .A1(n1035), .B0(data_out_1[23]), .B1(n1019), .Y(
        n776) );
  NAND2X1 U463 ( .A(n774), .B(n775), .Y(n943) );
  AOI222X1 U464 ( .A0(R0[24]), .A1(n1011), .B0(R2[24]), .B1(n1030), .C0(R1[24]), .C1(n1016), .Y(n775) );
  AOI22X1 U465 ( .A0(R3[24]), .A1(n1040), .B0(data_out_1[24]), .B1(n1020), .Y(
        n774) );
  NAND2X1 U466 ( .A(n772), .B(n773), .Y(n942) );
  AOI222X1 U467 ( .A0(R0[25]), .A1(n1011), .B0(R2[25]), .B1(n1030), .C0(R1[25]), .C1(n1015), .Y(n773) );
  AOI22X1 U468 ( .A0(R3[25]), .A1(n1041), .B0(data_out_1[25]), .B1(n1020), .Y(
        n772) );
  NAND2X1 U469 ( .A(n770), .B(n771), .Y(n941) );
  AOI222X1 U470 ( .A0(R0[26]), .A1(n1011), .B0(R2[26]), .B1(n1030), .C0(R1[26]), .C1(n1016), .Y(n771) );
  AOI22X1 U471 ( .A0(R3[26]), .A1(n1037), .B0(data_out_1[26]), .B1(n1020), .Y(
        n770) );
  NAND2X1 U472 ( .A(n768), .B(n769), .Y(n940) );
  AOI222X1 U473 ( .A0(R0[27]), .A1(n1011), .B0(R2[27]), .B1(n1030), .C0(R1[27]), .C1(n1016), .Y(n769) );
  AOI22X1 U474 ( .A0(R3[27]), .A1(n1036), .B0(data_out_1[27]), .B1(n1020), .Y(
        n768) );
  NAND2X1 U475 ( .A(n766), .B(n767), .Y(n939) );
  AOI222X1 U476 ( .A0(R0[28]), .A1(n1011), .B0(R2[28]), .B1(n1030), .C0(R1[28]), .C1(n1016), .Y(n767) );
  AOI22X1 U477 ( .A0(R3[28]), .A1(n1039), .B0(data_out_1[28]), .B1(n1020), .Y(
        n766) );
  NAND2X1 U478 ( .A(n764), .B(n765), .Y(n938) );
  AOI222X1 U479 ( .A0(R0[29]), .A1(n1011), .B0(R2[29]), .B1(n1029), .C0(R1[29]), .C1(n1015), .Y(n765) );
  AOI22X1 U480 ( .A0(R3[29]), .A1(n1038), .B0(data_out_1[29]), .B1(n1020), .Y(
        n764) );
  NAND2X1 U481 ( .A(n762), .B(n763), .Y(n937) );
  AOI222X1 U482 ( .A0(R0[30]), .A1(n1011), .B0(R2[30]), .B1(n1031), .C0(R1[30]), .C1(n1015), .Y(n763) );
  AOI22X1 U483 ( .A0(R3[30]), .A1(n1037), .B0(data_out_1[30]), .B1(n1020), .Y(
        n762) );
  NAND2X1 U484 ( .A(n760), .B(n761), .Y(n936) );
  AOI222X1 U485 ( .A0(R0[31]), .A1(n1009), .B0(R2[31]), .B1(n1029), .C0(R1[31]), .C1(n1015), .Y(n761) );
  AOI22X1 U486 ( .A0(R3[31]), .A1(n1036), .B0(data_out_1[31]), .B1(n1020), .Y(
        n760) );
  NAND2X1 U487 ( .A(n758), .B(n759), .Y(n935) );
  AOI222X1 U488 ( .A0(R0[32]), .A1(n1010), .B0(R2[32]), .B1(n1030), .C0(R1[32]), .C1(n1015), .Y(n759) );
  AOI22X1 U489 ( .A0(R3[32]), .A1(n1039), .B0(data_out_1[32]), .B1(n1020), .Y(
        n758) );
  NAND2X1 U490 ( .A(n756), .B(n757), .Y(n934) );
  AOI222X1 U491 ( .A0(R0[33]), .A1(n1011), .B0(R2[33]), .B1(n1030), .C0(R1[33]), .C1(n1015), .Y(n757) );
  AOI22X1 U492 ( .A0(R3[33]), .A1(n1040), .B0(data_out_1[33]), .B1(n1020), .Y(
        n756) );
  NAND2X1 U493 ( .A(n558), .B(n559), .Y(n835) );
  AOI222X1 U494 ( .A0(R12[30]), .A1(n1008), .B0(R14[30]), .B1(n1028), .C0(
        R13[30]), .C1(n1013), .Y(n559) );
  AOI22XL U495 ( .A0(R15[30]), .A1(n1033), .B0(data_out_1[132]), .B1(n1020), 
        .Y(n558) );
  NAND2X1 U496 ( .A(n556), .B(n557), .Y(n834) );
  AOI222X1 U497 ( .A0(R12[31]), .A1(n1008), .B0(R14[31]), .B1(n1028), .C0(
        R13[31]), .C1(n1013), .Y(n557) );
  NAND2X1 U498 ( .A(n554), .B(n555), .Y(n833) );
  AOI222X1 U499 ( .A0(R12[32]), .A1(n1008), .B0(R14[32]), .B1(n1028), .C0(
        R13[32]), .C1(n1013), .Y(n555) );
  NAND2X1 U500 ( .A(n551), .B(n552), .Y(n832) );
  AOI222X1 U501 ( .A0(R12[33]), .A1(n1010), .B0(R14[33]), .B1(n1029), .C0(
        R13[33]), .C1(n1014), .Y(n552) );
  AOI22XL U502 ( .A0(R15[33]), .A1(n1039), .B0(data_out_1[135]), .B1(n1027), 
        .Y(n551) );
  NAND2X1 U503 ( .A(counter[3]), .B(n1044), .Y(n827) );
  NAND2X1 U504 ( .A(counter[2]), .B(n1045), .Y(n829) );
  NOR2X1 U505 ( .A(n550), .B(n1043), .Y(n831) );
  OAI22X1 U506 ( .A0(n831), .A1(n1044), .B0(counter[2]), .B1(n826), .Y(N14) );
endmodule


module mux ( mux_flag, clk, rst_n, data_in_1, data_in_2, data_out, 
        data_in_3_33_, data_in_3_32_, data_in_3_31_, data_in_3_30_, 
        data_in_3_29_, data_in_3_28_, data_in_3_27_, data_in_3_26_, 
        data_in_3_25_, data_in_3_24_, data_in_3_23_, data_in_3_22_, 
        data_in_3_21_, data_in_3_20_, data_in_3_19_, data_in_3_18_, 
        data_in_3_17_, data_in_3_16_, data_in_3_15_, data_in_3_14_, 
        data_in_3_13_, data_in_3_12_, data_in_3_11_, data_in_3_10_, 
        data_in_3_9_, data_in_3_8_, data_in_3_7_, data_in_3_6_, data_in_3_5_, 
        data_in_3_4_, data_in_3_3_, data_in_3_2_, data_in_3_1_, data_in_3_0_
 );
  input [135:0] data_in_1;
  input [135:0] data_in_2;
  output [135:0] data_out;
  input mux_flag, clk, rst_n, data_in_3_33_, data_in_3_32_, data_in_3_31_,
         data_in_3_30_, data_in_3_29_, data_in_3_28_, data_in_3_27_,
         data_in_3_26_, data_in_3_25_, data_in_3_24_, data_in_3_23_,
         data_in_3_22_, data_in_3_21_, data_in_3_20_, data_in_3_19_,
         data_in_3_18_, data_in_3_17_, data_in_3_16_, data_in_3_15_,
         data_in_3_14_, data_in_3_13_, data_in_3_12_, data_in_3_11_,
         data_in_3_10_, data_in_3_9_, data_in_3_8_, data_in_3_7_, data_in_3_6_,
         data_in_3_5_, data_in_3_4_, data_in_3_3_, data_in_3_2_, data_in_3_1_,
         data_in_3_0_;
  wire   n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, N6, N7, N8, n140, n141, n281, n282, n285, n2, n3,
         n4, n5, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n51, n52, n53, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n211, n212,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n283, n284, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604;
  wire   [3:1] counter;
  wire   [32:0] R4;
  wire   [32:0] R3;
  wire   [32:0] R2;
  wire   [33:0] R1;

  JKFFRX4 counter_reg_0_ ( .J(1'b1), .K(1'b1), .CK(clk), .RN(rst_n), .Q(n35), 
        .QN(n140) );
  DFFRHQX4 counter_reg_1_ ( .D(N6), .CK(clk), .RN(rst_n), .Q(counter[1]) );
  DFFRHQX4 counter_reg_2_ ( .D(N7), .CK(clk), .RN(rst_n), .Q(counter[2]) );
  DFFRHQX4 counter_reg_3_ ( .D(N8), .CK(clk), .RN(rst_n), .Q(counter[3]) );
  TLATXL R3_reg_33_ ( .G(n253), .D(data_in_3_33_), .QN(n70) );
  TLATXL R1_reg_10_ ( .G(n251), .D(data_in_3_10_), .Q(R1[10]) );
  TLATXL R1_reg_9_ ( .G(n251), .D(data_in_3_9_), .Q(R1[9]) );
  TLATXL R1_reg_7_ ( .G(n251), .D(data_in_3_7_), .Q(R1[7]) );
  TLATXL R1_reg_4_ ( .G(n251), .D(data_in_3_4_), .Q(R1[4]) );
  TLATXL R1_reg_3_ ( .G(n251), .D(data_in_3_3_), .Q(R1[3]) );
  TLATXL R1_reg_1_ ( .G(n251), .D(data_in_3_1_), .Q(R1[1]) );
  TLATXL R4_reg_1_ ( .G(n254), .D(data_in_3_1_), .Q(R4[1]) );
  TLATXL R2_reg_16_ ( .G(n5), .D(data_in_3_16_), .Q(R2[16]) );
  TLATXL R2_reg_18_ ( .G(n5), .D(data_in_3_18_), .Q(R2[18]) );
  TLATXL R2_reg_33_ ( .G(n5), .D(data_in_3_33_), .QN(n9) );
  TLATXL R4_reg_16_ ( .G(n254), .D(data_in_3_16_), .Q(R4[16]) );
  TLATXL R1_reg_29_ ( .G(n251), .D(data_in_3_29_), .Q(R1[29]) );
  TLATXL R2_reg_32_ ( .G(n5), .D(data_in_3_32_), .Q(R2[32]) );
  TLATXL R2_reg_31_ ( .G(n5), .D(data_in_3_31_), .Q(R2[31]) );
  TLATXL R2_reg_30_ ( .G(n5), .D(data_in_3_30_), .Q(R2[30]) );
  TLATXL R2_reg_29_ ( .G(n5), .D(data_in_3_29_), .Q(R2[29]) );
  TLATXL R2_reg_28_ ( .G(n5), .D(data_in_3_28_), .Q(R2[28]) );
  TLATXL R2_reg_27_ ( .G(n5), .D(data_in_3_27_), .Q(R2[27]) );
  TLATXL R2_reg_26_ ( .G(n5), .D(data_in_3_26_), .Q(R2[26]) );
  TLATXL R2_reg_25_ ( .G(n5), .D(data_in_3_25_), .Q(R2[25]) );
  TLATXL R2_reg_24_ ( .G(n5), .D(data_in_3_24_), .Q(R2[24]) );
  TLATXL R3_reg_9_ ( .G(n253), .D(data_in_3_9_), .Q(R3[9]) );
  TLATXL R3_reg_8_ ( .G(n253), .D(data_in_3_8_), .Q(R3[8]) );
  TLATXL R3_reg_7_ ( .G(n253), .D(data_in_3_7_), .Q(R3[7]) );
  TLATXL R3_reg_6_ ( .G(n253), .D(data_in_3_6_), .Q(R3[6]) );
  TLATXL R3_reg_5_ ( .G(n253), .D(data_in_3_5_), .Q(R3[5]) );
  TLATXL R3_reg_4_ ( .G(n253), .D(data_in_3_4_), .Q(R3[4]) );
  TLATXL R3_reg_3_ ( .G(n253), .D(data_in_3_3_), .Q(R3[3]) );
  TLATXL R3_reg_2_ ( .G(n253), .D(data_in_3_2_), .Q(R3[2]) );
  TLATXL R4_reg_9_ ( .G(n254), .D(data_in_3_9_), .Q(R4[9]) );
  TLATXL R4_reg_8_ ( .G(n254), .D(data_in_3_8_), .Q(R4[8]) );
  TLATXL R4_reg_7_ ( .G(n254), .D(data_in_3_7_), .Q(R4[7]) );
  TLATXL R4_reg_6_ ( .G(n254), .D(data_in_3_6_), .Q(R4[6]) );
  TLATXL R4_reg_5_ ( .G(n254), .D(data_in_3_5_), .Q(R4[5]) );
  TLATXL R4_reg_4_ ( .G(n254), .D(data_in_3_4_), .Q(R4[4]) );
  TLATXL R4_reg_3_ ( .G(n254), .D(data_in_3_3_), .Q(R4[3]) );
  TLATXL R4_reg_2_ ( .G(n254), .D(data_in_3_2_), .Q(R4[2]) );
  TLATXL R1_reg_12_ ( .G(n251), .D(data_in_3_12_), .Q(R1[12]) );
  TLATXL R2_reg_23_ ( .G(n5), .D(data_in_3_23_), .Q(R2[23]) );
  TLATXL R2_reg_22_ ( .G(n5), .D(data_in_3_22_), .Q(R2[22]) );
  TLATXL R2_reg_21_ ( .G(n5), .D(data_in_3_21_), .Q(R2[21]) );
  TLATXL R2_reg_20_ ( .G(n5), .D(data_in_3_20_), .Q(R2[20]) );
  TLATXL R2_reg_19_ ( .G(n5), .D(data_in_3_19_), .Q(R2[19]) );
  TLATXL R2_reg_15_ ( .G(n5), .D(data_in_3_15_), .Q(R2[15]) );
  TLATXL R2_reg_14_ ( .G(n5), .D(data_in_3_14_), .Q(R2[14]) );
  TLATXL R2_reg_13_ ( .G(n5), .D(data_in_3_13_), .Q(R2[13]) );
  TLATXL R2_reg_12_ ( .G(n5), .D(data_in_3_12_), .Q(R2[12]) );
  TLATXL R2_reg_11_ ( .G(n5), .D(data_in_3_11_), .Q(R2[11]) );
  TLATXL R2_reg_10_ ( .G(n5), .D(data_in_3_10_), .Q(R2[10]) );
  TLATXL R2_reg_9_ ( .G(n5), .D(data_in_3_9_), .Q(R2[9]) );
  TLATXL R2_reg_8_ ( .G(n5), .D(data_in_3_8_), .Q(R2[8]) );
  TLATXL R2_reg_7_ ( .G(n5), .D(data_in_3_7_), .Q(R2[7]) );
  TLATXL R2_reg_6_ ( .G(n5), .D(data_in_3_6_), .Q(R2[6]) );
  TLATXL R2_reg_5_ ( .G(n5), .D(data_in_3_5_), .Q(R2[5]) );
  TLATXL R2_reg_4_ ( .G(n5), .D(data_in_3_4_), .Q(R2[4]) );
  TLATXL R2_reg_3_ ( .G(n5), .D(data_in_3_3_), .Q(R2[3]) );
  TLATXL R3_reg_32_ ( .G(n253), .D(data_in_3_32_), .Q(R3[32]) );
  TLATXL R3_reg_31_ ( .G(n253), .D(data_in_3_31_), .Q(R3[31]) );
  TLATXL R3_reg_30_ ( .G(n253), .D(data_in_3_30_), .Q(R3[30]) );
  TLATXL R3_reg_29_ ( .G(n253), .D(data_in_3_29_), .Q(R3[29]) );
  TLATXL R3_reg_28_ ( .G(n253), .D(data_in_3_28_), .Q(R3[28]) );
  TLATXL R3_reg_27_ ( .G(n253), .D(data_in_3_27_), .Q(R3[27]) );
  TLATXL R3_reg_26_ ( .G(n253), .D(data_in_3_26_), .Q(R3[26]) );
  TLATXL R3_reg_25_ ( .G(n253), .D(data_in_3_25_), .Q(R3[25]) );
  TLATXL R3_reg_24_ ( .G(n253), .D(data_in_3_24_), .Q(R3[24]) );
  TLATXL R3_reg_23_ ( .G(n253), .D(data_in_3_23_), .Q(R3[23]) );
  TLATXL R3_reg_22_ ( .G(n253), .D(data_in_3_22_), .Q(R3[22]) );
  TLATXL R3_reg_21_ ( .G(n253), .D(data_in_3_21_), .Q(R3[21]) );
  TLATXL R3_reg_20_ ( .G(n253), .D(data_in_3_20_), .Q(R3[20]) );
  TLATXL R3_reg_19_ ( .G(n253), .D(data_in_3_19_), .Q(R3[19]) );
  TLATXL R3_reg_16_ ( .G(n253), .D(data_in_3_16_), .Q(R3[16]) );
  TLATXL R3_reg_15_ ( .G(n253), .D(data_in_3_15_), .Q(R3[15]) );
  TLATXL R3_reg_14_ ( .G(n253), .D(data_in_3_14_), .Q(R3[14]) );
  TLATXL R3_reg_13_ ( .G(n253), .D(data_in_3_13_), .Q(R3[13]) );
  TLATXL R3_reg_12_ ( .G(n253), .D(data_in_3_12_), .Q(R3[12]) );
  TLATXL R3_reg_11_ ( .G(n253), .D(data_in_3_11_), .Q(R3[11]) );
  TLATXL R3_reg_10_ ( .G(n253), .D(data_in_3_10_), .Q(R3[10]) );
  TLATXL R4_reg_33_ ( .G(n254), .D(data_in_3_33_), .QN(n10) );
  TLATXL R4_reg_32_ ( .G(n254), .D(data_in_3_32_), .Q(R4[32]) );
  TLATXL R4_reg_31_ ( .G(n254), .D(data_in_3_31_), .Q(R4[31]) );
  TLATXL R4_reg_30_ ( .G(n254), .D(data_in_3_30_), .Q(R4[30]) );
  TLATXL R4_reg_29_ ( .G(n254), .D(data_in_3_29_), .Q(R4[29]) );
  TLATXL R4_reg_28_ ( .G(n254), .D(data_in_3_28_), .Q(R4[28]) );
  TLATXL R4_reg_27_ ( .G(n254), .D(data_in_3_27_), .Q(R4[27]) );
  TLATXL R4_reg_26_ ( .G(n254), .D(data_in_3_26_), .Q(R4[26]) );
  TLATXL R4_reg_25_ ( .G(n254), .D(data_in_3_25_), .Q(R4[25]) );
  TLATXL R4_reg_24_ ( .G(n254), .D(data_in_3_24_), .Q(R4[24]) );
  TLATXL R4_reg_23_ ( .G(n254), .D(data_in_3_23_), .Q(R4[23]) );
  TLATXL R4_reg_22_ ( .G(n254), .D(data_in_3_22_), .Q(R4[22]) );
  TLATXL R4_reg_21_ ( .G(n254), .D(data_in_3_21_), .Q(R4[21]) );
  TLATXL R4_reg_20_ ( .G(n254), .D(data_in_3_20_), .Q(R4[20]) );
  TLATXL R4_reg_19_ ( .G(n254), .D(data_in_3_19_), .Q(R4[19]) );
  TLATXL R4_reg_15_ ( .G(n254), .D(data_in_3_15_), .Q(R4[15]) );
  TLATXL R4_reg_14_ ( .G(n254), .D(data_in_3_14_), .Q(R4[14]) );
  TLATXL R4_reg_13_ ( .G(n254), .D(data_in_3_13_), .Q(R4[13]) );
  TLATXL R4_reg_12_ ( .G(n254), .D(data_in_3_12_), .Q(R4[12]) );
  TLATXL R4_reg_11_ ( .G(n254), .D(data_in_3_11_), .Q(R4[11]) );
  TLATXL R4_reg_10_ ( .G(n254), .D(data_in_3_10_), .Q(R4[10]) );
  TLATXL R3_reg_1_ ( .G(n253), .D(data_in_3_1_), .Q(R3[1]) );
  TLATXL R2_reg_1_ ( .G(n5), .D(data_in_3_1_), .Q(R2[1]) );
  TLATXL R3_reg_18_ ( .G(n253), .D(data_in_3_18_), .Q(R3[18]) );
  TLATXL R4_reg_18_ ( .G(n254), .D(data_in_3_18_), .Q(R4[18]) );
  TLATXL R1_reg_33_ ( .G(n251), .D(data_in_3_33_), .Q(R1[33]) );
  TLATXL R1_reg_32_ ( .G(n251), .D(data_in_3_32_), .Q(R1[32]) );
  TLATXL R1_reg_31_ ( .G(n251), .D(data_in_3_31_), .Q(R1[31]) );
  TLATXL R1_reg_30_ ( .G(n251), .D(data_in_3_30_), .Q(R1[30]) );
  TLATXL R1_reg_28_ ( .G(n285), .D(data_in_3_28_), .Q(R1[28]) );
  TLATXL R1_reg_27_ ( .G(n285), .D(data_in_3_27_), .Q(R1[27]) );
  TLATXL R1_reg_26_ ( .G(n285), .D(data_in_3_26_), .Q(R1[26]) );
  TLATXL R1_reg_25_ ( .G(n285), .D(data_in_3_25_), .Q(R1[25]) );
  TLATXL R1_reg_24_ ( .G(n285), .D(data_in_3_24_), .Q(R1[24]) );
  TLATXL R1_reg_23_ ( .G(n251), .D(data_in_3_23_), .Q(R1[23]) );
  TLATXL R1_reg_22_ ( .G(n251), .D(data_in_3_22_), .Q(R1[22]) );
  TLATXL R1_reg_21_ ( .G(n251), .D(data_in_3_21_), .Q(R1[21]) );
  TLATXL R1_reg_20_ ( .G(n251), .D(data_in_3_20_), .Q(R1[20]) );
  TLATXL R1_reg_19_ ( .G(n251), .D(data_in_3_19_), .Q(R1[19]) );
  TLATXL R1_reg_18_ ( .G(n251), .D(data_in_3_18_), .Q(R1[18]) );
  TLATXL R1_reg_16_ ( .G(n251), .D(data_in_3_16_), .Q(R1[16]) );
  TLATXL R1_reg_15_ ( .G(n251), .D(data_in_3_15_), .Q(R1[15]) );
  TLATXL R1_reg_14_ ( .G(n251), .D(data_in_3_14_), .Q(R1[14]) );
  TLATXL R1_reg_13_ ( .G(n251), .D(data_in_3_13_), .Q(R1[13]) );
  TLATXL R1_reg_11_ ( .G(n251), .D(data_in_3_11_), .Q(R1[11]) );
  TLATXL R1_reg_8_ ( .G(n251), .D(data_in_3_8_), .Q(R1[8]) );
  TLATXL R1_reg_6_ ( .G(n251), .D(data_in_3_6_), .Q(R1[6]) );
  TLATXL R1_reg_5_ ( .G(n251), .D(data_in_3_5_), .Q(R1[5]) );
  TLATXL R1_reg_2_ ( .G(n251), .D(data_in_3_2_), .Q(R1[2]) );
  TLATXL R2_reg_2_ ( .G(n5), .D(data_in_3_2_), .Q(n21) );
  TLATXL R3_reg_0_ ( .G(n253), .D(data_in_3_0_), .Q(R3[0]) );
  TLATXL R2_reg_17_ ( .G(n5), .D(data_in_3_17_), .Q(R2[17]) );
  TLATXL R2_reg_0_ ( .G(n5), .D(data_in_3_0_), .Q(R2[0]) );
  TLATXL R4_reg_0_ ( .G(n254), .D(data_in_3_0_), .Q(R4[0]) );
  TLATXL R1_reg_17_ ( .G(n251), .D(data_in_3_17_), .Q(R1[17]) );
  TLATXL R1_reg_0_ ( .G(n251), .D(data_in_3_0_), .Q(R1[0]) );
  TLATXL R3_reg_17_ ( .G(n253), .D(data_in_3_17_), .Q(R3[17]) );
  TLATXL R4_reg_17_ ( .G(n254), .D(data_in_3_17_), .Q(R4[17]) );
  CLKBUFX20 U4 ( .A(n611), .Y(data_out[85]) );
  CLKINVX8 U5 ( .A(n20), .Y(n4) );
  NAND2BX1 U6 ( .AN(n256), .B(data_in_2[119]), .Y(n556) );
  BUFX20 U7 ( .A(n41), .Y(n2) );
  BUFX12 U8 ( .A(n612), .Y(data_out[71]) );
  NAND2X4 U9 ( .A(n43), .B(R3[16]), .Y(n453) );
  AOI2BB2X4 U10 ( .B0(n557), .B1(n30), .A0N(n4), .A1N(n556), .Y(n558) );
  NAND3X1 U11 ( .A(n257), .B(data_in_2[121]), .C(n12), .Y(n563) );
  BUFX12 U12 ( .A(n599), .Y(n12) );
  AOI2BB2X4 U13 ( .B0(n456), .B1(n23), .A0N(n455), .A1N(n4), .Y(n457) );
  INVX4 U14 ( .A(n45), .Y(n3) );
  CLKINVX8 U15 ( .A(n245), .Y(n45) );
  INVX12 U16 ( .A(n248), .Y(n246) );
  NAND2X1 U17 ( .A(data_in_1[38]), .B(n240), .Y(n317) );
  INVX4 U18 ( .A(n243), .Y(n48) );
  NAND3X2 U19 ( .A(data_in_1[70]), .B(n255), .C(n48), .Y(n413) );
  NAND2BX1 U20 ( .AN(n256), .B(data_in_2[35]), .Y(n312) );
  INVX8 U21 ( .A(n599), .Y(n22) );
  NAND2X1 U22 ( .A(data_in_2[123]), .B(n17), .Y(n571) );
  NAND2X1 U23 ( .A(R4[21]), .B(n223), .Y(n569) );
  INVX20 U24 ( .A(n249), .Y(n29) );
  NOR2X2 U25 ( .A(n37), .B(n511), .Y(n513) );
  NAND2BX2 U26 ( .AN(n10), .B(n42), .Y(n600) );
  NAND3X2 U27 ( .A(n565), .B(n564), .C(n563), .Y(n606) );
  INVX8 U28 ( .A(n2), .Y(n47) );
  CLKINVX8 U29 ( .A(n47), .Y(n32) );
  AOI2BB2X4 U30 ( .B0(n43), .B1(R4[18]), .A0N(n247), .A1N(n559), .Y(n560) );
  AOI2BB2X4 U31 ( .B0(n310), .B1(n30), .A0N(n22), .A1N(n309), .Y(n311) );
  OR2X4 U32 ( .A(n66), .B(n212), .Y(n20) );
  OR3X4 U33 ( .A(n31), .B(n66), .C(n70), .Y(n504) );
  INVX12 U34 ( .A(n300), .Y(n594) );
  BUFX20 U35 ( .A(n300), .Y(n11) );
  INVX20 U36 ( .A(n11), .Y(n241) );
  INVX2 U37 ( .A(n222), .Y(n17) );
  BUFX20 U38 ( .A(n303), .Y(n222) );
  INVX12 U39 ( .A(n235), .Y(n231) );
  CLKINVX8 U40 ( .A(n236), .Y(n298) );
  CLKINVX3 U41 ( .A(n252), .Y(n251) );
  NOR3X4 U42 ( .A(n282), .B(n603), .C(n604), .Y(n5) );
  CLKINVX3 U43 ( .A(n8), .Y(n254) );
  CLKINVX3 U44 ( .A(n7), .Y(n253) );
  BUFX20 U45 ( .A(n616), .Y(data_out[35]) );
  NAND2XL U46 ( .A(R2[7]), .B(n32), .Y(n325) );
  NAND2XL U47 ( .A(R3[20]), .B(n41), .Y(n463) );
  NAND3BX4 U48 ( .AN(n256), .B(data_in_2[101]), .C(n52), .Y(n502) );
  NAND3X1 U49 ( .A(data_in_1[87]), .B(n255), .C(n28), .Y(n462) );
  AND2X2 U50 ( .A(n28), .B(n512), .Y(n68) );
  BUFX20 U51 ( .A(n561), .Y(n227) );
  BUFX8 U52 ( .A(n41), .Y(n37) );
  INVX3 U53 ( .A(n43), .Y(n44) );
  INVX8 U54 ( .A(n42), .Y(n28) );
  BUFX8 U55 ( .A(n606), .Y(data_out[121]) );
  NAND2X2 U56 ( .A(data_in_1[88]), .B(n240), .Y(n464) );
  INVX3 U57 ( .A(n234), .Y(n233) );
  INVX1 U58 ( .A(data_in_2[29]), .Y(n301) );
  OAI2BB1X1 U59 ( .A0N(data_in_2[11]), .A1N(n233), .B0(n272), .Y(data_out[11])
         );
  NAND2BX2 U60 ( .AN(n256), .B(data_in_2[69]), .Y(n409) );
  NAND2BX2 U61 ( .AN(n256), .B(data_in_2[120]), .Y(n559) );
  NAND2BX2 U62 ( .AN(n256), .B(data_in_2[68]), .Y(n406) );
  NAND2BX2 U63 ( .AN(n256), .B(data_in_2[52]), .Y(n358) );
  NAND2X2 U64 ( .A(data_in_2[56]), .B(n305), .Y(n372) );
  NAND2BX2 U65 ( .AN(n256), .B(data_in_2[84]), .Y(n451) );
  OR3XL U66 ( .A(n224), .B(n38), .C(n40), .Y(n141) );
  CLKINVX4 U67 ( .A(n41), .Y(n24) );
  OR2X2 U68 ( .A(n211), .B(n141), .Y(n7) );
  OR2XL U69 ( .A(n36), .B(n141), .Y(n8) );
  AND2X4 U70 ( .A(R4[2]), .B(n243), .Y(n69) );
  CLKINVX8 U71 ( .A(n593), .Y(n236) );
  CLKBUFX8 U72 ( .A(n53), .Y(n30) );
  AOI2BB2X4 U73 ( .B0(R4[0]), .B1(n19), .A0N(n4), .A1N(n505), .Y(n506) );
  NAND2BX1 U74 ( .AN(n256), .B(data_in_2[102]), .Y(n505) );
  CLKINVX3 U75 ( .A(n24), .Y(n13) );
  INVX12 U76 ( .A(n249), .Y(n223) );
  INVX12 U77 ( .A(n249), .Y(n226) );
  NAND2XL U78 ( .A(data_in_1[58]), .B(n237), .Y(n377) );
  BUFX16 U79 ( .A(n605), .Y(data_out[135]) );
  NAND3X1 U80 ( .A(n52), .B(data_in_1[121]), .C(n255), .Y(n564) );
  NAND2X4 U81 ( .A(data_in_1[55]), .B(n238), .Y(n368) );
  NAND2X4 U82 ( .A(n403), .B(n28), .Y(n404) );
  NAND2X2 U83 ( .A(data_in_1[56]), .B(n238), .Y(n371) );
  NAND2X4 U84 ( .A(data_in_2[54]), .B(n273), .Y(n366) );
  INVX8 U85 ( .A(n236), .Y(n273) );
  NAND2X1 U86 ( .A(R2[20]), .B(n2), .Y(n364) );
  NAND2X1 U87 ( .A(R4[7]), .B(n2), .Y(n526) );
  BUFX20 U88 ( .A(n613), .Y(data_out[67]) );
  INVX4 U89 ( .A(n245), .Y(n46) );
  AND2X1 U90 ( .A(data_in_1[127]), .B(n237), .Y(n78) );
  AND2X4 U91 ( .A(n502), .B(n504), .Y(n14) );
  NAND2BX4 U92 ( .AN(n15), .B(n14), .Y(data_out[101]) );
  AND3X2 U93 ( .A(n53), .B(n255), .C(data_in_1[101]), .Y(n15) );
  NAND2BX1 U94 ( .AN(n256), .B(data_in_2[34]), .Y(n309) );
  INVX8 U95 ( .A(n22), .Y(n23) );
  NOR3BX4 U96 ( .AN(data_in_2[135]), .B(n598), .C(n255), .Y(n602) );
  NAND2X2 U97 ( .A(R4[19]), .B(n2), .Y(n565) );
  NAND2X2 U98 ( .A(R4[4]), .B(n244), .Y(n517) );
  NAND2X2 U99 ( .A(R3[23]), .B(n244), .Y(n472) );
  AOI2BB2X2 U100 ( .B0(n356), .B1(n30), .A0N(n355), .A1N(n598), .Y(n357) );
  BUFX3 U101 ( .A(n618), .Y(data_out[13]) );
  AOI2BB2X4 U102 ( .B0(R2[18]), .B1(n19), .A0N(n247), .A1N(n358), .Y(n359) );
  OAI2BB1X4 U103 ( .A0N(R2[17]), .A1N(n247), .B0(n357), .Y(data_out[51]) );
  OAI2BB1X4 U104 ( .A0N(R4[17]), .A1N(n247), .B0(n558), .Y(n608) );
  OAI2BB2X4 U105 ( .B0(n28), .B1(n9), .A0N(n18), .A1N(n250), .Y(n405) );
  AND2X2 U106 ( .A(data_in_1[67]), .B(n255), .Y(n18) );
  INVX8 U107 ( .A(n12), .Y(n19) );
  NAND2X4 U108 ( .A(data_in_2[37]), .B(n273), .Y(n26) );
  AND2X2 U109 ( .A(R3[19]), .B(n2), .Y(n62) );
  NAND3X1 U110 ( .A(data_in_1[135]), .B(n255), .C(n599), .Y(n601) );
  INVX8 U111 ( .A(n235), .Y(n305) );
  CLKINVX8 U112 ( .A(n34), .Y(n250) );
  NAND3BX2 U113 ( .AN(n256), .B(data_in_2[70]), .C(n45), .Y(n412) );
  CLKINVX8 U114 ( .A(n234), .Y(n232) );
  AOI22X4 U115 ( .A0(data_in_2[36]), .A1(n230), .B0(n21), .B1(n29), .Y(n315)
         );
  NAND2X4 U116 ( .A(R3[3]), .B(n246), .Y(n415) );
  CLKINVX8 U117 ( .A(n34), .Y(n249) );
  NAND3XL U118 ( .A(n599), .B(data_in_1[53]), .C(n255), .Y(n362) );
  NAND3XL U119 ( .A(n258), .B(data_in_2[53]), .C(n599), .Y(n361) );
  NAND3X4 U120 ( .A(n26), .B(n27), .C(n25), .Y(data_out[37]) );
  CLKINVX20 U121 ( .A(n67), .Y(n25) );
  NAND2X4 U122 ( .A(data_in_1[37]), .B(n239), .Y(n27) );
  INVX8 U123 ( .A(n42), .Y(n248) );
  INVX8 U124 ( .A(n235), .Y(n280) );
  NAND2X2 U125 ( .A(data_in_2[122]), .B(n280), .Y(n568) );
  NAND2X2 U126 ( .A(data_in_2[57]), .B(n280), .Y(n375) );
  NAND2X2 U127 ( .A(data_in_2[59]), .B(n280), .Y(n381) );
  CLKINVX8 U128 ( .A(n258), .Y(n256) );
  INVX8 U129 ( .A(n11), .Y(n239) );
  NAND2X2 U130 ( .A(data_in_1[125]), .B(n239), .Y(n576) );
  NAND2X2 U131 ( .A(data_in_1[74]), .B(n239), .Y(n425) );
  NAND2X2 U132 ( .A(data_in_1[41]), .B(n239), .Y(n326) );
  NAND2X2 U133 ( .A(data_in_1[95]), .B(n239), .Y(n485) );
  INVX8 U134 ( .A(n227), .Y(n42) );
  NAND2XL U135 ( .A(R2[14]), .B(n37), .Y(n346) );
  NAND2XL U136 ( .A(R2[29]), .B(n37), .Y(n391) );
  NAND2XL U137 ( .A(R3[9]), .B(n37), .Y(n433) );
  INVXL U138 ( .A(n36), .Y(n31) );
  NAND2XL U139 ( .A(R3[4]), .B(n37), .Y(n418) );
  AND2X1 U140 ( .A(R4[25]), .B(n37), .Y(n79) );
  AOI2BB2X4 U141 ( .B0(n407), .B1(n23), .A0N(n43), .A1N(n406), .Y(n408) );
  BUFX20 U142 ( .A(n615), .Y(data_out[36]) );
  NAND2XL U143 ( .A(R3[13]), .B(n226), .Y(n445) );
  NAND2XL U144 ( .A(R3[28]), .B(n226), .Y(n487) );
  NAND2XL U145 ( .A(R2[25]), .B(n226), .Y(n379) );
  NAND2XL U146 ( .A(R3[6]), .B(n29), .Y(n424) );
  NAND2XL U147 ( .A(R4[20]), .B(n226), .Y(n566) );
  DLY1X1 U148 ( .A(counter[1]), .Y(n224) );
  NAND2X2 U149 ( .A(data_in_2[38]), .B(n296), .Y(n318) );
  NOR2X2 U150 ( .A(n503), .B(n35), .Y(n225) );
  NAND2X2 U151 ( .A(data_in_1[72]), .B(n237), .Y(n419) );
  NAND2XL U152 ( .A(R2[30]), .B(n37), .Y(n394) );
  NAND2X2 U153 ( .A(data_in_1[89]), .B(n241), .Y(n467) );
  NAND2XL U154 ( .A(data_in_1[54]), .B(n594), .Y(n365) );
  NAND2X2 U155 ( .A(R3[12]), .B(n29), .Y(n442) );
  NAND2X2 U156 ( .A(R3[14]), .B(n29), .Y(n448) );
  NAND2X2 U157 ( .A(R2[19]), .B(n243), .Y(n363) );
  INVX8 U158 ( .A(n11), .Y(n238) );
  BUFX20 U159 ( .A(n617), .Y(data_out[34]) );
  BUFX20 U160 ( .A(n607), .Y(data_out[120]) );
  AOI2BB2X2 U161 ( .B0(R2[1]), .B1(n41), .A0N(n598), .A1N(n312), .Y(n313) );
  NAND3X2 U162 ( .A(n540), .B(n539), .C(n538), .Y(data_out[113]) );
  OAI2BB1X1 U163 ( .A0N(data_in_2[28]), .A1N(n280), .B0(n297), .Y(data_out[28]) );
  NAND3X2 U164 ( .A(n396), .B(n395), .C(n394), .Y(data_out[64]) );
  OAI22X4 U165 ( .A0(n452), .A1(n598), .B0(n22), .B1(n451), .Y(n454) );
  INVX8 U166 ( .A(n71), .Y(data_out[88]) );
  CLKINVX8 U167 ( .A(n236), .Y(n228) );
  CLKINVX8 U168 ( .A(n593), .Y(n234) );
  INVX8 U169 ( .A(n227), .Y(n41) );
  BUFX20 U170 ( .A(n609), .Y(data_out[104]) );
  NAND2X2 U171 ( .A(R3[2]), .B(n2), .Y(n414) );
  NAND2X2 U172 ( .A(data_in_1[106]), .B(n240), .Y(n518) );
  INVX8 U173 ( .A(n11), .Y(n240) );
  OAI2BB1X4 U174 ( .A0N(n314), .A1N(n46), .B0(n313), .Y(n616) );
  BUFX20 U175 ( .A(n610), .Y(data_out[86]) );
  AOI2BB2X4 U176 ( .B0(R3[1]), .B1(n243), .A0N(n247), .A1N(n409), .Y(n410) );
  NAND2XL U177 ( .A(data_in_2[96]), .B(n231), .Y(n489) );
  NAND2XL U178 ( .A(data_in_2[94]), .B(n17), .Y(n483) );
  NAND2XL U179 ( .A(data_in_2[92]), .B(n231), .Y(n477) );
  NAND2X4 U180 ( .A(data_in_1[123]), .B(n237), .Y(n570) );
  INVX8 U181 ( .A(n11), .Y(n237) );
  AOI2BB2X4 U182 ( .B0(R3[18]), .B1(n245), .A0N(n247), .A1N(n458), .Y(n459) );
  NAND2X4 U183 ( .A(data_in_1[73]), .B(n240), .Y(n422) );
  OR2X4 U184 ( .A(n212), .B(n66), .Y(n49) );
  OAI2BB1X4 U185 ( .A0N(R3[0]), .A1N(n247), .B0(n408), .Y(data_out[68]) );
  NAND2X2 U186 ( .A(R2[21]), .B(n29), .Y(n367) );
  NAND2X2 U187 ( .A(R4[24]), .B(n226), .Y(n578) );
  NAND2X2 U188 ( .A(R2[27]), .B(n29), .Y(n385) );
  INVX8 U189 ( .A(n593), .Y(n235) );
  OAI2BB1X4 U190 ( .A0N(data_in_1[36]), .A1N(n594), .B0(n315), .Y(n615) );
  INVX8 U191 ( .A(n227), .Y(n34) );
  AOI22XL U192 ( .A0(data_in_1[18]), .A1(n241), .B0(R1[18]), .B1(n226), .Y(
        n286) );
  OAI2BB1X4 U193 ( .A0N(n460), .A1N(n44), .B0(n459), .Y(n610) );
  INVX8 U194 ( .A(n212), .Y(n36) );
  CLKINVX8 U195 ( .A(n260), .Y(n66) );
  DLY1X1 U196 ( .A(counter[2]), .Y(n38) );
  NAND3X4 U197 ( .A(n363), .B(n362), .C(n361), .Y(data_out[53]) );
  INVX8 U198 ( .A(mux_flag), .Y(n258) );
  NAND2BX1 U199 ( .AN(n256), .B(data_in_2[103]), .Y(n508) );
  CLKINVX20 U200 ( .A(n258), .Y(n255) );
  NOR2BX2 U201 ( .AN(data_in_2[67]), .B(n255), .Y(n403) );
  XOR2XL U202 ( .A(n224), .B(n211), .Y(N6) );
  NAND2X4 U203 ( .A(n39), .B(n555), .Y(data_out[118]) );
  AND2X4 U204 ( .A(n553), .B(n554), .Y(n39) );
  INVX20 U205 ( .A(n225), .Y(n599) );
  NAND3X2 U206 ( .A(n471), .B(n470), .C(n469), .Y(data_out[90]) );
  INVX1 U207 ( .A(n604), .Y(n40) );
  NAND3BX4 U208 ( .AN(n256), .B(data_in_2[87]), .C(n47), .Y(n461) );
  NAND2XL U209 ( .A(R4[3]), .B(n223), .Y(n514) );
  INVX8 U210 ( .A(n249), .Y(n243) );
  NAND2X4 U211 ( .A(n255), .B(n49), .Y(n300) );
  NAND3X4 U212 ( .A(n468), .B(n467), .C(n466), .Y(data_out[89]) );
  INVX8 U213 ( .A(n222), .Y(n230) );
  AOI2BB2X2 U214 ( .B0(n353), .B1(n23), .A0N(n352), .A1N(n598), .Y(n354) );
  NAND2BX4 U215 ( .AN(n599), .B(R4[16]), .Y(n553) );
  AOI2BB2X2 U216 ( .B0(n509), .B1(n12), .A0N(n508), .A1N(n598), .Y(n510) );
  INVX8 U217 ( .A(n503), .Y(n260) );
  NAND3X1 U218 ( .A(data_in_1[118]), .B(n255), .C(n20), .Y(n555) );
  INVX8 U219 ( .A(n248), .Y(n245) );
  BUFX20 U220 ( .A(n608), .Y(data_out[119]) );
  OR2X4 U221 ( .A(n66), .B(n212), .Y(n52) );
  INVX8 U222 ( .A(n72), .Y(data_out[54]) );
  NAND2X4 U223 ( .A(data_in_2[106]), .B(n228), .Y(n519) );
  NAND2X2 U224 ( .A(data_in_2[72]), .B(n229), .Y(n420) );
  CLKINVX8 U225 ( .A(n222), .Y(n229) );
  INVX8 U226 ( .A(n250), .Y(n43) );
  NAND2X4 U227 ( .A(n260), .B(n36), .Y(n561) );
  NAND3BX4 U228 ( .AN(n602), .B(n601), .C(n600), .Y(n605) );
  INVX8 U229 ( .A(n53), .Y(n598) );
  NAND3BX1 U230 ( .AN(n255), .B(n53), .C(data_in_2[118]), .Y(n554) );
  OR2X4 U231 ( .A(n503), .B(n212), .Y(n53) );
  INVX12 U232 ( .A(n235), .Y(n296) );
  INVX8 U233 ( .A(n222), .Y(n593) );
  NAND2X4 U234 ( .A(n49), .B(n257), .Y(n303) );
  INVXL U235 ( .A(n239), .Y(n51) );
  INVX16 U236 ( .A(n11), .Y(n242) );
  INVX8 U237 ( .A(n24), .Y(n244) );
  NAND2XL U238 ( .A(R3[21]), .B(n246), .Y(n466) );
  INVX8 U239 ( .A(n599), .Y(n247) );
  NAND3BX4 U240 ( .AN(n62), .B(n462), .C(n461), .Y(data_out[87]) );
  NAND3X4 U241 ( .A(n412), .B(n413), .C(n414), .Y(data_out[70]) );
  NAND2BX2 U242 ( .AN(n256), .B(data_in_2[86]), .Y(n458) );
  AND2X2 U243 ( .A(data_in_1[128]), .B(n237), .Y(n75) );
  NAND3BX1 U244 ( .AN(n73), .B(n63), .C(n64), .Y(data_out[129]) );
  NAND2XL U245 ( .A(data_in_1[129]), .B(n240), .Y(n63) );
  NAND2XL U246 ( .A(R4[27]), .B(n226), .Y(n64) );
  AOI22XL U247 ( .A0(data_in_1[19]), .A1(n237), .B0(R1[19]), .B1(n246), .Y(
        n287) );
  AOI22XL U248 ( .A0(data_in_1[2]), .A1(n240), .B0(R1[2]), .B1(n37), .Y(n263)
         );
  AOI22XL U249 ( .A0(data_in_1[21]), .A1(n241), .B0(R1[21]), .B1(n226), .Y(
        n289) );
  AOI22XL U250 ( .A0(data_in_1[22]), .A1(n239), .B0(R1[22]), .B1(n223), .Y(
        n290) );
  AOI22XL U251 ( .A0(data_in_1[24]), .A1(n241), .B0(R1[24]), .B1(n226), .Y(
        n292) );
  AOI22XL U252 ( .A0(data_in_1[5]), .A1(n240), .B0(R1[5]), .B1(n223), .Y(n266)
         );
  AOI22XL U253 ( .A0(data_in_1[6]), .A1(n241), .B0(R1[6]), .B1(n13), .Y(n267)
         );
  AOI22XL U254 ( .A0(data_in_1[8]), .A1(n242), .B0(R1[8]), .B1(n246), .Y(n269)
         );
  AOI22XL U255 ( .A0(data_in_1[14]), .A1(n240), .B0(R1[14]), .B1(n246), .Y(
        n278) );
  OAI2BB1X1 U256 ( .A0N(data_in_2[13]), .A1N(n296), .B0(n277), .Y(n618) );
  AOI22XL U257 ( .A0(data_in_1[11]), .A1(n241), .B0(R1[11]), .B1(n223), .Y(
        n272) );
  OR2X2 U258 ( .A(n276), .B(n65), .Y(data_out[12]) );
  AND2X1 U259 ( .A(R1[12]), .B(n13), .Y(n65) );
  AOI22XL U260 ( .A0(data_in_1[16]), .A1(n238), .B0(R1[16]), .B1(n37), .Y(n283) );
  OAI2BB1X1 U261 ( .A0N(data_in_2[15]), .A1N(n305), .B0(n279), .Y(data_out[15]) );
  AOI22XL U262 ( .A0(data_in_1[15]), .A1(n241), .B0(R1[15]), .B1(n29), .Y(n279) );
  INVX1 U263 ( .A(n285), .Y(n252) );
  INVXL U264 ( .A(mux_flag), .Y(n257) );
  XOR2X1 U265 ( .A(n603), .B(n282), .Y(N7) );
  AND2X1 U266 ( .A(n598), .B(R2[3]), .Y(n67) );
  OR3X4 U267 ( .A(n69), .B(n68), .C(n513), .Y(n609) );
  NAND2BXL U268 ( .AN(n256), .B(data_in_2[50]), .Y(n352) );
  AND3X4 U269 ( .A(n465), .B(n464), .C(n463), .Y(n71) );
  NAND2BXL U270 ( .AN(n256), .B(data_in_2[85]), .Y(n455) );
  AND3X4 U271 ( .A(n366), .B(n365), .C(n364), .Y(n72) );
  NAND2XL U272 ( .A(R2[22]), .B(n226), .Y(n370) );
  NAND2X2 U273 ( .A(data_in_2[88]), .B(n305), .Y(n465) );
  NAND2XL U274 ( .A(R2[4]), .B(n246), .Y(n316) );
  NAND2XL U275 ( .A(R3[7]), .B(n246), .Y(n427) );
  NAND2XL U276 ( .A(data_in_1[75]), .B(n240), .Y(n428) );
  NAND2XL U277 ( .A(data_in_2[75]), .B(n229), .Y(n429) );
  NAND2XL U278 ( .A(data_in_2[74]), .B(n296), .Y(n426) );
  NAND2XL U279 ( .A(R2[5]), .B(n4), .Y(n319) );
  NAND2XL U280 ( .A(data_in_1[39]), .B(n240), .Y(n320) );
  NAND2XL U281 ( .A(data_in_2[39]), .B(n296), .Y(n321) );
  NAND2XL U282 ( .A(data_in_1[126]), .B(n594), .Y(n579) );
  NAND2XL U283 ( .A(data_in_2[126]), .B(n233), .Y(n580) );
  NAND2XL U284 ( .A(data_in_1[109]), .B(n594), .Y(n527) );
  NAND2XL U285 ( .A(data_in_2[109]), .B(n231), .Y(n528) );
  NAND2XL U286 ( .A(R4[23]), .B(n42), .Y(n575) );
  NAND2XL U287 ( .A(data_in_2[125]), .B(n231), .Y(n577) );
  NAND2XL U288 ( .A(R2[24]), .B(n223), .Y(n376) );
  NAND2XL U289 ( .A(data_in_2[58]), .B(n229), .Y(n378) );
  NAND2XL U290 ( .A(R3[5]), .B(n223), .Y(n421) );
  NAND2XL U291 ( .A(data_in_2[73]), .B(n230), .Y(n423) );
  NAND2XL U292 ( .A(data_in_1[91]), .B(n241), .Y(n473) );
  NAND2XL U293 ( .A(data_in_2[91]), .B(n228), .Y(n474) );
  NAND2XL U294 ( .A(R3[22]), .B(n226), .Y(n469) );
  NAND2XL U295 ( .A(data_in_1[90]), .B(n242), .Y(n470) );
  NAND2XL U296 ( .A(data_in_2[90]), .B(n305), .Y(n471) );
  NAND2BXL U297 ( .AN(n256), .B(data_in_2[104]), .Y(n511) );
  NAND2XL U298 ( .A(R4[6]), .B(n29), .Y(n523) );
  NAND2XL U299 ( .A(data_in_1[108]), .B(n237), .Y(n524) );
  NAND2XL U300 ( .A(data_in_2[108]), .B(n228), .Y(n525) );
  NAND2XL U301 ( .A(R2[23]), .B(n246), .Y(n373) );
  NAND2XL U302 ( .A(data_in_1[57]), .B(n240), .Y(n374) );
  NAND2XL U303 ( .A(R4[5]), .B(n223), .Y(n520) );
  NAND2XL U304 ( .A(data_in_1[107]), .B(n242), .Y(n521) );
  NAND2XL U305 ( .A(data_in_2[107]), .B(n231), .Y(n522) );
  NAND2XL U306 ( .A(R2[6]), .B(n19), .Y(n322) );
  NAND2XL U307 ( .A(data_in_1[40]), .B(n240), .Y(n323) );
  NAND2XL U308 ( .A(data_in_2[40]), .B(n298), .Y(n324) );
  NAND2XL U309 ( .A(R4[22]), .B(n223), .Y(n572) );
  NAND2XL U310 ( .A(data_in_1[124]), .B(n241), .Y(n573) );
  NAND2XL U311 ( .A(data_in_2[124]), .B(n229), .Y(n574) );
  NAND2XL U312 ( .A(data_in_1[63]), .B(n241), .Y(n392) );
  NAND2XL U313 ( .A(data_in_2[63]), .B(n305), .Y(n393) );
  NAND2XL U314 ( .A(R2[28]), .B(n246), .Y(n388) );
  NAND2XL U315 ( .A(data_in_1[62]), .B(n241), .Y(n389) );
  NAND2XL U316 ( .A(data_in_2[62]), .B(n305), .Y(n390) );
  NAND2XL U317 ( .A(data_in_1[61]), .B(n238), .Y(n386) );
  NAND2XL U318 ( .A(data_in_2[61]), .B(n231), .Y(n387) );
  NAND2XL U319 ( .A(R2[26]), .B(n223), .Y(n382) );
  NAND2XL U320 ( .A(data_in_1[60]), .B(n242), .Y(n383) );
  NAND2XL U321 ( .A(data_in_2[60]), .B(n305), .Y(n384) );
  NAND2XL U322 ( .A(data_in_1[59]), .B(n241), .Y(n380) );
  NAND2XL U323 ( .A(data_in_1[77]), .B(n237), .Y(n434) );
  NAND2XL U324 ( .A(data_in_2[77]), .B(n305), .Y(n435) );
  NAND2XL U325 ( .A(R4[9]), .B(n2), .Y(n532) );
  NAND2XL U326 ( .A(data_in_1[111]), .B(n237), .Y(n533) );
  NAND2XL U327 ( .A(data_in_2[111]), .B(n298), .Y(n534) );
  NAND2XL U328 ( .A(R3[8]), .B(n29), .Y(n430) );
  NAND2XL U329 ( .A(data_in_1[76]), .B(n594), .Y(n431) );
  NAND2XL U330 ( .A(data_in_2[76]), .B(n298), .Y(n432) );
  NAND2XL U331 ( .A(R4[8]), .B(n13), .Y(n529) );
  NAND2XL U332 ( .A(data_in_1[110]), .B(n238), .Y(n530) );
  NAND2XL U333 ( .A(data_in_2[110]), .B(n228), .Y(n531) );
  NAND2XL U334 ( .A(R3[26]), .B(n246), .Y(n481) );
  NAND2XL U335 ( .A(data_in_1[94]), .B(n594), .Y(n482) );
  NAND2XL U336 ( .A(R3[25]), .B(n32), .Y(n478) );
  NAND2XL U337 ( .A(data_in_1[93]), .B(n240), .Y(n479) );
  NAND2XL U338 ( .A(data_in_2[93]), .B(n232), .Y(n480) );
  NAND2XL U339 ( .A(R3[24]), .B(n13), .Y(n475) );
  NAND2XL U340 ( .A(data_in_1[92]), .B(n241), .Y(n476) );
  NAND2XL U341 ( .A(R2[9]), .B(n223), .Y(n331) );
  NAND2XL U342 ( .A(data_in_1[43]), .B(n238), .Y(n332) );
  NAND2XL U343 ( .A(data_in_2[43]), .B(n233), .Y(n333) );
  NAND2XL U344 ( .A(R2[8]), .B(n246), .Y(n328) );
  NAND2XL U345 ( .A(data_in_1[42]), .B(n594), .Y(n329) );
  NAND2XL U346 ( .A(data_in_2[42]), .B(n229), .Y(n330) );
  NAND2XL U347 ( .A(data_in_2[41]), .B(n228), .Y(n327) );
  AND2X1 U348 ( .A(data_in_2[129]), .B(n298), .Y(n73) );
  OR3X4 U349 ( .A(n74), .B(n75), .C(n76), .Y(data_out[128]) );
  AND2X1 U350 ( .A(data_in_2[128]), .B(n296), .Y(n74) );
  AND2X1 U351 ( .A(R4[26]), .B(n244), .Y(n76) );
  OR3X4 U352 ( .A(n77), .B(n78), .C(n79), .Y(data_out[127]) );
  AND2X1 U353 ( .A(data_in_2[127]), .B(n232), .Y(n77) );
  NAND2XL U354 ( .A(R2[32]), .B(n223), .Y(n400) );
  NAND2XL U355 ( .A(data_in_1[66]), .B(n240), .Y(n401) );
  NAND2XL U356 ( .A(data_in_2[66]), .B(n233), .Y(n402) );
  NAND2XL U357 ( .A(data_in_1[80]), .B(n594), .Y(n443) );
  NAND2XL U358 ( .A(data_in_2[80]), .B(n228), .Y(n444) );
  NAND2XL U359 ( .A(R3[11]), .B(n244), .Y(n439) );
  NAND2XL U360 ( .A(data_in_1[79]), .B(n241), .Y(n440) );
  NAND2XL U361 ( .A(data_in_2[79]), .B(n298), .Y(n441) );
  NAND2XL U362 ( .A(R4[30]), .B(n246), .Y(n587) );
  NAND2XL U363 ( .A(data_in_1[132]), .B(n237), .Y(n588) );
  NAND2XL U364 ( .A(data_in_2[132]), .B(n298), .Y(n589) );
  NAND2XL U365 ( .A(R4[29]), .B(n223), .Y(n584) );
  NAND2XL U366 ( .A(data_in_1[131]), .B(n240), .Y(n585) );
  NAND2XL U367 ( .A(data_in_2[131]), .B(n231), .Y(n586) );
  NAND2XL U368 ( .A(R4[12]), .B(n13), .Y(n541) );
  NAND2XL U369 ( .A(data_in_1[114]), .B(n240), .Y(n542) );
  NAND2XL U370 ( .A(data_in_2[114]), .B(n280), .Y(n543) );
  NAND2XL U371 ( .A(data_in_1[64]), .B(n240), .Y(n395) );
  NAND2XL U372 ( .A(data_in_2[64]), .B(n298), .Y(n396) );
  NAND2XL U373 ( .A(R2[12]), .B(n223), .Y(n340) );
  NAND2XL U374 ( .A(data_in_1[46]), .B(n242), .Y(n341) );
  NAND2XL U375 ( .A(data_in_2[46]), .B(n296), .Y(n342) );
  NAND2XL U376 ( .A(R2[31]), .B(n246), .Y(n397) );
  NAND2XL U377 ( .A(data_in_1[65]), .B(n241), .Y(n398) );
  NAND2XL U378 ( .A(data_in_2[65]), .B(n232), .Y(n399) );
  NAND2XL U379 ( .A(R2[11]), .B(n223), .Y(n337) );
  NAND2XL U380 ( .A(data_in_1[45]), .B(n239), .Y(n338) );
  NAND2XL U381 ( .A(data_in_2[45]), .B(n298), .Y(n339) );
  NAND2XL U382 ( .A(R3[29]), .B(n246), .Y(n490) );
  NAND2XL U383 ( .A(data_in_1[97]), .B(n242), .Y(n491) );
  NAND2XL U384 ( .A(data_in_2[97]), .B(n229), .Y(n492) );
  NAND2XL U385 ( .A(data_in_1[96]), .B(n237), .Y(n488) );
  NAND2XL U386 ( .A(R3[10]), .B(n223), .Y(n436) );
  NAND2XL U387 ( .A(data_in_1[78]), .B(n241), .Y(n437) );
  NAND2XL U388 ( .A(data_in_2[78]), .B(n305), .Y(n438) );
  NAND2XL U389 ( .A(R4[11]), .B(n3), .Y(n538) );
  NAND2XL U390 ( .A(data_in_1[113]), .B(n242), .Y(n539) );
  NAND2XL U391 ( .A(data_in_2[113]), .B(n280), .Y(n540) );
  NAND2XL U392 ( .A(R4[10]), .B(n226), .Y(n535) );
  NAND2XL U393 ( .A(data_in_1[112]), .B(n241), .Y(n536) );
  NAND2XL U394 ( .A(data_in_2[112]), .B(n233), .Y(n537) );
  NAND2XL U395 ( .A(R3[27]), .B(n32), .Y(n484) );
  NAND2XL U396 ( .A(data_in_2[95]), .B(n229), .Y(n486) );
  NAND2XL U397 ( .A(R2[10]), .B(n29), .Y(n334) );
  NAND2XL U398 ( .A(data_in_1[44]), .B(n241), .Y(n335) );
  NAND2XL U399 ( .A(data_in_2[44]), .B(n231), .Y(n336) );
  NAND2XL U400 ( .A(R4[28]), .B(n2), .Y(n581) );
  NAND2XL U401 ( .A(data_in_1[130]), .B(n242), .Y(n582) );
  NAND2XL U402 ( .A(data_in_2[130]), .B(n232), .Y(n583) );
  OR3X4 U403 ( .A(n80), .B(n81), .C(n82), .Y(data_out[83]) );
  AND2X1 U404 ( .A(data_in_2[83]), .B(n296), .Y(n80) );
  AND2X1 U405 ( .A(data_in_1[83]), .B(n240), .Y(n81) );
  AND2X2 U406 ( .A(R3[15]), .B(n226), .Y(n82) );
  NAND2XL U407 ( .A(R4[15]), .B(n13), .Y(n550) );
  NAND2XL U408 ( .A(data_in_1[117]), .B(n237), .Y(n551) );
  NAND2XL U409 ( .A(data_in_2[117]), .B(n305), .Y(n552) );
  NAND2XL U410 ( .A(R3[32]), .B(n223), .Y(n499) );
  NAND2XL U411 ( .A(data_in_1[100]), .B(n239), .Y(n500) );
  NAND2XL U412 ( .A(data_in_2[100]), .B(n298), .Y(n501) );
  NAND2XL U413 ( .A(data_in_1[81]), .B(n238), .Y(n446) );
  NAND2XL U414 ( .A(data_in_2[81]), .B(n280), .Y(n447) );
  NAND2XL U415 ( .A(data_in_1[82]), .B(n241), .Y(n449) );
  NAND2XL U416 ( .A(data_in_2[82]), .B(n233), .Y(n450) );
  NAND2XL U417 ( .A(R4[31]), .B(n223), .Y(n590) );
  NAND2XL U418 ( .A(data_in_1[133]), .B(n241), .Y(n591) );
  NAND2XL U419 ( .A(data_in_2[133]), .B(n229), .Y(n592) );
  NAND2XL U420 ( .A(R4[13]), .B(n29), .Y(n544) );
  NAND2XL U421 ( .A(data_in_1[115]), .B(n238), .Y(n545) );
  NAND2XL U422 ( .A(data_in_2[115]), .B(n232), .Y(n546) );
  NAND2XL U423 ( .A(R4[14]), .B(n244), .Y(n547) );
  NAND2XL U424 ( .A(data_in_1[116]), .B(n237), .Y(n548) );
  NAND2XL U425 ( .A(data_in_2[116]), .B(n305), .Y(n549) );
  NAND2XL U426 ( .A(R2[13]), .B(n226), .Y(n343) );
  NAND2XL U427 ( .A(data_in_1[47]), .B(n594), .Y(n344) );
  NAND2XL U428 ( .A(data_in_2[47]), .B(n17), .Y(n345) );
  NAND2XL U429 ( .A(data_in_1[48]), .B(n238), .Y(n347) );
  NAND2XL U430 ( .A(data_in_2[48]), .B(n229), .Y(n348) );
  NAND2XL U431 ( .A(R3[30]), .B(n2), .Y(n493) );
  NAND2XL U432 ( .A(data_in_1[98]), .B(n240), .Y(n494) );
  NAND2XL U433 ( .A(data_in_2[98]), .B(n305), .Y(n495) );
  NAND2XL U434 ( .A(R3[31]), .B(n223), .Y(n496) );
  NAND2XL U435 ( .A(data_in_1[99]), .B(n239), .Y(n497) );
  NAND2XL U436 ( .A(data_in_2[99]), .B(n229), .Y(n498) );
  NAND2XL U437 ( .A(R2[15]), .B(n244), .Y(n349) );
  NAND2XL U438 ( .A(data_in_1[49]), .B(n242), .Y(n350) );
  NAND2XL U439 ( .A(data_in_2[49]), .B(n280), .Y(n351) );
  NAND2XL U440 ( .A(R4[32]), .B(n13), .Y(n595) );
  NAND2XL U441 ( .A(data_in_1[134]), .B(n238), .Y(n596) );
  NAND2XL U442 ( .A(data_in_2[134]), .B(n231), .Y(n597) );
  OAI2BB1X1 U443 ( .A0N(data_in_2[7]), .A1N(n228), .B0(n268), .Y(data_out[7])
         );
  OAI2BB1X1 U444 ( .A0N(data_in_2[4]), .A1N(n228), .B0(n265), .Y(data_out[4])
         );
  OAI2BB1X1 U445 ( .A0N(data_in_2[0]), .A1N(n229), .B0(n261), .Y(data_out[0])
         );
  OAI2BB1X1 U446 ( .A0N(data_in_2[1]), .A1N(n232), .B0(n262), .Y(data_out[1])
         );
  OAI2BB1X1 U447 ( .A0N(data_in_2[3]), .A1N(n228), .B0(n264), .Y(data_out[3])
         );
  OAI2BB1X1 U448 ( .A0N(data_in_2[6]), .A1N(n231), .B0(n267), .Y(data_out[6])
         );
  OAI2BB1X1 U449 ( .A0N(data_in_2[5]), .A1N(n231), .B0(n266), .Y(data_out[5])
         );
  OAI2BB1X1 U450 ( .A0N(data_in_2[2]), .A1N(n233), .B0(n263), .Y(data_out[2])
         );
  OAI2BB1X1 U451 ( .A0N(data_in_2[18]), .A1N(n229), .B0(n286), .Y(data_out[18]) );
  OAI2BB1X1 U452 ( .A0N(data_in_2[19]), .A1N(n305), .B0(n287), .Y(data_out[19]) );
  OAI2BB1X1 U453 ( .A0N(data_in_2[22]), .A1N(n296), .B0(n290), .Y(data_out[22]) );
  OAI2BB1X1 U454 ( .A0N(data_in_2[20]), .A1N(n298), .B0(n288), .Y(data_out[20]) );
  AOI22XL U455 ( .A0(data_in_1[20]), .A1(n242), .B0(R1[20]), .B1(n29), .Y(n288) );
  OAI2BB1X1 U456 ( .A0N(data_in_2[23]), .A1N(n305), .B0(n291), .Y(data_out[23]) );
  AOI22XL U457 ( .A0(data_in_1[23]), .A1(n594), .B0(R1[23]), .B1(n29), .Y(n291) );
  OAI2BB1X1 U458 ( .A0N(data_in_2[17]), .A1N(n231), .B0(n284), .Y(data_out[17]) );
  AOI22XL U459 ( .A0(data_in_1[17]), .A1(n240), .B0(R1[17]), .B1(n29), .Y(n284) );
  INVX1 U460 ( .A(data_in_2[12]), .Y(n275) );
  AOI22XL U461 ( .A0(data_in_1[28]), .A1(n237), .B0(R1[28]), .B1(n13), .Y(n297) );
  OAI2BB1X2 U462 ( .A0N(data_in_2[27]), .A1N(n229), .B0(n295), .Y(data_out[27]) );
  AOI22XL U463 ( .A0(data_in_1[27]), .A1(n241), .B0(R1[27]), .B1(n223), .Y(
        n295) );
  OAI2BB1X1 U464 ( .A0N(data_in_2[10]), .A1N(n298), .B0(n271), .Y(data_out[10]) );
  OAI2BB1X1 U465 ( .A0N(data_in_2[9]), .A1N(n229), .B0(n270), .Y(data_out[9])
         );
  OAI2BB1X1 U466 ( .A0N(data_in_2[8]), .A1N(n280), .B0(n269), .Y(data_out[8])
         );
  OAI2BB1X1 U467 ( .A0N(data_in_2[21]), .A1N(n17), .B0(n289), .Y(data_out[21])
         );
  OAI2BB1X1 U468 ( .A0N(data_in_2[24]), .A1N(n298), .B0(n292), .Y(data_out[24]) );
  OAI2BB1X1 U469 ( .A0N(data_in_2[26]), .A1N(n298), .B0(n294), .Y(data_out[26]) );
  AOI22XL U470 ( .A0(data_in_1[26]), .A1(n239), .B0(R1[26]), .B1(n37), .Y(n294) );
  OAI2BB1X1 U471 ( .A0N(data_in_2[25]), .A1N(n232), .B0(n293), .Y(data_out[25]) );
  AOI22XL U472 ( .A0(data_in_1[25]), .A1(n242), .B0(R1[25]), .B1(n246), .Y(
        n293) );
  OR2X2 U473 ( .A(n302), .B(n83), .Y(data_out[29]) );
  AND2X1 U474 ( .A(R1[29]), .B(n223), .Y(n83) );
  OAI2BB1X2 U475 ( .A0N(data_in_2[30]), .A1N(n296), .B0(n304), .Y(data_out[30]) );
  AOI22XL U476 ( .A0(data_in_1[30]), .A1(n238), .B0(R1[30]), .B1(n223), .Y(
        n304) );
  AOI22XL U477 ( .A0(data_in_1[13]), .A1(n242), .B0(R1[13]), .B1(n226), .Y(
        n277) );
  OAI2BB1X1 U478 ( .A0N(data_in_2[14]), .A1N(n231), .B0(n278), .Y(data_out[14]) );
  OAI2BB1X1 U479 ( .A0N(data_in_2[31]), .A1N(n228), .B0(n306), .Y(data_out[31]) );
  AOI22XL U480 ( .A0(data_in_1[31]), .A1(n237), .B0(R1[31]), .B1(n226), .Y(
        n306) );
  OAI2BB1X1 U481 ( .A0N(data_in_2[32]), .A1N(n298), .B0(n307), .Y(data_out[32]) );
  AOI22XL U482 ( .A0(data_in_1[32]), .A1(n594), .B0(R1[32]), .B1(n246), .Y(
        n307) );
  OAI2BB1X1 U483 ( .A0N(data_in_2[33]), .A1N(n228), .B0(n308), .Y(data_out[33]) );
  AOI22XL U484 ( .A0(data_in_1[33]), .A1(n242), .B0(R1[33]), .B1(n246), .Y(
        n308) );
  OAI2BB1X1 U485 ( .A0N(data_in_2[16]), .A1N(n17), .B0(n283), .Y(data_out[16])
         );
  INVX1 U486 ( .A(data_in_1[12]), .Y(n274) );
  INVX1 U487 ( .A(data_in_1[29]), .Y(n299) );
  NOR2X1 U488 ( .A(n603), .B(n282), .Y(n281) );
  INVXL U489 ( .A(n38), .Y(n603) );
  INVXL U490 ( .A(counter[3]), .Y(n604) );
  INVXL U491 ( .A(n36), .Y(n211) );
  CLKINVX8 U492 ( .A(n140), .Y(n212) );
  OAI22XL U493 ( .A0(n236), .A1(n301), .B0(n51), .B1(n299), .Y(n302) );
  OAI22XL U494 ( .A0(n222), .A1(n275), .B0(n51), .B1(n274), .Y(n276) );
  BUFX20 U495 ( .A(n614), .Y(data_out[50]) );
  AND2X4 U496 ( .A(data_in_1[68]), .B(n255), .Y(n407) );
  AOI22XL U497 ( .A0(data_in_1[10]), .A1(n240), .B0(R1[10]), .B1(n29), .Y(n271) );
  AOI22XL U498 ( .A0(data_in_1[9]), .A1(n238), .B0(R1[9]), .B1(n223), .Y(n270)
         );
  AOI22XL U499 ( .A0(data_in_1[7]), .A1(n237), .B0(R1[7]), .B1(n244), .Y(n268)
         );
  AOI22XL U500 ( .A0(data_in_1[4]), .A1(n241), .B0(R1[4]), .B1(n32), .Y(n265)
         );
  AOI22XL U501 ( .A0(data_in_1[3]), .A1(n238), .B0(R1[3]), .B1(n223), .Y(n264)
         );
  AOI22XL U502 ( .A0(data_in_1[0]), .A1(n240), .B0(R1[0]), .B1(n246), .Y(n261)
         );
  AOI22XL U503 ( .A0(data_in_1[1]), .A1(n594), .B0(R1[1]), .B1(n223), .Y(n262)
         );
  NOR4BXL U504 ( .AN(n224), .B(n603), .C(n604), .D(n211), .Y(n285) );
  NAND2XL U505 ( .A(n224), .B(n211), .Y(n282) );
  XOR2X1 U506 ( .A(n40), .B(n281), .Y(N8) );
  NOR2X4 U507 ( .A(counter[3]), .B(counter[2]), .Y(n259) );
  NAND2X4 U508 ( .A(n259), .B(counter[1]), .Y(n503) );
  AND2X2 U509 ( .A(data_in_1[34]), .B(n255), .Y(n310) );
  OAI2BB1X4 U510 ( .A0N(R2[0]), .A1N(n247), .B0(n311), .Y(n617) );
  AND2X2 U511 ( .A(data_in_1[35]), .B(n255), .Y(n314) );
  NAND3X4 U512 ( .A(n318), .B(n317), .C(n316), .Y(data_out[38]) );
  NAND3X4 U513 ( .A(n321), .B(n320), .C(n319), .Y(data_out[39]) );
  NAND3X4 U514 ( .A(n324), .B(n323), .C(n322), .Y(data_out[40]) );
  NAND3X4 U515 ( .A(n327), .B(n326), .C(n325), .Y(data_out[41]) );
  NAND3X4 U516 ( .A(n330), .B(n329), .C(n328), .Y(data_out[42]) );
  NAND3X4 U517 ( .A(n333), .B(n332), .C(n331), .Y(data_out[43]) );
  NAND3X4 U518 ( .A(n336), .B(n335), .C(n334), .Y(data_out[44]) );
  NAND3X4 U519 ( .A(n339), .B(n338), .C(n337), .Y(data_out[45]) );
  NAND3X4 U520 ( .A(n342), .B(n341), .C(n340), .Y(data_out[46]) );
  NAND3X4 U521 ( .A(n345), .B(n344), .C(n343), .Y(data_out[47]) );
  NAND3X4 U522 ( .A(n348), .B(n347), .C(n346), .Y(data_out[48]) );
  NAND3X4 U523 ( .A(n351), .B(n350), .C(n349), .Y(data_out[49]) );
  AND2X2 U524 ( .A(data_in_1[50]), .B(n255), .Y(n353) );
  OAI2BB1X4 U525 ( .A0N(R2[16]), .A1N(n247), .B0(n354), .Y(n614) );
  AND2X2 U526 ( .A(data_in_1[51]), .B(n255), .Y(n356) );
  NAND2BX4 U527 ( .AN(n256), .B(data_in_2[51]), .Y(n355) );
  AND2X2 U528 ( .A(data_in_1[52]), .B(n255), .Y(n360) );
  OAI2BB1X4 U529 ( .A0N(n360), .A1N(n44), .B0(n359), .Y(data_out[52]) );
  NAND2X4 U530 ( .A(data_in_2[55]), .B(n305), .Y(n369) );
  NAND3X4 U531 ( .A(n369), .B(n368), .C(n367), .Y(data_out[55]) );
  NAND3X4 U532 ( .A(n372), .B(n371), .C(n370), .Y(data_out[56]) );
  NAND3X4 U533 ( .A(n375), .B(n374), .C(n373), .Y(data_out[57]) );
  NAND3X4 U534 ( .A(n378), .B(n377), .C(n376), .Y(data_out[58]) );
  NAND3X4 U535 ( .A(n381), .B(n380), .C(n379), .Y(data_out[59]) );
  NAND3X4 U536 ( .A(n384), .B(n383), .C(n382), .Y(data_out[60]) );
  NAND3X4 U537 ( .A(n387), .B(n386), .C(n385), .Y(data_out[61]) );
  NAND3X4 U538 ( .A(n390), .B(n389), .C(n388), .Y(data_out[62]) );
  NAND3X4 U539 ( .A(n393), .B(n392), .C(n391), .Y(data_out[63]) );
  NAND3X4 U540 ( .A(n399), .B(n398), .C(n397), .Y(data_out[65]) );
  NAND3X4 U541 ( .A(n402), .B(n401), .C(n400), .Y(data_out[66]) );
  NAND2BX4 U542 ( .AN(n405), .B(n404), .Y(n613) );
  AND2X2 U543 ( .A(data_in_1[69]), .B(n256), .Y(n411) );
  OAI2BB1X4 U544 ( .A0N(n411), .A1N(n46), .B0(n410), .Y(data_out[69]) );
  NAND2X4 U545 ( .A(data_in_2[71]), .B(n232), .Y(n417) );
  NAND2X4 U546 ( .A(data_in_1[71]), .B(n242), .Y(n416) );
  NAND3X4 U547 ( .A(n417), .B(n416), .C(n415), .Y(n612) );
  NAND3X4 U548 ( .A(n420), .B(n419), .C(n418), .Y(data_out[72]) );
  NAND3X4 U549 ( .A(n423), .B(n422), .C(n421), .Y(data_out[73]) );
  NAND3X4 U550 ( .A(n426), .B(n425), .C(n424), .Y(data_out[74]) );
  NAND3X4 U551 ( .A(n429), .B(n428), .C(n427), .Y(data_out[75]) );
  NAND3X4 U552 ( .A(n432), .B(n431), .C(n430), .Y(data_out[76]) );
  NAND3X4 U553 ( .A(n435), .B(n434), .C(n433), .Y(data_out[77]) );
  NAND3X4 U554 ( .A(n438), .B(n437), .C(n436), .Y(data_out[78]) );
  NAND3X4 U555 ( .A(n441), .B(n440), .C(n439), .Y(data_out[79]) );
  NAND3X4 U556 ( .A(n444), .B(n443), .C(n442), .Y(data_out[80]) );
  NAND3X4 U557 ( .A(n447), .B(n446), .C(n445), .Y(data_out[81]) );
  NAND3X4 U558 ( .A(n450), .B(n449), .C(n448), .Y(data_out[82]) );
  NAND2X4 U559 ( .A(data_in_1[84]), .B(n255), .Y(n452) );
  NAND2BX4 U560 ( .AN(n454), .B(n453), .Y(data_out[84]) );
  AND2X2 U561 ( .A(data_in_1[85]), .B(n256), .Y(n456) );
  OAI2BB1X4 U562 ( .A0N(R3[17]), .A1N(n247), .B0(n457), .Y(n611) );
  AND2X2 U563 ( .A(data_in_1[86]), .B(n255), .Y(n460) );
  NAND2X4 U564 ( .A(data_in_2[89]), .B(n298), .Y(n468) );
  NAND3X4 U565 ( .A(n474), .B(n473), .C(n472), .Y(data_out[91]) );
  NAND3X4 U566 ( .A(n477), .B(n476), .C(n475), .Y(data_out[92]) );
  NAND3X4 U567 ( .A(n480), .B(n479), .C(n478), .Y(data_out[93]) );
  NAND3X4 U568 ( .A(n483), .B(n482), .C(n481), .Y(data_out[94]) );
  NAND3X4 U569 ( .A(n486), .B(n485), .C(n484), .Y(data_out[95]) );
  NAND3X4 U570 ( .A(n489), .B(n488), .C(n487), .Y(data_out[96]) );
  NAND3X4 U571 ( .A(n492), .B(n491), .C(n490), .Y(data_out[97]) );
  NAND3X4 U572 ( .A(n495), .B(n494), .C(n493), .Y(data_out[98]) );
  NAND3X4 U573 ( .A(n498), .B(n497), .C(n496), .Y(data_out[99]) );
  NAND3X4 U574 ( .A(n501), .B(n500), .C(n499), .Y(data_out[100]) );
  AND2X2 U575 ( .A(data_in_1[102]), .B(n255), .Y(n507) );
  OAI2BB1X4 U576 ( .A0N(n507), .A1N(n20), .B0(n506), .Y(data_out[102]) );
  AND2X2 U577 ( .A(data_in_1[103]), .B(n255), .Y(n509) );
  OAI2BB1X4 U578 ( .A0N(R4[1]), .A1N(n247), .B0(n510), .Y(data_out[103]) );
  AND2X2 U579 ( .A(data_in_1[104]), .B(n255), .Y(n512) );
  NAND2X4 U580 ( .A(data_in_2[105]), .B(n233), .Y(n516) );
  NAND2X4 U581 ( .A(data_in_1[105]), .B(n241), .Y(n515) );
  NAND3X4 U582 ( .A(n516), .B(n515), .C(n514), .Y(data_out[105]) );
  NAND3X4 U583 ( .A(n519), .B(n518), .C(n517), .Y(data_out[106]) );
  NAND3X4 U584 ( .A(n522), .B(n521), .C(n520), .Y(data_out[107]) );
  NAND3X4 U585 ( .A(n525), .B(n524), .C(n523), .Y(data_out[108]) );
  NAND3X4 U586 ( .A(n528), .B(n527), .C(n526), .Y(data_out[109]) );
  NAND3X4 U587 ( .A(n531), .B(n530), .C(n529), .Y(data_out[110]) );
  NAND3X4 U588 ( .A(n534), .B(n533), .C(n532), .Y(data_out[111]) );
  NAND3X4 U589 ( .A(n537), .B(n536), .C(n535), .Y(data_out[112]) );
  NAND3X4 U590 ( .A(n543), .B(n542), .C(n541), .Y(data_out[114]) );
  NAND3X4 U591 ( .A(n546), .B(n545), .C(n544), .Y(data_out[115]) );
  NAND3X4 U592 ( .A(n549), .B(n548), .C(n547), .Y(data_out[116]) );
  NAND3X4 U593 ( .A(n552), .B(n551), .C(n550), .Y(data_out[117]) );
  AND2X2 U594 ( .A(data_in_1[119]), .B(n255), .Y(n557) );
  AND2X2 U595 ( .A(data_in_1[120]), .B(n255), .Y(n562) );
  OAI2BB1X4 U596 ( .A0N(n562), .A1N(n47), .B0(n560), .Y(n607) );
  NAND2X4 U597 ( .A(data_in_1[122]), .B(n241), .Y(n567) );
  NAND3X4 U598 ( .A(n568), .B(n567), .C(n566), .Y(data_out[122]) );
  NAND3X4 U599 ( .A(n571), .B(n570), .C(n569), .Y(data_out[123]) );
  NAND3X4 U600 ( .A(n574), .B(n573), .C(n572), .Y(data_out[124]) );
  NAND3X4 U601 ( .A(n577), .B(n576), .C(n575), .Y(data_out[125]) );
  NAND3X4 U602 ( .A(n580), .B(n579), .C(n578), .Y(data_out[126]) );
  NAND3X4 U603 ( .A(n583), .B(n582), .C(n581), .Y(data_out[130]) );
  NAND3X4 U604 ( .A(n586), .B(n585), .C(n584), .Y(data_out[131]) );
  NAND3X4 U605 ( .A(n589), .B(n588), .C(n587), .Y(data_out[132]) );
  NAND3X4 U606 ( .A(n592), .B(n591), .C(n590), .Y(data_out[133]) );
  NAND3X4 U607 ( .A(n597), .B(n596), .C(n595), .Y(data_out[134]) );
endmodule


module multi16_11_DW01_add_5 ( A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, 
        A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, 
        B_20_, B_19_, B_18_, B_17_, B_16_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, 
        SUM_17_, SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, 
        SUM_9_, SUM_8_, SUM_7_, SUM_6_, SUM_5_ );
  input A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_,
         A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, B_20_, B_19_,
         B_18_, B_17_, B_16_;
  output SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, SUM_15_,
         SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, SUM_7_,
         SUM_6_, SUM_5_;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46;

  INVX4 U2 ( .A(n38), .Y(n1) );
  INVX8 U3 ( .A(n34), .Y(n38) );
  NAND2X4 U4 ( .A(B_18_), .B(A_18_), .Y(n34) );
  NOR2X4 U5 ( .A(A_18_), .B(B_18_), .Y(n2) );
  BUFX4 U6 ( .A(A_16_), .Y(n5) );
  OR2X1 U7 ( .A(n8), .B(n34), .Y(n6) );
  AND3X4 U8 ( .A(n44), .B(n5), .C(B_16_), .Y(n3) );
  NOR2X2 U9 ( .A(n8), .B(n2), .Y(n29) );
  NAND2BX4 U10 ( .AN(n38), .B(n37), .Y(n35) );
  NOR2X2 U11 ( .A(A_17_), .B(B_17_), .Y(n4) );
  NAND2X4 U12 ( .A(n32), .B(n41), .Y(n42) );
  BUFX12 U13 ( .A(A_12_), .Y(SUM_12_) );
  AOI21X2 U14 ( .A0(n28), .A1(n29), .B0(n30), .Y(n27) );
  NAND2X1 U15 ( .A(n24), .B(n25), .Y(n23) );
  BUFX12 U16 ( .A(A_15_), .Y(SUM_15_) );
  BUFX12 U17 ( .A(A_14_), .Y(SUM_14_) );
  AOI21XL U18 ( .A0(n32), .A1(n33), .B0(n4), .Y(n28) );
  OR2X4 U19 ( .A(A_16_), .B(B_16_), .Y(n7) );
  NAND2X4 U20 ( .A(B_16_), .B(A_16_), .Y(n33) );
  CLKINVX3 U21 ( .A(n33), .Y(n45) );
  NAND2X4 U22 ( .A(n1), .B(n39), .Y(n43) );
  NAND2X4 U23 ( .A(B_17_), .B(A_17_), .Y(n32) );
  BUFX8 U24 ( .A(A_6_), .Y(SUM_6_) );
  NOR2BX4 U25 ( .AN(n31), .B(n8), .Y(n36) );
  NOR2X4 U26 ( .A(A_19_), .B(B_19_), .Y(n8) );
  XNOR2X4 U27 ( .A(n42), .B(n43), .Y(SUM_18_) );
  OR2X4 U28 ( .A(A_18_), .B(B_18_), .Y(n39) );
  NAND2X4 U29 ( .A(B_19_), .B(A_19_), .Y(n31) );
  NAND2X2 U30 ( .A(B_20_), .B(A_20_), .Y(n22) );
  NOR2X2 U31 ( .A(n2), .B(n32), .Y(n40) );
  AND2X4 U32 ( .A(n22), .B(n25), .Y(n26) );
  NAND3X4 U33 ( .A(n44), .B(n5), .C(B_16_), .Y(n41) );
  AND2X4 U34 ( .A(n7), .B(n33), .Y(SUM_16_) );
  OR2X4 U35 ( .A(A_20_), .B(B_20_), .Y(n25) );
  BUFX8 U36 ( .A(A_9_), .Y(SUM_9_) );
  BUFX8 U37 ( .A(A_7_), .Y(SUM_7_) );
  INVX1 U38 ( .A(n31), .Y(n30) );
  BUFX8 U39 ( .A(A_11_), .Y(SUM_11_) );
  BUFX8 U40 ( .A(A_10_), .Y(SUM_10_) );
  BUFX8 U41 ( .A(A_5_), .Y(SUM_5_) );
  BUFX8 U42 ( .A(A_8_), .Y(SUM_8_) );
  BUFX8 U43 ( .A(A_13_), .Y(SUM_13_) );
  XOR3X2 U44 ( .A(B_21_), .B(A_21_), .C(n21), .Y(SUM_21_) );
  NAND2XL U45 ( .A(n22), .B(n23), .Y(n21) );
  XOR2X4 U46 ( .A(n24), .B(n26), .Y(SUM_20_) );
  NAND2X4 U47 ( .A(n6), .B(n27), .Y(n24) );
  XOR2X4 U48 ( .A(n35), .B(n36), .Y(SUM_19_) );
  AOI21X4 U49 ( .A0(n3), .A1(n39), .B0(n40), .Y(n37) );
  XOR2X4 U50 ( .A(n46), .B(n45), .Y(SUM_17_) );
  NOR2BX4 U51 ( .AN(n32), .B(n4), .Y(n46) );
  OR2X4 U52 ( .A(A_17_), .B(B_17_), .Y(n44) );
endmodule


module multi16_11_DW02_mult_0 ( A, B, PRODUCT_23_, PRODUCT_22_, PRODUCT_21_, 
        PRODUCT_20_, PRODUCT_19_, PRODUCT_18_, PRODUCT_17_, PRODUCT_16_, 
        PRODUCT_15_, PRODUCT_14_, PRODUCT_13_, PRODUCT_12_, PRODUCT_11_, 
        PRODUCT_10_, PRODUCT_9_, PRODUCT_8_, PRODUCT_7_ );
  input [16:0] A;
  input [7:0] B;
  output PRODUCT_23_, PRODUCT_22_, PRODUCT_21_, PRODUCT_20_, PRODUCT_19_,
         PRODUCT_18_, PRODUCT_17_, PRODUCT_16_, PRODUCT_15_, PRODUCT_14_,
         PRODUCT_13_, PRODUCT_12_, PRODUCT_11_, PRODUCT_10_, PRODUCT_9_,
         PRODUCT_8_, PRODUCT_7_;
  wire   ab_16__7_, ab_16__6_, ab_16__5_, ab_16__4_, ab_16__3_, ab_16__2_,
         ab_16__1_, ab_16__0_, ab_15__7_, ab_15__6_, ab_15__5_, ab_15__4_,
         ab_15__3_, ab_15__2_, ab_15__1_, ab_15__0_, ab_14__7_, ab_14__6_,
         ab_14__5_, ab_14__4_, ab_14__3_, ab_14__2_, ab_14__1_, ab_14__0_,
         ab_13__7_, ab_13__6_, ab_13__5_, ab_13__4_, ab_13__3_, ab_13__2_,
         ab_13__1_, ab_13__0_, ab_12__7_, ab_12__6_, ab_12__5_, ab_12__4_,
         ab_12__3_, ab_12__2_, ab_12__1_, ab_12__0_, ab_11__7_, ab_11__6_,
         ab_11__5_, ab_11__4_, ab_11__3_, ab_11__2_, ab_11__1_, ab_11__0_,
         ab_10__7_, ab_10__6_, ab_10__5_, ab_10__4_, ab_10__3_, ab_10__2_,
         ab_10__1_, ab_10__0_, ab_9__7_, ab_9__6_, ab_9__5_, ab_9__4_,
         ab_9__3_, ab_9__2_, ab_9__1_, ab_9__0_, ab_8__7_, ab_8__6_, ab_8__5_,
         ab_8__4_, ab_8__3_, ab_8__2_, ab_8__1_, ab_8__0_, ab_7__7_, ab_7__6_,
         ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_, ab_7__0_, ab_6__7_,
         ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_, ab_6__1_, ab_6__0_,
         ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_, ab_5__2_, ab_5__1_,
         ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_, ab_4__3_, ab_4__2_,
         ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_, ab_3__4_, ab_3__3_,
         ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_, ab_2__5_, ab_2__4_,
         ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_, ab_1__6_, ab_1__5_,
         ab_1__4_, ab_1__3_, ab_1__2_, ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_,
         ab_0__3_, ab_0__2_, CARRYB_16__6_, CARRYB_16__5_, CARRYB_16__4_,
         CARRYB_16__3_, CARRYB_16__2_, CARRYB_16__1_, CARRYB_16__0_,
         CARRYB_15__6_, CARRYB_15__5_, CARRYB_15__4_, CARRYB_15__3_,
         CARRYB_15__2_, CARRYB_15__1_, CARRYB_15__0_, CARRYB_14__6_,
         CARRYB_14__5_, CARRYB_14__4_, CARRYB_14__3_, CARRYB_14__2_,
         CARRYB_14__1_, CARRYB_14__0_, CARRYB_13__6_, CARRYB_13__5_,
         CARRYB_13__4_, CARRYB_13__3_, CARRYB_13__2_, CARRYB_13__1_,
         CARRYB_13__0_, CARRYB_12__6_, CARRYB_12__5_, CARRYB_12__4_,
         CARRYB_12__3_, CARRYB_12__2_, CARRYB_12__1_, CARRYB_12__0_,
         CARRYB_11__6_, CARRYB_11__5_, CARRYB_11__4_, CARRYB_11__3_,
         CARRYB_11__2_, CARRYB_11__1_, CARRYB_11__0_, CARRYB_10__6_,
         CARRYB_10__5_, CARRYB_10__4_, CARRYB_10__3_, CARRYB_10__2_,
         CARRYB_10__1_, CARRYB_10__0_, CARRYB_9__6_, CARRYB_9__5_,
         CARRYB_9__4_, CARRYB_9__3_, CARRYB_9__2_, CARRYB_9__1_, CARRYB_9__0_,
         CARRYB_8__6_, CARRYB_8__5_, CARRYB_8__4_, CARRYB_8__3_, CARRYB_8__2_,
         CARRYB_8__1_, CARRYB_8__0_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_,
         CARRYB_7__3_, CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_,
         CARRYB_6__5_, CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_,
         CARRYB_6__0_, CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_,
         CARRYB_5__2_, CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_,
         CARRYB_4__4_, CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_,
         CARRYB_3__6_, CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_,
         CARRYB_3__1_, CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_,
         CARRYB_2__3_, CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__4_,
         CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_16__6_, SUMB_16__5_,
         SUMB_16__4_, SUMB_16__3_, SUMB_16__2_, SUMB_16__1_, SUMB_16__0_,
         SUMB_15__6_, SUMB_15__5_, SUMB_15__4_, SUMB_15__3_, SUMB_15__2_,
         SUMB_15__1_, SUMB_14__6_, SUMB_14__5_, SUMB_14__4_, SUMB_14__3_,
         SUMB_14__2_, SUMB_14__1_, SUMB_13__6_, SUMB_13__5_, SUMB_13__4_,
         SUMB_13__3_, SUMB_13__2_, SUMB_13__1_, SUMB_12__6_, SUMB_12__5_,
         SUMB_12__4_, SUMB_12__3_, SUMB_12__2_, SUMB_12__1_, SUMB_11__6_,
         SUMB_11__5_, SUMB_11__4_, SUMB_11__3_, SUMB_11__2_, SUMB_11__1_,
         SUMB_10__6_, SUMB_10__5_, SUMB_10__4_, SUMB_10__3_, SUMB_10__2_,
         SUMB_10__1_, SUMB_9__6_, SUMB_9__5_, SUMB_9__4_, SUMB_9__3_,
         SUMB_9__2_, SUMB_9__1_, SUMB_8__6_, SUMB_8__5_, SUMB_8__4_,
         SUMB_8__3_, SUMB_8__2_, SUMB_8__1_, SUMB_7__6_, SUMB_7__5_,
         SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_, SUMB_6__6_,
         SUMB_6__5_, SUMB_6__4_, SUMB_6__3_, SUMB_6__2_, SUMB_6__1_,
         SUMB_5__6_, SUMB_5__5_, SUMB_5__4_, SUMB_5__3_, SUMB_5__2_,
         SUMB_5__1_, SUMB_4__6_, SUMB_4__5_, SUMB_4__4_, SUMB_4__3_,
         SUMB_4__2_, SUMB_4__1_, SUMB_3__6_, SUMB_3__5_, SUMB_3__4_,
         SUMB_3__3_, SUMB_3__2_, SUMB_3__1_, SUMB_2__6_, SUMB_2__5_,
         SUMB_2__4_, SUMB_2__3_, SUMB_2__2_, SUMB_2__1_, SUMB_1__6_,
         SUMB_1__5_, SUMB_1__4_, SUMB_1__3_, SUMB_1__2_, SUMB_1__1_, PROD1_7_,
         A1_21_, A1_20_, A1_19_, A1_18_, A1_17_, A1_16_, A1_15_, A1_13_,
         A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, A1_4_, A1_3_,
         A1_2_, A1_1_, A1_0_, A2_16_, n3, n4, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43;

  multi16_11_DW01_add_5 FS_1 ( .A_21_(A1_21_), .A_20_(A1_20_), .A_19_(A1_19_), 
        .A_18_(A1_18_), .A_17_(A1_17_), .A_16_(A1_16_), .A_15_(A1_15_), 
        .A_14_(SUMB_16__0_), .A_13_(A1_13_), .A_12_(A1_12_), .A_11_(A1_11_), 
        .A_10_(A1_10_), .A_9_(A1_9_), .A_8_(A1_8_), .A_7_(A1_7_), .A_6_(A1_6_), 
        .A_5_(PROD1_7_), .B_21_(n6), .B_20_(n17), .B_19_(n15), .B_18_(n14), 
        .B_17_(n16), .B_16_(A2_16_), .SUM_21_(PRODUCT_23_), .SUM_20_(
        PRODUCT_22_), .SUM_19_(PRODUCT_21_), .SUM_18_(PRODUCT_20_), .SUM_17_(
        PRODUCT_19_), .SUM_16_(PRODUCT_18_), .SUM_15_(PRODUCT_17_), .SUM_14_(
        PRODUCT_16_), .SUM_13_(PRODUCT_15_), .SUM_12_(PRODUCT_14_), .SUM_11_(
        PRODUCT_13_), .SUM_10_(PRODUCT_12_), .SUM_9_(PRODUCT_11_), .SUM_8_(
        PRODUCT_10_), .SUM_7_(PRODUCT_9_), .SUM_6_(PRODUCT_8_), .SUM_5_(
        PRODUCT_7_) );
  ADDFHX4 S2_13_1 ( .A(ab_13__1_), .B(CARRYB_12__1_), .CI(SUMB_12__2_), .CO(
        CARRYB_13__1_), .S(SUMB_13__1_) );
  ADDFHX4 S2_11_5 ( .A(ab_11__5_), .B(CARRYB_10__5_), .CI(SUMB_10__6_), .CO(
        CARRYB_11__5_), .S(SUMB_11__5_) );
  ADDFHX4 S2_8_4 ( .A(ab_8__4_), .B(CARRYB_7__4_), .CI(SUMB_7__5_), .CO(
        CARRYB_8__4_), .S(SUMB_8__4_) );
  ADDFHX4 S2_9_3 ( .A(ab_9__3_), .B(CARRYB_8__3_), .CI(SUMB_8__4_), .CO(
        CARRYB_9__3_), .S(SUMB_9__3_) );
  ADDFHX4 S2_8_3 ( .A(ab_8__3_), .B(CARRYB_7__3_), .CI(SUMB_7__4_), .CO(
        CARRYB_8__3_), .S(SUMB_8__3_) );
  ADDFHX4 S2_15_1 ( .A(ab_15__1_), .B(CARRYB_14__1_), .CI(SUMB_14__2_), .CO(
        CARRYB_15__1_), .S(SUMB_15__1_) );
  ADDFHX4 S4_1 ( .A(ab_16__1_), .B(CARRYB_15__1_), .CI(SUMB_15__2_), .CO(
        CARRYB_16__1_), .S(SUMB_16__1_) );
  ADDFHX4 S4_0 ( .A(ab_16__0_), .B(CARRYB_15__0_), .CI(SUMB_15__1_), .CO(
        CARRYB_16__0_), .S(SUMB_16__0_) );
  ADDFHX4 S1_10_0 ( .A(ab_10__0_), .B(CARRYB_9__0_), .CI(SUMB_9__1_), .CO(
        CARRYB_10__0_), .S(A1_8_) );
  ADDFHX4 S1_11_0 ( .A(ab_11__0_), .B(CARRYB_10__0_), .CI(SUMB_10__1_), .CO(
        CARRYB_11__0_), .S(A1_9_) );
  ADDFHX4 S2_9_2 ( .A(ab_9__2_), .B(CARRYB_8__2_), .CI(SUMB_8__3_), .CO(
        CARRYB_9__2_), .S(SUMB_9__2_) );
  ADDFHX4 S2_12_2 ( .A(ab_12__2_), .B(CARRYB_11__2_), .CI(SUMB_11__3_), .CO(
        CARRYB_12__2_), .S(SUMB_12__2_) );
  ADDFHX4 S2_12_4 ( .A(ab_12__4_), .B(CARRYB_11__4_), .CI(SUMB_11__5_), .CO(
        CARRYB_12__4_), .S(SUMB_12__4_) );
  ADDFHX4 S2_13_4 ( .A(ab_13__4_), .B(CARRYB_12__4_), .CI(SUMB_12__5_), .CO(
        CARRYB_13__4_), .S(SUMB_13__4_) );
  ADDFHX4 S2_15_2 ( .A(ab_15__2_), .B(CARRYB_14__2_), .CI(SUMB_14__3_), .CO(
        CARRYB_15__2_), .S(SUMB_15__2_) );
  ADDFHX4 S1_14_0 ( .A(ab_14__0_), .B(CARRYB_13__0_), .CI(SUMB_13__1_), .CO(
        CARRYB_14__0_), .S(A1_12_) );
  ADDFHX4 S1_15_0 ( .A(ab_15__0_), .B(CARRYB_14__0_), .CI(SUMB_14__1_), .CO(
        CARRYB_15__0_), .S(A1_13_) );
  ADDFHX4 S1_8_0 ( .A(ab_8__0_), .B(CARRYB_7__0_), .CI(SUMB_7__1_), .CO(
        CARRYB_8__0_), .S(A1_6_) );
  ADDFHX4 S1_9_0 ( .A(ab_9__0_), .B(CARRYB_8__0_), .CI(SUMB_8__1_), .CO(
        CARRYB_9__0_), .S(A1_7_) );
  ADDFHX4 S2_10_4 ( .A(ab_10__4_), .B(CARRYB_9__4_), .CI(SUMB_9__5_), .CO(
        CARRYB_10__4_), .S(SUMB_10__4_) );
  ADDFHX4 S2_11_4 ( .A(ab_11__4_), .B(CARRYB_10__4_), .CI(SUMB_10__5_), .CO(
        CARRYB_11__4_), .S(SUMB_11__4_) );
  ADDFHX4 S2_10_3 ( .A(ab_10__3_), .B(CARRYB_9__3_), .CI(SUMB_9__4_), .CO(
        CARRYB_10__3_), .S(SUMB_10__3_) );
  ADDFHX4 S2_13_2 ( .A(ab_13__2_), .B(CARRYB_12__2_), .CI(SUMB_12__3_), .CO(
        CARRYB_13__2_), .S(SUMB_13__2_) );
  ADDFHX4 S2_14_2 ( .A(ab_14__2_), .B(CARRYB_13__2_), .CI(SUMB_13__3_), .CO(
        CARRYB_14__2_), .S(SUMB_14__2_) );
  ADDFHX4 S2_14_1 ( .A(ab_14__1_), .B(CARRYB_13__1_), .CI(SUMB_13__2_), .CO(
        CARRYB_14__1_), .S(SUMB_14__1_) );
  ADDFHX4 S4_4 ( .A(ab_16__4_), .B(CARRYB_15__4_), .CI(SUMB_15__5_), .CO(
        CARRYB_16__4_), .S(SUMB_16__4_) );
  ADDFHX4 S4_3 ( .A(ab_16__3_), .B(CARRYB_15__3_), .CI(SUMB_15__4_), .CO(
        CARRYB_16__3_), .S(SUMB_16__3_) );
  ADDFHX4 S2_9_1 ( .A(ab_9__1_), .B(CARRYB_8__1_), .CI(SUMB_8__2_), .CO(
        CARRYB_9__1_), .S(SUMB_9__1_) );
  ADDFHX4 S2_8_1 ( .A(ab_8__1_), .B(CARRYB_7__1_), .CI(SUMB_7__2_), .CO(
        CARRYB_8__1_), .S(SUMB_8__1_) );
  ADDFHX4 S2_11_1 ( .A(ab_11__1_), .B(CARRYB_10__1_), .CI(SUMB_10__2_), .CO(
        CARRYB_11__1_), .S(SUMB_11__1_) );
  ADDFHX4 S2_10_2 ( .A(ab_10__2_), .B(CARRYB_9__2_), .CI(SUMB_9__3_), .CO(
        CARRYB_10__2_), .S(SUMB_10__2_) );
  ADDFHX4 S2_11_2 ( .A(ab_11__2_), .B(CARRYB_10__2_), .CI(SUMB_10__3_), .CO(
        CARRYB_11__2_), .S(SUMB_11__2_) );
  ADDFHX4 S2_10_1 ( .A(ab_10__1_), .B(CARRYB_9__1_), .CI(SUMB_9__2_), .CO(
        CARRYB_10__1_), .S(SUMB_10__1_) );
  ADDFHX4 S2_8_2 ( .A(ab_8__2_), .B(CARRYB_7__2_), .CI(SUMB_7__3_), .CO(
        CARRYB_8__2_), .S(SUMB_8__2_) );
  ADDFHX4 S2_12_3 ( .A(ab_12__3_), .B(CARRYB_11__3_), .CI(SUMB_11__4_), .CO(
        CARRYB_12__3_), .S(SUMB_12__3_) );
  ADDFHX4 S2_14_3 ( .A(ab_14__3_), .B(CARRYB_13__3_), .CI(SUMB_13__4_), .CO(
        CARRYB_14__3_), .S(SUMB_14__3_) );
  ADDFHX4 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  ADDFHX4 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  ADDFHX4 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  ADDFHX4 S3_7_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(
        CARRYB_7__6_), .S(SUMB_7__6_) );
  ADDFHX4 S3_9_6 ( .A(ab_9__6_), .B(CARRYB_8__6_), .CI(ab_8__7_), .CO(
        CARRYB_9__6_), .S(SUMB_9__6_) );
  ADDFHX4 S2_7_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  ADDFHX4 S2_8_5 ( .A(ab_8__5_), .B(CARRYB_7__5_), .CI(SUMB_7__6_), .CO(
        CARRYB_8__5_), .S(SUMB_8__5_) );
  ADDFHX4 S2_9_5 ( .A(ab_9__5_), .B(CARRYB_8__5_), .CI(SUMB_8__6_), .CO(
        CARRYB_9__5_), .S(SUMB_9__5_) );
  ADDFHX4 S2_10_5 ( .A(ab_10__5_), .B(CARRYB_9__5_), .CI(SUMB_9__6_), .CO(
        CARRYB_10__5_), .S(SUMB_10__5_) );
  ADDFHX4 S2_7_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  ADDFHX4 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  ADDFHX4 S1_12_0 ( .A(ab_12__0_), .B(CARRYB_11__0_), .CI(SUMB_11__1_), .CO(
        CARRYB_12__0_), .S(A1_10_) );
  ADDFHX4 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  ADDFHX4 S2_7_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  ADDFHX4 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  ADDFHX4 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  ADDFHX4 S1_7_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(PROD1_7_) );
  ADDFHX4 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  ADDFHX4 S2_7_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  ADDFHX4 S2_9_4 ( .A(ab_9__4_), .B(CARRYB_8__4_), .CI(SUMB_8__5_), .CO(
        CARRYB_9__4_), .S(SUMB_9__4_) );
  ADDFHX4 S3_8_6 ( .A(ab_8__6_), .B(CARRYB_7__6_), .CI(ab_7__7_), .CO(
        CARRYB_8__6_), .S(SUMB_8__6_) );
  ADDFHX4 S4_5 ( .A(ab_16__5_), .B(CARRYB_15__5_), .CI(SUMB_15__6_), .CO(
        CARRYB_16__5_), .S(SUMB_16__5_) );
  ADDFHX4 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  ADDFHX4 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  ADDFHX4 S1_13_0 ( .A(ab_13__0_), .B(CARRYB_12__0_), .CI(SUMB_12__1_), .CO(
        CARRYB_13__0_), .S(A1_11_) );
  ADDFHX4 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  ADDFHX4 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  ADDFHX4 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  ADDFHX4 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  ADDFHX4 S2_12_5 ( .A(ab_12__5_), .B(CARRYB_11__5_), .CI(SUMB_11__6_), .CO(
        CARRYB_12__5_), .S(SUMB_12__5_) );
  ADDFHX4 S2_13_5 ( .A(ab_13__5_), .B(CARRYB_12__5_), .CI(SUMB_12__6_), .CO(
        CARRYB_13__5_), .S(SUMB_13__5_) );
  ADDFHX4 S2_2_5 ( .A(ab_2__5_), .B(n10), .CI(SUMB_1__6_), .CO(CARRYB_2__5_), 
        .S(SUMB_2__5_) );
  ADDFHX4 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  ADDFHX4 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  ADDFHX4 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  ADDFHX4 S2_12_1 ( .A(ab_12__1_), .B(CARRYB_11__1_), .CI(SUMB_11__2_), .CO(
        CARRYB_12__1_), .S(SUMB_12__1_) );
  ADDFHX4 S4_2 ( .A(ab_16__2_), .B(CARRYB_15__2_), .CI(SUMB_15__3_), .CO(
        CARRYB_16__2_), .S(SUMB_16__2_) );
  ADDFHX4 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  ADDFHX4 S2_7_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  ADDFHX4 S2_11_3 ( .A(ab_11__3_), .B(CARRYB_10__3_), .CI(SUMB_10__4_), .CO(
        CARRYB_11__3_), .S(SUMB_11__3_) );
  ADDFHX4 S2_15_3 ( .A(ab_15__3_), .B(CARRYB_14__3_), .CI(SUMB_14__4_), .CO(
        CARRYB_15__3_), .S(SUMB_15__3_) );
  ADDFHX4 S3_12_6 ( .A(ab_12__6_), .B(CARRYB_11__6_), .CI(ab_11__7_), .CO(
        CARRYB_12__6_), .S(SUMB_12__6_) );
  ADDFHX4 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  ADDFHX4 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  ADDFHX4 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  ADDFHX4 S3_10_6 ( .A(ab_10__6_), .B(CARRYB_9__6_), .CI(ab_9__7_), .CO(
        CARRYB_10__6_), .S(SUMB_10__6_) );
  ADDFHX4 S3_11_6 ( .A(ab_11__6_), .B(CARRYB_10__6_), .CI(ab_10__7_), .CO(
        CARRYB_11__6_), .S(SUMB_11__6_) );
  ADDFHX4 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  ADDFHX4 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  ADDFHX4 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  ADDFHX4 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  ADDFHX4 S2_13_3 ( .A(ab_13__3_), .B(CARRYB_12__3_), .CI(SUMB_12__4_), .CO(
        CARRYB_13__3_), .S(SUMB_13__3_) );
  ADDFHX4 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  ADDFHX4 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  ADDFHX4 S2_14_5 ( .A(ab_14__5_), .B(CARRYB_13__5_), .CI(SUMB_13__6_), .CO(
        CARRYB_14__5_), .S(SUMB_14__5_) );
  ADDFHX4 S2_15_4 ( .A(ab_15__4_), .B(CARRYB_14__4_), .CI(SUMB_14__5_), .CO(
        CARRYB_15__4_), .S(SUMB_15__4_) );
  ADDFHX4 S2_14_4 ( .A(ab_14__4_), .B(CARRYB_13__4_), .CI(SUMB_13__5_), .CO(
        CARRYB_14__4_), .S(SUMB_14__4_) );
  ADDFHX4 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  ADDFHX4 S3_13_6 ( .A(ab_13__6_), .B(CARRYB_12__6_), .CI(ab_12__7_), .CO(
        CARRYB_13__6_), .S(SUMB_13__6_) );
  ADDFHX2 S3_14_6 ( .A(ab_14__6_), .B(CARRYB_13__6_), .CI(ab_13__7_), .CO(
        CARRYB_14__6_), .S(SUMB_14__6_) );
  ADDFHX4 S3_2_6 ( .A(ab_2__6_), .B(n4), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  ADDFHX4 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  ADDFHX4 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  ADDFHX4 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  ADDFHX4 S2_2_3 ( .A(ab_2__3_), .B(n11), .CI(SUMB_1__4_), .CO(CARRYB_2__3_), 
        .S(SUMB_2__3_) );
  ADDFHX4 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  ADDFHX2 S2_15_5 ( .A(ab_15__5_), .B(CARRYB_14__5_), .CI(SUMB_14__6_), .CO(
        CARRYB_15__5_), .S(SUMB_15__5_) );
  ADDFHX2 S3_15_6 ( .A(ab_15__6_), .B(CARRYB_14__6_), .CI(ab_14__7_), .CO(
        CARRYB_15__6_), .S(SUMB_15__6_) );
  ADDFHX4 S5_6 ( .A(ab_16__6_), .B(CARRYB_15__6_), .CI(ab_15__7_), .CO(
        CARRYB_16__6_), .S(SUMB_16__6_) );
  NAND2X2 U2 ( .A(ab_1__4_), .B(ab_0__5_), .Y(n18) );
  NOR2BX4 U3 ( .AN(ab_1__3_), .B(n3), .Y(n11) );
  CLKINVX20 U4 ( .A(ab_0__4_), .Y(n3) );
  XOR2X4 U5 ( .A(n43), .B(ab_0__2_), .Y(SUMB_1__1_) );
  AND2X4 U6 ( .A(ab_0__7_), .B(ab_1__6_), .Y(n4) );
  NOR2BX1 U7 ( .AN(A[5]), .B(n22), .Y(ab_5__5_) );
  NOR2BX2 U8 ( .AN(A[3]), .B(n31), .Y(ab_3__6_) );
  XOR2X2 U9 ( .A(ab_1__3_), .B(ab_0__4_), .Y(SUMB_1__3_) );
  AND2X4 U10 ( .A(A[1]), .B(B[3]), .Y(ab_1__3_) );
  NAND2X4 U11 ( .A(ab_1__2_), .B(ab_0__3_), .Y(n21) );
  NAND2X4 U12 ( .A(n43), .B(ab_0__2_), .Y(n20) );
  NOR2BX4 U13 ( .AN(n12), .B(n39), .Y(ab_2__3_) );
  INVX8 U14 ( .A(ab_0__3_), .Y(n7) );
  NOR2BX4 U15 ( .AN(B[3]), .B(n34), .Y(ab_0__3_) );
  INVX4 U16 ( .A(B[4]), .Y(n38) );
  NOR2BX1 U17 ( .AN(A[10]), .B(n23), .Y(ab_10__5_) );
  NOR2BX1 U18 ( .AN(A[14]), .B(n25), .Y(ab_14__4_) );
  NOR2BX2 U19 ( .AN(A[8]), .B(n22), .Y(ab_8__5_) );
  NOR2BX2 U20 ( .AN(A[8]), .B(n24), .Y(ab_8__4_) );
  NOR2BX1 U21 ( .AN(A[14]), .B(n28), .Y(ab_14__2_) );
  NOR2BX1 U22 ( .AN(A[12]), .B(n23), .Y(ab_12__5_) );
  NOR2BX1 U23 ( .AN(A[10]), .B(n25), .Y(ab_10__4_) );
  NOR2BX1 U24 ( .AN(A[10]), .B(n26), .Y(ab_10__3_) );
  NOR2BXL U25 ( .AN(A[16]), .B(n28), .Y(ab_16__2_) );
  NOR2BXL U26 ( .AN(A[16]), .B(n26), .Y(ab_16__3_) );
  INVX4 U27 ( .A(n20), .Y(CARRYB_1__1_) );
  INVX4 U28 ( .A(n21), .Y(CARRYB_1__2_) );
  NOR2BX2 U29 ( .AN(A[13]), .B(n33), .Y(ab_13__0_) );
  NOR2BXL U30 ( .AN(A[16]), .B(n25), .Y(ab_16__4_) );
  AND2X2 U32 ( .A(CARRYB_16__5_), .B(SUMB_16__6_), .Y(n6) );
  INVX3 U33 ( .A(B[3]), .Y(n39) );
  BUFX3 U34 ( .A(n39), .Y(n26) );
  CLKINVX2 U35 ( .A(A[1]), .Y(n8) );
  NOR2X4 U36 ( .A(n36), .B(n34), .Y(ab_0__6_) );
  XNOR2X4 U37 ( .A(ab_1__2_), .B(n7), .Y(SUMB_1__2_) );
  AND3X4 U38 ( .A(n9), .B(B[1]), .C(n35), .Y(CARRYB_1__0_) );
  CLKINVX4 U39 ( .A(n8), .Y(n9) );
  NOR2BX2 U40 ( .AN(A[3]), .B(n22), .Y(ab_3__5_) );
  NOR2BX2 U41 ( .AN(n9), .B(n42), .Y(ab_1__7_) );
  NOR2BX4 U42 ( .AN(n12), .B(n22), .Y(ab_2__5_) );
  NOR2BX2 U43 ( .AN(A[6]), .B(n24), .Y(ab_6__4_) );
  NOR2BX4 U44 ( .AN(n12), .B(n24), .Y(ab_2__4_) );
  BUFX16 U45 ( .A(A[2]), .Y(n12) );
  XOR2X4 U46 ( .A(CARRYB_16__5_), .B(SUMB_16__6_), .Y(A1_20_) );
  NOR2BX4 U47 ( .AN(n12), .B(n29), .Y(ab_2__1_) );
  AND2X4 U48 ( .A(SUMB_16__3_), .B(CARRYB_16__2_), .Y(n14) );
  XOR2X4 U49 ( .A(ab_1__6_), .B(ab_0__7_), .Y(SUMB_1__6_) );
  AND2X4 U50 ( .A(ab_0__6_), .B(ab_1__5_), .Y(n10) );
  NOR2BX4 U51 ( .AN(B[4]), .B(n34), .Y(ab_0__4_) );
  NOR2BXL U52 ( .AN(A[0]), .B(n32), .Y(n35) );
  INVX16 U53 ( .A(B[0]), .Y(n32) );
  INVX8 U54 ( .A(A[0]), .Y(n34) );
  INVX8 U55 ( .A(B[1]), .Y(n41) );
  NOR2BX2 U56 ( .AN(A[3]), .B(n32), .Y(ab_3__0_) );
  NOR2BX1 U57 ( .AN(A[5]), .B(n27), .Y(ab_5__2_) );
  BUFX20 U58 ( .A(n37), .Y(n22) );
  NOR2BX2 U59 ( .AN(A[3]), .B(n39), .Y(ab_3__3_) );
  NOR2BX2 U60 ( .AN(A[3]), .B(n27), .Y(ab_3__2_) );
  NOR2BX2 U61 ( .AN(A[3]), .B(n24), .Y(ab_3__4_) );
  NOR2BX2 U62 ( .AN(A[3]), .B(n29), .Y(ab_3__1_) );
  INVX4 U63 ( .A(n18), .Y(CARRYB_1__4_) );
  NAND2X4 U64 ( .A(CARRYB_16__0_), .B(SUMB_16__1_), .Y(n19) );
  INVX8 U65 ( .A(B[6]), .Y(n36) );
  INVX4 U66 ( .A(B[2]), .Y(n40) );
  XOR2X4 U67 ( .A(ab_1__5_), .B(ab_0__6_), .Y(SUMB_1__5_) );
  INVX8 U68 ( .A(B[5]), .Y(n37) );
  NOR2BX1 U69 ( .AN(A[3]), .B(n42), .Y(ab_3__7_) );
  XOR2X4 U70 ( .A(ab_1__4_), .B(ab_0__5_), .Y(SUMB_1__4_) );
  INVX8 U71 ( .A(n19), .Y(A2_16_) );
  NOR2BX4 U72 ( .AN(n13), .B(n34), .Y(ab_0__7_) );
  NOR2BX2 U73 ( .AN(n12), .B(n32), .Y(ab_2__0_) );
  NOR2BX4 U74 ( .AN(B[2]), .B(n34), .Y(ab_0__2_) );
  BUFX8 U75 ( .A(B[7]), .Y(n13) );
  INVX16 U76 ( .A(n13), .Y(n42) );
  NOR2BX4 U77 ( .AN(A[1]), .B(n29), .Y(n43) );
  NOR2BX4 U78 ( .AN(A[1]), .B(n27), .Y(ab_1__2_) );
  XOR2X4 U79 ( .A(CARRYB_16__0_), .B(SUMB_16__1_), .Y(A1_15_) );
  NOR2BX4 U80 ( .AN(A[1]), .B(n22), .Y(ab_1__5_) );
  NOR2BX4 U81 ( .AN(n12), .B(n27), .Y(ab_2__2_) );
  AND2X4 U82 ( .A(A[1]), .B(B[6]), .Y(ab_1__6_) );
  AND2X2 U83 ( .A(CARRYB_16__3_), .B(SUMB_16__4_), .Y(n15) );
  XOR2X4 U84 ( .A(SUMB_16__4_), .B(CARRYB_16__3_), .Y(A1_18_) );
  NOR2BXL U85 ( .AN(A[7]), .B(n22), .Y(ab_7__5_) );
  NOR2BX1 U86 ( .AN(A[4]), .B(n29), .Y(ab_4__1_) );
  NOR2BX1 U87 ( .AN(A[4]), .B(n22), .Y(ab_4__5_) );
  NOR2BX1 U88 ( .AN(A[8]), .B(n32), .Y(ab_8__0_) );
  NOR2BX1 U89 ( .AN(A[8]), .B(n39), .Y(ab_8__3_) );
  NOR2BXL U90 ( .AN(A[11]), .B(n31), .Y(ab_11__6_) );
  NOR2BX1 U91 ( .AN(A[8]), .B(n31), .Y(ab_8__6_) );
  NOR2BXL U92 ( .AN(A[14]), .B(n31), .Y(ab_14__6_) );
  NOR2BX2 U93 ( .AN(A[4]), .B(n31), .Y(ab_4__6_) );
  NOR2BX1 U94 ( .AN(A[9]), .B(n23), .Y(ab_9__5_) );
  NOR2BX1 U95 ( .AN(A[7]), .B(n27), .Y(ab_7__2_) );
  NOR2BX1 U96 ( .AN(A[6]), .B(n32), .Y(ab_6__0_) );
  NOR2BX1 U97 ( .AN(A[7]), .B(n32), .Y(ab_7__0_) );
  NOR2BX1 U98 ( .AN(A[6]), .B(n27), .Y(ab_6__2_) );
  NOR2BX1 U99 ( .AN(A[4]), .B(n39), .Y(ab_4__3_) );
  NOR2BX1 U100 ( .AN(A[8]), .B(n27), .Y(ab_8__2_) );
  NOR2BX1 U101 ( .AN(A[6]), .B(n31), .Y(ab_6__6_) );
  BUFX16 U102 ( .A(n36), .Y(n31) );
  INVXL U103 ( .A(B[0]), .Y(n33) );
  AND2X4 U104 ( .A(CARRYB_16__1_), .B(SUMB_16__2_), .Y(n16) );
  NOR2BXL U105 ( .AN(A[7]), .B(n24), .Y(ab_7__4_) );
  NOR2BX1 U106 ( .AN(A[14]), .B(n26), .Y(ab_14__3_) );
  NOR2BX1 U107 ( .AN(A[12]), .B(n26), .Y(ab_12__3_) );
  NOR2BXL U108 ( .AN(A[6]), .B(n22), .Y(ab_6__5_) );
  NOR2BX1 U109 ( .AN(A[6]), .B(n26), .Y(ab_6__3_) );
  NOR2BXL U110 ( .AN(A[5]), .B(n24), .Y(ab_5__4_) );
  NOR2BX1 U111 ( .AN(A[12]), .B(n28), .Y(ab_12__2_) );
  NOR2BX1 U112 ( .AN(A[12]), .B(n25), .Y(ab_12__4_) );
  NOR2BXL U113 ( .AN(A[10]), .B(n32), .Y(ab_10__0_) );
  NOR2BX1 U114 ( .AN(A[14]), .B(n30), .Y(ab_14__1_) );
  NOR2BX1 U115 ( .AN(A[10]), .B(n30), .Y(ab_10__1_) );
  NOR2BX1 U116 ( .AN(A[10]), .B(n28), .Y(ab_10__2_) );
  NOR2BX1 U117 ( .AN(A[12]), .B(n30), .Y(ab_12__1_) );
  CLKBUFXL U118 ( .A(n38), .Y(n25) );
  BUFX8 U119 ( .A(n41), .Y(n29) );
  NOR2BX1 U120 ( .AN(A[15]), .B(n25), .Y(ab_15__4_) );
  NOR2BX4 U121 ( .AN(n12), .B(n31), .Y(ab_2__6_) );
  NOR2BX1 U122 ( .AN(A[10]), .B(n31), .Y(ab_10__6_) );
  NOR2BX1 U123 ( .AN(A[6]), .B(n42), .Y(ab_6__7_) );
  NOR2BX1 U124 ( .AN(A[14]), .B(n42), .Y(ab_14__7_) );
  NOR2BX1 U125 ( .AN(A[15]), .B(n33), .Y(ab_15__0_) );
  CLKBUFXL U126 ( .A(n40), .Y(n28) );
  CLKBUFXL U127 ( .A(n41), .Y(n30) );
  NOR2BX1 U128 ( .AN(A[11]), .B(n26), .Y(ab_11__3_) );
  NOR2BX1 U129 ( .AN(A[9]), .B(n25), .Y(ab_9__4_) );
  NOR2BX1 U130 ( .AN(A[5]), .B(n29), .Y(ab_5__1_) );
  NOR2BX1 U131 ( .AN(A[13]), .B(n23), .Y(ab_13__5_) );
  NOR2BXL U132 ( .AN(A[12]), .B(n32), .Y(ab_12__0_) );
  NOR2BX2 U133 ( .AN(A[14]), .B(n23), .Y(ab_14__5_) );
  NOR2BX1 U134 ( .AN(A[14]), .B(n33), .Y(ab_14__0_) );
  NOR2BX1 U135 ( .AN(A[13]), .B(n30), .Y(ab_13__1_) );
  NOR2BX2 U136 ( .AN(A[6]), .B(n29), .Y(ab_6__1_) );
  NOR2BX1 U137 ( .AN(A[5]), .B(n39), .Y(ab_5__3_) );
  NOR2BX1 U138 ( .AN(A[4]), .B(n24), .Y(ab_4__4_) );
  NOR2BX1 U139 ( .AN(A[13]), .B(n28), .Y(ab_13__2_) );
  NOR2BX1 U140 ( .AN(A[11]), .B(n28), .Y(ab_11__2_) );
  NOR2BX1 U141 ( .AN(A[13]), .B(n26), .Y(ab_13__3_) );
  NOR2BXL U142 ( .AN(A[9]), .B(n32), .Y(ab_9__0_) );
  NOR2BX1 U143 ( .AN(A[11]), .B(n25), .Y(ab_11__4_) );
  NOR2BX1 U144 ( .AN(A[9]), .B(n28), .Y(ab_9__2_) );
  NOR2BX1 U145 ( .AN(A[9]), .B(n26), .Y(ab_9__3_) );
  NOR2BX1 U146 ( .AN(A[9]), .B(n30), .Y(ab_9__1_) );
  NOR2BX1 U147 ( .AN(A[8]), .B(n29), .Y(ab_8__1_) );
  NOR2BX1 U148 ( .AN(A[7]), .B(n29), .Y(ab_7__1_) );
  NOR2BX1 U149 ( .AN(A[7]), .B(n39), .Y(ab_7__3_) );
  NOR2BX1 U150 ( .AN(A[4]), .B(n27), .Y(ab_4__2_) );
  NOR2BX1 U151 ( .AN(A[11]), .B(n30), .Y(ab_11__1_) );
  NOR2BXL U152 ( .AN(A[11]), .B(n32), .Y(ab_11__0_) );
  NOR2BX1 U153 ( .AN(A[13]), .B(n25), .Y(ab_13__4_) );
  NOR2BX1 U154 ( .AN(A[11]), .B(n23), .Y(ab_11__5_) );
  BUFX12 U155 ( .A(n38), .Y(n24) );
  AND2X2 U156 ( .A(CARRYB_16__4_), .B(SUMB_16__5_), .Y(n17) );
  XOR2X1 U157 ( .A(CARRYB_16__6_), .B(ab_16__7_), .Y(A1_21_) );
  BUFX3 U158 ( .A(n37), .Y(n23) );
  NOR2BX1 U159 ( .AN(A[16]), .B(n23), .Y(ab_16__5_) );
  NOR2BX1 U160 ( .AN(A[16]), .B(n31), .Y(ab_16__6_) );
  NOR2BX1 U161 ( .AN(A[15]), .B(n42), .Y(ab_15__7_) );
  NOR2BXL U162 ( .AN(A[5]), .B(n42), .Y(ab_5__7_) );
  NOR2BXL U163 ( .AN(A[11]), .B(n42), .Y(ab_11__7_) );
  NOR2BX2 U164 ( .AN(A[12]), .B(n31), .Y(ab_12__6_) );
  NOR2BXL U165 ( .AN(A[4]), .B(n42), .Y(ab_4__7_) );
  NOR2BX1 U166 ( .AN(A[5]), .B(n31), .Y(ab_5__6_) );
  NOR2BXL U167 ( .AN(A[10]), .B(n42), .Y(ab_10__7_) );
  NOR2BX1 U168 ( .AN(A[16]), .B(n30), .Y(ab_16__1_) );
  NOR2BX1 U169 ( .AN(A[16]), .B(n33), .Y(ab_16__0_) );
  NOR2BXL U170 ( .AN(A[13]), .B(n42), .Y(ab_13__7_) );
  NOR2BX1 U171 ( .AN(A[15]), .B(n31), .Y(ab_15__6_) );
  NOR2BXL U172 ( .AN(A[12]), .B(n42), .Y(ab_12__7_) );
  NOR2BX1 U173 ( .AN(A[13]), .B(n31), .Y(ab_13__6_) );
  NOR2BX1 U174 ( .AN(n12), .B(n42), .Y(ab_2__7_) );
  NOR2BX1 U175 ( .AN(A[15]), .B(n30), .Y(ab_15__1_) );
  NOR2BXL U176 ( .AN(A[8]), .B(n42), .Y(ab_8__7_) );
  NOR2BX1 U177 ( .AN(A[9]), .B(n31), .Y(ab_9__6_) );
  NOR2BXL U178 ( .AN(A[7]), .B(n42), .Y(ab_7__7_) );
  NOR2BX1 U179 ( .AN(A[15]), .B(n28), .Y(ab_15__2_) );
  NOR2BXL U180 ( .AN(A[5]), .B(n32), .Y(ab_5__0_) );
  NOR2BX2 U181 ( .AN(A[4]), .B(n32), .Y(ab_4__0_) );
  NOR2BXL U182 ( .AN(A[9]), .B(n42), .Y(ab_9__7_) );
  BUFX12 U183 ( .A(n40), .Y(n27) );
  NOR2BXL U184 ( .AN(A[15]), .B(n23), .Y(ab_15__5_) );
  NOR2BX1 U185 ( .AN(A[7]), .B(n31), .Y(ab_7__6_) );
  NOR2BX1 U186 ( .AN(A[15]), .B(n26), .Y(ab_15__3_) );
  NOR2BXL U187 ( .AN(A[16]), .B(n42), .Y(ab_16__7_) );
  XOR2X4 U188 ( .A(CARRYB_16__4_), .B(SUMB_16__5_), .Y(A1_19_) );
  XOR2X4 U189 ( .A(SUMB_16__2_), .B(CARRYB_16__1_), .Y(A1_16_) );
  XOR2X4 U190 ( .A(SUMB_16__3_), .B(CARRYB_16__2_), .Y(A1_17_) );
  NOR2BX4 U191 ( .AN(B[5]), .B(n34), .Y(ab_0__5_) );
  NOR2BX4 U192 ( .AN(A[1]), .B(n24), .Y(ab_1__4_) );
endmodule


module multi16_11 ( in_17bit, in_8bit, out );
  input [16:0] in_17bit;
  input [7:0] in_8bit;
  output [16:0] out;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122;
  wire   [15:1] in_17bit_b;
  wire   [7:1] in_8bit_b;
  wire   [23:8] mul;

  multi16_11_DW02_mult_0 mult_55 ( .A({n12, in_17bit_b[15:2], n46, n23}), .B({
        in_8bit_b, n49}), .PRODUCT_23_(mul[23]), .PRODUCT_22_(mul[22]), 
        .PRODUCT_21_(mul[21]), .PRODUCT_20_(mul[20]), .PRODUCT_19_(mul[19]), 
        .PRODUCT_18_(mul[18]), .PRODUCT_17_(mul[17]), .PRODUCT_16_(mul[16]), 
        .PRODUCT_15_(mul[15]), .PRODUCT_14_(mul[14]), .PRODUCT_13_(mul[13]), 
        .PRODUCT_12_(mul[12]), .PRODUCT_11_(mul[11]), .PRODUCT_10_(mul[10]), 
        .PRODUCT_9_(mul[9]), .PRODUCT_8_(mul[8]), .PRODUCT_7_(out[0]) );
  OR2X4 U2 ( .A(mul[17]), .B(n8), .Y(n3) );
  INVXL U3 ( .A(n112), .Y(n1) );
  CLKINVX8 U4 ( .A(n19), .Y(n20) );
  INVX2 U5 ( .A(mul[20]), .Y(n19) );
  OR2X4 U6 ( .A(in_8bit[1]), .B(in_8bit[2]), .Y(n52) );
  INVX2 U7 ( .A(in_8bit[2]), .Y(n48) );
  NOR2XL U8 ( .A(n39), .B(n93), .Y(n70) );
  CLKINVX4 U9 ( .A(n93), .Y(n5) );
  OR2X2 U10 ( .A(n44), .B(n93), .Y(n38) );
  AND2X2 U11 ( .A(n47), .B(n66), .Y(n34) );
  BUFX16 U12 ( .A(in_17bit_b[1]), .Y(n46) );
  OR3X1 U13 ( .A(in_17bit[15]), .B(n94), .C(n93), .Y(n2) );
  NAND2X4 U14 ( .A(n18), .B(n4), .Y(n15) );
  OR2X4 U15 ( .A(in_17bit[1]), .B(in_17bit[0]), .Y(n4) );
  AOI21X4 U16 ( .A0(n116), .A1(n112), .B0(n119), .Y(n117) );
  CLKINVX3 U17 ( .A(n57), .Y(n13) );
  CLKINVX2 U18 ( .A(n106), .Y(n11) );
  INVX1 U19 ( .A(n83), .Y(n85) );
  NAND2X2 U20 ( .A(n42), .B(n87), .Y(n88) );
  CLKINVX2 U21 ( .A(in_17bit[5]), .Y(n69) );
  INVX8 U22 ( .A(in_17bit[4]), .Y(n67) );
  XNOR2X2 U23 ( .A(mul[8]), .B(n24), .Y(out[1]) );
  OR2X2 U24 ( .A(mul[8]), .B(out[0]), .Y(n96) );
  NAND2BX2 U25 ( .AN(mul[16]), .B(n11), .Y(n8) );
  OAI21X2 U26 ( .A0(n49), .A1(n52), .B0(in_8bit[7]), .Y(n51) );
  NOR2X4 U27 ( .A(in_17bit[1]), .B(in_17bit[0]), .Y(n6) );
  AOI2BB1X4 U28 ( .A0N(mul[19]), .A1N(n7), .B0(n119), .Y(n113) );
  OR2X4 U29 ( .A(n3), .B(mul[18]), .Y(n7) );
  BUFX20 U30 ( .A(in_8bit[0]), .Y(n49) );
  AND2X1 U31 ( .A(n47), .B(n68), .Y(n29) );
  CLKINVX8 U32 ( .A(n56), .Y(n58) );
  NOR2X4 U33 ( .A(mul[21]), .B(n118), .Y(n116) );
  CLKINVX4 U34 ( .A(in_8bit[5]), .Y(n57) );
  XNOR2X4 U35 ( .A(n70), .B(n71), .Y(in_17bit_b[6]) );
  XNOR2X2 U36 ( .A(in_8bit[1]), .B(n35), .Y(in_8bit_b[1]) );
  OR2X4 U37 ( .A(mul[12]), .B(n99), .Y(n100) );
  INVX2 U38 ( .A(n53), .Y(n9) );
  CLKINVX8 U39 ( .A(n9), .Y(n10) );
  INVXL U40 ( .A(in_8bit[3]), .Y(n53) );
  NAND2XL U41 ( .A(n5), .B(n72), .Y(n30) );
  AND3X4 U42 ( .A(in_17bit[1]), .B(n47), .C(in_17bit[0]), .Y(n63) );
  NAND2BX4 U43 ( .AN(mul[16]), .B(n11), .Y(n108) );
  CLKINVX4 U44 ( .A(n2), .Y(n12) );
  XOR2X4 U45 ( .A(mul[23]), .B(n122), .Y(out[16]) );
  AOI21X2 U46 ( .A0(n120), .A1(n121), .B0(n119), .Y(n122) );
  NOR2XL U47 ( .A(n42), .B(n93), .Y(n86) );
  NOR2XL U48 ( .A(n82), .B(n93), .Y(n80) );
  NOR2XL U49 ( .A(n43), .B(n93), .Y(n75) );
  XOR2X4 U50 ( .A(n112), .B(n111), .Y(out[12]) );
  BUFX20 U51 ( .A(in_17bit[16]), .Y(n47) );
  NAND2X4 U52 ( .A(n44), .B(n67), .Y(n68) );
  NAND2X4 U53 ( .A(n49), .B(in_8bit[7]), .Y(n35) );
  INVX8 U54 ( .A(in_17bit[2]), .Y(n65) );
  XOR2X4 U55 ( .A(n14), .B(n13), .Y(in_8bit_b[5]) );
  NOR2X4 U56 ( .A(n58), .B(n61), .Y(n14) );
  OR2X4 U57 ( .A(n47), .B(in_17bit[1]), .Y(n18) );
  NOR2X4 U58 ( .A(n15), .B(n63), .Y(in_17bit_b[1]) );
  OR2X4 U59 ( .A(mul[14]), .B(n102), .Y(n103) );
  NOR2X2 U60 ( .A(mul[20]), .B(n21), .Y(n16) );
  NOR3X2 U61 ( .A(n49), .B(n37), .C(n52), .Y(n17) );
  NOR2X2 U62 ( .A(n17), .B(n61), .Y(n54) );
  NAND2X4 U63 ( .A(n62), .B(in_8bit[7]), .Y(n60) );
  XOR2X4 U64 ( .A(n50), .B(n48), .Y(in_8bit_b[2]) );
  OAI21X2 U65 ( .A0(in_8bit[1]), .A1(n49), .B0(in_8bit[7]), .Y(n50) );
  XNOR2X4 U66 ( .A(n69), .B(n29), .Y(in_17bit_b[5]) );
  INVX8 U67 ( .A(mul[19]), .Y(n112) );
  XNOR2X4 U68 ( .A(n64), .B(n65), .Y(in_17bit_b[2]) );
  NAND2X4 U69 ( .A(n6), .B(n65), .Y(n66) );
  INVX8 U70 ( .A(n47), .Y(n93) );
  OR2X4 U71 ( .A(n3), .B(mul[18]), .Y(n21) );
  OR2X4 U72 ( .A(n21), .B(mul[20]), .Y(n118) );
  XOR2X4 U73 ( .A(n51), .B(n10), .Y(in_8bit_b[3]) );
  NOR3X4 U74 ( .A(in_8bit[6]), .B(n62), .C(n61), .Y(in_8bit_b[7]) );
  NOR2XL U75 ( .A(n1), .B(n118), .Y(n120) );
  NAND2X4 U76 ( .A(n39), .B(n71), .Y(n72) );
  NOR2X4 U77 ( .A(n68), .B(in_17bit[5]), .Y(n39) );
  INVX4 U78 ( .A(in_17bit[0]), .Y(n22) );
  CLKINVX4 U79 ( .A(n22), .Y(n23) );
  AOI21X4 U80 ( .A0(n16), .A1(n112), .B0(n119), .Y(n115) );
  OR2X4 U81 ( .A(mul[17]), .B(n8), .Y(n114) );
  XOR2X4 U82 ( .A(n113), .B(n20), .Y(out[13]) );
  XNOR2X2 U83 ( .A(mul[12]), .B(n27), .Y(out[5]) );
  NAND2X2 U84 ( .A(n99), .B(n110), .Y(n27) );
  XNOR2X4 U85 ( .A(mul[15]), .B(n31), .Y(out[8]) );
  OR2X4 U86 ( .A(mul[13]), .B(n100), .Y(n102) );
  NOR2X4 U87 ( .A(in_17bit[3]), .B(n66), .Y(n44) );
  XOR2X4 U88 ( .A(n38), .B(n67), .Y(in_17bit_b[4]) );
  NAND2X4 U89 ( .A(n58), .B(n57), .Y(n62) );
  NAND2XL U90 ( .A(n82), .B(n81), .Y(n83) );
  INVX2 U91 ( .A(in_17bit[6]), .Y(n71) );
  OR2X4 U92 ( .A(mul[9]), .B(n96), .Y(n97) );
  INVXL U93 ( .A(in_17bit[7]), .Y(n73) );
  XOR2X2 U94 ( .A(mul[11]), .B(n25), .Y(out[4]) );
  NAND2XL U95 ( .A(n5), .B(n77), .Y(n32) );
  NOR2XL U96 ( .A(n88), .B(in_17bit[13]), .Y(n41) );
  NAND2X2 U97 ( .A(n41), .B(n91), .Y(n94) );
  NAND2X4 U98 ( .A(n103), .B(n110), .Y(n31) );
  XNOR2X2 U99 ( .A(mul[10]), .B(n28), .Y(out[3]) );
  NAND2X2 U100 ( .A(n97), .B(n110), .Y(n28) );
  AND2X2 U101 ( .A(n98), .B(n110), .Y(n25) );
  OR2X4 U102 ( .A(mul[11]), .B(n98), .Y(n99) );
  INVX4 U103 ( .A(n10), .Y(n37) );
  XNOR2X4 U104 ( .A(mul[9]), .B(n95), .Y(out[2]) );
  NAND2X4 U105 ( .A(n96), .B(n110), .Y(n95) );
  NAND2XL U106 ( .A(out[0]), .B(n110), .Y(n24) );
  XNOR2X4 U107 ( .A(mul[13]), .B(n26), .Y(out[6]) );
  NAND2X4 U108 ( .A(n100), .B(n110), .Y(n26) );
  XOR2X2 U109 ( .A(n73), .B(n30), .Y(in_17bit_b[7]) );
  XOR2X2 U110 ( .A(n78), .B(n32), .Y(in_17bit_b[9]) );
  NAND2BXL U111 ( .AN(n77), .B(n78), .Y(n79) );
  AND2X4 U112 ( .A(n74), .B(n73), .Y(n43) );
  XOR2X2 U113 ( .A(n89), .B(n33), .Y(in_17bit_b[13]) );
  NAND2XL U114 ( .A(n5), .B(n88), .Y(n33) );
  AND2X4 U115 ( .A(n85), .B(n84), .Y(n42) );
  XOR2X4 U116 ( .A(in_17bit[3]), .B(n34), .Y(in_17bit_b[3]) );
  INVX4 U117 ( .A(in_17bit[8]), .Y(n76) );
  INVX4 U118 ( .A(n119), .Y(n110) );
  OR2X2 U119 ( .A(mul[10]), .B(n97), .Y(n98) );
  NOR3X4 U120 ( .A(n49), .B(n37), .C(n52), .Y(n36) );
  NOR2XL U121 ( .A(n41), .B(n93), .Y(n90) );
  XNOR2X2 U122 ( .A(n84), .B(n40), .Y(in_17bit_b[11]) );
  AND2X1 U123 ( .A(n5), .B(n83), .Y(n40) );
  NOR2XL U124 ( .A(mul[22]), .B(mul[21]), .Y(n121) );
  XNOR2X2 U125 ( .A(n92), .B(n45), .Y(in_17bit_b[15]) );
  AND2X1 U126 ( .A(n94), .B(n5), .Y(n45) );
  INVXL U127 ( .A(in_17bit[9]), .Y(n78) );
  INVXL U128 ( .A(in_17bit[12]), .Y(n87) );
  INVXL U129 ( .A(in_17bit[10]), .Y(n81) );
  INVXL U130 ( .A(in_17bit[11]), .Y(n84) );
  INVXL U131 ( .A(in_17bit[14]), .Y(n91) );
  INVXL U132 ( .A(in_17bit[13]), .Y(n89) );
  INVXL U133 ( .A(in_8bit[6]), .Y(n59) );
  XNOR2X1 U134 ( .A(n47), .B(in_8bit[7]), .Y(n119) );
  INVX1 U135 ( .A(in_8bit[7]), .Y(n61) );
  INVX1 U136 ( .A(in_8bit[4]), .Y(n55) );
  XNOR2X4 U137 ( .A(mul[18]), .B(n109), .Y(out[11]) );
  OAI21X2 U138 ( .A0(mul[18]), .A1(n3), .B0(n110), .Y(n111) );
  XNOR2X4 U139 ( .A(n54), .B(n55), .Y(in_8bit_b[4]) );
  NAND2X4 U140 ( .A(n55), .B(n36), .Y(n56) );
  XOR2X4 U141 ( .A(n60), .B(n59), .Y(in_8bit_b[6]) );
  NOR2X4 U142 ( .A(n93), .B(n6), .Y(n64) );
  CLKINVX3 U143 ( .A(n72), .Y(n74) );
  XNOR2X4 U144 ( .A(n75), .B(n76), .Y(in_17bit_b[8]) );
  NAND2X4 U145 ( .A(n43), .B(n76), .Y(n77) );
  CLKINVX3 U146 ( .A(n79), .Y(n82) );
  XNOR2X4 U147 ( .A(n80), .B(n81), .Y(in_17bit_b[10]) );
  XNOR2X4 U148 ( .A(n86), .B(n87), .Y(in_17bit_b[12]) );
  XNOR2X4 U149 ( .A(n90), .B(n91), .Y(in_17bit_b[14]) );
  CLKINVX3 U150 ( .A(in_17bit[15]), .Y(n92) );
  NAND2X4 U151 ( .A(n102), .B(n110), .Y(n101) );
  XNOR2X4 U152 ( .A(mul[14]), .B(n101), .Y(out[7]) );
  CLKINVX3 U153 ( .A(n103), .Y(n104) );
  NAND2BX4 U154 ( .AN(mul[15]), .B(n104), .Y(n106) );
  NAND2X4 U155 ( .A(n106), .B(n110), .Y(n105) );
  XNOR2X4 U156 ( .A(mul[16]), .B(n105), .Y(out[9]) );
  NAND2X4 U157 ( .A(n108), .B(n110), .Y(n107) );
  XNOR2X4 U158 ( .A(mul[17]), .B(n107), .Y(out[10]) );
  NAND2X4 U159 ( .A(n114), .B(n110), .Y(n109) );
  XOR2X4 U160 ( .A(n115), .B(mul[21]), .Y(out[14]) );
  XOR2X4 U161 ( .A(n117), .B(mul[22]), .Y(out[15]) );
endmodule


module multi16_10_DW01_add_0 ( A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, 
        A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, 
        B_20_, B_19_, B_18_, B_17_, B_16_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, 
        SUM_17_, SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, 
        SUM_9_, SUM_8_, SUM_7_, SUM_6_, SUM_5_ );
  input A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_,
         A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, B_20_, B_19_,
         B_18_, B_17_, B_16_;
  output SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, SUM_15_,
         SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, SUM_7_,
         SUM_6_, SUM_5_;
  wire   n1, n2, n3, n4, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40;

  OR2X4 U2 ( .A(A_17_), .B(B_17_), .Y(n1) );
  AOI21X1 U3 ( .A0(n24), .A1(n25), .B0(n16), .Y(n23) );
  NOR2X4 U4 ( .A(B_19_), .B(A_19_), .Y(n28) );
  XOR2X4 U5 ( .A(n2), .B(n24), .Y(SUM_20_) );
  AND2X4 U6 ( .A(n26), .B(n25), .Y(n2) );
  BUFX16 U7 ( .A(A_5_), .Y(SUM_5_) );
  NAND2BX4 U8 ( .AN(n18), .B(n17), .Y(n39) );
  INVX2 U9 ( .A(n33), .Y(n18) );
  AOI21X4 U10 ( .A0(n20), .A1(n1), .B0(n19), .Y(n3) );
  AOI21X2 U11 ( .A0(n20), .A1(n1), .B0(n19), .Y(n38) );
  OR2X2 U12 ( .A(B_20_), .B(A_20_), .Y(n25) );
  INVX8 U13 ( .A(n21), .Y(SUM_15_) );
  CLKINVX8 U14 ( .A(n34), .Y(n20) );
  XOR2X1 U15 ( .A(n22), .B(n23), .Y(SUM_21_) );
  NOR2BX4 U16 ( .AN(n29), .B(n28), .Y(n37) );
  BUFX12 U17 ( .A(A_14_), .Y(SUM_14_) );
  BUFX8 U18 ( .A(A_10_), .Y(SUM_10_) );
  NAND2X4 U19 ( .A(A_16_), .B(B_16_), .Y(n34) );
  CLKINVX8 U20 ( .A(A_15_), .Y(n21) );
  OAI21X4 U21 ( .A0(n27), .A1(n28), .B0(n29), .Y(n24) );
  NAND2X4 U22 ( .A(B_18_), .B(A_18_), .Y(n33) );
  NAND2X4 U23 ( .A(B_19_), .B(A_19_), .Y(n29) );
  AND2X4 U24 ( .A(n4), .B(n34), .Y(SUM_16_) );
  OAI21X1 U25 ( .A0(n30), .A1(n34), .B0(n35), .Y(n32) );
  INVXL U26 ( .A(n26), .Y(n16) );
  INVX4 U27 ( .A(n31), .Y(n17) );
  OR2X4 U28 ( .A(A_16_), .B(B_16_), .Y(n4) );
  AOI21X2 U29 ( .A0(n17), .A1(n32), .B0(n18), .Y(n27) );
  BUFX4 U30 ( .A(A_9_), .Y(SUM_9_) );
  BUFX4 U31 ( .A(A_7_), .Y(SUM_7_) );
  BUFX8 U32 ( .A(A_8_), .Y(SUM_8_) );
  BUFX4 U33 ( .A(A_6_), .Y(SUM_6_) );
  BUFX8 U34 ( .A(A_13_), .Y(SUM_13_) );
  BUFX8 U35 ( .A(A_12_), .Y(SUM_12_) );
  BUFX8 U36 ( .A(A_11_), .Y(SUM_11_) );
  OAI21X2 U37 ( .A0(n38), .A1(n31), .B0(n33), .Y(n36) );
  NOR2X4 U38 ( .A(B_18_), .B(A_18_), .Y(n31) );
  NAND2X4 U39 ( .A(A_17_), .B(B_17_), .Y(n35) );
  NOR2X4 U40 ( .A(n19), .B(n30), .Y(n40) );
  INVX8 U41 ( .A(n35), .Y(n19) );
  XOR2X4 U42 ( .A(n36), .B(n37), .Y(SUM_19_) );
  XOR2X4 U43 ( .A(n40), .B(n20), .Y(SUM_17_) );
  NOR2X4 U44 ( .A(A_17_), .B(B_17_), .Y(n30) );
  XOR2X4 U45 ( .A(n39), .B(n3), .Y(SUM_18_) );
  XNOR2X1 U46 ( .A(B_21_), .B(A_21_), .Y(n22) );
  NAND2X1 U47 ( .A(B_20_), .B(A_20_), .Y(n26) );
endmodule


module multi16_10_DW02_mult_0 ( A, B, PRODUCT_23_, PRODUCT_22_, PRODUCT_21_, 
        PRODUCT_20_, PRODUCT_19_, PRODUCT_18_, PRODUCT_17_, PRODUCT_16_, 
        PRODUCT_15_, PRODUCT_14_, PRODUCT_13_, PRODUCT_12_, PRODUCT_11_, 
        PRODUCT_10_, PRODUCT_9_, PRODUCT_8_, PRODUCT_7_ );
  input [16:0] A;
  input [7:0] B;
  output PRODUCT_23_, PRODUCT_22_, PRODUCT_21_, PRODUCT_20_, PRODUCT_19_,
         PRODUCT_18_, PRODUCT_17_, PRODUCT_16_, PRODUCT_15_, PRODUCT_14_,
         PRODUCT_13_, PRODUCT_12_, PRODUCT_11_, PRODUCT_10_, PRODUCT_9_,
         PRODUCT_8_, PRODUCT_7_;
  wire   ab_16__7_, ab_16__6_, ab_16__5_, ab_16__4_, ab_16__3_, ab_16__2_,
         ab_16__1_, ab_16__0_, ab_15__7_, ab_15__6_, ab_15__5_, ab_15__4_,
         ab_15__3_, ab_15__2_, ab_15__1_, ab_15__0_, ab_14__7_, ab_14__6_,
         ab_14__5_, ab_14__4_, ab_14__3_, ab_14__2_, ab_14__1_, ab_14__0_,
         ab_13__7_, ab_13__6_, ab_13__5_, ab_13__4_, ab_13__3_, ab_13__2_,
         ab_13__1_, ab_13__0_, ab_12__7_, ab_12__6_, ab_12__5_, ab_12__4_,
         ab_12__3_, ab_12__2_, ab_12__1_, ab_12__0_, ab_11__7_, ab_11__6_,
         ab_11__5_, ab_11__4_, ab_11__3_, ab_11__2_, ab_11__1_, ab_11__0_,
         ab_10__7_, ab_10__6_, ab_10__5_, ab_10__4_, ab_10__3_, ab_10__2_,
         ab_10__1_, ab_10__0_, ab_9__7_, ab_9__6_, ab_9__5_, ab_9__4_,
         ab_9__3_, ab_9__2_, ab_9__1_, ab_9__0_, ab_8__7_, ab_8__6_, ab_8__5_,
         ab_8__4_, ab_8__3_, ab_8__2_, ab_8__1_, ab_8__0_, ab_7__7_, ab_7__6_,
         ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_, ab_7__0_, ab_6__7_,
         ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_, ab_6__1_, ab_6__0_,
         ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_, ab_5__2_, ab_5__1_,
         ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_, ab_4__3_, ab_4__2_,
         ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_, ab_3__4_, ab_3__3_,
         ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_, ab_2__5_, ab_2__4_,
         ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_, ab_1__6_, ab_1__5_,
         ab_1__4_, ab_1__3_, ab_1__2_, ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_,
         ab_0__3_, ab_0__2_, CARRYB_16__6_, CARRYB_16__5_, CARRYB_16__4_,
         CARRYB_16__3_, CARRYB_16__2_, CARRYB_16__1_, CARRYB_16__0_,
         CARRYB_15__6_, CARRYB_15__5_, CARRYB_15__4_, CARRYB_15__3_,
         CARRYB_15__2_, CARRYB_15__1_, CARRYB_15__0_, CARRYB_14__6_,
         CARRYB_14__5_, CARRYB_14__4_, CARRYB_14__3_, CARRYB_14__2_,
         CARRYB_14__1_, CARRYB_14__0_, CARRYB_13__6_, CARRYB_13__5_,
         CARRYB_13__4_, CARRYB_13__3_, CARRYB_13__2_, CARRYB_13__1_,
         CARRYB_13__0_, CARRYB_12__6_, CARRYB_12__5_, CARRYB_12__4_,
         CARRYB_12__3_, CARRYB_12__2_, CARRYB_12__1_, CARRYB_12__0_,
         CARRYB_11__6_, CARRYB_11__5_, CARRYB_11__4_, CARRYB_11__3_,
         CARRYB_11__2_, CARRYB_11__1_, CARRYB_11__0_, CARRYB_10__6_,
         CARRYB_10__5_, CARRYB_10__4_, CARRYB_10__3_, CARRYB_10__2_,
         CARRYB_10__1_, CARRYB_10__0_, CARRYB_9__6_, CARRYB_9__5_,
         CARRYB_9__4_, CARRYB_9__3_, CARRYB_9__2_, CARRYB_9__1_, CARRYB_9__0_,
         CARRYB_8__6_, CARRYB_8__5_, CARRYB_8__4_, CARRYB_8__3_, CARRYB_8__2_,
         CARRYB_8__1_, CARRYB_8__0_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_,
         CARRYB_7__3_, CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_,
         CARRYB_6__5_, CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_,
         CARRYB_6__0_, CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_,
         CARRYB_5__2_, CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_,
         CARRYB_4__4_, CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_,
         CARRYB_3__6_, CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_,
         CARRYB_3__1_, CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_,
         CARRYB_2__3_, CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__6_,
         CARRYB_1__3_, CARRYB_1__0_, SUMB_16__6_, SUMB_16__5_, SUMB_16__4_,
         SUMB_16__3_, SUMB_16__2_, SUMB_16__1_, SUMB_16__0_, SUMB_15__6_,
         SUMB_15__5_, SUMB_15__4_, SUMB_15__3_, SUMB_15__2_, SUMB_15__1_,
         SUMB_14__6_, SUMB_14__5_, SUMB_14__4_, SUMB_14__3_, SUMB_14__2_,
         SUMB_14__1_, SUMB_13__6_, SUMB_13__5_, SUMB_13__4_, SUMB_13__3_,
         SUMB_13__2_, SUMB_13__1_, SUMB_12__6_, SUMB_12__5_, SUMB_12__4_,
         SUMB_12__3_, SUMB_12__2_, SUMB_12__1_, SUMB_11__6_, SUMB_11__5_,
         SUMB_11__4_, SUMB_11__3_, SUMB_11__2_, SUMB_11__1_, SUMB_10__6_,
         SUMB_10__5_, SUMB_10__4_, SUMB_10__3_, SUMB_10__2_, SUMB_10__1_,
         SUMB_9__6_, SUMB_9__5_, SUMB_9__4_, SUMB_9__3_, SUMB_9__2_,
         SUMB_9__1_, SUMB_8__6_, SUMB_8__5_, SUMB_8__4_, SUMB_8__3_,
         SUMB_8__2_, SUMB_8__1_, SUMB_7__6_, SUMB_7__5_, SUMB_7__4_,
         SUMB_7__3_, SUMB_7__2_, SUMB_7__1_, SUMB_6__6_, SUMB_6__5_,
         SUMB_6__4_, SUMB_6__3_, SUMB_6__2_, SUMB_6__1_, SUMB_5__6_,
         SUMB_5__5_, SUMB_5__4_, SUMB_5__3_, SUMB_5__2_, SUMB_5__1_,
         SUMB_4__6_, SUMB_4__5_, SUMB_4__4_, SUMB_4__3_, SUMB_4__2_,
         SUMB_4__1_, SUMB_3__6_, SUMB_3__5_, SUMB_3__4_, SUMB_3__3_,
         SUMB_3__2_, SUMB_3__1_, SUMB_2__6_, SUMB_2__5_, SUMB_2__4_,
         SUMB_2__3_, SUMB_2__2_, SUMB_2__1_, SUMB_1__6_, SUMB_1__5_,
         SUMB_1__4_, SUMB_1__3_, SUMB_1__2_, SUMB_1__1_, PROD1_7_, A1_21_,
         A1_20_, A1_19_, A1_18_, A1_17_, A1_16_, A1_15_, A1_13_, A1_12_,
         A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, A1_4_, A1_3_, A1_2_,
         A1_1_, A1_0_, n3, n4, n5, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47;

  multi16_10_DW01_add_0 FS_1 ( .A_21_(A1_21_), .A_20_(A1_20_), .A_19_(A1_19_), 
        .A_18_(A1_18_), .A_17_(A1_17_), .A_16_(A1_16_), .A_15_(A1_15_), 
        .A_14_(SUMB_16__0_), .A_13_(A1_13_), .A_12_(A1_12_), .A_11_(A1_11_), 
        .A_10_(A1_10_), .A_9_(A1_9_), .A_8_(A1_8_), .A_7_(A1_7_), .A_6_(A1_6_), 
        .A_5_(PROD1_7_), .B_21_(n19), .B_20_(n23), .B_19_(n22), .B_18_(n3), 
        .B_17_(n7), .B_16_(n21), .SUM_21_(PRODUCT_23_), .SUM_20_(PRODUCT_22_), 
        .SUM_19_(PRODUCT_21_), .SUM_18_(PRODUCT_20_), .SUM_17_(PRODUCT_19_), 
        .SUM_16_(PRODUCT_18_), .SUM_15_(PRODUCT_17_), .SUM_14_(PRODUCT_16_), 
        .SUM_13_(PRODUCT_15_), .SUM_12_(PRODUCT_14_), .SUM_11_(PRODUCT_13_), 
        .SUM_10_(PRODUCT_12_), .SUM_9_(PRODUCT_11_), .SUM_8_(PRODUCT_10_), 
        .SUM_7_(PRODUCT_9_), .SUM_6_(PRODUCT_8_), .SUM_5_(PRODUCT_7_) );
  ADDFHX4 S4_3 ( .A(ab_16__3_), .B(CARRYB_15__3_), .CI(SUMB_15__4_), .CO(
        CARRYB_16__3_), .S(SUMB_16__3_) );
  ADDFHX4 S2_9_4 ( .A(ab_9__4_), .B(CARRYB_8__4_), .CI(SUMB_8__5_), .CO(
        CARRYB_9__4_), .S(SUMB_9__4_) );
  ADDFHX4 S2_11_2 ( .A(ab_11__2_), .B(CARRYB_10__2_), .CI(SUMB_10__3_), .CO(
        CARRYB_11__2_), .S(SUMB_11__2_) );
  ADDFHX4 S2_12_2 ( .A(ab_12__2_), .B(CARRYB_11__2_), .CI(SUMB_11__3_), .CO(
        CARRYB_12__2_), .S(SUMB_12__2_) );
  ADDFHX4 S2_14_3 ( .A(ab_14__3_), .B(CARRYB_13__3_), .CI(SUMB_13__4_), .CO(
        CARRYB_14__3_), .S(SUMB_14__3_) );
  ADDFHX4 S2_8_3 ( .A(ab_8__3_), .B(CARRYB_7__3_), .CI(SUMB_7__4_), .CO(
        CARRYB_8__3_), .S(SUMB_8__3_) );
  ADDFHX4 S2_9_3 ( .A(ab_9__3_), .B(CARRYB_8__3_), .CI(SUMB_8__4_), .CO(
        CARRYB_9__3_), .S(SUMB_9__3_) );
  ADDFHX4 S2_10_4 ( .A(ab_10__4_), .B(CARRYB_9__4_), .CI(SUMB_9__5_), .CO(
        CARRYB_10__4_), .S(SUMB_10__4_) );
  ADDFHX4 S2_11_4 ( .A(ab_11__4_), .B(CARRYB_10__4_), .CI(SUMB_10__5_), .CO(
        CARRYB_11__4_), .S(SUMB_11__4_) );
  ADDFHX4 S4_0 ( .A(ab_16__0_), .B(CARRYB_15__0_), .CI(SUMB_15__1_), .CO(
        CARRYB_16__0_), .S(SUMB_16__0_) );
  ADDFHX4 S1_10_0 ( .A(ab_10__0_), .B(CARRYB_9__0_), .CI(SUMB_9__1_), .CO(
        CARRYB_10__0_), .S(A1_8_) );
  ADDFHX4 S1_11_0 ( .A(ab_11__0_), .B(CARRYB_10__0_), .CI(SUMB_10__1_), .CO(
        CARRYB_11__0_), .S(A1_9_) );
  ADDFHX4 S2_9_1 ( .A(ab_9__1_), .B(CARRYB_8__1_), .CI(SUMB_8__2_), .CO(
        CARRYB_9__1_), .S(SUMB_9__1_) );
  ADDFHX4 S2_9_2 ( .A(ab_9__2_), .B(CARRYB_8__2_), .CI(SUMB_8__3_), .CO(
        CARRYB_9__2_), .S(SUMB_9__2_) );
  ADDFHX4 S2_10_2 ( .A(ab_10__2_), .B(CARRYB_9__2_), .CI(SUMB_9__3_), .CO(
        CARRYB_10__2_), .S(SUMB_10__2_) );
  ADDFHX4 S2_15_1 ( .A(ab_15__1_), .B(CARRYB_14__1_), .CI(SUMB_14__2_), .CO(
        CARRYB_15__1_), .S(SUMB_15__1_) );
  ADDFHX4 S4_1 ( .A(ab_16__1_), .B(CARRYB_15__1_), .CI(SUMB_15__2_), .CO(
        CARRYB_16__1_), .S(SUMB_16__1_) );
  ADDFHX4 S2_8_1 ( .A(ab_8__1_), .B(CARRYB_7__1_), .CI(SUMB_7__2_), .CO(
        CARRYB_8__1_), .S(SUMB_8__1_) );
  ADDFHX4 S3_15_6 ( .A(ab_15__6_), .B(CARRYB_14__6_), .CI(ab_14__7_), .CO(
        CARRYB_15__6_), .S(SUMB_15__6_) );
  ADDFHX4 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  ADDFHX4 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  ADDFHX4 S4_2 ( .A(ab_16__2_), .B(CARRYB_15__2_), .CI(SUMB_15__3_), .CO(
        CARRYB_16__2_), .S(SUMB_16__2_) );
  ADDFHX4 S2_12_5 ( .A(ab_12__5_), .B(CARRYB_11__5_), .CI(SUMB_11__6_), .CO(
        CARRYB_12__5_), .S(SUMB_12__5_) );
  ADDFHX4 S3_13_6 ( .A(ab_13__6_), .B(CARRYB_12__6_), .CI(ab_12__7_), .CO(
        CARRYB_13__6_), .S(SUMB_13__6_) );
  ADDFHX4 S3_14_6 ( .A(ab_14__6_), .B(CARRYB_13__6_), .CI(ab_13__7_), .CO(
        CARRYB_14__6_), .S(SUMB_14__6_) );
  ADDFHX4 S2_11_5 ( .A(ab_11__5_), .B(SUMB_10__6_), .CI(CARRYB_10__5_), .CO(
        CARRYB_11__5_), .S(SUMB_11__5_) );
  ADDFHX4 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  ADDFHX4 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  ADDFHX4 S2_8_2 ( .A(ab_8__2_), .B(CARRYB_7__2_), .CI(SUMB_7__3_), .CO(
        CARRYB_8__2_), .S(SUMB_8__2_) );
  ADDFHX4 S3_11_6 ( .A(ab_11__6_), .B(CARRYB_10__6_), .CI(ab_10__7_), .CO(
        CARRYB_11__6_), .S(SUMB_11__6_) );
  ADDFHX4 S3_12_6 ( .A(ab_12__6_), .B(CARRYB_11__6_), .CI(ab_11__7_), .CO(
        CARRYB_12__6_), .S(SUMB_12__6_) );
  ADDFHX4 S2_15_5 ( .A(ab_15__5_), .B(CARRYB_14__5_), .CI(SUMB_14__6_), .CO(
        CARRYB_15__5_), .S(SUMB_15__5_) );
  ADDFHX4 S4_4 ( .A(ab_16__4_), .B(CARRYB_15__4_), .CI(SUMB_15__5_), .CO(
        CARRYB_16__4_), .S(SUMB_16__4_) );
  ADDFHX4 S2_7_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  ADDFHX4 S1_8_0 ( .A(ab_8__0_), .B(CARRYB_7__0_), .CI(SUMB_7__1_), .CO(
        CARRYB_8__0_), .S(A1_6_) );
  ADDFHX4 S1_9_0 ( .A(ab_9__0_), .B(CARRYB_8__0_), .CI(SUMB_8__1_), .CO(
        CARRYB_9__0_), .S(A1_7_) );
  ADDFHX4 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  ADDFHX4 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  ADDFHX4 S2_7_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  ADDFHX4 S2_8_4 ( .A(ab_8__4_), .B(CARRYB_7__4_), .CI(SUMB_7__5_), .CO(
        CARRYB_8__4_), .S(SUMB_8__4_) );
  ADDFHX4 S3_10_6 ( .A(ab_10__6_), .B(CARRYB_9__6_), .CI(ab_9__7_), .CO(
        CARRYB_10__6_), .S(SUMB_10__6_) );
  ADDFHX4 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  ADDFHX4 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  ADDFHX4 S2_15_2 ( .A(ab_15__2_), .B(CARRYB_14__2_), .CI(SUMB_14__3_), .CO(
        CARRYB_15__2_), .S(SUMB_15__2_) );
  ADDFHX4 S2_13_2 ( .A(ab_13__2_), .B(CARRYB_12__2_), .CI(SUMB_12__3_), .CO(
        CARRYB_13__2_), .S(SUMB_13__2_) );
  ADDFHX4 S2_14_2 ( .A(ab_14__2_), .B(CARRYB_13__2_), .CI(SUMB_13__3_), .CO(
        CARRYB_14__2_), .S(SUMB_14__2_) );
  ADDFHX4 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  ADDFHX4 S2_11_1 ( .A(ab_11__1_), .B(CARRYB_10__1_), .CI(SUMB_10__2_), .CO(
        CARRYB_11__1_), .S(SUMB_11__1_) );
  ADDFHX4 S2_12_1 ( .A(ab_12__1_), .B(CARRYB_11__1_), .CI(SUMB_11__2_), .CO(
        CARRYB_12__1_), .S(SUMB_12__1_) );
  ADDFHX4 S1_13_0 ( .A(ab_13__0_), .B(CARRYB_12__0_), .CI(SUMB_12__1_), .CO(
        CARRYB_13__0_), .S(A1_11_) );
  ADDFHX4 S1_14_0 ( .A(ab_14__0_), .B(CARRYB_13__0_), .CI(SUMB_13__1_), .CO(
        CARRYB_14__0_), .S(A1_12_) );
  ADDFHX4 S2_7_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  ADDFHX4 S3_9_6 ( .A(ab_9__6_), .B(CARRYB_8__6_), .CI(ab_8__7_), .CO(
        CARRYB_9__6_), .S(SUMB_9__6_) );
  ADDFHX4 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  ADDFHX4 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  ADDFHX4 S2_12_3 ( .A(ab_12__3_), .B(CARRYB_11__3_), .CI(SUMB_11__4_), .CO(
        CARRYB_12__3_), .S(SUMB_12__3_) );
  ADDFHX4 S2_2_2 ( .A(ab_2__2_), .B(n9), .CI(SUMB_1__3_), .CO(CARRYB_2__2_), 
        .S(SUMB_2__2_) );
  ADDFHX4 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  ADDFHX4 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  ADDFHX4 S2_13_1 ( .A(ab_13__1_), .B(CARRYB_12__1_), .CI(SUMB_12__2_), .CO(
        CARRYB_13__1_), .S(SUMB_13__1_) );
  ADDFHX4 S2_14_1 ( .A(ab_14__1_), .B(CARRYB_13__1_), .CI(SUMB_13__2_), .CO(
        CARRYB_14__1_), .S(SUMB_14__1_) );
  ADDFHX4 S2_10_1 ( .A(ab_10__1_), .B(CARRYB_9__1_), .CI(SUMB_9__2_), .CO(
        CARRYB_10__1_), .S(SUMB_10__1_) );
  ADDFHX4 S2_8_5 ( .A(ab_8__5_), .B(CARRYB_7__5_), .CI(SUMB_7__6_), .CO(
        CARRYB_8__5_), .S(SUMB_8__5_) );
  ADDFHX4 S3_7_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(
        CARRYB_7__6_), .S(SUMB_7__6_) );
  ADDFHX4 S3_8_6 ( .A(ab_8__6_), .B(CARRYB_7__6_), .CI(ab_7__7_), .CO(
        CARRYB_8__6_), .S(SUMB_8__6_) );
  ADDFHX4 S2_2_3 ( .A(CARRYB_1__3_), .B(ab_2__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  ADDFHX4 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  ADDFHX4 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  ADDFHX4 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  ADDFHX4 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  ADDFHX4 S1_7_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(PROD1_7_) );
  ADDFHX4 S2_2_1 ( .A(ab_2__1_), .B(n5), .CI(SUMB_1__2_), .CO(CARRYB_2__1_), 
        .S(SUMB_2__1_) );
  ADDFHX4 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  ADDFHX4 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  ADDFHX4 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  ADDFHX4 S2_7_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  ADDFHX4 S2_9_5 ( .A(ab_9__5_), .B(CARRYB_8__5_), .CI(SUMB_8__6_), .CO(
        CARRYB_9__5_), .S(SUMB_9__5_) );
  ADDFHX4 S2_7_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  ADDFHX4 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  ADDFHX4 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  ADDFHX4 S2_10_3 ( .A(ab_10__3_), .B(CARRYB_9__3_), .CI(SUMB_9__4_), .CO(
        CARRYB_10__3_), .S(SUMB_10__3_) );
  ADDFHX4 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  ADDFHX4 S1_12_0 ( .A(ab_12__0_), .B(CARRYB_11__0_), .CI(SUMB_11__1_), .CO(
        CARRYB_12__0_), .S(A1_10_) );
  ADDFHX4 S1_15_0 ( .A(ab_15__0_), .B(CARRYB_14__0_), .CI(SUMB_14__1_), .CO(
        CARRYB_15__0_), .S(A1_13_) );
  ADDFHX4 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  ADDFHX4 S2_13_4 ( .A(ab_13__4_), .B(CARRYB_12__4_), .CI(SUMB_12__5_), .CO(
        CARRYB_13__4_), .S(SUMB_13__4_) );
  ADDFHX4 S2_11_3 ( .A(ab_11__3_), .B(CARRYB_10__3_), .CI(SUMB_10__4_), .CO(
        CARRYB_11__3_), .S(SUMB_11__3_) );
  ADDFHX4 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  ADDFHX4 S2_12_4 ( .A(ab_12__4_), .B(CARRYB_11__4_), .CI(SUMB_11__5_), .CO(
        CARRYB_12__4_), .S(SUMB_12__4_) );
  ADDFHX4 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  ADDFHX4 S3_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(ab_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  ADDFHX4 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  ADDFHX4 S2_13_3 ( .A(ab_13__3_), .B(CARRYB_12__3_), .CI(SUMB_12__4_), .CO(
        CARRYB_13__3_), .S(SUMB_13__3_) );
  ADDFHX4 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  ADDFHX4 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  ADDFHX4 S2_14_4 ( .A(ab_14__4_), .B(CARRYB_13__4_), .CI(SUMB_13__5_), .CO(
        CARRYB_14__4_), .S(SUMB_14__4_) );
  ADDFHX4 S2_15_3 ( .A(ab_15__3_), .B(CARRYB_14__3_), .CI(SUMB_14__4_), .CO(
        CARRYB_15__3_), .S(SUMB_15__3_) );
  ADDFHX4 S2_13_5 ( .A(ab_13__5_), .B(CARRYB_12__5_), .CI(SUMB_12__6_), .CO(
        CARRYB_13__5_), .S(SUMB_13__5_) );
  ADDFHX4 S2_14_5 ( .A(ab_14__5_), .B(CARRYB_13__5_), .CI(SUMB_13__6_), .CO(
        CARRYB_14__5_), .S(SUMB_14__5_) );
  ADDFHX4 S2_15_4 ( .A(ab_15__4_), .B(CARRYB_14__4_), .CI(SUMB_14__5_), .CO(
        CARRYB_15__4_), .S(SUMB_15__4_) );
  ADDFHX4 S5_6 ( .A(ab_16__6_), .B(CARRYB_15__6_), .CI(ab_15__7_), .CO(
        CARRYB_16__6_), .S(SUMB_16__6_) );
  ADDFHX2 S2_10_5 ( .A(ab_10__5_), .B(CARRYB_9__5_), .CI(SUMB_9__6_), .CO(
        CARRYB_10__5_), .S(SUMB_10__5_) );
  ADDFHX2 S2_2_5 ( .A(ab_2__5_), .B(n8), .CI(SUMB_1__6_), .CO(CARRYB_2__5_), 
        .S(SUMB_2__5_) );
  ADDFHX2 S2_2_4 ( .A(ab_2__4_), .B(n10), .CI(SUMB_1__5_), .CO(CARRYB_2__4_), 
        .S(SUMB_2__4_) );
  BUFX8 U2 ( .A(n20), .Y(n3) );
  AND2X4 U3 ( .A(A[1]), .B(B[2]), .Y(ab_1__2_) );
  BUFX20 U4 ( .A(n43), .Y(n32) );
  AND3X2 U5 ( .A(A[1]), .B(B[1]), .C(n38), .Y(CARRYB_1__0_) );
  AND2X4 U6 ( .A(A[1]), .B(B[3]), .Y(n4) );
  NOR2BX4 U7 ( .AN(A[2]), .B(n40), .Y(ab_2__5_) );
  AND2X4 U8 ( .A(n11), .B(B[6]), .Y(ab_1__6_) );
  NOR2BX4 U9 ( .AN(B[4]), .B(n37), .Y(ab_0__4_) );
  NOR2BX2 U10 ( .AN(A[5]), .B(n29), .Y(ab_5__4_) );
  AND2X4 U11 ( .A(ab_0__2_), .B(n47), .Y(n5) );
  NOR2BX1 U12 ( .AN(A[8]), .B(n28), .Y(ab_8__5_) );
  NOR2BX2 U13 ( .AN(A[8]), .B(n29), .Y(ab_8__4_) );
  NOR2BX1 U14 ( .AN(A[11]), .B(n30), .Y(ab_11__4_) );
  NOR2BXL U15 ( .AN(A[8]), .B(n42), .Y(ab_8__3_) );
  NOR2BXL U16 ( .AN(A[11]), .B(n28), .Y(ab_11__5_) );
  NOR2BX1 U17 ( .AN(A[12]), .B(n33), .Y(ab_12__2_) );
  NOR2BX2 U18 ( .AN(A[8]), .B(n32), .Y(ab_8__2_) );
  NOR2BX2 U19 ( .AN(A[8]), .B(n34), .Y(ab_8__1_) );
  NOR2BX2 U20 ( .AN(A[8]), .B(n36), .Y(ab_8__0_) );
  NOR2BXL U21 ( .AN(A[9]), .B(n28), .Y(ab_9__5_) );
  NOR2BX1 U22 ( .AN(A[9]), .B(n30), .Y(ab_9__4_) );
  NOR2BX1 U23 ( .AN(A[9]), .B(n31), .Y(ab_9__3_) );
  NOR2BX1 U24 ( .AN(A[13]), .B(n30), .Y(ab_13__4_) );
  NOR2BX1 U25 ( .AN(A[13]), .B(n33), .Y(ab_13__2_) );
  INVX4 U26 ( .A(B[4]), .Y(n41) );
  NOR2BX1 U27 ( .AN(A[9]), .B(n35), .Y(ab_9__1_) );
  NOR2BXL U28 ( .AN(A[13]), .B(n28), .Y(ab_13__5_) );
  BUFX20 U29 ( .A(n45), .Y(n36) );
  NOR2BX2 U30 ( .AN(A[5]), .B(n34), .Y(ab_5__1_) );
  NOR2BX2 U31 ( .AN(A[5]), .B(n27), .Y(ab_5__6_) );
  NOR2BXL U32 ( .AN(A[10]), .B(n28), .Y(ab_10__5_) );
  NOR2BX1 U33 ( .AN(A[10]), .B(n31), .Y(ab_10__3_) );
  NOR2BX1 U34 ( .AN(A[14]), .B(n33), .Y(ab_14__2_) );
  NOR2BX1 U35 ( .AN(A[14]), .B(n30), .Y(ab_14__4_) );
  NOR2BX1 U36 ( .AN(A[10]), .B(n35), .Y(ab_10__1_) );
  NOR2BXL U37 ( .AN(A[14]), .B(n28), .Y(ab_14__5_) );
  NOR2BX2 U38 ( .AN(A[5]), .B(n36), .Y(ab_5__0_) );
  NOR2BX2 U39 ( .AN(A[6]), .B(n34), .Y(ab_6__1_) );
  NOR2BX1 U40 ( .AN(A[7]), .B(n28), .Y(ab_7__5_) );
  NOR2BX2 U41 ( .AN(A[3]), .B(n40), .Y(ab_3__5_) );
  NOR2BX1 U42 ( .AN(A[12]), .B(n30), .Y(ab_12__4_) );
  NOR2BX1 U43 ( .AN(A[11]), .B(n31), .Y(ab_11__3_) );
  NOR2BXL U44 ( .AN(A[7]), .B(n42), .Y(ab_7__3_) );
  NOR2BX2 U45 ( .AN(A[7]), .B(n32), .Y(ab_7__2_) );
  NOR2BX1 U46 ( .AN(A[11]), .B(n33), .Y(ab_11__2_) );
  NOR2BXL U47 ( .AN(A[12]), .B(n28), .Y(ab_12__5_) );
  INVX1 U48 ( .A(n34), .Y(n14) );
  NOR2BX1 U49 ( .AN(A[11]), .B(n35), .Y(ab_11__1_) );
  NOR2BX2 U50 ( .AN(A[7]), .B(n34), .Y(ab_7__1_) );
  NOR2BX1 U51 ( .AN(A[16]), .B(n35), .Y(ab_16__1_) );
  NOR2BX1 U52 ( .AN(A[16]), .B(n33), .Y(ab_16__2_) );
  NOR2BX1 U53 ( .AN(A[16]), .B(n30), .Y(ab_16__4_) );
  NAND3X2 U54 ( .A(n18), .B(n16), .C(n17), .Y(CARRYB_16__5_) );
  NOR2BX2 U55 ( .AN(A[7]), .B(n36), .Y(ab_7__0_) );
  NOR2BX2 U56 ( .AN(A[6]), .B(n36), .Y(ab_6__0_) );
  INVX2 U58 ( .A(B[3]), .Y(n42) );
  BUFX3 U59 ( .A(n42), .Y(n31) );
  INVX4 U60 ( .A(B[5]), .Y(n40) );
  CLKBUFX2 U61 ( .A(n40), .Y(n28) );
  AND2X4 U62 ( .A(CARRYB_16__1_), .B(SUMB_16__2_), .Y(n7) );
  AND2X4 U63 ( .A(ab_1__5_), .B(ab_0__6_), .Y(n8) );
  AND2X4 U64 ( .A(ab_1__2_), .B(ab_0__3_), .Y(n9) );
  AND2X4 U65 ( .A(ab_0__5_), .B(ab_1__4_), .Y(n10) );
  CLKINVX4 U66 ( .A(B[0]), .Y(n45) );
  NOR2BX2 U67 ( .AN(A[3]), .B(n29), .Y(ab_3__4_) );
  BUFX8 U68 ( .A(n39), .Y(n27) );
  BUFX8 U69 ( .A(A[1]), .Y(n11) );
  NOR2BX4 U70 ( .AN(A[2]), .B(n36), .Y(ab_2__0_) );
  BUFX20 U71 ( .A(n39), .Y(n26) );
  INVX12 U72 ( .A(A[0]), .Y(n37) );
  XOR2X4 U73 ( .A(ab_1__4_), .B(ab_0__5_), .Y(SUMB_1__4_) );
  XOR2X4 U74 ( .A(ab_1__2_), .B(ab_0__3_), .Y(SUMB_1__2_) );
  NAND2X4 U75 ( .A(ab_0__4_), .B(ab_1__3_), .Y(n24) );
  AND2X4 U76 ( .A(B[7]), .B(A[0]), .Y(n12) );
  AND2X2 U77 ( .A(B[7]), .B(A[0]), .Y(ab_0__7_) );
  NOR2BX4 U78 ( .AN(n11), .B(n46), .Y(ab_1__7_) );
  AND2X2 U79 ( .A(CARRYB_16__2_), .B(SUMB_16__3_), .Y(n20) );
  NAND2X4 U80 ( .A(n13), .B(ab_0__7_), .Y(n25) );
  NOR2X4 U81 ( .A(n40), .B(n37), .Y(ab_0__5_) );
  AND2X4 U82 ( .A(A[1]), .B(B[3]), .Y(ab_1__3_) );
  XOR2X2 U83 ( .A(n47), .B(ab_0__2_), .Y(SUMB_1__1_) );
  NOR2BX2 U84 ( .AN(B[2]), .B(n37), .Y(ab_0__2_) );
  NOR2BX4 U85 ( .AN(n11), .B(n26), .Y(n13) );
  AND2X4 U86 ( .A(A[1]), .B(n14), .Y(n47) );
  NOR2BX2 U87 ( .AN(A[3]), .B(n36), .Y(ab_3__0_) );
  NOR2BX4 U88 ( .AN(A[2]), .B(n34), .Y(ab_2__1_) );
  NOR2BX4 U89 ( .AN(A[2]), .B(n29), .Y(ab_2__4_) );
  INVX4 U90 ( .A(n24), .Y(CARRYB_1__3_) );
  XOR2X4 U91 ( .A(ab_1__5_), .B(ab_0__6_), .Y(SUMB_1__5_) );
  NOR2BX4 U92 ( .AN(A[2]), .B(n32), .Y(ab_2__2_) );
  NOR2BX2 U93 ( .AN(A[9]), .B(n33), .Y(ab_9__2_) );
  INVX4 U94 ( .A(n25), .Y(CARRYB_1__6_) );
  NOR2BX2 U95 ( .AN(A[3]), .B(n34), .Y(ab_3__1_) );
  NOR2BX2 U96 ( .AN(A[4]), .B(n32), .Y(ab_4__2_) );
  NOR2BX2 U97 ( .AN(A[3]), .B(n42), .Y(ab_3__3_) );
  NOR2BX2 U98 ( .AN(A[3]), .B(n32), .Y(ab_3__2_) );
  NOR2BX2 U99 ( .AN(A[4]), .B(n42), .Y(ab_4__3_) );
  NOR2BX2 U100 ( .AN(B[3]), .B(n37), .Y(ab_0__3_) );
  INVX8 U101 ( .A(B[6]), .Y(n39) );
  NOR2BX4 U102 ( .AN(A[2]), .B(n42), .Y(ab_2__3_) );
  XOR2X4 U103 ( .A(ab_1__6_), .B(n12), .Y(SUMB_1__6_) );
  NOR2BX4 U104 ( .AN(B[6]), .B(n37), .Y(ab_0__6_) );
  NOR2BX2 U105 ( .AN(A[4]), .B(n34), .Y(ab_4__1_) );
  NOR2BX2 U106 ( .AN(A[4]), .B(n29), .Y(ab_4__4_) );
  XOR2X2 U107 ( .A(n4), .B(ab_0__4_), .Y(SUMB_1__3_) );
  NOR2BX2 U108 ( .AN(A[8]), .B(n27), .Y(ab_8__6_) );
  NOR2BX2 U109 ( .AN(A[4]), .B(n26), .Y(ab_4__6_) );
  XOR2X4 U110 ( .A(SUMB_16__2_), .B(CARRYB_16__1_), .Y(A1_16_) );
  NOR2BX2 U111 ( .AN(A[3]), .B(n26), .Y(ab_3__6_) );
  BUFX20 U112 ( .A(n44), .Y(n34) );
  INVX8 U113 ( .A(B[1]), .Y(n44) );
  NOR2BX4 U114 ( .AN(A[1]), .B(n29), .Y(ab_1__4_) );
  BUFX20 U115 ( .A(n41), .Y(n29) );
  XOR2X4 U116 ( .A(SUMB_16__1_), .B(CARRYB_16__0_), .Y(A1_15_) );
  NOR2BX2 U117 ( .AN(A[2]), .B(n26), .Y(ab_2__6_) );
  XOR2X4 U118 ( .A(SUMB_15__6_), .B(ab_16__5_), .Y(n15) );
  XOR2X4 U119 ( .A(CARRYB_15__5_), .B(n15), .Y(SUMB_16__5_) );
  NAND2XL U120 ( .A(SUMB_15__6_), .B(CARRYB_15__5_), .Y(n16) );
  NAND2X1 U121 ( .A(ab_16__5_), .B(CARRYB_15__5_), .Y(n17) );
  NAND2XL U122 ( .A(ab_16__5_), .B(SUMB_15__6_), .Y(n18) );
  NOR2BXL U123 ( .AN(A[16]), .B(n28), .Y(ab_16__5_) );
  XOR2X4 U124 ( .A(CARRYB_16__4_), .B(SUMB_16__5_), .Y(A1_19_) );
  AND2X4 U125 ( .A(SUMB_16__1_), .B(CARRYB_16__0_), .Y(n21) );
  NOR2BX2 U126 ( .AN(A[12]), .B(n31), .Y(ab_12__3_) );
  NOR2BX1 U127 ( .AN(A[11]), .B(n36), .Y(ab_11__0_) );
  NOR2BXL U128 ( .AN(A[6]), .B(n28), .Y(ab_6__5_) );
  NOR2BX2 U129 ( .AN(A[14]), .B(n36), .Y(ab_14__0_) );
  NOR2BX2 U130 ( .AN(A[12]), .B(n35), .Y(ab_12__1_) );
  NOR2BX2 U131 ( .AN(A[13]), .B(n36), .Y(ab_13__0_) );
  NOR2BX2 U132 ( .AN(A[12]), .B(n36), .Y(ab_12__0_) );
  NOR2BX1 U133 ( .AN(A[3]), .B(n46), .Y(ab_3__7_) );
  NOR2BX1 U134 ( .AN(A[15]), .B(n27), .Y(ab_15__6_) );
  NOR2BX1 U135 ( .AN(A[15]), .B(n30), .Y(ab_15__4_) );
  INVX4 U136 ( .A(B[2]), .Y(n43) );
  NOR2BX1 U137 ( .AN(A[6]), .B(n32), .Y(ab_6__2_) );
  NOR2BX1 U138 ( .AN(A[9]), .B(n27), .Y(ab_9__6_) );
  NOR2BXL U139 ( .AN(A[7]), .B(n27), .Y(ab_7__6_) );
  NOR2BXL U140 ( .AN(A[6]), .B(n27), .Y(ab_6__6_) );
  NOR2BX1 U141 ( .AN(A[11]), .B(n27), .Y(ab_11__6_) );
  NOR2BX1 U142 ( .AN(A[12]), .B(n27), .Y(ab_12__6_) );
  INVX12 U143 ( .A(B[7]), .Y(n46) );
  XOR2X2 U144 ( .A(CARRYB_16__5_), .B(SUMB_16__6_), .Y(A1_20_) );
  NOR2BX1 U145 ( .AN(A[6]), .B(n29), .Y(ab_6__4_) );
  NOR2BX1 U146 ( .AN(A[6]), .B(n31), .Y(ab_6__3_) );
  NOR2BX1 U147 ( .AN(A[7]), .B(n29), .Y(ab_7__4_) );
  NOR2BXL U148 ( .AN(A[13]), .B(n46), .Y(ab_13__7_) );
  NOR2BX1 U149 ( .AN(A[10]), .B(n33), .Y(ab_10__2_) );
  NOR2BX1 U150 ( .AN(A[10]), .B(n36), .Y(ab_10__0_) );
  NOR2BX1 U151 ( .AN(A[10]), .B(n30), .Y(ab_10__4_) );
  AND2X1 U152 ( .A(CARRYB_16__5_), .B(SUMB_16__6_), .Y(n19) );
  NOR2BX4 U153 ( .AN(A[1]), .B(n40), .Y(ab_1__5_) );
  NOR2BX1 U154 ( .AN(A[2]), .B(n46), .Y(ab_2__7_) );
  NOR2BXL U155 ( .AN(A[14]), .B(n46), .Y(ab_14__7_) );
  NOR2BX1 U156 ( .AN(A[16]), .B(n31), .Y(ab_16__3_) );
  BUFX3 U157 ( .A(n43), .Y(n33) );
  BUFX3 U158 ( .A(n44), .Y(n35) );
  NOR2BX2 U159 ( .AN(A[14]), .B(n35), .Y(ab_14__1_) );
  NOR2BX2 U160 ( .AN(A[13]), .B(n31), .Y(ab_13__3_) );
  NOR2BX2 U161 ( .AN(A[9]), .B(n36), .Y(ab_9__0_) );
  NOR2BX1 U162 ( .AN(A[5]), .B(n42), .Y(ab_5__3_) );
  NOR2BX1 U163 ( .AN(A[5]), .B(n40), .Y(ab_5__5_) );
  NOR2BX2 U164 ( .AN(A[13]), .B(n35), .Y(ab_13__1_) );
  NOR2BX1 U165 ( .AN(A[12]), .B(n46), .Y(ab_12__7_) );
  NOR2BX1 U166 ( .AN(A[13]), .B(n27), .Y(ab_13__6_) );
  NOR2BX1 U167 ( .AN(A[11]), .B(n46), .Y(ab_11__7_) );
  NOR2BX1 U168 ( .AN(A[14]), .B(n27), .Y(ab_14__6_) );
  NOR2BX1 U169 ( .AN(A[10]), .B(n46), .Y(ab_10__7_) );
  AND2X2 U170 ( .A(CARRYB_16__3_), .B(SUMB_16__4_), .Y(n22) );
  NOR2BX1 U171 ( .AN(A[4]), .B(n36), .Y(ab_4__0_) );
  NOR2BX2 U172 ( .AN(A[14]), .B(n31), .Y(ab_14__3_) );
  NOR2BX1 U173 ( .AN(A[8]), .B(n46), .Y(ab_8__7_) );
  NOR2BX1 U174 ( .AN(A[5]), .B(n32), .Y(ab_5__2_) );
  NOR2BX1 U175 ( .AN(A[7]), .B(n46), .Y(ab_7__7_) );
  NOR2BX1 U176 ( .AN(A[6]), .B(n46), .Y(ab_6__7_) );
  NOR2BX1 U177 ( .AN(A[5]), .B(n46), .Y(ab_5__7_) );
  NOR2BX1 U178 ( .AN(A[4]), .B(n46), .Y(ab_4__7_) );
  NOR2BX1 U179 ( .AN(A[9]), .B(n46), .Y(ab_9__7_) );
  NOR2BX2 U180 ( .AN(A[10]), .B(n27), .Y(ab_10__6_) );
  NOR2BX1 U181 ( .AN(A[4]), .B(n40), .Y(ab_4__5_) );
  AND2X2 U182 ( .A(CARRYB_16__4_), .B(SUMB_16__5_), .Y(n23) );
  XOR2X1 U183 ( .A(CARRYB_16__6_), .B(ab_16__7_), .Y(A1_21_) );
  NOR2BX1 U184 ( .AN(A[16]), .B(n27), .Y(ab_16__6_) );
  NOR2BXL U185 ( .AN(A[15]), .B(n46), .Y(ab_15__7_) );
  NOR2BXL U186 ( .AN(A[15]), .B(n36), .Y(ab_15__0_) );
  NOR2BXL U187 ( .AN(A[15]), .B(n33), .Y(ab_15__2_) );
  NOR2BXL U188 ( .AN(A[15]), .B(n28), .Y(ab_15__5_) );
  NOR2BXL U189 ( .AN(A[16]), .B(n36), .Y(ab_16__0_) );
  NOR2BXL U190 ( .AN(A[15]), .B(n35), .Y(ab_15__1_) );
  NOR2BXL U191 ( .AN(A[15]), .B(n31), .Y(ab_15__3_) );
  BUFX1 U192 ( .A(n41), .Y(n30) );
  NOR2BXL U193 ( .AN(A[16]), .B(n46), .Y(ab_16__7_) );
  NOR2BX1 U194 ( .AN(A[0]), .B(n36), .Y(n38) );
  XOR2X4 U195 ( .A(SUMB_16__3_), .B(CARRYB_16__2_), .Y(A1_17_) );
  XOR2X4 U196 ( .A(CARRYB_16__3_), .B(SUMB_16__4_), .Y(A1_18_) );
endmodule


module multi16_10 ( in_17bit, in_8bit, out );
  input [16:0] in_17bit;
  input [7:0] in_8bit;
  output [16:0] out;
  wire   n119, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117;
  wire   [16:2] in_17bit_b;
  wire   [7:1] in_8bit_b;
  wire   [23:8] mul;

  multi16_10_DW02_mult_0 mult_55 ( .A({in_17bit_b, n18, in_17bit[0]}), .B({n17, 
        in_8bit_b[6:1], in_8bit[0]}), .PRODUCT_23_(mul[23]), .PRODUCT_22_(
        mul[22]), .PRODUCT_21_(mul[21]), .PRODUCT_20_(mul[20]), .PRODUCT_19_(
        mul[19]), .PRODUCT_18_(mul[18]), .PRODUCT_17_(mul[17]), .PRODUCT_16_(
        mul[16]), .PRODUCT_15_(mul[15]), .PRODUCT_14_(mul[14]), .PRODUCT_13_(
        mul[13]), .PRODUCT_12_(mul[12]), .PRODUCT_11_(mul[11]), .PRODUCT_10_(
        mul[10]), .PRODUCT_9_(mul[9]), .PRODUCT_8_(mul[8]), .PRODUCT_7_(out[0]) );
  BUFX8 U2 ( .A(mul[20]), .Y(n1) );
  AOI21X4 U3 ( .A0(n58), .A1(n57), .B0(n46), .Y(n59) );
  INVX8 U4 ( .A(n3), .Y(in_17bit_b[2]) );
  BUFX16 U5 ( .A(n26), .Y(n18) );
  BUFX12 U6 ( .A(n119), .Y(out[11]) );
  NOR2X2 U7 ( .A(in_8bit[3]), .B(in_8bit[4]), .Y(n6) );
  CLKINVX4 U8 ( .A(n50), .Y(n9) );
  BUFX16 U9 ( .A(in_8bit[2]), .Y(n50) );
  OR2X2 U10 ( .A(mul[17]), .B(n105), .Y(n2) );
  XOR2X4 U11 ( .A(n16), .B(in_17bit[2]), .Y(n3) );
  NOR2X2 U12 ( .A(n32), .B(n43), .Y(n73) );
  CLKINVX2 U13 ( .A(in_8bit[6]), .Y(n15) );
  NOR2X1 U14 ( .A(n36), .B(n43), .Y(n85) );
  CLKINVX2 U15 ( .A(in_8bit[5]), .Y(n60) );
  INVX2 U16 ( .A(n60), .Y(n8) );
  CLKINVX4 U17 ( .A(in_8bit[0]), .Y(n5) );
  NOR2X4 U18 ( .A(n41), .B(n45), .Y(n11) );
  NOR2X4 U19 ( .A(n39), .B(n43), .Y(n65) );
  OR2X4 U20 ( .A(in_17bit[0]), .B(in_17bit[1]), .Y(n4) );
  NAND3BX4 U21 ( .AN(n48), .B(n5), .C(n6), .Y(n42) );
  NOR2X4 U22 ( .A(n63), .B(n7), .Y(n26) );
  AND3X2 U23 ( .A(in_17bit[16]), .B(in_17bit[0]), .C(in_17bit[1]), .Y(n7) );
  INVX1 U24 ( .A(in_17bit[16]), .Y(n89) );
  NAND2XL U25 ( .A(n90), .B(in_17bit[16]), .Y(n27) );
  NAND2X4 U26 ( .A(n9), .B(n10), .Y(n62) );
  NOR2X4 U27 ( .A(n42), .B(n8), .Y(n10) );
  NAND2X4 U28 ( .A(in_8bit[0]), .B(n44), .Y(n51) );
  XOR2X4 U29 ( .A(n11), .B(n8), .Y(in_8bit_b[5]) );
  INVX4 U30 ( .A(mul[22]), .Y(n113) );
  NOR3XL U31 ( .A(mul[22]), .B(mul[21]), .C(n114), .Y(n115) );
  INVXL U32 ( .A(in_8bit[3]), .Y(n55) );
  XOR2X4 U33 ( .A(n108), .B(mul[21]), .Y(out[14]) );
  NAND2X4 U34 ( .A(n109), .B(n111), .Y(n14) );
  AND2X4 U35 ( .A(n31), .B(n76), .Y(n30) );
  AND2X4 U36 ( .A(n32), .B(n74), .Y(n31) );
  XOR2X2 U37 ( .A(mul[23]), .B(n117), .Y(out[16]) );
  AOI2BB1X4 U38 ( .A0N(n13), .A1N(n1), .B0(n116), .Y(n108) );
  OR2X4 U39 ( .A(n109), .B(mul[19]), .Y(n13) );
  XNOR2X4 U40 ( .A(n14), .B(mul[19]), .Y(out[12]) );
  XOR2X4 U41 ( .A(n61), .B(n15), .Y(in_8bit_b[6]) );
  NAND2X4 U42 ( .A(n106), .B(n111), .Y(n22) );
  NOR2X2 U43 ( .A(n64), .B(in_17bit[2]), .Y(n39) );
  XNOR2X4 U44 ( .A(n65), .B(in_17bit[3]), .Y(n40) );
  NAND2BX4 U45 ( .AN(n47), .B(n62), .Y(n61) );
  CLKINVX8 U46 ( .A(n47), .Y(n44) );
  NOR2XL U47 ( .A(in_8bit[0]), .B(in_8bit[3]), .Y(n57) );
  INVX8 U48 ( .A(n40), .Y(in_17bit_b[3]) );
  CLKINVX8 U49 ( .A(n66), .Y(n68) );
  XNOR2X2 U50 ( .A(mul[18]), .B(n22), .Y(n119) );
  OAI21X4 U51 ( .A0(n50), .A1(n54), .B0(n44), .Y(n56) );
  NAND2X4 U52 ( .A(n95), .B(n111), .Y(n20) );
  OR2X4 U53 ( .A(n48), .B(in_8bit[0]), .Y(n54) );
  XNOR2X2 U54 ( .A(mul[11]), .B(n21), .Y(out[4]) );
  NAND2BX4 U55 ( .AN(in_17bit[3]), .B(n39), .Y(n66) );
  NAND2X4 U56 ( .A(n4), .B(in_17bit[16]), .Y(n16) );
  AND2X2 U57 ( .A(n68), .B(n67), .Y(n34) );
  NOR3X2 U58 ( .A(in_17bit[15]), .B(n90), .C(n43), .Y(in_17bit_b[16]) );
  NAND2X4 U59 ( .A(n35), .B(n88), .Y(n90) );
  XNOR2X4 U60 ( .A(mul[12]), .B(n20), .Y(out[5]) );
  BUFX4 U61 ( .A(in_8bit_b[7]), .Y(n17) );
  NOR3X1 U62 ( .A(in_8bit[6]), .B(n62), .C(n46), .Y(in_8bit_b[7]) );
  OAI21X4 U63 ( .A0(n114), .A1(mul[21]), .B0(n111), .Y(n112) );
  NOR2X4 U64 ( .A(n50), .B(n48), .Y(n58) );
  XNOR2X4 U65 ( .A(mul[10]), .B(n24), .Y(out[3]) );
  NAND2X4 U66 ( .A(n93), .B(n111), .Y(n24) );
  NAND2BX4 U67 ( .AN(mul[13]), .B(n97), .Y(n99) );
  CLKINVX3 U68 ( .A(n96), .Y(n97) );
  NAND2X4 U69 ( .A(n100), .B(n111), .Y(n25) );
  XOR2X4 U70 ( .A(n49), .B(n51), .Y(in_8bit_b[1]) );
  INVX12 U71 ( .A(in_8bit[7]), .Y(n47) );
  AND2X4 U72 ( .A(n34), .B(n70), .Y(n33) );
  NOR2X2 U73 ( .A(n34), .B(n43), .Y(n69) );
  NAND2X4 U74 ( .A(n96), .B(n111), .Y(n23) );
  OR2X4 U75 ( .A(mul[12]), .B(n95), .Y(n96) );
  XOR2X4 U76 ( .A(n50), .B(n53), .Y(in_8bit_b[2]) );
  NOR2X4 U77 ( .A(n52), .B(n45), .Y(n53) );
  CLKINVX8 U78 ( .A(n49), .Y(n48) );
  NAND2BX4 U79 ( .AN(mul[20]), .B(n110), .Y(n114) );
  NOR2X2 U80 ( .A(n109), .B(mul[19]), .Y(n110) );
  INVX8 U81 ( .A(in_8bit[1]), .Y(n49) );
  AND2X1 U82 ( .A(n33), .B(n72), .Y(n32) );
  AND2X2 U83 ( .A(n30), .B(n78), .Y(n29) );
  AND2X4 U84 ( .A(n37), .B(n84), .Y(n36) );
  OR2X4 U85 ( .A(mul[18]), .B(n2), .Y(n109) );
  OR2X4 U86 ( .A(mul[9]), .B(n92), .Y(n93) );
  OR2X4 U87 ( .A(mul[11]), .B(n94), .Y(n95) );
  OR2X4 U88 ( .A(mul[14]), .B(n99), .Y(n100) );
  OR2X4 U89 ( .A(mul[16]), .B(n103), .Y(n105) );
  XOR2X4 U90 ( .A(mul[8]), .B(n19), .Y(out[1]) );
  AND2X4 U91 ( .A(out[0]), .B(n111), .Y(n19) );
  XNOR2X4 U92 ( .A(mul[9]), .B(n91), .Y(out[2]) );
  NAND2X4 U93 ( .A(n92), .B(n111), .Y(n91) );
  NAND2X1 U94 ( .A(n94), .B(n111), .Y(n21) );
  XNOR2X4 U95 ( .A(mul[13]), .B(n23), .Y(out[6]) );
  XNOR2X4 U96 ( .A(mul[15]), .B(n25), .Y(out[8]) );
  OR2X4 U97 ( .A(n68), .B(n43), .Y(n28) );
  AND2X4 U98 ( .A(n36), .B(n86), .Y(n35) );
  INVX4 U99 ( .A(n116), .Y(n111) );
  BUFX12 U100 ( .A(n89), .Y(n43) );
  XNOR2X2 U101 ( .A(n27), .B(in_17bit[15]), .Y(in_17bit_b[15]) );
  OR2X2 U102 ( .A(mul[10]), .B(n93), .Y(n94) );
  OR2X2 U103 ( .A(mul[8]), .B(out[0]), .Y(n92) );
  INVX1 U104 ( .A(n54), .Y(n52) );
  OR2X4 U105 ( .A(mul[17]), .B(n105), .Y(n106) );
  INVXL U106 ( .A(in_8bit[7]), .Y(n45) );
  INVXL U107 ( .A(in_8bit[7]), .Y(n46) );
  XOR2X4 U108 ( .A(n28), .B(n67), .Y(in_17bit_b[4]) );
  AND2X2 U109 ( .A(n38), .B(n82), .Y(n37) );
  AND2X2 U110 ( .A(n29), .B(n80), .Y(n38) );
  NOR2X1 U111 ( .A(n116), .B(n115), .Y(n117) );
  XNOR2X1 U112 ( .A(in_17bit[16]), .B(n44), .Y(n116) );
  NOR2X4 U113 ( .A(n50), .B(n42), .Y(n41) );
  XNOR2X4 U114 ( .A(n1), .B(n107), .Y(out[13]) );
  OAI21X4 U115 ( .A0(mul[19]), .A1(n109), .B0(n111), .Y(n107) );
  XOR2X4 U116 ( .A(n56), .B(n55), .Y(in_8bit_b[3]) );
  XOR2X4 U117 ( .A(n59), .B(in_8bit[4]), .Y(in_8bit_b[4]) );
  OR2X4 U118 ( .A(in_17bit[0]), .B(in_17bit[1]), .Y(n64) );
  OAI21X4 U119 ( .A0(in_17bit[16]), .A1(in_17bit[1]), .B0(n64), .Y(n63) );
  CLKINVX3 U120 ( .A(in_17bit[4]), .Y(n67) );
  CLKINVX3 U121 ( .A(in_17bit[5]), .Y(n70) );
  XNOR2X4 U122 ( .A(n69), .B(n70), .Y(in_17bit_b[5]) );
  NOR2X4 U123 ( .A(n33), .B(n43), .Y(n71) );
  CLKINVX3 U124 ( .A(in_17bit[6]), .Y(n72) );
  XNOR2X4 U125 ( .A(n71), .B(n72), .Y(in_17bit_b[6]) );
  CLKINVX3 U126 ( .A(in_17bit[7]), .Y(n74) );
  XNOR2X4 U127 ( .A(n73), .B(n74), .Y(in_17bit_b[7]) );
  NOR2X4 U128 ( .A(n31), .B(n43), .Y(n75) );
  CLKINVX3 U129 ( .A(in_17bit[8]), .Y(n76) );
  XNOR2X4 U130 ( .A(n75), .B(n76), .Y(in_17bit_b[8]) );
  NOR2X4 U131 ( .A(n30), .B(n43), .Y(n77) );
  CLKINVX3 U132 ( .A(in_17bit[9]), .Y(n78) );
  XNOR2X4 U133 ( .A(n77), .B(n78), .Y(in_17bit_b[9]) );
  NOR2X4 U134 ( .A(n29), .B(n43), .Y(n79) );
  CLKINVX3 U135 ( .A(in_17bit[10]), .Y(n80) );
  XNOR2X4 U136 ( .A(n79), .B(n80), .Y(in_17bit_b[10]) );
  NOR2X4 U137 ( .A(n38), .B(n43), .Y(n81) );
  CLKINVX3 U138 ( .A(in_17bit[11]), .Y(n82) );
  XNOR2X4 U139 ( .A(n81), .B(n82), .Y(in_17bit_b[11]) );
  NOR2X4 U140 ( .A(n37), .B(n43), .Y(n83) );
  CLKINVX3 U141 ( .A(in_17bit[12]), .Y(n84) );
  XNOR2X4 U142 ( .A(n83), .B(n84), .Y(in_17bit_b[12]) );
  CLKINVX3 U143 ( .A(in_17bit[13]), .Y(n86) );
  XNOR2X4 U144 ( .A(n85), .B(n86), .Y(in_17bit_b[13]) );
  NOR2X4 U145 ( .A(n35), .B(n43), .Y(n87) );
  CLKINVX3 U146 ( .A(in_17bit[14]), .Y(n88) );
  XNOR2X4 U147 ( .A(n87), .B(n88), .Y(in_17bit_b[14]) );
  NAND2X4 U148 ( .A(n99), .B(n111), .Y(n98) );
  XNOR2X4 U149 ( .A(mul[14]), .B(n98), .Y(out[7]) );
  CLKINVX3 U150 ( .A(n100), .Y(n101) );
  NAND2BX4 U151 ( .AN(mul[15]), .B(n101), .Y(n103) );
  NAND2X4 U152 ( .A(n103), .B(n111), .Y(n102) );
  XNOR2X4 U153 ( .A(mul[16]), .B(n102), .Y(out[9]) );
  NAND2X4 U154 ( .A(n105), .B(n111), .Y(n104) );
  XNOR2X4 U155 ( .A(n104), .B(mul[17]), .Y(out[10]) );
  XOR2X4 U156 ( .A(n113), .B(n112), .Y(out[15]) );
endmodule


module multi16_9_DW01_add_4 ( A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, 
        A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, 
        B_20_, B_19_, B_18_, B_17_, B_16_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, 
        SUM_17_, SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, 
        SUM_9_, SUM_8_, SUM_7_, SUM_6_, SUM_5_ );
  input A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_,
         A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, B_20_, B_19_,
         B_18_, B_17_, B_16_;
  output SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, SUM_15_,
         SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, SUM_7_,
         SUM_6_, SUM_5_;
  wire   n42, n1, n2, n3, n5, n6, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41;

  OAI2BB1X4 U2 ( .A0N(n35), .A1N(n1), .B0(n29), .Y(n33) );
  CLKINVX20 U3 ( .A(n6), .Y(n1) );
  NOR2X2 U4 ( .A(n5), .B(n6), .Y(n28) );
  AND2X4 U5 ( .A(A_16_), .B(B_16_), .Y(n2) );
  BUFX16 U6 ( .A(n42), .Y(SUM_17_) );
  NAND2X4 U7 ( .A(n38), .B(n2), .Y(n37) );
  OR2X2 U8 ( .A(A_17_), .B(B_17_), .Y(n38) );
  NOR2X2 U9 ( .A(A_17_), .B(B_17_), .Y(n3) );
  NAND2X1 U10 ( .A(n19), .B(n20), .Y(n18) );
  XNOR2X4 U11 ( .A(n40), .B(n31), .Y(n42) );
  BUFX8 U12 ( .A(A_6_), .Y(SUM_6_) );
  BUFX12 U13 ( .A(A_11_), .Y(SUM_11_) );
  OAI21X2 U14 ( .A0(n26), .A1(n27), .B0(n28), .Y(n25) );
  BUFX12 U15 ( .A(A_14_), .Y(SUM_14_) );
  BUFX12 U16 ( .A(A_15_), .Y(SUM_15_) );
  NAND2X4 U17 ( .A(n30), .B(n37), .Y(n35) );
  NAND2X4 U18 ( .A(A_17_), .B(B_17_), .Y(n30) );
  INVX8 U19 ( .A(n41), .Y(SUM_16_) );
  NAND2X4 U20 ( .A(n31), .B(n39), .Y(n41) );
  NAND2X4 U21 ( .A(B_16_), .B(A_16_), .Y(n31) );
  NOR2BX4 U22 ( .AN(n32), .B(n5), .Y(n34) );
  BUFX12 U23 ( .A(A_12_), .Y(SUM_12_) );
  NOR2X4 U24 ( .A(A_19_), .B(B_19_), .Y(n5) );
  NAND2X2 U25 ( .A(B_19_), .B(A_19_), .Y(n32) );
  NOR2BX4 U26 ( .AN(n30), .B(n3), .Y(n40) );
  NAND2X4 U27 ( .A(n32), .B(n25), .Y(n21) );
  OR2X4 U28 ( .A(A_16_), .B(B_16_), .Y(n39) );
  BUFX8 U29 ( .A(A_5_), .Y(SUM_5_) );
  NAND2X2 U30 ( .A(B_20_), .B(A_20_), .Y(n19) );
  NOR2XL U31 ( .A(n31), .B(n3), .Y(n26) );
  NAND2XL U32 ( .A(n29), .B(n30), .Y(n27) );
  NAND2XL U33 ( .A(n21), .B(n22), .Y(n20) );
  NOR2X4 U34 ( .A(A_18_), .B(B_18_), .Y(n6) );
  BUFX8 U35 ( .A(A_9_), .Y(SUM_9_) );
  BUFX8 U36 ( .A(A_10_), .Y(SUM_10_) );
  BUFX8 U37 ( .A(A_7_), .Y(SUM_7_) );
  BUFX8 U38 ( .A(A_8_), .Y(SUM_8_) );
  BUFX8 U39 ( .A(A_13_), .Y(SUM_13_) );
  XOR3X4 U40 ( .A(B_21_), .B(A_21_), .C(n18), .Y(SUM_21_) );
  XOR2X4 U41 ( .A(n21), .B(n23), .Y(SUM_20_) );
  NOR2BX4 U42 ( .AN(n19), .B(n24), .Y(n23) );
  CLKINVX3 U43 ( .A(n22), .Y(n24) );
  OR2X4 U44 ( .A(A_20_), .B(B_20_), .Y(n22) );
  XOR2X4 U45 ( .A(n33), .B(n34), .Y(SUM_19_) );
  XOR2X4 U46 ( .A(n35), .B(n36), .Y(SUM_18_) );
  NOR2BX4 U47 ( .AN(n29), .B(n6), .Y(n36) );
  NAND2X4 U48 ( .A(B_18_), .B(A_18_), .Y(n29) );
endmodule


module multi16_9_DW02_mult_0 ( A, B, PRODUCT_23_, PRODUCT_22_, PRODUCT_21_, 
        PRODUCT_20_, PRODUCT_19_, PRODUCT_18_, PRODUCT_17_, PRODUCT_16_, 
        PRODUCT_15_, PRODUCT_14_, PRODUCT_13_, PRODUCT_12_, PRODUCT_11_, 
        PRODUCT_10_, PRODUCT_9_, PRODUCT_8_, PRODUCT_7_ );
  input [16:0] A;
  input [7:0] B;
  output PRODUCT_23_, PRODUCT_22_, PRODUCT_21_, PRODUCT_20_, PRODUCT_19_,
         PRODUCT_18_, PRODUCT_17_, PRODUCT_16_, PRODUCT_15_, PRODUCT_14_,
         PRODUCT_13_, PRODUCT_12_, PRODUCT_11_, PRODUCT_10_, PRODUCT_9_,
         PRODUCT_8_, PRODUCT_7_;
  wire   ab_16__7_, ab_16__6_, ab_16__5_, ab_16__4_, ab_16__3_, ab_16__2_,
         ab_16__1_, ab_16__0_, ab_15__7_, ab_15__6_, ab_15__5_, ab_15__4_,
         ab_15__3_, ab_15__2_, ab_15__1_, ab_15__0_, ab_14__7_, ab_14__6_,
         ab_14__5_, ab_14__4_, ab_14__3_, ab_14__2_, ab_14__1_, ab_14__0_,
         ab_13__7_, ab_13__6_, ab_13__5_, ab_13__4_, ab_13__3_, ab_13__2_,
         ab_13__1_, ab_13__0_, ab_12__7_, ab_12__6_, ab_12__5_, ab_12__4_,
         ab_12__3_, ab_12__2_, ab_12__1_, ab_12__0_, ab_11__7_, ab_11__6_,
         ab_11__5_, ab_11__4_, ab_11__3_, ab_11__2_, ab_11__1_, ab_11__0_,
         ab_10__7_, ab_10__6_, ab_10__5_, ab_10__4_, ab_10__3_, ab_10__2_,
         ab_10__1_, ab_10__0_, ab_9__7_, ab_9__6_, ab_9__5_, ab_9__4_,
         ab_9__3_, ab_9__2_, ab_9__1_, ab_9__0_, ab_8__7_, ab_8__6_, ab_8__5_,
         ab_8__4_, ab_8__3_, ab_8__2_, ab_8__1_, ab_8__0_, ab_7__7_, ab_7__6_,
         ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_, ab_7__0_, ab_6__7_,
         ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_, ab_6__1_, ab_6__0_,
         ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_, ab_5__2_, ab_5__1_,
         ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_, ab_4__3_, ab_4__2_,
         ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_, ab_3__4_, ab_3__3_,
         ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_, ab_2__5_, ab_2__4_,
         ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_, ab_1__6_, ab_1__5_,
         ab_1__4_, ab_1__3_, ab_1__2_, ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_,
         ab_0__3_, ab_0__2_, CARRYB_16__6_, CARRYB_16__5_, CARRYB_16__4_,
         CARRYB_16__3_, CARRYB_16__2_, CARRYB_16__1_, CARRYB_16__0_,
         CARRYB_15__6_, CARRYB_15__5_, CARRYB_15__4_, CARRYB_15__3_,
         CARRYB_15__2_, CARRYB_15__1_, CARRYB_15__0_, CARRYB_14__6_,
         CARRYB_14__5_, CARRYB_14__4_, CARRYB_14__3_, CARRYB_14__2_,
         CARRYB_14__1_, CARRYB_14__0_, CARRYB_13__6_, CARRYB_13__5_,
         CARRYB_13__4_, CARRYB_13__3_, CARRYB_13__2_, CARRYB_13__1_,
         CARRYB_13__0_, CARRYB_12__6_, CARRYB_12__5_, CARRYB_12__4_,
         CARRYB_12__3_, CARRYB_12__2_, CARRYB_12__1_, CARRYB_12__0_,
         CARRYB_11__6_, CARRYB_11__5_, CARRYB_11__4_, CARRYB_11__3_,
         CARRYB_11__2_, CARRYB_11__1_, CARRYB_11__0_, CARRYB_10__6_,
         CARRYB_10__5_, CARRYB_10__4_, CARRYB_10__3_, CARRYB_10__2_,
         CARRYB_10__1_, CARRYB_10__0_, CARRYB_9__6_, CARRYB_9__5_,
         CARRYB_9__4_, CARRYB_9__3_, CARRYB_9__2_, CARRYB_9__1_, CARRYB_9__0_,
         CARRYB_8__6_, CARRYB_8__5_, CARRYB_8__4_, CARRYB_8__3_, CARRYB_8__2_,
         CARRYB_8__1_, CARRYB_8__0_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_,
         CARRYB_7__3_, CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_,
         CARRYB_6__5_, CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_,
         CARRYB_6__0_, CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_,
         CARRYB_5__2_, CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_,
         CARRYB_4__4_, CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_,
         CARRYB_3__6_, CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_,
         CARRYB_3__1_, CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_,
         CARRYB_2__3_, CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__0_,
         SUMB_16__6_, SUMB_16__5_, SUMB_16__4_, SUMB_16__3_, SUMB_16__2_,
         SUMB_16__1_, SUMB_16__0_, SUMB_15__6_, SUMB_15__5_, SUMB_15__4_,
         SUMB_15__3_, SUMB_15__2_, SUMB_15__1_, SUMB_14__6_, SUMB_14__5_,
         SUMB_14__4_, SUMB_14__3_, SUMB_14__2_, SUMB_14__1_, SUMB_13__6_,
         SUMB_13__5_, SUMB_13__4_, SUMB_13__3_, SUMB_13__2_, SUMB_13__1_,
         SUMB_12__6_, SUMB_12__5_, SUMB_12__4_, SUMB_12__3_, SUMB_12__2_,
         SUMB_12__1_, SUMB_11__6_, SUMB_11__5_, SUMB_11__4_, SUMB_11__3_,
         SUMB_11__2_, SUMB_11__1_, SUMB_10__6_, SUMB_10__5_, SUMB_10__4_,
         SUMB_10__3_, SUMB_10__2_, SUMB_10__1_, SUMB_9__6_, SUMB_9__5_,
         SUMB_9__4_, SUMB_9__3_, SUMB_9__2_, SUMB_9__1_, SUMB_8__6_,
         SUMB_8__5_, SUMB_8__4_, SUMB_8__3_, SUMB_8__2_, SUMB_8__1_,
         SUMB_7__6_, SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_,
         SUMB_7__1_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, PROD1_7_, A1_21_, A1_20_, A1_19_, A1_18_,
         A1_17_, A1_16_, A1_15_, A1_13_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_,
         A1_7_, A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, n3, n4, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41;

  ADDFHX2 S5_6 ( .A(ab_16__6_), .B(CARRYB_15__6_), .CI(ab_15__7_), .CO(
        CARRYB_16__6_), .S(SUMB_16__6_) );
  ADDFHX2 S2_15_5 ( .A(ab_15__5_), .B(CARRYB_14__5_), .CI(SUMB_14__6_), .CO(
        CARRYB_15__5_), .S(SUMB_15__5_) );
  ADDFHX2 S3_15_6 ( .A(ab_15__6_), .B(CARRYB_14__6_), .CI(ab_14__7_), .CO(
        CARRYB_15__6_), .S(SUMB_15__6_) );
  multi16_9_DW01_add_4 FS_1 ( .A_21_(A1_21_), .A_20_(A1_20_), .A_19_(A1_19_), 
        .A_18_(A1_18_), .A_17_(A1_17_), .A_16_(A1_16_), .A_15_(A1_15_), 
        .A_14_(SUMB_16__0_), .A_13_(A1_13_), .A_12_(A1_12_), .A_11_(A1_11_), 
        .A_10_(A1_10_), .A_9_(A1_9_), .A_8_(A1_8_), .A_7_(A1_7_), .A_6_(A1_6_), 
        .A_5_(PROD1_7_), .B_21_(n4), .B_20_(n19), .B_19_(n18), .B_18_(n17), 
        .B_17_(n8), .B_16_(n16), .SUM_21_(PRODUCT_23_), .SUM_20_(PRODUCT_22_), 
        .SUM_19_(PRODUCT_21_), .SUM_18_(PRODUCT_20_), .SUM_17_(PRODUCT_19_), 
        .SUM_16_(PRODUCT_18_), .SUM_15_(PRODUCT_17_), .SUM_14_(PRODUCT_16_), 
        .SUM_13_(PRODUCT_15_), .SUM_12_(PRODUCT_14_), .SUM_11_(PRODUCT_13_), 
        .SUM_10_(PRODUCT_12_), .SUM_9_(PRODUCT_11_), .SUM_8_(PRODUCT_10_), 
        .SUM_7_(PRODUCT_9_), .SUM_6_(PRODUCT_8_), .SUM_5_(PRODUCT_7_) );
  ADDFHX4 S2_12_1 ( .A(ab_12__1_), .B(CARRYB_11__1_), .CI(SUMB_11__2_), .CO(
        CARRYB_12__1_), .S(SUMB_12__1_) );
  ADDFHX4 S1_12_0 ( .A(ab_12__0_), .B(CARRYB_11__0_), .CI(SUMB_11__1_), .CO(
        CARRYB_12__0_), .S(A1_10_) );
  ADDFHX4 S2_10_5 ( .A(ab_10__5_), .B(CARRYB_9__5_), .CI(SUMB_9__6_), .CO(
        CARRYB_10__5_), .S(SUMB_10__5_) );
  ADDFHX4 S2_11_5 ( .A(ab_11__5_), .B(CARRYB_10__5_), .CI(SUMB_10__6_), .CO(
        CARRYB_11__5_), .S(SUMB_11__5_) );
  ADDFHX4 S4_1 ( .A(ab_16__1_), .B(CARRYB_15__1_), .CI(SUMB_15__2_), .CO(
        CARRYB_16__1_), .S(SUMB_16__1_) );
  ADDFHX4 S1_9_0 ( .A(ab_9__0_), .B(CARRYB_8__0_), .CI(SUMB_8__1_), .CO(
        CARRYB_9__0_), .S(A1_7_) );
  ADDFHX4 S1_10_0 ( .A(ab_10__0_), .B(CARRYB_9__0_), .CI(SUMB_9__1_), .CO(
        CARRYB_10__0_), .S(A1_8_) );
  ADDFHX4 S2_13_2 ( .A(ab_13__2_), .B(CARRYB_12__2_), .CI(SUMB_12__3_), .CO(
        CARRYB_13__2_), .S(SUMB_13__2_) );
  ADDFHX4 S2_14_2 ( .A(ab_14__2_), .B(CARRYB_13__2_), .CI(SUMB_13__3_), .CO(
        CARRYB_14__2_), .S(SUMB_14__2_) );
  ADDFHX4 S2_12_4 ( .A(ab_12__4_), .B(CARRYB_11__4_), .CI(SUMB_11__5_), .CO(
        CARRYB_12__4_), .S(SUMB_12__4_) );
  ADDFHX4 S2_13_4 ( .A(ab_13__4_), .B(CARRYB_12__4_), .CI(SUMB_12__5_), .CO(
        CARRYB_13__4_), .S(SUMB_13__4_) );
  ADDFHX4 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  ADDFHX4 S1_7_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(PROD1_7_) );
  ADDFHX4 S2_10_3 ( .A(ab_10__3_), .B(CARRYB_9__3_), .CI(SUMB_9__4_), .CO(
        CARRYB_10__3_), .S(SUMB_10__3_) );
  ADDFHX4 S2_13_3 ( .A(ab_13__3_), .B(CARRYB_12__3_), .CI(SUMB_12__4_), .CO(
        CARRYB_13__3_), .S(SUMB_13__3_) );
  ADDFHX4 S2_14_3 ( .A(ab_14__3_), .B(CARRYB_13__3_), .CI(SUMB_13__4_), .CO(
        CARRYB_14__3_), .S(SUMB_14__3_) );
  ADDFHX4 S2_12_5 ( .A(ab_12__5_), .B(CARRYB_11__5_), .CI(SUMB_11__6_), .CO(
        CARRYB_12__5_), .S(SUMB_12__5_) );
  ADDFHX4 S2_11_2 ( .A(ab_11__2_), .B(CARRYB_10__2_), .CI(SUMB_10__3_), .CO(
        CARRYB_11__2_), .S(SUMB_11__2_) );
  ADDFHX4 S2_8_2 ( .A(ab_8__2_), .B(CARRYB_7__2_), .CI(SUMB_7__3_), .CO(
        CARRYB_8__2_), .S(SUMB_8__2_) );
  ADDFHX4 S1_15_0 ( .A(ab_15__0_), .B(CARRYB_14__0_), .CI(SUMB_14__1_), .CO(
        CARRYB_15__0_), .S(A1_13_) );
  ADDFHX4 S4_0 ( .A(ab_16__0_), .B(CARRYB_15__0_), .CI(SUMB_15__1_), .CO(
        CARRYB_16__0_), .S(SUMB_16__0_) );
  ADDFHX4 S2_8_1 ( .A(ab_8__1_), .B(CARRYB_7__1_), .CI(SUMB_7__2_), .CO(
        CARRYB_8__1_), .S(SUMB_8__1_) );
  ADDFHX4 S2_11_1 ( .A(ab_11__1_), .B(CARRYB_10__1_), .CI(SUMB_10__2_), .CO(
        CARRYB_11__1_), .S(SUMB_11__1_) );
  ADDFHX4 S2_13_1 ( .A(ab_13__1_), .B(CARRYB_12__1_), .CI(SUMB_12__2_), .CO(
        CARRYB_13__1_), .S(SUMB_13__1_) );
  ADDFHX4 S2_11_4 ( .A(ab_11__4_), .B(CARRYB_10__4_), .CI(SUMB_10__5_), .CO(
        CARRYB_11__4_), .S(SUMB_11__4_) );
  ADDFHX4 S2_11_3 ( .A(ab_11__3_), .B(CARRYB_10__3_), .CI(SUMB_10__4_), .CO(
        CARRYB_11__3_), .S(SUMB_11__3_) );
  ADDFHX4 S1_13_0 ( .A(ab_13__0_), .B(CARRYB_12__0_), .CI(SUMB_12__1_), .CO(
        CARRYB_13__0_), .S(A1_11_) );
  ADDFHX4 S1_14_0 ( .A(ab_14__0_), .B(CARRYB_13__0_), .CI(SUMB_13__1_), .CO(
        CARRYB_14__0_), .S(A1_12_) );
  ADDFHX4 S4_2 ( .A(ab_16__2_), .B(CARRYB_15__2_), .CI(SUMB_15__3_), .CO(
        CARRYB_16__2_), .S(SUMB_16__2_) );
  ADDFHX4 S4_3 ( .A(ab_16__3_), .B(CARRYB_15__3_), .CI(SUMB_15__4_), .CO(
        CARRYB_16__3_), .S(SUMB_16__3_) );
  ADDFHX4 S3_7_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(
        CARRYB_7__6_), .S(SUMB_7__6_) );
  ADDFHX4 S3_8_6 ( .A(ab_8__6_), .B(CARRYB_7__6_), .CI(ab_7__7_), .CO(
        CARRYB_8__6_), .S(SUMB_8__6_) );
  ADDFHX4 S2_9_4 ( .A(ab_9__4_), .B(CARRYB_8__4_), .CI(SUMB_8__5_), .CO(
        CARRYB_9__4_), .S(SUMB_9__4_) );
  ADDFHX4 S2_10_4 ( .A(ab_10__4_), .B(CARRYB_9__4_), .CI(SUMB_9__5_), .CO(
        CARRYB_10__4_), .S(SUMB_10__4_) );
  ADDFHX4 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  ADDFHX4 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  ADDFHX4 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  ADDFHX4 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  ADDFHX4 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  ADDFHX4 S3_11_6 ( .A(ab_11__6_), .B(CARRYB_10__6_), .CI(ab_10__7_), .CO(
        CARRYB_11__6_), .S(SUMB_11__6_) );
  ADDFHX4 S3_12_6 ( .A(ab_12__6_), .B(CARRYB_11__6_), .CI(ab_11__7_), .CO(
        CARRYB_12__6_), .S(SUMB_12__6_) );
  ADDFHX4 S2_9_5 ( .A(ab_9__5_), .B(CARRYB_8__5_), .CI(SUMB_8__6_), .CO(
        CARRYB_9__5_), .S(SUMB_9__5_) );
  ADDFHX4 S2_15_1 ( .A(ab_15__1_), .B(CARRYB_14__1_), .CI(SUMB_14__2_), .CO(
        CARRYB_15__1_), .S(SUMB_15__1_) );
  ADDFHX4 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  ADDFHX4 S2_7_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  ADDFHX4 S2_9_1 ( .A(ab_9__1_), .B(CARRYB_8__1_), .CI(SUMB_8__2_), .CO(
        CARRYB_9__1_), .S(SUMB_9__1_) );
  ADDFHX4 S2_14_1 ( .A(ab_14__1_), .B(CARRYB_13__1_), .CI(SUMB_13__2_), .CO(
        CARRYB_14__1_), .S(SUMB_14__1_) );
  ADDFHX4 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  ADDFHX4 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  ADDFHX4 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  ADDFHX4 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  ADDFHX4 S2_12_3 ( .A(ab_12__3_), .B(CARRYB_11__3_), .CI(SUMB_11__4_), .CO(
        CARRYB_12__3_), .S(SUMB_12__3_) );
  ADDFHX4 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  ADDFHX4 S2_10_2 ( .A(ab_10__2_), .B(CARRYB_9__2_), .CI(SUMB_9__3_), .CO(
        CARRYB_10__2_), .S(SUMB_10__2_) );
  ADDFHX4 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  ADDFHX4 S2_2_1 ( .A(ab_2__1_), .B(n10), .CI(SUMB_1__2_), .CO(CARRYB_2__1_), 
        .S(SUMB_2__1_) );
  ADDFHX4 S1_11_0 ( .A(ab_11__0_), .B(CARRYB_10__0_), .CI(SUMB_10__1_), .CO(
        CARRYB_11__0_), .S(A1_9_) );
  ADDFHX4 S2_8_5 ( .A(ab_8__5_), .B(CARRYB_7__5_), .CI(SUMB_7__6_), .CO(
        CARRYB_8__5_), .S(SUMB_8__5_) );
  ADDFHX4 S3_9_6 ( .A(ab_9__6_), .B(CARRYB_8__6_), .CI(ab_8__7_), .CO(
        CARRYB_9__6_), .S(SUMB_9__6_) );
  ADDFHX4 S3_10_6 ( .A(ab_10__6_), .B(CARRYB_9__6_), .CI(ab_9__7_), .CO(
        CARRYB_10__6_), .S(SUMB_10__6_) );
  ADDFHX4 S4_5 ( .A(ab_16__5_), .B(CARRYB_15__5_), .CI(SUMB_15__6_), .CO(
        CARRYB_16__5_), .S(SUMB_16__5_) );
  ADDFHX4 S2_7_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  ADDFHX4 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  ADDFHX4 S2_9_3 ( .A(ab_9__3_), .B(CARRYB_8__3_), .CI(SUMB_8__4_), .CO(
        CARRYB_9__3_), .S(SUMB_9__3_) );
  ADDFHX4 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  ADDFHX4 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  ADDFHX4 S2_7_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  ADDFHX4 S2_2_4 ( .A(ab_2__4_), .B(n12), .CI(SUMB_1__5_), .CO(CARRYB_2__4_), 
        .S(SUMB_2__4_) );
  ADDFHX4 S2_14_4 ( .A(ab_14__4_), .B(CARRYB_13__4_), .CI(SUMB_13__5_), .CO(
        CARRYB_14__4_), .S(SUMB_14__4_) );
  ADDFHX4 S2_15_3 ( .A(ab_15__3_), .B(CARRYB_14__3_), .CI(SUMB_14__4_), .CO(
        CARRYB_15__3_), .S(SUMB_15__3_) );
  ADDFHX4 S2_7_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  ADDFHX4 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  ADDFHX4 S2_2_5 ( .A(ab_2__5_), .B(n7), .CI(SUMB_1__6_), .CO(CARRYB_2__5_), 
        .S(SUMB_2__5_) );
  ADDFHX4 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  ADDFHX4 S3_2_6 ( .A(ab_2__6_), .B(n6), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  ADDFHX4 S3_3_6 ( .A(ab_3__6_), .B(ab_2__7_), .CI(CARRYB_2__6_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  ADDFHX4 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  ADDFHX4 S2_2_3 ( .A(ab_2__3_), .B(n13), .CI(SUMB_1__4_), .CO(CARRYB_2__3_), 
        .S(SUMB_2__3_) );
  ADDFHX4 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  ADDFHX4 S2_7_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  ADDFHX4 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  ADDFHX4 S2_2_2 ( .A(ab_2__2_), .B(n9), .CI(SUMB_1__3_), .CO(CARRYB_2__2_), 
        .S(SUMB_2__2_) );
  ADDFHX4 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  ADDFHX4 S1_8_0 ( .A(ab_8__0_), .B(CARRYB_7__0_), .CI(SUMB_7__1_), .CO(
        CARRYB_8__0_), .S(A1_6_) );
  ADDFHX4 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  ADDFHX4 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  ADDFHX4 S4_4 ( .A(ab_16__4_), .B(CARRYB_15__4_), .CI(SUMB_15__5_), .CO(
        CARRYB_16__4_), .S(SUMB_16__4_) );
  ADDFHX4 S2_8_3 ( .A(ab_8__3_), .B(CARRYB_7__3_), .CI(SUMB_7__4_), .CO(
        CARRYB_8__3_), .S(SUMB_8__3_) );
  ADDFHX4 S2_12_2 ( .A(ab_12__2_), .B(CARRYB_11__2_), .CI(SUMB_11__3_), .CO(
        CARRYB_12__2_), .S(SUMB_12__2_) );
  ADDFHX4 S3_13_6 ( .A(ab_13__6_), .B(CARRYB_12__6_), .CI(ab_12__7_), .CO(
        CARRYB_13__6_), .S(SUMB_13__6_) );
  ADDFHX4 S3_14_6 ( .A(ab_14__6_), .B(CARRYB_13__6_), .CI(ab_13__7_), .CO(
        CARRYB_14__6_), .S(SUMB_14__6_) );
  ADDFHX4 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  ADDFHX4 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  ADDFHX4 S2_10_1 ( .A(ab_10__1_), .B(CARRYB_9__1_), .CI(SUMB_9__2_), .CO(
        CARRYB_10__1_), .S(SUMB_10__1_) );
  ADDFHX4 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  ADDFHX4 S2_8_4 ( .A(ab_8__4_), .B(CARRYB_7__4_), .CI(SUMB_7__5_), .CO(
        CARRYB_8__4_), .S(SUMB_8__4_) );
  ADDFHX4 S2_9_2 ( .A(ab_9__2_), .B(CARRYB_8__2_), .CI(SUMB_8__3_), .CO(
        CARRYB_9__2_), .S(SUMB_9__2_) );
  ADDFHX4 S2_13_5 ( .A(ab_13__5_), .B(CARRYB_12__5_), .CI(SUMB_12__6_), .CO(
        CARRYB_13__5_), .S(SUMB_13__5_) );
  ADDFHX4 S2_14_5 ( .A(ab_14__5_), .B(CARRYB_13__5_), .CI(SUMB_13__6_), .CO(
        CARRYB_14__5_), .S(SUMB_14__5_) );
  ADDFHX4 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  ADDFHX4 S2_15_2 ( .A(ab_15__2_), .B(CARRYB_14__2_), .CI(SUMB_14__3_), .CO(
        CARRYB_15__2_), .S(SUMB_15__2_) );
  ADDFHX4 S2_15_4 ( .A(ab_15__4_), .B(CARRYB_14__4_), .CI(SUMB_14__5_), .CO(
        CARRYB_15__4_), .S(SUMB_15__4_) );
  NOR2X4 U2 ( .A(n35), .B(n31), .Y(ab_0__4_) );
  AND2X4 U3 ( .A(A[1]), .B(B[5]), .Y(ab_1__5_) );
  AND2X4 U4 ( .A(n15), .B(B[3]), .Y(ab_2__3_) );
  BUFX16 U5 ( .A(n36), .Y(n24) );
  XOR2X4 U6 ( .A(n3), .B(ab_0__4_), .Y(SUMB_1__3_) );
  AND2X4 U7 ( .A(A[1]), .B(B[4]), .Y(ab_1__4_) );
  BUFX8 U8 ( .A(n35), .Y(n22) );
  BUFX20 U9 ( .A(n38), .Y(n28) );
  CLKBUFXL U10 ( .A(A[1]), .Y(n11) );
  NOR2BX4 U11 ( .AN(A[1]), .B(n24), .Y(n3) );
  NOR2BX2 U12 ( .AN(A[1]), .B(n24), .Y(ab_1__3_) );
  INVX3 U13 ( .A(n26), .Y(n14) );
  AND2X1 U14 ( .A(CARRYB_16__5_), .B(SUMB_16__6_), .Y(n4) );
  NOR2BX1 U15 ( .AN(A[0]), .B(n39), .Y(n32) );
  BUFX20 U16 ( .A(A[2]), .Y(n15) );
  NOR2BX1 U17 ( .AN(A[9]), .B(n23), .Y(ab_9__4_) );
  NOR2BX1 U18 ( .AN(A[9]), .B(n25), .Y(ab_9__3_) );
  NOR2BX1 U19 ( .AN(A[9]), .B(n27), .Y(ab_9__2_) );
  NOR2BX1 U20 ( .AN(A[9]), .B(n29), .Y(ab_9__1_) );
  NOR2BX1 U21 ( .AN(A[12]), .B(n25), .Y(ab_12__3_) );
  NOR2BX1 U22 ( .AN(A[12]), .B(n23), .Y(ab_12__4_) );
  NOR2BX1 U23 ( .AN(A[12]), .B(n27), .Y(ab_12__2_) );
  NOR2BX1 U24 ( .AN(A[12]), .B(n29), .Y(ab_12__1_) );
  NOR2BX1 U25 ( .AN(A[11]), .B(n23), .Y(ab_11__4_) );
  NOR2BX1 U26 ( .AN(A[11]), .B(n25), .Y(ab_11__3_) );
  NOR2BX1 U27 ( .AN(A[11]), .B(n27), .Y(ab_11__2_) );
  NOR2BX1 U28 ( .AN(A[11]), .B(n29), .Y(ab_11__1_) );
  NOR2BX1 U29 ( .AN(A[11]), .B(n39), .Y(ab_11__0_) );
  NOR2BX2 U30 ( .AN(A[11]), .B(n30), .Y(ab_11__6_) );
  AND2X4 U32 ( .A(ab_0__7_), .B(ab_1__6_), .Y(n6) );
  AND2X4 U33 ( .A(ab_0__6_), .B(ab_1__5_), .Y(n7) );
  AND2X4 U34 ( .A(CARRYB_16__1_), .B(SUMB_16__2_), .Y(n8) );
  AND2X4 U35 ( .A(ab_0__3_), .B(ab_1__2_), .Y(n9) );
  AND2X4 U36 ( .A(B[6]), .B(A[0]), .Y(ab_0__6_) );
  INVX16 U37 ( .A(A[0]), .Y(n31) );
  NOR2BXL U38 ( .AN(A[5]), .B(n22), .Y(ab_5__4_) );
  AND2X4 U39 ( .A(ab_0__2_), .B(n41), .Y(n10) );
  NOR2BX2 U40 ( .AN(A[5]), .B(n26), .Y(ab_5__2_) );
  NOR2BX1 U41 ( .AN(A[5]), .B(n30), .Y(ab_5__6_) );
  NOR2BX1 U42 ( .AN(A[5]), .B(n39), .Y(ab_5__0_) );
  NOR2BX2 U43 ( .AN(A[5]), .B(n24), .Y(ab_5__3_) );
  NOR2BX2 U44 ( .AN(n11), .B(n40), .Y(ab_1__7_) );
  NOR2BX1 U45 ( .AN(A[6]), .B(n28), .Y(ab_6__1_) );
  XOR2X4 U46 ( .A(ab_1__4_), .B(ab_0__5_), .Y(SUMB_1__4_) );
  CLKINVX8 U47 ( .A(B[0]), .Y(n39) );
  NOR2BX2 U48 ( .AN(A[8]), .B(n26), .Y(ab_8__2_) );
  NOR2BX1 U49 ( .AN(A[8]), .B(n24), .Y(ab_8__3_) );
  AND2X4 U50 ( .A(ab_1__4_), .B(ab_0__5_), .Y(n12) );
  BUFX16 U51 ( .A(n34), .Y(n20) );
  NOR2BX1 U52 ( .AN(A[6]), .B(n26), .Y(ab_6__2_) );
  AND2X4 U53 ( .A(ab_1__3_), .B(ab_0__4_), .Y(n13) );
  INVX4 U54 ( .A(B[3]), .Y(n36) );
  INVX3 U55 ( .A(B[6]), .Y(n33) );
  NOR2BX4 U56 ( .AN(n15), .B(n39), .Y(ab_2__0_) );
  NOR2BX2 U57 ( .AN(A[3]), .B(n28), .Y(ab_3__1_) );
  NOR2BX2 U58 ( .AN(A[3]), .B(n20), .Y(ab_3__5_) );
  NOR2BX2 U59 ( .AN(A[3]), .B(n24), .Y(ab_3__3_) );
  AND2X4 U60 ( .A(A[1]), .B(n14), .Y(ab_1__2_) );
  NOR2BX2 U61 ( .AN(A[3]), .B(n26), .Y(ab_3__2_) );
  NOR2BX2 U62 ( .AN(A[3]), .B(n39), .Y(ab_3__0_) );
  NOR2BX4 U63 ( .AN(n15), .B(n28), .Y(ab_2__1_) );
  XOR2X4 U64 ( .A(n41), .B(ab_0__2_), .Y(SUMB_1__1_) );
  NOR2BX2 U65 ( .AN(A[3]), .B(n22), .Y(ab_3__4_) );
  XOR2X4 U66 ( .A(ab_1__2_), .B(ab_0__3_), .Y(SUMB_1__2_) );
  BUFX16 U67 ( .A(n37), .Y(n26) );
  CLKINVX8 U68 ( .A(B[2]), .Y(n37) );
  NOR2BX4 U69 ( .AN(n15), .B(n20), .Y(ab_2__5_) );
  NOR2BX2 U70 ( .AN(A[10]), .B(n30), .Y(ab_10__6_) );
  NOR2BX2 U71 ( .AN(A[4]), .B(n22), .Y(ab_4__4_) );
  NOR2BX2 U72 ( .AN(A[4]), .B(n26), .Y(ab_4__2_) );
  NOR2BX4 U73 ( .AN(B[3]), .B(n31), .Y(ab_0__3_) );
  XOR2X2 U74 ( .A(ab_1__6_), .B(ab_0__7_), .Y(SUMB_1__6_) );
  NOR2BX4 U75 ( .AN(B[7]), .B(n31), .Y(ab_0__7_) );
  NOR2BX4 U76 ( .AN(B[2]), .B(n31), .Y(ab_0__2_) );
  NOR2BX4 U77 ( .AN(n15), .B(n22), .Y(ab_2__4_) );
  NOR2BX4 U78 ( .AN(B[5]), .B(n31), .Y(ab_0__5_) );
  NOR2BX1 U79 ( .AN(A[4]), .B(n20), .Y(ab_4__5_) );
  NOR2BX1 U80 ( .AN(A[4]), .B(n39), .Y(ab_4__0_) );
  NOR2BX1 U81 ( .AN(A[4]), .B(n28), .Y(ab_4__1_) );
  NOR2BX1 U82 ( .AN(A[4]), .B(n24), .Y(ab_4__3_) );
  XOR2X4 U83 ( .A(ab_1__5_), .B(ab_0__6_), .Y(SUMB_1__5_) );
  AND2X4 U84 ( .A(CARRYB_16__3_), .B(SUMB_16__4_), .Y(n18) );
  NOR2BX4 U85 ( .AN(n15), .B(n26), .Y(ab_2__2_) );
  BUFX20 U86 ( .A(n33), .Y(n30) );
  NOR2BX4 U87 ( .AN(A[1]), .B(n28), .Y(n41) );
  XOR2X4 U88 ( .A(CARRYB_16__4_), .B(SUMB_16__5_), .Y(A1_19_) );
  AND2X4 U89 ( .A(A[1]), .B(B[6]), .Y(ab_1__6_) );
  AND3X1 U90 ( .A(n32), .B(A[1]), .C(B[1]), .Y(CARRYB_1__0_) );
  AND2X4 U91 ( .A(CARRYB_16__0_), .B(SUMB_16__1_), .Y(n16) );
  INVX4 U92 ( .A(B[1]), .Y(n38) );
  INVX4 U93 ( .A(B[5]), .Y(n34) );
  AND2X2 U94 ( .A(CARRYB_16__2_), .B(SUMB_16__3_), .Y(n17) );
  NOR2BX4 U95 ( .AN(n15), .B(n30), .Y(ab_2__6_) );
  NOR2BX2 U96 ( .AN(A[4]), .B(n30), .Y(ab_4__6_) );
  NOR2BX2 U97 ( .AN(A[6]), .B(n30), .Y(ab_6__6_) );
  NOR2BX2 U98 ( .AN(A[7]), .B(n30), .Y(ab_7__6_) );
  NOR2BX1 U99 ( .AN(A[12]), .B(n39), .Y(ab_12__0_) );
  NOR2BX2 U100 ( .AN(A[3]), .B(n30), .Y(ab_3__6_) );
  NOR2BX1 U101 ( .AN(A[4]), .B(n40), .Y(ab_4__7_) );
  NOR2BX1 U102 ( .AN(A[9]), .B(n40), .Y(ab_9__7_) );
  CLKBUFXL U103 ( .A(n38), .Y(n29) );
  INVX12 U104 ( .A(B[7]), .Y(n40) );
  NOR2BXL U105 ( .AN(A[12]), .B(n40), .Y(ab_12__7_) );
  NOR2BX1 U106 ( .AN(A[7]), .B(n22), .Y(ab_7__4_) );
  NOR2BX1 U107 ( .AN(A[10]), .B(n29), .Y(ab_10__1_) );
  NOR2BX1 U108 ( .AN(A[9]), .B(n39), .Y(ab_9__0_) );
  NOR2BX1 U109 ( .AN(A[7]), .B(n39), .Y(ab_7__0_) );
  NOR2BX1 U110 ( .AN(A[10]), .B(n39), .Y(ab_10__0_) );
  NOR2BX1 U111 ( .AN(A[16]), .B(n39), .Y(ab_16__0_) );
  CLKBUFXL U112 ( .A(n36), .Y(n25) );
  NOR2BX1 U113 ( .AN(A[8]), .B(n28), .Y(ab_8__1_) );
  NOR2BX1 U114 ( .AN(A[10]), .B(n25), .Y(ab_10__3_) );
  NOR2BX1 U115 ( .AN(A[11]), .B(n40), .Y(ab_11__7_) );
  NOR2BXL U116 ( .AN(A[12]), .B(n30), .Y(ab_12__6_) );
  NOR2BX1 U117 ( .AN(A[10]), .B(n27), .Y(ab_10__2_) );
  NOR2BX1 U118 ( .AN(A[8]), .B(n39), .Y(ab_8__0_) );
  NOR2BX1 U119 ( .AN(A[9]), .B(n21), .Y(ab_9__5_) );
  NOR2BXL U120 ( .AN(A[14]), .B(n30), .Y(ab_14__6_) );
  NOR2BXL U121 ( .AN(A[9]), .B(n30), .Y(ab_9__6_) );
  NOR2BX1 U122 ( .AN(A[8]), .B(n40), .Y(ab_8__7_) );
  NOR2BX1 U123 ( .AN(A[6]), .B(n39), .Y(ab_6__0_) );
  NOR2BX1 U124 ( .AN(A[12]), .B(n21), .Y(ab_12__5_) );
  NOR2BX1 U125 ( .AN(A[5]), .B(n28), .Y(ab_5__1_) );
  NOR2BX1 U126 ( .AN(A[11]), .B(n21), .Y(ab_11__5_) );
  CLKBUFXL U127 ( .A(n34), .Y(n21) );
  NOR2BX1 U128 ( .AN(A[16]), .B(n25), .Y(ab_16__3_) );
  NOR2BX1 U129 ( .AN(A[15]), .B(n27), .Y(ab_15__2_) );
  NOR2BX1 U130 ( .AN(A[15]), .B(n25), .Y(ab_15__3_) );
  NOR2BX1 U131 ( .AN(A[3]), .B(n40), .Y(ab_3__7_) );
  NOR2BX1 U132 ( .AN(A[15]), .B(n21), .Y(ab_15__5_) );
  CLKBUFXL U133 ( .A(n35), .Y(n23) );
  BUFX3 U134 ( .A(n37), .Y(n27) );
  NOR2BX1 U135 ( .AN(A[6]), .B(n24), .Y(ab_6__3_) );
  NOR2BXL U136 ( .AN(A[6]), .B(n40), .Y(ab_6__7_) );
  NOR2BX1 U137 ( .AN(A[6]), .B(n22), .Y(ab_6__4_) );
  NOR2BXL U138 ( .AN(A[14]), .B(n29), .Y(ab_14__1_) );
  NOR2BX1 U139 ( .AN(A[8]), .B(n20), .Y(ab_8__5_) );
  NOR2BX1 U140 ( .AN(A[5]), .B(n40), .Y(ab_5__7_) );
  NOR2BX1 U141 ( .AN(A[14]), .B(n23), .Y(ab_14__4_) );
  NOR2BX1 U142 ( .AN(A[13]), .B(n21), .Y(ab_13__5_) );
  NOR2BX1 U143 ( .AN(A[7]), .B(n20), .Y(ab_7__5_) );
  NOR2BX1 U144 ( .AN(A[14]), .B(n21), .Y(ab_14__5_) );
  NOR2BXL U145 ( .AN(A[13]), .B(n40), .Y(ab_13__7_) );
  NOR2BXL U146 ( .AN(A[13]), .B(n27), .Y(ab_13__2_) );
  NOR2BXL U147 ( .AN(A[13]), .B(n25), .Y(ab_13__3_) );
  NOR2BX1 U148 ( .AN(A[10]), .B(n21), .Y(ab_10__5_) );
  NOR2BXL U149 ( .AN(A[7]), .B(n24), .Y(ab_7__3_) );
  NOR2BXL U150 ( .AN(A[14]), .B(n39), .Y(ab_14__0_) );
  NOR2BXL U151 ( .AN(A[13]), .B(n39), .Y(ab_13__0_) );
  NOR2BX1 U152 ( .AN(A[10]), .B(n23), .Y(ab_10__4_) );
  NOR2BXL U153 ( .AN(A[10]), .B(n40), .Y(ab_10__7_) );
  NOR2BXL U154 ( .AN(A[7]), .B(n26), .Y(ab_7__2_) );
  NOR2BX1 U155 ( .AN(A[8]), .B(n22), .Y(ab_8__4_) );
  NOR2BX1 U156 ( .AN(A[5]), .B(n20), .Y(ab_5__5_) );
  NOR2BXL U157 ( .AN(A[14]), .B(n25), .Y(ab_14__3_) );
  NOR2BXL U158 ( .AN(A[13]), .B(n29), .Y(ab_13__1_) );
  NOR2BX1 U159 ( .AN(A[13]), .B(n23), .Y(ab_13__4_) );
  NOR2BX1 U160 ( .AN(A[6]), .B(n20), .Y(ab_6__5_) );
  NOR2BXL U161 ( .AN(A[14]), .B(n27), .Y(ab_14__2_) );
  NOR2BXL U162 ( .AN(A[7]), .B(n28), .Y(ab_7__1_) );
  NOR2BXL U163 ( .AN(A[13]), .B(n30), .Y(ab_13__6_) );
  NOR2BXL U164 ( .AN(A[7]), .B(n40), .Y(ab_7__7_) );
  NOR2BXL U165 ( .AN(A[8]), .B(n30), .Y(ab_8__6_) );
  AND2X2 U166 ( .A(CARRYB_16__4_), .B(SUMB_16__5_), .Y(n19) );
  NOR2BX1 U167 ( .AN(A[16]), .B(n23), .Y(ab_16__4_) );
  NOR2BX1 U168 ( .AN(A[16]), .B(n21), .Y(ab_16__5_) );
  NOR2BX1 U169 ( .AN(A[16]), .B(n29), .Y(ab_16__1_) );
  NOR2BX1 U170 ( .AN(A[16]), .B(n27), .Y(ab_16__2_) );
  NOR2BX1 U171 ( .AN(A[15]), .B(n23), .Y(ab_15__4_) );
  NOR2BXL U172 ( .AN(A[15]), .B(n30), .Y(ab_15__6_) );
  NOR2BXL U173 ( .AN(A[14]), .B(n40), .Y(ab_14__7_) );
  NOR2BXL U174 ( .AN(A[15]), .B(n39), .Y(ab_15__0_) );
  NOR2BXL U175 ( .AN(A[15]), .B(n29), .Y(ab_15__1_) );
  NOR2BXL U176 ( .AN(A[15]), .B(n40), .Y(ab_15__7_) );
  NOR2BXL U177 ( .AN(A[16]), .B(n30), .Y(ab_16__6_) );
  NOR2BXL U178 ( .AN(A[16]), .B(n40), .Y(ab_16__7_) );
  XOR2X4 U179 ( .A(CARRYB_16__3_), .B(SUMB_16__4_), .Y(A1_18_) );
  XOR2X4 U180 ( .A(CARRYB_16__5_), .B(SUMB_16__6_), .Y(A1_20_) );
  XOR2X4 U181 ( .A(CARRYB_16__6_), .B(ab_16__7_), .Y(A1_21_) );
  XOR2X4 U182 ( .A(SUMB_16__2_), .B(CARRYB_16__1_), .Y(A1_16_) );
  XOR2X4 U183 ( .A(SUMB_16__3_), .B(CARRYB_16__2_), .Y(A1_17_) );
  XOR2X4 U184 ( .A(SUMB_16__1_), .B(CARRYB_16__0_), .Y(A1_15_) );
  NOR2BX1 U185 ( .AN(n15), .B(n40), .Y(ab_2__7_) );
  INVX8 U186 ( .A(B[4]), .Y(n35) );
endmodule


module multi16_9 ( in_17bit, in_8bit, out );
  input [16:0] in_17bit;
  input [7:0] in_8bit;
  output [16:0] out;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115;
  wire   [16:1] in_17bit_b;
  wire   [7:1] in_8bit_b;
  wire   [23:8] mul;

  multi16_9_DW02_mult_0 mult_55 ( .A({in_17bit_b[16:2], n35, n12}), .B({
        in_8bit_b, n14}), .PRODUCT_23_(mul[23]), .PRODUCT_22_(mul[22]), 
        .PRODUCT_21_(mul[21]), .PRODUCT_20_(mul[20]), .PRODUCT_19_(mul[19]), 
        .PRODUCT_18_(mul[18]), .PRODUCT_17_(mul[17]), .PRODUCT_16_(mul[16]), 
        .PRODUCT_15_(mul[15]), .PRODUCT_14_(mul[14]), .PRODUCT_13_(mul[13]), 
        .PRODUCT_12_(mul[12]), .PRODUCT_11_(mul[11]), .PRODUCT_10_(mul[10]), 
        .PRODUCT_9_(mul[9]), .PRODUCT_8_(mul[8]), .PRODUCT_7_(out[0]) );
  CLKINVX1 U2 ( .A(n82), .Y(n7) );
  INVX3 U3 ( .A(in_17bit[1]), .Y(n52) );
  XOR2X4 U4 ( .A(n1), .B(n2), .Y(in_8bit_b[6]) );
  CLKINVX20 U5 ( .A(in_8bit[6]), .Y(n1) );
  NAND2X4 U6 ( .A(n37), .B(n51), .Y(n2) );
  CLKINVX4 U7 ( .A(n101), .Y(n106) );
  INVX4 U8 ( .A(n82), .Y(n3) );
  NOR2XL U9 ( .A(mul[22]), .B(mul[21]), .Y(n114) );
  INVX2 U10 ( .A(mul[20]), .Y(n104) );
  BUFX20 U11 ( .A(in_17bit[16]), .Y(n36) );
  INVXL U12 ( .A(in_17bit[9]), .Y(n70) );
  CLKINVX2 U13 ( .A(in_17bit[5]), .Y(n61) );
  INVXL U14 ( .A(in_17bit[13]), .Y(n79) );
  INVX20 U15 ( .A(n112), .Y(n108) );
  INVX3 U16 ( .A(in_17bit[2]), .Y(n55) );
  INVX8 U17 ( .A(n3), .Y(n4) );
  INVX1 U18 ( .A(n97), .Y(n6) );
  INVX2 U19 ( .A(n75), .Y(n29) );
  NOR2X2 U20 ( .A(n78), .B(in_17bit[13]), .Y(n27) );
  NAND2X2 U21 ( .A(n89), .B(n108), .Y(n88) );
  INVX1 U22 ( .A(mul[18]), .Y(n105) );
  NOR2X4 U23 ( .A(n34), .B(n38), .Y(n23) );
  XNOR2X4 U24 ( .A(mul[17]), .B(n5), .Y(out[10]) );
  NAND2X4 U25 ( .A(n98), .B(n108), .Y(n5) );
  NOR2XL U26 ( .A(n24), .B(n4), .Y(n66) );
  AOI31X2 U27 ( .A0(n48), .A1(n41), .A2(n43), .B0(n40), .Y(n49) );
  INVX1 U28 ( .A(in_8bit[1]), .Y(n41) );
  NAND2X4 U29 ( .A(n7), .B(n60), .Y(n59) );
  NAND2BX4 U30 ( .AN(mul[16]), .B(n6), .Y(n98) );
  NOR4X4 U31 ( .A(in_8bit[1]), .B(in_8bit[0]), .C(in_8bit[4]), .D(in_8bit[3]), 
        .Y(n9) );
  INVX8 U32 ( .A(in_8bit[2]), .Y(n43) );
  INVX4 U33 ( .A(in_17bit[4]), .Y(n58) );
  XNOR2X4 U34 ( .A(n62), .B(n63), .Y(in_17bit_b[6]) );
  NOR2XL U35 ( .A(n26), .B(n4), .Y(n62) );
  INVX1 U36 ( .A(in_8bit[5]), .Y(n50) );
  BUFX1 U37 ( .A(n113), .Y(n8) );
  INVX4 U38 ( .A(n13), .Y(n14) );
  INVX8 U39 ( .A(n43), .Y(n42) );
  XNOR2X4 U40 ( .A(n66), .B(n67), .Y(in_17bit_b[8]) );
  NOR2X4 U41 ( .A(n64), .B(n25), .Y(n24) );
  NAND2X4 U42 ( .A(n26), .B(n63), .Y(n64) );
  XNOR2X2 U43 ( .A(n47), .B(in_8bit[3]), .Y(in_8bit_b[3]) );
  AND2X4 U44 ( .A(n9), .B(n43), .Y(n34) );
  CLKINVX8 U45 ( .A(n11), .Y(n12) );
  NOR2X4 U46 ( .A(n113), .B(n10), .Y(n107) );
  CLKINVX20 U47 ( .A(n108), .Y(n10) );
  NOR2XL U48 ( .A(n28), .B(n4), .Y(n76) );
  XOR2X2 U49 ( .A(mul[8]), .B(n16), .Y(out[1]) );
  XOR2X4 U50 ( .A(n42), .B(n45), .Y(in_8bit_b[2]) );
  NOR2X2 U51 ( .A(n32), .B(n82), .Y(n20) );
  AOI21X1 U52 ( .A0(n114), .A1(n8), .B0(n112), .Y(n115) );
  XNOR2X4 U53 ( .A(n71), .B(n72), .Y(in_17bit_b[10]) );
  NOR2XL U54 ( .A(n30), .B(n4), .Y(n71) );
  NAND2X2 U55 ( .A(n91), .B(n108), .Y(n17) );
  NAND2X2 U56 ( .A(n3), .B(n57), .Y(n56) );
  NOR2X4 U57 ( .A(n31), .B(n82), .Y(n54) );
  XNOR2X2 U58 ( .A(mul[10]), .B(n86), .Y(out[3]) );
  OAI21X4 U59 ( .A0(mul[21]), .A1(n109), .B0(n108), .Y(n110) );
  INVX8 U60 ( .A(n109), .Y(n113) );
  NOR2X4 U61 ( .A(in_17bit[3]), .B(n57), .Y(n32) );
  NAND2X4 U62 ( .A(n31), .B(n55), .Y(n57) );
  NAND2X4 U63 ( .A(n32), .B(n58), .Y(n60) );
  NOR2X4 U64 ( .A(n44), .B(n38), .Y(n45) );
  INVX4 U65 ( .A(n46), .Y(n44) );
  INVX12 U66 ( .A(in_8bit[7]), .Y(n38) );
  INVX2 U67 ( .A(in_17bit[0]), .Y(n11) );
  XOR2X2 U68 ( .A(mul[23]), .B(n115), .Y(out[16]) );
  INVXL U69 ( .A(in_8bit[0]), .Y(n13) );
  NOR2XL U70 ( .A(in_8bit[0]), .B(in_8bit[3]), .Y(n48) );
  NOR3X2 U71 ( .A(n51), .B(in_8bit[6]), .C(n39), .Y(in_8bit_b[7]) );
  NOR2X4 U72 ( .A(in_17bit[0]), .B(in_17bit[1]), .Y(n31) );
  OAI21X2 U73 ( .A0(mul[18]), .A1(n101), .B0(n108), .Y(n100) );
  NAND2X4 U74 ( .A(n36), .B(in_17bit[0]), .Y(n53) );
  XNOR2X4 U75 ( .A(mul[9]), .B(n84), .Y(out[2]) );
  NAND2X2 U76 ( .A(n85), .B(n108), .Y(n84) );
  BUFX12 U77 ( .A(in_17bit_b[1]), .Y(n35) );
  XNOR2X2 U78 ( .A(mul[13]), .B(n17), .Y(out[6]) );
  OAI21X4 U79 ( .A0(n102), .A1(mul[19]), .B0(n108), .Y(n103) );
  XOR2X4 U80 ( .A(n41), .B(n19), .Y(in_8bit_b[1]) );
  NAND2X2 U81 ( .A(n14), .B(n37), .Y(n19) );
  INVX8 U82 ( .A(in_8bit[7]), .Y(n39) );
  INVX8 U83 ( .A(n36), .Y(n82) );
  XNOR2X2 U84 ( .A(mul[11]), .B(n88), .Y(out[4]) );
  XNOR2X4 U85 ( .A(in_17bit[3]), .B(n56), .Y(in_17bit_b[3]) );
  OR2X4 U86 ( .A(in_8bit[1]), .B(in_8bit[0]), .Y(n46) );
  XOR2X2 U87 ( .A(mul[12]), .B(n15), .Y(out[5]) );
  XNOR2X4 U88 ( .A(n23), .B(n50), .Y(in_8bit_b[5]) );
  XNOR2X4 U89 ( .A(mul[15]), .B(n18), .Y(out[8]) );
  OR2X4 U90 ( .A(mul[14]), .B(n93), .Y(n94) );
  AOI32X2 U91 ( .A0(n36), .A1(in_17bit[0]), .A2(in_17bit[1]), .B0(n53), .B1(
        n52), .Y(in_17bit_b[1]) );
  NOR3X1 U92 ( .A(in_17bit[15]), .B(n83), .C(n4), .Y(in_17bit_b[16]) );
  XNOR2X4 U93 ( .A(mul[14]), .B(n92), .Y(out[7]) );
  NOR2X4 U94 ( .A(n60), .B(in_17bit[5]), .Y(n26) );
  NAND2X4 U95 ( .A(n101), .B(n108), .Y(n99) );
  NOR2X1 U96 ( .A(n69), .B(in_17bit[9]), .Y(n30) );
  NAND2X4 U97 ( .A(n93), .B(n108), .Y(n92) );
  NAND2X2 U98 ( .A(n94), .B(n108), .Y(n18) );
  XNOR2X4 U99 ( .A(n20), .B(n58), .Y(in_17bit_b[4]) );
  NAND2XL U100 ( .A(n7), .B(n78), .Y(n22) );
  OR2X4 U101 ( .A(mul[11]), .B(n89), .Y(n90) );
  AND2X4 U102 ( .A(n90), .B(n108), .Y(n15) );
  AND2X1 U103 ( .A(out[0]), .B(n108), .Y(n16) );
  NOR2X4 U104 ( .A(n74), .B(n29), .Y(n28) );
  XNOR2X4 U105 ( .A(n80), .B(n81), .Y(in_17bit_b[14]) );
  NAND2XL U106 ( .A(n24), .B(n67), .Y(n69) );
  OR2X4 U107 ( .A(mul[10]), .B(n87), .Y(n89) );
  OR2X4 U108 ( .A(mul[9]), .B(n85), .Y(n87) );
  OR2X4 U109 ( .A(mul[13]), .B(n91), .Y(n93) );
  OR2X4 U110 ( .A(mul[8]), .B(out[0]), .Y(n85) );
  OR2X4 U111 ( .A(mul[12]), .B(n90), .Y(n91) );
  OR2X4 U112 ( .A(mul[17]), .B(n98), .Y(n101) );
  INVX4 U113 ( .A(n39), .Y(n37) );
  XOR2X2 U114 ( .A(n65), .B(n21), .Y(in_17bit_b[7]) );
  NAND2XL U115 ( .A(n7), .B(n64), .Y(n21) );
  CLKINVX3 U116 ( .A(n65), .Y(n25) );
  XOR2X2 U117 ( .A(n79), .B(n22), .Y(in_17bit_b[13]) );
  INVX2 U118 ( .A(mul[22]), .Y(n111) );
  NAND2X1 U119 ( .A(n87), .B(n108), .Y(n86) );
  XNOR2X1 U120 ( .A(n3), .B(n37), .Y(n112) );
  NAND2XL U121 ( .A(n7), .B(n74), .Y(n73) );
  NAND2XL U122 ( .A(n3), .B(n69), .Y(n68) );
  NAND2XL U123 ( .A(n28), .B(n77), .Y(n78) );
  NAND2X2 U124 ( .A(n30), .B(n72), .Y(n74) );
  XOR2X2 U125 ( .A(in_17bit[15]), .B(n33), .Y(in_17bit_b[15]) );
  AND2X1 U126 ( .A(n3), .B(n83), .Y(n33) );
  INVXL U127 ( .A(in_8bit[7]), .Y(n40) );
  NAND2BX2 U128 ( .AN(mul[18]), .B(n106), .Y(n102) );
  NOR2XL U129 ( .A(n27), .B(n4), .Y(n80) );
  OAI21X4 U130 ( .A0(n42), .A1(n46), .B0(n37), .Y(n47) );
  XOR2X4 U131 ( .A(n49), .B(in_8bit[4]), .Y(in_8bit_b[4]) );
  NAND2X4 U132 ( .A(n34), .B(n50), .Y(n51) );
  XNOR2X4 U133 ( .A(n54), .B(n55), .Y(in_17bit_b[2]) );
  XOR2X4 U134 ( .A(n61), .B(n59), .Y(in_17bit_b[5]) );
  CLKINVX3 U135 ( .A(in_17bit[6]), .Y(n63) );
  CLKINVX3 U136 ( .A(in_17bit[7]), .Y(n65) );
  CLKINVX3 U137 ( .A(in_17bit[8]), .Y(n67) );
  XOR2X4 U138 ( .A(n70), .B(n68), .Y(in_17bit_b[9]) );
  CLKINVX3 U139 ( .A(in_17bit[10]), .Y(n72) );
  CLKINVX3 U140 ( .A(in_17bit[11]), .Y(n75) );
  XOR2X4 U141 ( .A(n75), .B(n73), .Y(in_17bit_b[11]) );
  CLKINVX3 U142 ( .A(in_17bit[12]), .Y(n77) );
  XNOR2X4 U143 ( .A(n76), .B(n77), .Y(in_17bit_b[12]) );
  CLKINVX3 U144 ( .A(in_17bit[14]), .Y(n81) );
  NAND2X4 U145 ( .A(n27), .B(n81), .Y(n83) );
  CLKINVX3 U146 ( .A(n94), .Y(n95) );
  NAND2BX4 U147 ( .AN(mul[15]), .B(n95), .Y(n97) );
  NAND2X4 U148 ( .A(n97), .B(n108), .Y(n96) );
  XNOR2X4 U149 ( .A(mul[16]), .B(n96), .Y(out[9]) );
  XNOR2X4 U150 ( .A(n99), .B(mul[18]), .Y(out[11]) );
  XNOR2X4 U151 ( .A(mul[19]), .B(n100), .Y(out[12]) );
  XOR2X4 U152 ( .A(n104), .B(n103), .Y(out[13]) );
  NAND4BBX4 U153 ( .AN(mul[20]), .BN(mul[19]), .C(n106), .D(n105), .Y(n109) );
  XOR2X4 U154 ( .A(n107), .B(mul[21]), .Y(out[14]) );
  XOR2X4 U155 ( .A(n111), .B(n110), .Y(out[15]) );
endmodule


module multi16_8_DW01_add_5 ( A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, 
        A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, 
        B_20_, B_19_, B_18_, B_17_, B_16_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, 
        SUM_17_, SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, 
        SUM_9_, SUM_8_, SUM_7_, SUM_6_, SUM_5_ );
  input A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_,
         A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, B_20_, B_19_,
         B_18_, B_17_, B_16_;
  output SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, SUM_15_,
         SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, SUM_7_,
         SUM_6_, SUM_5_;
  wire   n1, n2, n3, n4, n6, n7, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44;

  INVX2 U2 ( .A(n33), .Y(n43) );
  NOR2X2 U3 ( .A(A_17_), .B(B_17_), .Y(n3) );
  NAND2X2 U4 ( .A(n20), .B(n21), .Y(n19) );
  AND2X4 U5 ( .A(A_16_), .B(B_16_), .Y(n2) );
  CLKBUFX8 U6 ( .A(n32), .Y(n1) );
  NOR2X2 U7 ( .A(n7), .B(n6), .Y(n30) );
  BUFX12 U8 ( .A(A_15_), .Y(SUM_15_) );
  NAND2X4 U9 ( .A(B_16_), .B(A_16_), .Y(n33) );
  OR2X4 U10 ( .A(A_16_), .B(B_16_), .Y(n4) );
  INVX4 U11 ( .A(n39), .Y(n38) );
  NAND2XL U12 ( .A(n31), .B(n1), .Y(n29) );
  BUFX12 U13 ( .A(A_14_), .Y(SUM_14_) );
  NAND2X4 U14 ( .A(n2), .B(n42), .Y(n41) );
  OAI21X4 U15 ( .A0(n38), .A1(n6), .B0(n31), .Y(n36) );
  NAND2X4 U16 ( .A(B_17_), .B(A_17_), .Y(n32) );
  NOR2BX4 U17 ( .AN(n35), .B(n7), .Y(n37) );
  XOR2X4 U18 ( .A(n36), .B(n37), .Y(SUM_19_) );
  XOR2X4 U19 ( .A(n39), .B(n40), .Y(SUM_18_) );
  BUFX12 U20 ( .A(A_10_), .Y(SUM_10_) );
  NOR2BX4 U21 ( .AN(n31), .B(n6), .Y(n40) );
  NOR2X4 U22 ( .A(A_19_), .B(B_19_), .Y(n7) );
  NAND2X2 U23 ( .A(B_19_), .B(A_19_), .Y(n35) );
  NOR2X4 U24 ( .A(A_18_), .B(B_18_), .Y(n6) );
  AND2X4 U25 ( .A(n33), .B(n4), .Y(SUM_16_) );
  NAND2X4 U26 ( .A(B_18_), .B(A_18_), .Y(n31) );
  INVX1 U27 ( .A(n34), .Y(n26) );
  OAI21X2 U28 ( .A0(n28), .A1(n29), .B0(n30), .Y(n27) );
  INVX1 U29 ( .A(n35), .Y(n34) );
  NAND2XL U30 ( .A(n22), .B(n23), .Y(n21) );
  NAND2X4 U31 ( .A(n1), .B(n41), .Y(n39) );
  BUFX4 U32 ( .A(A_7_), .Y(SUM_7_) );
  BUFX8 U33 ( .A(A_12_), .Y(SUM_12_) );
  BUFX8 U34 ( .A(A_11_), .Y(SUM_11_) );
  BUFX8 U35 ( .A(A_9_), .Y(SUM_9_) );
  BUFX8 U36 ( .A(A_8_), .Y(SUM_8_) );
  NAND2X2 U37 ( .A(B_20_), .B(A_20_), .Y(n20) );
  BUFX8 U38 ( .A(A_5_), .Y(SUM_5_) );
  BUFX4 U39 ( .A(A_6_), .Y(SUM_6_) );
  BUFX8 U40 ( .A(A_13_), .Y(SUM_13_) );
  NOR2XL U41 ( .A(n33), .B(n3), .Y(n28) );
  XOR3X4 U42 ( .A(B_21_), .B(A_21_), .C(n19), .Y(SUM_21_) );
  XOR2X4 U43 ( .A(n22), .B(n24), .Y(SUM_20_) );
  NOR2BX4 U44 ( .AN(n20), .B(n25), .Y(n24) );
  CLKINVX3 U45 ( .A(n23), .Y(n25) );
  OR2X4 U46 ( .A(A_20_), .B(B_20_), .Y(n23) );
  NAND2X4 U47 ( .A(n26), .B(n27), .Y(n22) );
  XOR2X4 U48 ( .A(n44), .B(n43), .Y(SUM_17_) );
  NOR2BX4 U49 ( .AN(n32), .B(n3), .Y(n44) );
  OR2X4 U50 ( .A(A_17_), .B(B_17_), .Y(n42) );
endmodule


module multi16_8_DW02_mult_0 ( A, B, PRODUCT_23_, PRODUCT_22_, PRODUCT_21_, 
        PRODUCT_20_, PRODUCT_19_, PRODUCT_18_, PRODUCT_17_, PRODUCT_16_, 
        PRODUCT_15_, PRODUCT_14_, PRODUCT_13_, PRODUCT_12_, PRODUCT_11_, 
        PRODUCT_10_, PRODUCT_9_, PRODUCT_8_, PRODUCT_7_ );
  input [16:0] A;
  input [7:0] B;
  output PRODUCT_23_, PRODUCT_22_, PRODUCT_21_, PRODUCT_20_, PRODUCT_19_,
         PRODUCT_18_, PRODUCT_17_, PRODUCT_16_, PRODUCT_15_, PRODUCT_14_,
         PRODUCT_13_, PRODUCT_12_, PRODUCT_11_, PRODUCT_10_, PRODUCT_9_,
         PRODUCT_8_, PRODUCT_7_;
  wire   ab_16__7_, ab_16__6_, ab_16__5_, ab_16__4_, ab_16__3_, ab_16__2_,
         ab_16__1_, ab_16__0_, ab_15__7_, ab_15__6_, ab_15__5_, ab_15__4_,
         ab_15__3_, ab_15__2_, ab_15__1_, ab_15__0_, ab_14__7_, ab_14__6_,
         ab_14__5_, ab_14__4_, ab_14__3_, ab_14__2_, ab_14__1_, ab_14__0_,
         ab_13__7_, ab_13__6_, ab_13__5_, ab_13__4_, ab_13__3_, ab_13__2_,
         ab_13__1_, ab_13__0_, ab_12__7_, ab_12__6_, ab_12__5_, ab_12__4_,
         ab_12__3_, ab_12__2_, ab_12__1_, ab_12__0_, ab_11__7_, ab_11__6_,
         ab_11__5_, ab_11__4_, ab_11__3_, ab_11__2_, ab_11__1_, ab_11__0_,
         ab_10__7_, ab_10__6_, ab_10__5_, ab_10__4_, ab_10__3_, ab_10__2_,
         ab_10__1_, ab_10__0_, ab_9__7_, ab_9__6_, ab_9__5_, ab_9__4_,
         ab_9__3_, ab_9__2_, ab_9__1_, ab_9__0_, ab_8__7_, ab_8__6_, ab_8__5_,
         ab_8__4_, ab_8__3_, ab_8__2_, ab_8__1_, ab_8__0_, ab_7__7_, ab_7__6_,
         ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_, ab_7__0_, ab_6__7_,
         ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_, ab_6__1_, ab_6__0_,
         ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_, ab_5__2_, ab_5__1_,
         ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_, ab_4__3_, ab_4__2_,
         ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_, ab_3__4_, ab_3__3_,
         ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_, ab_2__5_, ab_2__4_,
         ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_, ab_1__6_, ab_1__5_,
         ab_1__4_, ab_1__3_, ab_1__2_, ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_,
         ab_0__3_, ab_0__2_, CARRYB_16__6_, CARRYB_16__5_, CARRYB_16__4_,
         CARRYB_16__3_, CARRYB_16__2_, CARRYB_16__1_, CARRYB_16__0_,
         CARRYB_15__6_, CARRYB_15__5_, CARRYB_15__4_, CARRYB_15__3_,
         CARRYB_15__2_, CARRYB_15__1_, CARRYB_15__0_, CARRYB_14__6_,
         CARRYB_14__5_, CARRYB_14__4_, CARRYB_14__3_, CARRYB_14__2_,
         CARRYB_14__1_, CARRYB_14__0_, CARRYB_13__6_, CARRYB_13__5_,
         CARRYB_13__4_, CARRYB_13__3_, CARRYB_13__2_, CARRYB_13__1_,
         CARRYB_13__0_, CARRYB_12__6_, CARRYB_12__5_, CARRYB_12__4_,
         CARRYB_12__3_, CARRYB_12__2_, CARRYB_12__1_, CARRYB_12__0_,
         CARRYB_11__6_, CARRYB_11__5_, CARRYB_11__4_, CARRYB_11__3_,
         CARRYB_11__2_, CARRYB_11__1_, CARRYB_11__0_, CARRYB_10__6_,
         CARRYB_10__5_, CARRYB_10__4_, CARRYB_10__3_, CARRYB_10__2_,
         CARRYB_10__1_, CARRYB_10__0_, CARRYB_9__6_, CARRYB_9__5_,
         CARRYB_9__4_, CARRYB_9__3_, CARRYB_9__2_, CARRYB_9__1_, CARRYB_9__0_,
         CARRYB_8__6_, CARRYB_8__5_, CARRYB_8__4_, CARRYB_8__3_, CARRYB_8__2_,
         CARRYB_8__1_, CARRYB_8__0_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_,
         CARRYB_7__3_, CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_,
         CARRYB_6__5_, CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_,
         CARRYB_6__0_, CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_,
         CARRYB_5__2_, CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_,
         CARRYB_4__4_, CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_,
         CARRYB_3__6_, CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_,
         CARRYB_3__1_, CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_,
         CARRYB_2__3_, CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__1_,
         CARRYB_1__0_, SUMB_16__6_, SUMB_16__5_, SUMB_16__4_, SUMB_16__3_,
         SUMB_16__2_, SUMB_16__1_, SUMB_16__0_, SUMB_15__6_, SUMB_15__5_,
         SUMB_15__4_, SUMB_15__3_, SUMB_15__2_, SUMB_15__1_, SUMB_14__6_,
         SUMB_14__5_, SUMB_14__4_, SUMB_14__3_, SUMB_14__2_, SUMB_14__1_,
         SUMB_13__6_, SUMB_13__5_, SUMB_13__4_, SUMB_13__3_, SUMB_13__2_,
         SUMB_13__1_, SUMB_12__6_, SUMB_12__5_, SUMB_12__4_, SUMB_12__3_,
         SUMB_12__2_, SUMB_12__1_, SUMB_11__6_, SUMB_11__5_, SUMB_11__4_,
         SUMB_11__3_, SUMB_11__2_, SUMB_11__1_, SUMB_10__6_, SUMB_10__5_,
         SUMB_10__4_, SUMB_10__3_, SUMB_10__2_, SUMB_10__1_, SUMB_9__6_,
         SUMB_9__5_, SUMB_9__4_, SUMB_9__3_, SUMB_9__2_, SUMB_9__1_,
         SUMB_8__6_, SUMB_8__5_, SUMB_8__4_, SUMB_8__3_, SUMB_8__2_,
         SUMB_8__1_, SUMB_7__6_, SUMB_7__5_, SUMB_7__4_, SUMB_7__3_,
         SUMB_7__2_, SUMB_7__1_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_,
         SUMB_6__3_, SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_,
         SUMB_5__4_, SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_,
         SUMB_4__5_, SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_,
         SUMB_3__6_, SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_,
         SUMB_3__1_, SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_,
         SUMB_2__2_, SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_,
         SUMB_1__3_, SUMB_1__2_, SUMB_1__1_, PROD1_7_, A1_21_, A1_20_, A1_19_,
         A1_18_, A1_17_, A1_16_, A1_15_, A1_13_, A1_12_, A1_11_, A1_10_, A1_9_,
         A1_8_, A1_7_, A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, n3, n4, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43;

  ADDFHX2 S5_6 ( .A(ab_16__6_), .B(CARRYB_15__6_), .CI(ab_15__7_), .CO(
        CARRYB_16__6_), .S(SUMB_16__6_) );
  ADDFHX2 S2_15_5 ( .A(ab_15__5_), .B(CARRYB_14__5_), .CI(SUMB_14__6_), .CO(
        CARRYB_15__5_), .S(SUMB_15__5_) );
  multi16_8_DW01_add_5 FS_1 ( .A_21_(A1_21_), .A_20_(A1_20_), .A_19_(A1_19_), 
        .A_18_(A1_18_), .A_17_(A1_17_), .A_16_(A1_16_), .A_15_(A1_15_), 
        .A_14_(SUMB_16__0_), .A_13_(A1_13_), .A_12_(A1_12_), .A_11_(A1_11_), 
        .A_10_(A1_10_), .A_9_(A1_9_), .A_8_(A1_8_), .A_7_(A1_7_), .A_6_(A1_6_), 
        .A_5_(PROD1_7_), .B_21_(n20), .B_20_(n19), .B_19_(n17), .B_18_(n18), 
        .B_17_(n7), .B_16_(n16), .SUM_21_(PRODUCT_23_), .SUM_20_(PRODUCT_22_), 
        .SUM_19_(PRODUCT_21_), .SUM_18_(PRODUCT_20_), .SUM_17_(PRODUCT_19_), 
        .SUM_16_(PRODUCT_18_), .SUM_15_(PRODUCT_17_), .SUM_14_(PRODUCT_16_), 
        .SUM_13_(PRODUCT_15_), .SUM_12_(PRODUCT_14_), .SUM_11_(PRODUCT_13_), 
        .SUM_10_(PRODUCT_12_), .SUM_9_(PRODUCT_11_), .SUM_8_(PRODUCT_10_), 
        .SUM_7_(PRODUCT_9_), .SUM_6_(PRODUCT_8_), .SUM_5_(PRODUCT_7_) );
  ADDFHX4 S4_1 ( .A(ab_16__1_), .B(CARRYB_15__1_), .CI(SUMB_15__2_), .CO(
        CARRYB_16__1_), .S(SUMB_16__1_) );
  ADDFHX4 S4_2 ( .A(ab_16__2_), .B(CARRYB_15__2_), .CI(SUMB_15__3_), .CO(
        CARRYB_16__2_), .S(SUMB_16__2_) );
  ADDFHX4 S4_3 ( .A(ab_16__3_), .B(SUMB_15__4_), .CI(CARRYB_15__3_), .CO(
        CARRYB_16__3_), .S(SUMB_16__3_) );
  ADDFHX4 S2_11_1 ( .A(ab_11__1_), .B(CARRYB_10__1_), .CI(SUMB_10__2_), .CO(
        CARRYB_11__1_), .S(SUMB_11__1_) );
  ADDFHX4 S2_12_2 ( .A(ab_12__2_), .B(CARRYB_11__2_), .CI(SUMB_11__3_), .CO(
        CARRYB_12__2_), .S(SUMB_12__2_) );
  ADDFHX4 S2_13_2 ( .A(ab_13__2_), .B(CARRYB_12__2_), .CI(SUMB_12__3_), .CO(
        CARRYB_13__2_), .S(SUMB_13__2_) );
  ADDFHX4 S2_14_3 ( .A(ab_14__3_), .B(CARRYB_13__3_), .CI(SUMB_13__4_), .CO(
        CARRYB_14__3_), .S(SUMB_14__3_) );
  ADDFHX4 S2_15_2 ( .A(ab_15__2_), .B(CARRYB_14__2_), .CI(SUMB_14__3_), .CO(
        CARRYB_15__2_), .S(SUMB_15__2_) );
  ADDFHX4 S2_9_2 ( .A(ab_9__2_), .B(CARRYB_8__2_), .CI(SUMB_8__3_), .CO(
        CARRYB_9__2_), .S(SUMB_9__2_) );
  ADDFHX4 S1_14_0 ( .A(ab_14__0_), .B(CARRYB_13__0_), .CI(SUMB_13__1_), .CO(
        CARRYB_14__0_), .S(A1_12_) );
  ADDFHX4 S1_15_0 ( .A(ab_15__0_), .B(CARRYB_14__0_), .CI(SUMB_14__1_), .CO(
        CARRYB_15__0_), .S(A1_13_) );
  ADDFHX4 S2_12_1 ( .A(ab_12__1_), .B(CARRYB_11__1_), .CI(SUMB_11__2_), .CO(
        CARRYB_12__1_), .S(SUMB_12__1_) );
  ADDFHX4 S2_13_1 ( .A(ab_13__1_), .B(CARRYB_12__1_), .CI(SUMB_12__2_), .CO(
        CARRYB_13__1_), .S(SUMB_13__1_) );
  ADDFHX4 S1_12_0 ( .A(ab_12__0_), .B(CARRYB_11__0_), .CI(SUMB_11__1_), .CO(
        CARRYB_12__0_), .S(A1_10_) );
  ADDFHX4 S1_13_0 ( .A(ab_13__0_), .B(CARRYB_12__0_), .CI(SUMB_12__1_), .CO(
        CARRYB_13__0_), .S(A1_11_) );
  ADDFHX4 S2_12_4 ( .A(ab_12__4_), .B(CARRYB_11__4_), .CI(SUMB_11__5_), .CO(
        CARRYB_12__4_), .S(SUMB_12__4_) );
  ADDFHX4 S2_10_4 ( .A(ab_10__4_), .B(CARRYB_9__4_), .CI(SUMB_9__5_), .CO(
        CARRYB_10__4_), .S(SUMB_10__4_) );
  ADDFHX4 S2_11_4 ( .A(ab_11__4_), .B(CARRYB_10__4_), .CI(SUMB_10__5_), .CO(
        CARRYB_11__4_), .S(SUMB_11__4_) );
  ADDFHX4 S4_0 ( .A(ab_16__0_), .B(CARRYB_15__0_), .CI(SUMB_15__1_), .CO(
        CARRYB_16__0_), .S(SUMB_16__0_) );
  ADDFHX4 S2_10_3 ( .A(ab_10__3_), .B(CARRYB_9__3_), .CI(SUMB_9__4_), .CO(
        CARRYB_10__3_), .S(SUMB_10__3_) );
  ADDFHX4 S2_11_3 ( .A(ab_11__3_), .B(CARRYB_10__3_), .CI(SUMB_10__4_), .CO(
        CARRYB_11__3_), .S(SUMB_11__3_) );
  ADDFHX4 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  ADDFHX4 S1_11_0 ( .A(ab_11__0_), .B(SUMB_10__1_), .CI(CARRYB_10__0_), .CO(
        CARRYB_11__0_), .S(A1_9_) );
  ADDFHX4 S1_7_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(PROD1_7_) );
  ADDFHX4 S1_8_0 ( .A(ab_8__0_), .B(CARRYB_7__0_), .CI(SUMB_7__1_), .CO(
        CARRYB_8__0_), .S(A1_6_) );
  ADDFHX4 S2_12_3 ( .A(ab_12__3_), .B(CARRYB_11__3_), .CI(SUMB_11__4_), .CO(
        CARRYB_12__3_), .S(SUMB_12__3_) );
  ADDFHX4 S2_10_1 ( .A(ab_10__1_), .B(CARRYB_9__1_), .CI(SUMB_9__2_), .CO(
        CARRYB_10__1_), .S(SUMB_10__1_) );
  ADDFHX1 S3_15_6 ( .A(ab_15__6_), .B(CARRYB_14__6_), .CI(ab_14__7_), .CO(
        CARRYB_15__6_), .S(SUMB_15__6_) );
  ADDFHX4 S2_8_2 ( .A(ab_8__2_), .B(CARRYB_7__2_), .CI(SUMB_7__3_), .CO(
        CARRYB_8__2_), .S(SUMB_8__2_) );
  ADDFHX4 S2_11_5 ( .A(ab_11__5_), .B(CARRYB_10__5_), .CI(SUMB_10__6_), .CO(
        CARRYB_11__5_), .S(SUMB_11__5_) );
  ADDFHX4 S4_4 ( .A(ab_16__4_), .B(CARRYB_15__4_), .CI(SUMB_15__5_), .CO(
        CARRYB_16__4_), .S(SUMB_16__4_) );
  ADDFHX4 S3_9_6 ( .A(ab_9__6_), .B(CARRYB_8__6_), .CI(ab_8__7_), .CO(
        CARRYB_9__6_), .S(SUMB_9__6_) );
  ADDFHX4 S3_8_6 ( .A(ab_8__6_), .B(CARRYB_7__6_), .CI(ab_7__7_), .CO(
        CARRYB_8__6_), .S(SUMB_8__6_) );
  ADDFHX4 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  ADDFHX4 S2_7_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  ADDFHX4 S2_7_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  ADDFHX4 S2_10_5 ( .A(ab_10__5_), .B(CARRYB_9__5_), .CI(SUMB_9__6_), .CO(
        CARRYB_10__5_), .S(SUMB_10__5_) );
  ADDFHX4 S2_13_4 ( .A(ab_13__4_), .B(CARRYB_12__4_), .CI(SUMB_12__5_), .CO(
        CARRYB_13__4_), .S(SUMB_13__4_) );
  ADDFHX4 S2_15_3 ( .A(ab_15__3_), .B(CARRYB_14__3_), .CI(SUMB_14__4_), .CO(
        CARRYB_15__3_), .S(SUMB_15__3_) );
  ADDFHX4 S2_2_3 ( .A(ab_2__3_), .B(n9), .CI(SUMB_1__4_), .CO(CARRYB_2__3_), 
        .S(SUMB_2__3_) );
  ADDFHX4 S2_7_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  ADDFHX4 S2_8_4 ( .A(ab_8__4_), .B(CARRYB_7__4_), .CI(SUMB_7__5_), .CO(
        CARRYB_8__4_), .S(SUMB_8__4_) );
  ADDFHX4 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  ADDFHX4 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  ADDFHX4 S3_7_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(
        CARRYB_7__6_), .S(SUMB_7__6_) );
  ADDFHX4 S3_12_6 ( .A(ab_12__6_), .B(CARRYB_11__6_), .CI(ab_11__7_), .CO(
        CARRYB_12__6_), .S(SUMB_12__6_) );
  ADDFHX4 S3_11_6 ( .A(ab_11__6_), .B(CARRYB_10__6_), .CI(ab_10__7_), .CO(
        CARRYB_11__6_), .S(SUMB_11__6_) );
  ADDFHX4 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  ADDFHX4 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  ADDFHX4 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  ADDFHX4 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  ADDFHX4 S2_2_4 ( .A(ab_2__4_), .B(n4), .CI(SUMB_1__5_), .CO(CARRYB_2__4_), 
        .S(SUMB_2__4_) );
  ADDFHX4 S2_8_3 ( .A(ab_8__3_), .B(CARRYB_7__3_), .CI(SUMB_7__4_), .CO(
        CARRYB_8__3_), .S(SUMB_8__3_) );
  ADDFHX4 S2_9_3 ( .A(ab_9__3_), .B(CARRYB_8__3_), .CI(SUMB_8__4_), .CO(
        CARRYB_9__3_), .S(SUMB_9__3_) );
  ADDFHX4 S2_13_3 ( .A(ab_13__3_), .B(CARRYB_12__3_), .CI(SUMB_12__4_), .CO(
        CARRYB_13__3_), .S(SUMB_13__3_) );
  ADDFHX4 S3_10_6 ( .A(ab_10__6_), .B(CARRYB_9__6_), .CI(ab_9__7_), .CO(
        CARRYB_10__6_), .S(SUMB_10__6_) );
  ADDFHX4 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  ADDFHX4 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  ADDFHX4 S2_14_1 ( .A(ab_14__1_), .B(CARRYB_13__1_), .CI(SUMB_13__2_), .CO(
        CARRYB_14__1_), .S(SUMB_14__1_) );
  ADDFHX4 S2_15_1 ( .A(ab_15__1_), .B(CARRYB_14__1_), .CI(SUMB_14__2_), .CO(
        CARRYB_15__1_), .S(SUMB_15__1_) );
  ADDFHX4 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  ADDFHX4 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  ADDFHX4 S2_9_4 ( .A(ab_9__4_), .B(CARRYB_8__4_), .CI(SUMB_8__5_), .CO(
        CARRYB_9__4_), .S(SUMB_9__4_) );
  ADDFHX4 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  ADDFHX4 S2_7_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  ADDFHX4 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  ADDFHX4 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  ADDFHX4 S1_9_0 ( .A(ab_9__0_), .B(CARRYB_8__0_), .CI(SUMB_8__1_), .CO(
        CARRYB_9__0_), .S(A1_7_) );
  ADDFHX4 S2_8_5 ( .A(ab_8__5_), .B(CARRYB_7__5_), .CI(SUMB_7__6_), .CO(
        CARRYB_8__5_), .S(SUMB_8__5_) );
  ADDFHX4 S2_9_5 ( .A(ab_9__5_), .B(CARRYB_8__5_), .CI(SUMB_8__6_), .CO(
        CARRYB_9__5_), .S(SUMB_9__5_) );
  ADDFHX4 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  ADDFHX4 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  ADDFHX4 S3_4_6 ( .A(ab_4__6_), .B(ab_3__7_), .CI(CARRYB_3__6_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  ADDFHX4 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  ADDFHX4 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  ADDFHX4 S2_2_1 ( .A(CARRYB_1__1_), .B(ab_2__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  ADDFHX4 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  ADDFHX4 S2_2_5 ( .A(ab_2__5_), .B(n8), .CI(SUMB_1__6_), .CO(CARRYB_2__5_), 
        .S(SUMB_2__5_) );
  ADDFHX4 S2_8_1 ( .A(ab_8__1_), .B(CARRYB_7__1_), .CI(SUMB_7__2_), .CO(
        CARRYB_8__1_), .S(SUMB_8__1_) );
  ADDFHX4 S2_9_1 ( .A(ab_9__1_), .B(CARRYB_8__1_), .CI(SUMB_8__2_), .CO(
        CARRYB_9__1_), .S(SUMB_9__1_) );
  ADDFHX4 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  ADDFHX4 S2_10_2 ( .A(ab_10__2_), .B(CARRYB_9__2_), .CI(SUMB_9__3_), .CO(
        CARRYB_10__2_), .S(SUMB_10__2_) );
  ADDFHX4 S2_11_2 ( .A(ab_11__2_), .B(CARRYB_10__2_), .CI(SUMB_10__3_), .CO(
        CARRYB_11__2_), .S(SUMB_11__2_) );
  ADDFHX4 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  ADDFHX4 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  ADDFHX4 S2_2_2 ( .A(ab_2__2_), .B(n10), .CI(SUMB_1__3_), .CO(CARRYB_2__2_), 
        .S(SUMB_2__2_) );
  ADDFHX4 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  ADDFHX4 S2_7_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  ADDFHX4 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  ADDFHX4 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  ADDFHX4 S2_14_2 ( .A(ab_14__2_), .B(CARRYB_13__2_), .CI(SUMB_13__3_), .CO(
        CARRYB_14__2_), .S(SUMB_14__2_) );
  ADDFHX4 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  ADDFHX2 S3_2_6 ( .A(ab_2__6_), .B(n6), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  ADDFHX4 S4_5 ( .A(ab_16__5_), .B(CARRYB_15__5_), .CI(SUMB_15__6_), .CO(
        CARRYB_16__5_), .S(SUMB_16__5_) );
  ADDFHX2 S2_12_5 ( .A(ab_12__5_), .B(CARRYB_11__5_), .CI(SUMB_11__6_), .CO(
        CARRYB_12__5_), .S(SUMB_12__5_) );
  ADDFHX4 S3_13_6 ( .A(ab_13__6_), .B(CARRYB_12__6_), .CI(ab_12__7_), .CO(
        CARRYB_13__6_), .S(SUMB_13__6_) );
  ADDFHX4 S2_15_4 ( .A(ab_15__4_), .B(SUMB_14__5_), .CI(CARRYB_14__4_), .CO(
        CARRYB_15__4_), .S(SUMB_15__4_) );
  ADDFHX2 S3_14_6 ( .A(ab_14__6_), .B(CARRYB_13__6_), .CI(ab_13__7_), .CO(
        CARRYB_14__6_), .S(SUMB_14__6_) );
  ADDFHX2 S1_10_0 ( .A(ab_10__0_), .B(CARRYB_9__0_), .CI(SUMB_9__1_), .CO(
        CARRYB_10__0_), .S(A1_8_) );
  ADDFHX2 S3_3_6 ( .A(ab_3__6_), .B(ab_2__7_), .CI(CARRYB_2__6_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  ADDFHX2 S2_13_5 ( .A(ab_13__5_), .B(SUMB_12__6_), .CI(CARRYB_12__5_), .CO(
        CARRYB_13__5_), .S(SUMB_13__5_) );
  ADDFHX4 S2_14_5 ( .A(ab_14__5_), .B(SUMB_13__6_), .CI(CARRYB_13__5_), .CO(
        CARRYB_14__5_), .S(SUMB_14__5_) );
  ADDFHX4 S2_14_4 ( .A(ab_14__4_), .B(CARRYB_13__4_), .CI(SUMB_13__5_), .CO(
        CARRYB_14__4_), .S(SUMB_14__4_) );
  AND3X2 U2 ( .A(n15), .B(B[1]), .C(n35), .Y(CARRYB_1__0_) );
  NOR2BX2 U3 ( .AN(n15), .B(n30), .Y(n3) );
  BUFX20 U4 ( .A(A[1]), .Y(n15) );
  AND2X4 U5 ( .A(ab_0__5_), .B(ab_1__4_), .Y(n4) );
  XOR2X2 U6 ( .A(n3), .B(ab_0__2_), .Y(SUMB_1__1_) );
  DLY1X1 U7 ( .A(n22), .Y(n23) );
  NOR2BX2 U8 ( .AN(A[8]), .B(n28), .Y(ab_8__2_) );
  NOR2BX1 U9 ( .AN(A[14]), .B(n31), .Y(ab_14__1_) );
  NOR2BX2 U10 ( .AN(A[7]), .B(n28), .Y(ab_7__2_) );
  NOR2BX1 U11 ( .AN(A[11]), .B(n31), .Y(ab_11__1_) );
  NOR2BX2 U12 ( .AN(A[7]), .B(n30), .Y(ab_7__1_) );
  NOR2BX1 U13 ( .AN(A[9]), .B(n27), .Y(ab_9__3_) );
  NOR2BX1 U14 ( .AN(A[13]), .B(n27), .Y(ab_13__3_) );
  NOR2BX1 U15 ( .AN(A[13]), .B(n25), .Y(ab_13__4_) );
  NOR2BX1 U16 ( .AN(A[9]), .B(n29), .Y(ab_9__2_) );
  NOR2BX2 U17 ( .AN(A[8]), .B(n30), .Y(ab_8__1_) );
  NOR2BX1 U18 ( .AN(A[13]), .B(n31), .Y(ab_13__1_) );
  NOR2BX1 U19 ( .AN(A[13]), .B(n23), .Y(ab_13__5_) );
  NOR2BX1 U20 ( .AN(A[11]), .B(n23), .Y(ab_11__5_) );
  NOR2BX1 U21 ( .AN(A[11]), .B(n29), .Y(ab_11__2_) );
  NOR2BX1 U22 ( .AN(A[9]), .B(n31), .Y(ab_9__1_) );
  NOR2BX1 U23 ( .AN(A[16]), .B(n27), .Y(ab_16__3_) );
  NOR2BXL U24 ( .AN(A[16]), .B(n33), .Y(ab_16__0_) );
  NOR2BX2 U25 ( .AN(A[4]), .B(n26), .Y(ab_4__3_) );
  NOR2BX2 U26 ( .AN(A[5]), .B(n30), .Y(ab_5__1_) );
  NOR2BX2 U27 ( .AN(A[12]), .B(n32), .Y(ab_12__6_) );
  NOR2BX1 U28 ( .AN(A[9]), .B(n25), .Y(ab_9__4_) );
  NOR2BX1 U29 ( .AN(A[10]), .B(n23), .Y(ab_10__5_) );
  NOR2BX2 U30 ( .AN(A[8]), .B(n26), .Y(ab_8__3_) );
  NOR2BX1 U31 ( .AN(A[14]), .B(n27), .Y(ab_14__3_) );
  BUFX3 U32 ( .A(n40), .Y(n29) );
  NOR2BX1 U33 ( .AN(A[14]), .B(n25), .Y(ab_14__4_) );
  NOR2BX1 U34 ( .AN(A[12]), .B(n31), .Y(ab_12__1_) );
  INVX4 U35 ( .A(B[2]), .Y(n40) );
  NOR2BX1 U36 ( .AN(A[14]), .B(n23), .Y(ab_14__5_) );
  NOR2BX2 U37 ( .AN(A[6]), .B(n30), .Y(ab_6__1_) );
  AND2X4 U39 ( .A(ab_0__7_), .B(ab_1__6_), .Y(n6) );
  AND2X4 U40 ( .A(CARRYB_16__1_), .B(SUMB_16__2_), .Y(n7) );
  AND2X4 U41 ( .A(ab_1__5_), .B(ab_0__6_), .Y(n8) );
  AND2X4 U42 ( .A(ab_0__4_), .B(ab_1__3_), .Y(n9) );
  AND2X4 U43 ( .A(ab_1__2_), .B(ab_0__3_), .Y(n10) );
  CLKINVX8 U44 ( .A(B[0]), .Y(n33) );
  NOR2BX2 U45 ( .AN(A[2]), .B(n33), .Y(ab_2__0_) );
  BUFX16 U46 ( .A(A[3]), .Y(n11) );
  NOR2BX1 U47 ( .AN(n15), .B(n42), .Y(ab_1__7_) );
  INVX12 U48 ( .A(A[0]), .Y(n34) );
  INVX4 U49 ( .A(n21), .Y(CARRYB_1__1_) );
  XOR2X4 U50 ( .A(ab_1__2_), .B(ab_0__3_), .Y(SUMB_1__2_) );
  XOR2X4 U51 ( .A(ab_1__3_), .B(ab_0__4_), .Y(SUMB_1__3_) );
  INVX4 U52 ( .A(B[6]), .Y(n36) );
  BUFX20 U53 ( .A(n36), .Y(n32) );
  AND2X4 U54 ( .A(B[6]), .B(n15), .Y(ab_1__6_) );
  XOR2X4 U55 ( .A(ab_1__5_), .B(ab_0__6_), .Y(SUMB_1__5_) );
  BUFX20 U56 ( .A(n41), .Y(n30) );
  CLKINVX8 U57 ( .A(B[1]), .Y(n41) );
  XOR2X4 U58 ( .A(CARRYB_16__4_), .B(SUMB_16__5_), .Y(A1_19_) );
  NOR2BX2 U59 ( .AN(A[6]), .B(n32), .Y(ab_6__6_) );
  XOR2X4 U60 ( .A(ab_1__6_), .B(ab_0__7_), .Y(SUMB_1__6_) );
  NAND2X4 U61 ( .A(n43), .B(ab_0__2_), .Y(n21) );
  DLY1X1 U62 ( .A(n24), .Y(n12) );
  NOR2BX4 U63 ( .AN(n11), .B(n24), .Y(ab_3__4_) );
  NOR2BX4 U64 ( .AN(n11), .B(n30), .Y(ab_3__1_) );
  NOR2BX2 U65 ( .AN(A[4]), .B(n32), .Y(ab_4__6_) );
  NOR2BX4 U66 ( .AN(n11), .B(n28), .Y(ab_3__2_) );
  DLY1X1 U67 ( .A(n24), .Y(n25) );
  NOR2BX2 U68 ( .AN(A[5]), .B(n22), .Y(ab_5__5_) );
  CLKINVX4 U69 ( .A(n37), .Y(n13) );
  AND2X4 U70 ( .A(B[6]), .B(A[0]), .Y(ab_0__6_) );
  INVX3 U71 ( .A(B[3]), .Y(n39) );
  CLKINVX4 U72 ( .A(n38), .Y(n14) );
  NOR2BX4 U73 ( .AN(A[4]), .B(n24), .Y(ab_4__4_) );
  NOR2BX2 U74 ( .AN(A[5]), .B(n24), .Y(ab_5__4_) );
  NOR2BX2 U75 ( .AN(A[5]), .B(n26), .Y(ab_5__3_) );
  INVX8 U76 ( .A(B[5]), .Y(n37) );
  NOR2BX2 U77 ( .AN(A[5]), .B(n32), .Y(ab_5__6_) );
  INVX8 U78 ( .A(B[4]), .Y(n38) );
  NOR2BX4 U79 ( .AN(n14), .B(n34), .Y(ab_0__4_) );
  BUFX20 U80 ( .A(n37), .Y(n22) );
  BUFX20 U81 ( .A(n38), .Y(n24) );
  NOR2BX4 U82 ( .AN(n13), .B(n34), .Y(ab_0__5_) );
  NOR2BX4 U83 ( .AN(n11), .B(n26), .Y(ab_3__3_) );
  NOR2BX4 U84 ( .AN(A[2]), .B(n30), .Y(ab_2__1_) );
  XOR2X4 U85 ( .A(ab_1__4_), .B(ab_0__5_), .Y(SUMB_1__4_) );
  BUFX20 U86 ( .A(n40), .Y(n28) );
  NOR2BX2 U87 ( .AN(n11), .B(n32), .Y(ab_3__6_) );
  NOR2BX4 U88 ( .AN(A[2]), .B(n32), .Y(ab_2__6_) );
  NOR2BX4 U89 ( .AN(A[2]), .B(n28), .Y(ab_2__2_) );
  NOR2BX2 U90 ( .AN(A[4]), .B(n22), .Y(ab_4__5_) );
  INVX20 U91 ( .A(B[7]), .Y(n42) );
  NOR2BX2 U92 ( .AN(A[2]), .B(n42), .Y(ab_2__7_) );
  NOR2BX2 U93 ( .AN(n11), .B(n42), .Y(ab_3__7_) );
  NOR2BX2 U94 ( .AN(A[4]), .B(n42), .Y(ab_4__7_) );
  NOR2BX2 U95 ( .AN(A[6]), .B(n42), .Y(ab_6__7_) );
  NOR2BX2 U96 ( .AN(A[7]), .B(n42), .Y(ab_7__7_) );
  NOR2BX2 U97 ( .AN(A[8]), .B(n42), .Y(ab_8__7_) );
  NOR2BX2 U98 ( .AN(A[9]), .B(n42), .Y(ab_9__7_) );
  NOR2BX2 U99 ( .AN(n11), .B(n22), .Y(ab_3__5_) );
  NOR2BX2 U100 ( .AN(A[5]), .B(n28), .Y(ab_5__2_) );
  NOR2BX2 U101 ( .AN(A[7]), .B(n26), .Y(ab_7__3_) );
  NOR2BX1 U102 ( .AN(A[15]), .B(n25), .Y(ab_15__4_) );
  NOR2BX1 U103 ( .AN(A[7]), .B(n32), .Y(ab_7__6_) );
  NOR2BX2 U104 ( .AN(n11), .B(n33), .Y(ab_3__0_) );
  NOR2BX2 U105 ( .AN(A[4]), .B(n33), .Y(ab_4__0_) );
  NOR2BX2 U106 ( .AN(A[5]), .B(n33), .Y(ab_5__0_) );
  NOR2BX2 U107 ( .AN(A[6]), .B(n33), .Y(ab_6__0_) );
  NOR2BX2 U108 ( .AN(A[7]), .B(n33), .Y(ab_7__0_) );
  NOR2BX2 U109 ( .AN(A[8]), .B(n33), .Y(ab_8__0_) );
  NOR2BX1 U110 ( .AN(A[0]), .B(n33), .Y(n35) );
  NOR2BX2 U111 ( .AN(A[4]), .B(n28), .Y(ab_4__2_) );
  NOR2BX2 U112 ( .AN(A[4]), .B(n30), .Y(ab_4__1_) );
  NOR2BX4 U113 ( .AN(B[7]), .B(n34), .Y(ab_0__7_) );
  NOR2BX1 U114 ( .AN(A[7]), .B(n12), .Y(ab_7__4_) );
  NOR2BX4 U115 ( .AN(A[2]), .B(n26), .Y(ab_2__3_) );
  NOR2BXL U116 ( .AN(A[12]), .B(n33), .Y(ab_12__0_) );
  NOR2BXL U117 ( .AN(A[11]), .B(n33), .Y(ab_11__0_) );
  NOR2BXL U118 ( .AN(A[10]), .B(n33), .Y(ab_10__0_) );
  NOR2BXL U119 ( .AN(A[9]), .B(n33), .Y(ab_9__0_) );
  NOR2BX4 U120 ( .AN(A[2]), .B(n24), .Y(ab_2__4_) );
  NOR2BX4 U121 ( .AN(n15), .B(n30), .Y(n43) );
  NOR2BX4 U122 ( .AN(n15), .B(n24), .Y(ab_1__4_) );
  NOR2BX4 U123 ( .AN(n15), .B(n28), .Y(ab_1__2_) );
  NOR2BX4 U124 ( .AN(A[2]), .B(n22), .Y(ab_2__5_) );
  NOR2BX4 U125 ( .AN(n15), .B(n26), .Y(ab_1__3_) );
  AND2X2 U126 ( .A(CARRYB_16__2_), .B(SUMB_16__3_), .Y(n18) );
  NOR2BX1 U127 ( .AN(A[13]), .B(n33), .Y(ab_13__0_) );
  NOR2BX1 U128 ( .AN(A[11]), .B(n42), .Y(ab_11__7_) );
  NOR2BX1 U129 ( .AN(A[10]), .B(n42), .Y(ab_10__7_) );
  NOR2BX1 U130 ( .AN(A[12]), .B(n42), .Y(ab_12__7_) );
  NOR2BX1 U131 ( .AN(A[6]), .B(n22), .Y(ab_6__5_) );
  NOR2BX1 U132 ( .AN(A[6]), .B(n28), .Y(ab_6__2_) );
  NOR2BX1 U133 ( .AN(A[8]), .B(n12), .Y(ab_8__4_) );
  NOR2BX1 U134 ( .AN(A[6]), .B(n24), .Y(ab_6__4_) );
  NOR2BX1 U135 ( .AN(A[14]), .B(n33), .Y(ab_14__0_) );
  NOR2BX1 U136 ( .AN(A[6]), .B(n26), .Y(ab_6__3_) );
  NOR2BX1 U137 ( .AN(A[10]), .B(n31), .Y(ab_10__1_) );
  AND2X4 U138 ( .A(CARRYB_16__0_), .B(SUMB_16__1_), .Y(n16) );
  AND2X1 U139 ( .A(CARRYB_16__4_), .B(SUMB_16__5_), .Y(n19) );
  NOR2BX1 U140 ( .AN(A[9]), .B(n23), .Y(ab_9__5_) );
  NOR2BXL U141 ( .AN(A[8]), .B(n22), .Y(ab_8__5_) );
  NOR2BX1 U142 ( .AN(A[12]), .B(n23), .Y(ab_12__5_) );
  NOR2BX1 U143 ( .AN(A[13]), .B(n29), .Y(ab_13__2_) );
  NOR2BX1 U144 ( .AN(A[12]), .B(n27), .Y(ab_12__3_) );
  NOR2BX1 U145 ( .AN(A[12]), .B(n25), .Y(ab_12__4_) );
  NOR2BX1 U146 ( .AN(A[11]), .B(n25), .Y(ab_11__4_) );
  NOR2BX1 U147 ( .AN(A[10]), .B(n25), .Y(ab_10__4_) );
  NOR2BX1 U148 ( .AN(A[11]), .B(n27), .Y(ab_11__3_) );
  NOR2BX1 U149 ( .AN(A[12]), .B(n29), .Y(ab_12__2_) );
  NOR2BX1 U150 ( .AN(A[10]), .B(n27), .Y(ab_10__3_) );
  NOR2BX4 U151 ( .AN(n15), .B(n22), .Y(ab_1__5_) );
  BUFX8 U152 ( .A(n39), .Y(n26) );
  NOR2BX1 U153 ( .AN(A[13]), .B(n42), .Y(ab_13__7_) );
  NOR2BXL U154 ( .AN(A[14]), .B(n32), .Y(ab_14__6_) );
  NOR2BXL U155 ( .AN(A[10]), .B(n32), .Y(ab_10__6_) );
  NOR2BXL U156 ( .AN(A[8]), .B(n32), .Y(ab_8__6_) );
  NOR2BX2 U157 ( .AN(A[16]), .B(n29), .Y(ab_16__2_) );
  NOR2BXL U158 ( .AN(A[9]), .B(n32), .Y(ab_9__6_) );
  NOR2BXL U159 ( .AN(A[13]), .B(n32), .Y(ab_13__6_) );
  NOR2BX1 U160 ( .AN(A[14]), .B(n42), .Y(ab_14__7_) );
  NOR2BXL U161 ( .AN(A[15]), .B(n32), .Y(ab_15__6_) );
  NOR2BXL U162 ( .AN(A[11]), .B(n32), .Y(ab_11__6_) );
  NOR2BXL U163 ( .AN(A[16]), .B(n32), .Y(ab_16__6_) );
  DLY1X1 U164 ( .A(n41), .Y(n31) );
  CLKBUFXL U165 ( .A(n39), .Y(n27) );
  AND2X2 U166 ( .A(CARRYB_16__3_), .B(SUMB_16__4_), .Y(n17) );
  NOR2BX1 U167 ( .AN(A[7]), .B(n22), .Y(ab_7__5_) );
  NOR2BX1 U168 ( .AN(A[14]), .B(n29), .Y(ab_14__2_) );
  AND2X2 U169 ( .A(CARRYB_16__5_), .B(SUMB_16__6_), .Y(n20) );
  NOR2BX1 U170 ( .AN(A[16]), .B(n25), .Y(ab_16__4_) );
  NOR2BX1 U171 ( .AN(A[16]), .B(n23), .Y(ab_16__5_) );
  NOR2BX1 U172 ( .AN(A[15]), .B(n27), .Y(ab_15__3_) );
  NOR2BX1 U173 ( .AN(A[5]), .B(n42), .Y(ab_5__7_) );
  NOR2BX1 U174 ( .AN(A[16]), .B(n31), .Y(ab_16__1_) );
  NOR2BXL U175 ( .AN(A[15]), .B(n23), .Y(ab_15__5_) );
  NOR2BXL U176 ( .AN(A[15]), .B(n33), .Y(ab_15__0_) );
  NOR2BX1 U177 ( .AN(A[15]), .B(n29), .Y(ab_15__2_) );
  NOR2BX1 U178 ( .AN(A[15]), .B(n31), .Y(ab_15__1_) );
  NOR2BXL U179 ( .AN(A[15]), .B(n42), .Y(ab_15__7_) );
  NOR2BXL U180 ( .AN(A[16]), .B(n42), .Y(ab_16__7_) );
  XOR2X4 U181 ( .A(CARRYB_16__3_), .B(SUMB_16__4_), .Y(A1_18_) );
  XOR2X4 U182 ( .A(CARRYB_16__5_), .B(SUMB_16__6_), .Y(A1_20_) );
  XOR2X4 U183 ( .A(CARRYB_16__6_), .B(ab_16__7_), .Y(A1_21_) );
  XOR2X4 U184 ( .A(SUMB_16__2_), .B(CARRYB_16__1_), .Y(A1_16_) );
  XOR2X4 U185 ( .A(SUMB_16__1_), .B(CARRYB_16__0_), .Y(A1_15_) );
  XOR2X4 U186 ( .A(SUMB_16__3_), .B(CARRYB_16__2_), .Y(A1_17_) );
  NOR2BX4 U187 ( .AN(B[3]), .B(n34), .Y(ab_0__3_) );
  NOR2BX4 U188 ( .AN(B[2]), .B(n34), .Y(ab_0__2_) );
  NOR2BX4 U189 ( .AN(A[10]), .B(n29), .Y(ab_10__2_) );
endmodule


module multi16_8 ( in_17bit, in_8bit, out );
  input [16:0] in_17bit;
  input [7:0] in_8bit;
  output [16:0] out;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107;
  wire   [16:1] in_17bit_b;
  wire   [7:1] in_8bit_b;
  wire   [23:8] mul;

  multi16_8_DW02_mult_0 mult_55 ( .A({in_17bit_b[16:3], n15, in_17bit_b[1], 
        in_17bit[0]}), .B({in_8bit_b, n10}), .PRODUCT_23_(mul[23]), 
        .PRODUCT_22_(mul[22]), .PRODUCT_21_(mul[21]), .PRODUCT_20_(mul[20]), 
        .PRODUCT_19_(mul[19]), .PRODUCT_18_(mul[18]), .PRODUCT_17_(mul[17]), 
        .PRODUCT_16_(mul[16]), .PRODUCT_15_(mul[15]), .PRODUCT_14_(mul[14]), 
        .PRODUCT_13_(mul[13]), .PRODUCT_12_(mul[12]), .PRODUCT_11_(mul[11]), 
        .PRODUCT_10_(mul[10]), .PRODUCT_9_(mul[9]), .PRODUCT_8_(mul[8]), 
        .PRODUCT_7_(out[0]) );
  BUFX20 U2 ( .A(in_8bit[0]), .Y(n42) );
  AOI21X2 U3 ( .A0(n106), .A1(n12), .B0(n104), .Y(n107) );
  NOR2X1 U4 ( .A(mul[22]), .B(mul[21]), .Y(n106) );
  XOR2X4 U5 ( .A(n46), .B(n1), .Y(in_8bit_b[5]) );
  CLKINVX20 U6 ( .A(n47), .Y(n1) );
  XOR2X4 U7 ( .A(n50), .B(n2), .Y(in_8bit_b[6]) );
  CLKINVX20 U8 ( .A(in_8bit[6]), .Y(n2) );
  BUFX8 U9 ( .A(mul[20]), .Y(n3) );
  INVX20 U10 ( .A(n104), .Y(n101) );
  XNOR2X4 U11 ( .A(n97), .B(n3), .Y(out[13]) );
  BUFX12 U12 ( .A(n49), .Y(n9) );
  XNOR2X4 U13 ( .A(in_8bit[1]), .B(n28), .Y(in_8bit_b[1]) );
  CLKBUFX8 U14 ( .A(n42), .Y(n10) );
  NOR2X2 U15 ( .A(n35), .B(n40), .Y(n76) );
  CLKINVX3 U16 ( .A(n55), .Y(n57) );
  INVX1 U17 ( .A(n91), .Y(n8) );
  CLKINVX3 U18 ( .A(n95), .Y(n99) );
  AND2X4 U19 ( .A(n48), .B(n47), .Y(n4) );
  AOI21X2 U20 ( .A0(in_17bit[16]), .A1(in_17bit[0]), .B0(in_17bit[1]), .Y(n53)
         );
  INVX8 U21 ( .A(n19), .Y(out[8]) );
  XOR2X4 U22 ( .A(mul[15]), .B(n20), .Y(n19) );
  NOR2X4 U23 ( .A(n9), .B(n51), .Y(n25) );
  NAND2BX4 U24 ( .AN(in_8bit[1]), .B(n41), .Y(n5) );
  AND3X4 U25 ( .A(in_17bit[0]), .B(in_17bit[16]), .C(in_17bit[1]), .Y(n6) );
  NOR2X4 U26 ( .A(n53), .B(n6), .Y(in_17bit_b[1]) );
  INVXL U27 ( .A(n78), .Y(n7) );
  INVX3 U28 ( .A(in_17bit[16]), .Y(n78) );
  INVX8 U29 ( .A(n102), .Y(n105) );
  BUFX20 U30 ( .A(n78), .Y(n40) );
  NAND2X4 U31 ( .A(n93), .B(n101), .Y(n92) );
  INVX4 U32 ( .A(in_8bit[5]), .Y(n47) );
  NOR3X4 U33 ( .A(in_8bit[6]), .B(n51), .C(n52), .Y(in_8bit_b[7]) );
  CLKINVX8 U34 ( .A(mul[18]), .Y(n98) );
  BUFX20 U35 ( .A(in_17bit_b[2]), .Y(n15) );
  NAND2BX4 U36 ( .AN(mul[16]), .B(n8), .Y(n93) );
  XNOR2X4 U37 ( .A(mul[13]), .B(n85), .Y(out[6]) );
  NAND2X4 U38 ( .A(n86), .B(n101), .Y(n85) );
  NAND2BX4 U39 ( .AN(mul[18]), .B(n99), .Y(n96) );
  OAI2BB1X4 U40 ( .A0N(n98), .A1N(n99), .B0(n101), .Y(n94) );
  NAND2BX2 U41 ( .AN(in_17bit[3]), .B(n39), .Y(n55) );
  NAND2X4 U42 ( .A(n54), .B(in_17bit[16]), .Y(n26) );
  NAND2BX4 U43 ( .AN(n51), .B(n52), .Y(n50) );
  XOR2X4 U44 ( .A(n43), .B(n41), .Y(in_8bit_b[2]) );
  NOR2X4 U45 ( .A(n105), .B(n104), .Y(n100) );
  NOR2X4 U46 ( .A(n57), .B(n40), .Y(n14) );
  INVXL U47 ( .A(n105), .Y(n11) );
  INVX2 U48 ( .A(n11), .Y(n12) );
  NAND2X2 U49 ( .A(n81), .B(n101), .Y(n21) );
  XOR2X2 U50 ( .A(mul[23]), .B(n107), .Y(out[16]) );
  XOR2X4 U51 ( .A(n25), .B(in_8bit[4]), .Y(in_8bit_b[4]) );
  AOI21X4 U52 ( .A0(n9), .A1(n48), .B0(n51), .Y(n46) );
  NAND2X4 U53 ( .A(n4), .B(n9), .Y(n52) );
  NAND2X4 U54 ( .A(n10), .B(in_8bit[7]), .Y(n28) );
  XNOR2X2 U55 ( .A(n44), .B(in_8bit[3]), .Y(in_8bit_b[3]) );
  XNOR2X4 U56 ( .A(n26), .B(in_17bit[2]), .Y(in_17bit_b[2]) );
  OR2X4 U57 ( .A(n39), .B(n40), .Y(n24) );
  XOR2X4 U58 ( .A(n14), .B(n13), .Y(in_17bit_b[4]) );
  CLKINVX20 U59 ( .A(n56), .Y(n13) );
  AND2X2 U60 ( .A(n57), .B(n56), .Y(n34) );
  AND2X4 U61 ( .A(n33), .B(n61), .Y(n32) );
  AND2X2 U62 ( .A(n34), .B(n59), .Y(n33) );
  XNOR2X4 U63 ( .A(n27), .B(in_17bit[15]), .Y(in_17bit_b[15]) );
  XNOR2X2 U64 ( .A(mul[10]), .B(n21), .Y(out[3]) );
  OAI21X2 U65 ( .A0(mul[21]), .A1(n102), .B0(n101), .Y(n103) );
  XNOR2X2 U66 ( .A(mul[9]), .B(n16), .Y(out[2]) );
  NAND4BBX4 U67 ( .AN(mul[20]), .BN(mul[19]), .C(n99), .D(n98), .Y(n102) );
  OR2X4 U68 ( .A(mul[17]), .B(n93), .Y(n95) );
  NAND2BX4 U69 ( .AN(in_8bit[1]), .B(n41), .Y(n45) );
  CLKINVX8 U70 ( .A(in_8bit[2]), .Y(n41) );
  OR2X4 U71 ( .A(mul[10]), .B(n81), .Y(n83) );
  XNOR2X2 U72 ( .A(mul[11]), .B(n82), .Y(out[4]) );
  NOR2X4 U73 ( .A(in_17bit[2]), .B(n54), .Y(n39) );
  OAI21X4 U74 ( .A0(n42), .A1(n5), .B0(in_8bit[7]), .Y(n44) );
  XOR2X4 U75 ( .A(mul[12]), .B(n17), .Y(out[5]) );
  NAND2X2 U76 ( .A(n83), .B(n101), .Y(n82) );
  AND2X2 U77 ( .A(n38), .B(n71), .Y(n37) );
  NAND2X2 U78 ( .A(n88), .B(n101), .Y(n20) );
  OR2X4 U79 ( .A(in_17bit[1]), .B(in_17bit[0]), .Y(n54) );
  OR2X2 U80 ( .A(mul[14]), .B(n87), .Y(n88) );
  OR2X4 U81 ( .A(mul[13]), .B(n86), .Y(n87) );
  OR2X4 U82 ( .A(mul[9]), .B(n80), .Y(n81) );
  OR2X4 U83 ( .A(mul[8]), .B(out[0]), .Y(n80) );
  OR2X4 U84 ( .A(mul[12]), .B(n84), .Y(n86) );
  OR2X4 U85 ( .A(mul[11]), .B(n83), .Y(n84) );
  NAND2XL U86 ( .A(n80), .B(n101), .Y(n16) );
  AND2X2 U87 ( .A(n84), .B(n101), .Y(n17) );
  XNOR2X1 U88 ( .A(mul[8]), .B(n18), .Y(out[1]) );
  NAND2XL U89 ( .A(out[0]), .B(n101), .Y(n18) );
  XNOR2X4 U90 ( .A(mul[18]), .B(n22), .Y(out[11]) );
  NAND2X4 U91 ( .A(n95), .B(n101), .Y(n22) );
  XNOR2X4 U92 ( .A(mul[14]), .B(n23), .Y(out[7]) );
  NAND2X4 U93 ( .A(n87), .B(n101), .Y(n23) );
  AND2X4 U94 ( .A(n37), .B(n73), .Y(n36) );
  AND2X4 U95 ( .A(n36), .B(n75), .Y(n35) );
  XNOR2X4 U96 ( .A(in_17bit[3]), .B(n24), .Y(in_17bit_b[3]) );
  NAND2XL U97 ( .A(n79), .B(n7), .Y(n27) );
  XNOR2X4 U98 ( .A(n103), .B(mul[22]), .Y(out[15]) );
  AND2X2 U99 ( .A(n30), .B(n67), .Y(n29) );
  AND2X2 U100 ( .A(n31), .B(n65), .Y(n30) );
  AND2X2 U101 ( .A(n32), .B(n63), .Y(n31) );
  AND2X2 U102 ( .A(n29), .B(n69), .Y(n38) );
  NAND2XL U103 ( .A(n35), .B(n77), .Y(n79) );
  XNOR2X1 U104 ( .A(in_17bit[16]), .B(in_8bit[7]), .Y(n104) );
  INVX1 U105 ( .A(in_8bit[4]), .Y(n48) );
  INVX1 U106 ( .A(in_8bit[7]), .Y(n51) );
  OAI21X4 U107 ( .A0(n96), .A1(mul[19]), .B0(n101), .Y(n97) );
  OAI21X2 U108 ( .A0(in_8bit[1]), .A1(n42), .B0(in_8bit[7]), .Y(n43) );
  NOR3X4 U109 ( .A(n42), .B(in_8bit[3]), .C(n45), .Y(n49) );
  CLKINVX3 U110 ( .A(in_17bit[4]), .Y(n56) );
  NOR2X4 U111 ( .A(n34), .B(n40), .Y(n58) );
  CLKINVX3 U112 ( .A(in_17bit[5]), .Y(n59) );
  XNOR2X4 U113 ( .A(n58), .B(n59), .Y(in_17bit_b[5]) );
  NOR2X4 U114 ( .A(n33), .B(n40), .Y(n60) );
  CLKINVX3 U115 ( .A(in_17bit[6]), .Y(n61) );
  XNOR2X4 U116 ( .A(n60), .B(n61), .Y(in_17bit_b[6]) );
  NOR2X4 U117 ( .A(n32), .B(n40), .Y(n62) );
  CLKINVX3 U118 ( .A(in_17bit[7]), .Y(n63) );
  XNOR2X4 U119 ( .A(n62), .B(n63), .Y(in_17bit_b[7]) );
  NOR2X4 U120 ( .A(n31), .B(n40), .Y(n64) );
  CLKINVX3 U121 ( .A(in_17bit[8]), .Y(n65) );
  XNOR2X4 U122 ( .A(n64), .B(n65), .Y(in_17bit_b[8]) );
  NOR2X4 U123 ( .A(n30), .B(n40), .Y(n66) );
  CLKINVX3 U124 ( .A(in_17bit[9]), .Y(n67) );
  XNOR2X4 U125 ( .A(n66), .B(n67), .Y(in_17bit_b[9]) );
  NOR2X4 U126 ( .A(n29), .B(n40), .Y(n68) );
  CLKINVX3 U127 ( .A(in_17bit[10]), .Y(n69) );
  XNOR2X4 U128 ( .A(n68), .B(n69), .Y(in_17bit_b[10]) );
  NOR2X4 U129 ( .A(n38), .B(n40), .Y(n70) );
  CLKINVX3 U130 ( .A(in_17bit[11]), .Y(n71) );
  XNOR2X4 U131 ( .A(n70), .B(n71), .Y(in_17bit_b[11]) );
  NOR2X4 U132 ( .A(n37), .B(n40), .Y(n72) );
  CLKINVX3 U133 ( .A(in_17bit[12]), .Y(n73) );
  XNOR2X4 U134 ( .A(n72), .B(n73), .Y(in_17bit_b[12]) );
  NOR2X4 U135 ( .A(n36), .B(n40), .Y(n74) );
  CLKINVX3 U136 ( .A(in_17bit[13]), .Y(n75) );
  XNOR2X4 U137 ( .A(n74), .B(n75), .Y(in_17bit_b[13]) );
  CLKINVX3 U138 ( .A(in_17bit[14]), .Y(n77) );
  XNOR2X4 U139 ( .A(n76), .B(n77), .Y(in_17bit_b[14]) );
  NOR3X4 U140 ( .A(in_17bit[15]), .B(n79), .C(n40), .Y(in_17bit_b[16]) );
  CLKINVX3 U141 ( .A(n88), .Y(n89) );
  NAND2BX4 U142 ( .AN(mul[15]), .B(n89), .Y(n91) );
  NAND2X4 U143 ( .A(n91), .B(n101), .Y(n90) );
  XNOR2X4 U144 ( .A(mul[16]), .B(n90), .Y(out[9]) );
  XNOR2X4 U145 ( .A(mul[17]), .B(n92), .Y(out[10]) );
  XNOR2X4 U146 ( .A(mul[19]), .B(n94), .Y(out[12]) );
  XOR2X4 U147 ( .A(n100), .B(mul[21]), .Y(out[14]) );
endmodule


module multi16_7_DW01_add_5 ( A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, 
        A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, 
        B_20_, B_19_, B_18_, B_17_, B_16_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, 
        SUM_17_, SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, 
        SUM_9_, SUM_8_, SUM_7_, SUM_6_, SUM_5_ );
  input A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_,
         A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, B_20_, B_19_,
         B_18_, B_17_, B_16_;
  output SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, SUM_15_,
         SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, SUM_7_,
         SUM_6_, SUM_5_;
  wire   n1, n2, n3, n4, n5, n6, n7, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43;

  BUFX4 U2 ( .A(n33), .Y(n3) );
  XOR2X4 U3 ( .A(n1), .B(n2), .Y(SUM_18_) );
  NAND2X2 U4 ( .A(n3), .B(n40), .Y(n1) );
  AND2X4 U5 ( .A(n41), .B(n28), .Y(n2) );
  NOR2X2 U6 ( .A(n34), .B(n4), .Y(n29) );
  OR2X2 U7 ( .A(A_17_), .B(B_17_), .Y(n26) );
  AOI21X2 U8 ( .A0(n29), .A1(n30), .B0(n31), .Y(n24) );
  BUFX12 U9 ( .A(A_10_), .Y(SUM_10_) );
  INVX2 U10 ( .A(n32), .Y(n5) );
  NAND2XL U11 ( .A(n32), .B(n33), .Y(n30) );
  NOR2X4 U12 ( .A(A_17_), .B(B_17_), .Y(n4) );
  NAND2BX4 U13 ( .AN(n32), .B(n26), .Y(n40) );
  BUFX12 U14 ( .A(A_14_), .Y(SUM_14_) );
  XOR2X4 U15 ( .A(n42), .B(n5), .Y(SUM_17_) );
  BUFX12 U16 ( .A(A_15_), .Y(SUM_15_) );
  NAND2X4 U17 ( .A(n37), .B(n38), .Y(n35) );
  AOI2BB1X4 U18 ( .A0N(n34), .A1N(n3), .B0(n31), .Y(n37) );
  NAND2X4 U19 ( .A(n39), .B(n28), .Y(n38) );
  CLKINVX4 U20 ( .A(n41), .Y(n31) );
  BUFX12 U21 ( .A(A_12_), .Y(SUM_12_) );
  XNOR3X4 U22 ( .A(B_21_), .B(A_21_), .C(n6), .Y(SUM_21_) );
  NAND2X2 U23 ( .A(B_18_), .B(A_18_), .Y(n41) );
  NAND2X4 U24 ( .A(A_17_), .B(B_17_), .Y(n33) );
  INVX2 U25 ( .A(n40), .Y(n39) );
  INVX8 U26 ( .A(n43), .Y(SUM_16_) );
  NAND2X4 U27 ( .A(B_19_), .B(A_19_), .Y(n25) );
  NOR2X4 U28 ( .A(A_19_), .B(B_19_), .Y(n7) );
  INVX4 U29 ( .A(n28), .Y(n34) );
  NAND2X2 U30 ( .A(B_20_), .B(A_20_), .Y(n19) );
  AND2X4 U31 ( .A(n19), .B(n22), .Y(n23) );
  AND2X2 U32 ( .A(n19), .B(n20), .Y(n6) );
  NOR2BX2 U33 ( .AN(n25), .B(n7), .Y(n36) );
  OR2X4 U34 ( .A(A_18_), .B(B_18_), .Y(n28) );
  OR2X4 U35 ( .A(A_20_), .B(B_20_), .Y(n22) );
  NAND2XL U36 ( .A(n21), .B(n22), .Y(n20) );
  BUFX8 U37 ( .A(A_5_), .Y(SUM_5_) );
  BUFX4 U38 ( .A(A_9_), .Y(SUM_9_) );
  BUFX8 U39 ( .A(A_11_), .Y(SUM_11_) );
  BUFX4 U40 ( .A(A_6_), .Y(SUM_6_) );
  BUFX4 U41 ( .A(A_7_), .Y(SUM_7_) );
  BUFX4 U42 ( .A(A_8_), .Y(SUM_8_) );
  BUFX8 U43 ( .A(A_13_), .Y(SUM_13_) );
  XOR2X4 U44 ( .A(n21), .B(n23), .Y(SUM_20_) );
  OAI21X4 U45 ( .A0(n24), .A1(n7), .B0(n25), .Y(n21) );
  XOR2X4 U46 ( .A(n35), .B(n36), .Y(SUM_19_) );
  NOR2BX4 U47 ( .AN(n33), .B(n4), .Y(n42) );
  NAND2X4 U48 ( .A(n32), .B(n27), .Y(n43) );
  OR2X4 U49 ( .A(A_16_), .B(B_16_), .Y(n27) );
  NAND2X4 U50 ( .A(B_16_), .B(A_16_), .Y(n32) );
endmodule


module multi16_7_DW02_mult_0 ( A, B, PRODUCT_23_, PRODUCT_22_, PRODUCT_21_, 
        PRODUCT_20_, PRODUCT_19_, PRODUCT_18_, PRODUCT_17_, PRODUCT_16_, 
        PRODUCT_15_, PRODUCT_14_, PRODUCT_13_, PRODUCT_12_, PRODUCT_11_, 
        PRODUCT_10_, PRODUCT_9_, PRODUCT_8_, PRODUCT_7_ );
  input [16:0] A;
  input [7:0] B;
  output PRODUCT_23_, PRODUCT_22_, PRODUCT_21_, PRODUCT_20_, PRODUCT_19_,
         PRODUCT_18_, PRODUCT_17_, PRODUCT_16_, PRODUCT_15_, PRODUCT_14_,
         PRODUCT_13_, PRODUCT_12_, PRODUCT_11_, PRODUCT_10_, PRODUCT_9_,
         PRODUCT_8_, PRODUCT_7_;
  wire   ab_16__7_, ab_16__6_, ab_16__5_, ab_16__4_, ab_16__3_, ab_16__2_,
         ab_16__1_, ab_16__0_, ab_15__7_, ab_15__6_, ab_15__5_, ab_15__4_,
         ab_15__3_, ab_15__2_, ab_15__1_, ab_15__0_, ab_14__7_, ab_14__6_,
         ab_14__5_, ab_14__4_, ab_14__3_, ab_14__2_, ab_14__1_, ab_14__0_,
         ab_13__7_, ab_13__6_, ab_13__5_, ab_13__4_, ab_13__3_, ab_13__2_,
         ab_13__1_, ab_13__0_, ab_12__7_, ab_12__6_, ab_12__5_, ab_12__4_,
         ab_12__3_, ab_12__2_, ab_12__1_, ab_12__0_, ab_11__7_, ab_11__6_,
         ab_11__5_, ab_11__4_, ab_11__3_, ab_11__2_, ab_11__1_, ab_11__0_,
         ab_10__7_, ab_10__6_, ab_10__5_, ab_10__4_, ab_10__3_, ab_10__2_,
         ab_10__1_, ab_10__0_, ab_9__7_, ab_9__6_, ab_9__5_, ab_9__4_,
         ab_9__3_, ab_9__2_, ab_9__1_, ab_9__0_, ab_8__7_, ab_8__6_, ab_8__5_,
         ab_8__4_, ab_8__3_, ab_8__2_, ab_8__1_, ab_8__0_, ab_7__7_, ab_7__6_,
         ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_, ab_7__0_, ab_6__7_,
         ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_, ab_6__1_, ab_6__0_,
         ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_, ab_5__2_, ab_5__1_,
         ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_, ab_4__3_, ab_4__2_,
         ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_, ab_3__4_, ab_3__3_,
         ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_, ab_2__5_, ab_2__4_,
         ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_, ab_1__6_, ab_1__5_,
         ab_1__4_, ab_1__3_, ab_1__2_, ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_,
         ab_0__3_, ab_0__2_, CARRYB_16__6_, CARRYB_16__5_, CARRYB_16__4_,
         CARRYB_16__3_, CARRYB_16__2_, CARRYB_16__1_, CARRYB_16__0_,
         CARRYB_15__6_, CARRYB_15__5_, CARRYB_15__4_, CARRYB_15__3_,
         CARRYB_15__2_, CARRYB_15__1_, CARRYB_15__0_, CARRYB_14__6_,
         CARRYB_14__5_, CARRYB_14__4_, CARRYB_14__3_, CARRYB_14__2_,
         CARRYB_14__1_, CARRYB_14__0_, CARRYB_13__6_, CARRYB_13__5_,
         CARRYB_13__4_, CARRYB_13__3_, CARRYB_13__2_, CARRYB_13__1_,
         CARRYB_13__0_, CARRYB_12__6_, CARRYB_12__5_, CARRYB_12__4_,
         CARRYB_12__3_, CARRYB_12__2_, CARRYB_12__1_, CARRYB_12__0_,
         CARRYB_11__6_, CARRYB_11__5_, CARRYB_11__4_, CARRYB_11__3_,
         CARRYB_11__2_, CARRYB_11__1_, CARRYB_11__0_, CARRYB_10__6_,
         CARRYB_10__5_, CARRYB_10__4_, CARRYB_10__3_, CARRYB_10__2_,
         CARRYB_10__1_, CARRYB_10__0_, CARRYB_9__6_, CARRYB_9__5_,
         CARRYB_9__4_, CARRYB_9__3_, CARRYB_9__2_, CARRYB_9__1_, CARRYB_9__0_,
         CARRYB_8__6_, CARRYB_8__5_, CARRYB_8__4_, CARRYB_8__3_, CARRYB_8__2_,
         CARRYB_8__1_, CARRYB_8__0_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_,
         CARRYB_7__3_, CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_,
         CARRYB_6__5_, CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_,
         CARRYB_6__0_, CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_,
         CARRYB_5__2_, CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_,
         CARRYB_4__4_, CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_,
         CARRYB_3__6_, CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_,
         CARRYB_3__1_, CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_,
         CARRYB_2__3_, CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__3_,
         CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_16__6_, SUMB_16__5_,
         SUMB_16__4_, SUMB_16__3_, SUMB_16__2_, SUMB_16__1_, SUMB_16__0_,
         SUMB_15__6_, SUMB_15__5_, SUMB_15__4_, SUMB_15__3_, SUMB_15__2_,
         SUMB_15__1_, SUMB_14__6_, SUMB_14__5_, SUMB_14__4_, SUMB_14__3_,
         SUMB_14__2_, SUMB_14__1_, SUMB_13__6_, SUMB_13__5_, SUMB_13__4_,
         SUMB_13__3_, SUMB_13__2_, SUMB_13__1_, SUMB_12__6_, SUMB_12__5_,
         SUMB_12__4_, SUMB_12__3_, SUMB_12__2_, SUMB_12__1_, SUMB_11__6_,
         SUMB_11__5_, SUMB_11__4_, SUMB_11__3_, SUMB_11__2_, SUMB_11__1_,
         SUMB_10__6_, SUMB_10__5_, SUMB_10__4_, SUMB_10__3_, SUMB_10__2_,
         SUMB_10__1_, SUMB_9__6_, SUMB_9__5_, SUMB_9__4_, SUMB_9__3_,
         SUMB_9__2_, SUMB_9__1_, SUMB_8__6_, SUMB_8__5_, SUMB_8__4_,
         SUMB_8__3_, SUMB_8__2_, SUMB_8__1_, SUMB_7__6_, SUMB_7__5_,
         SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_, SUMB_6__6_,
         SUMB_6__5_, SUMB_6__4_, SUMB_6__3_, SUMB_6__2_, SUMB_6__1_,
         SUMB_5__6_, SUMB_5__5_, SUMB_5__4_, SUMB_5__3_, SUMB_5__2_,
         SUMB_5__1_, SUMB_4__6_, SUMB_4__5_, SUMB_4__4_, SUMB_4__3_,
         SUMB_4__2_, SUMB_4__1_, SUMB_3__6_, SUMB_3__5_, SUMB_3__4_,
         SUMB_3__3_, SUMB_3__2_, SUMB_3__1_, SUMB_2__6_, SUMB_2__5_,
         SUMB_2__4_, SUMB_2__3_, SUMB_2__2_, SUMB_2__1_, SUMB_1__6_,
         SUMB_1__5_, SUMB_1__4_, SUMB_1__3_, SUMB_1__2_, SUMB_1__1_, PROD1_7_,
         A1_21_, A1_20_, A1_19_, A1_18_, A1_17_, A1_16_, A1_15_, A1_13_,
         A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, A1_4_, A1_3_,
         A1_2_, A1_1_, A1_0_, n3, n4, n5, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51;

  ADDFHX2 S5_6 ( .A(ab_16__6_), .B(CARRYB_15__6_), .CI(ab_15__7_), .CO(
        CARRYB_16__6_), .S(SUMB_16__6_) );
  multi16_7_DW01_add_5 FS_1 ( .A_21_(A1_21_), .A_20_(A1_20_), .A_19_(A1_19_), 
        .A_18_(A1_18_), .A_17_(A1_17_), .A_16_(A1_16_), .A_15_(A1_15_), 
        .A_14_(SUMB_16__0_), .A_13_(A1_13_), .A_12_(A1_12_), .A_11_(A1_11_), 
        .A_10_(A1_10_), .A_9_(A1_9_), .A_8_(A1_8_), .A_7_(A1_7_), .A_6_(A1_6_), 
        .A_5_(PROD1_7_), .B_21_(n5), .B_20_(n25), .B_19_(n23), .B_18_(n22), 
        .B_17_(n8), .B_16_(n24), .SUM_21_(PRODUCT_23_), .SUM_20_(PRODUCT_22_), 
        .SUM_19_(PRODUCT_21_), .SUM_18_(PRODUCT_20_), .SUM_17_(PRODUCT_19_), 
        .SUM_16_(PRODUCT_18_), .SUM_15_(PRODUCT_17_), .SUM_14_(PRODUCT_16_), 
        .SUM_13_(PRODUCT_15_), .SUM_12_(PRODUCT_14_), .SUM_11_(PRODUCT_13_), 
        .SUM_10_(PRODUCT_12_), .SUM_9_(PRODUCT_11_), .SUM_8_(PRODUCT_10_), 
        .SUM_7_(PRODUCT_9_), .SUM_6_(PRODUCT_8_), .SUM_5_(PRODUCT_7_) );
  ADDFHX4 S4_2 ( .A(ab_16__2_), .B(CARRYB_15__2_), .CI(SUMB_15__3_), .CO(
        CARRYB_16__2_), .S(SUMB_16__2_) );
  ADDFHX4 S2_15_2 ( .A(ab_15__2_), .B(CARRYB_14__2_), .CI(SUMB_14__3_), .CO(
        CARRYB_15__2_), .S(SUMB_15__2_) );
  ADDFHX4 S2_15_1 ( .A(ab_15__1_), .B(CARRYB_14__1_), .CI(SUMB_14__2_), .CO(
        CARRYB_15__1_), .S(SUMB_15__1_) );
  ADDFHX4 S4_1 ( .A(ab_16__1_), .B(CARRYB_15__1_), .CI(SUMB_15__2_), .CO(
        CARRYB_16__1_), .S(SUMB_16__1_) );
  ADDFHX4 S4_0 ( .A(ab_16__0_), .B(CARRYB_15__0_), .CI(SUMB_15__1_), .CO(
        CARRYB_16__0_), .S(SUMB_16__0_) );
  ADDFHX4 S1_9_0 ( .A(ab_9__0_), .B(CARRYB_8__0_), .CI(SUMB_8__1_), .CO(
        CARRYB_9__0_), .S(A1_7_) );
  ADDFHX4 S1_10_0 ( .A(ab_10__0_), .B(CARRYB_9__0_), .CI(SUMB_9__1_), .CO(
        CARRYB_10__0_), .S(A1_8_) );
  ADDFHX4 S2_13_2 ( .A(ab_13__2_), .B(CARRYB_12__2_), .CI(SUMB_12__3_), .CO(
        CARRYB_13__2_), .S(SUMB_13__2_) );
  ADDFHX4 S1_7_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(PROD1_7_) );
  ADDFHX4 S1_8_0 ( .A(ab_8__0_), .B(CARRYB_7__0_), .CI(SUMB_7__1_), .CO(
        CARRYB_8__0_), .S(A1_6_) );
  ADDFHX4 S1_14_0 ( .A(ab_14__0_), .B(CARRYB_13__0_), .CI(SUMB_13__1_), .CO(
        CARRYB_14__0_), .S(A1_12_) );
  ADDFHX4 S1_15_0 ( .A(ab_15__0_), .B(SUMB_14__1_), .CI(CARRYB_14__0_), .CO(
        CARRYB_15__0_), .S(A1_13_) );
  ADDFHX4 S1_12_0 ( .A(ab_12__0_), .B(CARRYB_11__0_), .CI(SUMB_11__1_), .CO(
        CARRYB_12__0_), .S(A1_10_) );
  ADDFHX4 S1_13_0 ( .A(ab_13__0_), .B(CARRYB_12__0_), .CI(SUMB_12__1_), .CO(
        CARRYB_13__0_), .S(A1_11_) );
  ADDFHX4 S2_13_1 ( .A(ab_13__1_), .B(CARRYB_12__1_), .CI(SUMB_12__2_), .CO(
        CARRYB_13__1_), .S(SUMB_13__1_) );
  ADDFHX4 S2_14_3 ( .A(ab_14__3_), .B(CARRYB_13__3_), .CI(SUMB_13__4_), .CO(
        CARRYB_14__3_), .S(SUMB_14__3_) );
  ADDFHX4 S2_15_3 ( .A(ab_15__3_), .B(CARRYB_14__3_), .CI(SUMB_14__4_), .CO(
        CARRYB_15__3_), .S(SUMB_15__3_) );
  ADDFHX4 S2_14_1 ( .A(ab_14__1_), .B(CARRYB_13__1_), .CI(SUMB_13__2_), .CO(
        CARRYB_14__1_), .S(SUMB_14__1_) );
  ADDFHX4 S2_14_2 ( .A(ab_14__2_), .B(CARRYB_13__2_), .CI(SUMB_13__3_), .CO(
        CARRYB_14__2_), .S(SUMB_14__2_) );
  ADDFHX1 S3_15_6 ( .A(ab_15__6_), .B(CARRYB_14__6_), .CI(ab_14__7_), .CO(
        CARRYB_15__6_), .S(SUMB_15__6_) );
  ADDFHX4 S2_12_1 ( .A(ab_12__1_), .B(CARRYB_11__1_), .CI(SUMB_11__2_), .CO(
        CARRYB_12__1_), .S(SUMB_12__1_) );
  ADDFHX4 S4_3 ( .A(ab_16__3_), .B(CARRYB_15__3_), .CI(SUMB_15__4_), .CO(
        CARRYB_16__3_), .S(SUMB_16__3_) );
  ADDFHX4 S4_5 ( .A(ab_16__5_), .B(CARRYB_15__5_), .CI(SUMB_15__6_), .CO(
        CARRYB_16__5_), .S(SUMB_16__5_) );
  ADDFHX4 S4_4 ( .A(ab_16__4_), .B(CARRYB_15__4_), .CI(SUMB_15__5_), .CO(
        CARRYB_16__4_), .S(SUMB_16__4_) );
  ADDFHX4 S2_10_5 ( .A(ab_10__5_), .B(CARRYB_9__5_), .CI(SUMB_9__6_), .CO(
        CARRYB_10__5_), .S(SUMB_10__5_) );
  ADDFHX4 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  ADDFHX4 S2_13_4 ( .A(ab_13__4_), .B(CARRYB_12__4_), .CI(SUMB_12__5_), .CO(
        CARRYB_13__4_), .S(SUMB_13__4_) );
  ADDFHX4 S2_14_4 ( .A(ab_14__4_), .B(CARRYB_13__4_), .CI(SUMB_13__5_), .CO(
        CARRYB_14__4_), .S(SUMB_14__4_) );
  ADDFHX4 S2_11_4 ( .A(ab_11__4_), .B(CARRYB_10__4_), .CI(SUMB_10__5_), .CO(
        CARRYB_11__4_), .S(SUMB_11__4_) );
  ADDFHX4 S3_2_6 ( .A(ab_2__6_), .B(n9), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  ADDFHX4 S2_11_1 ( .A(ab_11__1_), .B(CARRYB_10__1_), .CI(SUMB_10__2_), .CO(
        CARRYB_11__1_), .S(SUMB_11__1_) );
  ADDFHX4 S2_9_5 ( .A(ab_9__5_), .B(CARRYB_8__5_), .CI(SUMB_8__6_), .CO(
        CARRYB_9__5_), .S(SUMB_9__5_) );
  ADDFHX4 S2_11_2 ( .A(ab_11__2_), .B(CARRYB_10__2_), .CI(SUMB_10__3_), .CO(
        CARRYB_11__2_), .S(SUMB_11__2_) );
  ADDFHX4 S2_12_2 ( .A(ab_12__2_), .B(CARRYB_11__2_), .CI(SUMB_11__3_), .CO(
        CARRYB_12__2_), .S(SUMB_12__2_) );
  ADDFHX4 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  ADDFHX4 S2_7_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  ADDFHX4 S2_11_5 ( .A(ab_11__5_), .B(CARRYB_10__5_), .CI(SUMB_10__6_), .CO(
        CARRYB_11__5_), .S(SUMB_11__5_) );
  ADDFHX4 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  ADDFHX4 S2_10_2 ( .A(ab_10__2_), .B(CARRYB_9__2_), .CI(SUMB_9__3_), .CO(
        CARRYB_10__2_), .S(SUMB_10__2_) );
  ADDFHX4 S3_9_6 ( .A(ab_9__6_), .B(CARRYB_8__6_), .CI(ab_8__7_), .CO(
        CARRYB_9__6_), .S(SUMB_9__6_) );
  ADDFHX4 S3_8_6 ( .A(ab_8__6_), .B(CARRYB_7__6_), .CI(ab_7__7_), .CO(
        CARRYB_8__6_), .S(SUMB_8__6_) );
  ADDFHX4 S2_9_4 ( .A(ab_9__4_), .B(CARRYB_8__4_), .CI(SUMB_8__5_), .CO(
        CARRYB_9__4_), .S(SUMB_9__4_) );
  ADDFHX4 S2_10_4 ( .A(ab_10__4_), .B(CARRYB_9__4_), .CI(SUMB_9__5_), .CO(
        CARRYB_10__4_), .S(SUMB_10__4_) );
  ADDFHX4 S2_7_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  ADDFHX4 S2_7_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  ADDFHX4 S2_8_3 ( .A(ab_8__3_), .B(CARRYB_7__3_), .CI(SUMB_7__4_), .CO(
        CARRYB_8__3_), .S(SUMB_8__3_) );
  ADDFHX4 S2_12_3 ( .A(ab_12__3_), .B(CARRYB_11__3_), .CI(SUMB_11__4_), .CO(
        CARRYB_12__3_), .S(SUMB_12__3_) );
  ADDFHX4 S2_13_3 ( .A(ab_13__3_), .B(CARRYB_12__3_), .CI(SUMB_12__4_), .CO(
        CARRYB_13__3_), .S(SUMB_13__3_) );
  ADDFHX4 S2_9_2 ( .A(ab_9__2_), .B(CARRYB_8__2_), .CI(SUMB_8__3_), .CO(
        CARRYB_9__2_), .S(SUMB_9__2_) );
  ADDFHX4 S3_11_6 ( .A(ab_11__6_), .B(CARRYB_10__6_), .CI(ab_10__7_), .CO(
        CARRYB_11__6_), .S(SUMB_11__6_) );
  ADDFHX4 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  ADDFHX4 S2_10_3 ( .A(ab_10__3_), .B(CARRYB_9__3_), .CI(SUMB_9__4_), .CO(
        CARRYB_10__3_), .S(SUMB_10__3_) );
  ADDFHX4 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  ADDFHX2 S2_15_5 ( .A(ab_15__5_), .B(CARRYB_14__5_), .CI(SUMB_14__6_), .CO(
        CARRYB_15__5_), .S(SUMB_15__5_) );
  ADDFHX4 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  ADDFHX4 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  ADDFHX4 S2_8_5 ( .A(ab_8__5_), .B(CARRYB_7__5_), .CI(SUMB_7__6_), .CO(
        CARRYB_8__5_), .S(SUMB_8__5_) );
  ADDFHX4 S2_8_2 ( .A(ab_8__2_), .B(CARRYB_7__2_), .CI(SUMB_7__3_), .CO(
        CARRYB_8__2_), .S(SUMB_8__2_) );
  ADDFHX4 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  ADDFHX4 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  ADDFHX4 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  ADDFHX4 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  ADDFHX4 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  ADDFHX4 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  ADDFHX4 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  ADDFHX4 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  ADDFHX4 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  ADDFHX4 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  ADDFHX4 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  ADDFHX4 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  ADDFHX4 S3_7_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(
        CARRYB_7__6_), .S(SUMB_7__6_) );
  ADDFHX4 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  ADDFHX4 S2_2_5 ( .A(ab_2__5_), .B(n7), .CI(SUMB_1__6_), .CO(CARRYB_2__5_), 
        .S(SUMB_2__5_) );
  ADDFHX4 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  ADDFHX4 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  ADDFHX4 S3_10_6 ( .A(ab_10__6_), .B(CARRYB_9__6_), .CI(ab_9__7_), .CO(
        CARRYB_10__6_), .S(SUMB_10__6_) );
  ADDFHX4 S2_7_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  ADDFHX4 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  ADDFHX4 S2_9_1 ( .A(ab_9__1_), .B(CARRYB_8__1_), .CI(SUMB_8__2_), .CO(
        CARRYB_9__1_), .S(SUMB_9__1_) );
  ADDFHX4 S2_10_1 ( .A(ab_10__1_), .B(CARRYB_9__1_), .CI(SUMB_9__2_), .CO(
        CARRYB_10__1_), .S(SUMB_10__1_) );
  ADDFHX4 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  ADDFHX4 S2_8_4 ( .A(ab_8__4_), .B(CARRYB_7__4_), .CI(SUMB_7__5_), .CO(
        CARRYB_8__4_), .S(SUMB_8__4_) );
  ADDFHX4 S2_12_4 ( .A(ab_12__4_), .B(CARRYB_11__4_), .CI(SUMB_11__5_), .CO(
        CARRYB_12__4_), .S(SUMB_12__4_) );
  ADDFHX4 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  ADDFHX4 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  ADDFHX4 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  ADDFHX4 S2_11_3 ( .A(ab_11__3_), .B(CARRYB_10__3_), .CI(SUMB_10__4_), .CO(
        CARRYB_11__3_), .S(SUMB_11__3_) );
  ADDFHX4 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  ADDFHX2 S3_14_6 ( .A(ab_14__6_), .B(CARRYB_13__6_), .CI(ab_13__7_), .CO(
        CARRYB_14__6_), .S(SUMB_14__6_) );
  ADDFHX4 S2_12_5 ( .A(ab_12__5_), .B(CARRYB_11__5_), .CI(SUMB_11__6_), .CO(
        CARRYB_12__5_), .S(SUMB_12__5_) );
  ADDFHX4 S2_13_5 ( .A(ab_13__5_), .B(CARRYB_12__5_), .CI(SUMB_12__6_), .CO(
        CARRYB_13__5_), .S(SUMB_13__5_) );
  ADDFHX4 S2_9_3 ( .A(ab_9__3_), .B(CARRYB_8__3_), .CI(SUMB_8__4_), .CO(
        CARRYB_9__3_), .S(SUMB_9__3_) );
  ADDFHX4 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  ADDFHX4 S2_2_4 ( .A(ab_2__4_), .B(n10), .CI(SUMB_1__5_), .CO(CARRYB_2__4_), 
        .S(SUMB_2__4_) );
  ADDFHX4 S2_8_1 ( .A(ab_8__1_), .B(CARRYB_7__1_), .CI(SUMB_7__2_), .CO(
        CARRYB_8__1_), .S(SUMB_8__1_) );
  ADDFHX4 S2_7_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  ADDFHX4 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  ADDFHX4 S3_13_6 ( .A(ab_13__6_), .B(ab_12__7_), .CI(CARRYB_12__6_), .CO(
        CARRYB_13__6_), .S(SUMB_13__6_) );
  ADDFHX4 S1_11_0 ( .A(ab_11__0_), .B(CARRYB_10__0_), .CI(SUMB_10__1_), .CO(
        CARRYB_11__0_), .S(A1_9_) );
  ADDFHX4 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  ADDFHX4 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  ADDFHX2 S3_12_6 ( .A(ab_12__6_), .B(CARRYB_11__6_), .CI(ab_11__7_), .CO(
        CARRYB_12__6_), .S(SUMB_12__6_) );
  ADDFHX4 S2_15_4 ( .A(ab_15__4_), .B(CARRYB_14__4_), .CI(SUMB_14__5_), .CO(
        CARRYB_15__4_), .S(SUMB_15__4_) );
  ADDFHX4 S2_14_5 ( .A(ab_14__5_), .B(CARRYB_13__5_), .CI(SUMB_13__6_), .CO(
        CARRYB_14__5_), .S(SUMB_14__5_) );
  BUFX20 U2 ( .A(n44), .Y(n29) );
  AND2X4 U3 ( .A(A[1]), .B(B[2]), .Y(ab_1__2_) );
  AND2X4 U4 ( .A(A[1]), .B(B[3]), .Y(ab_1__3_) );
  BUFX12 U5 ( .A(n46), .Y(n33) );
  NOR2BX4 U6 ( .AN(A[3]), .B(n31), .Y(ab_3__4_) );
  AND2X2 U7 ( .A(A[3]), .B(B[0]), .Y(ab_3__0_) );
  NOR2BX1 U8 ( .AN(n13), .B(n31), .Y(ab_7__4_) );
  BUFX12 U9 ( .A(A[7]), .Y(n13) );
  NOR2BX2 U10 ( .AN(A[4]), .B(n39), .Y(ab_4__6_) );
  NOR2BX2 U11 ( .AN(A[4]), .B(n37), .Y(ab_4__1_) );
  NOR2BXL U12 ( .AN(A[4]), .B(n40), .Y(ab_4__0_) );
  BUFX16 U13 ( .A(n44), .Y(n30) );
  INVX8 U14 ( .A(B[5]), .Y(n44) );
  BUFX20 U15 ( .A(n47), .Y(n35) );
  INVX8 U16 ( .A(B[2]), .Y(n47) );
  NOR2BX1 U17 ( .AN(A[8]), .B(n37), .Y(ab_8__1_) );
  NAND2X4 U18 ( .A(n18), .B(SUMB_16__3_), .Y(n21) );
  CLKINVX4 U19 ( .A(n46), .Y(n3) );
  BUFX16 U20 ( .A(A[2]), .Y(n4) );
  AND2X1 U21 ( .A(CARRYB_16__5_), .B(SUMB_16__6_), .Y(n5) );
  INVX8 U22 ( .A(B[4]), .Y(n45) );
  CLKBUFX20 U23 ( .A(n45), .Y(n31) );
  NOR2BX2 U24 ( .AN(A[14]), .B(n34), .Y(ab_14__3_) );
  NOR2BX2 U25 ( .AN(A[16]), .B(n34), .Y(ab_16__3_) );
  NOR2BX2 U26 ( .AN(A[3]), .B(n35), .Y(ab_3__2_) );
  NOR2BX1 U27 ( .AN(A[16]), .B(n38), .Y(ab_16__1_) );
  NAND2X2 U28 ( .A(n14), .B(SUMB_16__5_), .Y(n17) );
  NOR2BX1 U29 ( .AN(n4), .B(n40), .Y(ab_2__0_) );
  NOR2BX2 U30 ( .AN(A[12]), .B(n34), .Y(ab_12__3_) );
  NOR2BX1 U31 ( .AN(A[13]), .B(n32), .Y(ab_13__4_) );
  INVX1 U32 ( .A(n41), .Y(n11) );
  NOR2BX1 U33 ( .AN(A[11]), .B(n36), .Y(ab_11__2_) );
  NOR2BX1 U34 ( .AN(A[9]), .B(n38), .Y(ab_9__1_) );
  AND2X4 U36 ( .A(ab_0__6_), .B(ab_1__5_), .Y(n7) );
  AND2X4 U37 ( .A(CARRYB_16__1_), .B(SUMB_16__2_), .Y(n8) );
  AND2X4 U38 ( .A(ab_0__7_), .B(ab_1__6_), .Y(n9) );
  NOR2BX1 U39 ( .AN(A[3]), .B(n50), .Y(ab_3__7_) );
  NOR2BXL U40 ( .AN(A[6]), .B(n39), .Y(ab_6__6_) );
  NOR2BX1 U41 ( .AN(n13), .B(n37), .Y(ab_7__1_) );
  NOR2BX4 U42 ( .AN(n3), .B(n41), .Y(ab_0__3_) );
  NAND2X4 U43 ( .A(ab_1__3_), .B(ab_0__4_), .Y(n28) );
  AND2X4 U44 ( .A(ab_1__4_), .B(ab_0__5_), .Y(n10) );
  INVX4 U45 ( .A(B[6]), .Y(n43) );
  XOR2X4 U46 ( .A(ab_1__2_), .B(ab_0__3_), .Y(SUMB_1__2_) );
  NOR2BX1 U47 ( .AN(A[0]), .B(n40), .Y(n42) );
  INVX12 U48 ( .A(A[0]), .Y(n41) );
  NOR2BX1 U49 ( .AN(A[8]), .B(n35), .Y(ab_8__2_) );
  NOR2BX2 U50 ( .AN(A[4]), .B(n33), .Y(ab_4__3_) );
  NAND2X4 U51 ( .A(ab_1__2_), .B(ab_0__3_), .Y(n27) );
  NOR2BX1 U52 ( .AN(n13), .B(n35), .Y(ab_7__2_) );
  INVX4 U53 ( .A(n27), .Y(CARRYB_1__2_) );
  NOR2BX1 U54 ( .AN(A[6]), .B(n35), .Y(ab_6__2_) );
  INVX4 U55 ( .A(ab_0__4_), .Y(n12) );
  NOR2BX1 U56 ( .AN(A[8]), .B(n33), .Y(ab_8__3_) );
  INVX4 U57 ( .A(SUMB_16__3_), .Y(n19) );
  AND2X4 U58 ( .A(B[6]), .B(n11), .Y(ab_0__6_) );
  NOR2BX1 U59 ( .AN(n13), .B(n33), .Y(ab_7__3_) );
  AND2X4 U60 ( .A(A[1]), .B(B[6]), .Y(ab_1__6_) );
  XOR2X4 U61 ( .A(ab_1__5_), .B(ab_0__6_), .Y(SUMB_1__5_) );
  AND2X4 U62 ( .A(CARRYB_16__0_), .B(SUMB_16__1_), .Y(n24) );
  XOR2X2 U63 ( .A(n51), .B(ab_0__2_), .Y(SUMB_1__1_) );
  NAND2X4 U64 ( .A(ab_0__2_), .B(n51), .Y(n26) );
  INVX4 U65 ( .A(n26), .Y(CARRYB_1__1_) );
  XNOR2X4 U66 ( .A(ab_1__3_), .B(n12), .Y(SUMB_1__3_) );
  NOR2BX1 U67 ( .AN(A[1]), .B(n50), .Y(ab_1__7_) );
  AND3X1 U68 ( .A(A[1]), .B(B[1]), .C(n42), .Y(CARRYB_1__0_) );
  NOR2BX2 U69 ( .AN(A[3]), .B(n37), .Y(ab_3__1_) );
  NOR2BX2 U70 ( .AN(n4), .B(n35), .Y(ab_2__2_) );
  NOR2BX2 U71 ( .AN(n4), .B(n31), .Y(ab_2__4_) );
  NOR2BX2 U72 ( .AN(n4), .B(n37), .Y(ab_2__1_) );
  NOR2BX2 U73 ( .AN(n4), .B(n33), .Y(ab_2__3_) );
  BUFX20 U74 ( .A(n46), .Y(n34) );
  CLKINVX4 U75 ( .A(CARRYB_16__2_), .Y(n18) );
  INVX8 U76 ( .A(B[3]), .Y(n46) );
  BUFX20 U77 ( .A(n43), .Y(n39) );
  NOR2BX2 U78 ( .AN(A[3]), .B(n33), .Y(ab_3__3_) );
  NAND2X4 U79 ( .A(n19), .B(CARRYB_16__2_), .Y(n20) );
  XOR2X4 U80 ( .A(ab_1__4_), .B(ab_0__5_), .Y(SUMB_1__4_) );
  INVX20 U81 ( .A(B[7]), .Y(n50) );
  NOR2BX2 U82 ( .AN(A[5]), .B(n39), .Y(ab_5__6_) );
  NOR2BX2 U83 ( .AN(A[5]), .B(n29), .Y(ab_5__5_) );
  NOR2BX2 U84 ( .AN(A[5]), .B(n31), .Y(ab_5__4_) );
  NOR2BX2 U85 ( .AN(A[5]), .B(n33), .Y(ab_5__3_) );
  NOR2BX2 U86 ( .AN(A[5]), .B(n37), .Y(ab_5__1_) );
  NOR2BX4 U87 ( .AN(n4), .B(n39), .Y(ab_2__6_) );
  NOR2BX2 U88 ( .AN(B[2]), .B(n41), .Y(ab_0__2_) );
  INVX4 U89 ( .A(n28), .Y(CARRYB_1__3_) );
  NOR2BX2 U90 ( .AN(A[3]), .B(n29), .Y(ab_3__5_) );
  NOR2BX1 U91 ( .AN(A[6]), .B(n30), .Y(ab_6__5_) );
  XOR2X4 U92 ( .A(SUMB_16__1_), .B(CARRYB_16__0_), .Y(A1_15_) );
  NOR2BX4 U93 ( .AN(B[5]), .B(n41), .Y(ab_0__5_) );
  XOR2X4 U94 ( .A(CARRYB_16__3_), .B(SUMB_16__4_), .Y(A1_18_) );
  NOR2BX2 U95 ( .AN(A[3]), .B(n39), .Y(ab_3__6_) );
  XOR2X4 U96 ( .A(ab_1__6_), .B(ab_0__7_), .Y(SUMB_1__6_) );
  NOR2BX4 U97 ( .AN(B[4]), .B(n41), .Y(ab_0__4_) );
  NOR2BX2 U98 ( .AN(n4), .B(n30), .Y(ab_2__5_) );
  NOR2BX4 U99 ( .AN(B[7]), .B(n41), .Y(ab_0__7_) );
  NOR2BX2 U100 ( .AN(A[4]), .B(n30), .Y(ab_4__5_) );
  NOR2BX2 U101 ( .AN(A[5]), .B(n35), .Y(ab_5__2_) );
  NAND2X4 U102 ( .A(CARRYB_16__4_), .B(n15), .Y(n16) );
  NAND2X4 U103 ( .A(n16), .B(n17), .Y(A1_19_) );
  INVX1 U104 ( .A(CARRYB_16__4_), .Y(n14) );
  INVX4 U105 ( .A(SUMB_16__5_), .Y(n15) );
  NAND2X4 U106 ( .A(n20), .B(n21), .Y(A1_17_) );
  NOR2BX2 U107 ( .AN(A[4]), .B(n35), .Y(ab_4__2_) );
  NOR2BX1 U108 ( .AN(A[14]), .B(n40), .Y(ab_14__0_) );
  NOR2BXL U109 ( .AN(A[10]), .B(n39), .Y(ab_10__6_) );
  NOR2BX1 U110 ( .AN(A[9]), .B(n32), .Y(ab_9__4_) );
  NOR2BX1 U111 ( .AN(n4), .B(n50), .Y(ab_2__7_) );
  NOR2BX1 U112 ( .AN(A[15]), .B(n40), .Y(ab_15__0_) );
  NOR2BXL U113 ( .AN(A[16]), .B(n40), .Y(ab_16__0_) );
  CLKBUFXL U114 ( .A(n47), .Y(n36) );
  BUFX8 U115 ( .A(n48), .Y(n37) );
  CLKBUFXL U116 ( .A(n48), .Y(n38) );
  NOR2BX1 U117 ( .AN(A[10]), .B(n38), .Y(ab_10__1_) );
  NOR2BX1 U118 ( .AN(A[12]), .B(n30), .Y(ab_12__5_) );
  NOR2BX1 U119 ( .AN(A[9]), .B(n39), .Y(ab_9__6_) );
  NOR2BX1 U120 ( .AN(A[10]), .B(n36), .Y(ab_10__2_) );
  NOR2BXL U121 ( .AN(A[10]), .B(n50), .Y(ab_10__7_) );
  NOR2BX1 U122 ( .AN(A[11]), .B(n39), .Y(ab_11__6_) );
  NOR2BX1 U123 ( .AN(A[13]), .B(n34), .Y(ab_13__3_) );
  NOR2BX1 U124 ( .AN(A[9]), .B(n36), .Y(ab_9__2_) );
  NOR2BX1 U125 ( .AN(A[12]), .B(n32), .Y(ab_12__4_) );
  NOR2BX1 U126 ( .AN(A[11]), .B(n32), .Y(ab_11__4_) );
  NOR2BX1 U127 ( .AN(A[10]), .B(n32), .Y(ab_10__4_) );
  NOR2BX1 U128 ( .AN(A[10]), .B(n30), .Y(ab_10__5_) );
  NOR2BX1 U129 ( .AN(n13), .B(n29), .Y(ab_7__5_) );
  NOR2BXL U130 ( .AN(A[8]), .B(n30), .Y(ab_8__5_) );
  NOR2BX1 U131 ( .AN(A[5]), .B(n50), .Y(ab_5__7_) );
  NOR2BX2 U132 ( .AN(A[9]), .B(n34), .Y(ab_9__3_) );
  NOR2BX1 U133 ( .AN(A[9]), .B(n50), .Y(ab_9__7_) );
  NOR2BX1 U134 ( .AN(A[11]), .B(n29), .Y(ab_11__5_) );
  NOR2BX1 U135 ( .AN(n13), .B(n50), .Y(ab_7__7_) );
  NOR2BX1 U136 ( .AN(A[13]), .B(n38), .Y(ab_13__1_) );
  NOR2BX1 U137 ( .AN(A[13]), .B(n36), .Y(ab_13__2_) );
  NOR2BX1 U138 ( .AN(A[14]), .B(n32), .Y(ab_14__4_) );
  NOR2BXL U139 ( .AN(A[12]), .B(n39), .Y(ab_12__6_) );
  NOR2BXL U140 ( .AN(A[8]), .B(n40), .Y(ab_8__0_) );
  NOR2BXL U141 ( .AN(A[12]), .B(n50), .Y(ab_12__7_) );
  NOR2BX4 U142 ( .AN(A[1]), .B(n29), .Y(ab_1__5_) );
  NOR2BX4 U143 ( .AN(A[1]), .B(n31), .Y(ab_1__4_) );
  NOR2BX1 U144 ( .AN(A[15]), .B(n38), .Y(ab_15__1_) );
  NOR2BX1 U145 ( .AN(A[15]), .B(n36), .Y(ab_15__2_) );
  NOR2BX4 U146 ( .AN(A[1]), .B(n37), .Y(n51) );
  NOR2BX1 U147 ( .AN(A[15]), .B(n34), .Y(ab_15__3_) );
  CLKBUFXL U148 ( .A(n45), .Y(n32) );
  NOR2BX1 U149 ( .AN(A[6]), .B(n50), .Y(ab_6__7_) );
  NOR2BX1 U150 ( .AN(n13), .B(n39), .Y(ab_7__6_) );
  NOR2BX1 U151 ( .AN(A[11]), .B(n40), .Y(ab_11__0_) );
  NOR2BXL U152 ( .AN(A[11]), .B(n38), .Y(ab_11__1_) );
  NOR2BX1 U153 ( .AN(A[5]), .B(n40), .Y(ab_5__0_) );
  NOR2BX1 U154 ( .AN(A[4]), .B(n50), .Y(ab_4__7_) );
  NOR2BX1 U155 ( .AN(A[13]), .B(n29), .Y(ab_13__5_) );
  NOR2BXL U156 ( .AN(A[11]), .B(n50), .Y(ab_11__7_) );
  AND2X2 U157 ( .A(SUMB_16__3_), .B(CARRYB_16__2_), .Y(n22) );
  AND2X2 U158 ( .A(CARRYB_16__3_), .B(SUMB_16__4_), .Y(n23) );
  NOR2BX1 U159 ( .AN(A[14]), .B(n30), .Y(ab_14__5_) );
  NOR2BXL U160 ( .AN(A[13]), .B(n50), .Y(ab_13__7_) );
  NOR2BXL U161 ( .AN(A[14]), .B(n39), .Y(ab_14__6_) );
  NOR2BXL U162 ( .AN(A[13]), .B(n39), .Y(ab_13__6_) );
  NOR2BX1 U163 ( .AN(A[12]), .B(n40), .Y(ab_12__0_) );
  NOR2BX1 U164 ( .AN(n13), .B(n40), .Y(ab_7__0_) );
  NOR2BX1 U165 ( .AN(A[6]), .B(n40), .Y(ab_6__0_) );
  NOR2BX1 U166 ( .AN(A[12]), .B(n38), .Y(ab_12__1_) );
  NOR2BXL U167 ( .AN(A[10]), .B(n34), .Y(ab_10__3_) );
  NOR2BXL U168 ( .AN(A[8]), .B(n39), .Y(ab_8__6_) );
  NOR2BX1 U169 ( .AN(A[4]), .B(n31), .Y(ab_4__4_) );
  NOR2BX1 U170 ( .AN(A[13]), .B(n40), .Y(ab_13__0_) );
  NOR2BX1 U171 ( .AN(A[14]), .B(n38), .Y(ab_14__1_) );
  NOR2BX1 U172 ( .AN(A[14]), .B(n36), .Y(ab_14__2_) );
  NOR2BX1 U173 ( .AN(A[9]), .B(n40), .Y(ab_9__0_) );
  NOR2BX1 U174 ( .AN(A[12]), .B(n36), .Y(ab_12__2_) );
  NOR2BXL U175 ( .AN(A[6]), .B(n37), .Y(ab_6__1_) );
  NOR2BXL U176 ( .AN(A[11]), .B(n34), .Y(ab_11__3_) );
  NOR2BX1 U177 ( .AN(A[9]), .B(n29), .Y(ab_9__5_) );
  NOR2BXL U178 ( .AN(A[8]), .B(n31), .Y(ab_8__4_) );
  NOR2BXL U179 ( .AN(A[8]), .B(n50), .Y(ab_8__7_) );
  NOR2BXL U180 ( .AN(A[6]), .B(n31), .Y(ab_6__4_) );
  NOR2BXL U181 ( .AN(A[6]), .B(n33), .Y(ab_6__3_) );
  NOR2BX1 U182 ( .AN(A[10]), .B(n40), .Y(ab_10__0_) );
  XOR2X2 U183 ( .A(CARRYB_16__5_), .B(SUMB_16__6_), .Y(A1_20_) );
  AND2X2 U184 ( .A(CARRYB_16__4_), .B(SUMB_16__5_), .Y(n25) );
  BUFX3 U185 ( .A(n49), .Y(n40) );
  INVX1 U186 ( .A(B[0]), .Y(n49) );
  INVX1 U187 ( .A(B[1]), .Y(n48) );
  NOR2BX1 U188 ( .AN(A[16]), .B(n30), .Y(ab_16__5_) );
  NOR2BX1 U189 ( .AN(A[16]), .B(n32), .Y(ab_16__4_) );
  NOR2BX1 U190 ( .AN(A[16]), .B(n36), .Y(ab_16__2_) );
  NOR2BXL U191 ( .AN(A[15]), .B(n32), .Y(ab_15__4_) );
  NOR2BXL U192 ( .AN(A[15]), .B(n29), .Y(ab_15__5_) );
  NOR2BXL U193 ( .AN(A[14]), .B(n50), .Y(ab_14__7_) );
  NOR2BXL U194 ( .AN(A[15]), .B(n39), .Y(ab_15__6_) );
  NOR2BXL U195 ( .AN(A[16]), .B(n39), .Y(ab_16__6_) );
  NOR2BXL U196 ( .AN(A[15]), .B(n50), .Y(ab_15__7_) );
  NOR2BXL U197 ( .AN(A[16]), .B(n50), .Y(ab_16__7_) );
  XOR2X4 U198 ( .A(CARRYB_16__6_), .B(ab_16__7_), .Y(A1_21_) );
  XOR2X4 U199 ( .A(CARRYB_16__1_), .B(SUMB_16__2_), .Y(A1_16_) );
endmodule


module multi16_7 ( in_17bit, in_8bit, out );
  input [16:0] in_17bit;
  input [7:0] in_8bit;
  output [16:0] out;
  wire   n121, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119;
  wire   [16:1] in_17bit_b;
  wire   [7:1] in_8bit_b;
  wire   [23:8] mul;

  multi16_7_DW02_mult_0 mult_55 ( .A({in_17bit_b, in_17bit[0]}), .B({in_8bit_b, 
        in_8bit[0]}), .PRODUCT_23_(mul[23]), .PRODUCT_22_(mul[22]), 
        .PRODUCT_21_(mul[21]), .PRODUCT_20_(mul[20]), .PRODUCT_19_(mul[19]), 
        .PRODUCT_18_(mul[18]), .PRODUCT_17_(mul[17]), .PRODUCT_16_(mul[16]), 
        .PRODUCT_15_(mul[15]), .PRODUCT_14_(mul[14]), .PRODUCT_13_(mul[13]), 
        .PRODUCT_12_(mul[12]), .PRODUCT_11_(mul[11]), .PRODUCT_10_(mul[10]), 
        .PRODUCT_9_(mul[9]), .PRODUCT_8_(mul[8]), .PRODUCT_7_(out[0]) );
  INVX8 U2 ( .A(mul[21]), .Y(n115) );
  BUFX8 U3 ( .A(n65), .Y(n1) );
  CLKINVX2 U4 ( .A(n52), .Y(n92) );
  XNOR2X1 U5 ( .A(n52), .B(in_8bit[7]), .Y(n117) );
  XNOR2X2 U6 ( .A(n74), .B(n47), .Y(in_17bit_b[7]) );
  AND2X4 U7 ( .A(n111), .B(n110), .Y(n2) );
  NOR2X1 U8 ( .A(n1), .B(in_17bit[3]), .Y(n3) );
  INVX3 U9 ( .A(in_8bit[2]), .Y(n16) );
  NAND3BX4 U10 ( .AN(n4), .B(n50), .C(n15), .Y(n49) );
  NOR2X4 U11 ( .A(in_17bit[1]), .B(n52), .Y(n4) );
  OAI21X4 U12 ( .A0(n17), .A1(n55), .B0(in_8bit[7]), .Y(n56) );
  INVX3 U13 ( .A(in_8bit[5]), .Y(n54) );
  INVX4 U14 ( .A(n54), .Y(n14) );
  XNOR2X2 U15 ( .A(mul[11]), .B(n30), .Y(out[4]) );
  NOR2X4 U16 ( .A(n12), .B(n61), .Y(n57) );
  NAND2X2 U17 ( .A(n27), .B(mul[18]), .Y(n7) );
  NAND2X4 U18 ( .A(n5), .B(n6), .Y(n8) );
  NAND2X4 U19 ( .A(n7), .B(n8), .Y(out[11]) );
  INVX4 U20 ( .A(n27), .Y(n5) );
  INVX8 U21 ( .A(mul[18]), .Y(n6) );
  NAND2X2 U22 ( .A(n53), .B(n54), .Y(n9) );
  NAND2X4 U23 ( .A(n10), .B(n12), .Y(n62) );
  CLKINVX4 U24 ( .A(n9), .Y(n10) );
  XOR2X4 U25 ( .A(n60), .B(n11), .Y(in_8bit_b[6]) );
  CLKINVX20 U26 ( .A(in_8bit[6]), .Y(n11) );
  INVXL U27 ( .A(n112), .Y(n13) );
  INVX1 U28 ( .A(n87), .Y(n89) );
  XNOR2X2 U29 ( .A(mul[8]), .B(n94), .Y(out[1]) );
  NAND2X4 U30 ( .A(n52), .B(n65), .Y(n36) );
  OR2X4 U31 ( .A(mul[12]), .B(n98), .Y(n99) );
  BUFX8 U32 ( .A(n59), .Y(n12) );
  NOR2BX4 U33 ( .AN(n105), .B(n13), .Y(n23) );
  AOI21X1 U34 ( .A0(n118), .A1(n2), .B0(n117), .Y(n119) );
  NAND2X4 U35 ( .A(n112), .B(n109), .Y(n38) );
  INVX8 U36 ( .A(n16), .Y(n17) );
  CLKINVX4 U37 ( .A(n107), .Y(n19) );
  NAND2X4 U38 ( .A(n107), .B(n37), .Y(n109) );
  INVX8 U39 ( .A(mul[19]), .Y(n107) );
  BUFX20 U40 ( .A(in_17bit[16]), .Y(n52) );
  AOI21X4 U41 ( .A0(n12), .A1(n53), .B0(n61), .Y(n58) );
  NAND3X2 U42 ( .A(in_17bit[1]), .B(n52), .C(in_17bit[0]), .Y(n15) );
  XOR2X4 U43 ( .A(n58), .B(n14), .Y(in_8bit_b[5]) );
  NOR3X4 U44 ( .A(in_8bit[6]), .B(n62), .C(n61), .Y(in_8bit_b[7]) );
  XNOR2X2 U45 ( .A(mul[9]), .B(n31), .Y(out[2]) );
  NAND2X2 U46 ( .A(n95), .B(n112), .Y(n31) );
  NOR2X2 U47 ( .A(mul[22]), .B(mul[21]), .Y(n118) );
  OR2X4 U48 ( .A(in_17bit[0]), .B(in_17bit[1]), .Y(n50) );
  OR2X4 U49 ( .A(mul[14]), .B(n100), .Y(n101) );
  XOR2X4 U50 ( .A(mul[10]), .B(n29), .Y(out[3]) );
  AND2X4 U51 ( .A(n96), .B(n112), .Y(n29) );
  NAND2BX4 U52 ( .AN(in_17bit[2]), .B(n64), .Y(n65) );
  INVX4 U53 ( .A(n109), .Y(n111) );
  NAND2X2 U54 ( .A(n3), .B(n67), .Y(n69) );
  NAND2X2 U55 ( .A(in_8bit[0]), .B(in_8bit[7]), .Y(n35) );
  INVX8 U56 ( .A(in_8bit[7]), .Y(n61) );
  XNOR2X2 U57 ( .A(in_8bit[1]), .B(n35), .Y(in_8bit_b[1]) );
  OR2X4 U58 ( .A(n39), .B(n92), .Y(n33) );
  AND2X4 U59 ( .A(n71), .B(n70), .Y(n39) );
  CLKINVX4 U60 ( .A(n108), .Y(n18) );
  XNOR2X4 U61 ( .A(mul[14]), .B(n24), .Y(out[7]) );
  NAND2X4 U62 ( .A(n100), .B(n112), .Y(n24) );
  INVX8 U63 ( .A(in_8bit[4]), .Y(n53) );
  XOR2X4 U64 ( .A(mul[17]), .B(n23), .Y(out[10]) );
  NOR2X2 U65 ( .A(in_17bit[0]), .B(in_17bit[1]), .Y(n64) );
  XOR2X2 U66 ( .A(mul[23]), .B(n119), .Y(out[16]) );
  NOR2X4 U67 ( .A(n1), .B(in_17bit[3]), .Y(n48) );
  XNOR2X2 U68 ( .A(mul[12]), .B(n26), .Y(out[5]) );
  NAND2X2 U69 ( .A(n98), .B(n112), .Y(n26) );
  XNOR2X4 U70 ( .A(mul[13]), .B(n28), .Y(out[6]) );
  NAND2X2 U71 ( .A(n99), .B(n112), .Y(n28) );
  OAI21X4 U72 ( .A0(in_17bit[0]), .A1(in_17bit[1]), .B0(n52), .Y(n63) );
  BUFX20 U73 ( .A(n121), .Y(out[13]) );
  NOR2X4 U74 ( .A(mul[18]), .B(n106), .Y(n37) );
  NOR2X2 U75 ( .A(n37), .B(n117), .Y(n108) );
  XOR2X4 U76 ( .A(n70), .B(n68), .Y(in_17bit_b[5]) );
  NAND2X2 U77 ( .A(n101), .B(n112), .Y(n25) );
  XNOR2X4 U78 ( .A(n17), .B(n32), .Y(in_8bit_b[2]) );
  NAND2X4 U79 ( .A(in_8bit[7]), .B(n55), .Y(n32) );
  XNOR2X4 U80 ( .A(mul[15]), .B(n25), .Y(out[8]) );
  INVX8 U81 ( .A(mul[20]), .Y(n110) );
  NAND2X2 U82 ( .A(n107), .B(n108), .Y(n20) );
  NAND2X4 U83 ( .A(n18), .B(n19), .Y(n21) );
  NAND2X4 U84 ( .A(n21), .B(n20), .Y(out[12]) );
  INVX8 U85 ( .A(n49), .Y(in_17bit_b[1]) );
  OR2X4 U86 ( .A(mul[17]), .B(n105), .Y(n106) );
  XNOR2X4 U87 ( .A(n34), .B(n76), .Y(in_17bit_b[8]) );
  NOR2XL U88 ( .A(n43), .B(n92), .Y(n34) );
  NAND2X1 U89 ( .A(n40), .B(n91), .Y(n93) );
  OR2X4 U90 ( .A(in_8bit[1]), .B(in_8bit[0]), .Y(n55) );
  NAND2X2 U91 ( .A(n52), .B(n69), .Y(n68) );
  NAND2XL U92 ( .A(n43), .B(n76), .Y(n77) );
  NAND2XL U93 ( .A(n42), .B(n81), .Y(n82) );
  NAND2XL U94 ( .A(n41), .B(n86), .Y(n87) );
  OR2X4 U95 ( .A(mul[11]), .B(n97), .Y(n98) );
  OR2X4 U96 ( .A(mul[10]), .B(n96), .Y(n97) );
  OR2X4 U97 ( .A(mul[9]), .B(n95), .Y(n96) );
  OR2X4 U98 ( .A(mul[8]), .B(out[0]), .Y(n95) );
  OR2X4 U99 ( .A(mul[16]), .B(n104), .Y(n105) );
  NAND2X4 U100 ( .A(n106), .B(n112), .Y(n27) );
  NAND2XL U101 ( .A(out[0]), .B(n112), .Y(n94) );
  NAND2XL U102 ( .A(n97), .B(n112), .Y(n30) );
  XNOR2X4 U103 ( .A(n56), .B(in_8bit[3]), .Y(in_8bit_b[3]) );
  INVX4 U104 ( .A(n117), .Y(n112) );
  XOR2X4 U105 ( .A(n33), .B(n72), .Y(in_17bit_b[6]) );
  NAND2X4 U106 ( .A(n39), .B(n72), .Y(n73) );
  AND2X4 U107 ( .A(n75), .B(n74), .Y(n43) );
  AND2X4 U108 ( .A(n79), .B(n78), .Y(n42) );
  AND2X4 U109 ( .A(n89), .B(n88), .Y(n40) );
  AND2X4 U110 ( .A(n84), .B(n83), .Y(n41) );
  XNOR2X4 U111 ( .A(in_17bit[3]), .B(n36), .Y(in_17bit_b[3]) );
  INVX4 U112 ( .A(in_17bit[4]), .Y(n67) );
  OR2X4 U113 ( .A(mul[13]), .B(n99), .Y(n100) );
  XOR2X4 U114 ( .A(n38), .B(n110), .Y(n121) );
  NOR2XL U115 ( .A(n40), .B(n92), .Y(n90) );
  NOR2XL U116 ( .A(n41), .B(n92), .Y(n85) );
  NOR2XL U117 ( .A(n42), .B(n92), .Y(n80) );
  XNOR2X2 U118 ( .A(n88), .B(n44), .Y(in_17bit_b[13]) );
  AND2X1 U119 ( .A(n52), .B(n87), .Y(n44) );
  XNOR2X2 U120 ( .A(n83), .B(n45), .Y(in_17bit_b[11]) );
  AND2X1 U121 ( .A(n52), .B(n82), .Y(n45) );
  XNOR2X2 U122 ( .A(n78), .B(n46), .Y(in_17bit_b[9]) );
  AND2X1 U123 ( .A(n52), .B(n77), .Y(n46) );
  AND2X1 U124 ( .A(n52), .B(n73), .Y(n47) );
  XNOR2X4 U125 ( .A(n63), .B(in_17bit[2]), .Y(in_17bit_b[2]) );
  XOR2X2 U126 ( .A(in_17bit[15]), .B(n51), .Y(in_17bit_b[15]) );
  AND2X1 U127 ( .A(n52), .B(n93), .Y(n51) );
  INVX1 U128 ( .A(in_17bit[5]), .Y(n70) );
  NOR4X4 U129 ( .A(in_8bit[2]), .B(in_8bit[1]), .C(in_8bit[0]), .D(in_8bit[3]), 
        .Y(n59) );
  XNOR2X4 U130 ( .A(n57), .B(n53), .Y(in_8bit_b[4]) );
  NAND2X4 U131 ( .A(n62), .B(in_8bit[7]), .Y(n60) );
  NOR2X4 U132 ( .A(n48), .B(n92), .Y(n66) );
  XNOR2X4 U133 ( .A(n66), .B(n67), .Y(in_17bit_b[4]) );
  CLKINVX3 U134 ( .A(n69), .Y(n71) );
  CLKINVX3 U135 ( .A(in_17bit[6]), .Y(n72) );
  CLKINVX3 U136 ( .A(in_17bit[7]), .Y(n74) );
  CLKINVX3 U137 ( .A(n73), .Y(n75) );
  CLKINVX3 U138 ( .A(in_17bit[8]), .Y(n76) );
  CLKINVX3 U139 ( .A(in_17bit[9]), .Y(n78) );
  CLKINVX3 U140 ( .A(n77), .Y(n79) );
  CLKINVX3 U141 ( .A(in_17bit[10]), .Y(n81) );
  XNOR2X4 U142 ( .A(n80), .B(n81), .Y(in_17bit_b[10]) );
  CLKINVX3 U143 ( .A(in_17bit[11]), .Y(n83) );
  CLKINVX3 U144 ( .A(n82), .Y(n84) );
  CLKINVX3 U145 ( .A(in_17bit[12]), .Y(n86) );
  XNOR2X4 U146 ( .A(n85), .B(n86), .Y(in_17bit_b[12]) );
  CLKINVX3 U147 ( .A(in_17bit[13]), .Y(n88) );
  CLKINVX3 U148 ( .A(in_17bit[14]), .Y(n91) );
  XNOR2X4 U149 ( .A(n90), .B(n91), .Y(in_17bit_b[14]) );
  NOR3X4 U150 ( .A(in_17bit[15]), .B(n93), .C(n92), .Y(in_17bit_b[16]) );
  CLKINVX3 U151 ( .A(n101), .Y(n102) );
  NAND2BX4 U152 ( .AN(mul[15]), .B(n102), .Y(n104) );
  NAND2X4 U153 ( .A(n104), .B(n112), .Y(n103) );
  XNOR2X4 U154 ( .A(mul[16]), .B(n103), .Y(out[9]) );
  NAND2X4 U155 ( .A(n111), .B(n110), .Y(n114) );
  NAND2X4 U156 ( .A(n114), .B(n112), .Y(n113) );
  XOR2X4 U157 ( .A(n113), .B(n115), .Y(out[14]) );
  AOI21X4 U158 ( .A0(n2), .A1(n115), .B0(n117), .Y(n116) );
  XOR2X4 U159 ( .A(n116), .B(mul[22]), .Y(out[15]) );
endmodule


module multi16_6_DW01_add_0 ( A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, 
        A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, 
        B_20_, B_19_, B_18_, B_17_, B_16_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, 
        SUM_17_, SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, 
        SUM_9_, SUM_8_, SUM_7_, SUM_6_, SUM_5_ );
  input A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_,
         A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, B_20_, B_19_,
         B_18_, B_17_, B_16_;
  output SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, SUM_15_,
         SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, SUM_7_,
         SUM_6_, SUM_5_;
  wire   n1, n2, n3, n4, n5, n6, n7, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44;

  INVX4 U2 ( .A(n34), .Y(n19) );
  INVX2 U3 ( .A(n36), .Y(n20) );
  NOR2X2 U4 ( .A(n30), .B(n31), .Y(n4) );
  OAI21X4 U5 ( .A0(n41), .A1(n34), .B0(n36), .Y(n39) );
  BUFX4 U6 ( .A(n21), .Y(n3) );
  BUFX12 U7 ( .A(A_12_), .Y(SUM_12_) );
  CLKINVX3 U8 ( .A(n21), .Y(n1) );
  INVX4 U9 ( .A(n33), .Y(n22) );
  NAND2X2 U10 ( .A(B_18_), .B(A_18_), .Y(n36) );
  AOI21X4 U11 ( .A0(n23), .A1(n22), .B0(n3), .Y(n2) );
  INVX8 U12 ( .A(n38), .Y(n21) );
  INVX8 U13 ( .A(n37), .Y(n23) );
  BUFX12 U14 ( .A(A_14_), .Y(SUM_14_) );
  XOR2X4 U15 ( .A(n27), .B(n7), .Y(SUM_20_) );
  NOR2BX4 U16 ( .AN(n32), .B(n31), .Y(n40) );
  OAI21X1 U17 ( .A0(n37), .A1(n33), .B0(n1), .Y(n35) );
  AOI21X4 U18 ( .A0(n23), .A1(n22), .B0(n3), .Y(n41) );
  XOR2X4 U19 ( .A(n39), .B(n40), .Y(SUM_19_) );
  OR2X4 U20 ( .A(B_20_), .B(A_20_), .Y(n28) );
  NOR2X4 U21 ( .A(B_18_), .B(A_18_), .Y(n34) );
  NAND2X4 U22 ( .A(n36), .B(n19), .Y(n42) );
  BUFX8 U23 ( .A(A_6_), .Y(SUM_6_) );
  CLKINVX8 U24 ( .A(A_15_), .Y(n24) );
  NOR2X4 U25 ( .A(A_17_), .B(B_17_), .Y(n33) );
  NAND2X2 U26 ( .A(B_19_), .B(A_19_), .Y(n32) );
  NOR2X4 U27 ( .A(B_19_), .B(A_19_), .Y(n31) );
  BUFX12 U28 ( .A(A_10_), .Y(SUM_10_) );
  INVX8 U29 ( .A(n24), .Y(SUM_15_) );
  INVXL U30 ( .A(n32), .Y(n5) );
  OR2X4 U31 ( .A(n4), .B(n5), .Y(n27) );
  AOI21X2 U32 ( .A0(n19), .A1(n35), .B0(n20), .Y(n30) );
  AOI21X2 U33 ( .A0(n27), .A1(n28), .B0(n18), .Y(n26) );
  XOR2X4 U34 ( .A(n6), .B(n23), .Y(SUM_17_) );
  NOR2X4 U35 ( .A(n21), .B(n33), .Y(n6) );
  AND2X2 U36 ( .A(n29), .B(n28), .Y(n7) );
  INVXL U37 ( .A(n29), .Y(n18) );
  BUFX4 U38 ( .A(A_9_), .Y(SUM_9_) );
  BUFX8 U39 ( .A(A_11_), .Y(SUM_11_) );
  BUFX8 U40 ( .A(A_5_), .Y(SUM_5_) );
  BUFX4 U41 ( .A(A_8_), .Y(SUM_8_) );
  BUFX4 U42 ( .A(A_7_), .Y(SUM_7_) );
  BUFX8 U43 ( .A(A_13_), .Y(SUM_13_) );
  INVX8 U44 ( .A(n44), .Y(SUM_16_) );
  NAND2X4 U45 ( .A(n43), .B(n37), .Y(n44) );
  OR2X4 U46 ( .A(A_16_), .B(B_16_), .Y(n43) );
  NAND2X4 U47 ( .A(B_16_), .B(A_16_), .Y(n37) );
  NAND2X4 U48 ( .A(A_17_), .B(B_17_), .Y(n38) );
  XOR2X4 U49 ( .A(n2), .B(n42), .Y(SUM_18_) );
  XOR2X1 U50 ( .A(n25), .B(n26), .Y(SUM_21_) );
  XNOR2X1 U51 ( .A(B_21_), .B(A_21_), .Y(n25) );
  NAND2X1 U52 ( .A(B_20_), .B(A_20_), .Y(n29) );
endmodule


module multi16_6_DW02_mult_0 ( A, B, PRODUCT_23_, PRODUCT_22_, PRODUCT_21_, 
        PRODUCT_20_, PRODUCT_19_, PRODUCT_18_, PRODUCT_17_, PRODUCT_16_, 
        PRODUCT_15_, PRODUCT_14_, PRODUCT_13_, PRODUCT_12_, PRODUCT_11_, 
        PRODUCT_10_, PRODUCT_9_, PRODUCT_8_, PRODUCT_7_ );
  input [16:0] A;
  input [7:0] B;
  output PRODUCT_23_, PRODUCT_22_, PRODUCT_21_, PRODUCT_20_, PRODUCT_19_,
         PRODUCT_18_, PRODUCT_17_, PRODUCT_16_, PRODUCT_15_, PRODUCT_14_,
         PRODUCT_13_, PRODUCT_12_, PRODUCT_11_, PRODUCT_10_, PRODUCT_9_,
         PRODUCT_8_, PRODUCT_7_;
  wire   n47, ab_16__7_, ab_16__6_, ab_16__5_, ab_16__4_, ab_16__3_, ab_16__2_,
         ab_16__1_, ab_16__0_, ab_15__7_, ab_15__6_, ab_15__5_, ab_15__4_,
         ab_15__3_, ab_15__2_, ab_15__1_, ab_15__0_, ab_14__7_, ab_14__6_,
         ab_14__5_, ab_14__4_, ab_14__3_, ab_14__2_, ab_14__1_, ab_14__0_,
         ab_13__7_, ab_13__6_, ab_13__5_, ab_13__4_, ab_13__3_, ab_13__2_,
         ab_13__1_, ab_13__0_, ab_12__7_, ab_12__6_, ab_12__5_, ab_12__4_,
         ab_12__3_, ab_12__2_, ab_12__1_, ab_12__0_, ab_11__7_, ab_11__6_,
         ab_11__5_, ab_11__4_, ab_11__3_, ab_11__2_, ab_11__1_, ab_11__0_,
         ab_10__7_, ab_10__6_, ab_10__5_, ab_10__4_, ab_10__3_, ab_10__2_,
         ab_10__1_, ab_10__0_, ab_9__7_, ab_9__6_, ab_9__5_, ab_9__4_,
         ab_9__3_, ab_9__2_, ab_9__1_, ab_9__0_, ab_8__7_, ab_8__6_, ab_8__5_,
         ab_8__4_, ab_8__3_, ab_8__2_, ab_8__1_, ab_8__0_, ab_7__7_, ab_7__6_,
         ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_, ab_7__0_, ab_6__7_,
         ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_, ab_6__1_, ab_6__0_,
         ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_, ab_5__2_, ab_5__1_,
         ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_, ab_4__3_, ab_4__2_,
         ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_, ab_3__4_, ab_3__3_,
         ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_, ab_2__5_, ab_2__4_,
         ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_, ab_1__6_, ab_1__5_,
         ab_1__4_, ab_1__3_, ab_1__2_, ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_,
         ab_0__3_, ab_0__2_, CARRYB_16__6_, CARRYB_16__5_, CARRYB_16__4_,
         CARRYB_16__3_, CARRYB_16__2_, CARRYB_16__1_, CARRYB_16__0_,
         CARRYB_15__6_, CARRYB_15__5_, CARRYB_15__4_, CARRYB_15__3_,
         CARRYB_15__2_, CARRYB_15__1_, CARRYB_15__0_, CARRYB_14__6_,
         CARRYB_14__5_, CARRYB_14__4_, CARRYB_14__3_, CARRYB_14__2_,
         CARRYB_14__1_, CARRYB_14__0_, CARRYB_13__6_, CARRYB_13__5_,
         CARRYB_13__4_, CARRYB_13__3_, CARRYB_13__2_, CARRYB_13__1_,
         CARRYB_13__0_, CARRYB_12__6_, CARRYB_12__5_, CARRYB_12__4_,
         CARRYB_12__3_, CARRYB_12__2_, CARRYB_12__1_, CARRYB_12__0_,
         CARRYB_11__6_, CARRYB_11__5_, CARRYB_11__4_, CARRYB_11__3_,
         CARRYB_11__2_, CARRYB_11__1_, CARRYB_11__0_, CARRYB_10__6_,
         CARRYB_10__5_, CARRYB_10__4_, CARRYB_10__3_, CARRYB_10__2_,
         CARRYB_10__1_, CARRYB_10__0_, CARRYB_9__6_, CARRYB_9__5_,
         CARRYB_9__4_, CARRYB_9__3_, CARRYB_9__2_, CARRYB_9__1_, CARRYB_9__0_,
         CARRYB_8__6_, CARRYB_8__5_, CARRYB_8__4_, CARRYB_8__3_, CARRYB_8__2_,
         CARRYB_8__1_, CARRYB_8__0_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_,
         CARRYB_7__3_, CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_,
         CARRYB_6__5_, CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_,
         CARRYB_6__0_, CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_,
         CARRYB_5__2_, CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_,
         CARRYB_4__4_, CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_,
         CARRYB_3__6_, CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_,
         CARRYB_3__1_, CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_,
         CARRYB_2__3_, CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__0_,
         SUMB_16__6_, SUMB_16__5_, SUMB_16__4_, SUMB_16__3_, SUMB_16__2_,
         SUMB_16__1_, SUMB_16__0_, SUMB_15__6_, SUMB_15__5_, SUMB_15__4_,
         SUMB_15__3_, SUMB_15__2_, SUMB_15__1_, SUMB_14__6_, SUMB_14__5_,
         SUMB_14__4_, SUMB_14__3_, SUMB_14__2_, SUMB_14__1_, SUMB_13__6_,
         SUMB_13__5_, SUMB_13__4_, SUMB_13__3_, SUMB_13__2_, SUMB_13__1_,
         SUMB_12__6_, SUMB_12__5_, SUMB_12__4_, SUMB_12__3_, SUMB_12__2_,
         SUMB_12__1_, SUMB_11__6_, SUMB_11__5_, SUMB_11__4_, SUMB_11__3_,
         SUMB_11__2_, SUMB_11__1_, SUMB_10__6_, SUMB_10__5_, SUMB_10__4_,
         SUMB_10__3_, SUMB_10__2_, SUMB_10__1_, SUMB_9__6_, SUMB_9__5_,
         SUMB_9__4_, SUMB_9__3_, SUMB_9__2_, SUMB_9__1_, SUMB_8__6_,
         SUMB_8__5_, SUMB_8__4_, SUMB_8__3_, SUMB_8__2_, SUMB_8__1_,
         SUMB_7__6_, SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_,
         SUMB_7__1_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, PROD1_7_, A1_21_, A1_20_, A1_19_, A1_18_,
         A1_17_, A1_16_, A1_15_, A1_13_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_,
         A1_7_, A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, n3, n4, n5, n6, n8,
         n9, n10, n11, n12, n13, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44;

  ADDFHX2 S3_13_6 ( .A(ab_13__6_), .B(CARRYB_12__6_), .CI(ab_12__7_), .CO(
        CARRYB_13__6_), .S(SUMB_13__6_) );
  multi16_6_DW01_add_0 FS_1 ( .A_21_(A1_21_), .A_20_(A1_20_), .A_19_(A1_19_), 
        .A_18_(A1_18_), .A_17_(A1_17_), .A_16_(A1_16_), .A_15_(A1_15_), 
        .A_14_(SUMB_16__0_), .A_13_(A1_13_), .A_12_(A1_12_), .A_11_(A1_11_), 
        .A_10_(A1_10_), .A_9_(A1_9_), .A_8_(A1_8_), .A_7_(A1_7_), .A_6_(A1_6_), 
        .A_5_(PROD1_7_), .B_21_(n23), .B_20_(n22), .B_19_(n21), .B_18_(n19), 
        .B_17_(n8), .B_16_(n20), .SUM_21_(PRODUCT_23_), .SUM_20_(PRODUCT_22_), 
        .SUM_19_(PRODUCT_21_), .SUM_18_(n47), .SUM_17_(PRODUCT_19_), .SUM_16_(
        PRODUCT_18_), .SUM_15_(PRODUCT_17_), .SUM_14_(PRODUCT_16_), .SUM_13_(
        PRODUCT_15_), .SUM_12_(PRODUCT_14_), .SUM_11_(PRODUCT_13_), .SUM_10_(
        PRODUCT_12_), .SUM_9_(PRODUCT_11_), .SUM_8_(PRODUCT_10_), .SUM_7_(
        PRODUCT_9_), .SUM_6_(PRODUCT_8_), .SUM_5_(PRODUCT_7_) );
  ADDFHX4 S2_9_2 ( .A(ab_9__2_), .B(CARRYB_8__2_), .CI(SUMB_8__3_), .CO(
        CARRYB_9__2_), .S(SUMB_9__2_) );
  ADDFHX4 S2_9_1 ( .A(ab_9__1_), .B(CARRYB_8__1_), .CI(SUMB_8__2_), .CO(
        CARRYB_9__1_), .S(SUMB_9__1_) );
  ADDFHX4 S4_2 ( .A(ab_16__2_), .B(CARRYB_15__2_), .CI(SUMB_15__3_), .CO(
        CARRYB_16__2_), .S(SUMB_16__2_) );
  ADDFHX4 S2_13_4 ( .A(ab_13__4_), .B(CARRYB_12__4_), .CI(SUMB_12__5_), .CO(
        CARRYB_13__4_), .S(SUMB_13__4_) );
  ADDFHX4 S2_12_5 ( .A(ab_12__5_), .B(CARRYB_11__5_), .CI(SUMB_11__6_), .CO(
        CARRYB_12__5_), .S(SUMB_12__5_) );
  ADDFHX4 S2_14_1 ( .A(ab_14__1_), .B(CARRYB_13__1_), .CI(SUMB_13__2_), .CO(
        CARRYB_14__1_), .S(SUMB_14__1_) );
  ADDFHX4 S2_11_3 ( .A(ab_11__3_), .B(CARRYB_10__3_), .CI(SUMB_10__4_), .CO(
        CARRYB_11__3_), .S(SUMB_11__3_) );
  ADDFHX4 S2_12_2 ( .A(ab_12__2_), .B(CARRYB_11__2_), .CI(SUMB_11__3_), .CO(
        CARRYB_12__2_), .S(SUMB_12__2_) );
  ADDFHX4 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  ADDFHX4 S1_15_0 ( .A(ab_15__0_), .B(CARRYB_14__0_), .CI(SUMB_14__1_), .CO(
        CARRYB_15__0_), .S(A1_13_) );
  ADDFHX4 S1_13_0 ( .A(ab_13__0_), .B(CARRYB_12__0_), .CI(SUMB_12__1_), .CO(
        CARRYB_13__0_), .S(A1_11_) );
  ADDFHX4 S1_14_0 ( .A(ab_14__0_), .B(CARRYB_13__0_), .CI(SUMB_13__1_), .CO(
        CARRYB_14__0_), .S(A1_12_) );
  ADDFHX4 S2_15_2 ( .A(ab_15__2_), .B(CARRYB_14__2_), .CI(SUMB_14__3_), .CO(
        CARRYB_15__2_), .S(SUMB_15__2_) );
  ADDFHX4 S2_10_3 ( .A(ab_10__3_), .B(CARRYB_9__3_), .CI(SUMB_9__4_), .CO(
        CARRYB_10__3_), .S(SUMB_10__3_) );
  ADDFHX4 S3_10_6 ( .A(ab_10__6_), .B(CARRYB_9__6_), .CI(ab_9__7_), .CO(
        CARRYB_10__6_), .S(SUMB_10__6_) );
  ADDFHX4 S3_11_6 ( .A(ab_11__6_), .B(CARRYB_10__6_), .CI(ab_10__7_), .CO(
        CARRYB_11__6_), .S(SUMB_11__6_) );
  ADDFHX4 S2_11_4 ( .A(ab_11__4_), .B(CARRYB_10__4_), .CI(SUMB_10__5_), .CO(
        CARRYB_11__4_), .S(SUMB_11__4_) );
  ADDFHX4 S2_12_4 ( .A(ab_12__4_), .B(CARRYB_11__4_), .CI(SUMB_11__5_), .CO(
        CARRYB_12__4_), .S(SUMB_12__4_) );
  ADDFHX4 S2_12_3 ( .A(ab_12__3_), .B(CARRYB_11__3_), .CI(SUMB_11__4_), .CO(
        CARRYB_12__3_), .S(SUMB_12__3_) );
  ADDFHX4 S2_13_2 ( .A(ab_13__2_), .B(CARRYB_12__2_), .CI(SUMB_12__3_), .CO(
        CARRYB_13__2_), .S(SUMB_13__2_) );
  ADDFHX4 S2_10_2 ( .A(ab_10__2_), .B(CARRYB_9__2_), .CI(SUMB_9__3_), .CO(
        CARRYB_10__2_), .S(SUMB_10__2_) );
  ADDFHX4 S2_15_1 ( .A(ab_15__1_), .B(CARRYB_14__1_), .CI(SUMB_14__2_), .CO(
        CARRYB_15__1_), .S(SUMB_15__1_) );
  ADDFHX4 S4_1 ( .A(ab_16__1_), .B(CARRYB_15__1_), .CI(SUMB_15__2_), .CO(
        CARRYB_16__1_), .S(SUMB_16__1_) );
  ADDFHX4 S2_12_1 ( .A(ab_12__1_), .B(CARRYB_11__1_), .CI(SUMB_11__2_), .CO(
        CARRYB_12__1_), .S(SUMB_12__1_) );
  ADDFHX4 S2_13_1 ( .A(ab_13__1_), .B(CARRYB_12__1_), .CI(SUMB_12__2_), .CO(
        CARRYB_13__1_), .S(SUMB_13__1_) );
  ADDFX2 S3_15_6 ( .A(ab_15__6_), .B(CARRYB_14__6_), .CI(ab_14__7_), .CO(
        CARRYB_15__6_), .S(SUMB_15__6_) );
  ADDFHX4 S2_2_4 ( .A(ab_2__4_), .B(n13), .CI(SUMB_1__5_), .CO(CARRYB_2__4_), 
        .S(SUMB_2__4_) );
  ADDFHX4 S2_8_4 ( .A(ab_8__4_), .B(CARRYB_7__4_), .CI(SUMB_7__5_), .CO(
        CARRYB_8__4_), .S(SUMB_8__4_) );
  ADDFHX4 S2_8_2 ( .A(ab_8__2_), .B(CARRYB_7__2_), .CI(SUMB_7__3_), .CO(
        CARRYB_8__2_), .S(SUMB_8__2_) );
  ADDFHX4 S2_14_2 ( .A(ab_14__2_), .B(CARRYB_13__2_), .CI(SUMB_13__3_), .CO(
        CARRYB_14__2_), .S(SUMB_14__2_) );
  ADDFHX4 S4_5 ( .A(ab_16__5_), .B(CARRYB_15__5_), .CI(SUMB_15__6_), .CO(
        CARRYB_16__5_), .S(SUMB_16__5_) );
  ADDFHX4 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  ADDFHX4 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  ADDFHX4 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  ADDFHX4 S1_10_0 ( .A(ab_10__0_), .B(CARRYB_9__0_), .CI(SUMB_9__1_), .CO(
        CARRYB_10__0_), .S(A1_8_) );
  ADDFHX4 S4_3 ( .A(ab_16__3_), .B(CARRYB_15__3_), .CI(SUMB_15__4_), .CO(
        CARRYB_16__3_), .S(SUMB_16__3_) );
  ADDFHX4 S2_10_1 ( .A(ab_10__1_), .B(CARRYB_9__1_), .CI(SUMB_9__2_), .CO(
        CARRYB_10__1_), .S(SUMB_10__1_) );
  ADDFHX4 S2_11_1 ( .A(ab_11__1_), .B(CARRYB_10__1_), .CI(SUMB_10__2_), .CO(
        CARRYB_11__1_), .S(SUMB_11__1_) );
  ADDFHX4 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  ADDFHX4 S2_9_3 ( .A(ab_9__3_), .B(CARRYB_8__3_), .CI(SUMB_8__4_), .CO(
        CARRYB_9__3_), .S(SUMB_9__3_) );
  ADDFHX4 S2_7_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  ADDFHX4 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  ADDFHX4 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  ADDFHX4 S2_7_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  ADDFHX4 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  ADDFHX4 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  ADDFHX4 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  ADDFHX4 S2_11_5 ( .A(ab_11__5_), .B(CARRYB_10__5_), .CI(SUMB_10__6_), .CO(
        CARRYB_11__5_), .S(SUMB_11__5_) );
  ADDFHX4 S1_11_0 ( .A(ab_11__0_), .B(CARRYB_10__0_), .CI(SUMB_10__1_), .CO(
        CARRYB_11__0_), .S(A1_9_) );
  ADDFHX4 S1_12_0 ( .A(ab_12__0_), .B(CARRYB_11__0_), .CI(SUMB_11__1_), .CO(
        CARRYB_12__0_), .S(A1_10_) );
  ADDFHX4 S1_8_0 ( .A(ab_8__0_), .B(CARRYB_7__0_), .CI(SUMB_7__1_), .CO(
        CARRYB_8__0_), .S(A1_6_) );
  ADDFHX4 S1_9_0 ( .A(ab_9__0_), .B(CARRYB_8__0_), .CI(SUMB_8__1_), .CO(
        CARRYB_9__0_), .S(A1_7_) );
  ADDFHX4 S3_9_6 ( .A(ab_9__6_), .B(CARRYB_8__6_), .CI(ab_8__7_), .CO(
        CARRYB_9__6_), .S(SUMB_9__6_) );
  ADDFHX4 S3_8_6 ( .A(ab_8__6_), .B(CARRYB_7__6_), .CI(ab_7__7_), .CO(
        CARRYB_8__6_), .S(SUMB_8__6_) );
  ADDFHX4 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  ADDFHX4 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  ADDFHX4 S2_10_5 ( .A(ab_10__5_), .B(CARRYB_9__5_), .CI(SUMB_9__6_), .CO(
        CARRYB_10__5_), .S(SUMB_10__5_) );
  ADDFHX4 S2_8_5 ( .A(ab_8__5_), .B(CARRYB_7__5_), .CI(SUMB_7__6_), .CO(
        CARRYB_8__5_), .S(SUMB_8__5_) );
  ADDFHX4 S2_9_5 ( .A(ab_9__5_), .B(CARRYB_8__5_), .CI(SUMB_8__6_), .CO(
        CARRYB_9__5_), .S(SUMB_9__5_) );
  ADDFHX4 S2_7_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  ADDFHX4 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  ADDFHX4 S2_2_3 ( .A(ab_2__3_), .B(n10), .CI(SUMB_1__4_), .CO(CARRYB_2__3_), 
        .S(SUMB_2__3_) );
  ADDFHX4 S2_2_2 ( .A(ab_2__2_), .B(n12), .CI(SUMB_1__3_), .CO(CARRYB_2__2_), 
        .S(SUMB_2__2_) );
  ADDFHX4 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  ADDFHX4 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  ADDFHX4 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  ADDFHX4 S1_7_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(PROD1_7_) );
  ADDFHX4 S2_8_3 ( .A(ab_8__3_), .B(CARRYB_7__3_), .CI(SUMB_7__4_), .CO(
        CARRYB_8__3_), .S(SUMB_8__3_) );
  ADDFHX4 S2_14_3 ( .A(ab_14__3_), .B(CARRYB_13__3_), .CI(SUMB_13__4_), .CO(
        CARRYB_14__3_), .S(SUMB_14__3_) );
  ADDFHX4 S2_14_4 ( .A(ab_14__4_), .B(CARRYB_13__4_), .CI(SUMB_13__5_), .CO(
        CARRYB_14__4_), .S(SUMB_14__4_) );
  ADDFHX4 S2_10_4 ( .A(ab_10__4_), .B(CARRYB_9__4_), .CI(SUMB_9__5_), .CO(
        CARRYB_10__4_), .S(SUMB_10__4_) );
  ADDFHX4 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  ADDFHX4 S2_13_3 ( .A(ab_13__3_), .B(CARRYB_12__3_), .CI(SUMB_12__4_), .CO(
        CARRYB_13__3_), .S(SUMB_13__3_) );
  ADDFHX4 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  ADDFHX4 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  ADDFHX4 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  ADDFHX4 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  ADDFHX4 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  ADDFHX4 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  ADDFHX4 S2_2_5 ( .A(ab_2__5_), .B(n16), .CI(SUMB_1__6_), .CO(CARRYB_2__5_), 
        .S(SUMB_2__5_) );
  ADDFHX4 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  ADDFHX4 S2_2_1 ( .A(ab_2__1_), .B(n9), .CI(SUMB_1__2_), .CO(CARRYB_2__1_), 
        .S(SUMB_2__1_) );
  ADDFHX4 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  ADDFHX4 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  ADDFHX4 S3_2_6 ( .A(ab_2__6_), .B(n11), .CI(ab_1__7_), .CO(CARRYB_2__6_), 
        .S(SUMB_2__6_) );
  ADDFHX4 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  ADDFHX4 S2_7_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  ADDFHX4 S3_7_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(
        CARRYB_7__6_), .S(SUMB_7__6_) );
  ADDFHX4 S4_4 ( .A(ab_16__4_), .B(CARRYB_15__4_), .CI(SUMB_15__5_), .CO(
        CARRYB_16__4_), .S(SUMB_16__4_) );
  ADDFHX4 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  ADDFHX4 S2_11_2 ( .A(ab_11__2_), .B(CARRYB_10__2_), .CI(SUMB_10__3_), .CO(
        CARRYB_11__2_), .S(SUMB_11__2_) );
  ADDFHX4 S2_7_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  ADDFHX4 S2_8_1 ( .A(ab_8__1_), .B(CARRYB_7__1_), .CI(SUMB_7__2_), .CO(
        CARRYB_8__1_), .S(SUMB_8__1_) );
  ADDFHX4 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  ADDFHX4 S4_0 ( .A(ab_16__0_), .B(CARRYB_15__0_), .CI(SUMB_15__1_), .CO(
        CARRYB_16__0_), .S(SUMB_16__0_) );
  ADDFHX4 S2_13_5 ( .A(ab_13__5_), .B(CARRYB_12__5_), .CI(SUMB_12__6_), .CO(
        CARRYB_13__5_), .S(SUMB_13__5_) );
  ADDFHX4 S5_6 ( .A(ab_16__6_), .B(CARRYB_15__6_), .CI(ab_15__7_), .CO(
        CARRYB_16__6_), .S(SUMB_16__6_) );
  ADDFHX4 S2_15_3 ( .A(ab_15__3_), .B(CARRYB_14__3_), .CI(SUMB_14__4_), .CO(
        CARRYB_15__3_), .S(SUMB_15__3_) );
  ADDFHX4 S2_9_4 ( .A(ab_9__4_), .B(CARRYB_8__4_), .CI(SUMB_8__5_), .CO(
        CARRYB_9__4_), .S(SUMB_9__4_) );
  ADDFHX4 S3_12_6 ( .A(ab_12__6_), .B(CARRYB_11__6_), .CI(ab_11__7_), .CO(
        CARRYB_12__6_), .S(SUMB_12__6_) );
  ADDFHX2 S3_14_6 ( .A(ab_14__6_), .B(CARRYB_13__6_), .CI(ab_13__7_), .CO(
        CARRYB_14__6_), .S(SUMB_14__6_) );
  ADDFHX4 S2_15_4 ( .A(ab_15__4_), .B(CARRYB_14__4_), .CI(SUMB_14__5_), .CO(
        CARRYB_15__4_), .S(SUMB_15__4_) );
  ADDFHX4 S2_15_5 ( .A(ab_15__5_), .B(CARRYB_14__5_), .CI(SUMB_14__6_), .CO(
        CARRYB_15__5_), .S(SUMB_15__5_) );
  ADDFHX4 S2_14_5 ( .A(ab_14__5_), .B(CARRYB_13__5_), .CI(SUMB_13__6_), .CO(
        CARRYB_14__5_), .S(SUMB_14__5_) );
  BUFX8 U2 ( .A(ab_0__6_), .Y(n3) );
  BUFX20 U3 ( .A(A[1]), .Y(n18) );
  CLKINVX3 U4 ( .A(n18), .Y(n4) );
  INVX4 U5 ( .A(n4), .Y(n5) );
  NAND2BX2 U6 ( .AN(n38), .B(A[0]), .Y(n6) );
  CLKINVX20 U7 ( .A(n6), .Y(ab_0__4_) );
  INVX8 U8 ( .A(B[4]), .Y(n38) );
  NOR2BX4 U9 ( .AN(A[3]), .B(n29), .Y(ab_3__2_) );
  NOR2BX4 U10 ( .AN(A[3]), .B(n31), .Y(ab_3__1_) );
  NOR2BX4 U11 ( .AN(A[3]), .B(n27), .Y(ab_3__3_) );
  NOR2BX4 U12 ( .AN(A[3]), .B(n38), .Y(ab_3__4_) );
  NOR2BX4 U13 ( .AN(A[3]), .B(n37), .Y(ab_3__5_) );
  XOR2X4 U14 ( .A(n44), .B(ab_0__2_), .Y(SUMB_1__1_) );
  NOR2BX1 U15 ( .AN(A[8]), .B(n38), .Y(ab_8__4_) );
  NOR2BXL U16 ( .AN(A[9]), .B(n25), .Y(ab_9__5_) );
  NOR2BX1 U17 ( .AN(A[9]), .B(n26), .Y(ab_9__4_) );
  NOR2BX2 U18 ( .AN(A[9]), .B(n28), .Y(ab_9__3_) );
  NOR2BX1 U19 ( .AN(A[5]), .B(n24), .Y(ab_5__6_) );
  NOR2BX2 U20 ( .AN(A[12]), .B(n28), .Y(ab_12__3_) );
  NOR2BX2 U21 ( .AN(A[8]), .B(n27), .Y(ab_8__3_) );
  NOR2BX1 U22 ( .AN(A[12]), .B(n30), .Y(ab_12__2_) );
  NOR2BX2 U23 ( .AN(A[8]), .B(n31), .Y(ab_8__1_) );
  NOR2BX1 U24 ( .AN(A[6]), .B(n24), .Y(ab_6__6_) );
  NOR2BX1 U25 ( .AN(A[14]), .B(n30), .Y(ab_14__2_) );
  NOR2BX1 U26 ( .AN(A[10]), .B(n32), .Y(ab_10__1_) );
  NOR2BX1 U27 ( .AN(A[16]), .B(n28), .Y(ab_16__3_) );
  NOR2BX1 U28 ( .AN(A[7]), .B(n38), .Y(ab_7__4_) );
  NOR2BX1 U29 ( .AN(A[11]), .B(n30), .Y(ab_11__2_) );
  NOR2BX1 U30 ( .AN(A[7]), .B(n36), .Y(ab_7__6_) );
  NOR2BX2 U31 ( .AN(A[14]), .B(n28), .Y(ab_14__3_) );
  INVX1 U32 ( .A(n29), .Y(n15) );
  BUFX16 U33 ( .A(A[2]), .Y(n17) );
  CLKINVX4 U34 ( .A(B[2]), .Y(n40) );
  NOR2BX2 U35 ( .AN(A[7]), .B(n31), .Y(ab_7__1_) );
  NOR2BX1 U36 ( .AN(A[15]), .B(n32), .Y(ab_15__1_) );
  INVX4 U37 ( .A(B[1]), .Y(n41) );
  CLKBUFX8 U38 ( .A(n42), .Y(n33) );
  AND2X4 U40 ( .A(CARRYB_16__1_), .B(SUMB_16__2_), .Y(n8) );
  BUFX3 U41 ( .A(n38), .Y(n26) );
  AND2X4 U42 ( .A(n44), .B(ab_0__2_), .Y(n9) );
  AND2X4 U43 ( .A(ab_0__4_), .B(ab_1__3_), .Y(n10) );
  AND2X4 U44 ( .A(ab_0__7_), .B(ab_1__6_), .Y(n11) );
  AND2X4 U45 ( .A(ab_1__2_), .B(ab_0__3_), .Y(n12) );
  AND2X4 U46 ( .A(ab_0__5_), .B(ab_1__4_), .Y(n13) );
  INVX4 U47 ( .A(B[6]), .Y(n36) );
  CLKBUFX2 U48 ( .A(n36), .Y(n24) );
  BUFX1 U49 ( .A(n37), .Y(n25) );
  INVX4 U50 ( .A(B[3]), .Y(n39) );
  NOR2BX2 U51 ( .AN(A[5]), .B(n29), .Y(ab_5__2_) );
  NOR2BX2 U52 ( .AN(A[4]), .B(n33), .Y(ab_4__0_) );
  XOR2X4 U53 ( .A(ab_1__2_), .B(ab_0__3_), .Y(SUMB_1__2_) );
  BUFX12 U54 ( .A(n47), .Y(PRODUCT_20_) );
  XOR2X4 U55 ( .A(ab_1__3_), .B(ab_0__4_), .Y(SUMB_1__3_) );
  NOR2BX2 U56 ( .AN(B[2]), .B(n34), .Y(ab_0__2_) );
  AND2X4 U57 ( .A(n17), .B(n15), .Y(ab_2__2_) );
  NOR2BX4 U58 ( .AN(n17), .B(n33), .Y(ab_2__0_) );
  NOR2BX4 U59 ( .AN(n17), .B(n37), .Y(ab_2__5_) );
  NOR2BX4 U60 ( .AN(n17), .B(n31), .Y(ab_2__1_) );
  NOR2BX2 U61 ( .AN(A[5]), .B(n33), .Y(ab_5__0_) );
  XOR2X2 U62 ( .A(ab_1__6_), .B(ab_0__7_), .Y(SUMB_1__6_) );
  AND2X4 U63 ( .A(n3), .B(ab_1__5_), .Y(n16) );
  AND3X2 U64 ( .A(n5), .B(B[1]), .C(n35), .Y(CARRYB_1__0_) );
  NOR2BX2 U65 ( .AN(A[3]), .B(n33), .Y(ab_3__0_) );
  NOR2BX2 U66 ( .AN(A[3]), .B(n36), .Y(ab_3__6_) );
  NOR2BX4 U67 ( .AN(B[3]), .B(n34), .Y(ab_0__3_) );
  NOR2BX4 U68 ( .AN(n17), .B(n27), .Y(ab_2__3_) );
  XOR2X4 U69 ( .A(ab_1__5_), .B(n3), .Y(SUMB_1__5_) );
  XOR2X4 U70 ( .A(ab_1__4_), .B(ab_0__5_), .Y(SUMB_1__4_) );
  NOR2BX4 U71 ( .AN(B[5]), .B(n34), .Y(ab_0__5_) );
  BUFX16 U72 ( .A(n39), .Y(n27) );
  BUFX20 U73 ( .A(n39), .Y(n28) );
  BUFX16 U74 ( .A(n41), .Y(n31) );
  NOR2BX4 U75 ( .AN(n17), .B(n38), .Y(ab_2__4_) );
  NOR2BX4 U76 ( .AN(n18), .B(n29), .Y(ab_1__2_) );
  XOR2X2 U77 ( .A(CARRYB_16__5_), .B(SUMB_16__6_), .Y(A1_20_) );
  NOR2BX4 U78 ( .AN(n18), .B(n38), .Y(ab_1__4_) );
  AND2X4 U79 ( .A(CARRYB_16__0_), .B(SUMB_16__1_), .Y(n20) );
  AND2X4 U80 ( .A(CARRYB_16__3_), .B(SUMB_16__4_), .Y(n21) );
  NOR2BX4 U81 ( .AN(n17), .B(n36), .Y(ab_2__6_) );
  NOR2BX2 U82 ( .AN(A[5]), .B(n31), .Y(ab_5__1_) );
  NOR2BX2 U83 ( .AN(A[4]), .B(n31), .Y(ab_4__1_) );
  NOR2BX2 U84 ( .AN(A[6]), .B(n31), .Y(ab_6__1_) );
  NOR2BX2 U85 ( .AN(B[7]), .B(n34), .Y(ab_0__7_) );
  INVX8 U86 ( .A(A[0]), .Y(n34) );
  NOR2BX4 U87 ( .AN(n18), .B(n31), .Y(n44) );
  NOR2BX4 U88 ( .AN(n18), .B(n37), .Y(ab_1__5_) );
  NOR2BX4 U89 ( .AN(n18), .B(n27), .Y(ab_1__3_) );
  XOR2X4 U90 ( .A(CARRYB_16__4_), .B(SUMB_16__5_), .Y(A1_19_) );
  NOR2BX4 U91 ( .AN(n18), .B(n36), .Y(ab_1__6_) );
  NOR2BXL U92 ( .AN(A[16]), .B(n33), .Y(ab_16__0_) );
  NOR2BX1 U93 ( .AN(A[9]), .B(n32), .Y(ab_9__1_) );
  NOR2BX2 U94 ( .AN(A[15]), .B(n33), .Y(ab_15__0_) );
  NOR2BX4 U95 ( .AN(A[15]), .B(n30), .Y(ab_15__2_) );
  NOR2BX2 U96 ( .AN(A[12]), .B(n33), .Y(ab_12__0_) );
  NOR2BX2 U97 ( .AN(A[7]), .B(n29), .Y(ab_7__2_) );
  NOR2BX2 U98 ( .AN(A[14]), .B(n32), .Y(ab_14__1_) );
  AND2X2 U99 ( .A(CARRYB_16__2_), .B(SUMB_16__3_), .Y(n19) );
  NOR2BX1 U100 ( .AN(A[8]), .B(n29), .Y(ab_8__2_) );
  BUFX12 U101 ( .A(n40), .Y(n29) );
  NOR2BX1 U102 ( .AN(A[8]), .B(n37), .Y(ab_8__5_) );
  NOR2BX1 U103 ( .AN(A[10]), .B(n25), .Y(ab_10__5_) );
  NOR2BX1 U104 ( .AN(A[8]), .B(n33), .Y(ab_8__0_) );
  NOR2BX1 U105 ( .AN(A[7]), .B(n33), .Y(ab_7__0_) );
  NOR2BX1 U106 ( .AN(A[6]), .B(n33), .Y(ab_6__0_) );
  NOR2BX1 U107 ( .AN(A[6]), .B(n29), .Y(ab_6__2_) );
  NOR2BX1 U108 ( .AN(A[5]), .B(n37), .Y(ab_5__5_) );
  NOR2BX1 U109 ( .AN(A[4]), .B(n37), .Y(ab_4__5_) );
  NOR2BX1 U110 ( .AN(A[7]), .B(n27), .Y(ab_7__3_) );
  NOR2BX1 U111 ( .AN(A[6]), .B(n25), .Y(ab_6__5_) );
  NOR2BX1 U112 ( .AN(A[7]), .B(n25), .Y(ab_7__5_) );
  NOR2BX1 U113 ( .AN(A[14]), .B(n26), .Y(ab_14__4_) );
  NOR2BX2 U114 ( .AN(A[14]), .B(n33), .Y(ab_14__0_) );
  NOR2BX1 U115 ( .AN(A[12]), .B(n25), .Y(ab_12__5_) );
  NOR2BX1 U116 ( .AN(A[12]), .B(n26), .Y(ab_12__4_) );
  NOR2BX1 U117 ( .AN(A[3]), .B(n43), .Y(ab_3__7_) );
  NOR2BX1 U118 ( .AN(A[4]), .B(n36), .Y(ab_4__6_) );
  NOR2BX1 U119 ( .AN(A[9]), .B(n24), .Y(ab_9__6_) );
  NOR2BX1 U120 ( .AN(A[8]), .B(n43), .Y(ab_8__7_) );
  NOR2BX1 U121 ( .AN(A[8]), .B(n36), .Y(ab_8__6_) );
  NOR2BX1 U122 ( .AN(A[7]), .B(n43), .Y(ab_7__7_) );
  NOR2BX1 U123 ( .AN(A[5]), .B(n43), .Y(ab_5__7_) );
  NOR2BX1 U124 ( .AN(A[15]), .B(n28), .Y(ab_15__3_) );
  NOR2BX1 U125 ( .AN(A[9]), .B(n43), .Y(ab_9__7_) );
  NOR2BX1 U126 ( .AN(A[15]), .B(n25), .Y(ab_15__5_) );
  NOR2BX1 U127 ( .AN(A[11]), .B(n43), .Y(ab_11__7_) );
  NOR2BX1 U128 ( .AN(A[12]), .B(n24), .Y(ab_12__6_) );
  NOR2BX1 U129 ( .AN(A[13]), .B(n43), .Y(ab_13__7_) );
  NOR2BX1 U130 ( .AN(A[12]), .B(n43), .Y(ab_12__7_) );
  BUFX3 U131 ( .A(n41), .Y(n32) );
  CLKBUFXL U132 ( .A(n40), .Y(n30) );
  NOR2BXL U133 ( .AN(A[11]), .B(n25), .Y(ab_11__5_) );
  NOR2BX1 U134 ( .AN(A[10]), .B(n26), .Y(ab_10__4_) );
  NOR2BXL U135 ( .AN(A[11]), .B(n32), .Y(ab_11__1_) );
  NOR2BXL U136 ( .AN(A[11]), .B(n33), .Y(ab_11__0_) );
  NOR2BXL U137 ( .AN(A[10]), .B(n33), .Y(ab_10__0_) );
  NOR2BX2 U138 ( .AN(A[9]), .B(n33), .Y(ab_9__0_) );
  NOR2BX1 U139 ( .AN(A[13]), .B(n28), .Y(ab_13__3_) );
  NOR2BX1 U140 ( .AN(A[14]), .B(n25), .Y(ab_14__5_) );
  NOR2BX1 U141 ( .AN(A[11]), .B(n26), .Y(ab_11__4_) );
  NOR2BXL U142 ( .AN(A[13]), .B(n33), .Y(ab_13__0_) );
  NOR2BX1 U143 ( .AN(A[12]), .B(n32), .Y(ab_12__1_) );
  NOR2BX1 U144 ( .AN(A[10]), .B(n28), .Y(ab_10__3_) );
  NOR2BX1 U145 ( .AN(A[4]), .B(n27), .Y(ab_4__3_) );
  NOR2BX1 U146 ( .AN(A[13]), .B(n26), .Y(ab_13__4_) );
  NOR2BXL U147 ( .AN(A[13]), .B(n32), .Y(ab_13__1_) );
  NOR2BX1 U148 ( .AN(A[11]), .B(n28), .Y(ab_11__3_) );
  NOR2BX1 U149 ( .AN(A[9]), .B(n30), .Y(ab_9__2_) );
  NOR2BX1 U150 ( .AN(A[5]), .B(n38), .Y(ab_5__4_) );
  NOR2BX1 U151 ( .AN(A[5]), .B(n27), .Y(ab_5__3_) );
  NOR2BXL U152 ( .AN(A[13]), .B(n25), .Y(ab_13__5_) );
  NOR2BXL U153 ( .AN(A[13]), .B(n30), .Y(ab_13__2_) );
  NOR2BXL U154 ( .AN(A[10]), .B(n30), .Y(ab_10__2_) );
  NOR2BX1 U155 ( .AN(A[6]), .B(n26), .Y(ab_6__4_) );
  NOR2BX1 U156 ( .AN(A[4]), .B(n29), .Y(ab_4__2_) );
  NOR2BX1 U157 ( .AN(A[6]), .B(n27), .Y(ab_6__3_) );
  AND2X2 U158 ( .A(CARRYB_16__4_), .B(SUMB_16__5_), .Y(n22) );
  NOR2BX1 U159 ( .AN(A[4]), .B(n38), .Y(ab_4__4_) );
  INVXL U160 ( .A(B[0]), .Y(n42) );
  XOR2X1 U161 ( .A(CARRYB_16__6_), .B(ab_16__7_), .Y(A1_21_) );
  AND2X2 U162 ( .A(CARRYB_16__5_), .B(SUMB_16__6_), .Y(n23) );
  NOR2BX1 U163 ( .AN(A[16]), .B(n24), .Y(ab_16__6_) );
  NOR2BXL U164 ( .AN(A[15]), .B(n43), .Y(ab_15__7_) );
  NOR2BX1 U165 ( .AN(A[16]), .B(n25), .Y(ab_16__5_) );
  NOR2BX1 U166 ( .AN(A[16]), .B(n26), .Y(ab_16__4_) );
  NOR2BX1 U167 ( .AN(A[6]), .B(n43), .Y(ab_6__7_) );
  NOR2BX1 U168 ( .AN(A[16]), .B(n32), .Y(ab_16__1_) );
  NOR2BX1 U169 ( .AN(A[16]), .B(n30), .Y(ab_16__2_) );
  NOR2BX1 U170 ( .AN(A[13]), .B(n24), .Y(ab_13__6_) );
  NOR2BXL U171 ( .AN(A[14]), .B(n43), .Y(ab_14__7_) );
  NOR2BX1 U172 ( .AN(A[15]), .B(n24), .Y(ab_15__6_) );
  NOR2BX1 U173 ( .AN(A[14]), .B(n24), .Y(ab_14__6_) );
  NOR2BX1 U174 ( .AN(A[10]), .B(n24), .Y(ab_10__6_) );
  NOR2BXL U175 ( .AN(A[10]), .B(n43), .Y(ab_10__7_) );
  NOR2BX1 U176 ( .AN(A[11]), .B(n24), .Y(ab_11__6_) );
  NOR2BX1 U177 ( .AN(n17), .B(n43), .Y(ab_2__7_) );
  NOR2BX1 U178 ( .AN(A[15]), .B(n26), .Y(ab_15__4_) );
  NOR2BX1 U179 ( .AN(A[4]), .B(n43), .Y(ab_4__7_) );
  NOR2BXL U180 ( .AN(A[16]), .B(n43), .Y(ab_16__7_) );
  NOR2BX1 U181 ( .AN(A[0]), .B(n33), .Y(n35) );
  NOR2BX2 U182 ( .AN(B[6]), .B(n34), .Y(ab_0__6_) );
  XOR2X4 U183 ( .A(SUMB_16__3_), .B(CARRYB_16__2_), .Y(A1_17_) );
  XOR2X4 U184 ( .A(SUMB_16__2_), .B(CARRYB_16__1_), .Y(A1_16_) );
  XOR2X4 U185 ( .A(CARRYB_16__3_), .B(SUMB_16__4_), .Y(A1_18_) );
  XOR2X4 U186 ( .A(SUMB_16__1_), .B(CARRYB_16__0_), .Y(A1_15_) );
  NOR2BX1 U187 ( .AN(n5), .B(n43), .Y(ab_1__7_) );
  INVX8 U188 ( .A(B[5]), .Y(n37) );
  INVX20 U189 ( .A(B[7]), .Y(n43) );
endmodule


module multi16_6 ( in_17bit, in_8bit, out );
  input [16:0] in_17bit;
  input [7:0] in_8bit;
  output [16:0] out;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114;
  wire   [16:1] in_17bit_b;
  wire   [7:1] in_8bit_b;
  wire   [23:8] mul;

  multi16_6_DW02_mult_0 mult_55 ( .A({in_17bit_b[16:4], n2, in_17bit_b[2:1], 
        n13}), .B({in_8bit_b, in_8bit[0]}), .PRODUCT_23_(mul[23]), 
        .PRODUCT_22_(mul[22]), .PRODUCT_21_(mul[21]), .PRODUCT_20_(mul[20]), 
        .PRODUCT_19_(mul[19]), .PRODUCT_18_(mul[18]), .PRODUCT_17_(mul[17]), 
        .PRODUCT_16_(mul[16]), .PRODUCT_15_(mul[15]), .PRODUCT_14_(mul[14]), 
        .PRODUCT_13_(mul[13]), .PRODUCT_12_(mul[12]), .PRODUCT_11_(mul[11]), 
        .PRODUCT_10_(mul[10]), .PRODUCT_9_(mul[9]), .PRODUCT_8_(mul[8]), 
        .PRODUCT_7_(out[0]) );
  BUFX4 U2 ( .A(n10), .Y(n1) );
  INVX20 U3 ( .A(in_17bit[0]), .Y(n12) );
  NAND2X2 U4 ( .A(n5), .B(n60), .Y(n59) );
  NAND2X2 U5 ( .A(n33), .B(n58), .Y(n60) );
  BUFX12 U6 ( .A(in_17bit[16]), .Y(n38) );
  NAND2BX4 U7 ( .AN(in_8bit[0]), .B(n25), .Y(n43) );
  BUFX12 U8 ( .A(in_17bit_b[3]), .Y(n2) );
  INVX4 U9 ( .A(in_17bit[2]), .Y(n56) );
  NOR2BX4 U10 ( .AN(n38), .B(n10), .Y(n55) );
  INVX12 U11 ( .A(n38), .Y(n83) );
  CLKINVX2 U12 ( .A(n83), .Y(n5) );
  OR2X1 U13 ( .A(n28), .B(n83), .Y(n26) );
  OR2XL U14 ( .A(n31), .B(n83), .Y(n21) );
  OR2X2 U15 ( .A(n33), .B(n83), .Y(n27) );
  OR2X4 U16 ( .A(in_17bit[1]), .B(in_17bit[0]), .Y(n54) );
  XOR2X4 U17 ( .A(mul[13]), .B(n3), .Y(out[6]) );
  AND2X2 U18 ( .A(n93), .B(n106), .Y(n3) );
  NAND2X2 U19 ( .A(n38), .B(n64), .Y(n63) );
  INVXL U20 ( .A(in_17bit[13]), .Y(n79) );
  INVXL U21 ( .A(in_17bit[7]), .Y(n65) );
  INVX2 U22 ( .A(n70), .Y(n32) );
  NAND2X2 U23 ( .A(n31), .B(n71), .Y(n72) );
  XNOR2X4 U24 ( .A(mul[8]), .B(n85), .Y(out[1]) );
  CLKINVX2 U25 ( .A(n98), .Y(n4) );
  OR2X4 U26 ( .A(in_17bit[1]), .B(n38), .Y(n36) );
  NAND3X2 U27 ( .A(in_17bit[0]), .B(n38), .C(in_17bit[1]), .Y(n37) );
  XNOR2X4 U28 ( .A(n46), .B(n34), .Y(in_8bit_b[3]) );
  INVX4 U29 ( .A(n48), .Y(n50) );
  NAND4BX4 U30 ( .AN(in_8bit[0]), .B(n25), .C(n46), .D(n45), .Y(n48) );
  NOR3X1 U31 ( .A(in_17bit[15]), .B(n84), .C(n83), .Y(in_17bit_b[16]) );
  OAI21XL U32 ( .A0(in_8bit[1]), .A1(in_8bit[0]), .B0(n39), .Y(n42) );
  OR2X4 U33 ( .A(mul[14]), .B(n94), .Y(n95) );
  NAND2X4 U34 ( .A(n95), .B(n106), .Y(n15) );
  NAND2BX4 U35 ( .AN(mul[16]), .B(n4), .Y(n99) );
  XOR2X4 U36 ( .A(mul[23]), .B(n114), .Y(out[16]) );
  XNOR2X4 U37 ( .A(mul[10]), .B(n87), .Y(out[3]) );
  NAND2X4 U38 ( .A(n88), .B(n106), .Y(n87) );
  BUFX4 U39 ( .A(n105), .Y(n6) );
  OR2X4 U40 ( .A(mul[10]), .B(n88), .Y(n90) );
  XNOR2X2 U41 ( .A(mul[11]), .B(n89), .Y(out[4]) );
  NAND2X2 U42 ( .A(n39), .B(n48), .Y(n47) );
  INVX4 U43 ( .A(mul[22]), .Y(n109) );
  NOR2BX4 U44 ( .AN(n106), .B(n23), .Y(n102) );
  NOR2X1 U45 ( .A(mul[20]), .B(n11), .Y(n112) );
  NAND2BX4 U46 ( .AN(mul[20]), .B(n6), .Y(n107) );
  NAND2X2 U47 ( .A(n38), .B(n57), .Y(n8) );
  NOR2X4 U48 ( .A(n105), .B(n7), .Y(n103) );
  CLKINVX20 U49 ( .A(n106), .Y(n7) );
  INVX2 U50 ( .A(in_8bit[5]), .Y(n49) );
  INVXL U51 ( .A(in_8bit[2]), .Y(n41) );
  XNOR2X4 U52 ( .A(in_17bit[3]), .B(n8), .Y(in_17bit_b[3]) );
  XOR2X2 U53 ( .A(n42), .B(n41), .Y(in_8bit_b[2]) );
  NAND2X2 U54 ( .A(n86), .B(n106), .Y(n16) );
  XNOR2X4 U55 ( .A(mul[9]), .B(n16), .Y(out[2]) );
  NOR2X4 U56 ( .A(n60), .B(n29), .Y(n28) );
  NAND2X4 U57 ( .A(n28), .B(n62), .Y(n64) );
  CLKINVX8 U58 ( .A(in_17bit[6]), .Y(n62) );
  OR2X2 U59 ( .A(mul[17]), .B(n99), .Y(n9) );
  NOR2X4 U60 ( .A(in_17bit[0]), .B(in_17bit[1]), .Y(n10) );
  XOR2X4 U61 ( .A(mul[14]), .B(n14), .Y(out[7]) );
  XOR2X4 U62 ( .A(n55), .B(in_17bit[2]), .Y(in_17bit_b[2]) );
  INVX3 U63 ( .A(mul[19]), .Y(n101) );
  AND2X1 U64 ( .A(in_8bit[0]), .B(n39), .Y(n24) );
  XOR2X4 U65 ( .A(n26), .B(n62), .Y(in_17bit_b[6]) );
  NOR2X1 U66 ( .A(mul[21]), .B(mul[22]), .Y(n113) );
  XNOR2X4 U67 ( .A(mul[15]), .B(n15), .Y(out[8]) );
  XNOR2X4 U68 ( .A(mul[12]), .B(n91), .Y(out[5]) );
  OAI21X4 U69 ( .A0(mul[21]), .A1(n107), .B0(n106), .Y(n108) );
  AND2X4 U70 ( .A(n39), .B(n43), .Y(n34) );
  XOR2X4 U71 ( .A(n61), .B(n59), .Y(in_17bit_b[5]) );
  OAI21X4 U72 ( .A0(mul[20]), .A1(n11), .B0(n106), .Y(n104) );
  XOR2X4 U73 ( .A(n109), .B(n108), .Y(out[15]) );
  NOR2X2 U74 ( .A(n64), .B(in_17bit[7]), .Y(n22) );
  NAND2BX2 U75 ( .AN(mul[19]), .B(n23), .Y(n11) );
  INVX8 U76 ( .A(n110), .Y(n105) );
  CLKINVX4 U77 ( .A(n12), .Y(n13) );
  AND2X4 U78 ( .A(n94), .B(n106), .Y(n14) );
  NOR2X4 U79 ( .A(in_8bit[2]), .B(in_8bit[1]), .Y(n25) );
  OR2X4 U80 ( .A(mul[8]), .B(out[0]), .Y(n86) );
  XNOR2X4 U81 ( .A(mul[18]), .B(n18), .Y(out[11]) );
  XOR2X4 U82 ( .A(n27), .B(n58), .Y(in_17bit_b[4]) );
  NOR2X4 U83 ( .A(in_17bit[3]), .B(n57), .Y(n33) );
  NAND2X4 U84 ( .A(n1), .B(n56), .Y(n57) );
  NAND2X2 U85 ( .A(n92), .B(n106), .Y(n91) );
  XNOR2X4 U86 ( .A(mul[17]), .B(n17), .Y(out[10]) );
  CLKINVX3 U87 ( .A(n61), .Y(n29) );
  NAND2X2 U88 ( .A(n22), .B(n67), .Y(n69) );
  NAND2X4 U89 ( .A(n53), .B(n39), .Y(n52) );
  NAND2X4 U90 ( .A(n99), .B(n106), .Y(n17) );
  NAND2X4 U91 ( .A(n100), .B(n106), .Y(n18) );
  NAND2X2 U92 ( .A(n30), .B(n81), .Y(n84) );
  OR2X4 U93 ( .A(mul[17]), .B(n99), .Y(n100) );
  CLKINVX8 U94 ( .A(n40), .Y(n39) );
  NOR2XL U95 ( .A(n78), .B(in_17bit[13]), .Y(n30) );
  NAND2BXL U96 ( .AN(n72), .B(n73), .Y(n74) );
  NAND2BX4 U97 ( .AN(mul[19]), .B(n23), .Y(n110) );
  OR2X4 U98 ( .A(mul[12]), .B(n92), .Y(n93) );
  OR2X4 U99 ( .A(mul[11]), .B(n90), .Y(n92) );
  OR2X4 U100 ( .A(mul[9]), .B(n86), .Y(n88) );
  AOI21X2 U101 ( .A0(n113), .A1(n112), .B0(n111), .Y(n114) );
  INVX4 U102 ( .A(n111), .Y(n106) );
  NOR2X4 U103 ( .A(n69), .B(n32), .Y(n31) );
  XOR2X2 U104 ( .A(n73), .B(n19), .Y(in_17bit_b[11]) );
  NAND2XL U105 ( .A(n5), .B(n72), .Y(n19) );
  XOR2X2 U106 ( .A(n79), .B(n20), .Y(in_17bit_b[13]) );
  NAND2XL U107 ( .A(n5), .B(n78), .Y(n20) );
  XOR2X2 U108 ( .A(n21), .B(n71), .Y(in_17bit_b[10]) );
  NOR2X4 U109 ( .A(mul[18]), .B(n9), .Y(n23) );
  OR2X2 U110 ( .A(mul[13]), .B(n93), .Y(n94) );
  NAND2XL U111 ( .A(n90), .B(n106), .Y(n89) );
  NAND2X1 U112 ( .A(out[0]), .B(n106), .Y(n85) );
  XOR2X2 U113 ( .A(in_8bit[1]), .B(n24), .Y(in_8bit_b[1]) );
  INVX8 U114 ( .A(in_8bit[7]), .Y(n40) );
  NOR2XL U115 ( .A(n22), .B(n83), .Y(n66) );
  NOR2XL U116 ( .A(n30), .B(n83), .Y(n80) );
  NAND2XL U117 ( .A(n38), .B(n69), .Y(n68) );
  NOR2XL U118 ( .A(n77), .B(n83), .Y(n75) );
  XNOR2X1 U119 ( .A(n38), .B(n39), .Y(n111) );
  XNOR2X2 U120 ( .A(n82), .B(n35), .Y(in_17bit_b[15]) );
  AND2X1 U121 ( .A(n5), .B(n84), .Y(n35) );
  INVX1 U122 ( .A(in_8bit[6]), .Y(n51) );
  INVX1 U123 ( .A(in_8bit[4]), .Y(n45) );
  INVX1 U124 ( .A(in_8bit[3]), .Y(n46) );
  AND3X4 U125 ( .A(n36), .B(n54), .C(n37), .Y(in_17bit_b[1]) );
  OAI21X4 U126 ( .A0(in_8bit[3]), .A1(n43), .B0(n39), .Y(n44) );
  XOR2X4 U127 ( .A(n44), .B(n45), .Y(in_8bit_b[4]) );
  XOR2X4 U128 ( .A(n49), .B(n47), .Y(in_8bit_b[5]) );
  NAND2X4 U129 ( .A(n50), .B(n49), .Y(n53) );
  XOR2X4 U130 ( .A(n52), .B(n51), .Y(in_8bit_b[6]) );
  NOR3X4 U131 ( .A(in_8bit[6]), .B(n53), .C(n40), .Y(in_8bit_b[7]) );
  CLKINVX3 U132 ( .A(in_17bit[4]), .Y(n58) );
  CLKINVX3 U133 ( .A(in_17bit[5]), .Y(n61) );
  XOR2X4 U134 ( .A(n65), .B(n63), .Y(in_17bit_b[7]) );
  CLKINVX3 U135 ( .A(in_17bit[8]), .Y(n67) );
  XNOR2X4 U136 ( .A(n66), .B(n67), .Y(in_17bit_b[8]) );
  CLKINVX3 U137 ( .A(in_17bit[9]), .Y(n70) );
  XOR2X4 U138 ( .A(n70), .B(n68), .Y(in_17bit_b[9]) );
  CLKINVX3 U139 ( .A(in_17bit[10]), .Y(n71) );
  CLKINVX3 U140 ( .A(in_17bit[11]), .Y(n73) );
  CLKINVX3 U141 ( .A(n74), .Y(n77) );
  CLKINVX3 U142 ( .A(in_17bit[12]), .Y(n76) );
  XNOR2X4 U143 ( .A(n75), .B(n76), .Y(in_17bit_b[12]) );
  NAND2X4 U144 ( .A(n77), .B(n76), .Y(n78) );
  CLKINVX3 U145 ( .A(in_17bit[14]), .Y(n81) );
  XNOR2X4 U146 ( .A(n80), .B(n81), .Y(in_17bit_b[14]) );
  CLKINVX3 U147 ( .A(in_17bit[15]), .Y(n82) );
  CLKINVX3 U148 ( .A(n95), .Y(n96) );
  NAND2BX4 U149 ( .AN(mul[15]), .B(n96), .Y(n98) );
  NAND2X4 U150 ( .A(n98), .B(n106), .Y(n97) );
  XNOR2X4 U151 ( .A(mul[16]), .B(n97), .Y(out[9]) );
  XNOR2X4 U152 ( .A(n102), .B(n101), .Y(out[12]) );
  XOR2X4 U153 ( .A(n103), .B(mul[20]), .Y(out[13]) );
  XNOR2X4 U154 ( .A(n104), .B(mul[21]), .Y(out[14]) );
endmodule


module multi16_5_DW01_add_4 ( A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, 
        A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, 
        B_20_, B_19_, B_18_, B_17_, B_16_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, 
        SUM_17_, SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, 
        SUM_9_, SUM_8_, SUM_7_, SUM_6_, SUM_5_ );
  input A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_,
         A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, B_20_, B_19_,
         B_18_, B_17_, B_16_;
  output SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, SUM_15_,
         SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, SUM_7_,
         SUM_6_, SUM_5_;
  wire   n1, n2, n3, n4, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42;

  AOI2BB1X4 U2 ( .A0N(n1), .A1N(n2), .B0(n29), .Y(n22) );
  OR2X2 U3 ( .A(n32), .B(n33), .Y(n1) );
  AND2X2 U4 ( .A(n30), .B(n31), .Y(n2) );
  BUFX12 U5 ( .A(A_14_), .Y(SUM_14_) );
  AOI2BB1X4 U6 ( .A0N(n32), .A1N(n31), .B0(n29), .Y(n37) );
  NAND2X2 U7 ( .A(B_19_), .B(A_19_), .Y(n25) );
  BUFX8 U8 ( .A(A_6_), .Y(SUM_6_) );
  XOR3X4 U9 ( .A(B_21_), .B(A_21_), .C(n16), .Y(SUM_21_) );
  XNOR2X4 U10 ( .A(n41), .B(n30), .Y(SUM_17_) );
  NAND2X4 U11 ( .A(n38), .B(n26), .Y(n40) );
  NAND2X4 U12 ( .A(n36), .B(n37), .Y(n34) );
  NAND2X4 U13 ( .A(n31), .B(n3), .Y(n39) );
  OR2X4 U14 ( .A(A_16_), .B(B_16_), .Y(n28) );
  NAND2X4 U15 ( .A(A_16_), .B(B_16_), .Y(n30) );
  BUFX12 U16 ( .A(A_15_), .Y(SUM_15_) );
  NAND2X2 U17 ( .A(n17), .B(n18), .Y(n16) );
  NAND2X4 U18 ( .A(n28), .B(n30), .Y(n42) );
  INVX4 U19 ( .A(n27), .Y(n33) );
  INVX4 U20 ( .A(n38), .Y(n29) );
  NAND2X2 U21 ( .A(B_18_), .B(A_18_), .Y(n38) );
  NOR2X4 U22 ( .A(A_19_), .B(B_19_), .Y(n4) );
  INVX8 U23 ( .A(n42), .Y(SUM_16_) );
  NAND2BX2 U24 ( .AN(n3), .B(n26), .Y(n36) );
  INVX4 U25 ( .A(n26), .Y(n32) );
  XNOR2X4 U26 ( .A(n39), .B(n40), .Y(SUM_18_) );
  NOR2BX4 U27 ( .AN(n25), .B(n4), .Y(n35) );
  NAND2X2 U28 ( .A(B_20_), .B(A_20_), .Y(n17) );
  AND2X2 U29 ( .A(n17), .B(n20), .Y(n21) );
  BUFX4 U30 ( .A(A_9_), .Y(SUM_9_) );
  OR2X4 U31 ( .A(B_18_), .B(A_18_), .Y(n26) );
  NAND3X4 U32 ( .A(n27), .B(B_16_), .C(A_16_), .Y(n3) );
  OR2X4 U33 ( .A(A_20_), .B(B_20_), .Y(n20) );
  INVX1 U34 ( .A(n24), .Y(n23) );
  INVX1 U35 ( .A(n25), .Y(n24) );
  NAND2XL U36 ( .A(n19), .B(n20), .Y(n18) );
  BUFX8 U37 ( .A(A_12_), .Y(SUM_12_) );
  BUFX8 U38 ( .A(A_5_), .Y(SUM_5_) );
  BUFX8 U39 ( .A(A_11_), .Y(SUM_11_) );
  BUFX8 U40 ( .A(A_10_), .Y(SUM_10_) );
  BUFX4 U41 ( .A(A_8_), .Y(SUM_8_) );
  BUFX4 U42 ( .A(A_7_), .Y(SUM_7_) );
  BUFX8 U43 ( .A(A_13_), .Y(SUM_13_) );
  XOR2X4 U44 ( .A(n19), .B(n21), .Y(SUM_20_) );
  OAI21X4 U45 ( .A0(n22), .A1(n4), .B0(n23), .Y(n19) );
  XOR2X4 U46 ( .A(n34), .B(n35), .Y(SUM_19_) );
  NOR2BX4 U47 ( .AN(n31), .B(n33), .Y(n41) );
  OR2X4 U48 ( .A(A_17_), .B(B_17_), .Y(n27) );
  NAND2X4 U49 ( .A(B_17_), .B(A_17_), .Y(n31) );
endmodule


module multi16_5_DW02_mult_0 ( A, B, PRODUCT_23_, PRODUCT_22_, PRODUCT_21_, 
        PRODUCT_20_, PRODUCT_19_, PRODUCT_18_, PRODUCT_17_, PRODUCT_16_, 
        PRODUCT_15_, PRODUCT_14_, PRODUCT_13_, PRODUCT_12_, PRODUCT_11_, 
        PRODUCT_10_, PRODUCT_9_, PRODUCT_8_, PRODUCT_7_ );
  input [16:0] A;
  input [7:0] B;
  output PRODUCT_23_, PRODUCT_22_, PRODUCT_21_, PRODUCT_20_, PRODUCT_19_,
         PRODUCT_18_, PRODUCT_17_, PRODUCT_16_, PRODUCT_15_, PRODUCT_14_,
         PRODUCT_13_, PRODUCT_12_, PRODUCT_11_, PRODUCT_10_, PRODUCT_9_,
         PRODUCT_8_, PRODUCT_7_;
  wire   ab_16__7_, ab_16__6_, ab_16__5_, ab_16__4_, ab_16__3_, ab_16__2_,
         ab_16__1_, ab_16__0_, ab_15__7_, ab_15__6_, ab_15__5_, ab_15__4_,
         ab_15__3_, ab_15__2_, ab_15__1_, ab_15__0_, ab_14__7_, ab_14__6_,
         ab_14__5_, ab_14__4_, ab_14__3_, ab_14__2_, ab_14__1_, ab_14__0_,
         ab_13__7_, ab_13__6_, ab_13__5_, ab_13__4_, ab_13__3_, ab_13__2_,
         ab_13__1_, ab_13__0_, ab_12__7_, ab_12__6_, ab_12__5_, ab_12__4_,
         ab_12__3_, ab_12__2_, ab_12__1_, ab_12__0_, ab_11__7_, ab_11__6_,
         ab_11__5_, ab_11__4_, ab_11__3_, ab_11__2_, ab_11__1_, ab_11__0_,
         ab_10__7_, ab_10__6_, ab_10__5_, ab_10__4_, ab_10__3_, ab_10__2_,
         ab_10__1_, ab_10__0_, ab_9__7_, ab_9__6_, ab_9__5_, ab_9__4_,
         ab_9__3_, ab_9__2_, ab_9__1_, ab_9__0_, ab_8__7_, ab_8__6_, ab_8__5_,
         ab_8__4_, ab_8__3_, ab_8__2_, ab_8__1_, ab_8__0_, ab_7__7_, ab_7__6_,
         ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_, ab_7__0_, ab_6__7_,
         ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_, ab_6__1_, ab_6__0_,
         ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_, ab_5__2_, ab_5__1_,
         ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_, ab_4__3_, ab_4__2_,
         ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_, ab_3__4_, ab_3__3_,
         ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_, ab_2__5_, ab_2__4_,
         ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_, ab_1__6_, ab_1__5_,
         ab_1__4_, ab_1__3_, ab_1__2_, ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_,
         ab_0__3_, ab_0__2_, CARRYB_16__6_, CARRYB_16__5_, CARRYB_16__4_,
         CARRYB_16__3_, CARRYB_16__2_, CARRYB_16__1_, CARRYB_16__0_,
         CARRYB_15__6_, CARRYB_15__5_, CARRYB_15__4_, CARRYB_15__3_,
         CARRYB_15__2_, CARRYB_15__1_, CARRYB_15__0_, CARRYB_14__6_,
         CARRYB_14__5_, CARRYB_14__4_, CARRYB_14__3_, CARRYB_14__2_,
         CARRYB_14__1_, CARRYB_14__0_, CARRYB_13__6_, CARRYB_13__5_,
         CARRYB_13__4_, CARRYB_13__3_, CARRYB_13__2_, CARRYB_13__1_,
         CARRYB_13__0_, CARRYB_12__6_, CARRYB_12__5_, CARRYB_12__4_,
         CARRYB_12__3_, CARRYB_12__2_, CARRYB_12__1_, CARRYB_12__0_,
         CARRYB_11__6_, CARRYB_11__5_, CARRYB_11__4_, CARRYB_11__3_,
         CARRYB_11__2_, CARRYB_11__1_, CARRYB_11__0_, CARRYB_10__6_,
         CARRYB_10__5_, CARRYB_10__4_, CARRYB_10__3_, CARRYB_10__2_,
         CARRYB_10__1_, CARRYB_10__0_, CARRYB_9__6_, CARRYB_9__5_,
         CARRYB_9__4_, CARRYB_9__3_, CARRYB_9__2_, CARRYB_9__1_, CARRYB_9__0_,
         CARRYB_8__6_, CARRYB_8__5_, CARRYB_8__4_, CARRYB_8__3_, CARRYB_8__2_,
         CARRYB_8__1_, CARRYB_8__0_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_,
         CARRYB_7__3_, CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_,
         CARRYB_6__5_, CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_,
         CARRYB_6__0_, CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_,
         CARRYB_5__2_, CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_,
         CARRYB_4__4_, CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_,
         CARRYB_3__6_, CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_,
         CARRYB_3__1_, CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_,
         CARRYB_2__3_, CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__0_,
         SUMB_16__6_, SUMB_16__5_, SUMB_16__4_, SUMB_16__3_, SUMB_16__2_,
         SUMB_16__1_, SUMB_16__0_, SUMB_15__6_, SUMB_15__5_, SUMB_15__4_,
         SUMB_15__3_, SUMB_15__2_, SUMB_15__1_, SUMB_14__6_, SUMB_14__5_,
         SUMB_14__4_, SUMB_14__3_, SUMB_14__2_, SUMB_14__1_, SUMB_13__6_,
         SUMB_13__5_, SUMB_13__4_, SUMB_13__3_, SUMB_13__2_, SUMB_13__1_,
         SUMB_12__6_, SUMB_12__5_, SUMB_12__4_, SUMB_12__3_, SUMB_12__2_,
         SUMB_12__1_, SUMB_11__6_, SUMB_11__5_, SUMB_11__4_, SUMB_11__3_,
         SUMB_11__2_, SUMB_11__1_, SUMB_10__6_, SUMB_10__5_, SUMB_10__4_,
         SUMB_10__3_, SUMB_10__2_, SUMB_10__1_, SUMB_9__6_, SUMB_9__5_,
         SUMB_9__4_, SUMB_9__3_, SUMB_9__2_, SUMB_9__1_, SUMB_8__6_,
         SUMB_8__5_, SUMB_8__4_, SUMB_8__3_, SUMB_8__2_, SUMB_8__1_,
         SUMB_7__6_, SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_,
         SUMB_7__1_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, PROD1_7_, A1_21_, A1_20_, A1_19_, A1_18_,
         A1_17_, A1_16_, A1_15_, A1_13_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_,
         A1_7_, A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_17_, n3, n5, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39;

  multi16_5_DW01_add_4 FS_1 ( .A_21_(A1_21_), .A_20_(A1_20_), .A_19_(A1_19_), 
        .A_18_(A1_18_), .A_17_(A1_17_), .A_16_(A1_16_), .A_15_(A1_15_), 
        .A_14_(SUMB_16__0_), .A_13_(A1_13_), .A_12_(A1_12_), .A_11_(A1_11_), 
        .A_10_(A1_10_), .A_9_(A1_9_), .A_8_(A1_8_), .A_7_(A1_7_), .A_6_(A1_6_), 
        .A_5_(PROD1_7_), .B_21_(n10), .B_20_(n17), .B_19_(n16), .B_18_(n15), 
        .B_17_(A2_17_), .B_16_(n14), .SUM_21_(PRODUCT_23_), .SUM_20_(
        PRODUCT_22_), .SUM_19_(PRODUCT_21_), .SUM_18_(PRODUCT_20_), .SUM_17_(
        PRODUCT_19_), .SUM_16_(PRODUCT_18_), .SUM_15_(PRODUCT_17_), .SUM_14_(
        PRODUCT_16_), .SUM_13_(PRODUCT_15_), .SUM_12_(PRODUCT_14_), .SUM_11_(
        PRODUCT_13_), .SUM_10_(PRODUCT_12_), .SUM_9_(PRODUCT_11_), .SUM_8_(
        PRODUCT_10_), .SUM_7_(PRODUCT_9_), .SUM_6_(PRODUCT_8_), .SUM_5_(
        PRODUCT_7_) );
  ADDFHX4 S4_3 ( .A(ab_16__3_), .B(CARRYB_15__3_), .CI(SUMB_15__4_), .CO(
        CARRYB_16__3_), .S(SUMB_16__3_) );
  ADDFHX4 S4_1 ( .A(ab_16__1_), .B(CARRYB_15__1_), .CI(SUMB_15__2_), .CO(
        CARRYB_16__1_), .S(SUMB_16__1_) );
  ADDFHX4 S4_0 ( .A(ab_16__0_), .B(CARRYB_15__0_), .CI(SUMB_15__1_), .CO(
        CARRYB_16__0_), .S(SUMB_16__0_) );
  ADDFHX4 S1_9_0 ( .A(ab_9__0_), .B(CARRYB_8__0_), .CI(SUMB_8__1_), .CO(
        CARRYB_9__0_), .S(A1_7_) );
  ADDFHX4 S1_10_0 ( .A(ab_10__0_), .B(CARRYB_9__0_), .CI(SUMB_9__1_), .CO(
        CARRYB_10__0_), .S(A1_8_) );
  ADDFHX4 S2_14_2 ( .A(ab_14__2_), .B(CARRYB_13__2_), .CI(SUMB_13__3_), .CO(
        CARRYB_14__2_), .S(SUMB_14__2_) );
  ADDFHX4 S2_15_2 ( .A(ab_15__2_), .B(CARRYB_14__2_), .CI(SUMB_14__3_), .CO(
        CARRYB_15__2_), .S(SUMB_15__2_) );
  ADDFHX4 S2_12_1 ( .A(ab_12__1_), .B(CARRYB_11__1_), .CI(SUMB_11__2_), .CO(
        CARRYB_12__1_), .S(SUMB_12__1_) );
  ADDFHX4 S2_13_1 ( .A(ab_13__1_), .B(CARRYB_12__1_), .CI(SUMB_12__2_), .CO(
        CARRYB_13__1_), .S(SUMB_13__1_) );
  ADDFHX4 S2_12_4 ( .A(ab_12__4_), .B(CARRYB_11__4_), .CI(SUMB_11__5_), .CO(
        CARRYB_12__4_), .S(SUMB_12__4_) );
  ADDFHX4 S2_13_4 ( .A(ab_13__4_), .B(CARRYB_12__4_), .CI(SUMB_12__5_), .CO(
        CARRYB_13__4_), .S(SUMB_13__4_) );
  ADDFHX4 S1_8_0 ( .A(ab_8__0_), .B(CARRYB_7__0_), .CI(SUMB_7__1_), .CO(
        CARRYB_8__0_), .S(A1_6_) );
  ADDFHX4 S2_13_3 ( .A(ab_13__3_), .B(CARRYB_12__3_), .CI(SUMB_12__4_), .CO(
        CARRYB_13__3_), .S(SUMB_13__3_) );
  ADDFHX4 S2_14_3 ( .A(ab_14__3_), .B(CARRYB_13__3_), .CI(SUMB_13__4_), .CO(
        CARRYB_14__3_), .S(SUMB_14__3_) );
  ADDFHX4 S2_11_3 ( .A(ab_11__3_), .B(CARRYB_10__3_), .CI(SUMB_10__4_), .CO(
        CARRYB_11__3_), .S(SUMB_11__3_) );
  ADDFHX4 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  ADDFHX4 S1_7_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(PROD1_7_) );
  ADDFHX4 S1_14_0 ( .A(ab_14__0_), .B(CARRYB_13__0_), .CI(SUMB_13__1_), .CO(
        CARRYB_14__0_), .S(A1_12_) );
  ADDFHX4 S1_15_0 ( .A(ab_15__0_), .B(CARRYB_14__0_), .CI(SUMB_14__1_), .CO(
        CARRYB_15__0_), .S(A1_13_) );
  ADDFHX4 S1_11_0 ( .A(ab_11__0_), .B(CARRYB_10__0_), .CI(SUMB_10__1_), .CO(
        CARRYB_11__0_), .S(A1_9_) );
  ADDFHX4 S2_13_5 ( .A(ab_13__5_), .B(CARRYB_12__5_), .CI(SUMB_12__6_), .CO(
        CARRYB_13__5_), .S(SUMB_13__5_) );
  ADDFHX4 S2_14_4 ( .A(ab_14__4_), .B(CARRYB_13__4_), .CI(SUMB_13__5_), .CO(
        CARRYB_14__4_), .S(SUMB_14__4_) );
  ADDFHX4 S2_12_2 ( .A(ab_12__2_), .B(CARRYB_11__2_), .CI(SUMB_11__3_), .CO(
        CARRYB_12__2_), .S(SUMB_12__2_) );
  ADDFHX4 S2_12_3 ( .A(ab_12__3_), .B(CARRYB_11__3_), .CI(SUMB_11__4_), .CO(
        CARRYB_12__3_), .S(SUMB_12__3_) );
  ADDFHX4 S2_13_2 ( .A(ab_13__2_), .B(CARRYB_12__2_), .CI(SUMB_12__3_), .CO(
        CARRYB_13__2_), .S(SUMB_13__2_) );
  ADDFHX4 S2_10_2 ( .A(ab_10__2_), .B(CARRYB_9__2_), .CI(SUMB_9__3_), .CO(
        CARRYB_10__2_), .S(SUMB_10__2_) );
  ADDFHX4 S2_11_2 ( .A(ab_11__2_), .B(CARRYB_10__2_), .CI(SUMB_10__3_), .CO(
        CARRYB_11__2_), .S(SUMB_11__2_) );
  ADDFHX4 S2_12_5 ( .A(ab_12__5_), .B(CARRYB_11__5_), .CI(SUMB_11__6_), .CO(
        CARRYB_12__5_), .S(SUMB_12__5_) );
  ADDFHX4 S2_11_5 ( .A(ab_11__5_), .B(CARRYB_10__5_), .CI(SUMB_10__6_), .CO(
        CARRYB_11__5_), .S(SUMB_11__5_) );
  ADDFHX4 S2_11_1 ( .A(ab_11__1_), .B(CARRYB_10__1_), .CI(SUMB_10__2_), .CO(
        CARRYB_11__1_), .S(SUMB_11__1_) );
  ADDFHX4 S2_10_1 ( .A(ab_10__1_), .B(CARRYB_9__1_), .CI(SUMB_9__2_), .CO(
        CARRYB_10__1_), .S(SUMB_10__1_) );
  ADDFHX4 S1_12_0 ( .A(ab_12__0_), .B(CARRYB_11__0_), .CI(SUMB_11__1_), .CO(
        CARRYB_12__0_), .S(A1_10_) );
  ADDFHX4 S1_13_0 ( .A(ab_13__0_), .B(CARRYB_12__0_), .CI(SUMB_12__1_), .CO(
        CARRYB_13__0_), .S(A1_11_) );
  ADDFHX4 S4_2 ( .A(ab_16__2_), .B(CARRYB_15__2_), .CI(SUMB_15__3_), .CO(
        CARRYB_16__2_), .S(SUMB_16__2_) );
  ADDFHX4 S2_14_1 ( .A(ab_14__1_), .B(CARRYB_13__1_), .CI(SUMB_13__2_), .CO(
        CARRYB_14__1_), .S(SUMB_14__1_) );
  ADDFHX4 S2_9_1 ( .A(ab_9__1_), .B(CARRYB_8__1_), .CI(SUMB_8__2_), .CO(
        CARRYB_9__1_), .S(SUMB_9__1_) );
  ADDFHX4 S2_11_4 ( .A(ab_11__4_), .B(CARRYB_10__4_), .CI(SUMB_10__5_), .CO(
        CARRYB_11__4_), .S(SUMB_11__4_) );
  ADDFHX4 S2_10_3 ( .A(ab_10__3_), .B(CARRYB_9__3_), .CI(SUMB_9__4_), .CO(
        CARRYB_10__3_), .S(SUMB_10__3_) );
  ADDFHX4 S2_9_4 ( .A(ab_9__4_), .B(CARRYB_8__4_), .CI(SUMB_8__5_), .CO(
        CARRYB_9__4_), .S(SUMB_9__4_) );
  ADDFHX4 S2_9_2 ( .A(ab_9__2_), .B(CARRYB_8__2_), .CI(SUMB_8__3_), .CO(
        CARRYB_9__2_), .S(SUMB_9__2_) );
  ADDFHX4 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  ADDFHX4 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  ADDFHX4 S4_4 ( .A(ab_16__4_), .B(CARRYB_15__4_), .CI(SUMB_15__5_), .CO(
        CARRYB_16__4_), .S(SUMB_16__4_) );
  ADDFHX4 S2_10_5 ( .A(ab_10__5_), .B(CARRYB_9__5_), .CI(SUMB_9__6_), .CO(
        CARRYB_10__5_), .S(SUMB_10__5_) );
  ADDFHX4 S2_8_5 ( .A(ab_8__5_), .B(CARRYB_7__5_), .CI(SUMB_7__6_), .CO(
        CARRYB_8__5_), .S(SUMB_8__5_) );
  ADDFHX4 S2_9_5 ( .A(ab_9__5_), .B(CARRYB_8__5_), .CI(SUMB_8__6_), .CO(
        CARRYB_9__5_), .S(SUMB_9__5_) );
  ADDFHX4 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  ADDFHX4 S2_8_1 ( .A(ab_8__1_), .B(CARRYB_7__1_), .CI(SUMB_7__2_), .CO(
        CARRYB_8__1_), .S(SUMB_8__1_) );
  ADDFHX4 S2_15_1 ( .A(ab_15__1_), .B(CARRYB_14__1_), .CI(SUMB_14__2_), .CO(
        CARRYB_15__1_), .S(SUMB_15__1_) );
  ADDFHX4 S3_2_6 ( .A(ab_2__6_), .B(n7), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  ADDFHX4 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  ADDFHX4 S3_9_6 ( .A(ab_9__6_), .B(CARRYB_8__6_), .CI(ab_8__7_), .CO(
        CARRYB_9__6_), .S(SUMB_9__6_) );
  ADDFHX4 S3_10_6 ( .A(ab_10__6_), .B(CARRYB_9__6_), .CI(ab_9__7_), .CO(
        CARRYB_10__6_), .S(SUMB_10__6_) );
  ADDFHX4 S2_7_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  ADDFHX4 S2_7_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  ADDFHX4 S2_8_4 ( .A(ab_8__4_), .B(CARRYB_7__4_), .CI(SUMB_7__5_), .CO(
        CARRYB_8__4_), .S(SUMB_8__4_) );
  ADDFHX4 S2_9_3 ( .A(ab_9__3_), .B(CARRYB_8__3_), .CI(SUMB_8__4_), .CO(
        CARRYB_9__3_), .S(SUMB_9__3_) );
  ADDFHX4 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  ADDFHX4 S2_8_2 ( .A(ab_8__2_), .B(CARRYB_7__2_), .CI(SUMB_7__3_), .CO(
        CARRYB_8__2_), .S(SUMB_8__2_) );
  ADDFHX4 S3_7_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(
        CARRYB_7__6_), .S(SUMB_7__6_) );
  ADDFHX4 S3_8_6 ( .A(ab_8__6_), .B(CARRYB_7__6_), .CI(ab_7__7_), .CO(
        CARRYB_8__6_), .S(SUMB_8__6_) );
  ADDFHX4 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  ADDFHX4 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  ADDFHX4 S2_10_4 ( .A(ab_10__4_), .B(CARRYB_9__4_), .CI(SUMB_9__5_), .CO(
        CARRYB_10__4_), .S(SUMB_10__4_) );
  ADDFHX4 S2_8_3 ( .A(ab_8__3_), .B(CARRYB_7__3_), .CI(SUMB_7__4_), .CO(
        CARRYB_8__3_), .S(SUMB_8__3_) );
  ADDFHX4 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  ADDFHX4 S3_12_6 ( .A(ab_12__6_), .B(CARRYB_11__6_), .CI(ab_11__7_), .CO(
        CARRYB_12__6_), .S(SUMB_12__6_) );
  ADDFHX4 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  ADDFHX4 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  ADDFHX4 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  ADDFHX4 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  ADDFHX4 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  ADDFHX4 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  ADDFHX4 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  ADDFHX4 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  ADDFHX4 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  ADDFHX4 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  ADDFHX4 S2_2_3 ( .A(ab_2__3_), .B(n9), .CI(SUMB_1__4_), .CO(CARRYB_2__3_), 
        .S(SUMB_2__3_) );
  ADDFHX4 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  ADDFHX4 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  ADDFHX4 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  ADDFHX4 S2_7_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  ADDFHX4 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  ADDFHX4 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  ADDFHX4 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  ADDFHX4 S2_2_1 ( .A(ab_2__1_), .B(n8), .CI(SUMB_1__2_), .CO(CARRYB_2__1_), 
        .S(SUMB_2__1_) );
  ADDFHX4 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  ADDFHX4 S2_14_5 ( .A(ab_14__5_), .B(CARRYB_13__5_), .CI(SUMB_13__6_), .CO(
        CARRYB_14__5_), .S(SUMB_14__5_) );
  ADDFHX2 S3_14_6 ( .A(ab_14__6_), .B(CARRYB_13__6_), .CI(ab_13__7_), .CO(
        CARRYB_14__6_), .S(SUMB_14__6_) );
  ADDFHX2 S2_15_5 ( .A(ab_15__5_), .B(CARRYB_14__5_), .CI(SUMB_14__6_), .CO(
        CARRYB_15__5_), .S(SUMB_15__5_) );
  ADDFHX4 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  ADDFHX4 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  ADDFHX4 S2_7_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  ADDFHX4 S2_15_3 ( .A(ab_15__3_), .B(CARRYB_14__3_), .CI(SUMB_14__4_), .CO(
        CARRYB_15__3_), .S(SUMB_15__3_) );
  ADDFHX4 S2_7_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  ADDFHX4 S5_6 ( .A(ab_16__6_), .B(CARRYB_15__6_), .CI(ab_15__7_), .CO(
        CARRYB_16__6_), .S(SUMB_16__6_) );
  ADDFHX4 S3_11_6 ( .A(ab_11__6_), .B(CARRYB_10__6_), .CI(ab_10__7_), .CO(
        CARRYB_11__6_), .S(SUMB_11__6_) );
  ADDFHX4 S2_2_5 ( .A(ab_2__5_), .B(n3), .CI(SUMB_1__6_), .CO(CARRYB_2__5_), 
        .S(SUMB_2__5_) );
  ADDFHX4 S2_2_2 ( .A(ab_2__2_), .B(n6), .CI(SUMB_1__3_), .CO(CARRYB_2__2_), 
        .S(SUMB_2__2_) );
  ADDFHX4 S4_5 ( .A(ab_16__5_), .B(CARRYB_15__5_), .CI(SUMB_15__6_), .CO(
        CARRYB_16__5_), .S(SUMB_16__5_) );
  ADDFHX4 S3_13_6 ( .A(ab_13__6_), .B(CARRYB_12__6_), .CI(ab_12__7_), .CO(
        CARRYB_13__6_), .S(SUMB_13__6_) );
  ADDFHX2 S3_15_6 ( .A(ab_15__6_), .B(CARRYB_14__6_), .CI(ab_14__7_), .CO(
        CARRYB_15__6_), .S(SUMB_15__6_) );
  ADDFHX4 S2_15_4 ( .A(ab_15__4_), .B(CARRYB_14__4_), .CI(SUMB_14__5_), .CO(
        CARRYB_15__4_), .S(SUMB_15__4_) );
  ADDFHX4 S2_2_4 ( .A(ab_2__4_), .B(n5), .CI(SUMB_1__5_), .CO(CARRYB_2__4_), 
        .S(SUMB_2__4_) );
  ADDFHX4 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  INVX2 U2 ( .A(n34), .Y(n12) );
  INVX8 U3 ( .A(B[3]), .Y(n34) );
  NOR2BX2 U4 ( .AN(B[4]), .B(n29), .Y(ab_0__4_) );
  XOR2X4 U5 ( .A(ab_1__4_), .B(ab_0__5_), .Y(SUMB_1__4_) );
  AND2X4 U6 ( .A(ab_0__6_), .B(ab_1__5_), .Y(n3) );
  NAND2X4 U7 ( .A(CARRYB_16__1_), .B(SUMB_16__2_), .Y(n18) );
  NOR2BX1 U8 ( .AN(A[12]), .B(n23), .Y(ab_12__3_) );
  NOR2BX1 U9 ( .AN(A[9]), .B(n26), .Y(ab_9__1_) );
  NOR2BX2 U10 ( .AN(A[9]), .B(n20), .Y(ab_9__5_) );
  NOR2BXL U11 ( .AN(A[14]), .B(n23), .Y(ab_14__3_) );
  NOR2BX1 U12 ( .AN(A[9]), .B(n24), .Y(ab_9__2_) );
  NOR2BX2 U13 ( .AN(A[8]), .B(n25), .Y(ab_8__1_) );
  BUFX16 U14 ( .A(A[2]), .Y(n13) );
  NOR2BX1 U15 ( .AN(A[10]), .B(n22), .Y(ab_10__4_) );
  NOR2BX2 U16 ( .AN(A[10]), .B(n20), .Y(ab_10__5_) );
  NOR2BX1 U17 ( .AN(A[10]), .B(n23), .Y(ab_10__3_) );
  INVX4 U18 ( .A(B[4]), .Y(n33) );
  NOR2BXL U19 ( .AN(A[16]), .B(n23), .Y(ab_16__3_) );
  NOR2BX1 U20 ( .AN(A[10]), .B(n26), .Y(ab_10__1_) );
  NOR2BXL U21 ( .AN(A[16]), .B(n24), .Y(ab_16__2_) );
  NOR2BX1 U22 ( .AN(A[16]), .B(n26), .Y(ab_16__1_) );
  INVX1 U23 ( .A(n35), .Y(n11) );
  NOR2BX2 U24 ( .AN(A[5]), .B(n25), .Y(ab_5__1_) );
  AND2X4 U26 ( .A(ab_1__4_), .B(ab_0__5_), .Y(n5) );
  AND2X4 U27 ( .A(ab_1__2_), .B(ab_0__3_), .Y(n6) );
  CLKINVX8 U28 ( .A(B[2]), .Y(n35) );
  BUFX1 U29 ( .A(n35), .Y(n24) );
  AND2X4 U30 ( .A(ab_0__7_), .B(ab_1__6_), .Y(n7) );
  AND2X4 U31 ( .A(ab_0__2_), .B(n39), .Y(n8) );
  AND2X4 U32 ( .A(ab_0__4_), .B(ab_1__3_), .Y(n9) );
  CLKBUFX2 U33 ( .A(n34), .Y(n23) );
  AND2X2 U34 ( .A(CARRYB_16__5_), .B(SUMB_16__6_), .Y(n10) );
  AND2X4 U35 ( .A(n13), .B(n11), .Y(ab_2__2_) );
  NOR2BX1 U36 ( .AN(A[0]), .B(n28), .Y(n30) );
  INVX3 U37 ( .A(B[6]), .Y(n31) );
  NOR2BX4 U38 ( .AN(B[5]), .B(n29), .Y(ab_0__5_) );
  INVX4 U39 ( .A(B[5]), .Y(n32) );
  XOR2X4 U40 ( .A(ab_1__3_), .B(ab_0__4_), .Y(SUMB_1__3_) );
  BUFX16 U41 ( .A(n32), .Y(n20) );
  BUFX20 U42 ( .A(n32), .Y(n19) );
  XOR2X2 U43 ( .A(ab_1__6_), .B(ab_0__7_), .Y(SUMB_1__6_) );
  XOR2X2 U44 ( .A(n39), .B(ab_0__2_), .Y(SUMB_1__1_) );
  NOR2BX2 U45 ( .AN(A[5]), .B(n19), .Y(ab_5__5_) );
  NOR2BX4 U46 ( .AN(n13), .B(n19), .Y(ab_2__5_) );
  NOR2BX2 U47 ( .AN(A[4]), .B(n28), .Y(ab_4__0_) );
  NOR2BX4 U48 ( .AN(n13), .B(n25), .Y(ab_2__1_) );
  NOR2BX4 U49 ( .AN(n13), .B(n27), .Y(ab_2__6_) );
  AND2X4 U50 ( .A(n13), .B(n12), .Y(ab_2__3_) );
  NOR2BX4 U51 ( .AN(n13), .B(n38), .Y(ab_2__7_) );
  NOR2BX2 U52 ( .AN(A[3]), .B(n38), .Y(ab_3__7_) );
  NOR2BX2 U53 ( .AN(A[4]), .B(n38), .Y(ab_4__7_) );
  INVX20 U54 ( .A(B[7]), .Y(n38) );
  NOR2BX2 U55 ( .AN(A[3]), .B(n19), .Y(ab_3__5_) );
  XOR2X4 U56 ( .A(ab_1__5_), .B(ab_0__6_), .Y(SUMB_1__5_) );
  NOR2BX2 U57 ( .AN(A[5]), .B(n28), .Y(ab_5__0_) );
  NOR2BX2 U58 ( .AN(A[5]), .B(n24), .Y(ab_5__2_) );
  NOR2BX2 U59 ( .AN(A[5]), .B(n23), .Y(ab_5__3_) );
  NOR2BX2 U60 ( .AN(A[5]), .B(n21), .Y(ab_5__4_) );
  NOR2BX2 U61 ( .AN(A[4]), .B(n35), .Y(ab_4__2_) );
  NOR2BX2 U62 ( .AN(A[4]), .B(n34), .Y(ab_4__3_) );
  NOR2BX2 U63 ( .AN(A[4]), .B(n21), .Y(ab_4__4_) );
  NOR2BX2 U64 ( .AN(A[4]), .B(n25), .Y(ab_4__1_) );
  XOR2X4 U65 ( .A(ab_1__2_), .B(ab_0__3_), .Y(SUMB_1__2_) );
  NOR2BX4 U66 ( .AN(A[1]), .B(n35), .Y(ab_1__2_) );
  NOR2BX2 U67 ( .AN(A[3]), .B(n21), .Y(ab_3__4_) );
  NOR2BX2 U68 ( .AN(A[3]), .B(n25), .Y(ab_3__1_) );
  NOR2BX2 U69 ( .AN(A[3]), .B(n28), .Y(ab_3__0_) );
  NOR2BX2 U70 ( .AN(A[3]), .B(n27), .Y(ab_3__6_) );
  INVX4 U71 ( .A(n18), .Y(A2_17_) );
  XOR2X4 U72 ( .A(CARRYB_16__0_), .B(SUMB_16__1_), .Y(A1_15_) );
  NOR2BX2 U73 ( .AN(A[3]), .B(n35), .Y(ab_3__2_) );
  NOR2BX4 U74 ( .AN(A[1]), .B(n34), .Y(ab_1__3_) );
  NOR2BX2 U75 ( .AN(n13), .B(n28), .Y(ab_2__0_) );
  XOR2X4 U76 ( .A(CARRYB_16__5_), .B(SUMB_16__6_), .Y(A1_20_) );
  NOR2BX2 U77 ( .AN(A[5]), .B(n27), .Y(ab_5__6_) );
  AND2X4 U78 ( .A(CARRYB_16__0_), .B(SUMB_16__1_), .Y(n14) );
  NOR2BX2 U79 ( .AN(A[3]), .B(n34), .Y(ab_3__3_) );
  NOR2BX4 U80 ( .AN(n13), .B(n21), .Y(ab_2__4_) );
  BUFX20 U81 ( .A(n31), .Y(n27) );
  NOR2BX4 U82 ( .AN(B[2]), .B(n29), .Y(ab_0__2_) );
  NOR2BX4 U83 ( .AN(B[3]), .B(n29), .Y(ab_0__3_) );
  INVX12 U84 ( .A(A[0]), .Y(n29) );
  NOR2BX4 U85 ( .AN(A[1]), .B(n21), .Y(ab_1__4_) );
  NOR2BX4 U86 ( .AN(A[1]), .B(n25), .Y(n39) );
  NOR2BX4 U87 ( .AN(A[1]), .B(n19), .Y(ab_1__5_) );
  XOR2X4 U88 ( .A(SUMB_16__4_), .B(CARRYB_16__3_), .Y(A1_18_) );
  BUFX12 U89 ( .A(n36), .Y(n25) );
  AND2X4 U90 ( .A(B[6]), .B(A[1]), .Y(ab_1__6_) );
  NOR2BX2 U91 ( .AN(A[12]), .B(n28), .Y(ab_12__0_) );
  NOR2BX1 U92 ( .AN(A[14]), .B(n28), .Y(ab_14__0_) );
  NOR2BXL U93 ( .AN(A[16]), .B(n28), .Y(ab_16__0_) );
  NOR2BX2 U94 ( .AN(A[4]), .B(n27), .Y(ab_4__6_) );
  NOR2BX1 U95 ( .AN(A[12]), .B(n27), .Y(ab_12__6_) );
  AND2X2 U96 ( .A(CARRYB_16__2_), .B(SUMB_16__3_), .Y(n15) );
  NOR2BX1 U97 ( .AN(A[8]), .B(n21), .Y(ab_8__4_) );
  NOR2BX1 U98 ( .AN(A[14]), .B(n26), .Y(ab_14__1_) );
  NOR2BXL U99 ( .AN(A[6]), .B(n27), .Y(ab_6__6_) );
  NOR2BXL U100 ( .AN(A[10]), .B(n27), .Y(ab_10__6_) );
  INVX4 U101 ( .A(B[1]), .Y(n36) );
  NOR2BX1 U102 ( .AN(A[7]), .B(n21), .Y(ab_7__4_) );
  NOR2BX1 U103 ( .AN(A[8]), .B(n35), .Y(ab_8__2_) );
  NOR2BX1 U104 ( .AN(A[7]), .B(n25), .Y(ab_7__1_) );
  NOR2BX1 U105 ( .AN(A[8]), .B(n34), .Y(ab_8__3_) );
  NOR2BX1 U106 ( .AN(A[7]), .B(n19), .Y(ab_7__5_) );
  NOR2BX1 U107 ( .AN(A[12]), .B(n26), .Y(ab_12__1_) );
  NOR2BX1 U108 ( .AN(A[10]), .B(n28), .Y(ab_10__0_) );
  NOR2BX1 U109 ( .AN(A[8]), .B(n28), .Y(ab_8__0_) );
  NOR2BX1 U110 ( .AN(A[12]), .B(n24), .Y(ab_12__2_) );
  NOR2BX1 U111 ( .AN(A[12]), .B(n20), .Y(ab_12__5_) );
  NOR2BX1 U112 ( .AN(A[12]), .B(n22), .Y(ab_12__4_) );
  NOR2BX1 U113 ( .AN(A[10]), .B(n24), .Y(ab_10__2_) );
  NOR2BX1 U114 ( .AN(A[14]), .B(n24), .Y(ab_14__2_) );
  AND2X1 U115 ( .A(CARRYB_16__3_), .B(SUMB_16__4_), .Y(n16) );
  NOR2BX1 U116 ( .AN(A[14]), .B(n20), .Y(ab_14__5_) );
  NOR2BX1 U117 ( .AN(A[7]), .B(n28), .Y(ab_7__0_) );
  NOR2BX1 U118 ( .AN(A[14]), .B(n22), .Y(ab_14__4_) );
  BUFX12 U119 ( .A(n33), .Y(n21) );
  CLKBUFXL U120 ( .A(n33), .Y(n22) );
  NOR2BXL U121 ( .AN(A[11]), .B(n27), .Y(ab_11__6_) );
  NOR2BX1 U122 ( .AN(A[8]), .B(n27), .Y(ab_8__6_) );
  NOR2BX1 U123 ( .AN(A[15]), .B(n28), .Y(ab_15__0_) );
  NOR2BX1 U124 ( .AN(A[15]), .B(n24), .Y(ab_15__2_) );
  NOR2BXL U125 ( .AN(A[13]), .B(n27), .Y(ab_13__6_) );
  NOR2BXL U126 ( .AN(A[14]), .B(n27), .Y(ab_14__6_) );
  NOR2BX1 U127 ( .AN(A[15]), .B(n22), .Y(ab_15__4_) );
  BUFX3 U128 ( .A(n36), .Y(n26) );
  NOR2BX1 U129 ( .AN(A[9]), .B(n23), .Y(ab_9__3_) );
  BUFX20 U130 ( .A(n37), .Y(n28) );
  CLKINVX4 U131 ( .A(B[0]), .Y(n37) );
  NOR2BXL U132 ( .AN(A[13]), .B(n28), .Y(ab_13__0_) );
  NOR2BXL U133 ( .AN(A[13]), .B(n24), .Y(ab_13__2_) );
  NOR2BXL U134 ( .AN(A[13]), .B(n26), .Y(ab_13__1_) );
  NOR2BX1 U135 ( .AN(A[13]), .B(n23), .Y(ab_13__3_) );
  NOR2BXL U136 ( .AN(A[11]), .B(n28), .Y(ab_11__0_) );
  NOR2BX1 U137 ( .AN(A[13]), .B(n22), .Y(ab_13__4_) );
  NOR2BXL U138 ( .AN(A[6]), .B(n28), .Y(ab_6__0_) );
  NOR2BXL U139 ( .AN(A[11]), .B(n26), .Y(ab_11__1_) );
  NOR2BXL U140 ( .AN(A[11]), .B(n24), .Y(ab_11__2_) );
  NOR2BX1 U141 ( .AN(A[11]), .B(n23), .Y(ab_11__3_) );
  NOR2BXL U142 ( .AN(A[9]), .B(n28), .Y(ab_9__0_) );
  NOR2BX1 U143 ( .AN(A[11]), .B(n22), .Y(ab_11__4_) );
  NOR2BXL U144 ( .AN(A[11]), .B(n20), .Y(ab_11__5_) );
  NOR2BX1 U145 ( .AN(A[9]), .B(n22), .Y(ab_9__4_) );
  NOR2BXL U146 ( .AN(A[6]), .B(n25), .Y(ab_6__1_) );
  NOR2BX2 U147 ( .AN(A[8]), .B(n19), .Y(ab_8__5_) );
  NOR2BXL U148 ( .AN(A[7]), .B(n35), .Y(ab_7__2_) );
  NOR2BXL U149 ( .AN(A[6]), .B(n35), .Y(ab_6__2_) );
  NOR2BX1 U150 ( .AN(A[6]), .B(n34), .Y(ab_6__3_) );
  NOR2BXL U151 ( .AN(A[13]), .B(n20), .Y(ab_13__5_) );
  NOR2BX1 U152 ( .AN(A[7]), .B(n34), .Y(ab_7__3_) );
  NOR2BX2 U153 ( .AN(A[4]), .B(n19), .Y(ab_4__5_) );
  NOR2BXL U154 ( .AN(A[6]), .B(n21), .Y(ab_6__4_) );
  NOR2BXL U155 ( .AN(A[6]), .B(n19), .Y(ab_6__5_) );
  AND2X2 U156 ( .A(CARRYB_16__4_), .B(SUMB_16__5_), .Y(n17) );
  XOR2X1 U157 ( .A(CARRYB_16__6_), .B(ab_16__7_), .Y(A1_21_) );
  NOR2BX1 U158 ( .AN(A[16]), .B(n22), .Y(ab_16__4_) );
  NOR2BX1 U159 ( .AN(A[16]), .B(n20), .Y(ab_16__5_) );
  NOR2BX1 U160 ( .AN(A[15]), .B(n23), .Y(ab_15__3_) );
  NOR2BX1 U161 ( .AN(A[11]), .B(n38), .Y(ab_11__7_) );
  NOR2BXL U162 ( .AN(A[15]), .B(n20), .Y(ab_15__5_) );
  NOR2BX1 U163 ( .AN(A[12]), .B(n38), .Y(ab_12__7_) );
  NOR2BX1 U164 ( .AN(A[14]), .B(n38), .Y(ab_14__7_) );
  NOR2BX1 U165 ( .AN(A[15]), .B(n27), .Y(ab_15__6_) );
  NOR2BX1 U166 ( .AN(A[13]), .B(n38), .Y(ab_13__7_) );
  NOR2BX1 U167 ( .AN(A[9]), .B(n38), .Y(ab_9__7_) );
  NOR2BX1 U168 ( .AN(A[8]), .B(n38), .Y(ab_8__7_) );
  NOR2BX1 U169 ( .AN(A[9]), .B(n27), .Y(ab_9__6_) );
  NOR2BX1 U170 ( .AN(A[7]), .B(n38), .Y(ab_7__7_) );
  NOR2BX1 U171 ( .AN(A[6]), .B(n38), .Y(ab_6__7_) );
  NOR2BX1 U172 ( .AN(A[7]), .B(n27), .Y(ab_7__6_) );
  NOR2BX1 U173 ( .AN(A[5]), .B(n38), .Y(ab_5__7_) );
  NOR2BX1 U174 ( .AN(A[10]), .B(n38), .Y(ab_10__7_) );
  NOR2BXL U175 ( .AN(A[15]), .B(n26), .Y(ab_15__1_) );
  NOR2BX1 U176 ( .AN(A[16]), .B(n27), .Y(ab_16__6_) );
  NOR2BX1 U177 ( .AN(A[15]), .B(n38), .Y(ab_15__7_) );
  NOR2BX1 U178 ( .AN(A[16]), .B(n38), .Y(ab_16__7_) );
  XOR2X4 U179 ( .A(CARRYB_16__4_), .B(SUMB_16__5_), .Y(A1_19_) );
  XOR2X4 U180 ( .A(SUMB_16__3_), .B(CARRYB_16__2_), .Y(A1_17_) );
  XOR2X4 U181 ( .A(CARRYB_16__1_), .B(SUMB_16__2_), .Y(A1_16_) );
  AND3X1 U182 ( .A(A[1]), .B(B[1]), .C(n30), .Y(CARRYB_1__0_) );
  NOR2BXL U183 ( .AN(A[1]), .B(n38), .Y(ab_1__7_) );
  NOR2BX4 U184 ( .AN(B[7]), .B(n29), .Y(ab_0__7_) );
  NOR2BX4 U185 ( .AN(B[6]), .B(n29), .Y(ab_0__6_) );
endmodule


module multi16_5 ( in_17bit, in_8bit, out );
  input [16:0] in_17bit;
  input [7:0] in_8bit;
  output [16:0] out;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113;
  wire   [16:1] in_17bit_b;
  wire   [7:1] in_8bit_b;
  wire   [23:8] mul;

  multi16_5_DW02_mult_0 mult_55 ( .A({in_17bit_b[16:2], n35, in_17bit[0]}), 
        .B({in_8bit_b, n38}), .PRODUCT_23_(mul[23]), .PRODUCT_22_(mul[22]), 
        .PRODUCT_21_(mul[21]), .PRODUCT_20_(mul[20]), .PRODUCT_19_(mul[19]), 
        .PRODUCT_18_(mul[18]), .PRODUCT_17_(mul[17]), .PRODUCT_16_(mul[16]), 
        .PRODUCT_15_(mul[15]), .PRODUCT_14_(mul[14]), .PRODUCT_13_(mul[13]), 
        .PRODUCT_12_(mul[12]), .PRODUCT_11_(mul[11]), .PRODUCT_10_(mul[10]), 
        .PRODUCT_9_(mul[9]), .PRODUCT_8_(mul[8]), .PRODUCT_7_(out[0]) );
  NAND2X2 U2 ( .A(n9), .B(n108), .Y(n109) );
  INVX8 U3 ( .A(mul[21]), .Y(n9) );
  INVX2 U4 ( .A(mul[20]), .Y(n105) );
  INVX2 U5 ( .A(n110), .Y(n2) );
  XNOR2X4 U6 ( .A(mul[17]), .B(n1), .Y(out[10]) );
  NAND2X2 U7 ( .A(n98), .B(n102), .Y(n1) );
  NOR4X4 U8 ( .A(in_8bit[0]), .B(in_8bit[1]), .C(in_8bit[3]), .D(n3), .Y(n48)
         );
  INVX8 U9 ( .A(n44), .Y(n3) );
  NOR4X4 U10 ( .A(in_8bit[0]), .B(in_8bit[1]), .C(in_8bit[2]), .D(in_8bit[3]), 
        .Y(n7) );
  AND2X4 U11 ( .A(n106), .B(n2), .Y(n100) );
  INVX8 U12 ( .A(in_8bit[2]), .Y(n44) );
  INVX8 U13 ( .A(n6), .Y(n4) );
  NAND2X1 U14 ( .A(n39), .B(n70), .Y(n19) );
  BUFX12 U15 ( .A(n85), .Y(n6) );
  INVX3 U16 ( .A(n99), .Y(n101) );
  NAND2X2 U17 ( .A(n75), .B(n74), .Y(n76) );
  XNOR2X4 U18 ( .A(mul[13]), .B(n10), .Y(out[6]) );
  XNOR2X4 U19 ( .A(mul[16]), .B(n15), .Y(out[9]) );
  NAND2X4 U20 ( .A(n99), .B(n102), .Y(n14) );
  AND2X1 U21 ( .A(n39), .B(n64), .Y(n31) );
  INVX2 U22 ( .A(n109), .Y(n112) );
  NAND2X4 U23 ( .A(n109), .B(n102), .Y(n5) );
  AND2X2 U24 ( .A(n39), .B(n60), .Y(n17) );
  INVX4 U25 ( .A(in_8bit[5]), .Y(n49) );
  OAI21X2 U26 ( .A0(in_8bit[1]), .A1(in_8bit[0]), .B0(n40), .Y(n45) );
  AND2X1 U27 ( .A(in_8bit[0]), .B(n40), .Y(n26) );
  XOR2X4 U28 ( .A(n5), .B(n111), .Y(out[15]) );
  BUFX12 U29 ( .A(in_17bit[16]), .Y(n39) );
  XNOR2X4 U30 ( .A(n107), .B(n9), .Y(out[14]) );
  NOR2X4 U31 ( .A(n28), .B(n6), .Y(n18) );
  NOR2X2 U32 ( .A(n69), .B(n6), .Y(n67) );
  NOR2X1 U33 ( .A(n75), .B(n6), .Y(n73) );
  NOR2X4 U34 ( .A(n33), .B(n41), .Y(n20) );
  NAND3BX2 U35 ( .AN(in_8bit[0]), .B(n44), .C(n43), .Y(n36) );
  NOR2X2 U36 ( .A(n41), .B(n48), .Y(n46) );
  INVX2 U37 ( .A(in_8bit[1]), .Y(n43) );
  CLKINVX8 U38 ( .A(n42), .Y(n40) );
  NAND2X4 U39 ( .A(n94), .B(n102), .Y(n16) );
  NOR2X4 U40 ( .A(in_17bit[1]), .B(in_17bit[0]), .Y(n8) );
  INVX4 U41 ( .A(in_17bit[0]), .Y(n55) );
  XOR2X2 U42 ( .A(n113), .B(mul[23]), .Y(out[16]) );
  OAI22X4 U43 ( .A0(in_17bit[0]), .A1(in_17bit[1]), .B0(n39), .B1(in_17bit[1]), 
        .Y(n53) );
  CLKINVX8 U44 ( .A(in_17bit[4]), .Y(n59) );
  XNOR2X4 U45 ( .A(n20), .B(n49), .Y(in_8bit_b[5]) );
  AOI21X4 U46 ( .A0(n54), .A1(n39), .B0(n53), .Y(in_17bit_b[1]) );
  BUFX16 U47 ( .A(in_17bit_b[1]), .Y(n35) );
  AOI21X1 U48 ( .A0(n112), .A1(n111), .B0(n110), .Y(n113) );
  CLKINVX8 U49 ( .A(in_17bit[2]), .Y(n57) );
  NOR2X4 U50 ( .A(n8), .B(n85), .Y(n56) );
  NAND2X4 U51 ( .A(n28), .B(n63), .Y(n64) );
  XNOR2X4 U52 ( .A(n65), .B(n31), .Y(in_17bit_b[7]) );
  NOR2BX4 U53 ( .AN(in_17bit[1]), .B(n55), .Y(n54) );
  NAND2X2 U54 ( .A(n52), .B(n40), .Y(n51) );
  AND2X4 U55 ( .A(n40), .B(n36), .Y(n24) );
  INVX4 U56 ( .A(in_8bit[7]), .Y(n41) );
  XOR2X4 U57 ( .A(n27), .B(n59), .Y(in_17bit_b[4]) );
  AND2X4 U58 ( .A(n39), .B(n58), .Y(n23) );
  XOR2X4 U59 ( .A(in_17bit[3]), .B(n23), .Y(in_17bit_b[3]) );
  XNOR2X2 U60 ( .A(mul[11]), .B(n11), .Y(out[4]) );
  INVX8 U61 ( .A(mul[22]), .Y(n111) );
  NAND2X2 U62 ( .A(n92), .B(n102), .Y(n91) );
  NAND2BX4 U63 ( .AN(mul[18]), .B(n101), .Y(n103) );
  NAND2X2 U64 ( .A(n32), .B(n59), .Y(n60) );
  NOR2X2 U65 ( .A(in_17bit[3]), .B(n58), .Y(n32) );
  NOR2X4 U66 ( .A(n108), .B(n110), .Y(n107) );
  XNOR2X4 U67 ( .A(mul[15]), .B(n12), .Y(out[8]) );
  NAND2X4 U68 ( .A(n95), .B(n102), .Y(n12) );
  XOR2X4 U69 ( .A(n24), .B(in_8bit[3]), .Y(in_8bit_b[3]) );
  NAND2X2 U70 ( .A(n93), .B(n102), .Y(n10) );
  XNOR2X2 U71 ( .A(n26), .B(n43), .Y(in_8bit_b[1]) );
  XOR2X2 U72 ( .A(mul[9]), .B(n25), .Y(out[2]) );
  INVX8 U73 ( .A(in_8bit[7]), .Y(n42) );
  XNOR2X4 U74 ( .A(mul[18]), .B(n14), .Y(out[11]) );
  NOR3X4 U75 ( .A(mul[19]), .B(mul[20]), .C(n106), .Y(n108) );
  XNOR2X4 U76 ( .A(mul[14]), .B(n16), .Y(out[7]) );
  OR2X4 U77 ( .A(n32), .B(n85), .Y(n27) );
  NAND2X2 U78 ( .A(n97), .B(n102), .Y(n15) );
  NAND2XL U79 ( .A(n90), .B(n102), .Y(n11) );
  NAND2X4 U80 ( .A(n57), .B(n8), .Y(n58) );
  XNOR2X4 U81 ( .A(n18), .B(n63), .Y(in_17bit_b[6]) );
  XOR2X2 U82 ( .A(n77), .B(n22), .Y(in_17bit_b[11]) );
  NAND2X2 U83 ( .A(n29), .B(n84), .Y(n86) );
  OR2X4 U84 ( .A(mul[10]), .B(n89), .Y(n90) );
  OR2X4 U85 ( .A(mul[17]), .B(n98), .Y(n99) );
  XOR2X1 U86 ( .A(mul[8]), .B(n13), .Y(out[1]) );
  AND2X2 U87 ( .A(out[0]), .B(n102), .Y(n13) );
  OR2X4 U88 ( .A(mul[9]), .B(n87), .Y(n89) );
  OR2X4 U89 ( .A(mul[14]), .B(n94), .Y(n95) );
  OR2X4 U90 ( .A(mul[13]), .B(n93), .Y(n94) );
  OR2X4 U91 ( .A(mul[12]), .B(n92), .Y(n93) );
  OR2X4 U92 ( .A(mul[8]), .B(out[0]), .Y(n87) );
  INVX4 U93 ( .A(n110), .Y(n102) );
  XNOR2X4 U94 ( .A(n61), .B(n17), .Y(in_17bit_b[5]) );
  AND2X4 U95 ( .A(n62), .B(n61), .Y(n28) );
  XOR2X2 U96 ( .A(n71), .B(n19), .Y(in_17bit_b[9]) );
  NAND2BXL U97 ( .AN(n64), .B(n65), .Y(n66) );
  XOR2X2 U98 ( .A(n82), .B(n21), .Y(in_17bit_b[13]) );
  NAND2XL U99 ( .A(n4), .B(n81), .Y(n21) );
  NAND2XL U100 ( .A(n4), .B(n76), .Y(n22) );
  NOR2XL U101 ( .A(n81), .B(in_17bit[13]), .Y(n29) );
  NAND2BXL U102 ( .AN(n70), .B(n71), .Y(n72) );
  AND2X4 U103 ( .A(n78), .B(n77), .Y(n30) );
  AND2X4 U104 ( .A(n7), .B(n47), .Y(n33) );
  INVXL U105 ( .A(in_17bit[11]), .Y(n77) );
  OR2X2 U106 ( .A(mul[11]), .B(n90), .Y(n92) );
  OR2X4 U107 ( .A(mul[16]), .B(n97), .Y(n98) );
  AND2X2 U108 ( .A(n87), .B(n102), .Y(n25) );
  XOR2X4 U109 ( .A(n100), .B(mul[19]), .Y(out[12]) );
  INVXL U110 ( .A(in_8bit[0]), .Y(n37) );
  NOR2XL U111 ( .A(n29), .B(n6), .Y(n83) );
  NOR2XL U112 ( .A(n30), .B(n6), .Y(n79) );
  XNOR2X1 U113 ( .A(n39), .B(n40), .Y(n110) );
  XOR2X2 U114 ( .A(in_17bit[15]), .B(n34), .Y(in_17bit_b[15]) );
  AND2X1 U115 ( .A(n4), .B(n86), .Y(n34) );
  INVX1 U116 ( .A(in_17bit[5]), .Y(n61) );
  INVX1 U117 ( .A(in_8bit[6]), .Y(n50) );
  INVX1 U118 ( .A(in_8bit[4]), .Y(n47) );
  INVX2 U119 ( .A(n37), .Y(n38) );
  INVX8 U120 ( .A(n39), .Y(n85) );
  XOR2X4 U121 ( .A(n45), .B(n44), .Y(in_8bit_b[2]) );
  XNOR2X4 U122 ( .A(n46), .B(n47), .Y(in_8bit_b[4]) );
  NAND2X4 U123 ( .A(n33), .B(n49), .Y(n52) );
  XOR2X4 U124 ( .A(n51), .B(n50), .Y(in_8bit_b[6]) );
  NOR3X4 U125 ( .A(in_8bit[6]), .B(n52), .C(n42), .Y(in_8bit_b[7]) );
  XNOR2X4 U126 ( .A(n56), .B(n57), .Y(in_17bit_b[2]) );
  CLKINVX3 U127 ( .A(n60), .Y(n62) );
  CLKINVX3 U128 ( .A(in_17bit[6]), .Y(n63) );
  CLKINVX3 U129 ( .A(in_17bit[7]), .Y(n65) );
  CLKINVX3 U130 ( .A(n66), .Y(n69) );
  CLKINVX3 U131 ( .A(in_17bit[8]), .Y(n68) );
  XNOR2X4 U132 ( .A(n67), .B(n68), .Y(in_17bit_b[8]) );
  CLKINVX3 U133 ( .A(in_17bit[9]), .Y(n71) );
  NAND2X4 U134 ( .A(n69), .B(n68), .Y(n70) );
  CLKINVX3 U135 ( .A(n72), .Y(n75) );
  CLKINVX3 U136 ( .A(in_17bit[10]), .Y(n74) );
  XNOR2X4 U137 ( .A(n73), .B(n74), .Y(in_17bit_b[10]) );
  CLKINVX3 U138 ( .A(n76), .Y(n78) );
  CLKINVX3 U139 ( .A(in_17bit[12]), .Y(n80) );
  XNOR2X4 U140 ( .A(n79), .B(n80), .Y(in_17bit_b[12]) );
  CLKINVX3 U141 ( .A(in_17bit[13]), .Y(n82) );
  NAND2X4 U142 ( .A(n30), .B(n80), .Y(n81) );
  CLKINVX3 U143 ( .A(in_17bit[14]), .Y(n84) );
  XNOR2X4 U144 ( .A(n83), .B(n84), .Y(in_17bit_b[14]) );
  NOR3X4 U145 ( .A(in_17bit[15]), .B(n86), .C(n6), .Y(in_17bit_b[16]) );
  NAND2X4 U146 ( .A(n89), .B(n102), .Y(n88) );
  XNOR2X4 U147 ( .A(mul[10]), .B(n88), .Y(out[3]) );
  XNOR2X4 U148 ( .A(mul[12]), .B(n91), .Y(out[5]) );
  CLKINVX3 U149 ( .A(n95), .Y(n96) );
  NAND2BX4 U150 ( .AN(mul[15]), .B(n96), .Y(n97) );
  NAND2BX4 U151 ( .AN(mul[18]), .B(n101), .Y(n106) );
  OAI21X4 U152 ( .A0(mul[19]), .A1(n103), .B0(n102), .Y(n104) );
  XOR2X4 U153 ( .A(n104), .B(n105), .Y(out[13]) );
endmodule


module multi16_4_DW01_add_0 ( A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, 
        A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, 
        B_20_, B_19_, B_18_, B_17_, B_16_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, 
        SUM_17_, SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, 
        SUM_9_, SUM_8_, SUM_7_, SUM_6_, SUM_5_ );
  input A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_,
         A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, B_20_, B_19_,
         B_18_, B_17_, B_16_;
  output SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, SUM_15_,
         SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, SUM_7_,
         SUM_6_, SUM_5_;
  wire   n49, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48;

  CLKINVX8 U2 ( .A(n28), .Y(n7) );
  BUFX12 U3 ( .A(n49), .Y(SUM_18_) );
  INVX8 U4 ( .A(n6), .Y(n5) );
  OR2X4 U5 ( .A(B_16_), .B(A_16_), .Y(n47) );
  INVX3 U6 ( .A(n37), .Y(n27) );
  INVXL U7 ( .A(n2), .Y(n3) );
  AND2X4 U8 ( .A(B_19_), .B(A_19_), .Y(n2) );
  BUFX8 U9 ( .A(A_6_), .Y(SUM_6_) );
  NAND2X4 U10 ( .A(n4), .B(n3), .Y(n32) );
  OR2X4 U11 ( .A(n35), .B(n36), .Y(n4) );
  INVX8 U12 ( .A(n26), .Y(n6) );
  AOI21X2 U13 ( .A0(n32), .A1(n33), .B0(n23), .Y(n31) );
  XOR2X2 U14 ( .A(n30), .B(n31), .Y(SUM_21_) );
  OR2X4 U15 ( .A(B_20_), .B(A_20_), .Y(n33) );
  NAND2BX4 U16 ( .AN(n7), .B(n8), .Y(n9) );
  BUFX8 U17 ( .A(A_8_), .Y(SUM_8_) );
  NOR2X4 U18 ( .A(n2), .B(n36), .Y(n44) );
  OAI21X1 U19 ( .A0(n37), .A1(n41), .B0(n6), .Y(n39) );
  BUFX12 U20 ( .A(A_11_), .Y(SUM_11_) );
  INVX8 U21 ( .A(n41), .Y(n28) );
  INVX8 U22 ( .A(n29), .Y(SUM_15_) );
  NAND2X4 U23 ( .A(n40), .B(n24), .Y(n46) );
  BUFX12 U24 ( .A(A_14_), .Y(SUM_14_) );
  AOI21X2 U25 ( .A0(n24), .A1(n39), .B0(n25), .Y(n35) );
  XOR2X4 U26 ( .A(n32), .B(n12), .Y(SUM_20_) );
  OAI21X2 U27 ( .A0(n45), .A1(n38), .B0(n40), .Y(n43) );
  XOR2X4 U28 ( .A(n43), .B(n44), .Y(SUM_19_) );
  NAND2X4 U29 ( .A(B_18_), .B(A_18_), .Y(n40) );
  BUFX12 U30 ( .A(A_13_), .Y(SUM_13_) );
  INVX8 U31 ( .A(n48), .Y(SUM_16_) );
  NAND2X2 U32 ( .A(n11), .B(n7), .Y(n10) );
  NAND2X4 U33 ( .A(n9), .B(n10), .Y(SUM_17_) );
  INVX4 U34 ( .A(n11), .Y(n8) );
  NOR2X4 U35 ( .A(n26), .B(n37), .Y(n11) );
  INVX4 U36 ( .A(n38), .Y(n24) );
  NOR2X2 U37 ( .A(B_19_), .B(A_19_), .Y(n36) );
  AND2X2 U38 ( .A(n34), .B(n33), .Y(n12) );
  INVXL U39 ( .A(n40), .Y(n25) );
  NAND2X4 U40 ( .A(n47), .B(n41), .Y(n48) );
  INVXL U41 ( .A(n34), .Y(n23) );
  BUFX8 U42 ( .A(A_12_), .Y(SUM_12_) );
  BUFX8 U43 ( .A(A_5_), .Y(SUM_5_) );
  BUFX8 U44 ( .A(A_10_), .Y(SUM_10_) );
  BUFX8 U45 ( .A(A_9_), .Y(SUM_9_) );
  BUFX4 U46 ( .A(A_7_), .Y(SUM_7_) );
  AOI21X4 U47 ( .A0(n27), .A1(n28), .B0(n5), .Y(n45) );
  CLKINVX8 U48 ( .A(A_15_), .Y(n29) );
  INVX8 U49 ( .A(n42), .Y(n26) );
  NAND2X4 U50 ( .A(B_16_), .B(A_16_), .Y(n41) );
  NOR2X4 U51 ( .A(B_18_), .B(A_18_), .Y(n38) );
  NOR2X4 U52 ( .A(A_17_), .B(B_17_), .Y(n37) );
  NAND2X4 U53 ( .A(A_17_), .B(B_17_), .Y(n42) );
  XOR2X4 U54 ( .A(n45), .B(n46), .Y(n49) );
  XNOR2X1 U55 ( .A(B_21_), .B(A_21_), .Y(n30) );
  NAND2X1 U56 ( .A(B_20_), .B(A_20_), .Y(n34) );
endmodule


module multi16_4_DW02_mult_0 ( A, B, PRODUCT_23_, PRODUCT_22_, PRODUCT_21_, 
        PRODUCT_20_, PRODUCT_19_, PRODUCT_18_, PRODUCT_17_, PRODUCT_16_, 
        PRODUCT_15_, PRODUCT_14_, PRODUCT_13_, PRODUCT_12_, PRODUCT_11_, 
        PRODUCT_10_, PRODUCT_9_, PRODUCT_8_, PRODUCT_7_ );
  input [16:0] A;
  input [7:0] B;
  output PRODUCT_23_, PRODUCT_22_, PRODUCT_21_, PRODUCT_20_, PRODUCT_19_,
         PRODUCT_18_, PRODUCT_17_, PRODUCT_16_, PRODUCT_15_, PRODUCT_14_,
         PRODUCT_13_, PRODUCT_12_, PRODUCT_11_, PRODUCT_10_, PRODUCT_9_,
         PRODUCT_8_, PRODUCT_7_;
  wire   ab_16__7_, ab_16__6_, ab_16__5_, ab_16__4_, ab_16__3_, ab_16__2_,
         ab_16__1_, ab_16__0_, ab_15__7_, ab_15__6_, ab_15__5_, ab_15__4_,
         ab_15__3_, ab_15__2_, ab_15__1_, ab_15__0_, ab_14__7_, ab_14__6_,
         ab_14__5_, ab_14__4_, ab_14__3_, ab_14__2_, ab_14__1_, ab_14__0_,
         ab_13__7_, ab_13__6_, ab_13__5_, ab_13__4_, ab_13__3_, ab_13__2_,
         ab_13__1_, ab_13__0_, ab_12__7_, ab_12__6_, ab_12__5_, ab_12__4_,
         ab_12__3_, ab_12__2_, ab_12__1_, ab_12__0_, ab_11__7_, ab_11__6_,
         ab_11__5_, ab_11__4_, ab_11__3_, ab_11__2_, ab_11__1_, ab_11__0_,
         ab_10__7_, ab_10__6_, ab_10__5_, ab_10__4_, ab_10__3_, ab_10__2_,
         ab_10__1_, ab_10__0_, ab_9__7_, ab_9__6_, ab_9__5_, ab_9__4_,
         ab_9__3_, ab_9__2_, ab_9__1_, ab_9__0_, ab_8__7_, ab_8__6_, ab_8__5_,
         ab_8__4_, ab_8__3_, ab_8__2_, ab_8__1_, ab_8__0_, ab_7__7_, ab_7__6_,
         ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_, ab_7__0_, ab_6__7_,
         ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_, ab_6__1_, ab_6__0_,
         ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_, ab_5__2_, ab_5__1_,
         ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_, ab_4__3_, ab_4__2_,
         ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_, ab_3__4_, ab_3__3_,
         ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_, ab_2__5_, ab_2__4_,
         ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_, ab_1__6_, ab_1__5_,
         ab_1__4_, ab_1__3_, ab_1__2_, ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_,
         ab_0__3_, ab_0__2_, CARRYB_16__6_, CARRYB_16__5_, CARRYB_16__4_,
         CARRYB_16__3_, CARRYB_16__2_, CARRYB_16__1_, CARRYB_16__0_,
         CARRYB_15__6_, CARRYB_15__5_, CARRYB_15__4_, CARRYB_15__3_,
         CARRYB_15__2_, CARRYB_15__1_, CARRYB_15__0_, CARRYB_14__6_,
         CARRYB_14__5_, CARRYB_14__4_, CARRYB_14__3_, CARRYB_14__2_,
         CARRYB_14__1_, CARRYB_14__0_, CARRYB_13__6_, CARRYB_13__5_,
         CARRYB_13__4_, CARRYB_13__3_, CARRYB_13__2_, CARRYB_13__1_,
         CARRYB_13__0_, CARRYB_12__6_, CARRYB_12__5_, CARRYB_12__4_,
         CARRYB_12__3_, CARRYB_12__2_, CARRYB_12__1_, CARRYB_12__0_,
         CARRYB_11__6_, CARRYB_11__5_, CARRYB_11__4_, CARRYB_11__3_,
         CARRYB_11__2_, CARRYB_11__1_, CARRYB_11__0_, CARRYB_10__6_,
         CARRYB_10__5_, CARRYB_10__4_, CARRYB_10__3_, CARRYB_10__2_,
         CARRYB_10__1_, CARRYB_10__0_, CARRYB_9__6_, CARRYB_9__5_,
         CARRYB_9__4_, CARRYB_9__3_, CARRYB_9__2_, CARRYB_9__1_, CARRYB_9__0_,
         CARRYB_8__6_, CARRYB_8__5_, CARRYB_8__4_, CARRYB_8__3_, CARRYB_8__2_,
         CARRYB_8__1_, CARRYB_8__0_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_,
         CARRYB_7__3_, CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_,
         CARRYB_6__5_, CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_,
         CARRYB_6__0_, CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_,
         CARRYB_5__2_, CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_,
         CARRYB_4__4_, CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_,
         CARRYB_3__6_, CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_,
         CARRYB_3__1_, CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_,
         CARRYB_2__3_, CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__0_,
         SUMB_16__6_, SUMB_16__5_, SUMB_16__4_, SUMB_16__3_, SUMB_16__2_,
         SUMB_16__1_, SUMB_16__0_, SUMB_15__6_, SUMB_15__5_, SUMB_15__4_,
         SUMB_15__3_, SUMB_15__2_, SUMB_15__1_, SUMB_14__6_, SUMB_14__5_,
         SUMB_14__4_, SUMB_14__3_, SUMB_14__2_, SUMB_14__1_, SUMB_13__6_,
         SUMB_13__5_, SUMB_13__4_, SUMB_13__3_, SUMB_13__2_, SUMB_13__1_,
         SUMB_12__6_, SUMB_12__5_, SUMB_12__4_, SUMB_12__3_, SUMB_12__2_,
         SUMB_12__1_, SUMB_11__6_, SUMB_11__5_, SUMB_11__4_, SUMB_11__3_,
         SUMB_11__2_, SUMB_11__1_, SUMB_10__6_, SUMB_10__5_, SUMB_10__4_,
         SUMB_10__3_, SUMB_10__2_, SUMB_10__1_, SUMB_9__6_, SUMB_9__5_,
         SUMB_9__4_, SUMB_9__3_, SUMB_9__2_, SUMB_9__1_, SUMB_8__6_,
         SUMB_8__5_, SUMB_8__4_, SUMB_8__3_, SUMB_8__2_, SUMB_8__1_,
         SUMB_7__6_, SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_,
         SUMB_7__1_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, PROD1_7_, A1_21_, A1_20_, A1_19_, A1_18_,
         A1_17_, A1_16_, A1_15_, A1_13_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_,
         A1_7_, A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, n3, n4, n5, n6, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47;

  multi16_4_DW01_add_0 FS_1 ( .A_21_(A1_21_), .A_20_(A1_20_), .A_19_(A1_19_), 
        .A_18_(A1_18_), .A_17_(A1_17_), .A_16_(A1_16_), .A_15_(A1_15_), 
        .A_14_(SUMB_16__0_), .A_13_(A1_13_), .A_12_(A1_12_), .A_11_(A1_11_), 
        .A_10_(A1_10_), .A_9_(A1_9_), .A_8_(A1_8_), .A_7_(A1_7_), .A_6_(A1_6_), 
        .A_5_(PROD1_7_), .B_21_(n26), .B_20_(n25), .B_19_(n24), .B_18_(n22), 
        .B_17_(n12), .B_16_(n23), .SUM_21_(PRODUCT_23_), .SUM_20_(PRODUCT_22_), 
        .SUM_19_(PRODUCT_21_), .SUM_18_(PRODUCT_20_), .SUM_17_(PRODUCT_19_), 
        .SUM_16_(PRODUCT_18_), .SUM_15_(PRODUCT_17_), .SUM_14_(PRODUCT_16_), 
        .SUM_13_(PRODUCT_15_), .SUM_12_(PRODUCT_14_), .SUM_11_(PRODUCT_13_), 
        .SUM_10_(PRODUCT_12_), .SUM_9_(PRODUCT_11_), .SUM_8_(PRODUCT_10_), 
        .SUM_7_(PRODUCT_9_), .SUM_6_(PRODUCT_8_), .SUM_5_(PRODUCT_7_) );
  ADDFHX4 S2_10_4 ( .A(ab_10__4_), .B(CARRYB_9__4_), .CI(SUMB_9__5_), .CO(
        CARRYB_10__4_), .S(SUMB_10__4_) );
  ADDFHX4 S2_11_4 ( .A(ab_11__4_), .B(CARRYB_10__4_), .CI(SUMB_10__5_), .CO(
        CARRYB_11__4_), .S(SUMB_11__4_) );
  ADDFHX4 S2_12_3 ( .A(ab_12__3_), .B(CARRYB_11__3_), .CI(SUMB_11__4_), .CO(
        CARRYB_12__3_), .S(SUMB_12__3_) );
  ADDFHX4 S2_12_2 ( .A(ab_12__2_), .B(CARRYB_11__2_), .CI(SUMB_11__3_), .CO(
        CARRYB_12__2_), .S(SUMB_12__2_) );
  ADDFHX4 S2_13_2 ( .A(ab_13__2_), .B(CARRYB_12__2_), .CI(SUMB_12__3_), .CO(
        CARRYB_13__2_), .S(SUMB_13__2_) );
  ADDFHX4 S4_1 ( .A(ab_16__1_), .B(CARRYB_15__1_), .CI(SUMB_15__2_), .CO(
        CARRYB_16__1_), .S(SUMB_16__1_) );
  ADDFHX4 S4_2 ( .A(ab_16__2_), .B(CARRYB_15__2_), .CI(SUMB_15__3_), .CO(
        CARRYB_16__2_), .S(SUMB_16__2_) );
  ADDFHX4 S2_11_2 ( .A(ab_11__2_), .B(CARRYB_10__2_), .CI(SUMB_10__3_), .CO(
        CARRYB_11__2_), .S(SUMB_11__2_) );
  ADDFHX4 S2_14_3 ( .A(ab_14__3_), .B(CARRYB_13__3_), .CI(SUMB_13__4_), .CO(
        CARRYB_14__3_), .S(SUMB_14__3_) );
  ADDFHX4 S2_13_3 ( .A(ab_13__3_), .B(CARRYB_12__3_), .CI(SUMB_12__4_), .CO(
        CARRYB_13__3_), .S(SUMB_13__3_) );
  ADDFHX4 S2_14_1 ( .A(ab_14__1_), .B(CARRYB_13__1_), .CI(SUMB_13__2_), .CO(
        CARRYB_14__1_), .S(SUMB_14__1_) );
  ADDFHX4 S2_13_1 ( .A(ab_13__1_), .B(SUMB_12__2_), .CI(CARRYB_12__1_), .CO(
        CARRYB_13__1_), .S(SUMB_13__1_) );
  ADDFHX4 S2_10_2 ( .A(ab_10__2_), .B(CARRYB_9__2_), .CI(SUMB_9__3_), .CO(
        CARRYB_10__2_), .S(SUMB_10__2_) );
  ADDFHX4 S1_10_0 ( .A(ab_10__0_), .B(SUMB_9__1_), .CI(CARRYB_9__0_), .CO(
        CARRYB_10__0_), .S(A1_8_) );
  ADDFHX4 S1_12_0 ( .A(ab_12__0_), .B(CARRYB_11__0_), .CI(SUMB_11__1_), .CO(
        CARRYB_12__0_), .S(A1_10_) );
  ADDFHX4 S1_13_0 ( .A(ab_13__0_), .B(CARRYB_12__0_), .CI(SUMB_12__1_), .CO(
        CARRYB_13__0_), .S(A1_11_) );
  ADDFHX4 S4_4 ( .A(ab_16__4_), .B(CARRYB_15__4_), .CI(SUMB_15__5_), .CO(
        CARRYB_16__4_), .S(SUMB_16__4_) );
  ADDFHX4 S2_11_1 ( .A(ab_11__1_), .B(CARRYB_10__1_), .CI(SUMB_10__2_), .CO(
        CARRYB_11__1_), .S(SUMB_11__1_) );
  ADDFHX4 S2_14_2 ( .A(ab_14__2_), .B(CARRYB_13__2_), .CI(SUMB_13__3_), .CO(
        CARRYB_14__2_), .S(SUMB_14__2_) );
  ADDFHX4 S2_13_5 ( .A(ab_13__5_), .B(CARRYB_12__5_), .CI(SUMB_12__6_), .CO(
        CARRYB_13__5_), .S(SUMB_13__5_) );
  ADDFHX4 S4_0 ( .A(ab_16__0_), .B(SUMB_15__1_), .CI(CARRYB_15__0_), .CO(
        CARRYB_16__0_), .S(SUMB_16__0_) );
  ADDFHX4 S1_14_0 ( .A(ab_14__0_), .B(CARRYB_13__0_), .CI(SUMB_13__1_), .CO(
        CARRYB_14__0_), .S(A1_12_) );
  ADDFHX4 S1_15_0 ( .A(ab_15__0_), .B(CARRYB_14__0_), .CI(SUMB_14__1_), .CO(
        CARRYB_15__0_), .S(A1_13_) );
  ADDFHX4 S2_13_4 ( .A(ab_13__4_), .B(CARRYB_12__4_), .CI(SUMB_12__5_), .CO(
        CARRYB_13__4_), .S(SUMB_13__4_) );
  ADDFHX4 S2_14_4 ( .A(ab_14__4_), .B(CARRYB_13__4_), .CI(SUMB_13__5_), .CO(
        CARRYB_14__4_), .S(SUMB_14__4_) );
  ADDFHX4 S2_10_3 ( .A(ab_10__3_), .B(CARRYB_9__3_), .CI(SUMB_9__4_), .CO(
        CARRYB_10__3_), .S(SUMB_10__3_) );
  ADDFHX4 S1_7_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(PROD1_7_) );
  ADDFHX4 S1_8_0 ( .A(ab_8__0_), .B(CARRYB_7__0_), .CI(SUMB_7__1_), .CO(
        CARRYB_8__0_), .S(A1_6_) );
  ADDFHX4 S1_11_0 ( .A(ab_11__0_), .B(CARRYB_10__0_), .CI(SUMB_10__1_), .CO(
        CARRYB_11__0_), .S(A1_9_) );
  ADDFHX4 S2_12_5 ( .A(ab_12__5_), .B(CARRYB_11__5_), .CI(SUMB_11__6_), .CO(
        CARRYB_12__5_), .S(SUMB_12__5_) );
  ADDFHX4 S2_11_5 ( .A(ab_11__5_), .B(CARRYB_10__5_), .CI(SUMB_10__6_), .CO(
        CARRYB_11__5_), .S(SUMB_11__5_) );
  ADDFHX4 S2_15_2 ( .A(ab_15__2_), .B(CARRYB_14__2_), .CI(SUMB_14__3_), .CO(
        CARRYB_15__2_), .S(SUMB_15__2_) );
  ADDFHX4 S2_15_3 ( .A(ab_15__3_), .B(CARRYB_14__3_), .CI(SUMB_14__4_), .CO(
        CARRYB_15__3_), .S(SUMB_15__3_) );
  ADDFHX4 S2_12_4 ( .A(ab_12__4_), .B(CARRYB_11__4_), .CI(SUMB_11__5_), .CO(
        CARRYB_12__4_), .S(SUMB_12__4_) );
  ADDFHX4 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  ADDFHX4 S2_11_3 ( .A(ab_11__3_), .B(CARRYB_10__3_), .CI(SUMB_10__4_), .CO(
        CARRYB_11__3_), .S(SUMB_11__3_) );
  ADDFHX4 S4_5 ( .A(ab_16__5_), .B(CARRYB_15__5_), .CI(SUMB_15__6_), .CO(
        CARRYB_16__5_), .S(SUMB_16__5_) );
  ADDFHX4 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  ADDFHX4 S2_9_4 ( .A(ab_9__4_), .B(CARRYB_8__4_), .CI(SUMB_8__5_), .CO(
        CARRYB_9__4_), .S(SUMB_9__4_) );
  ADDFHX4 S3_14_6 ( .A(ab_14__6_), .B(CARRYB_13__6_), .CI(ab_13__7_), .CO(
        CARRYB_14__6_), .S(SUMB_14__6_) );
  ADDFHX4 S2_15_5 ( .A(ab_15__5_), .B(CARRYB_14__5_), .CI(SUMB_14__6_), .CO(
        CARRYB_15__5_), .S(SUMB_15__5_) );
  ADDFHX4 S3_10_6 ( .A(ab_10__6_), .B(CARRYB_9__6_), .CI(ab_9__7_), .CO(
        CARRYB_10__6_), .S(SUMB_10__6_) );
  ADDFHX4 S2_9_2 ( .A(ab_9__2_), .B(CARRYB_8__2_), .CI(SUMB_8__3_), .CO(
        CARRYB_9__2_), .S(SUMB_9__2_) );
  ADDFHX4 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  ADDFHX4 S2_10_5 ( .A(ab_10__5_), .B(CARRYB_9__5_), .CI(SUMB_9__6_), .CO(
        CARRYB_10__5_), .S(SUMB_10__5_) );
  ADDFHX4 S2_15_1 ( .A(ab_15__1_), .B(CARRYB_14__1_), .CI(SUMB_14__2_), .CO(
        CARRYB_15__1_), .S(SUMB_15__1_) );
  ADDFHX4 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  ADDFHX4 S2_8_5 ( .A(ab_8__5_), .B(CARRYB_7__5_), .CI(SUMB_7__6_), .CO(
        CARRYB_8__5_), .S(SUMB_8__5_) );
  ADDFHX4 S2_9_5 ( .A(ab_9__5_), .B(CARRYB_8__5_), .CI(SUMB_8__6_), .CO(
        CARRYB_9__5_), .S(SUMB_9__5_) );
  ADDFHX4 S2_8_3 ( .A(ab_8__3_), .B(CARRYB_7__3_), .CI(SUMB_7__4_), .CO(
        CARRYB_8__3_), .S(SUMB_8__3_) );
  ADDFHX4 S2_9_3 ( .A(ab_9__3_), .B(CARRYB_8__3_), .CI(SUMB_8__4_), .CO(
        CARRYB_9__3_), .S(SUMB_9__3_) );
  ADDFHX4 S2_7_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  ADDFHX4 S3_8_6 ( .A(ab_8__6_), .B(CARRYB_7__6_), .CI(ab_7__7_), .CO(
        CARRYB_8__6_), .S(SUMB_8__6_) );
  ADDFHX4 S3_9_6 ( .A(ab_9__6_), .B(CARRYB_8__6_), .CI(ab_8__7_), .CO(
        CARRYB_9__6_), .S(SUMB_9__6_) );
  ADDFHX4 S4_3 ( .A(ab_16__3_), .B(CARRYB_15__3_), .CI(SUMB_15__4_), .CO(
        CARRYB_16__3_), .S(SUMB_16__3_) );
  ADDFHX4 S2_8_2 ( .A(ab_8__2_), .B(CARRYB_7__2_), .CI(SUMB_7__3_), .CO(
        CARRYB_8__2_), .S(SUMB_8__2_) );
  ADDFHX4 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  ADDFHX4 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  ADDFHX4 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  ADDFHX4 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  ADDFHX4 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  ADDFHX4 S2_8_4 ( .A(ab_8__4_), .B(CARRYB_7__4_), .CI(SUMB_7__5_), .CO(
        CARRYB_8__4_), .S(SUMB_8__4_) );
  ADDFHX4 S3_12_6 ( .A(ab_12__6_), .B(CARRYB_11__6_), .CI(ab_11__7_), .CO(
        CARRYB_12__6_), .S(SUMB_12__6_) );
  ADDFHX4 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  ADDFHX4 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  ADDFHX4 S2_7_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  ADDFHX4 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  ADDFHX4 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  ADDFHX4 S2_8_1 ( .A(ab_8__1_), .B(CARRYB_7__1_), .CI(SUMB_7__2_), .CO(
        CARRYB_8__1_), .S(SUMB_8__1_) );
  ADDFHX4 S2_2_4 ( .A(ab_2__4_), .B(n10), .CI(SUMB_1__5_), .CO(CARRYB_2__4_), 
        .S(SUMB_2__4_) );
  ADDFHX4 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  ADDFHX4 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  ADDFHX4 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  ADDFHX4 S2_2_5 ( .A(ab_2__5_), .B(n8), .CI(SUMB_1__6_), .CO(CARRYB_2__5_), 
        .S(SUMB_2__5_) );
  ADDFHX4 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  ADDFHX4 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  ADDFHX4 S2_7_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  ADDFHX4 S3_7_6 ( .A(ab_7__6_), .B(ab_6__7_), .CI(CARRYB_6__6_), .CO(
        CARRYB_7__6_), .S(SUMB_7__6_) );
  ADDFHX4 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  ADDFHX4 S3_2_6 ( .A(ab_2__6_), .B(n11), .CI(ab_1__7_), .CO(CARRYB_2__6_), 
        .S(SUMB_2__6_) );
  ADDFHX4 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  ADDFHX4 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  ADDFHX4 S2_15_4 ( .A(ab_15__4_), .B(CARRYB_14__4_), .CI(SUMB_14__5_), .CO(
        CARRYB_15__4_), .S(SUMB_15__4_) );
  ADDFHX4 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  ADDFHX4 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  ADDFHX4 S2_7_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  ADDFHX4 S2_9_1 ( .A(ab_9__1_), .B(CARRYB_8__1_), .CI(SUMB_8__2_), .CO(
        CARRYB_9__1_), .S(SUMB_9__1_) );
  ADDFHX4 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  ADDFHX4 S2_7_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  ADDFHX4 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  ADDFHX4 S2_2_2 ( .A(ab_2__2_), .B(n14), .CI(SUMB_1__3_), .CO(CARRYB_2__2_), 
        .S(SUMB_2__2_) );
  ADDFHX4 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  ADDFHX4 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  ADDFHX4 S2_2_3 ( .A(ab_2__3_), .B(n13), .CI(SUMB_1__4_), .CO(CARRYB_2__3_), 
        .S(SUMB_2__3_) );
  ADDFHX4 S2_2_1 ( .A(ab_2__1_), .B(n9), .CI(SUMB_1__2_), .CO(CARRYB_2__1_), 
        .S(SUMB_2__1_) );
  ADDFHX4 S3_11_6 ( .A(ab_11__6_), .B(CARRYB_10__6_), .CI(ab_10__7_), .CO(
        CARRYB_11__6_), .S(SUMB_11__6_) );
  ADDFHX2 S1_9_0 ( .A(ab_9__0_), .B(CARRYB_8__0_), .CI(SUMB_8__1_), .CO(
        CARRYB_9__0_), .S(A1_7_) );
  ADDFHX4 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  ADDFHX4 S3_15_6 ( .A(ab_15__6_), .B(CARRYB_14__6_), .CI(ab_14__7_), .CO(
        CARRYB_15__6_), .S(SUMB_15__6_) );
  ADDFHX4 S5_6 ( .A(ab_16__6_), .B(CARRYB_15__6_), .CI(ab_15__7_), .CO(
        CARRYB_16__6_), .S(SUMB_16__6_) );
  ADDFHX4 S2_14_5 ( .A(ab_14__5_), .B(CARRYB_13__5_), .CI(SUMB_13__6_), .CO(
        CARRYB_14__5_), .S(SUMB_14__5_) );
  ADDFHX2 S3_13_6 ( .A(ab_13__6_), .B(CARRYB_12__6_), .CI(ab_12__7_), .CO(
        CARRYB_13__6_), .S(SUMB_13__6_) );
  ADDFHX2 S2_12_1 ( .A(ab_12__1_), .B(CARRYB_11__1_), .CI(SUMB_11__2_), .CO(
        CARRYB_12__1_), .S(SUMB_12__1_) );
  INVX2 U2 ( .A(n37), .Y(n18) );
  NOR2BX4 U3 ( .AN(A[2]), .B(n33), .Y(ab_2__2_) );
  NOR2X4 U4 ( .A(n27), .B(n37), .Y(ab_0__6_) );
  AND2X2 U5 ( .A(A[2]), .B(B[4]), .Y(ab_2__4_) );
  CLKINVX4 U6 ( .A(B[4]), .Y(n41) );
  XOR2X2 U7 ( .A(ab_1__3_), .B(ab_0__4_), .Y(SUMB_1__3_) );
  AND2X2 U8 ( .A(A[3]), .B(n3), .Y(ab_3__4_) );
  CLKINVX20 U9 ( .A(n41), .Y(n3) );
  NOR2BX4 U10 ( .AN(n16), .B(n46), .Y(ab_1__7_) );
  XOR3X4 U11 ( .A(CARRYB_9__1_), .B(ab_10__1_), .C(SUMB_9__2_), .Y(SUMB_10__1_) );
  NAND2X2 U12 ( .A(SUMB_9__2_), .B(CARRYB_9__1_), .Y(n4) );
  NAND2X2 U13 ( .A(ab_10__1_), .B(CARRYB_9__1_), .Y(n5) );
  NAND2X4 U14 ( .A(ab_10__1_), .B(SUMB_9__2_), .Y(n6) );
  NAND3X4 U15 ( .A(n6), .B(n4), .C(n5), .Y(CARRYB_10__1_) );
  NOR2BX4 U16 ( .AN(A[10]), .B(n35), .Y(ab_10__1_) );
  CLKINVX1 U17 ( .A(A[1]), .Y(n15) );
  XOR2X2 U18 ( .A(ab_1__2_), .B(ab_0__3_), .Y(SUMB_1__2_) );
  AND2X4 U19 ( .A(A[1]), .B(B[4]), .Y(ab_1__4_) );
  NOR2BX2 U20 ( .AN(A[5]), .B(n27), .Y(ab_5__6_) );
  AND2X4 U21 ( .A(A[1]), .B(B[3]), .Y(ab_1__3_) );
  CLKINVX4 U22 ( .A(B[3]), .Y(n42) );
  NOR2BX4 U23 ( .AN(A[5]), .B(n46), .Y(ab_5__7_) );
  NOR2BXL U24 ( .AN(A[11]), .B(n31), .Y(ab_11__4_) );
  NOR2BX1 U25 ( .AN(A[11]), .B(n32), .Y(ab_11__3_) );
  NOR2BX2 U26 ( .AN(A[8]), .B(n33), .Y(ab_8__2_) );
  NOR2BX1 U27 ( .AN(A[7]), .B(n35), .Y(ab_7__1_) );
  NOR2BX1 U28 ( .AN(A[9]), .B(n28), .Y(ab_9__6_) );
  NOR2BX1 U29 ( .AN(A[9]), .B(n30), .Y(ab_9__5_) );
  NOR2BX1 U30 ( .AN(A[8]), .B(n41), .Y(ab_8__4_) );
  NOR2BX1 U31 ( .AN(A[14]), .B(n32), .Y(ab_14__3_) );
  NOR2BX1 U32 ( .AN(A[15]), .B(n35), .Y(ab_15__1_) );
  INVX12 U33 ( .A(A[0]), .Y(n37) );
  NOR2BX1 U34 ( .AN(A[9]), .B(n35), .Y(ab_9__1_) );
  NOR2BX1 U35 ( .AN(A[9]), .B(n46), .Y(ab_9__7_) );
  NOR2BX1 U36 ( .AN(A[10]), .B(n28), .Y(ab_10__6_) );
  NOR2BXL U37 ( .AN(A[9]), .B(n31), .Y(ab_9__4_) );
  NOR2BX1 U38 ( .AN(A[11]), .B(n30), .Y(ab_11__5_) );
  NOR2BX2 U39 ( .AN(A[9]), .B(n34), .Y(ab_9__2_) );
  NOR2BX1 U40 ( .AN(A[14]), .B(n35), .Y(ab_14__1_) );
  NOR2BXL U41 ( .AN(A[16]), .B(n32), .Y(ab_16__3_) );
  NOR2BXL U42 ( .AN(A[3]), .B(n36), .Y(ab_3__0_) );
  NOR2BX1 U43 ( .AN(A[11]), .B(n28), .Y(ab_11__6_) );
  NOR2BX1 U44 ( .AN(A[6]), .B(n35), .Y(ab_6__1_) );
  NOR2BX1 U45 ( .AN(A[5]), .B(n31), .Y(ab_5__4_) );
  NOR2BXL U46 ( .AN(A[10]), .B(n31), .Y(ab_10__4_) );
  NOR2BX1 U47 ( .AN(A[10]), .B(n30), .Y(ab_10__5_) );
  NOR2BX1 U48 ( .AN(A[10]), .B(n32), .Y(ab_10__3_) );
  NOR2BXL U49 ( .AN(A[14]), .B(n31), .Y(ab_14__4_) );
  NOR2BXL U50 ( .AN(A[16]), .B(n35), .Y(ab_16__1_) );
  NOR2BX1 U51 ( .AN(A[14]), .B(n30), .Y(ab_14__5_) );
  NOR2BX1 U52 ( .AN(A[7]), .B(n36), .Y(ab_7__0_) );
  AND2X4 U54 ( .A(ab_0__6_), .B(ab_1__5_), .Y(n8) );
  AND2X4 U55 ( .A(ab_0__2_), .B(n47), .Y(n9) );
  AND2X4 U56 ( .A(ab_1__4_), .B(ab_0__5_), .Y(n10) );
  AND2X4 U57 ( .A(ab_1__6_), .B(ab_0__7_), .Y(n11) );
  CLKBUFX2 U58 ( .A(n41), .Y(n31) );
  AND2X4 U59 ( .A(CARRYB_16__1_), .B(SUMB_16__2_), .Y(n12) );
  BUFX3 U60 ( .A(n42), .Y(n32) );
  INVX4 U61 ( .A(B[1]), .Y(n44) );
  CLKBUFX2 U62 ( .A(n44), .Y(n35) );
  NOR2BX1 U63 ( .AN(A[5]), .B(n29), .Y(ab_5__5_) );
  NOR2BX2 U64 ( .AN(A[4]), .B(n27), .Y(ab_4__6_) );
  NAND2X1 U65 ( .A(ab_5__7_), .B(ab_6__6_), .Y(n21) );
  AND2X4 U66 ( .A(ab_1__3_), .B(ab_0__4_), .Y(n13) );
  AND2X4 U67 ( .A(n17), .B(n18), .Y(ab_0__7_) );
  AND2X4 U68 ( .A(ab_1__2_), .B(ab_0__3_), .Y(n14) );
  BUFX4 U69 ( .A(n43), .Y(n34) );
  BUFX16 U70 ( .A(n43), .Y(n33) );
  AND3X4 U71 ( .A(B[1]), .B(n16), .C(n38), .Y(CARRYB_1__0_) );
  XOR2X4 U72 ( .A(ab_1__6_), .B(ab_0__7_), .Y(SUMB_1__6_) );
  DLY1X1 U73 ( .A(n39), .Y(n28) );
  BUFX20 U74 ( .A(n39), .Y(n27) );
  NOR2BX4 U75 ( .AN(A[2]), .B(n27), .Y(ab_2__6_) );
  NOR2BX4 U76 ( .AN(A[3]), .B(n42), .Y(ab_3__3_) );
  NOR2BX4 U77 ( .AN(A[2]), .B(n42), .Y(ab_2__3_) );
  NOR2BX4 U78 ( .AN(A[3]), .B(n44), .Y(ab_3__1_) );
  NOR2BX4 U79 ( .AN(A[3]), .B(n27), .Y(ab_3__6_) );
  NOR2BX4 U80 ( .AN(A[3]), .B(n33), .Y(ab_3__2_) );
  INVX4 U81 ( .A(n15), .Y(n16) );
  XOR2X4 U82 ( .A(ab_0__6_), .B(ab_1__5_), .Y(SUMB_1__5_) );
  NOR2BX1 U83 ( .AN(A[4]), .B(n44), .Y(ab_4__1_) );
  NOR2BX1 U84 ( .AN(A[4]), .B(n41), .Y(ab_4__4_) );
  AND2X2 U85 ( .A(CARRYB_16__2_), .B(SUMB_16__3_), .Y(n22) );
  XOR2X4 U86 ( .A(ab_1__4_), .B(ab_0__5_), .Y(SUMB_1__4_) );
  NOR2BX1 U87 ( .AN(A[7]), .B(n33), .Y(ab_7__2_) );
  NOR2BX1 U88 ( .AN(A[2]), .B(n36), .Y(ab_2__0_) );
  NOR2BX2 U89 ( .AN(A[3]), .B(n29), .Y(ab_3__5_) );
  NOR2BX1 U90 ( .AN(A[6]), .B(n27), .Y(ab_6__6_) );
  XOR3X4 U91 ( .A(CARRYB_5__6_), .B(ab_5__7_), .C(ab_6__6_), .Y(SUMB_6__6_) );
  BUFX8 U92 ( .A(B[7]), .Y(n17) );
  NOR2BX2 U93 ( .AN(A[4]), .B(n42), .Y(ab_4__3_) );
  NOR2BXL U94 ( .AN(A[8]), .B(n27), .Y(ab_8__6_) );
  NOR2BXL U95 ( .AN(A[7]), .B(n27), .Y(ab_7__6_) );
  NOR2BX2 U96 ( .AN(B[3]), .B(n37), .Y(ab_0__3_) );
  NOR2BX4 U97 ( .AN(A[1]), .B(n29), .Y(ab_1__5_) );
  BUFX20 U98 ( .A(n40), .Y(n29) );
  NOR2BX2 U99 ( .AN(A[2]), .B(n29), .Y(ab_2__5_) );
  NOR2BX2 U100 ( .AN(A[2]), .B(n46), .Y(ab_2__7_) );
  NOR2BX2 U101 ( .AN(A[2]), .B(n44), .Y(ab_2__1_) );
  NOR2BX2 U102 ( .AN(A[4]), .B(n33), .Y(ab_4__2_) );
  XOR2X4 U103 ( .A(CARRYB_16__4_), .B(SUMB_16__5_), .Y(A1_19_) );
  AND2X4 U104 ( .A(CARRYB_16__0_), .B(SUMB_16__1_), .Y(n23) );
  NOR2BX4 U105 ( .AN(A[1]), .B(n44), .Y(n47) );
  NAND3X4 U106 ( .A(n21), .B(n19), .C(n20), .Y(CARRYB_6__6_) );
  INVX4 U107 ( .A(B[6]), .Y(n39) );
  NOR2BX4 U108 ( .AN(A[1]), .B(n33), .Y(ab_1__2_) );
  NOR2BX4 U109 ( .AN(B[2]), .B(n37), .Y(ab_0__2_) );
  NOR2BX4 U110 ( .AN(B[4]), .B(n37), .Y(ab_0__4_) );
  NOR2BX4 U111 ( .AN(B[5]), .B(n37), .Y(ab_0__5_) );
  NAND2X1 U112 ( .A(ab_6__6_), .B(CARRYB_5__6_), .Y(n19) );
  NAND2X1 U113 ( .A(ab_5__7_), .B(CARRYB_5__6_), .Y(n20) );
  NOR2BX2 U114 ( .AN(A[6]), .B(n29), .Y(ab_6__5_) );
  NOR2BX2 U115 ( .AN(A[6]), .B(n33), .Y(ab_6__2_) );
  NOR2BX2 U116 ( .AN(A[6]), .B(n41), .Y(ab_6__4_) );
  NOR2BX2 U117 ( .AN(A[6]), .B(n46), .Y(ab_6__7_) );
  NOR2BX2 U118 ( .AN(A[6]), .B(n32), .Y(ab_6__3_) );
  NOR2BX1 U119 ( .AN(A[14]), .B(n36), .Y(ab_14__0_) );
  NOR2BX1 U120 ( .AN(A[13]), .B(n35), .Y(ab_13__1_) );
  NOR2BX1 U121 ( .AN(A[15]), .B(n34), .Y(ab_15__2_) );
  NOR2BX1 U122 ( .AN(A[16]), .B(n36), .Y(ab_16__0_) );
  NOR2BX1 U123 ( .AN(A[13]), .B(n36), .Y(ab_13__0_) );
  NOR2BX1 U124 ( .AN(A[15]), .B(n36), .Y(ab_15__0_) );
  NOR2BX1 U125 ( .AN(A[5]), .B(n33), .Y(ab_5__2_) );
  NOR2BX1 U126 ( .AN(A[8]), .B(n29), .Y(ab_8__5_) );
  NOR2BX1 U127 ( .AN(A[7]), .B(n32), .Y(ab_7__3_) );
  NOR2BX1 U128 ( .AN(A[4]), .B(n46), .Y(ab_4__7_) );
  NOR2BX1 U129 ( .AN(A[4]), .B(n29), .Y(ab_4__5_) );
  NOR2BX1 U130 ( .AN(A[11]), .B(n36), .Y(ab_11__0_) );
  NOR2BX1 U131 ( .AN(A[9]), .B(n36), .Y(ab_9__0_) );
  NOR2BX1 U132 ( .AN(A[11]), .B(n35), .Y(ab_11__1_) );
  NOR2BX1 U133 ( .AN(A[11]), .B(n34), .Y(ab_11__2_) );
  NOR2BX1 U134 ( .AN(A[3]), .B(n46), .Y(ab_3__7_) );
  INVX4 U135 ( .A(B[2]), .Y(n43) );
  NOR2BXL U136 ( .AN(A[10]), .B(n46), .Y(ab_10__7_) );
  NOR2BXL U137 ( .AN(A[8]), .B(n32), .Y(ab_8__3_) );
  NOR2BX1 U138 ( .AN(A[8]), .B(n46), .Y(ab_8__7_) );
  NOR2BXL U139 ( .AN(A[7]), .B(n29), .Y(ab_7__5_) );
  NOR2BX1 U140 ( .AN(A[10]), .B(n34), .Y(ab_10__2_) );
  NOR2BXL U141 ( .AN(A[12]), .B(n36), .Y(ab_12__0_) );
  NOR2BX1 U142 ( .AN(A[13]), .B(n34), .Y(ab_13__2_) );
  NOR2BX1 U143 ( .AN(A[13]), .B(n31), .Y(ab_13__4_) );
  NOR2BX1 U144 ( .AN(A[13]), .B(n32), .Y(ab_13__3_) );
  XOR2X2 U145 ( .A(CARRYB_16__5_), .B(SUMB_16__6_), .Y(A1_20_) );
  NOR2BX1 U146 ( .AN(A[8]), .B(n35), .Y(ab_8__1_) );
  NOR2BXL U147 ( .AN(A[7]), .B(n41), .Y(ab_7__4_) );
  NOR2BX1 U148 ( .AN(A[10]), .B(n36), .Y(ab_10__0_) );
  NOR2BX1 U149 ( .AN(A[13]), .B(n30), .Y(ab_13__5_) );
  AND2X1 U150 ( .A(CARRYB_16__5_), .B(SUMB_16__6_), .Y(n26) );
  NOR2BX4 U151 ( .AN(A[1]), .B(n27), .Y(ab_1__6_) );
  NOR2BX1 U152 ( .AN(A[16]), .B(n30), .Y(ab_16__5_) );
  NOR2BX1 U153 ( .AN(A[15]), .B(n31), .Y(ab_15__4_) );
  NOR2BX1 U154 ( .AN(A[15]), .B(n32), .Y(ab_15__3_) );
  INVX8 U155 ( .A(n17), .Y(n46) );
  BUFX1 U156 ( .A(n40), .Y(n30) );
  NOR2BXL U157 ( .AN(A[13]), .B(n46), .Y(ab_13__7_) );
  NOR2BX1 U158 ( .AN(A[14]), .B(n28), .Y(ab_14__6_) );
  NOR2BX1 U159 ( .AN(A[5]), .B(n36), .Y(ab_5__0_) );
  NOR2BX1 U160 ( .AN(A[4]), .B(n36), .Y(ab_4__0_) );
  NOR2BX2 U161 ( .AN(A[14]), .B(n34), .Y(ab_14__2_) );
  NOR2BXL U162 ( .AN(A[12]), .B(n35), .Y(ab_12__1_) );
  NOR2BXL U163 ( .AN(A[12]), .B(n34), .Y(ab_12__2_) );
  NOR2BXL U164 ( .AN(A[12]), .B(n32), .Y(ab_12__3_) );
  NOR2BXL U165 ( .AN(A[12]), .B(n31), .Y(ab_12__4_) );
  NOR2BX1 U166 ( .AN(A[6]), .B(n36), .Y(ab_6__0_) );
  NOR2BX1 U167 ( .AN(A[8]), .B(n36), .Y(ab_8__0_) );
  NOR2BXL U168 ( .AN(A[12]), .B(n30), .Y(ab_12__5_) );
  NOR2BX2 U169 ( .AN(A[9]), .B(n32), .Y(ab_9__3_) );
  NOR2BX1 U170 ( .AN(A[11]), .B(n46), .Y(ab_11__7_) );
  NOR2BXL U171 ( .AN(A[12]), .B(n28), .Y(ab_12__6_) );
  NOR2BX1 U172 ( .AN(A[7]), .B(n46), .Y(ab_7__7_) );
  NOR2BX1 U173 ( .AN(A[5]), .B(n42), .Y(ab_5__3_) );
  AND2X2 U174 ( .A(CARRYB_16__3_), .B(SUMB_16__4_), .Y(n24) );
  AND2X2 U175 ( .A(CARRYB_16__4_), .B(SUMB_16__5_), .Y(n25) );
  NOR2BX2 U176 ( .AN(A[5]), .B(n44), .Y(ab_5__1_) );
  NOR2BXL U177 ( .AN(A[12]), .B(n46), .Y(ab_12__7_) );
  NOR2BXL U178 ( .AN(A[13]), .B(n28), .Y(ab_13__6_) );
  XOR2X1 U179 ( .A(n47), .B(ab_0__2_), .Y(SUMB_1__1_) );
  BUFX3 U180 ( .A(n45), .Y(n36) );
  INVX1 U181 ( .A(B[0]), .Y(n45) );
  XOR2X1 U182 ( .A(CARRYB_16__6_), .B(ab_16__7_), .Y(A1_21_) );
  NOR2BX1 U183 ( .AN(A[16]), .B(n28), .Y(ab_16__6_) );
  NOR2BXL U184 ( .AN(A[15]), .B(n46), .Y(ab_15__7_) );
  NOR2BXL U185 ( .AN(A[15]), .B(n30), .Y(ab_15__5_) );
  NOR2BX1 U186 ( .AN(A[16]), .B(n34), .Y(ab_16__2_) );
  NOR2BX1 U187 ( .AN(A[16]), .B(n31), .Y(ab_16__4_) );
  NOR2BX1 U188 ( .AN(A[14]), .B(n46), .Y(ab_14__7_) );
  NOR2BXL U189 ( .AN(A[15]), .B(n28), .Y(ab_15__6_) );
  NOR2BXL U190 ( .AN(A[16]), .B(n46), .Y(ab_16__7_) );
  NOR2BX1 U191 ( .AN(A[0]), .B(n36), .Y(n38) );
  XOR2X4 U192 ( .A(SUMB_16__3_), .B(CARRYB_16__2_), .Y(A1_17_) );
  XOR2X4 U193 ( .A(SUMB_16__1_), .B(CARRYB_16__0_), .Y(A1_15_) );
  XOR2X4 U194 ( .A(CARRYB_16__3_), .B(SUMB_16__4_), .Y(A1_18_) );
  XOR2X4 U195 ( .A(SUMB_16__2_), .B(CARRYB_16__1_), .Y(A1_16_) );
  INVX8 U196 ( .A(B[5]), .Y(n40) );
endmodule


module multi16_4 ( in_17bit, in_8bit, out );
  input [16:0] in_17bit;
  input [7:0] in_8bit;
  output [16:0] out;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123;
  wire   [16:1] in_17bit_b;
  wire   [7:1] in_8bit_b;
  wire   [23:8] mul;

  multi16_4_DW02_mult_0 mult_55 ( .A({in_17bit_b[16:4], n27, in_17bit_b[2:1], 
        in_17bit[0]}), .B({in_8bit_b, in_8bit[0]}), .PRODUCT_23_(mul[23]), 
        .PRODUCT_22_(mul[22]), .PRODUCT_21_(mul[21]), .PRODUCT_20_(mul[20]), 
        .PRODUCT_19_(mul[19]), .PRODUCT_18_(mul[18]), .PRODUCT_17_(mul[17]), 
        .PRODUCT_16_(mul[16]), .PRODUCT_15_(mul[15]), .PRODUCT_14_(mul[14]), 
        .PRODUCT_13_(mul[13]), .PRODUCT_12_(mul[12]), .PRODUCT_11_(mul[11]), 
        .PRODUCT_10_(mul[10]), .PRODUCT_9_(mul[9]), .PRODUCT_8_(mul[8]), 
        .PRODUCT_7_(out[0]) );
  NOR2X4 U2 ( .A(n62), .B(n64), .Y(n38) );
  BUFX16 U3 ( .A(in_17bit[16]), .Y(n53) );
  NAND2BX4 U4 ( .AN(n64), .B(n59), .Y(n58) );
  BUFX12 U5 ( .A(n55), .Y(n8) );
  BUFX12 U6 ( .A(in_8bit[5]), .Y(n55) );
  CLKINVX8 U7 ( .A(in_8bit[4]), .Y(n54) );
  AND2X4 U8 ( .A(n53), .B(n66), .Y(n14) );
  INVX16 U9 ( .A(n53), .Y(n96) );
  INVX8 U10 ( .A(n18), .Y(n19) );
  NAND2X1 U11 ( .A(mul[15]), .B(n36), .Y(n22) );
  NAND2X4 U12 ( .A(n63), .B(n62), .Y(n9) );
  NAND3X4 U13 ( .A(n1), .B(n2), .C(n3), .Y(n50) );
  NAND3X2 U14 ( .A(in_17bit[1]), .B(n53), .C(in_17bit[0]), .Y(n1) );
  OR2X4 U15 ( .A(in_17bit[1]), .B(n53), .Y(n2) );
  OR2X4 U16 ( .A(in_17bit[1]), .B(in_17bit[0]), .Y(n3) );
  CLKINVX8 U17 ( .A(in_17bit[6]), .Y(n73) );
  CLKINVX1 U18 ( .A(n119), .Y(n122) );
  XOR2X2 U19 ( .A(n70), .B(n68), .Y(in_17bit_b[5]) );
  NAND2X2 U20 ( .A(n53), .B(n69), .Y(n68) );
  INVX8 U21 ( .A(n44), .Y(n62) );
  CLKINVX8 U22 ( .A(in_8bit[2]), .Y(n57) );
  INVX4 U23 ( .A(in_17bit[2]), .Y(n18) );
  INVX1 U24 ( .A(n109), .Y(n13) );
  INVX1 U25 ( .A(in_8bit[3]), .Y(n17) );
  NAND2X2 U26 ( .A(n106), .B(n114), .Y(n36) );
  INVXL U27 ( .A(n114), .Y(n7) );
  CLKINVX2 U28 ( .A(in_8bit[6]), .Y(n11) );
  NAND2X4 U29 ( .A(n103), .B(n114), .Y(n33) );
  CLKBUFXL U30 ( .A(n53), .Y(n4) );
  BUFX16 U31 ( .A(in_17bit_b[3]), .Y(n27) );
  XOR2X4 U32 ( .A(in_17bit[3]), .B(n14), .Y(in_17bit_b[3]) );
  XOR2X4 U33 ( .A(mul[23]), .B(n123), .Y(out[16]) );
  OR2X2 U34 ( .A(mul[14]), .B(n105), .Y(n106) );
  NAND2X4 U35 ( .A(n9), .B(in_8bit[7]), .Y(n37) );
  NAND2BX4 U36 ( .AN(mul[18]), .B(n5), .Y(n118) );
  NOR2X1 U37 ( .A(mul[17]), .B(n110), .Y(n5) );
  XOR2X4 U38 ( .A(n6), .B(n121), .Y(out[15]) );
  NAND2X4 U39 ( .A(n114), .B(n119), .Y(n6) );
  INVX3 U40 ( .A(mul[21]), .Y(n116) );
  XNOR2X4 U41 ( .A(mul[17]), .B(n31), .Y(out[10]) );
  OAI21X2 U42 ( .A0(n56), .A1(n59), .B0(in_8bit[7]), .Y(n60) );
  XOR2X2 U43 ( .A(n57), .B(n58), .Y(in_8bit_b[2]) );
  INVX2 U44 ( .A(n57), .Y(n56) );
  XNOR2X4 U45 ( .A(in_8bit[1]), .B(n41), .Y(in_8bit_b[1]) );
  INVX3 U46 ( .A(in_8bit[0]), .Y(n16) );
  OAI21X4 U47 ( .A0(in_17bit[0]), .A1(in_17bit[1]), .B0(n53), .Y(n65) );
  XNOR2X4 U48 ( .A(mul[13]), .B(n33), .Y(out[6]) );
  NOR2BX4 U49 ( .AN(n118), .B(n7), .Y(n113) );
  AND2X1 U50 ( .A(n53), .B(n80), .Y(n40) );
  NAND2XL U51 ( .A(n53), .B(n75), .Y(n74) );
  NAND2XL U52 ( .A(n4), .B(n91), .Y(n90) );
  XNOR2X1 U53 ( .A(n53), .B(in_8bit[7]), .Y(n120) );
  XOR2X2 U54 ( .A(mul[11]), .B(n35), .Y(out[4]) );
  XOR2X2 U55 ( .A(n76), .B(n74), .Y(in_17bit_b[7]) );
  NAND2X4 U56 ( .A(n45), .B(n73), .Y(n75) );
  NOR2X4 U57 ( .A(n55), .B(in_8bit[4]), .Y(n63) );
  AOI2BB1X4 U58 ( .A0N(n10), .A1N(mul[20]), .B0(n120), .Y(n117) );
  OR2X4 U59 ( .A(mul[19]), .B(n118), .Y(n10) );
  OR2X4 U60 ( .A(n111), .B(mul[18]), .Y(n26) );
  XOR2X4 U61 ( .A(n37), .B(n11), .Y(in_8bit_b[6]) );
  AND2X4 U62 ( .A(n98), .B(n114), .Y(n43) );
  CLKINVX1 U63 ( .A(mul[15]), .Y(n20) );
  BUFX8 U64 ( .A(mul[19]), .Y(n12) );
  NAND2BX4 U65 ( .AN(mul[16]), .B(n13), .Y(n110) );
  OAI21X2 U66 ( .A0(n118), .A1(mul[19]), .B0(n114), .Y(n115) );
  XOR2X4 U67 ( .A(mul[9]), .B(n43), .Y(out[2]) );
  INVX8 U68 ( .A(n50), .Y(in_17bit_b[1]) );
  NAND4X4 U69 ( .A(n57), .B(n15), .C(n16), .D(n17), .Y(n44) );
  CLKINVX20 U70 ( .A(in_8bit[1]), .Y(n15) );
  CLKINVX2 U71 ( .A(in_17bit[5]), .Y(n70) );
  NAND2X2 U72 ( .A(in_8bit[0]), .B(in_8bit[7]), .Y(n41) );
  XOR2X4 U73 ( .A(n39), .B(n67), .Y(in_17bit_b[4]) );
  NOR3X2 U74 ( .A(n9), .B(in_8bit[6]), .C(n64), .Y(in_8bit_b[7]) );
  XNOR2X4 U75 ( .A(n78), .B(n79), .Y(in_17bit_b[8]) );
  XOR2X4 U76 ( .A(mul[8]), .B(n32), .Y(out[1]) );
  OR2X4 U77 ( .A(in_8bit[1]), .B(in_8bit[0]), .Y(n59) );
  NAND2X4 U78 ( .A(n51), .B(n67), .Y(n69) );
  NOR2X4 U79 ( .A(in_17bit[3]), .B(n66), .Y(n51) );
  XNOR2X4 U80 ( .A(n65), .B(n19), .Y(in_17bit_b[2]) );
  OR3X4 U81 ( .A(in_17bit[2]), .B(in_17bit[1]), .C(in_17bit[0]), .Y(n66) );
  XNOR2X4 U82 ( .A(n60), .B(in_8bit[3]), .Y(in_8bit_b[3]) );
  XOR2X4 U83 ( .A(n113), .B(n12), .Y(out[12]) );
  NAND2X2 U84 ( .A(n111), .B(mul[18]), .Y(n25) );
  NAND2X4 U85 ( .A(n112), .B(n114), .Y(n111) );
  INVX8 U86 ( .A(in_8bit[7]), .Y(n64) );
  OR3X4 U87 ( .A(mul[21]), .B(n10), .C(mul[20]), .Y(n119) );
  XNOR2X4 U88 ( .A(n38), .B(n54), .Y(in_8bit_b[4]) );
  XNOR2X4 U89 ( .A(mul[12]), .B(n34), .Y(out[5]) );
  NAND2X4 U90 ( .A(n102), .B(n114), .Y(n34) );
  NOR2X4 U91 ( .A(n45), .B(n96), .Y(n72) );
  NAND2X2 U92 ( .A(n20), .B(n21), .Y(n23) );
  NAND2X4 U93 ( .A(n22), .B(n23), .Y(out[8]) );
  INVX1 U94 ( .A(n36), .Y(n21) );
  NAND2X2 U95 ( .A(n122), .B(n121), .Y(n24) );
  AND2X4 U96 ( .A(n24), .B(n114), .Y(n123) );
  INVX8 U97 ( .A(mul[22]), .Y(n121) );
  NAND2X4 U98 ( .A(n26), .B(n25), .Y(out[11]) );
  CLKINVX4 U99 ( .A(in_17bit[4]), .Y(n67) );
  NAND2X2 U100 ( .A(n72), .B(n73), .Y(n29) );
  NAND2X4 U101 ( .A(n28), .B(in_17bit[6]), .Y(n30) );
  NAND2X4 U102 ( .A(n29), .B(n30), .Y(in_17bit_b[6]) );
  INVX2 U103 ( .A(n72), .Y(n28) );
  NAND2X4 U104 ( .A(n110), .B(n114), .Y(n31) );
  OR2X4 U105 ( .A(mul[17]), .B(n110), .Y(n112) );
  NAND2X1 U106 ( .A(n47), .B(n89), .Y(n91) );
  AND2X4 U107 ( .A(out[0]), .B(n114), .Y(n32) );
  OR2X4 U108 ( .A(mul[10]), .B(n100), .Y(n101) );
  AND2X2 U109 ( .A(n101), .B(n114), .Y(n35) );
  XNOR2X2 U110 ( .A(n42), .B(n89), .Y(in_17bit_b[12]) );
  OR2X4 U111 ( .A(mul[13]), .B(n103), .Y(n105) );
  OR2X4 U112 ( .A(mul[9]), .B(n98), .Y(n100) );
  OR2X4 U113 ( .A(mul[12]), .B(n102), .Y(n103) );
  OR2X4 U114 ( .A(mul[8]), .B(out[0]), .Y(n98) );
  INVX4 U115 ( .A(n120), .Y(n114) );
  OR2X4 U116 ( .A(n51), .B(n96), .Y(n39) );
  AND2X4 U117 ( .A(n71), .B(n70), .Y(n45) );
  XNOR2X4 U118 ( .A(n81), .B(n40), .Y(in_17bit_b[9]) );
  AND2X4 U119 ( .A(n77), .B(n76), .Y(n49) );
  NAND2X4 U120 ( .A(n46), .B(n95), .Y(n97) );
  NOR2XL U121 ( .A(n47), .B(n96), .Y(n42) );
  AND2X4 U122 ( .A(n88), .B(n87), .Y(n47) );
  AND2X4 U123 ( .A(n82), .B(n81), .Y(n48) );
  AND2X4 U124 ( .A(n93), .B(n92), .Y(n46) );
  NAND2XL U125 ( .A(n4), .B(n86), .Y(n85) );
  INVXL U126 ( .A(in_17bit[8]), .Y(n79) );
  INVXL U127 ( .A(in_17bit[10]), .Y(n84) );
  INVXL U128 ( .A(in_17bit[11]), .Y(n87) );
  INVXL U129 ( .A(in_17bit[13]), .Y(n92) );
  OR2X2 U130 ( .A(mul[11]), .B(n101), .Y(n102) );
  NOR2X1 U131 ( .A(n49), .B(n96), .Y(n78) );
  XOR2X1 U132 ( .A(n92), .B(n90), .Y(in_17bit_b[13]) );
  NAND2X1 U133 ( .A(n48), .B(n84), .Y(n86) );
  NAND2X1 U134 ( .A(n49), .B(n79), .Y(n80) );
  XOR2X2 U135 ( .A(in_17bit[15]), .B(n52), .Y(in_17bit_b[15]) );
  AND2X1 U136 ( .A(n4), .B(n97), .Y(n52) );
  INVXL U137 ( .A(in_17bit[9]), .Y(n81) );
  INVXL U138 ( .A(in_17bit[7]), .Y(n76) );
  AOI21X4 U139 ( .A0(n62), .A1(n54), .B0(n64), .Y(n61) );
  XOR2X4 U140 ( .A(n61), .B(n8), .Y(in_8bit_b[5]) );
  CLKINVX3 U141 ( .A(n69), .Y(n71) );
  CLKINVX3 U142 ( .A(n75), .Y(n77) );
  CLKINVX3 U143 ( .A(n80), .Y(n82) );
  NOR2X4 U144 ( .A(n48), .B(n96), .Y(n83) );
  XNOR2X4 U145 ( .A(n83), .B(n84), .Y(in_17bit_b[10]) );
  XOR2X4 U146 ( .A(n87), .B(n85), .Y(in_17bit_b[11]) );
  CLKINVX3 U147 ( .A(n86), .Y(n88) );
  CLKINVX3 U148 ( .A(in_17bit[12]), .Y(n89) );
  CLKINVX3 U149 ( .A(n91), .Y(n93) );
  NOR2X4 U150 ( .A(n46), .B(n96), .Y(n94) );
  CLKINVX3 U151 ( .A(in_17bit[14]), .Y(n95) );
  XNOR2X4 U152 ( .A(n94), .B(n95), .Y(in_17bit_b[14]) );
  NOR3X4 U153 ( .A(in_17bit[15]), .B(n97), .C(n96), .Y(in_17bit_b[16]) );
  NAND2X4 U154 ( .A(n100), .B(n114), .Y(n99) );
  XNOR2X4 U155 ( .A(mul[10]), .B(n99), .Y(out[3]) );
  NAND2X4 U156 ( .A(n105), .B(n114), .Y(n104) );
  XNOR2X4 U157 ( .A(mul[14]), .B(n104), .Y(out[7]) );
  CLKINVX3 U158 ( .A(n106), .Y(n107) );
  NAND2BX4 U159 ( .AN(mul[15]), .B(n107), .Y(n109) );
  NAND2X4 U160 ( .A(n109), .B(n114), .Y(n108) );
  XNOR2X4 U161 ( .A(mul[16]), .B(n108), .Y(out[9]) );
  XNOR2X4 U162 ( .A(n115), .B(mul[20]), .Y(out[13]) );
  XNOR2X4 U163 ( .A(n117), .B(n116), .Y(out[14]) );
endmodule


module multi16_3_DW01_add_0 ( A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, 
        A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, 
        B_20_, B_19_, B_18_, B_17_, B_16_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, 
        SUM_17_, SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, 
        SUM_9_, SUM_8_, SUM_7_, SUM_6_, SUM_5_ );
  input A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_,
         A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, B_20_, B_19_,
         B_18_, B_17_, B_16_;
  output SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, SUM_15_,
         SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, SUM_7_,
         SUM_6_, SUM_5_;
  wire   n1, n2, n3, n4, n5, n7, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42;

  XOR2X2 U2 ( .A(n25), .B(n26), .Y(SUM_21_) );
  BUFX8 U3 ( .A(n23), .Y(n1) );
  INVX2 U4 ( .A(n21), .Y(n2) );
  AOI21X1 U5 ( .A0(n27), .A1(n28), .B0(n18), .Y(n26) );
  BUFX12 U6 ( .A(A_9_), .Y(SUM_9_) );
  BUFX12 U7 ( .A(A_12_), .Y(SUM_12_) );
  OAI21X1 U8 ( .A0(n37), .A1(n33), .B0(n2), .Y(n35) );
  OAI21X4 U9 ( .A0(n41), .A1(n3), .B0(n36), .Y(n39) );
  NOR2X4 U10 ( .A(n23), .B(n7), .Y(SUM_16_) );
  INVX8 U11 ( .A(n37), .Y(n23) );
  BUFX12 U12 ( .A(A_8_), .Y(SUM_8_) );
  XOR2X4 U13 ( .A(n5), .B(n27), .Y(SUM_20_) );
  BUFX12 U14 ( .A(A_11_), .Y(SUM_11_) );
  BUFX12 U15 ( .A(A_14_), .Y(SUM_14_) );
  INVX8 U16 ( .A(n24), .Y(SUM_15_) );
  INVX8 U17 ( .A(A_15_), .Y(n24) );
  INVX8 U18 ( .A(n38), .Y(n21) );
  NAND2X4 U19 ( .A(B_19_), .B(A_19_), .Y(n32) );
  AOI21X2 U20 ( .A0(n19), .A1(n35), .B0(n20), .Y(n30) );
  INVX3 U21 ( .A(n19), .Y(n3) );
  INVX8 U22 ( .A(n34), .Y(n19) );
  OAI21X4 U23 ( .A0(n30), .A1(n31), .B0(n32), .Y(n27) );
  NOR2X4 U24 ( .A(B_19_), .B(A_19_), .Y(n31) );
  NOR2X2 U25 ( .A(A_16_), .B(B_16_), .Y(n7) );
  NAND2X2 U26 ( .A(n36), .B(n19), .Y(n42) );
  BUFX12 U27 ( .A(A_6_), .Y(SUM_6_) );
  OR2X4 U28 ( .A(B_20_), .B(A_20_), .Y(n28) );
  INVX4 U29 ( .A(n33), .Y(n22) );
  NOR2X4 U30 ( .A(A_17_), .B(B_17_), .Y(n33) );
  NOR2BX4 U31 ( .AN(n32), .B(n31), .Y(n40) );
  NAND2X4 U32 ( .A(A_16_), .B(B_16_), .Y(n37) );
  AOI21X4 U33 ( .A0(n22), .A1(n23), .B0(n21), .Y(n41) );
  INVXL U34 ( .A(n36), .Y(n20) );
  NAND2X4 U35 ( .A(A_17_), .B(B_17_), .Y(n38) );
  NOR2X4 U36 ( .A(n21), .B(n33), .Y(n4) );
  XOR2X4 U37 ( .A(n1), .B(n4), .Y(SUM_17_) );
  INVXL U38 ( .A(n29), .Y(n18) );
  NAND2X4 U39 ( .A(B_18_), .B(A_18_), .Y(n36) );
  AND2X2 U40 ( .A(n29), .B(n28), .Y(n5) );
  BUFX8 U41 ( .A(A_5_), .Y(SUM_5_) );
  BUFX8 U42 ( .A(A_7_), .Y(SUM_7_) );
  BUFX8 U43 ( .A(A_13_), .Y(SUM_13_) );
  BUFX8 U44 ( .A(A_10_), .Y(SUM_10_) );
  XOR2X4 U45 ( .A(n39), .B(n40), .Y(SUM_19_) );
  NOR2X4 U46 ( .A(B_18_), .B(A_18_), .Y(n34) );
  XOR2X4 U47 ( .A(n41), .B(n42), .Y(SUM_18_) );
  XNOR2X1 U48 ( .A(B_21_), .B(A_21_), .Y(n25) );
  NAND2X1 U49 ( .A(B_20_), .B(A_20_), .Y(n29) );
endmodule


module multi16_3_DW02_mult_0 ( A, B, PRODUCT_23_, PRODUCT_22_, PRODUCT_21_, 
        PRODUCT_20_, PRODUCT_19_, PRODUCT_18_, PRODUCT_17_, PRODUCT_16_, 
        PRODUCT_15_, PRODUCT_14_, PRODUCT_13_, PRODUCT_12_, PRODUCT_11_, 
        PRODUCT_10_, PRODUCT_9_, PRODUCT_8_, PRODUCT_7_ );
  input [16:0] A;
  input [7:0] B;
  output PRODUCT_23_, PRODUCT_22_, PRODUCT_21_, PRODUCT_20_, PRODUCT_19_,
         PRODUCT_18_, PRODUCT_17_, PRODUCT_16_, PRODUCT_15_, PRODUCT_14_,
         PRODUCT_13_, PRODUCT_12_, PRODUCT_11_, PRODUCT_10_, PRODUCT_9_,
         PRODUCT_8_, PRODUCT_7_;
  wire   ab_16__7_, ab_16__6_, ab_16__5_, ab_16__4_, ab_16__3_, ab_16__2_,
         ab_16__1_, ab_16__0_, ab_15__7_, ab_15__6_, ab_15__5_, ab_15__4_,
         ab_15__3_, ab_15__2_, ab_15__1_, ab_15__0_, ab_14__7_, ab_14__6_,
         ab_14__5_, ab_14__4_, ab_14__3_, ab_14__2_, ab_14__1_, ab_14__0_,
         ab_13__7_, ab_13__6_, ab_13__5_, ab_13__4_, ab_13__3_, ab_13__2_,
         ab_13__1_, ab_13__0_, ab_12__7_, ab_12__6_, ab_12__5_, ab_12__4_,
         ab_12__3_, ab_12__2_, ab_12__1_, ab_12__0_, ab_11__7_, ab_11__6_,
         ab_11__5_, ab_11__4_, ab_11__3_, ab_11__2_, ab_11__1_, ab_11__0_,
         ab_10__7_, ab_10__6_, ab_10__5_, ab_10__4_, ab_10__3_, ab_10__2_,
         ab_10__1_, ab_10__0_, ab_9__7_, ab_9__6_, ab_9__5_, ab_9__4_,
         ab_9__3_, ab_9__2_, ab_9__1_, ab_9__0_, ab_8__7_, ab_8__6_, ab_8__5_,
         ab_8__4_, ab_8__3_, ab_8__2_, ab_8__1_, ab_8__0_, ab_7__7_, ab_7__6_,
         ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_, ab_7__0_, ab_6__7_,
         ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_, ab_6__1_, ab_6__0_,
         ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_, ab_5__2_, ab_5__1_,
         ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_, ab_4__3_, ab_4__2_,
         ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_, ab_3__4_, ab_3__3_,
         ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_, ab_2__5_, ab_2__4_,
         ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_, ab_1__6_, ab_1__5_,
         ab_1__4_, ab_1__3_, ab_1__2_, ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_,
         ab_0__3_, ab_0__2_, CARRYB_16__6_, CARRYB_16__5_, CARRYB_16__4_,
         CARRYB_16__3_, CARRYB_16__2_, CARRYB_16__1_, CARRYB_16__0_,
         CARRYB_15__6_, CARRYB_15__5_, CARRYB_15__4_, CARRYB_15__3_,
         CARRYB_15__2_, CARRYB_15__1_, CARRYB_15__0_, CARRYB_14__6_,
         CARRYB_14__5_, CARRYB_14__4_, CARRYB_14__3_, CARRYB_14__2_,
         CARRYB_14__1_, CARRYB_14__0_, CARRYB_13__6_, CARRYB_13__5_,
         CARRYB_13__4_, CARRYB_13__3_, CARRYB_13__2_, CARRYB_13__1_,
         CARRYB_13__0_, CARRYB_12__6_, CARRYB_12__5_, CARRYB_12__4_,
         CARRYB_12__3_, CARRYB_12__2_, CARRYB_12__1_, CARRYB_12__0_,
         CARRYB_11__6_, CARRYB_11__5_, CARRYB_11__4_, CARRYB_11__3_,
         CARRYB_11__2_, CARRYB_11__1_, CARRYB_11__0_, CARRYB_10__6_,
         CARRYB_10__5_, CARRYB_10__4_, CARRYB_10__3_, CARRYB_10__2_,
         CARRYB_10__1_, CARRYB_10__0_, CARRYB_9__6_, CARRYB_9__5_,
         CARRYB_9__4_, CARRYB_9__3_, CARRYB_9__2_, CARRYB_9__1_, CARRYB_9__0_,
         CARRYB_8__6_, CARRYB_8__5_, CARRYB_8__4_, CARRYB_8__3_, CARRYB_8__2_,
         CARRYB_8__1_, CARRYB_8__0_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_,
         CARRYB_7__3_, CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_,
         CARRYB_6__5_, CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_,
         CARRYB_6__0_, CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_,
         CARRYB_5__2_, CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_,
         CARRYB_4__4_, CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_,
         CARRYB_3__6_, CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_,
         CARRYB_3__1_, CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_,
         CARRYB_2__3_, CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__2_,
         CARRYB_1__0_, SUMB_16__6_, SUMB_16__5_, SUMB_16__4_, SUMB_16__3_,
         SUMB_16__2_, SUMB_16__1_, SUMB_16__0_, SUMB_15__6_, SUMB_15__5_,
         SUMB_15__4_, SUMB_15__3_, SUMB_15__2_, SUMB_15__1_, SUMB_14__6_,
         SUMB_14__5_, SUMB_14__4_, SUMB_14__3_, SUMB_14__2_, SUMB_14__1_,
         SUMB_13__6_, SUMB_13__5_, SUMB_13__4_, SUMB_13__3_, SUMB_13__2_,
         SUMB_13__1_, SUMB_12__6_, SUMB_12__5_, SUMB_12__4_, SUMB_12__3_,
         SUMB_12__2_, SUMB_12__1_, SUMB_11__6_, SUMB_11__5_, SUMB_11__4_,
         SUMB_11__3_, SUMB_11__2_, SUMB_11__1_, SUMB_10__6_, SUMB_10__5_,
         SUMB_10__4_, SUMB_10__3_, SUMB_10__2_, SUMB_10__1_, SUMB_9__6_,
         SUMB_9__5_, SUMB_9__4_, SUMB_9__3_, SUMB_9__2_, SUMB_9__1_,
         SUMB_8__6_, SUMB_8__5_, SUMB_8__4_, SUMB_8__3_, SUMB_8__2_,
         SUMB_8__1_, SUMB_7__6_, SUMB_7__5_, SUMB_7__4_, SUMB_7__3_,
         SUMB_7__2_, SUMB_7__1_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_,
         SUMB_6__3_, SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_,
         SUMB_5__4_, SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_,
         SUMB_4__5_, SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_,
         SUMB_3__6_, SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_,
         SUMB_3__1_, SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_,
         SUMB_2__2_, SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_,
         SUMB_1__3_, SUMB_1__2_, SUMB_1__1_, PROD1_7_, A1_21_, A1_20_, A1_19_,
         A1_18_, A1_17_, A1_16_, A1_15_, A1_13_, A1_12_, A1_11_, A1_10_, A1_9_,
         A1_8_, A1_7_, A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, n3, n5, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38;

  multi16_3_DW01_add_0 FS_1 ( .A_21_(A1_21_), .A_20_(A1_20_), .A_19_(A1_19_), 
        .A_18_(A1_18_), .A_17_(A1_17_), .A_16_(A1_16_), .A_15_(A1_15_), 
        .A_14_(SUMB_16__0_), .A_13_(A1_13_), .A_12_(A1_12_), .A_11_(A1_11_), 
        .A_10_(A1_10_), .A_9_(A1_9_), .A_8_(A1_8_), .A_7_(A1_7_), .A_6_(A1_6_), 
        .A_5_(PROD1_7_), .B_21_(n16), .B_20_(n15), .B_19_(n14), .B_18_(n11), 
        .B_17_(n12), .B_16_(n13), .SUM_21_(PRODUCT_23_), .SUM_20_(PRODUCT_22_), 
        .SUM_19_(PRODUCT_21_), .SUM_18_(PRODUCT_20_), .SUM_17_(PRODUCT_19_), 
        .SUM_16_(PRODUCT_18_), .SUM_15_(PRODUCT_17_), .SUM_14_(PRODUCT_16_), 
        .SUM_13_(PRODUCT_15_), .SUM_12_(PRODUCT_14_), .SUM_11_(PRODUCT_13_), 
        .SUM_10_(PRODUCT_12_), .SUM_9_(PRODUCT_11_), .SUM_8_(PRODUCT_10_), 
        .SUM_7_(PRODUCT_9_), .SUM_6_(PRODUCT_8_), .SUM_5_(PRODUCT_7_) );
  ADDFHX4 S2_9_2 ( .A(ab_9__2_), .B(CARRYB_8__2_), .CI(SUMB_8__3_), .CO(
        CARRYB_9__2_), .S(SUMB_9__2_) );
  ADDFHX4 S2_15_1 ( .A(ab_15__1_), .B(CARRYB_14__1_), .CI(SUMB_14__2_), .CO(
        CARRYB_15__1_), .S(SUMB_15__1_) );
  ADDFHX4 S2_7_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  ADDFHX4 S2_11_4 ( .A(ab_11__4_), .B(CARRYB_10__4_), .CI(SUMB_10__5_), .CO(
        CARRYB_11__4_), .S(SUMB_11__4_) );
  ADDFHX4 S2_12_4 ( .A(ab_12__4_), .B(CARRYB_11__4_), .CI(SUMB_11__5_), .CO(
        CARRYB_12__4_), .S(SUMB_12__4_) );
  ADDFHX4 S2_8_1 ( .A(ab_8__1_), .B(CARRYB_7__1_), .CI(SUMB_7__2_), .CO(
        CARRYB_8__1_), .S(SUMB_8__1_) );
  ADDFHX4 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  ADDFHX4 S2_15_3 ( .A(ab_15__3_), .B(CARRYB_14__3_), .CI(SUMB_14__4_), .CO(
        CARRYB_15__3_), .S(SUMB_15__3_) );
  ADDFHX4 S2_8_5 ( .A(ab_8__5_), .B(CARRYB_7__5_), .CI(SUMB_7__6_), .CO(
        CARRYB_8__5_), .S(SUMB_8__5_) );
  ADDFHX4 S2_9_5 ( .A(ab_9__5_), .B(CARRYB_8__5_), .CI(SUMB_8__6_), .CO(
        CARRYB_9__5_), .S(SUMB_9__5_) );
  ADDFHX4 S4_2 ( .A(ab_16__2_), .B(CARRYB_15__2_), .CI(SUMB_15__3_), .CO(
        CARRYB_16__2_), .S(SUMB_16__2_) );
  ADDFHX4 S2_10_1 ( .A(ab_10__1_), .B(CARRYB_9__1_), .CI(SUMB_9__2_), .CO(
        CARRYB_10__1_), .S(SUMB_10__1_) );
  ADDFHX4 S2_11_1 ( .A(ab_11__1_), .B(CARRYB_10__1_), .CI(SUMB_10__2_), .CO(
        CARRYB_11__1_), .S(SUMB_11__1_) );
  ADDFHX4 S2_13_3 ( .A(ab_13__3_), .B(CARRYB_12__3_), .CI(SUMB_12__4_), .CO(
        CARRYB_13__3_), .S(SUMB_13__3_) );
  ADDFHX4 S2_14_3 ( .A(ab_14__3_), .B(CARRYB_13__3_), .CI(SUMB_13__4_), .CO(
        CARRYB_14__3_), .S(SUMB_14__3_) );
  ADDFHX4 S2_10_4 ( .A(ab_10__4_), .B(CARRYB_9__4_), .CI(SUMB_9__5_), .CO(
        CARRYB_10__4_), .S(SUMB_10__4_) );
  ADDFHX4 S1_9_0 ( .A(ab_9__0_), .B(CARRYB_8__0_), .CI(SUMB_8__1_), .CO(
        CARRYB_9__0_), .S(A1_7_) );
  ADDFHX4 S1_7_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(PROD1_7_) );
  ADDFHX4 S1_8_0 ( .A(ab_8__0_), .B(CARRYB_7__0_), .CI(SUMB_7__1_), .CO(
        CARRYB_8__0_), .S(A1_6_) );
  ADDFHX4 S2_14_2 ( .A(ab_14__2_), .B(CARRYB_13__2_), .CI(SUMB_13__3_), .CO(
        CARRYB_14__2_), .S(SUMB_14__2_) );
  ADDFHX4 S3_10_6 ( .A(ab_10__6_), .B(CARRYB_9__6_), .CI(ab_9__7_), .CO(
        CARRYB_10__6_), .S(SUMB_10__6_) );
  ADDFHX4 S5_6 ( .A(ab_16__6_), .B(CARRYB_15__6_), .CI(ab_15__7_), .CO(
        CARRYB_16__6_), .S(SUMB_16__6_) );
  ADDFHX4 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  ADDFHX4 S3_2_6 ( .A(ab_2__6_), .B(n6), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  ADDFHX4 S2_15_5 ( .A(ab_15__5_), .B(CARRYB_14__5_), .CI(SUMB_14__6_), .CO(
        CARRYB_15__5_), .S(SUMB_15__5_) );
  ADDFHX4 S4_4 ( .A(ab_16__4_), .B(CARRYB_15__4_), .CI(SUMB_15__5_), .CO(
        CARRYB_16__4_), .S(SUMB_16__4_) );
  ADDFHX4 S2_7_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  ADDFHX4 S3_8_6 ( .A(ab_8__6_), .B(CARRYB_7__6_), .CI(ab_7__7_), .CO(
        CARRYB_8__6_), .S(SUMB_8__6_) );
  ADDFHX4 S4_5 ( .A(ab_16__5_), .B(CARRYB_15__5_), .CI(SUMB_15__6_), .CO(
        CARRYB_16__5_), .S(SUMB_16__5_) );
  ADDFHX4 S4_1 ( .A(ab_16__1_), .B(CARRYB_15__1_), .CI(SUMB_15__2_), .CO(
        CARRYB_16__1_), .S(SUMB_16__1_) );
  ADDFHX4 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  ADDFHX4 S3_7_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(
        CARRYB_7__6_), .S(SUMB_7__6_) );
  ADDFHX4 S3_9_6 ( .A(ab_9__6_), .B(CARRYB_8__6_), .CI(ab_8__7_), .CO(
        CARRYB_9__6_), .S(SUMB_9__6_) );
  ADDFHX4 S4_3 ( .A(ab_16__3_), .B(CARRYB_15__3_), .CI(SUMB_15__4_), .CO(
        CARRYB_16__3_), .S(SUMB_16__3_) );
  ADDFHX4 S1_12_0 ( .A(ab_12__0_), .B(CARRYB_11__0_), .CI(SUMB_11__1_), .CO(
        CARRYB_12__0_), .S(A1_10_) );
  ADDFHX4 S1_15_0 ( .A(ab_15__0_), .B(CARRYB_14__0_), .CI(SUMB_14__1_), .CO(
        CARRYB_15__0_), .S(A1_13_) );
  ADDFHX4 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  ADDFHX4 S2_12_3 ( .A(ab_12__3_), .B(CARRYB_11__3_), .CI(SUMB_11__4_), .CO(
        CARRYB_12__3_), .S(SUMB_12__3_) );
  ADDFHX4 S2_11_5 ( .A(ab_11__5_), .B(CARRYB_10__5_), .CI(SUMB_10__6_), .CO(
        CARRYB_11__5_), .S(SUMB_11__5_) );
  ADDFHX4 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  ADDFHX4 S2_2_4 ( .A(ab_2__4_), .B(n9), .CI(SUMB_1__5_), .CO(CARRYB_2__4_), 
        .S(SUMB_2__4_) );
  ADDFHX4 S2_2_3 ( .A(ab_2__3_), .B(n10), .CI(SUMB_1__4_), .CO(CARRYB_2__3_), 
        .S(SUMB_2__3_) );
  ADDFHX4 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  ADDFHX4 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  ADDFHX4 S2_12_2 ( .A(ab_12__2_), .B(CARRYB_11__2_), .CI(SUMB_11__3_), .CO(
        CARRYB_12__2_), .S(SUMB_12__2_) );
  ADDFHX4 S2_13_2 ( .A(ab_13__2_), .B(CARRYB_12__2_), .CI(SUMB_12__3_), .CO(
        CARRYB_13__2_), .S(SUMB_13__2_) );
  ADDFHX4 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  ADDFHX4 S2_14_1 ( .A(ab_14__1_), .B(SUMB_13__2_), .CI(CARRYB_13__1_), .CO(
        CARRYB_14__1_), .S(SUMB_14__1_) );
  ADDFHX4 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  ADDFHX4 S2_11_3 ( .A(ab_11__3_), .B(CARRYB_10__3_), .CI(SUMB_10__4_), .CO(
        CARRYB_11__3_), .S(SUMB_11__3_) );
  ADDFHX4 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  ADDFHX4 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  ADDFHX4 S2_10_5 ( .A(ab_10__5_), .B(CARRYB_9__5_), .CI(SUMB_9__6_), .CO(
        CARRYB_10__5_), .S(SUMB_10__5_) );
  ADDFHX4 S2_8_3 ( .A(ab_8__3_), .B(CARRYB_7__3_), .CI(SUMB_7__4_), .CO(
        CARRYB_8__3_), .S(SUMB_8__3_) );
  ADDFHX4 S2_9_3 ( .A(ab_9__3_), .B(CARRYB_8__3_), .CI(SUMB_8__4_), .CO(
        CARRYB_9__3_), .S(SUMB_9__3_) );
  ADDFHX4 S2_9_4 ( .A(ab_9__4_), .B(CARRYB_8__4_), .CI(SUMB_8__5_), .CO(
        CARRYB_9__4_), .S(SUMB_9__4_) );
  ADDFHX4 S2_8_2 ( .A(ab_8__2_), .B(CARRYB_7__2_), .CI(SUMB_7__3_), .CO(
        CARRYB_8__2_), .S(SUMB_8__2_) );
  ADDFHX2 S2_14_5 ( .A(ab_14__5_), .B(CARRYB_13__5_), .CI(SUMB_13__6_), .CO(
        CARRYB_14__5_), .S(SUMB_14__5_) );
  ADDFHX4 S2_7_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  ADDFHX4 S2_8_4 ( .A(ab_8__4_), .B(CARRYB_7__4_), .CI(SUMB_7__5_), .CO(
        CARRYB_8__4_), .S(SUMB_8__4_) );
  ADDFHX4 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  ADDFHX4 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  ADDFHX4 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  ADDFHX4 S1_10_0 ( .A(ab_10__0_), .B(CARRYB_9__0_), .CI(SUMB_9__1_), .CO(
        CARRYB_10__0_), .S(A1_8_) );
  ADDFHX4 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  ADDFHX4 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  ADDFHX4 S2_10_2 ( .A(ab_10__2_), .B(CARRYB_9__2_), .CI(SUMB_9__3_), .CO(
        CARRYB_10__2_), .S(SUMB_10__2_) );
  ADDFHX4 S3_4_6 ( .A(ab_4__6_), .B(ab_3__7_), .CI(CARRYB_3__6_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  ADDFHX4 S2_2_5 ( .A(ab_2__5_), .B(n3), .CI(SUMB_1__6_), .CO(CARRYB_2__5_), 
        .S(SUMB_2__5_) );
  ADDFHX4 S2_13_5 ( .A(ab_13__5_), .B(CARRYB_12__5_), .CI(SUMB_12__6_), .CO(
        CARRYB_13__5_), .S(SUMB_13__5_) );
  ADDFHX4 S2_13_4 ( .A(ab_13__4_), .B(CARRYB_12__4_), .CI(SUMB_12__5_), .CO(
        CARRYB_13__4_), .S(SUMB_13__4_) );
  ADDFHX4 S2_14_4 ( .A(ab_14__4_), .B(CARRYB_13__4_), .CI(SUMB_13__5_), .CO(
        CARRYB_14__4_), .S(SUMB_14__4_) );
  ADDFHX4 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  ADDFHX4 S2_7_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  ADDFHX4 S3_11_6 ( .A(ab_11__6_), .B(CARRYB_10__6_), .CI(ab_10__7_), .CO(
        CARRYB_11__6_), .S(SUMB_11__6_) );
  ADDFHX4 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  ADDFHX4 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  ADDFHX4 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  ADDFHX4 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  ADDFHX4 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  ADDFHX4 S3_12_6 ( .A(ab_12__6_), .B(CARRYB_11__6_), .CI(ab_11__7_), .CO(
        CARRYB_12__6_), .S(SUMB_12__6_) );
  ADDFHX2 S3_13_6 ( .A(ab_13__6_), .B(CARRYB_12__6_), .CI(ab_12__7_), .CO(
        CARRYB_13__6_), .S(SUMB_13__6_) );
  ADDFHX4 S2_12_1 ( .A(ab_12__1_), .B(CARRYB_11__1_), .CI(SUMB_11__2_), .CO(
        CARRYB_12__1_), .S(SUMB_12__1_) );
  ADDFHX4 S2_9_1 ( .A(ab_9__1_), .B(CARRYB_8__1_), .CI(SUMB_8__2_), .CO(
        CARRYB_9__1_), .S(SUMB_9__1_) );
  ADDFHX4 S2_11_2 ( .A(ab_11__2_), .B(CARRYB_10__2_), .CI(SUMB_10__3_), .CO(
        CARRYB_11__2_), .S(SUMB_11__2_) );
  ADDFHX4 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  ADDFHX4 S4_0 ( .A(ab_16__0_), .B(CARRYB_15__0_), .CI(SUMB_15__1_), .CO(
        CARRYB_16__0_), .S(SUMB_16__0_) );
  ADDFHX4 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  ADDFHX4 S1_13_0 ( .A(ab_13__0_), .B(CARRYB_12__0_), .CI(SUMB_12__1_), .CO(
        CARRYB_13__0_), .S(A1_11_) );
  ADDFHX4 S1_14_0 ( .A(ab_14__0_), .B(CARRYB_13__0_), .CI(SUMB_13__1_), .CO(
        CARRYB_14__0_), .S(A1_12_) );
  ADDFHX4 S2_15_2 ( .A(ab_15__2_), .B(CARRYB_14__2_), .CI(SUMB_14__3_), .CO(
        CARRYB_15__2_), .S(SUMB_15__2_) );
  ADDFHX4 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  ADDFHX4 S2_7_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  ADDFHX4 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  ADDFHX4 S2_10_3 ( .A(ab_10__3_), .B(CARRYB_9__3_), .CI(SUMB_9__4_), .CO(
        CARRYB_10__3_), .S(SUMB_10__3_) );
  ADDFHX4 S2_2_1 ( .A(ab_2__1_), .B(n5), .CI(SUMB_1__2_), .CO(CARRYB_2__1_), 
        .S(SUMB_2__1_) );
  ADDFHX4 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  ADDFHX4 S1_11_0 ( .A(ab_11__0_), .B(CARRYB_10__0_), .CI(SUMB_10__1_), .CO(
        CARRYB_11__0_), .S(A1_9_) );
  ADDFHX4 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  ADDFHX4 S2_12_5 ( .A(ab_12__5_), .B(CARRYB_11__5_), .CI(SUMB_11__6_), .CO(
        CARRYB_12__5_), .S(SUMB_12__5_) );
  ADDFHX2 S2_15_4 ( .A(ab_15__4_), .B(CARRYB_14__4_), .CI(SUMB_14__5_), .CO(
        CARRYB_15__4_), .S(SUMB_15__4_) );
  ADDFHX2 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  ADDFHX4 S3_14_6 ( .A(ab_14__6_), .B(CARRYB_13__6_), .CI(ab_13__7_), .CO(
        CARRYB_14__6_), .S(SUMB_14__6_) );
  ADDFHX4 S3_15_6 ( .A(ab_15__6_), .B(CARRYB_14__6_), .CI(ab_14__7_), .CO(
        CARRYB_15__6_), .S(SUMB_15__6_) );
  ADDFHX2 S2_13_1 ( .A(ab_13__1_), .B(CARRYB_12__1_), .CI(SUMB_12__2_), .CO(
        CARRYB_13__1_), .S(SUMB_13__1_) );
  NOR2BX1 U2 ( .AN(A[5]), .B(n18), .Y(ab_5__5_) );
  NOR2BX2 U3 ( .AN(A[5]), .B(n33), .Y(ab_5__4_) );
  AND2X4 U4 ( .A(ab_1__5_), .B(ab_0__6_), .Y(n3) );
  NOR2BX1 U5 ( .AN(A[7]), .B(n36), .Y(ab_7__1_) );
  NOR2BX2 U6 ( .AN(A[9]), .B(n19), .Y(ab_9__5_) );
  NOR2BX2 U7 ( .AN(A[8]), .B(n23), .Y(ab_8__2_) );
  NOR2BX1 U8 ( .AN(A[8]), .B(n27), .Y(ab_8__0_) );
  NOR2BX2 U9 ( .AN(A[7]), .B(n21), .Y(ab_7__3_) );
  NOR2BX2 U10 ( .AN(A[6]), .B(n26), .Y(ab_6__6_) );
  NOR2BX2 U11 ( .AN(A[6]), .B(n23), .Y(ab_6__2_) );
  CLKINVX3 U12 ( .A(B[2]), .Y(n35) );
  NOR2BX1 U13 ( .AN(A[10]), .B(n27), .Y(ab_10__0_) );
  NOR2BX2 U14 ( .AN(A[4]), .B(n26), .Y(ab_4__6_) );
  NOR2BX2 U15 ( .AN(A[8]), .B(n21), .Y(ab_8__3_) );
  NOR2BX2 U16 ( .AN(A[9]), .B(n25), .Y(ab_9__1_) );
  NOR2BX1 U17 ( .AN(A[16]), .B(n24), .Y(ab_16__2_) );
  NOR2BX1 U18 ( .AN(A[9]), .B(n27), .Y(ab_9__0_) );
  NOR2BX2 U19 ( .AN(A[13]), .B(n28), .Y(ab_13__0_) );
  NOR2BXL U20 ( .AN(A[16]), .B(n25), .Y(ab_16__1_) );
  NOR2BX1 U21 ( .AN(A[5]), .B(n36), .Y(ab_5__1_) );
  INVX4 U23 ( .A(B[1]), .Y(n36) );
  BUFX1 U24 ( .A(n36), .Y(n25) );
  AND2X4 U25 ( .A(ab_0__2_), .B(n38), .Y(n5) );
  INVX2 U26 ( .A(B[4]), .Y(n33) );
  CLKBUFX2 U27 ( .A(n33), .Y(n20) );
  AND2X4 U28 ( .A(ab_0__7_), .B(ab_1__6_), .Y(n6) );
  NAND2X4 U29 ( .A(ab_0__3_), .B(ab_1__2_), .Y(n17) );
  NOR2BX2 U30 ( .AN(B[3]), .B(n29), .Y(ab_0__3_) );
  CLKINVX4 U31 ( .A(B[3]), .Y(n34) );
  INVX4 U32 ( .A(B[5]), .Y(n32) );
  AND2X4 U33 ( .A(B[5]), .B(n7), .Y(ab_0__5_) );
  NOR2BX2 U34 ( .AN(A[4]), .B(n21), .Y(ab_4__3_) );
  NOR2BX2 U35 ( .AN(A[4]), .B(n23), .Y(ab_4__2_) );
  NOR2BX2 U36 ( .AN(A[4]), .B(n33), .Y(ab_4__4_) );
  NOR2BX2 U37 ( .AN(A[4]), .B(n36), .Y(ab_4__1_) );
  INVX12 U38 ( .A(A[0]), .Y(n29) );
  NOR2BX2 U39 ( .AN(B[2]), .B(n29), .Y(ab_0__2_) );
  BUFX16 U40 ( .A(n35), .Y(n23) );
  BUFX20 U41 ( .A(n31), .Y(n26) );
  NOR2BX2 U42 ( .AN(A[2]), .B(n18), .Y(ab_2__5_) );
  NOR2BX2 U43 ( .AN(A[2]), .B(n26), .Y(ab_2__6_) );
  NOR2BX4 U44 ( .AN(A[2]), .B(n23), .Y(ab_2__2_) );
  NOR2BX4 U45 ( .AN(A[2]), .B(n21), .Y(ab_2__3_) );
  NOR2BX4 U46 ( .AN(A[2]), .B(n33), .Y(ab_2__4_) );
  AND2X4 U47 ( .A(A[1]), .B(B[4]), .Y(ab_1__4_) );
  NOR2BXL U48 ( .AN(A[0]), .B(n27), .Y(n30) );
  AND3X1 U49 ( .A(A[1]), .B(B[1]), .C(n30), .Y(CARRYB_1__0_) );
  NOR2BX4 U50 ( .AN(B[7]), .B(n29), .Y(ab_0__7_) );
  INVX4 U51 ( .A(n21), .Y(n8) );
  BUFX16 U52 ( .A(n34), .Y(n21) );
  NOR2BX4 U53 ( .AN(B[4]), .B(n29), .Y(ab_0__4_) );
  NOR2BX2 U54 ( .AN(A[3]), .B(n23), .Y(ab_3__2_) );
  CLKINVX20 U55 ( .A(n29), .Y(n7) );
  AND2X4 U56 ( .A(A[1]), .B(n8), .Y(ab_1__3_) );
  NOR2BX2 U57 ( .AN(A[2]), .B(n27), .Y(ab_2__0_) );
  XOR2X4 U58 ( .A(n38), .B(ab_0__2_), .Y(SUMB_1__1_) );
  AND2X4 U59 ( .A(ab_1__4_), .B(ab_0__5_), .Y(n9) );
  NOR2BX1 U60 ( .AN(A[6]), .B(n21), .Y(ab_6__3_) );
  XOR2X4 U61 ( .A(ab_1__4_), .B(ab_0__5_), .Y(SUMB_1__4_) );
  NOR2BX1 U62 ( .AN(A[3]), .B(n37), .Y(ab_3__7_) );
  NOR2BX1 U63 ( .AN(A[3]), .B(n26), .Y(ab_3__6_) );
  NOR2BX1 U64 ( .AN(A[3]), .B(n27), .Y(ab_3__0_) );
  NOR2BX1 U65 ( .AN(A[3]), .B(n21), .Y(ab_3__3_) );
  NOR2BX1 U66 ( .AN(A[3]), .B(n33), .Y(ab_3__4_) );
  NOR2BX2 U67 ( .AN(A[3]), .B(n18), .Y(ab_3__5_) );
  XOR2X4 U68 ( .A(ab_1__2_), .B(ab_0__3_), .Y(SUMB_1__2_) );
  INVX4 U69 ( .A(n17), .Y(CARRYB_1__2_) );
  AND2X4 U70 ( .A(ab_0__4_), .B(ab_1__3_), .Y(n10) );
  XOR2X4 U71 ( .A(ab_1__3_), .B(ab_0__4_), .Y(SUMB_1__3_) );
  XOR2X4 U72 ( .A(ab_1__5_), .B(ab_0__6_), .Y(SUMB_1__5_) );
  NOR2BX4 U73 ( .AN(B[6]), .B(n29), .Y(ab_0__6_) );
  NOR2BX2 U74 ( .AN(A[2]), .B(n36), .Y(ab_2__1_) );
  NOR2BX1 U75 ( .AN(A[3]), .B(n36), .Y(ab_3__1_) );
  XOR2X4 U76 ( .A(ab_1__6_), .B(ab_0__7_), .Y(SUMB_1__6_) );
  AND2X4 U77 ( .A(A[1]), .B(B[6]), .Y(ab_1__6_) );
  XOR2X4 U78 ( .A(CARRYB_16__4_), .B(SUMB_16__5_), .Y(A1_19_) );
  NOR2BX4 U79 ( .AN(A[1]), .B(n36), .Y(n38) );
  NOR2BX2 U80 ( .AN(A[5]), .B(n26), .Y(ab_5__6_) );
  NOR2BX1 U81 ( .AN(A[4]), .B(n27), .Y(ab_4__0_) );
  NOR2BX4 U82 ( .AN(A[1]), .B(n23), .Y(ab_1__2_) );
  NOR2BX4 U83 ( .AN(A[1]), .B(n18), .Y(ab_1__5_) );
  AND2X4 U84 ( .A(SUMB_16__1_), .B(CARRYB_16__0_), .Y(n13) );
  AND2X4 U85 ( .A(SUMB_16__2_), .B(CARRYB_16__1_), .Y(n12) );
  INVX8 U86 ( .A(B[0]), .Y(n27) );
  NOR2BXL U87 ( .AN(A[7]), .B(n23), .Y(ab_7__2_) );
  NOR2BX4 U88 ( .AN(A[9]), .B(n26), .Y(ab_9__6_) );
  NOR2BX1 U89 ( .AN(A[8]), .B(n37), .Y(ab_8__7_) );
  NOR2BX1 U90 ( .AN(A[6]), .B(n27), .Y(ab_6__0_) );
  NOR2BX2 U91 ( .AN(A[8]), .B(n36), .Y(ab_8__1_) );
  NOR2BXL U92 ( .AN(A[7]), .B(n27), .Y(ab_7__0_) );
  NOR2BX1 U93 ( .AN(A[5]), .B(n21), .Y(ab_5__3_) );
  NOR2BX1 U94 ( .AN(A[4]), .B(n37), .Y(ab_4__7_) );
  NOR2BX1 U95 ( .AN(A[2]), .B(n37), .Y(ab_2__7_) );
  INVXL U96 ( .A(B[0]), .Y(n28) );
  CLKBUFXL U97 ( .A(n34), .Y(n22) );
  INVX16 U98 ( .A(B[7]), .Y(n37) );
  NOR2BX1 U99 ( .AN(A[11]), .B(n19), .Y(ab_11__5_) );
  NOR2BX1 U100 ( .AN(A[10]), .B(n19), .Y(ab_10__5_) );
  NOR2BX1 U101 ( .AN(A[7]), .B(n26), .Y(ab_7__6_) );
  NOR2BX1 U102 ( .AN(A[4]), .B(n18), .Y(ab_4__5_) );
  NOR2BX1 U103 ( .AN(A[5]), .B(n23), .Y(ab_5__2_) );
  NOR2BX1 U104 ( .AN(A[11]), .B(n22), .Y(ab_11__3_) );
  NOR2BX1 U105 ( .AN(A[11]), .B(n20), .Y(ab_11__4_) );
  NOR2BX1 U106 ( .AN(A[11]), .B(n24), .Y(ab_11__2_) );
  NOR2BX1 U107 ( .AN(A[10]), .B(n24), .Y(ab_10__2_) );
  NOR2BX1 U108 ( .AN(A[10]), .B(n22), .Y(ab_10__3_) );
  NOR2BX1 U109 ( .AN(A[10]), .B(n25), .Y(ab_10__1_) );
  NOR2BX1 U110 ( .AN(A[11]), .B(n25), .Y(ab_11__1_) );
  NOR2BX1 U111 ( .AN(A[16]), .B(n22), .Y(ab_16__3_) );
  NOR2BX1 U112 ( .AN(A[15]), .B(n19), .Y(ab_15__5_) );
  NOR2BX1 U113 ( .AN(A[15]), .B(n20), .Y(ab_15__4_) );
  NOR2BX1 U114 ( .AN(A[15]), .B(n25), .Y(ab_15__1_) );
  NOR2BX1 U115 ( .AN(A[15]), .B(n22), .Y(ab_15__3_) );
  NOR2BX1 U116 ( .AN(A[15]), .B(n28), .Y(ab_15__0_) );
  BUFX12 U117 ( .A(n32), .Y(n18) );
  CLKBUFXL U118 ( .A(n32), .Y(n19) );
  INVX4 U119 ( .A(B[6]), .Y(n31) );
  BUFX3 U120 ( .A(n35), .Y(n24) );
  NOR2BXL U121 ( .AN(A[14]), .B(n25), .Y(ab_14__1_) );
  NOR2BXL U122 ( .AN(A[13]), .B(n24), .Y(ab_13__2_) );
  NOR2BXL U123 ( .AN(A[12]), .B(n22), .Y(ab_12__3_) );
  NOR2BXL U124 ( .AN(A[9]), .B(n37), .Y(ab_9__7_) );
  NOR2BX1 U125 ( .AN(A[10]), .B(n26), .Y(ab_10__6_) );
  NOR2BXL U126 ( .AN(A[7]), .B(n18), .Y(ab_7__5_) );
  NOR2BXL U127 ( .AN(A[14]), .B(n28), .Y(ab_14__0_) );
  NOR2BXL U128 ( .AN(A[13]), .B(n25), .Y(ab_13__1_) );
  NOR2BXL U129 ( .AN(A[12]), .B(n24), .Y(ab_12__2_) );
  NOR2BXL U130 ( .AN(A[12]), .B(n27), .Y(ab_12__0_) );
  NOR2BXL U131 ( .AN(A[11]), .B(n27), .Y(ab_11__0_) );
  NOR2BXL U132 ( .AN(A[8]), .B(n20), .Y(ab_8__4_) );
  NOR2BXL U133 ( .AN(A[14]), .B(n20), .Y(ab_14__4_) );
  NOR2BXL U134 ( .AN(A[7]), .B(n37), .Y(ab_7__7_) );
  NOR2BX2 U135 ( .AN(A[8]), .B(n26), .Y(ab_8__6_) );
  NOR2BXL U136 ( .AN(A[6]), .B(n37), .Y(ab_6__7_) );
  NOR2BXL U137 ( .AN(A[6]), .B(n18), .Y(ab_6__5_) );
  NOR2BXL U138 ( .AN(A[5]), .B(n37), .Y(ab_5__7_) );
  NOR2BXL U139 ( .AN(A[13]), .B(n37), .Y(ab_13__7_) );
  NOR2BXL U140 ( .AN(A[14]), .B(n26), .Y(ab_14__6_) );
  NOR2BXL U141 ( .AN(A[12]), .B(n25), .Y(ab_12__1_) );
  NOR2BXL U142 ( .AN(A[13]), .B(n20), .Y(ab_13__4_) );
  NOR2BXL U143 ( .AN(A[7]), .B(n20), .Y(ab_7__4_) );
  NOR2BXL U144 ( .AN(A[14]), .B(n19), .Y(ab_14__5_) );
  NOR2BXL U145 ( .AN(A[6]), .B(n25), .Y(ab_6__1_) );
  NOR2BXL U146 ( .AN(A[12]), .B(n37), .Y(ab_12__7_) );
  NOR2BXL U147 ( .AN(A[13]), .B(n26), .Y(ab_13__6_) );
  AND2X2 U148 ( .A(CARRYB_16__2_), .B(SUMB_16__3_), .Y(n11) );
  XOR2X2 U149 ( .A(CARRYB_16__5_), .B(SUMB_16__6_), .Y(A1_20_) );
  NOR2BXL U150 ( .AN(A[14]), .B(n24), .Y(ab_14__2_) );
  NOR2BXL U151 ( .AN(A[13]), .B(n22), .Y(ab_13__3_) );
  NOR2BX1 U152 ( .AN(A[10]), .B(n20), .Y(ab_10__4_) );
  NOR2BXL U153 ( .AN(A[8]), .B(n18), .Y(ab_8__5_) );
  NOR2BXL U154 ( .AN(A[12]), .B(n20), .Y(ab_12__4_) );
  NOR2BXL U155 ( .AN(A[13]), .B(n19), .Y(ab_13__5_) );
  NOR2BXL U156 ( .AN(A[6]), .B(n33), .Y(ab_6__4_) );
  NOR2BXL U157 ( .AN(A[11]), .B(n37), .Y(ab_11__7_) );
  NOR2BXL U158 ( .AN(A[12]), .B(n26), .Y(ab_12__6_) );
  AND2X2 U159 ( .A(CARRYB_16__3_), .B(SUMB_16__4_), .Y(n14) );
  AND2X2 U160 ( .A(CARRYB_16__4_), .B(SUMB_16__5_), .Y(n15) );
  NOR2BXL U161 ( .AN(A[14]), .B(n22), .Y(ab_14__3_) );
  NOR2BXL U162 ( .AN(A[10]), .B(n37), .Y(ab_10__7_) );
  NOR2BXL U163 ( .AN(A[11]), .B(n26), .Y(ab_11__6_) );
  NOR2BXL U164 ( .AN(A[12]), .B(n19), .Y(ab_12__5_) );
  XOR2X1 U165 ( .A(CARRYB_16__6_), .B(ab_16__7_), .Y(A1_21_) );
  AND2X2 U166 ( .A(CARRYB_16__5_), .B(SUMB_16__6_), .Y(n16) );
  NOR2BX1 U167 ( .AN(A[16]), .B(n20), .Y(ab_16__4_) );
  NOR2BX1 U168 ( .AN(A[16]), .B(n19), .Y(ab_16__5_) );
  NOR2BXL U169 ( .AN(A[16]), .B(n26), .Y(ab_16__6_) );
  NOR2BXL U170 ( .AN(A[15]), .B(n37), .Y(ab_15__7_) );
  NOR2BX2 U171 ( .AN(A[16]), .B(n28), .Y(ab_16__0_) );
  NOR2BXL U172 ( .AN(A[14]), .B(n37), .Y(ab_14__7_) );
  NOR2BXL U173 ( .AN(A[15]), .B(n26), .Y(ab_15__6_) );
  NOR2BXL U174 ( .AN(A[15]), .B(n24), .Y(ab_15__2_) );
  NOR2BXL U175 ( .AN(A[16]), .B(n37), .Y(ab_16__7_) );
  XOR2X4 U176 ( .A(CARRYB_16__1_), .B(SUMB_16__2_), .Y(A1_16_) );
  XOR2X4 U177 ( .A(SUMB_16__3_), .B(CARRYB_16__2_), .Y(A1_17_) );
  XOR2X4 U178 ( .A(SUMB_16__4_), .B(CARRYB_16__3_), .Y(A1_18_) );
  XOR2X4 U179 ( .A(CARRYB_16__0_), .B(SUMB_16__1_), .Y(A1_15_) );
  NOR2BX1 U180 ( .AN(A[1]), .B(n37), .Y(ab_1__7_) );
  NOR2BX4 U181 ( .AN(A[5]), .B(n27), .Y(ab_5__0_) );
  NOR2BX4 U182 ( .AN(A[9]), .B(n20), .Y(ab_9__4_) );
  NOR2BX4 U183 ( .AN(A[9]), .B(n22), .Y(ab_9__3_) );
  NOR2BX4 U184 ( .AN(A[9]), .B(n24), .Y(ab_9__2_) );
endmodule


module multi16_3 ( in_17bit, in_8bit, out );
  input [16:0] in_17bit;
  input [7:0] in_8bit;
  output [16:0] out;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120;
  wire   [16:1] in_17bit_b;
  wire   [7:1] in_8bit_b;
  wire   [23:8] mul;

  multi16_3_DW02_mult_0 mult_55 ( .A({in_17bit_b[16:3], n3, n40, in_17bit[0]}), 
        .B({in_8bit_b, n41}), .PRODUCT_23_(mul[23]), .PRODUCT_22_(mul[22]), 
        .PRODUCT_21_(mul[21]), .PRODUCT_20_(mul[20]), .PRODUCT_19_(mul[19]), 
        .PRODUCT_18_(mul[18]), .PRODUCT_17_(mul[17]), .PRODUCT_16_(mul[16]), 
        .PRODUCT_15_(mul[15]), .PRODUCT_14_(mul[14]), .PRODUCT_13_(mul[13]), 
        .PRODUCT_12_(mul[12]), .PRODUCT_11_(mul[11]), .PRODUCT_10_(mul[10]), 
        .PRODUCT_9_(mul[9]), .PRODUCT_8_(mul[8]), .PRODUCT_7_(out[0]) );
  BUFX16 U2 ( .A(n17), .Y(n1) );
  BUFX8 U3 ( .A(n17), .Y(n20) );
  BUFX16 U4 ( .A(in_17bit[16]), .Y(n17) );
  INVX8 U5 ( .A(n115), .Y(n119) );
  OR2X4 U6 ( .A(n38), .B(n92), .Y(n30) );
  NOR2X1 U7 ( .A(n37), .B(n92), .Y(n79) );
  INVX12 U8 ( .A(n17), .Y(n92) );
  CLKINVX2 U9 ( .A(mul[17]), .Y(n9) );
  NOR2X4 U10 ( .A(mul[16]), .B(n105), .Y(n2) );
  INVXL U11 ( .A(in_17bit[9]), .Y(n78) );
  NAND2X2 U12 ( .A(n1), .B(n63), .Y(n19) );
  BUFX12 U13 ( .A(in_17bit_b[2]), .Y(n3) );
  AND2X2 U14 ( .A(out[0]), .B(n111), .Y(n21) );
  AOI21X2 U15 ( .A0(n4), .A1(n46), .B0(n44), .Y(n53) );
  INVX4 U16 ( .A(n42), .Y(n41) );
  INVX2 U17 ( .A(n67), .Y(n32) );
  NOR2X4 U18 ( .A(in_8bit[3]), .B(n51), .Y(n4) );
  NOR2X4 U19 ( .A(in_17bit[1]), .B(in_17bit[0]), .Y(n5) );
  XNOR2X2 U20 ( .A(in_8bit[3]), .B(n26), .Y(in_8bit_b[3]) );
  NAND2X1 U21 ( .A(n1), .B(n66), .Y(n65) );
  NAND2X2 U22 ( .A(n43), .B(n51), .Y(n26) );
  CLKINVX4 U23 ( .A(in_8bit[5]), .Y(n54) );
  BUFX16 U24 ( .A(in_17bit_b[1]), .Y(n40) );
  OR2X4 U25 ( .A(in_17bit[1]), .B(in_17bit[0]), .Y(n6) );
  INVX8 U26 ( .A(in_17bit[1]), .Y(n14) );
  CLKINVX8 U27 ( .A(n14), .Y(n15) );
  NOR2BX4 U28 ( .AN(n16), .B(mul[20]), .Y(n114) );
  CLKINVX8 U29 ( .A(in_8bit[2]), .Y(n50) );
  AOI21X1 U30 ( .A0(n119), .A1(n118), .B0(n117), .Y(n120) );
  INVX8 U31 ( .A(in_8bit[4]), .Y(n46) );
  XOR2X2 U32 ( .A(mul[23]), .B(n120), .Y(out[16]) );
  NAND2BX4 U33 ( .AN(mul[21]), .B(n114), .Y(n115) );
  XOR2X4 U34 ( .A(n7), .B(mul[21]), .Y(out[14]) );
  NOR2X4 U35 ( .A(n114), .B(n117), .Y(n7) );
  XNOR2X2 U36 ( .A(n52), .B(n46), .Y(in_8bit_b[4]) );
  INVX8 U37 ( .A(in_17bit[2]), .Y(n62) );
  NOR3X2 U38 ( .A(in_8bit[6]), .B(n57), .C(n45), .Y(in_8bit_b[7]) );
  NAND2X4 U39 ( .A(n101), .B(n111), .Y(n100) );
  NOR2X4 U40 ( .A(n58), .B(n14), .Y(n60) );
  BUFX8 U41 ( .A(mul[19]), .Y(n8) );
  NAND2X2 U42 ( .A(mul[17]), .B(n106), .Y(n11) );
  NAND2X4 U43 ( .A(n9), .B(n10), .Y(n12) );
  NAND2X4 U44 ( .A(n11), .B(n12), .Y(out[10]) );
  INVX4 U45 ( .A(n106), .Y(n10) );
  XOR2X4 U46 ( .A(mul[15]), .B(n27), .Y(out[8]) );
  AND2X4 U47 ( .A(n113), .B(n111), .Y(n110) );
  NAND2XL U48 ( .A(n1), .B(n82), .Y(n81) );
  XNOR2X1 U49 ( .A(n1), .B(n43), .Y(n117) );
  NAND2XL U50 ( .A(n1), .B(n77), .Y(n76) );
  NAND2XL U51 ( .A(n1), .B(n70), .Y(n69) );
  BUFX4 U52 ( .A(mul[20]), .Y(n13) );
  OR2X4 U53 ( .A(mul[10]), .B(n95), .Y(n96) );
  CLKINVX2 U54 ( .A(n98), .Y(n99) );
  CLKINVX8 U55 ( .A(n18), .Y(in_17bit_b[3]) );
  NAND2X4 U56 ( .A(n17), .B(in_17bit[0]), .Y(n58) );
  CLKINVX8 U57 ( .A(in_8bit[0]), .Y(n42) );
  XNOR2X4 U58 ( .A(n13), .B(n112), .Y(out[13]) );
  OAI21X2 U59 ( .A0(n113), .A1(mul[19]), .B0(n111), .Y(n112) );
  NAND2X4 U60 ( .A(n38), .B(n64), .Y(n66) );
  NOR2X4 U61 ( .A(in_17bit[3]), .B(n63), .Y(n38) );
  NOR2X4 U62 ( .A(n20), .B(n15), .Y(n59) );
  NAND2X4 U63 ( .A(n1), .B(n6), .Y(n61) );
  XOR2X4 U64 ( .A(in_17bit[3]), .B(n19), .Y(n18) );
  NAND2X4 U65 ( .A(n62), .B(n5), .Y(n63) );
  NOR2X4 U66 ( .A(mul[19]), .B(n113), .Y(n16) );
  OAI21X2 U67 ( .A0(n41), .A1(in_8bit[1]), .B0(n43), .Y(n49) );
  NAND2X4 U68 ( .A(n43), .B(n57), .Y(n55) );
  XOR2X4 U69 ( .A(mul[8]), .B(n21), .Y(out[1]) );
  INVX8 U70 ( .A(n45), .Y(n43) );
  INVX8 U71 ( .A(in_8bit[7]), .Y(n45) );
  OR2X4 U72 ( .A(mul[18]), .B(n109), .Y(n113) );
  NOR3X4 U73 ( .A(n59), .B(n60), .C(n5), .Y(in_17bit_b[1]) );
  NAND2X1 U74 ( .A(n35), .B(n90), .Y(n93) );
  CLKINVX8 U75 ( .A(in_17bit[8]), .Y(n74) );
  CLKINVX4 U76 ( .A(in_17bit[13]), .Y(n88) );
  OR2X4 U77 ( .A(mul[8]), .B(out[0]), .Y(n94) );
  OR2X4 U78 ( .A(mul[14]), .B(n101), .Y(n102) );
  CLKINVX3 U79 ( .A(in_17bit[11]), .Y(n83) );
  CLKINVX8 U80 ( .A(in_17bit[12]), .Y(n85) );
  XNOR2X4 U81 ( .A(mul[13]), .B(n24), .Y(out[6]) );
  XNOR2X4 U82 ( .A(mul[9]), .B(n23), .Y(out[2]) );
  XOR2X4 U83 ( .A(n29), .B(n68), .Y(in_17bit_b[6]) );
  OR2X4 U84 ( .A(n31), .B(n92), .Y(n29) );
  NAND2X4 U85 ( .A(n94), .B(n111), .Y(n23) );
  XNOR2X2 U86 ( .A(mul[11]), .B(n22), .Y(out[4]) );
  NAND2X2 U87 ( .A(n96), .B(n111), .Y(n22) );
  AND2X4 U88 ( .A(n102), .B(n111), .Y(n27) );
  NAND2X4 U89 ( .A(n98), .B(n111), .Y(n24) );
  INVXL U90 ( .A(in_8bit[6]), .Y(n56) );
  XOR2X2 U91 ( .A(n33), .B(n90), .Y(in_17bit_b[14]) );
  NAND2X2 U92 ( .A(n37), .B(n80), .Y(n82) );
  OR2X4 U93 ( .A(mul[9]), .B(n94), .Y(n95) );
  OR2X4 U94 ( .A(mul[11]), .B(n96), .Y(n97) );
  OR2X4 U95 ( .A(mul[16]), .B(n105), .Y(n107) );
  XNOR2X4 U96 ( .A(mul[12]), .B(n25), .Y(out[5]) );
  NAND2X4 U97 ( .A(n97), .B(n111), .Y(n25) );
  NAND3X4 U98 ( .A(n4), .B(n46), .C(n54), .Y(n57) );
  INVXL U99 ( .A(in_8bit[7]), .Y(n44) );
  INVX4 U100 ( .A(n117), .Y(n111) );
  XOR2X4 U101 ( .A(n61), .B(n62), .Y(in_17bit_b[2]) );
  NOR2X4 U102 ( .A(n66), .B(n32), .Y(n31) );
  NAND2X4 U103 ( .A(n75), .B(n74), .Y(n77) );
  NOR2XL U104 ( .A(n77), .B(in_17bit[9]), .Y(n37) );
  NAND2XL U105 ( .A(n41), .B(n43), .Y(n47) );
  XOR2X2 U106 ( .A(n88), .B(n86), .Y(in_17bit_b[13]) );
  NAND2XL U107 ( .A(n1), .B(n87), .Y(n86) );
  XOR2X2 U108 ( .A(n34), .B(n85), .Y(in_17bit_b[12]) );
  AND2X4 U109 ( .A(n89), .B(n88), .Y(n35) );
  AND2X4 U110 ( .A(n84), .B(n83), .Y(n36) );
  OR2X4 U111 ( .A(mul[12]), .B(n97), .Y(n98) );
  XOR2X4 U112 ( .A(mul[10]), .B(n28), .Y(out[3]) );
  AND2X4 U113 ( .A(n95), .B(n111), .Y(n28) );
  XOR2X4 U114 ( .A(n30), .B(n64), .Y(in_17bit_b[4]) );
  XOR2X2 U115 ( .A(n49), .B(n50), .Y(in_8bit_b[2]) );
  NAND2X2 U116 ( .A(n31), .B(n68), .Y(n70) );
  INVXL U117 ( .A(in_8bit[1]), .Y(n48) );
  NAND2BX4 U118 ( .AN(n70), .B(n71), .Y(n72) );
  OR2XL U119 ( .A(n35), .B(n92), .Y(n33) );
  OR2XL U120 ( .A(n36), .B(n92), .Y(n34) );
  XOR2X1 U121 ( .A(n83), .B(n81), .Y(in_17bit_b[11]) );
  XOR2X1 U122 ( .A(n78), .B(n76), .Y(in_17bit_b[9]) );
  NAND2X1 U123 ( .A(n36), .B(n85), .Y(n87) );
  XNOR2X2 U124 ( .A(n91), .B(n39), .Y(in_17bit_b[15]) );
  AND2X1 U125 ( .A(n1), .B(n93), .Y(n39) );
  INVX1 U126 ( .A(in_17bit[10]), .Y(n80) );
  XNOR2X4 U127 ( .A(mul[18]), .B(n108), .Y(out[11]) );
  NOR2X4 U128 ( .A(n119), .B(n117), .Y(n116) );
  INVX8 U129 ( .A(mul[22]), .Y(n118) );
  XOR2X4 U130 ( .A(n48), .B(n47), .Y(in_8bit_b[1]) );
  NAND3BX4 U131 ( .AN(in_8bit[1]), .B(n50), .C(n42), .Y(n51) );
  NOR2X4 U132 ( .A(n4), .B(n44), .Y(n52) );
  XNOR2X4 U133 ( .A(n53), .B(n54), .Y(in_8bit_b[5]) );
  XOR2X4 U134 ( .A(n56), .B(n55), .Y(in_8bit_b[6]) );
  CLKINVX3 U135 ( .A(in_17bit[4]), .Y(n64) );
  CLKINVX3 U136 ( .A(in_17bit[5]), .Y(n67) );
  XOR2X4 U137 ( .A(n67), .B(n65), .Y(in_17bit_b[5]) );
  CLKINVX3 U138 ( .A(in_17bit[6]), .Y(n68) );
  CLKINVX3 U139 ( .A(in_17bit[7]), .Y(n71) );
  XOR2X4 U140 ( .A(n71), .B(n69), .Y(in_17bit_b[7]) );
  CLKINVX3 U141 ( .A(n72), .Y(n75) );
  NOR2X4 U142 ( .A(n75), .B(n92), .Y(n73) );
  XNOR2X4 U143 ( .A(n73), .B(n74), .Y(in_17bit_b[8]) );
  XNOR2X4 U144 ( .A(n79), .B(n80), .Y(in_17bit_b[10]) );
  CLKINVX3 U145 ( .A(n82), .Y(n84) );
  CLKINVX3 U146 ( .A(n87), .Y(n89) );
  CLKINVX3 U147 ( .A(in_17bit[14]), .Y(n90) );
  CLKINVX3 U148 ( .A(in_17bit[15]), .Y(n91) );
  NOR3X4 U149 ( .A(in_17bit[15]), .B(n93), .C(n92), .Y(in_17bit_b[16]) );
  NAND2BX4 U150 ( .AN(mul[13]), .B(n99), .Y(n101) );
  XNOR2X4 U151 ( .A(mul[14]), .B(n100), .Y(out[7]) );
  CLKINVX3 U152 ( .A(n102), .Y(n103) );
  NAND2BX4 U153 ( .AN(mul[15]), .B(n103), .Y(n105) );
  NAND2X4 U154 ( .A(n105), .B(n111), .Y(n104) );
  XNOR2X4 U155 ( .A(mul[16]), .B(n104), .Y(out[9]) );
  NAND2X4 U156 ( .A(n107), .B(n111), .Y(n106) );
  NAND2BX4 U157 ( .AN(mul[17]), .B(n2), .Y(n109) );
  NAND2X4 U158 ( .A(n109), .B(n111), .Y(n108) );
  XOR2X4 U159 ( .A(n110), .B(n8), .Y(out[12]) );
  XNOR2X4 U160 ( .A(n116), .B(n118), .Y(out[15]) );
endmodule


module multi16_2_DW01_add_0 ( A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, 
        A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, 
        B_20_, B_19_, B_18_, B_17_, B_16_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, 
        SUM_17_, SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, 
        SUM_9_, SUM_8_, SUM_7_, SUM_6_, SUM_5_ );
  input A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_,
         A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, B_20_, B_19_,
         B_18_, B_17_, B_16_;
  output SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, SUM_15_,
         SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, SUM_7_,
         SUM_6_, SUM_5_;
  wire   n43, n1, n3, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42;

  OAI21X1 U2 ( .A0(n30), .A1(n34), .B0(n3), .Y(n32) );
  BUFX8 U3 ( .A(B_19_), .Y(n1) );
  BUFX8 U4 ( .A(A_14_), .Y(SUM_14_) );
  INVX1 U5 ( .A(n33), .Y(n17) );
  BUFX8 U6 ( .A(A_15_), .Y(SUM_15_) );
  CLKINVX3 U7 ( .A(n18), .Y(n3) );
  NAND2X4 U8 ( .A(n33), .B(n16), .Y(n39) );
  BUFX12 U9 ( .A(A_13_), .Y(SUM_13_) );
  INVX4 U10 ( .A(n34), .Y(n20) );
  BUFX16 U11 ( .A(n43), .Y(SUM_17_) );
  OAI21X4 U12 ( .A0(n27), .A1(n28), .B0(n29), .Y(n23) );
  INVX8 U13 ( .A(n35), .Y(n18) );
  XNOR2X4 U14 ( .A(n26), .B(n23), .Y(SUM_20_) );
  NAND2X4 U15 ( .A(n1), .B(A_19_), .Y(n29) );
  INVX8 U16 ( .A(n42), .Y(SUM_16_) );
  OAI21X2 U17 ( .A0(n38), .A1(n31), .B0(n33), .Y(n36) );
  NAND2X2 U18 ( .A(B_20_), .B(A_20_), .Y(n25) );
  OR2X4 U19 ( .A(B_20_), .B(A_20_), .Y(n24) );
  AOI21X2 U20 ( .A0(n16), .A1(n32), .B0(n17), .Y(n27) );
  BUFX12 U21 ( .A(A_7_), .Y(SUM_7_) );
  BUFX12 U22 ( .A(A_8_), .Y(SUM_8_) );
  XOR2X4 U23 ( .A(n36), .B(n37), .Y(SUM_19_) );
  XOR2X4 U24 ( .A(n38), .B(n39), .Y(SUM_18_) );
  NOR2BX4 U25 ( .AN(n29), .B(n28), .Y(n37) );
  NOR2X4 U26 ( .A(n1), .B(A_19_), .Y(n28) );
  AOI21X4 U27 ( .A0(n19), .A1(n20), .B0(n18), .Y(n38) );
  NAND2X2 U28 ( .A(B_18_), .B(A_18_), .Y(n33) );
  INVX4 U29 ( .A(n31), .Y(n16) );
  INVXL U30 ( .A(n25), .Y(n15) );
  BUFX8 U31 ( .A(A_12_), .Y(SUM_12_) );
  BUFX8 U32 ( .A(A_11_), .Y(SUM_11_) );
  BUFX8 U33 ( .A(A_10_), .Y(SUM_10_) );
  BUFX8 U34 ( .A(A_9_), .Y(SUM_9_) );
  BUFX8 U35 ( .A(A_5_), .Y(SUM_5_) );
  BUFX8 U36 ( .A(A_6_), .Y(SUM_6_) );
  INVX4 U37 ( .A(n30), .Y(n19) );
  NOR2X4 U38 ( .A(A_17_), .B(B_17_), .Y(n30) );
  NAND2X4 U39 ( .A(n41), .B(n34), .Y(n42) );
  OR2X4 U40 ( .A(B_16_), .B(A_16_), .Y(n41) );
  NOR2X4 U41 ( .A(B_18_), .B(A_18_), .Y(n31) );
  NAND2X4 U42 ( .A(B_16_), .B(A_16_), .Y(n34) );
  XOR2X4 U43 ( .A(n40), .B(n20), .Y(n43) );
  NOR2X4 U44 ( .A(n18), .B(n30), .Y(n40) );
  NAND2X4 U45 ( .A(B_17_), .B(A_17_), .Y(n35) );
  XOR2X1 U46 ( .A(n21), .B(n22), .Y(SUM_21_) );
  AOI21X1 U47 ( .A0(n23), .A1(n24), .B0(n15), .Y(n22) );
  XNOR2X1 U48 ( .A(B_21_), .B(A_21_), .Y(n21) );
  NAND2X1 U49 ( .A(n25), .B(n24), .Y(n26) );
endmodule


module multi16_2_DW02_mult_0 ( A, B, PRODUCT_23_, PRODUCT_22_, PRODUCT_21_, 
        PRODUCT_20_, PRODUCT_19_, PRODUCT_18_, PRODUCT_17_, PRODUCT_16_, 
        PRODUCT_15_, PRODUCT_14_, PRODUCT_13_, PRODUCT_12_, PRODUCT_11_, 
        PRODUCT_10_, PRODUCT_9_, PRODUCT_8_, PRODUCT_7_ );
  input [16:0] A;
  input [7:0] B;
  output PRODUCT_23_, PRODUCT_22_, PRODUCT_21_, PRODUCT_20_, PRODUCT_19_,
         PRODUCT_18_, PRODUCT_17_, PRODUCT_16_, PRODUCT_15_, PRODUCT_14_,
         PRODUCT_13_, PRODUCT_12_, PRODUCT_11_, PRODUCT_10_, PRODUCT_9_,
         PRODUCT_8_, PRODUCT_7_;
  wire   ab_16__7_, ab_16__6_, ab_16__5_, ab_16__4_, ab_16__3_, ab_16__2_,
         ab_16__1_, ab_16__0_, ab_15__7_, ab_15__6_, ab_15__5_, ab_15__4_,
         ab_15__3_, ab_15__2_, ab_15__1_, ab_15__0_, ab_14__7_, ab_14__6_,
         ab_14__5_, ab_14__4_, ab_14__3_, ab_14__2_, ab_14__1_, ab_14__0_,
         ab_13__7_, ab_13__6_, ab_13__5_, ab_13__4_, ab_13__3_, ab_13__2_,
         ab_13__1_, ab_13__0_, ab_12__7_, ab_12__6_, ab_12__5_, ab_12__4_,
         ab_12__3_, ab_12__2_, ab_12__1_, ab_12__0_, ab_11__7_, ab_11__6_,
         ab_11__5_, ab_11__4_, ab_11__3_, ab_11__2_, ab_11__1_, ab_11__0_,
         ab_10__7_, ab_10__6_, ab_10__5_, ab_10__4_, ab_10__3_, ab_10__2_,
         ab_10__1_, ab_10__0_, ab_9__7_, ab_9__6_, ab_9__5_, ab_9__4_,
         ab_9__3_, ab_9__2_, ab_9__1_, ab_9__0_, ab_8__7_, ab_8__6_, ab_8__5_,
         ab_8__4_, ab_8__3_, ab_8__2_, ab_8__1_, ab_8__0_, ab_7__7_, ab_7__6_,
         ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_, ab_7__0_, ab_6__7_,
         ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_, ab_6__1_, ab_6__0_,
         ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_, ab_5__2_, ab_5__1_,
         ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_, ab_4__3_, ab_4__2_,
         ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_, ab_3__4_, ab_3__3_,
         ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_, ab_2__5_, ab_2__4_,
         ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_, ab_1__6_, ab_1__5_,
         ab_1__4_, ab_1__3_, ab_1__2_, ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_,
         ab_0__3_, ab_0__2_, CARRYB_16__6_, CARRYB_16__5_, CARRYB_16__4_,
         CARRYB_16__3_, CARRYB_16__2_, CARRYB_16__1_, CARRYB_16__0_,
         CARRYB_15__6_, CARRYB_15__5_, CARRYB_15__4_, CARRYB_15__3_,
         CARRYB_15__2_, CARRYB_15__1_, CARRYB_15__0_, CARRYB_14__6_,
         CARRYB_14__5_, CARRYB_14__4_, CARRYB_14__3_, CARRYB_14__2_,
         CARRYB_14__1_, CARRYB_14__0_, CARRYB_13__6_, CARRYB_13__5_,
         CARRYB_13__4_, CARRYB_13__3_, CARRYB_13__2_, CARRYB_13__1_,
         CARRYB_13__0_, CARRYB_12__6_, CARRYB_12__5_, CARRYB_12__4_,
         CARRYB_12__3_, CARRYB_12__2_, CARRYB_12__1_, CARRYB_12__0_,
         CARRYB_11__6_, CARRYB_11__5_, CARRYB_11__4_, CARRYB_11__3_,
         CARRYB_11__2_, CARRYB_11__1_, CARRYB_11__0_, CARRYB_10__6_,
         CARRYB_10__5_, CARRYB_10__4_, CARRYB_10__3_, CARRYB_10__2_,
         CARRYB_10__1_, CARRYB_10__0_, CARRYB_9__6_, CARRYB_9__5_,
         CARRYB_9__4_, CARRYB_9__3_, CARRYB_9__2_, CARRYB_9__1_, CARRYB_9__0_,
         CARRYB_8__6_, CARRYB_8__5_, CARRYB_8__4_, CARRYB_8__3_, CARRYB_8__2_,
         CARRYB_8__1_, CARRYB_8__0_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_,
         CARRYB_7__3_, CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_,
         CARRYB_6__5_, CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_,
         CARRYB_6__0_, CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_,
         CARRYB_5__2_, CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_,
         CARRYB_4__4_, CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_,
         CARRYB_3__6_, CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_,
         CARRYB_3__1_, CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_,
         CARRYB_2__3_, CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__6_,
         CARRYB_1__1_, CARRYB_1__0_, SUMB_16__6_, SUMB_16__5_, SUMB_16__4_,
         SUMB_16__3_, SUMB_16__2_, SUMB_16__1_, SUMB_16__0_, SUMB_15__6_,
         SUMB_15__5_, SUMB_15__4_, SUMB_15__3_, SUMB_15__2_, SUMB_15__1_,
         SUMB_14__6_, SUMB_14__5_, SUMB_14__4_, SUMB_14__3_, SUMB_14__2_,
         SUMB_14__1_, SUMB_13__6_, SUMB_13__5_, SUMB_13__4_, SUMB_13__3_,
         SUMB_13__2_, SUMB_13__1_, SUMB_12__6_, SUMB_12__5_, SUMB_12__4_,
         SUMB_12__3_, SUMB_12__2_, SUMB_12__1_, SUMB_11__6_, SUMB_11__5_,
         SUMB_11__4_, SUMB_11__3_, SUMB_11__2_, SUMB_11__1_, SUMB_10__6_,
         SUMB_10__5_, SUMB_10__4_, SUMB_10__3_, SUMB_10__2_, SUMB_10__1_,
         SUMB_9__6_, SUMB_9__5_, SUMB_9__4_, SUMB_9__3_, SUMB_9__2_,
         SUMB_9__1_, SUMB_8__6_, SUMB_8__5_, SUMB_8__4_, SUMB_8__3_,
         SUMB_8__2_, SUMB_8__1_, SUMB_7__6_, SUMB_7__5_, SUMB_7__4_,
         SUMB_7__3_, SUMB_7__2_, SUMB_7__1_, SUMB_6__6_, SUMB_6__5_,
         SUMB_6__4_, SUMB_6__3_, SUMB_6__2_, SUMB_6__1_, SUMB_5__6_,
         SUMB_5__5_, SUMB_5__4_, SUMB_5__3_, SUMB_5__2_, SUMB_5__1_,
         SUMB_4__6_, SUMB_4__5_, SUMB_4__4_, SUMB_4__3_, SUMB_4__2_,
         SUMB_4__1_, SUMB_3__6_, SUMB_3__5_, SUMB_3__4_, SUMB_3__3_,
         SUMB_3__2_, SUMB_3__1_, SUMB_2__6_, SUMB_2__5_, SUMB_2__4_,
         SUMB_2__3_, SUMB_2__2_, SUMB_2__1_, SUMB_1__6_, SUMB_1__5_,
         SUMB_1__4_, SUMB_1__3_, SUMB_1__2_, SUMB_1__1_, PROD1_7_, A1_21_,
         A1_20_, A1_19_, A1_18_, A1_17_, A1_16_, A1_15_, A1_13_, A1_12_,
         A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, A1_4_, A1_3_, A1_2_,
         A1_1_, A1_0_, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43;

  multi16_2_DW01_add_0 FS_1 ( .A_21_(A1_21_), .A_20_(A1_20_), .A_19_(A1_19_), 
        .A_18_(A1_18_), .A_17_(A1_17_), .A_16_(A1_16_), .A_15_(A1_15_), 
        .A_14_(SUMB_16__0_), .A_13_(A1_13_), .A_12_(A1_12_), .A_11_(A1_11_), 
        .A_10_(A1_10_), .A_9_(A1_9_), .A_8_(A1_8_), .A_7_(A1_7_), .A_6_(A1_6_), 
        .A_5_(PROD1_7_), .B_21_(n4), .B_20_(n21), .B_19_(n19), .B_18_(n18), 
        .B_17_(n17), .B_16_(n20), .SUM_21_(PRODUCT_23_), .SUM_20_(PRODUCT_22_), 
        .SUM_19_(PRODUCT_21_), .SUM_18_(PRODUCT_20_), .SUM_17_(PRODUCT_19_), 
        .SUM_16_(PRODUCT_18_), .SUM_15_(PRODUCT_17_), .SUM_14_(PRODUCT_16_), 
        .SUM_13_(PRODUCT_15_), .SUM_12_(PRODUCT_14_), .SUM_11_(PRODUCT_13_), 
        .SUM_10_(PRODUCT_12_), .SUM_9_(PRODUCT_11_), .SUM_8_(PRODUCT_10_), 
        .SUM_7_(PRODUCT_9_), .SUM_6_(PRODUCT_8_), .SUM_5_(PRODUCT_7_) );
  ADDFHX4 S2_9_2 ( .A(ab_9__2_), .B(CARRYB_8__2_), .CI(SUMB_8__3_), .CO(
        CARRYB_9__2_), .S(SUMB_9__2_) );
  ADDFHX4 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  ADDFHX4 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  ADDFHX4 S4_1 ( .A(ab_16__1_), .B(CARRYB_15__1_), .CI(SUMB_15__2_), .CO(
        CARRYB_16__1_), .S(SUMB_16__1_) );
  ADDFHX4 S4_2 ( .A(ab_16__2_), .B(CARRYB_15__2_), .CI(SUMB_15__3_), .CO(
        CARRYB_16__2_), .S(SUMB_16__2_) );
  ADDFHX4 S2_7_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  ADDFHX4 S2_8_1 ( .A(ab_8__1_), .B(CARRYB_7__1_), .CI(SUMB_7__2_), .CO(
        CARRYB_8__1_), .S(SUMB_8__1_) );
  ADDFHX4 S2_9_3 ( .A(ab_9__3_), .B(CARRYB_8__3_), .CI(SUMB_8__4_), .CO(
        CARRYB_9__3_), .S(SUMB_9__3_) );
  ADDFHX4 S1_7_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(PROD1_7_) );
  ADDFHX4 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  ADDFHX4 S2_10_2 ( .A(ab_10__2_), .B(CARRYB_9__2_), .CI(SUMB_9__3_), .CO(
        CARRYB_10__2_), .S(SUMB_10__2_) );
  ADDFHX4 S2_11_2 ( .A(ab_11__2_), .B(CARRYB_10__2_), .CI(SUMB_10__3_), .CO(
        CARRYB_11__2_), .S(SUMB_11__2_) );
  ADDFHX4 S1_11_0 ( .A(ab_11__0_), .B(CARRYB_10__0_), .CI(SUMB_10__1_), .CO(
        CARRYB_11__0_), .S(A1_9_) );
  ADDFHX4 S1_10_0 ( .A(ab_10__0_), .B(CARRYB_9__0_), .CI(SUMB_9__1_), .CO(
        CARRYB_10__0_), .S(A1_8_) );
  ADDFHX4 S4_3 ( .A(ab_16__3_), .B(CARRYB_15__3_), .CI(SUMB_15__4_), .CO(
        CARRYB_16__3_), .S(SUMB_16__3_) );
  ADDFHX4 S4_4 ( .A(ab_16__4_), .B(CARRYB_15__4_), .CI(SUMB_15__5_), .CO(
        CARRYB_16__4_), .S(SUMB_16__4_) );
  ADDFHX4 S2_14_1 ( .A(ab_14__1_), .B(CARRYB_13__1_), .CI(SUMB_13__2_), .CO(
        CARRYB_14__1_), .S(SUMB_14__1_) );
  ADDFHX4 S2_15_1 ( .A(ab_15__1_), .B(CARRYB_14__1_), .CI(SUMB_14__2_), .CO(
        CARRYB_15__1_), .S(SUMB_15__1_) );
  ADDFHX4 S2_7_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  ADDFHX4 S1_8_0 ( .A(ab_8__0_), .B(CARRYB_7__0_), .CI(SUMB_7__1_), .CO(
        CARRYB_8__0_), .S(A1_6_) );
  ADDFHX4 S1_9_0 ( .A(ab_9__0_), .B(CARRYB_8__0_), .CI(SUMB_8__1_), .CO(
        CARRYB_9__0_), .S(A1_7_) );
  ADDFHX4 S1_15_0 ( .A(ab_15__0_), .B(CARRYB_14__0_), .CI(SUMB_14__1_), .CO(
        CARRYB_15__0_), .S(A1_13_) );
  ADDFHX4 S4_0 ( .A(ab_16__0_), .B(CARRYB_15__0_), .CI(SUMB_15__1_), .CO(
        CARRYB_16__0_), .S(SUMB_16__0_) );
  ADDFHX4 S2_10_3 ( .A(ab_10__3_), .B(CARRYB_9__3_), .CI(SUMB_9__4_), .CO(
        CARRYB_10__3_), .S(SUMB_10__3_) );
  ADDFHX4 S2_11_3 ( .A(ab_11__3_), .B(CARRYB_10__3_), .CI(SUMB_10__4_), .CO(
        CARRYB_11__3_), .S(SUMB_11__3_) );
  ADDFHX4 S2_10_4 ( .A(ab_10__4_), .B(CARRYB_9__4_), .CI(SUMB_9__5_), .CO(
        CARRYB_10__4_), .S(SUMB_10__4_) );
  ADDFHX4 S2_11_4 ( .A(ab_11__4_), .B(CARRYB_10__4_), .CI(SUMB_10__5_), .CO(
        CARRYB_11__4_), .S(SUMB_11__4_) );
  ADDFHX1 S2_15_5 ( .A(ab_15__5_), .B(CARRYB_14__5_), .CI(SUMB_14__6_), .CO(
        CARRYB_15__5_), .S(SUMB_15__5_) );
  ADDFHX4 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  ADDFHX4 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  ADDFX2 S5_6 ( .A(ab_16__6_), .B(CARRYB_15__6_), .CI(ab_15__7_), .CO(
        CARRYB_16__6_), .S(SUMB_16__6_) );
  ADDFHX4 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  ADDFHX4 S2_7_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  ADDFHX4 S2_8_4 ( .A(ab_8__4_), .B(CARRYB_7__4_), .CI(SUMB_7__5_), .CO(
        CARRYB_8__4_), .S(SUMB_8__4_) );
  ADDFHX4 S2_9_4 ( .A(ab_9__4_), .B(CARRYB_8__4_), .CI(SUMB_8__5_), .CO(
        CARRYB_9__4_), .S(SUMB_9__4_) );
  ADDFHX4 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  ADDFHX4 S3_4_6 ( .A(ab_4__6_), .B(ab_3__7_), .CI(CARRYB_3__6_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  ADDFHX4 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  ADDFHX4 S3_10_6 ( .A(ab_10__6_), .B(CARRYB_9__6_), .CI(ab_9__7_), .CO(
        CARRYB_10__6_), .S(SUMB_10__6_) );
  ADDFHX4 S3_11_6 ( .A(ab_11__6_), .B(CARRYB_10__6_), .CI(ab_10__7_), .CO(
        CARRYB_11__6_), .S(SUMB_11__6_) );
  ADDFHX4 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  ADDFHX4 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  ADDFHX4 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  ADDFHX4 S2_13_1 ( .A(ab_13__1_), .B(CARRYB_12__1_), .CI(SUMB_12__2_), .CO(
        CARRYB_13__1_), .S(SUMB_13__1_) );
  ADDFHX4 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  ADDFHX4 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  ADDFHX4 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  ADDFHX4 S2_13_3 ( .A(ab_13__3_), .B(CARRYB_12__3_), .CI(SUMB_12__4_), .CO(
        CARRYB_13__3_), .S(SUMB_13__3_) );
  ADDFHX4 S2_14_2 ( .A(ab_14__2_), .B(CARRYB_13__2_), .CI(SUMB_13__3_), .CO(
        CARRYB_14__2_), .S(SUMB_14__2_) );
  ADDFHX4 S2_12_2 ( .A(ab_12__2_), .B(CARRYB_11__2_), .CI(SUMB_11__3_), .CO(
        CARRYB_12__2_), .S(SUMB_12__2_) );
  ADDFHX4 S2_13_2 ( .A(ab_13__2_), .B(CARRYB_12__2_), .CI(SUMB_12__3_), .CO(
        CARRYB_13__2_), .S(SUMB_13__2_) );
  ADDFHX4 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  ADDFHX4 S2_13_5 ( .A(ab_13__5_), .B(CARRYB_12__5_), .CI(SUMB_12__6_), .CO(
        CARRYB_13__5_), .S(SUMB_13__5_) );
  ADDFHX4 S2_12_5 ( .A(ab_12__5_), .B(CARRYB_11__5_), .CI(SUMB_11__6_), .CO(
        CARRYB_12__5_), .S(SUMB_12__5_) );
  ADDFHX4 S2_2_5 ( .A(ab_2__5_), .B(n8), .CI(SUMB_1__6_), .CO(CARRYB_2__5_), 
        .S(SUMB_2__5_) );
  ADDFHX4 S3_9_6 ( .A(ab_9__6_), .B(CARRYB_8__6_), .CI(ab_8__7_), .CO(
        CARRYB_9__6_), .S(SUMB_9__6_) );
  ADDFHX4 S2_11_5 ( .A(ab_11__5_), .B(CARRYB_10__5_), .CI(SUMB_10__6_), .CO(
        CARRYB_11__5_), .S(SUMB_11__5_) );
  ADDFHX4 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  ADDFHX4 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  ADDFHX4 S2_9_1 ( .A(ab_9__1_), .B(CARRYB_8__1_), .CI(SUMB_8__2_), .CO(
        CARRYB_9__1_), .S(SUMB_9__1_) );
  ADDFHX4 S2_11_1 ( .A(ab_11__1_), .B(CARRYB_10__1_), .CI(SUMB_10__2_), .CO(
        CARRYB_11__1_), .S(SUMB_11__1_) );
  ADDFHX4 S2_7_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  ADDFHX4 S2_14_3 ( .A(ab_14__3_), .B(CARRYB_13__3_), .CI(SUMB_13__4_), .CO(
        CARRYB_14__3_), .S(SUMB_14__3_) );
  ADDFHX4 S2_15_3 ( .A(ab_15__3_), .B(CARRYB_14__3_), .CI(SUMB_14__4_), .CO(
        CARRYB_15__3_), .S(SUMB_15__3_) );
  ADDFHX4 S2_12_3 ( .A(ab_12__3_), .B(CARRYB_11__3_), .CI(SUMB_11__4_), .CO(
        CARRYB_12__3_), .S(SUMB_12__3_) );
  ADDFHX4 S2_12_1 ( .A(ab_12__1_), .B(CARRYB_11__1_), .CI(SUMB_11__2_), .CO(
        CARRYB_12__1_), .S(SUMB_12__1_) );
  ADDFHX4 S2_10_5 ( .A(ab_10__5_), .B(CARRYB_9__5_), .CI(SUMB_9__6_), .CO(
        CARRYB_10__5_), .S(SUMB_10__5_) );
  ADDFHX4 S2_12_4 ( .A(ab_12__4_), .B(CARRYB_11__4_), .CI(SUMB_11__5_), .CO(
        CARRYB_12__4_), .S(SUMB_12__4_) );
  ADDFHX4 S2_13_4 ( .A(ab_13__4_), .B(CARRYB_12__4_), .CI(SUMB_12__5_), .CO(
        CARRYB_13__4_), .S(SUMB_13__4_) );
  ADDFHX2 S3_13_6 ( .A(ab_13__6_), .B(CARRYB_12__6_), .CI(ab_12__7_), .CO(
        CARRYB_13__6_), .S(SUMB_13__6_) );
  ADDFHX2 S3_14_6 ( .A(ab_14__6_), .B(CARRYB_13__6_), .CI(ab_13__7_), .CO(
        CARRYB_14__6_), .S(SUMB_14__6_) );
  ADDFHX2 S3_15_6 ( .A(ab_15__6_), .B(CARRYB_14__6_), .CI(ab_14__7_), .CO(
        CARRYB_15__6_), .S(SUMB_15__6_) );
  ADDFHX4 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  ADDFHX4 S1_13_0 ( .A(ab_13__0_), .B(CARRYB_12__0_), .CI(SUMB_12__1_), .CO(
        CARRYB_13__0_), .S(A1_11_) );
  ADDFHX4 S1_14_0 ( .A(ab_14__0_), .B(CARRYB_13__0_), .CI(SUMB_13__1_), .CO(
        CARRYB_14__0_), .S(A1_12_) );
  ADDFHX4 S2_15_2 ( .A(ab_15__2_), .B(CARRYB_14__2_), .CI(SUMB_14__3_), .CO(
        CARRYB_15__2_), .S(SUMB_15__2_) );
  ADDFHX4 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  ADDFHX4 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  ADDFHX4 S2_9_5 ( .A(ab_9__5_), .B(CARRYB_8__5_), .CI(SUMB_8__6_), .CO(
        CARRYB_9__5_), .S(SUMB_9__5_) );
  ADDFHX4 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  ADDFHX4 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  ADDFHX4 S3_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(ab_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  ADDFHX4 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  ADDFHX4 S1_12_0 ( .A(ab_12__0_), .B(CARRYB_11__0_), .CI(SUMB_11__1_), .CO(
        CARRYB_12__0_), .S(A1_10_) );
  ADDFHX4 S2_2_4 ( .A(ab_2__4_), .B(n7), .CI(SUMB_1__5_), .CO(CARRYB_2__4_), 
        .S(SUMB_2__4_) );
  ADDFHX4 S2_8_3 ( .A(ab_8__3_), .B(CARRYB_7__3_), .CI(SUMB_7__4_), .CO(
        CARRYB_8__3_), .S(SUMB_8__3_) );
  ADDFHX4 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  ADDFHX4 S2_10_1 ( .A(ab_10__1_), .B(CARRYB_9__1_), .CI(SUMB_9__2_), .CO(
        CARRYB_10__1_), .S(SUMB_10__1_) );
  ADDFHX4 S2_14_4 ( .A(ab_14__4_), .B(CARRYB_13__4_), .CI(SUMB_13__5_), .CO(
        CARRYB_14__4_), .S(SUMB_14__4_) );
  ADDFHX4 S2_2_2 ( .A(ab_2__2_), .B(n5), .CI(SUMB_1__3_), .CO(CARRYB_2__2_), 
        .S(SUMB_2__2_) );
  ADDFHX4 S2_8_2 ( .A(ab_8__2_), .B(CARRYB_7__2_), .CI(SUMB_7__3_), .CO(
        CARRYB_8__2_), .S(SUMB_8__2_) );
  ADDFHX4 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  ADDFHX4 S3_8_6 ( .A(ab_8__6_), .B(CARRYB_7__6_), .CI(ab_7__7_), .CO(
        CARRYB_8__6_), .S(SUMB_8__6_) );
  ADDFHX4 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  ADDFHX4 S2_8_5 ( .A(ab_8__5_), .B(CARRYB_7__5_), .CI(SUMB_7__6_), .CO(
        CARRYB_8__5_), .S(SUMB_8__5_) );
  ADDFHX4 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  ADDFHX4 S3_12_6 ( .A(ab_12__6_), .B(CARRYB_11__6_), .CI(ab_11__7_), .CO(
        CARRYB_12__6_), .S(SUMB_12__6_) );
  ADDFHX4 S2_2_3 ( .A(ab_2__3_), .B(n6), .CI(SUMB_1__4_), .CO(CARRYB_2__3_), 
        .S(SUMB_2__3_) );
  ADDFHX2 S2_15_4 ( .A(ab_15__4_), .B(CARRYB_14__4_), .CI(SUMB_14__5_), .CO(
        CARRYB_15__4_), .S(SUMB_15__4_) );
  ADDFHX4 S3_7_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(
        CARRYB_7__6_), .S(SUMB_7__6_) );
  ADDFHX2 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  ADDFHX4 S4_5 ( .A(ab_16__5_), .B(CARRYB_15__5_), .CI(SUMB_15__6_), .CO(
        CARRYB_16__5_), .S(SUMB_16__5_) );
  ADDFHX4 S2_14_5 ( .A(ab_14__5_), .B(CARRYB_13__5_), .CI(SUMB_13__6_), .CO(
        CARRYB_14__5_), .S(SUMB_14__5_) );
  XOR2X2 U2 ( .A(ab_1__2_), .B(ab_0__3_), .Y(SUMB_1__2_) );
  NAND2X2 U3 ( .A(ab_0__2_), .B(n43), .Y(n23) );
  NOR2BX2 U4 ( .AN(A[1]), .B(n42), .Y(ab_1__7_) );
  NOR2BX4 U5 ( .AN(A[3]), .B(n38), .Y(ab_3__3_) );
  NOR2BX4 U6 ( .AN(A[3]), .B(n30), .Y(ab_3__1_) );
  NOR2BX4 U7 ( .AN(A[3]), .B(n39), .Y(ab_3__2_) );
  NOR2BX4 U8 ( .AN(A[3]), .B(n37), .Y(ab_3__4_) );
  NOR2BX4 U9 ( .AN(A[2]), .B(n24), .Y(ab_2__5_) );
  NOR2BX1 U10 ( .AN(A[6]), .B(n26), .Y(ab_6__4_) );
  NOR2BXL U11 ( .AN(A[12]), .B(n28), .Y(ab_12__2_) );
  NOR2BX1 U12 ( .AN(A[7]), .B(n39), .Y(ab_7__2_) );
  NOR2BX2 U13 ( .AN(A[7]), .B(n37), .Y(ab_7__4_) );
  NOR2BXL U14 ( .AN(A[11]), .B(n28), .Y(ab_11__2_) );
  NOR2BX1 U15 ( .AN(A[6]), .B(n39), .Y(ab_6__2_) );
  NOR2BX1 U16 ( .AN(A[9]), .B(n28), .Y(ab_9__2_) );
  NOR2BX1 U17 ( .AN(A[13]), .B(n30), .Y(ab_13__1_) );
  NOR2BX2 U18 ( .AN(A[7]), .B(n30), .Y(ab_7__1_) );
  NOR2BX1 U19 ( .AN(A[9]), .B(n25), .Y(ab_9__5_) );
  NOR2BX1 U20 ( .AN(A[9]), .B(n27), .Y(ab_9__3_) );
  NOR2BX2 U21 ( .AN(A[10]), .B(n30), .Y(ab_10__1_) );
  NOR2BX1 U22 ( .AN(A[14]), .B(n31), .Y(ab_14__0_) );
  NOR2BX2 U23 ( .AN(A[2]), .B(n31), .Y(ab_2__0_) );
  NOR2BX1 U24 ( .AN(A[9]), .B(n31), .Y(ab_9__0_) );
  NOR2BX1 U25 ( .AN(A[9]), .B(n26), .Y(ab_9__4_) );
  NOR2BX1 U26 ( .AN(A[7]), .B(n38), .Y(ab_7__3_) );
  NOR2BX1 U27 ( .AN(A[14]), .B(n28), .Y(ab_14__2_) );
  NOR2BX2 U28 ( .AN(A[11]), .B(n30), .Y(ab_11__1_) );
  NOR2BX1 U29 ( .AN(A[5]), .B(n28), .Y(ab_5__2_) );
  CLKBUFX8 U30 ( .A(n41), .Y(n31) );
  NOR2BX2 U31 ( .AN(A[5]), .B(n30), .Y(ab_5__1_) );
  BUFX12 U32 ( .A(n35), .Y(n29) );
  AND2X2 U34 ( .A(CARRYB_16__5_), .B(SUMB_16__6_), .Y(n4) );
  AND2X4 U35 ( .A(ab_0__3_), .B(ab_1__2_), .Y(n5) );
  AND2X4 U36 ( .A(ab_0__4_), .B(ab_1__3_), .Y(n6) );
  AND2X4 U37 ( .A(ab_0__5_), .B(ab_1__4_), .Y(n7) );
  AND2X4 U38 ( .A(ab_0__6_), .B(ab_1__5_), .Y(n8) );
  INVX4 U39 ( .A(B[2]), .Y(n39) );
  CLKBUFX2 U40 ( .A(n39), .Y(n28) );
  CLKINVX8 U41 ( .A(B[4]), .Y(n37) );
  CLKBUFX2 U42 ( .A(n37), .Y(n26) );
  INVX4 U43 ( .A(B[3]), .Y(n38) );
  BUFX3 U44 ( .A(n38), .Y(n27) );
  INVX8 U45 ( .A(n34), .Y(n43) );
  NOR2X2 U46 ( .A(n34), .B(n33), .Y(CARRYB_1__0_) );
  XOR2X4 U47 ( .A(ab_1__6_), .B(ab_0__7_), .Y(SUMB_1__6_) );
  AND2X4 U48 ( .A(B[7]), .B(A[0]), .Y(ab_0__7_) );
  XOR2X4 U49 ( .A(ab_6__6_), .B(ab_5__7_), .Y(n9) );
  XOR2X4 U50 ( .A(CARRYB_5__6_), .B(n9), .Y(SUMB_6__6_) );
  NAND2X1 U51 ( .A(ab_6__6_), .B(CARRYB_5__6_), .Y(n10) );
  NAND2X1 U52 ( .A(ab_5__7_), .B(CARRYB_5__6_), .Y(n11) );
  NAND2X2 U53 ( .A(ab_5__7_), .B(ab_6__6_), .Y(n12) );
  NAND3X4 U54 ( .A(n12), .B(n10), .C(n11), .Y(CARRYB_6__6_) );
  NOR2BX4 U55 ( .AN(A[6]), .B(n29), .Y(ab_6__6_) );
  NOR2BX2 U56 ( .AN(A[5]), .B(n42), .Y(ab_5__7_) );
  XOR2X4 U57 ( .A(CARRYB_16__4_), .B(SUMB_16__5_), .Y(A1_19_) );
  AND2X4 U58 ( .A(B[6]), .B(A[0]), .Y(ab_0__6_) );
  CLKINVX3 U59 ( .A(B[6]), .Y(n35) );
  NOR2BX4 U60 ( .AN(A[2]), .B(n37), .Y(ab_2__4_) );
  NOR2BX4 U61 ( .AN(A[2]), .B(n38), .Y(ab_2__3_) );
  NOR2BX4 U62 ( .AN(A[2]), .B(n39), .Y(ab_2__2_) );
  XOR2X2 U63 ( .A(ab_1__3_), .B(ab_0__4_), .Y(SUMB_1__3_) );
  NOR2BX4 U64 ( .AN(A[2]), .B(n30), .Y(ab_2__1_) );
  XOR2X4 U65 ( .A(ab_1__5_), .B(ab_0__6_), .Y(SUMB_1__5_) );
  NOR2BX2 U66 ( .AN(A[4]), .B(n29), .Y(ab_4__6_) );
  AND2X2 U67 ( .A(A[2]), .B(B[6]), .Y(ab_2__6_) );
  NOR2BX1 U68 ( .AN(A[4]), .B(n37), .Y(ab_4__4_) );
  NAND2X4 U69 ( .A(ab_0__7_), .B(ab_1__6_), .Y(n22) );
  NAND2X4 U70 ( .A(ab_7__5_), .B(CARRYB_6__5_), .Y(n15) );
  NAND2X4 U71 ( .A(SUMB_6__6_), .B(CARRYB_6__5_), .Y(n14) );
  NAND2X4 U72 ( .A(A[1]), .B(B[1]), .Y(n34) );
  NOR2BX1 U73 ( .AN(A[6]), .B(n27), .Y(ab_6__3_) );
  NOR2BXL U74 ( .AN(A[16]), .B(n29), .Y(ab_16__6_) );
  NOR2BXL U75 ( .AN(A[15]), .B(n29), .Y(ab_15__6_) );
  NOR2BXL U76 ( .AN(A[14]), .B(n29), .Y(ab_14__6_) );
  NOR2BXL U77 ( .AN(A[13]), .B(n29), .Y(ab_13__6_) );
  NOR2BXL U78 ( .AN(A[12]), .B(n29), .Y(ab_12__6_) );
  NOR2BXL U79 ( .AN(A[11]), .B(n29), .Y(ab_11__6_) );
  NOR2BXL U80 ( .AN(A[9]), .B(n29), .Y(ab_9__6_) );
  NOR2BX2 U81 ( .AN(A[3]), .B(n29), .Y(ab_3__6_) );
  XOR2X4 U82 ( .A(ab_1__4_), .B(ab_0__5_), .Y(SUMB_1__4_) );
  NOR2BXL U83 ( .AN(A[10]), .B(n29), .Y(ab_10__6_) );
  XOR2X4 U84 ( .A(CARRYB_6__5_), .B(n13), .Y(SUMB_7__5_) );
  XOR2X2 U85 ( .A(n43), .B(ab_0__2_), .Y(SUMB_1__1_) );
  AND2X4 U86 ( .A(B[6]), .B(A[1]), .Y(ab_1__6_) );
  BUFX20 U87 ( .A(n36), .Y(n24) );
  NOR2BX2 U88 ( .AN(B[2]), .B(n32), .Y(ab_0__2_) );
  AND2X4 U89 ( .A(CARRYB_16__1_), .B(SUMB_16__2_), .Y(n17) );
  INVX8 U90 ( .A(B[5]), .Y(n36) );
  CLKINVX8 U91 ( .A(B[1]), .Y(n40) );
  NOR2BX2 U92 ( .AN(A[3]), .B(n24), .Y(ab_3__5_) );
  NOR2BX2 U93 ( .AN(A[3]), .B(n31), .Y(ab_3__0_) );
  INVX8 U94 ( .A(A[0]), .Y(n32) );
  INVX4 U95 ( .A(n22), .Y(CARRYB_1__6_) );
  XOR2X4 U96 ( .A(SUMB_6__6_), .B(ab_7__5_), .Y(n13) );
  NOR2BX4 U97 ( .AN(A[1]), .B(n39), .Y(ab_1__2_) );
  INVX4 U98 ( .A(n23), .Y(CARRYB_1__1_) );
  NOR2BX2 U99 ( .AN(B[4]), .B(n32), .Y(ab_0__4_) );
  NAND2X1 U100 ( .A(ab_7__5_), .B(SUMB_6__6_), .Y(n16) );
  NOR2BX4 U101 ( .AN(A[7]), .B(n24), .Y(ab_7__5_) );
  INVX20 U102 ( .A(B[7]), .Y(n42) );
  NOR2BX4 U103 ( .AN(B[5]), .B(n32), .Y(ab_0__5_) );
  AND2X4 U104 ( .A(CARRYB_16__0_), .B(SUMB_16__1_), .Y(n20) );
  NOR2BX4 U105 ( .AN(A[1]), .B(n38), .Y(ab_1__3_) );
  NOR2BX4 U106 ( .AN(A[1]), .B(n37), .Y(ab_1__4_) );
  NOR2BX4 U107 ( .AN(A[1]), .B(n24), .Y(ab_1__5_) );
  NAND3X4 U108 ( .A(n16), .B(n14), .C(n15), .Y(CARRYB_7__5_) );
  NOR2BX1 U109 ( .AN(A[13]), .B(n31), .Y(ab_13__0_) );
  NOR2BX1 U110 ( .AN(A[13]), .B(n28), .Y(ab_13__2_) );
  NOR2BX1 U111 ( .AN(A[10]), .B(n31), .Y(ab_10__0_) );
  NOR2BXL U112 ( .AN(A[14]), .B(n30), .Y(ab_14__1_) );
  NOR2BX1 U113 ( .AN(A[15]), .B(n31), .Y(ab_15__0_) );
  NOR2BX2 U114 ( .AN(B[3]), .B(n32), .Y(ab_0__3_) );
  NOR2BX1 U115 ( .AN(A[7]), .B(n31), .Y(ab_7__0_) );
  BUFX12 U116 ( .A(n40), .Y(n30) );
  NOR2BX2 U117 ( .AN(A[12]), .B(n30), .Y(ab_12__1_) );
  NOR2BX1 U118 ( .AN(A[4]), .B(n39), .Y(ab_4__2_) );
  NOR2BX1 U119 ( .AN(A[5]), .B(n37), .Y(ab_5__4_) );
  NOR2BX1 U120 ( .AN(A[9]), .B(n30), .Y(ab_9__1_) );
  NOR2BX1 U121 ( .AN(A[6]), .B(n31), .Y(ab_6__0_) );
  CLKBUFXL U122 ( .A(n36), .Y(n25) );
  NOR2BX1 U123 ( .AN(A[5]), .B(n31), .Y(ab_5__0_) );
  NOR2BX1 U124 ( .AN(A[4]), .B(n31), .Y(ab_4__0_) );
  AND2X1 U125 ( .A(CARRYB_16__3_), .B(SUMB_16__4_), .Y(n19) );
  NOR2BX1 U126 ( .AN(A[4]), .B(n24), .Y(ab_4__5_) );
  NOR2BX1 U127 ( .AN(A[4]), .B(n38), .Y(ab_4__3_) );
  NOR2BX1 U128 ( .AN(A[5]), .B(n38), .Y(ab_5__3_) );
  NOR2BX1 U129 ( .AN(A[10]), .B(n25), .Y(ab_10__5_) );
  NOR2BX1 U130 ( .AN(A[13]), .B(n27), .Y(ab_13__3_) );
  NOR2BX1 U131 ( .AN(A[12]), .B(n26), .Y(ab_12__4_) );
  NOR2BX1 U132 ( .AN(A[14]), .B(n27), .Y(ab_14__3_) );
  NOR2BX1 U133 ( .AN(A[12]), .B(n27), .Y(ab_12__3_) );
  NOR2BX1 U134 ( .AN(A[13]), .B(n26), .Y(ab_13__4_) );
  NOR2BX1 U135 ( .AN(A[6]), .B(n30), .Y(ab_6__1_) );
  NOR2BX1 U136 ( .AN(A[11]), .B(n26), .Y(ab_11__4_) );
  NOR2BX1 U137 ( .AN(A[10]), .B(n27), .Y(ab_10__3_) );
  NOR2BX1 U138 ( .AN(A[11]), .B(n27), .Y(ab_11__3_) );
  NOR2BX1 U139 ( .AN(A[10]), .B(n28), .Y(ab_10__2_) );
  NOR2BX1 U140 ( .AN(A[16]), .B(n25), .Y(ab_16__5_) );
  NOR2BX1 U141 ( .AN(A[8]), .B(n29), .Y(ab_8__6_) );
  NOR2BX1 U142 ( .AN(A[16]), .B(n28), .Y(ab_16__2_) );
  NOR2BX1 U143 ( .AN(A[15]), .B(n27), .Y(ab_15__3_) );
  NOR2BX1 U144 ( .AN(A[15]), .B(n28), .Y(ab_15__2_) );
  NOR2BX1 U145 ( .AN(A[15]), .B(n26), .Y(ab_15__4_) );
  NOR2BX1 U146 ( .AN(A[11]), .B(n25), .Y(ab_11__5_) );
  NOR2BXL U147 ( .AN(A[8]), .B(n27), .Y(ab_8__3_) );
  NOR2BX1 U148 ( .AN(A[4]), .B(n30), .Y(ab_4__1_) );
  NOR2BXL U149 ( .AN(A[8]), .B(n39), .Y(ab_8__2_) );
  NOR2BX1 U150 ( .AN(A[5]), .B(n24), .Y(ab_5__5_) );
  NOR2BX2 U151 ( .AN(A[12]), .B(n31), .Y(ab_12__0_) );
  NOR2BXL U152 ( .AN(A[8]), .B(n37), .Y(ab_8__4_) );
  AND2X2 U153 ( .A(CARRYB_16__2_), .B(SUMB_16__3_), .Y(n18) );
  NOR2BX1 U154 ( .AN(A[14]), .B(n26), .Y(ab_14__4_) );
  NOR2BX1 U155 ( .AN(A[14]), .B(n25), .Y(ab_14__5_) );
  XOR2X1 U156 ( .A(CARRYB_16__5_), .B(SUMB_16__6_), .Y(A1_20_) );
  NOR2BX1 U157 ( .AN(A[10]), .B(n26), .Y(ab_10__4_) );
  NOR2BXL U158 ( .AN(A[8]), .B(n31), .Y(ab_8__0_) );
  NOR2BX2 U159 ( .AN(A[11]), .B(n31), .Y(ab_11__0_) );
  NOR2BXL U160 ( .AN(A[8]), .B(n30), .Y(ab_8__1_) );
  NOR2BXL U161 ( .AN(A[8]), .B(n24), .Y(ab_8__5_) );
  AND2X2 U162 ( .A(CARRYB_16__4_), .B(SUMB_16__5_), .Y(n21) );
  NOR2BXL U163 ( .AN(A[6]), .B(n24), .Y(ab_6__5_) );
  NOR2BX1 U164 ( .AN(A[12]), .B(n25), .Y(ab_12__5_) );
  NOR2BXL U165 ( .AN(A[13]), .B(n25), .Y(ab_13__5_) );
  XOR2X1 U166 ( .A(CARRYB_16__6_), .B(ab_16__7_), .Y(A1_21_) );
  NOR2BX1 U167 ( .AN(A[15]), .B(n42), .Y(ab_15__7_) );
  NOR2BX1 U168 ( .AN(A[6]), .B(n42), .Y(ab_6__7_) );
  NOR2BX1 U169 ( .AN(A[7]), .B(n29), .Y(ab_7__6_) );
  NOR2BXL U170 ( .AN(A[15]), .B(n25), .Y(ab_15__5_) );
  NOR2BX1 U171 ( .AN(A[13]), .B(n42), .Y(ab_13__7_) );
  NOR2BX1 U172 ( .AN(A[9]), .B(n42), .Y(ab_9__7_) );
  NOR2BXL U173 ( .AN(A[16]), .B(n30), .Y(ab_16__1_) );
  NOR2BX1 U174 ( .AN(A[16]), .B(n27), .Y(ab_16__3_) );
  NOR2BX1 U175 ( .AN(A[16]), .B(n26), .Y(ab_16__4_) );
  NOR2BXL U176 ( .AN(A[16]), .B(n31), .Y(ab_16__0_) );
  NOR2BX1 U177 ( .AN(A[10]), .B(n42), .Y(ab_10__7_) );
  NOR2BX1 U178 ( .AN(A[11]), .B(n42), .Y(ab_11__7_) );
  NOR2BX1 U179 ( .AN(A[12]), .B(n42), .Y(ab_12__7_) );
  NOR2BX1 U180 ( .AN(A[14]), .B(n42), .Y(ab_14__7_) );
  NOR2BXL U181 ( .AN(A[15]), .B(n30), .Y(ab_15__1_) );
  NOR2BX1 U182 ( .AN(A[8]), .B(n42), .Y(ab_8__7_) );
  NOR2BX1 U183 ( .AN(A[4]), .B(n42), .Y(ab_4__7_) );
  NOR2BX2 U184 ( .AN(A[5]), .B(n29), .Y(ab_5__6_) );
  NOR2BX1 U185 ( .AN(A[2]), .B(n42), .Y(ab_2__7_) );
  NOR2BX1 U186 ( .AN(A[7]), .B(n42), .Y(ab_7__7_) );
  NOR2BX1 U187 ( .AN(A[3]), .B(n42), .Y(ab_3__7_) );
  INVXL U188 ( .A(B[0]), .Y(n41) );
  NOR2BX1 U189 ( .AN(A[16]), .B(n42), .Y(ab_16__7_) );
  NAND2XL U190 ( .A(A[0]), .B(B[0]), .Y(n33) );
  XOR2X4 U191 ( .A(SUMB_16__2_), .B(CARRYB_16__1_), .Y(A1_16_) );
  XOR2X4 U192 ( .A(CARRYB_16__3_), .B(SUMB_16__4_), .Y(A1_18_) );
  XOR2X4 U193 ( .A(CARRYB_16__0_), .B(SUMB_16__1_), .Y(A1_15_) );
  XOR2X4 U194 ( .A(CARRYB_16__2_), .B(SUMB_16__3_), .Y(A1_17_) );
endmodule


module multi16_2 ( in_17bit, in_8bit, out );
  input [16:0] in_17bit;
  input [7:0] in_8bit;
  output [16:0] out;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121;
  wire   [16:1] in_17bit_b;
  wire   [7:1] in_8bit_b;
  wire   [23:8] mul;

  multi16_2_DW02_mult_0 mult_55 ( .A({in_17bit_b[16:2], n10, n17}), .B({
        in_8bit_b, n15}), .PRODUCT_23_(mul[23]), .PRODUCT_22_(mul[22]), 
        .PRODUCT_21_(mul[21]), .PRODUCT_20_(mul[20]), .PRODUCT_19_(mul[19]), 
        .PRODUCT_18_(mul[18]), .PRODUCT_17_(mul[17]), .PRODUCT_16_(mul[16]), 
        .PRODUCT_15_(mul[15]), .PRODUCT_14_(mul[14]), .PRODUCT_13_(mul[13]), 
        .PRODUCT_12_(mul[12]), .PRODUCT_11_(mul[11]), .PRODUCT_10_(mul[10]), 
        .PRODUCT_9_(mul[9]), .PRODUCT_8_(mul[8]), .PRODUCT_7_(out[0]) );
  INVX16 U2 ( .A(in_17bit[0]), .Y(n16) );
  INVX3 U3 ( .A(mul[20]), .Y(n1) );
  INVX4 U4 ( .A(n1), .Y(n2) );
  AND2X2 U5 ( .A(n41), .B(n61), .Y(n36) );
  NAND2XL U6 ( .A(n41), .B(n80), .Y(n79) );
  NAND3X2 U7 ( .A(in_17bit[1]), .B(n41), .C(in_17bit[0]), .Y(n40) );
  XOR2X2 U8 ( .A(n81), .B(n79), .Y(in_17bit_b[11]) );
  NAND2BX4 U9 ( .AN(mul[19]), .B(n114), .Y(n7) );
  NAND2BX2 U10 ( .AN(mul[19]), .B(n114), .Y(n117) );
  NOR2X2 U11 ( .A(n2), .B(n117), .Y(n3) );
  BUFX16 U12 ( .A(in_17bit[16]), .Y(n41) );
  CLKINVX8 U13 ( .A(n55), .Y(n21) );
  BUFX4 U14 ( .A(n63), .Y(n4) );
  XNOR2X2 U15 ( .A(mul[11]), .B(n95), .Y(out[4]) );
  NAND2X2 U16 ( .A(n68), .B(n67), .Y(n70) );
  NAND2X2 U17 ( .A(n32), .B(n89), .Y(n91) );
  CLKINVX3 U18 ( .A(in_8bit[3]), .Y(n53) );
  BUFX20 U19 ( .A(in_17bit_b[1]), .Y(n10) );
  NOR2BX4 U20 ( .AN(n41), .B(n13), .Y(n60) );
  INVX12 U21 ( .A(n41), .Y(n5) );
  NAND2XL U22 ( .A(n41), .B(n64), .Y(n63) );
  XNOR2X4 U23 ( .A(mul[16]), .B(n104), .Y(out[9]) );
  INVX8 U24 ( .A(in_8bit[0]), .Y(n50) );
  NOR2XL U25 ( .A(mul[21]), .B(n2), .Y(n119) );
  AND2X2 U26 ( .A(in_8bit[0]), .B(n43), .Y(n29) );
  OAI21X4 U27 ( .A0(n46), .A1(n14), .B0(n43), .Y(n51) );
  OR2X4 U28 ( .A(n38), .B(n5), .Y(n28) );
  OR2X2 U29 ( .A(n68), .B(n5), .Y(n30) );
  NOR2X1 U30 ( .A(n31), .B(n5), .Y(n25) );
  OR2X4 U31 ( .A(in_17bit[0]), .B(in_17bit[1]), .Y(n59) );
  INVXL U32 ( .A(n5), .Y(n6) );
  AOI21X2 U33 ( .A0(n120), .A1(n119), .B0(n118), .Y(n121) );
  NAND2X4 U34 ( .A(n38), .B(n62), .Y(n64) );
  NAND2XL U35 ( .A(n6), .B(n85), .Y(n84) );
  NAND2XL U36 ( .A(n41), .B(n74), .Y(n73) );
  NAND2XL U37 ( .A(n6), .B(n70), .Y(n69) );
  NOR2X1 U38 ( .A(mul[22]), .B(n117), .Y(n120) );
  XOR2X4 U39 ( .A(n113), .B(mul[21]), .Y(out[14]) );
  AOI2BB1X4 U40 ( .A0N(mul[20]), .A1N(n7), .B0(n118), .Y(n113) );
  NOR2X4 U41 ( .A(n114), .B(n8), .Y(n110) );
  CLKINVX20 U42 ( .A(n115), .Y(n8) );
  NAND3BX4 U43 ( .AN(n46), .B(n21), .C(n56), .Y(n9) );
  NAND2X4 U44 ( .A(n58), .B(n12), .Y(n11) );
  XOR2X4 U45 ( .A(mul[8]), .B(n23), .Y(out[1]) );
  NOR2X4 U46 ( .A(in_17bit[0]), .B(in_17bit[1]), .Y(n13) );
  NAND2BX2 U47 ( .AN(n64), .B(n65), .Y(n66) );
  CLKINVX8 U48 ( .A(in_17bit[5]), .Y(n65) );
  OAI21X2 U49 ( .A0(n46), .A1(in_8bit[0]), .B0(n43), .Y(n49) );
  XOR2X4 U50 ( .A(n11), .B(n42), .Y(in_8bit_b[5]) );
  XNOR2X1 U51 ( .A(n6), .B(n43), .Y(n118) );
  CLKBUFX3 U52 ( .A(n52), .Y(n14) );
  INVX8 U53 ( .A(in_8bit[1]), .Y(n47) );
  INVX8 U54 ( .A(in_8bit[7]), .Y(n45) );
  CLKINVX8 U55 ( .A(in_8bit[7]), .Y(n44) );
  CLKINVX20 U56 ( .A(n44), .Y(n12) );
  NAND2X4 U57 ( .A(n22), .B(n43), .Y(n54) );
  INVX2 U58 ( .A(n46), .Y(n20) );
  INVX8 U59 ( .A(n47), .Y(n46) );
  NOR4BX2 U60 ( .AN(n43), .B(n9), .C(in_8bit[6]), .D(in_8bit[5]), .Y(
        in_8bit_b[7]) );
  CLKINVX3 U61 ( .A(in_8bit[5]), .Y(n42) );
  CLKINVX8 U62 ( .A(n112), .Y(n114) );
  INVX4 U63 ( .A(mul[21]), .Y(n18) );
  AOI2BB1X4 U64 ( .A0N(n9), .A1N(in_8bit[5]), .B0(n44), .Y(n57) );
  XNOR2X4 U65 ( .A(n47), .B(n29), .Y(in_8bit_b[1]) );
  INVX8 U66 ( .A(in_8bit[4]), .Y(n56) );
  INVXL U67 ( .A(n50), .Y(n15) );
  OAI21X4 U68 ( .A0(n112), .A1(mul[19]), .B0(n115), .Y(n111) );
  OR2X4 U69 ( .A(mul[12]), .B(n97), .Y(n99) );
  XNOR2X4 U70 ( .A(mul[20]), .B(n111), .Y(out[13]) );
  CLKINVX4 U71 ( .A(n16), .Y(n17) );
  XOR2X2 U72 ( .A(mul[23]), .B(n121), .Y(out[16]) );
  NOR2X4 U73 ( .A(in_17bit[3]), .B(n61), .Y(n38) );
  NAND2BX4 U74 ( .AN(in_17bit[2]), .B(n13), .Y(n61) );
  OR2X4 U75 ( .A(n41), .B(in_17bit[1]), .Y(n37) );
  NOR2X1 U76 ( .A(n70), .B(in_17bit[7]), .Y(n31) );
  XOR2X2 U77 ( .A(n75), .B(n73), .Y(in_17bit_b[9]) );
  OR2X4 U78 ( .A(mul[8]), .B(out[0]), .Y(n93) );
  OR2X4 U79 ( .A(mul[9]), .B(n93), .Y(n94) );
  XNOR2X4 U80 ( .A(mul[17]), .B(n24), .Y(out[10]) );
  XOR2X4 U81 ( .A(n54), .B(n56), .Y(in_8bit_b[4]) );
  OR2X4 U82 ( .A(mul[11]), .B(n96), .Y(n97) );
  NAND2X4 U83 ( .A(n18), .B(n3), .Y(n19) );
  NAND2X4 U84 ( .A(n19), .B(n115), .Y(n116) );
  NAND2X2 U85 ( .A(n20), .B(n21), .Y(n22) );
  INVX8 U86 ( .A(n45), .Y(n43) );
  XOR2X4 U87 ( .A(in_17bit[3]), .B(n36), .Y(in_17bit_b[3]) );
  NAND2X2 U88 ( .A(n31), .B(n72), .Y(n74) );
  INVXL U89 ( .A(in_17bit[13]), .Y(n86) );
  INVXL U90 ( .A(in_17bit[14]), .Y(n89) );
  OR2X4 U91 ( .A(mul[16]), .B(n105), .Y(n106) );
  NAND2X4 U92 ( .A(n105), .B(n115), .Y(n104) );
  INVXL U93 ( .A(in_17bit[9]), .Y(n75) );
  NAND2X4 U94 ( .A(n106), .B(n115), .Y(n24) );
  NAND2X4 U95 ( .A(n33), .B(n83), .Y(n85) );
  INVXL U96 ( .A(in_17bit[7]), .Y(n71) );
  INVXL U97 ( .A(in_17bit[11]), .Y(n81) );
  OR2X4 U98 ( .A(mul[18]), .B(n109), .Y(n112) );
  OR2X4 U99 ( .A(mul[14]), .B(n101), .Y(n103) );
  OR2X4 U100 ( .A(mul[13]), .B(n99), .Y(n101) );
  OR2XL U101 ( .A(mul[10]), .B(n94), .Y(n96) );
  AND2X4 U102 ( .A(out[0]), .B(n115), .Y(n23) );
  XOR2X4 U103 ( .A(mul[12]), .B(n26), .Y(out[5]) );
  AND2X4 U104 ( .A(n97), .B(n115), .Y(n26) );
  NAND2X4 U105 ( .A(n93), .B(n115), .Y(n92) );
  INVX4 U106 ( .A(n118), .Y(n115) );
  XNOR2X2 U107 ( .A(n25), .B(n72), .Y(in_17bit_b[8]) );
  AND2X4 U108 ( .A(n76), .B(n75), .Y(n35) );
  NOR2X4 U109 ( .A(n80), .B(n34), .Y(n33) );
  INVX1 U110 ( .A(n81), .Y(n34) );
  AND2X4 U111 ( .A(n87), .B(n86), .Y(n32) );
  XNOR2X4 U112 ( .A(n116), .B(mul[22]), .Y(out[15]) );
  OR2X4 U113 ( .A(mul[15]), .B(n103), .Y(n105) );
  NAND2X1 U114 ( .A(n96), .B(n115), .Y(n95) );
  XOR2X4 U115 ( .A(mul[10]), .B(n27), .Y(out[3]) );
  AND2X4 U116 ( .A(n94), .B(n115), .Y(n27) );
  XOR2X4 U117 ( .A(n110), .B(mul[19]), .Y(out[12]) );
  NAND2BX4 U118 ( .AN(n52), .B(n53), .Y(n55) );
  XOR2X4 U119 ( .A(n28), .B(n62), .Y(in_17bit_b[4]) );
  INVXL U120 ( .A(in_8bit[2]), .Y(n48) );
  XOR2X4 U121 ( .A(n30), .B(n67), .Y(in_17bit_b[6]) );
  NOR2XL U122 ( .A(n33), .B(n5), .Y(n82) );
  XOR2X1 U123 ( .A(n86), .B(n84), .Y(in_17bit_b[13]) );
  NOR2XL U124 ( .A(n32), .B(n5), .Y(n88) );
  NOR2XL U125 ( .A(n35), .B(n5), .Y(n77) );
  XNOR2X2 U126 ( .A(n90), .B(n39), .Y(in_17bit_b[15]) );
  AND2X1 U127 ( .A(n41), .B(n91), .Y(n39) );
  AND3X4 U128 ( .A(n37), .B(n59), .C(n40), .Y(in_17bit_b[1]) );
  XOR2X4 U129 ( .A(n49), .B(n48), .Y(in_8bit_b[2]) );
  NAND2BX4 U130 ( .AN(in_8bit[2]), .B(n50), .Y(n52) );
  XOR2X4 U131 ( .A(n51), .B(n53), .Y(in_8bit_b[3]) );
  NAND3BX4 U132 ( .AN(n46), .B(n21), .C(n56), .Y(n58) );
  XOR2X4 U133 ( .A(n57), .B(in_8bit[6]), .Y(in_8bit_b[6]) );
  XOR2X4 U134 ( .A(n60), .B(in_17bit[2]), .Y(in_17bit_b[2]) );
  CLKINVX3 U135 ( .A(in_17bit[4]), .Y(n62) );
  XOR2X4 U136 ( .A(n65), .B(n4), .Y(in_17bit_b[5]) );
  CLKINVX3 U137 ( .A(n66), .Y(n68) );
  CLKINVX3 U138 ( .A(in_17bit[6]), .Y(n67) );
  XOR2X4 U139 ( .A(n71), .B(n69), .Y(in_17bit_b[7]) );
  CLKINVX3 U140 ( .A(in_17bit[8]), .Y(n72) );
  CLKINVX3 U141 ( .A(n74), .Y(n76) );
  CLKINVX3 U142 ( .A(in_17bit[10]), .Y(n78) );
  XNOR2X4 U143 ( .A(n77), .B(n78), .Y(in_17bit_b[10]) );
  NAND2X4 U144 ( .A(n35), .B(n78), .Y(n80) );
  CLKINVX3 U145 ( .A(in_17bit[12]), .Y(n83) );
  XNOR2X4 U146 ( .A(n82), .B(n83), .Y(in_17bit_b[12]) );
  CLKINVX3 U147 ( .A(n85), .Y(n87) );
  XNOR2X4 U148 ( .A(n88), .B(n89), .Y(in_17bit_b[14]) );
  CLKINVX3 U149 ( .A(in_17bit[15]), .Y(n90) );
  NOR3X4 U150 ( .A(in_17bit[15]), .B(n91), .C(n5), .Y(in_17bit_b[16]) );
  XNOR2X4 U151 ( .A(mul[9]), .B(n92), .Y(out[2]) );
  NAND2X4 U152 ( .A(n99), .B(n115), .Y(n98) );
  XNOR2X4 U153 ( .A(mul[13]), .B(n98), .Y(out[6]) );
  NAND2X4 U154 ( .A(n101), .B(n115), .Y(n100) );
  XNOR2X4 U155 ( .A(mul[14]), .B(n100), .Y(out[7]) );
  NAND2X4 U156 ( .A(n103), .B(n115), .Y(n102) );
  XNOR2X4 U157 ( .A(mul[15]), .B(n102), .Y(out[8]) );
  CLKINVX3 U158 ( .A(n106), .Y(n107) );
  NAND2BX4 U159 ( .AN(mul[17]), .B(n107), .Y(n109) );
  NAND2X4 U160 ( .A(n109), .B(n115), .Y(n108) );
  XNOR2X4 U161 ( .A(mul[18]), .B(n108), .Y(out[11]) );
endmodule


module multi16_1_DW01_add_0 ( A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, 
        A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, 
        B_20_, B_19_, B_18_, B_17_, B_16_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, 
        SUM_17_, SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, 
        SUM_9_, SUM_8_, SUM_7_, SUM_6_, SUM_5_ );
  input A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_,
         A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, B_20_, B_19_,
         B_18_, B_17_, B_16_;
  output SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, SUM_15_,
         SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, SUM_7_,
         SUM_6_, SUM_5_;
  wire   n1, n2, n3, n5, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41;

  INVX8 U2 ( .A(n32), .Y(n20) );
  NAND2X4 U3 ( .A(B_16_), .B(A_16_), .Y(n1) );
  AOI21X2 U4 ( .A0(n17), .A1(n34), .B0(n18), .Y(n29) );
  OAI21X4 U5 ( .A0(n29), .A1(n30), .B0(n31), .Y(n25) );
  BUFX12 U6 ( .A(A_11_), .Y(SUM_11_) );
  XNOR2X4 U7 ( .A(n2), .B(n3), .Y(SUM_18_) );
  AND2X4 U8 ( .A(n35), .B(n17), .Y(n2) );
  BUFX8 U9 ( .A(A_6_), .Y(SUM_6_) );
  CLKINVX8 U10 ( .A(n1), .Y(n21) );
  AOI21X2 U11 ( .A0(n21), .A1(n20), .B0(n19), .Y(n40) );
  AOI21X4 U12 ( .A0(n20), .A1(n21), .B0(n19), .Y(n3) );
  AOI21X1 U13 ( .A0(n25), .A1(n26), .B0(n16), .Y(n24) );
  OAI21X1 U14 ( .A0(n32), .A1(n36), .B0(n37), .Y(n34) );
  INVX8 U15 ( .A(n22), .Y(SUM_15_) );
  INVX8 U16 ( .A(n37), .Y(n19) );
  BUFX12 U17 ( .A(A_14_), .Y(SUM_14_) );
  INVX8 U18 ( .A(A_15_), .Y(n22) );
  NOR2BX4 U19 ( .AN(n31), .B(n30), .Y(n39) );
  NOR2X4 U20 ( .A(B_18_), .B(A_18_), .Y(n33) );
  NAND2X4 U21 ( .A(B_19_), .B(A_19_), .Y(n31) );
  NAND2X4 U22 ( .A(B_17_), .B(A_17_), .Y(n37) );
  NAND2X2 U23 ( .A(n27), .B(n26), .Y(n28) );
  OR2X4 U24 ( .A(B_20_), .B(A_20_), .Y(n26) );
  NOR2X2 U25 ( .A(A_16_), .B(B_16_), .Y(n5) );
  BUFX8 U26 ( .A(A_7_), .Y(SUM_7_) );
  NOR2X2 U27 ( .A(B_19_), .B(A_19_), .Y(n30) );
  BUFX12 U28 ( .A(A_10_), .Y(SUM_10_) );
  XNOR2X4 U29 ( .A(n28), .B(n25), .Y(SUM_20_) );
  OAI21X2 U30 ( .A0(n40), .A1(n33), .B0(n35), .Y(n38) );
  CLKINVX3 U31 ( .A(n35), .Y(n18) );
  NAND2X4 U32 ( .A(B_18_), .B(A_18_), .Y(n35) );
  NOR2BX4 U33 ( .AN(n36), .B(n5), .Y(SUM_16_) );
  INVX4 U34 ( .A(n33), .Y(n17) );
  INVXL U35 ( .A(n27), .Y(n16) );
  BUFX4 U36 ( .A(A_8_), .Y(SUM_8_) );
  BUFX8 U37 ( .A(A_12_), .Y(SUM_12_) );
  BUFX4 U38 ( .A(A_9_), .Y(SUM_9_) );
  BUFX8 U39 ( .A(A_5_), .Y(SUM_5_) );
  BUFX8 U40 ( .A(A_13_), .Y(SUM_13_) );
  NAND2X4 U41 ( .A(A_16_), .B(B_16_), .Y(n36) );
  XOR2X4 U42 ( .A(n38), .B(n39), .Y(SUM_19_) );
  XOR2X4 U43 ( .A(n41), .B(n21), .Y(SUM_17_) );
  NOR2X4 U44 ( .A(n19), .B(n32), .Y(n41) );
  NOR2X4 U45 ( .A(A_17_), .B(B_17_), .Y(n32) );
  XOR2X1 U46 ( .A(n23), .B(n24), .Y(SUM_21_) );
  XNOR2X1 U47 ( .A(B_21_), .B(A_21_), .Y(n23) );
  NAND2X1 U48 ( .A(B_20_), .B(A_20_), .Y(n27) );
endmodule


module multi16_1_DW02_mult_0 ( A, B, PRODUCT_23_, PRODUCT_22_, PRODUCT_21_, 
        PRODUCT_20_, PRODUCT_19_, PRODUCT_18_, PRODUCT_17_, PRODUCT_16_, 
        PRODUCT_15_, PRODUCT_14_, PRODUCT_13_, PRODUCT_12_, PRODUCT_11_, 
        PRODUCT_10_, PRODUCT_9_, PRODUCT_8_, PRODUCT_7_ );
  input [16:0] A;
  input [7:0] B;
  output PRODUCT_23_, PRODUCT_22_, PRODUCT_21_, PRODUCT_20_, PRODUCT_19_,
         PRODUCT_18_, PRODUCT_17_, PRODUCT_16_, PRODUCT_15_, PRODUCT_14_,
         PRODUCT_13_, PRODUCT_12_, PRODUCT_11_, PRODUCT_10_, PRODUCT_9_,
         PRODUCT_8_, PRODUCT_7_;
  wire   ab_16__7_, ab_16__6_, ab_16__5_, ab_16__4_, ab_16__3_, ab_16__2_,
         ab_16__1_, ab_16__0_, ab_15__7_, ab_15__6_, ab_15__5_, ab_15__4_,
         ab_15__3_, ab_15__2_, ab_15__1_, ab_15__0_, ab_14__7_, ab_14__6_,
         ab_14__5_, ab_14__4_, ab_14__3_, ab_14__2_, ab_14__1_, ab_14__0_,
         ab_13__7_, ab_13__6_, ab_13__5_, ab_13__4_, ab_13__3_, ab_13__2_,
         ab_13__1_, ab_13__0_, ab_12__7_, ab_12__6_, ab_12__5_, ab_12__4_,
         ab_12__3_, ab_12__2_, ab_12__1_, ab_12__0_, ab_11__7_, ab_11__6_,
         ab_11__5_, ab_11__4_, ab_11__3_, ab_11__2_, ab_11__1_, ab_11__0_,
         ab_10__7_, ab_10__6_, ab_10__5_, ab_10__4_, ab_10__3_, ab_10__2_,
         ab_10__1_, ab_10__0_, ab_9__7_, ab_9__6_, ab_9__5_, ab_9__4_,
         ab_9__3_, ab_9__2_, ab_9__1_, ab_9__0_, ab_8__7_, ab_8__6_, ab_8__5_,
         ab_8__4_, ab_8__3_, ab_8__2_, ab_8__1_, ab_8__0_, ab_7__7_, ab_7__6_,
         ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_, ab_7__0_, ab_6__7_,
         ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_, ab_6__1_, ab_6__0_,
         ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_, ab_5__2_, ab_5__1_,
         ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_, ab_4__3_, ab_4__2_,
         ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_, ab_3__4_, ab_3__3_,
         ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_, ab_2__5_, ab_2__4_,
         ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_, ab_1__6_, ab_1__5_,
         ab_1__4_, ab_1__3_, ab_1__2_, ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_,
         ab_0__3_, ab_0__2_, CARRYB_16__6_, CARRYB_16__5_, CARRYB_16__4_,
         CARRYB_16__3_, CARRYB_16__2_, CARRYB_16__1_, CARRYB_16__0_,
         CARRYB_15__6_, CARRYB_15__5_, CARRYB_15__4_, CARRYB_15__3_,
         CARRYB_15__2_, CARRYB_15__1_, CARRYB_15__0_, CARRYB_14__6_,
         CARRYB_14__5_, CARRYB_14__4_, CARRYB_14__3_, CARRYB_14__2_,
         CARRYB_14__1_, CARRYB_14__0_, CARRYB_13__6_, CARRYB_13__5_,
         CARRYB_13__4_, CARRYB_13__3_, CARRYB_13__2_, CARRYB_13__1_,
         CARRYB_13__0_, CARRYB_12__6_, CARRYB_12__5_, CARRYB_12__4_,
         CARRYB_12__3_, CARRYB_12__2_, CARRYB_12__1_, CARRYB_12__0_,
         CARRYB_11__6_, CARRYB_11__5_, CARRYB_11__4_, CARRYB_11__3_,
         CARRYB_11__2_, CARRYB_11__1_, CARRYB_11__0_, CARRYB_10__6_,
         CARRYB_10__5_, CARRYB_10__4_, CARRYB_10__3_, CARRYB_10__2_,
         CARRYB_10__1_, CARRYB_10__0_, CARRYB_9__6_, CARRYB_9__5_,
         CARRYB_9__4_, CARRYB_9__3_, CARRYB_9__2_, CARRYB_9__1_, CARRYB_9__0_,
         CARRYB_8__6_, CARRYB_8__5_, CARRYB_8__4_, CARRYB_8__3_, CARRYB_8__2_,
         CARRYB_8__1_, CARRYB_8__0_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_,
         CARRYB_7__3_, CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_,
         CARRYB_6__5_, CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_,
         CARRYB_6__0_, CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_,
         CARRYB_5__2_, CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_,
         CARRYB_4__4_, CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_,
         CARRYB_3__6_, CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_,
         CARRYB_3__1_, CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_,
         CARRYB_2__3_, CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__0_,
         SUMB_16__6_, SUMB_16__5_, SUMB_16__4_, SUMB_16__3_, SUMB_16__2_,
         SUMB_16__1_, SUMB_16__0_, SUMB_15__6_, SUMB_15__5_, SUMB_15__4_,
         SUMB_15__3_, SUMB_15__2_, SUMB_15__1_, SUMB_14__6_, SUMB_14__5_,
         SUMB_14__4_, SUMB_14__3_, SUMB_14__2_, SUMB_14__1_, SUMB_13__6_,
         SUMB_13__5_, SUMB_13__4_, SUMB_13__3_, SUMB_13__2_, SUMB_13__1_,
         SUMB_12__6_, SUMB_12__5_, SUMB_12__4_, SUMB_12__3_, SUMB_12__2_,
         SUMB_12__1_, SUMB_11__6_, SUMB_11__5_, SUMB_11__4_, SUMB_11__3_,
         SUMB_11__2_, SUMB_11__1_, SUMB_10__6_, SUMB_10__5_, SUMB_10__4_,
         SUMB_10__3_, SUMB_10__2_, SUMB_10__1_, SUMB_9__6_, SUMB_9__5_,
         SUMB_9__4_, SUMB_9__3_, SUMB_9__2_, SUMB_9__1_, SUMB_8__6_,
         SUMB_8__5_, SUMB_8__4_, SUMB_8__3_, SUMB_8__2_, SUMB_8__1_,
         SUMB_7__6_, SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_,
         SUMB_7__1_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, PROD1_7_, A1_21_, A1_20_, A1_19_, A1_18_,
         A1_17_, A1_16_, A1_15_, A1_13_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_,
         A1_7_, A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_16_, n3, n4, n5,
         n6, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45;

  multi16_1_DW01_add_0 FS_1 ( .A_21_(A1_21_), .A_20_(A1_20_), .A_19_(A1_19_), 
        .A_18_(A1_18_), .A_17_(A1_17_), .A_16_(A1_16_), .A_15_(A1_15_), 
        .A_14_(SUMB_16__0_), .A_13_(A1_13_), .A_12_(A1_12_), .A_11_(A1_11_), 
        .A_10_(A1_10_), .A_9_(A1_9_), .A_8_(A1_8_), .A_7_(A1_7_), .A_6_(A1_6_), 
        .A_5_(PROD1_7_), .B_21_(n18), .B_20_(n22), .B_19_(n21), .B_18_(n20), 
        .B_17_(n19), .B_16_(A2_16_), .SUM_21_(PRODUCT_23_), .SUM_20_(
        PRODUCT_22_), .SUM_19_(PRODUCT_21_), .SUM_18_(PRODUCT_20_), .SUM_17_(
        PRODUCT_19_), .SUM_16_(PRODUCT_18_), .SUM_15_(PRODUCT_17_), .SUM_14_(
        PRODUCT_16_), .SUM_13_(PRODUCT_15_), .SUM_12_(PRODUCT_14_), .SUM_11_(
        PRODUCT_13_), .SUM_10_(PRODUCT_12_), .SUM_9_(PRODUCT_11_), .SUM_8_(
        PRODUCT_10_), .SUM_7_(PRODUCT_9_), .SUM_6_(PRODUCT_8_), .SUM_5_(
        PRODUCT_7_) );
  ADDFHX4 S1_14_0 ( .A(ab_14__0_), .B(CARRYB_13__0_), .CI(SUMB_13__1_), .CO(
        CARRYB_14__0_), .S(A1_12_) );
  ADDFHX4 S1_15_0 ( .A(ab_15__0_), .B(CARRYB_14__0_), .CI(SUMB_14__1_), .CO(
        CARRYB_15__0_), .S(A1_13_) );
  ADDFHX4 S4_2 ( .A(ab_16__2_), .B(SUMB_15__3_), .CI(CARRYB_15__2_), .CO(
        CARRYB_16__2_), .S(SUMB_16__2_) );
  ADDFHX4 S1_8_0 ( .A(ab_8__0_), .B(CARRYB_7__0_), .CI(SUMB_7__1_), .CO(
        CARRYB_8__0_), .S(A1_6_) );
  ADDFHX4 S1_9_0 ( .A(ab_9__0_), .B(CARRYB_8__0_), .CI(SUMB_8__1_), .CO(
        CARRYB_9__0_), .S(A1_7_) );
  ADDFHX4 S2_14_3 ( .A(ab_14__3_), .B(SUMB_13__4_), .CI(CARRYB_13__3_), .CO(
        CARRYB_14__3_), .S(SUMB_14__3_) );
  ADDFHX4 S2_10_2 ( .A(ab_10__2_), .B(CARRYB_9__2_), .CI(SUMB_9__3_), .CO(
        CARRYB_10__2_), .S(SUMB_10__2_) );
  ADDFHX4 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  ADDFHX4 S1_7_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(PROD1_7_) );
  ADDFHX4 S1_11_0 ( .A(ab_11__0_), .B(CARRYB_10__0_), .CI(SUMB_10__1_), .CO(
        CARRYB_11__0_), .S(A1_9_) );
  ADDFHX4 S1_12_0 ( .A(ab_12__0_), .B(CARRYB_11__0_), .CI(SUMB_11__1_), .CO(
        CARRYB_12__0_), .S(A1_10_) );
  ADDFHX4 S2_15_1 ( .A(ab_15__1_), .B(CARRYB_14__1_), .CI(SUMB_14__2_), .CO(
        CARRYB_15__1_), .S(SUMB_15__1_) );
  ADDFHX4 S4_1 ( .A(ab_16__1_), .B(CARRYB_15__1_), .CI(SUMB_15__2_), .CO(
        CARRYB_16__1_), .S(SUMB_16__1_) );
  ADDFHX4 S2_11_5 ( .A(ab_11__5_), .B(CARRYB_10__5_), .CI(SUMB_10__6_), .CO(
        CARRYB_11__5_), .S(SUMB_11__5_) );
  ADDFHX4 S2_13_1 ( .A(ab_13__1_), .B(CARRYB_12__1_), .CI(SUMB_12__2_), .CO(
        CARRYB_13__1_), .S(SUMB_13__1_) );
  ADDFHX1 S3_14_6 ( .A(ab_14__6_), .B(CARRYB_13__6_), .CI(ab_13__7_), .CO(
        CARRYB_14__6_), .S(SUMB_14__6_) );
  ADDFHX4 S4_4 ( .A(ab_16__4_), .B(CARRYB_15__4_), .CI(SUMB_15__5_), .CO(
        CARRYB_16__4_), .S(SUMB_16__4_) );
  ADDFHX4 S2_12_5 ( .A(ab_12__5_), .B(CARRYB_11__5_), .CI(SUMB_11__6_), .CO(
        CARRYB_12__5_), .S(SUMB_12__5_) );
  ADDFHX4 S2_11_3 ( .A(ab_11__3_), .B(CARRYB_10__3_), .CI(SUMB_10__4_), .CO(
        CARRYB_11__3_), .S(SUMB_11__3_) );
  ADDFHX4 S2_10_1 ( .A(ab_10__1_), .B(CARRYB_9__1_), .CI(SUMB_9__2_), .CO(
        CARRYB_10__1_), .S(SUMB_10__1_) );
  ADDFHX4 S2_13_4 ( .A(ab_13__4_), .B(SUMB_12__5_), .CI(CARRYB_12__4_), .CO(
        CARRYB_13__4_), .S(SUMB_13__4_) );
  ADDFHX4 S2_8_5 ( .A(ab_8__5_), .B(SUMB_7__6_), .CI(CARRYB_7__5_), .CO(
        CARRYB_8__5_), .S(SUMB_8__5_) );
  ADDFHX4 S2_8_4 ( .A(ab_8__4_), .B(CARRYB_7__4_), .CI(SUMB_7__5_), .CO(
        CARRYB_8__4_), .S(SUMB_8__4_) );
  ADDFHX4 S2_2_3 ( .A(ab_2__3_), .B(n10), .CI(SUMB_1__4_), .CO(CARRYB_2__3_), 
        .S(SUMB_2__3_) );
  ADDFHX4 S2_9_3 ( .A(ab_9__3_), .B(CARRYB_8__3_), .CI(SUMB_8__4_), .CO(
        CARRYB_9__3_), .S(SUMB_9__3_) );
  ADDFHX4 S2_10_3 ( .A(ab_10__3_), .B(CARRYB_9__3_), .CI(SUMB_9__4_), .CO(
        CARRYB_10__3_), .S(SUMB_10__3_) );
  ADDFHX4 S2_11_2 ( .A(ab_11__2_), .B(CARRYB_10__2_), .CI(SUMB_10__3_), .CO(
        CARRYB_11__2_), .S(SUMB_11__2_) );
  ADDFHX4 S2_12_2 ( .A(ab_12__2_), .B(CARRYB_11__2_), .CI(SUMB_11__3_), .CO(
        CARRYB_12__2_), .S(SUMB_12__2_) );
  ADDFHX4 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  ADDFHX4 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  ADDFHX4 S2_8_1 ( .A(ab_8__1_), .B(CARRYB_7__1_), .CI(SUMB_7__2_), .CO(
        CARRYB_8__1_), .S(SUMB_8__1_) );
  ADDFHX4 S2_11_1 ( .A(ab_11__1_), .B(CARRYB_10__1_), .CI(SUMB_10__2_), .CO(
        CARRYB_11__1_), .S(SUMB_11__1_) );
  ADDFHX4 S2_7_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  ADDFHX4 S2_9_5 ( .A(ab_9__5_), .B(CARRYB_8__5_), .CI(SUMB_8__6_), .CO(
        CARRYB_9__5_), .S(SUMB_9__5_) );
  ADDFHX4 S2_10_5 ( .A(ab_10__5_), .B(SUMB_9__6_), .CI(CARRYB_9__5_), .CO(
        CARRYB_10__5_), .S(SUMB_10__5_) );
  ADDFHX2 S2_15_5 ( .A(ab_15__5_), .B(CARRYB_14__5_), .CI(SUMB_14__6_), .CO(
        CARRYB_15__5_), .S(SUMB_15__5_) );
  ADDFHX4 S4_5 ( .A(ab_16__5_), .B(CARRYB_15__5_), .CI(SUMB_15__6_), .CO(
        CARRYB_16__5_), .S(SUMB_16__5_) );
  ADDFHX4 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  ADDFHX4 S2_15_4 ( .A(ab_15__4_), .B(CARRYB_14__4_), .CI(SUMB_14__5_), .CO(
        CARRYB_15__4_), .S(SUMB_15__4_) );
  ADDFHX4 S4_3 ( .A(ab_16__3_), .B(CARRYB_15__3_), .CI(SUMB_15__4_), .CO(
        CARRYB_16__3_), .S(SUMB_16__3_) );
  ADDFHX4 S3_3_6 ( .A(ab_3__6_), .B(ab_2__7_), .CI(CARRYB_2__6_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  ADDFHX4 S2_9_2 ( .A(ab_9__2_), .B(CARRYB_8__2_), .CI(SUMB_8__3_), .CO(
        CARRYB_9__2_), .S(SUMB_9__2_) );
  ADDFHX4 S2_12_1 ( .A(ab_12__1_), .B(CARRYB_11__1_), .CI(SUMB_11__2_), .CO(
        CARRYB_12__1_), .S(SUMB_12__1_) );
  ADDFHX4 S2_7_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  ADDFHX4 S2_13_2 ( .A(ab_13__2_), .B(CARRYB_12__2_), .CI(SUMB_12__3_), .CO(
        CARRYB_13__2_), .S(SUMB_13__2_) );
  ADDFHX4 S2_14_1 ( .A(ab_14__1_), .B(CARRYB_13__1_), .CI(SUMB_13__2_), .CO(
        CARRYB_14__1_), .S(SUMB_14__1_) );
  ADDFHX4 S2_7_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  ADDFHX4 S2_8_3 ( .A(ab_8__3_), .B(CARRYB_7__3_), .CI(SUMB_7__4_), .CO(
        CARRYB_8__3_), .S(SUMB_8__3_) );
  ADDFHX4 S1_13_0 ( .A(ab_13__0_), .B(CARRYB_12__0_), .CI(SUMB_12__1_), .CO(
        CARRYB_13__0_), .S(A1_11_) );
  ADDFHX4 S4_0 ( .A(ab_16__0_), .B(CARRYB_15__0_), .CI(SUMB_15__1_), .CO(
        CARRYB_16__0_), .S(SUMB_16__0_) );
  ADDFHX4 S3_10_6 ( .A(ab_10__6_), .B(CARRYB_9__6_), .CI(ab_9__7_), .CO(
        CARRYB_10__6_), .S(SUMB_10__6_) );
  ADDFHX4 S3_11_6 ( .A(ab_11__6_), .B(CARRYB_10__6_), .CI(ab_10__7_), .CO(
        CARRYB_11__6_), .S(SUMB_11__6_) );
  ADDFHX2 S3_12_6 ( .A(ab_12__6_), .B(CARRYB_11__6_), .CI(ab_11__7_), .CO(
        CARRYB_12__6_), .S(SUMB_12__6_) );
  ADDFHX4 S2_6_5 ( .A(ab_6__5_), .B(SUMB_5__6_), .CI(CARRYB_5__5_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  ADDFHX2 S2_14_5 ( .A(ab_14__5_), .B(CARRYB_13__5_), .CI(SUMB_13__6_), .CO(
        CARRYB_14__5_), .S(SUMB_14__5_) );
  ADDFHX4 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  ADDFHX4 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  ADDFHX4 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  ADDFHX4 S2_14_4 ( .A(ab_14__4_), .B(CARRYB_13__4_), .CI(SUMB_13__5_), .CO(
        CARRYB_14__4_), .S(SUMB_14__4_) );
  ADDFHX4 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  ADDFHX4 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  ADDFHX4 S2_12_3 ( .A(ab_12__3_), .B(CARRYB_11__3_), .CI(SUMB_11__4_), .CO(
        CARRYB_12__3_), .S(SUMB_12__3_) );
  ADDFHX4 S2_14_2 ( .A(ab_14__2_), .B(CARRYB_13__2_), .CI(SUMB_13__3_), .CO(
        CARRYB_14__2_), .S(SUMB_14__2_) );
  ADDFHX4 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  ADDFHX4 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  ADDFHX4 S2_7_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  ADDFHX4 S2_11_4 ( .A(ab_11__4_), .B(SUMB_10__5_), .CI(CARRYB_10__4_), .CO(
        CARRYB_11__4_), .S(SUMB_11__4_) );
  ADDFHX4 S2_13_5 ( .A(ab_13__5_), .B(CARRYB_12__5_), .CI(SUMB_12__6_), .CO(
        CARRYB_13__5_), .S(SUMB_13__5_) );
  ADDFHX4 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  ADDFHX4 S2_9_1 ( .A(ab_9__1_), .B(CARRYB_8__1_), .CI(SUMB_8__2_), .CO(
        CARRYB_9__1_), .S(SUMB_9__1_) );
  ADDFHX4 S1_10_0 ( .A(ab_10__0_), .B(CARRYB_9__0_), .CI(SUMB_9__1_), .CO(
        CARRYB_10__0_), .S(A1_8_) );
  ADDFHX4 S3_9_6 ( .A(ab_9__6_), .B(CARRYB_8__6_), .CI(ab_8__7_), .CO(
        CARRYB_9__6_), .S(SUMB_9__6_) );
  ADDFHX4 S3_13_6 ( .A(ab_13__6_), .B(CARRYB_12__6_), .CI(ab_12__7_), .CO(
        CARRYB_13__6_), .S(SUMB_13__6_) );
  ADDFHX4 S2_2_5 ( .A(ab_2__5_), .B(n12), .CI(SUMB_1__6_), .CO(CARRYB_2__5_), 
        .S(SUMB_2__5_) );
  ADDFHX4 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  ADDFHX4 S2_15_3 ( .A(ab_15__3_), .B(CARRYB_14__3_), .CI(SUMB_14__4_), .CO(
        CARRYB_15__3_), .S(SUMB_15__3_) );
  ADDFHX4 S2_8_2 ( .A(ab_8__2_), .B(CARRYB_7__2_), .CI(SUMB_7__3_), .CO(
        CARRYB_8__2_), .S(SUMB_8__2_) );
  ADDFHX4 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  ADDFHX4 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  ADDFHX4 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  ADDFHX4 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  ADDFHX4 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  ADDFHX4 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  ADDFHX4 S2_2_4 ( .A(ab_2__4_), .B(n8), .CI(SUMB_1__5_), .CO(CARRYB_2__4_), 
        .S(SUMB_2__4_) );
  ADDFHX4 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  ADDFHX4 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  ADDFHX4 S3_8_6 ( .A(ab_8__6_), .B(CARRYB_7__6_), .CI(ab_7__7_), .CO(
        CARRYB_8__6_), .S(SUMB_8__6_) );
  ADDFHX4 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  ADDFHX4 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  ADDFHX4 S2_2_2 ( .A(ab_2__2_), .B(n6), .CI(SUMB_1__3_), .CO(CARRYB_2__2_), 
        .S(SUMB_2__2_) );
  ADDFHX4 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  ADDFHX4 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  ADDFHX4 S2_2_1 ( .A(ab_2__1_), .B(n9), .CI(SUMB_1__2_), .CO(CARRYB_2__1_), 
        .S(SUMB_2__1_) );
  ADDFHX4 S3_15_6 ( .A(ab_15__6_), .B(CARRYB_14__6_), .CI(ab_14__7_), .CO(
        CARRYB_15__6_), .S(SUMB_15__6_) );
  ADDFHX4 S5_6 ( .A(ab_16__6_), .B(CARRYB_15__6_), .CI(ab_15__7_), .CO(
        CARRYB_16__6_), .S(SUMB_16__6_) );
  ADDFHX4 S3_7_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(
        CARRYB_7__6_), .S(SUMB_7__6_) );
  ADDFHX2 S2_12_4 ( .A(ab_12__4_), .B(CARRYB_11__4_), .CI(SUMB_11__5_), .CO(
        CARRYB_12__4_), .S(SUMB_12__4_) );
  ADDFHX4 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  ADDFHX4 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  ADDFHX2 S2_15_2 ( .A(ab_15__2_), .B(CARRYB_14__2_), .CI(SUMB_14__3_), .CO(
        CARRYB_15__2_), .S(SUMB_15__2_) );
  ADDFHX2 S2_10_4 ( .A(ab_10__4_), .B(SUMB_9__5_), .CI(CARRYB_9__4_), .CO(
        CARRYB_10__4_), .S(SUMB_10__4_) );
  ADDFHX2 S3_2_6 ( .A(ab_2__6_), .B(n11), .CI(ab_1__7_), .CO(CARRYB_2__6_), 
        .S(SUMB_2__6_) );
  ADDFHX2 S2_13_3 ( .A(ab_13__3_), .B(CARRYB_12__3_), .CI(SUMB_12__4_), .CO(
        CARRYB_13__3_), .S(SUMB_13__3_) );
  ADDFHX4 S2_7_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  NOR2BX4 U2 ( .AN(A[1]), .B(n30), .Y(n3) );
  NOR2BX2 U3 ( .AN(A[1]), .B(n30), .Y(ab_1__2_) );
  AND2X4 U4 ( .A(A[1]), .B(B[1]), .Y(n45) );
  NOR2BX1 U5 ( .AN(n13), .B(n44), .Y(ab_2__7_) );
  NOR2BX2 U6 ( .AN(n13), .B(n24), .Y(ab_2__5_) );
  AND2X2 U7 ( .A(n13), .B(n4), .Y(ab_2__0_) );
  XOR2X4 U8 ( .A(ab_1__4_), .B(ab_0__5_), .Y(SUMB_1__4_) );
  CLKINVX20 U9 ( .A(n43), .Y(n4) );
  XOR2X4 U10 ( .A(n45), .B(ab_0__2_), .Y(SUMB_1__1_) );
  BUFX12 U11 ( .A(A[3]), .Y(n5) );
  AND2X4 U12 ( .A(ab_1__2_), .B(ab_0__3_), .Y(n6) );
  BUFX20 U13 ( .A(A[2]), .Y(n13) );
  NOR2BX2 U14 ( .AN(n5), .B(n26), .Y(ab_3__4_) );
  NOR2BX1 U15 ( .AN(A[9]), .B(n29), .Y(ab_9__3_) );
  NOR2BX1 U16 ( .AN(A[13]), .B(n31), .Y(ab_13__2_) );
  NOR2BX1 U17 ( .AN(A[11]), .B(n31), .Y(ab_11__2_) );
  NOR2BX2 U18 ( .AN(A[4]), .B(n32), .Y(ab_4__1_) );
  NOR2BX1 U19 ( .AN(A[10]), .B(n29), .Y(ab_10__3_) );
  NOR2BX1 U20 ( .AN(A[9]), .B(n31), .Y(ab_9__2_) );
  NOR2BX1 U21 ( .AN(A[14]), .B(n29), .Y(ab_14__3_) );
  NOR2BX1 U22 ( .AN(A[14]), .B(n33), .Y(ab_14__1_) );
  NOR2BX1 U23 ( .AN(A[9]), .B(n33), .Y(ab_9__1_) );
  NOR2BX1 U24 ( .AN(A[14]), .B(n43), .Y(ab_14__0_) );
  NOR2BX1 U25 ( .AN(A[3]), .B(n43), .Y(ab_3__0_) );
  NOR2BX2 U26 ( .AN(A[5]), .B(n32), .Y(ab_5__1_) );
  NOR2BX1 U27 ( .AN(A[9]), .B(n25), .Y(ab_9__5_) );
  NOR2BX1 U28 ( .AN(A[10]), .B(n31), .Y(ab_10__2_) );
  NOR2BX1 U29 ( .AN(A[14]), .B(n31), .Y(ab_14__2_) );
  NOR2BX1 U30 ( .AN(A[10]), .B(n33), .Y(ab_10__1_) );
  NOR2BX1 U31 ( .AN(A[15]), .B(n43), .Y(ab_15__0_) );
  NOR2BX1 U32 ( .AN(A[4]), .B(n43), .Y(ab_4__0_) );
  NOR2BX2 U33 ( .AN(A[6]), .B(n32), .Y(ab_6__1_) );
  AND2X4 U35 ( .A(ab_0__5_), .B(ab_1__4_), .Y(n8) );
  AND2X4 U36 ( .A(n45), .B(ab_0__2_), .Y(n9) );
  AND2X4 U37 ( .A(ab_0__4_), .B(ab_1__3_), .Y(n10) );
  AND2X4 U38 ( .A(ab_0__7_), .B(ab_1__6_), .Y(n11) );
  AND2X4 U39 ( .A(ab_0__6_), .B(ab_1__5_), .Y(n12) );
  BUFX20 U40 ( .A(n42), .Y(n32) );
  NOR2BX4 U41 ( .AN(B[4]), .B(n35), .Y(ab_0__4_) );
  INVX4 U42 ( .A(B[0]), .Y(n43) );
  NAND2X4 U43 ( .A(CARRYB_16__0_), .B(SUMB_16__1_), .Y(n23) );
  XOR2X4 U44 ( .A(ab_1__3_), .B(ab_0__4_), .Y(SUMB_1__3_) );
  INVX12 U45 ( .A(A[0]), .Y(n35) );
  NOR2BX4 U46 ( .AN(n5), .B(n34), .Y(ab_3__6_) );
  INVX4 U47 ( .A(B[6]), .Y(n37) );
  XOR2X2 U48 ( .A(ab_1__5_), .B(ab_0__6_), .Y(SUMB_1__5_) );
  NAND2X2 U49 ( .A(ab_9__4_), .B(CARRYB_8__4_), .Y(n16) );
  NOR2BX1 U50 ( .AN(A[7]), .B(n44), .Y(ab_7__7_) );
  NOR2BX1 U51 ( .AN(A[7]), .B(n32), .Y(ab_7__1_) );
  NOR2BX1 U52 ( .AN(A[7]), .B(n26), .Y(ab_7__4_) );
  NOR2BX1 U53 ( .AN(A[7]), .B(n28), .Y(ab_7__3_) );
  NOR2BX1 U54 ( .AN(A[7]), .B(n30), .Y(ab_7__2_) );
  NOR2BX1 U55 ( .AN(A[7]), .B(n24), .Y(ab_7__5_) );
  NOR2BX1 U56 ( .AN(A[7]), .B(n34), .Y(ab_7__6_) );
  BUFX20 U57 ( .A(n38), .Y(n24) );
  NOR2BX2 U58 ( .AN(n5), .B(n28), .Y(ab_3__3_) );
  NOR2BX1 U59 ( .AN(A[5]), .B(n24), .Y(ab_5__5_) );
  BUFX16 U60 ( .A(n40), .Y(n28) );
  NOR2BX4 U61 ( .AN(n13), .B(n28), .Y(ab_2__3_) );
  NOR2BX2 U62 ( .AN(A[4]), .B(n24), .Y(ab_4__5_) );
  NOR2BX2 U63 ( .AN(A[4]), .B(n34), .Y(ab_4__6_) );
  NOR2BX2 U64 ( .AN(B[2]), .B(n35), .Y(ab_0__2_) );
  CLKINVX8 U65 ( .A(B[1]), .Y(n42) );
  NOR2BX2 U66 ( .AN(n5), .B(n30), .Y(ab_3__2_) );
  BUFX20 U67 ( .A(n41), .Y(n30) );
  NAND2X2 U68 ( .A(ab_9__4_), .B(SUMB_8__5_), .Y(n17) );
  NOR2BX4 U69 ( .AN(n13), .B(n30), .Y(ab_2__2_) );
  NOR2BX2 U70 ( .AN(A[4]), .B(n28), .Y(ab_4__3_) );
  NOR2BX2 U71 ( .AN(A[4]), .B(n26), .Y(ab_4__4_) );
  NOR2BX2 U72 ( .AN(B[3]), .B(n35), .Y(ab_0__3_) );
  NOR2BX2 U73 ( .AN(n5), .B(n32), .Y(ab_3__1_) );
  NOR2BX2 U74 ( .AN(A[4]), .B(n30), .Y(ab_4__2_) );
  INVX4 U75 ( .A(B[5]), .Y(n38) );
  NOR2BX2 U76 ( .AN(B[5]), .B(n35), .Y(ab_0__5_) );
  NAND2X2 U77 ( .A(SUMB_8__5_), .B(CARRYB_8__4_), .Y(n15) );
  XOR2X4 U78 ( .A(CARRYB_8__4_), .B(n14), .Y(SUMB_9__4_) );
  NOR2BX4 U79 ( .AN(n13), .B(n32), .Y(ab_2__1_) );
  XOR2X4 U80 ( .A(n3), .B(ab_0__3_), .Y(SUMB_1__2_) );
  NOR2BX1 U81 ( .AN(n5), .B(n44), .Y(ab_3__7_) );
  AND2X4 U82 ( .A(CARRYB_16__1_), .B(SUMB_16__2_), .Y(n19) );
  NOR2BX2 U83 ( .AN(n5), .B(n24), .Y(ab_3__5_) );
  INVX4 U84 ( .A(B[3]), .Y(n40) );
  NOR2BX2 U85 ( .AN(A[6]), .B(n24), .Y(ab_6__5_) );
  AND2X4 U86 ( .A(A[1]), .B(B[6]), .Y(ab_1__6_) );
  NOR2BX1 U87 ( .AN(A[6]), .B(n34), .Y(ab_6__6_) );
  NOR2BX4 U88 ( .AN(n13), .B(n34), .Y(ab_2__6_) );
  NOR2BX2 U89 ( .AN(A[8]), .B(n32), .Y(ab_8__1_) );
  NOR2BX4 U90 ( .AN(A[9]), .B(n27), .Y(ab_9__4_) );
  XOR2X4 U91 ( .A(CARRYB_16__5_), .B(SUMB_16__6_), .Y(A1_20_) );
  INVX20 U92 ( .A(B[7]), .Y(n44) );
  NOR2BX2 U93 ( .AN(A[5]), .B(n44), .Y(ab_5__7_) );
  NOR2BX2 U94 ( .AN(A[6]), .B(n44), .Y(ab_6__7_) );
  NOR2BX2 U95 ( .AN(A[8]), .B(n44), .Y(ab_8__7_) );
  BUFX20 U96 ( .A(n39), .Y(n26) );
  INVX8 U97 ( .A(B[4]), .Y(n39) );
  INVX4 U98 ( .A(n23), .Y(A2_16_) );
  NOR2BX2 U99 ( .AN(n13), .B(n26), .Y(ab_2__4_) );
  XOR2X2 U100 ( .A(ab_1__6_), .B(ab_0__7_), .Y(SUMB_1__6_) );
  NOR2BX4 U101 ( .AN(A[1]), .B(n24), .Y(ab_1__5_) );
  BUFX20 U102 ( .A(n37), .Y(n34) );
  XOR2X4 U103 ( .A(SUMB_16__1_), .B(CARRYB_16__0_), .Y(A1_15_) );
  NOR2BX2 U104 ( .AN(A[5]), .B(n34), .Y(ab_5__6_) );
  XOR2X4 U105 ( .A(CARRYB_16__4_), .B(SUMB_16__5_), .Y(A1_19_) );
  XOR2X4 U106 ( .A(SUMB_8__5_), .B(ab_9__4_), .Y(n14) );
  NAND3X4 U107 ( .A(n17), .B(n15), .C(n16), .Y(CARRYB_9__4_) );
  NOR2BX4 U108 ( .AN(B[6]), .B(n35), .Y(ab_0__6_) );
  NOR2BX1 U109 ( .AN(A[13]), .B(n43), .Y(ab_13__0_) );
  NOR2BX1 U110 ( .AN(A[13]), .B(n33), .Y(ab_13__1_) );
  NOR2BX1 U111 ( .AN(A[15]), .B(n33), .Y(ab_15__1_) );
  NOR2BX1 U112 ( .AN(A[10]), .B(n43), .Y(ab_10__0_) );
  NOR2BXL U113 ( .AN(A[8]), .B(n24), .Y(ab_8__5_) );
  NOR2BX1 U114 ( .AN(A[11]), .B(n43), .Y(ab_11__0_) );
  NOR2BX1 U115 ( .AN(A[15]), .B(n29), .Y(ab_15__3_) );
  CLKBUFXL U116 ( .A(n40), .Y(n29) );
  NOR2BX1 U117 ( .AN(A[13]), .B(n29), .Y(ab_13__3_) );
  NOR2BX1 U118 ( .AN(A[11]), .B(n29), .Y(ab_11__3_) );
  NOR2BX1 U119 ( .AN(A[12]), .B(n31), .Y(ab_12__2_) );
  NOR2BX1 U120 ( .AN(A[10]), .B(n25), .Y(ab_10__5_) );
  NOR2BX1 U121 ( .AN(A[12]), .B(n33), .Y(ab_12__1_) );
  NOR2BX1 U122 ( .AN(A[12]), .B(n25), .Y(ab_12__5_) );
  NOR2BX1 U123 ( .AN(A[8]), .B(n43), .Y(ab_8__0_) );
  AND2X1 U124 ( .A(CARRYB_16__4_), .B(SUMB_16__5_), .Y(n22) );
  NOR2BX1 U125 ( .AN(A[11]), .B(n33), .Y(ab_11__1_) );
  NOR2BX1 U126 ( .AN(A[6]), .B(n43), .Y(ab_6__0_) );
  NOR2BX1 U127 ( .AN(A[7]), .B(n43), .Y(ab_7__0_) );
  NOR2BX1 U128 ( .AN(A[12]), .B(n43), .Y(ab_12__0_) );
  AND2X1 U129 ( .A(CARRYB_16__5_), .B(SUMB_16__6_), .Y(n18) );
  NOR2BX1 U130 ( .AN(A[16]), .B(n27), .Y(ab_16__4_) );
  NOR2BX1 U131 ( .AN(A[16]), .B(n29), .Y(ab_16__3_) );
  NOR2BXL U132 ( .AN(A[11]), .B(n34), .Y(ab_11__6_) );
  NOR2BXL U133 ( .AN(A[10]), .B(n34), .Y(ab_10__6_) );
  NOR2BXL U134 ( .AN(A[9]), .B(n34), .Y(ab_9__6_) );
  NOR2BXL U135 ( .AN(A[12]), .B(n34), .Y(ab_12__6_) );
  NOR2BX1 U136 ( .AN(A[16]), .B(n33), .Y(ab_16__1_) );
  NOR2BX1 U137 ( .AN(A[15]), .B(n31), .Y(ab_15__2_) );
  AND3X1 U138 ( .A(A[1]), .B(B[1]), .C(n36), .Y(CARRYB_1__0_) );
  NOR2BXL U139 ( .AN(A[14]), .B(n34), .Y(ab_14__6_) );
  BUFX3 U140 ( .A(n39), .Y(n27) );
  CLKBUFXL U141 ( .A(n38), .Y(n25) );
  BUFX3 U142 ( .A(n42), .Y(n33) );
  BUFX1 U143 ( .A(n41), .Y(n31) );
  NOR2BXL U144 ( .AN(A[6]), .B(n26), .Y(ab_6__4_) );
  NOR2BXL U145 ( .AN(A[8]), .B(n26), .Y(ab_8__4_) );
  NOR2BXL U146 ( .AN(A[5]), .B(n43), .Y(ab_5__0_) );
  NOR2BXL U147 ( .AN(A[8]), .B(n28), .Y(ab_8__3_) );
  NOR2BXL U148 ( .AN(A[6]), .B(n28), .Y(ab_6__3_) );
  NOR2BXL U149 ( .AN(A[5]), .B(n26), .Y(ab_5__4_) );
  NOR2BXL U150 ( .AN(A[5]), .B(n28), .Y(ab_5__3_) );
  AND2X2 U151 ( .A(CARRYB_16__2_), .B(SUMB_16__3_), .Y(n20) );
  AND2X2 U152 ( .A(CARRYB_16__3_), .B(SUMB_16__4_), .Y(n21) );
  NOR2BX1 U153 ( .AN(A[11]), .B(n27), .Y(ab_11__4_) );
  NOR2BXL U154 ( .AN(A[12]), .B(n27), .Y(ab_12__4_) );
  NOR2BX1 U155 ( .AN(A[13]), .B(n27), .Y(ab_13__4_) );
  NOR2BX1 U156 ( .AN(A[11]), .B(n25), .Y(ab_11__5_) );
  NOR2BXL U157 ( .AN(A[8]), .B(n30), .Y(ab_8__2_) );
  NOR2BXL U158 ( .AN(A[6]), .B(n30), .Y(ab_6__2_) );
  NOR2BXL U159 ( .AN(A[5]), .B(n30), .Y(ab_5__2_) );
  NOR2BXL U160 ( .AN(A[9]), .B(n43), .Y(ab_9__0_) );
  NOR2BX1 U161 ( .AN(A[10]), .B(n27), .Y(ab_10__4_) );
  NOR2BX1 U162 ( .AN(A[13]), .B(n25), .Y(ab_13__5_) );
  NOR2BX1 U163 ( .AN(A[14]), .B(n25), .Y(ab_14__5_) );
  NOR2BX2 U164 ( .AN(A[14]), .B(n27), .Y(ab_14__4_) );
  NOR2BXL U165 ( .AN(A[12]), .B(n29), .Y(ab_12__3_) );
  XOR2X1 U166 ( .A(CARRYB_16__6_), .B(ab_16__7_), .Y(A1_21_) );
  NOR2BXL U167 ( .AN(A[16]), .B(n25), .Y(ab_16__5_) );
  NOR2BX1 U168 ( .AN(A[16]), .B(n34), .Y(ab_16__6_) );
  NOR2BX1 U169 ( .AN(A[15]), .B(n44), .Y(ab_15__7_) );
  NOR2BX1 U170 ( .AN(A[9]), .B(n44), .Y(ab_9__7_) );
  NOR2BX1 U171 ( .AN(A[13]), .B(n34), .Y(ab_13__6_) );
  NOR2BX1 U172 ( .AN(A[12]), .B(n44), .Y(ab_12__7_) );
  NOR2BX1 U173 ( .AN(A[15]), .B(n34), .Y(ab_15__6_) );
  NOR2BX1 U174 ( .AN(A[14]), .B(n44), .Y(ab_14__7_) );
  NOR2BX1 U175 ( .AN(A[8]), .B(n34), .Y(ab_8__6_) );
  NOR2BX1 U176 ( .AN(A[11]), .B(n44), .Y(ab_11__7_) );
  NOR2BXL U177 ( .AN(A[16]), .B(n31), .Y(ab_16__2_) );
  NOR2BXL U178 ( .AN(A[16]), .B(n43), .Y(ab_16__0_) );
  NOR2BX1 U179 ( .AN(A[1]), .B(n44), .Y(ab_1__7_) );
  NOR2BXL U180 ( .AN(A[15]), .B(n25), .Y(ab_15__5_) );
  NOR2BX1 U181 ( .AN(A[13]), .B(n44), .Y(ab_13__7_) );
  NOR2BX1 U182 ( .AN(A[4]), .B(n44), .Y(ab_4__7_) );
  NOR2BX1 U183 ( .AN(A[10]), .B(n44), .Y(ab_10__7_) );
  NOR2BXL U184 ( .AN(A[15]), .B(n27), .Y(ab_15__4_) );
  NOR2BX1 U185 ( .AN(A[16]), .B(n44), .Y(ab_16__7_) );
  NOR2BX1 U186 ( .AN(A[0]), .B(n43), .Y(n36) );
  XOR2X4 U187 ( .A(CARRYB_16__2_), .B(SUMB_16__3_), .Y(A1_17_) );
  XOR2X4 U188 ( .A(SUMB_16__2_), .B(CARRYB_16__1_), .Y(A1_16_) );
  XOR2X4 U189 ( .A(CARRYB_16__3_), .B(SUMB_16__4_), .Y(A1_18_) );
  INVX8 U190 ( .A(B[2]), .Y(n41) );
  NOR2BX4 U191 ( .AN(B[7]), .B(n35), .Y(ab_0__7_) );
  NOR2BX4 U192 ( .AN(A[1]), .B(n26), .Y(ab_1__4_) );
  NOR2BX4 U193 ( .AN(A[1]), .B(n28), .Y(ab_1__3_) );
endmodule


module multi16_1 ( in_17bit, in_8bit, out );
  input [16:0] in_17bit;
  input [7:0] in_8bit;
  output [16:0] out;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124;
  wire   [16:1] in_17bit_b;
  wire   [7:1] in_8bit_b;
  wire   [23:8] mul;

  multi16_1_DW02_mult_0 mult_55 ( .A({in_17bit_b[16:8], n3, in_17bit_b[6:2], 
        n44, in_17bit[0]}), .B({in_8bit_b, in_8bit[0]}), .PRODUCT_23_(mul[23]), 
        .PRODUCT_22_(mul[22]), .PRODUCT_21_(mul[21]), .PRODUCT_20_(mul[20]), 
        .PRODUCT_19_(mul[19]), .PRODUCT_18_(mul[18]), .PRODUCT_17_(mul[17]), 
        .PRODUCT_16_(mul[16]), .PRODUCT_15_(mul[15]), .PRODUCT_14_(mul[14]), 
        .PRODUCT_13_(mul[13]), .PRODUCT_12_(mul[12]), .PRODUCT_11_(mul[11]), 
        .PRODUCT_10_(mul[10]), .PRODUCT_9_(mul[9]), .PRODUCT_8_(mul[8]), 
        .PRODUCT_7_(out[0]) );
  BUFX20 U2 ( .A(in_17bit_b[1]), .Y(n44) );
  NOR2X4 U3 ( .A(in_17bit[1]), .B(in_17bit[0]), .Y(n1) );
  NAND3X1 U4 ( .A(n51), .B(n62), .C(n46), .Y(n2) );
  INVX8 U5 ( .A(in_8bit[5]), .Y(n46) );
  INVXL U6 ( .A(in_8bit[7]), .Y(n48) );
  BUFX8 U7 ( .A(in_17bit_b[7]), .Y(n3) );
  INVX3 U8 ( .A(n112), .Y(n5) );
  AND2X1 U9 ( .A(n45), .B(n76), .Y(n39) );
  INVX12 U10 ( .A(n45), .Y(n94) );
  INVX1 U11 ( .A(in_8bit[7]), .Y(n49) );
  NOR2X4 U12 ( .A(mul[16]), .B(n108), .Y(n4) );
  INVXL U13 ( .A(in_17bit[9]), .Y(n81) );
  INVX16 U14 ( .A(n49), .Y(n47) );
  AND2X4 U15 ( .A(in_17bit[1]), .B(in_17bit[0]), .Y(n67) );
  CLKINVX2 U16 ( .A(n11), .Y(n6) );
  INVX2 U17 ( .A(in_17bit[13]), .Y(n91) );
  INVX4 U18 ( .A(in_8bit[3]), .Y(n10) );
  NOR2X4 U19 ( .A(in_8bit[3]), .B(in_8bit[2]), .Y(n58) );
  BUFX20 U20 ( .A(in_17bit[16]), .Y(n45) );
  INVX4 U21 ( .A(n10), .Y(n11) );
  NOR2X1 U22 ( .A(mul[22]), .B(mul[21]), .Y(n123) );
  CLKINVX8 U23 ( .A(n116), .Y(n112) );
  BUFX8 U24 ( .A(mul[19]), .Y(n12) );
  AOI21X2 U25 ( .A0(n117), .A1(n118), .B0(n121), .Y(n119) );
  NOR2XL U26 ( .A(n40), .B(n94), .Y(n82) );
  OR2X2 U27 ( .A(n41), .B(n94), .Y(n36) );
  NAND2X2 U28 ( .A(n45), .B(n70), .Y(n69) );
  XNOR2X2 U29 ( .A(mul[11]), .B(n99), .Y(out[4]) );
  INVX8 U30 ( .A(in_17bit[2]), .Y(n68) );
  XOR2X4 U31 ( .A(n54), .B(n6), .Y(in_8bit_b[3]) );
  INVX8 U32 ( .A(n45), .Y(n7) );
  CLKINVX8 U33 ( .A(n61), .Y(n62) );
  OR2X4 U34 ( .A(in_8bit[2]), .B(in_8bit[0]), .Y(n55) );
  OAI21X4 U35 ( .A0(n21), .A1(in_8bit[0]), .B0(n47), .Y(n53) );
  XOR2X4 U36 ( .A(in_8bit[1]), .B(n33), .Y(in_8bit_b[1]) );
  AND2X4 U37 ( .A(in_8bit[0]), .B(n47), .Y(n33) );
  AOI21X4 U38 ( .A0(n67), .A1(n45), .B0(n66), .Y(in_17bit_b[1]) );
  INVX3 U39 ( .A(mul[17]), .Y(n17) );
  NAND3X4 U40 ( .A(n51), .B(n62), .C(n46), .Y(n65) );
  NOR2X1 U41 ( .A(n38), .B(n94), .Y(n87) );
  OAI21X4 U42 ( .A0(n21), .A1(n55), .B0(n47), .Y(n54) );
  XNOR2X4 U43 ( .A(mul[13]), .B(n25), .Y(out[6]) );
  NAND2X2 U44 ( .A(n103), .B(n113), .Y(n25) );
  XOR2X4 U45 ( .A(mul[14]), .B(n23), .Y(out[7]) );
  AOI21X2 U46 ( .A0(n122), .A1(n123), .B0(n121), .Y(n124) );
  AND2X4 U47 ( .A(n116), .B(n113), .Y(n111) );
  NOR2X4 U48 ( .A(in_8bit[4]), .B(in_8bit[0]), .Y(n59) );
  INVX3 U49 ( .A(in_8bit[1]), .Y(n51) );
  NAND2BX4 U50 ( .AN(mul[19]), .B(n112), .Y(n114) );
  XOR2X4 U51 ( .A(n60), .B(n46), .Y(in_8bit_b[5]) );
  NAND2X4 U52 ( .A(n109), .B(n113), .Y(n26) );
  NAND2X2 U53 ( .A(n45), .B(n72), .Y(n31) );
  NAND2X4 U54 ( .A(n18), .B(n17), .Y(n20) );
  INVX4 U55 ( .A(n26), .Y(n18) );
  NAND2X2 U56 ( .A(n26), .B(mul[17]), .Y(n19) );
  XOR2X4 U57 ( .A(mul[10]), .B(n24), .Y(out[3]) );
  NOR2X4 U58 ( .A(in_17bit[1]), .B(in_17bit[0]), .Y(n8) );
  XNOR2X4 U59 ( .A(n9), .B(mul[20]), .Y(out[13]) );
  NAND2X4 U60 ( .A(n120), .B(n113), .Y(n9) );
  NOR2X4 U61 ( .A(n11), .B(n55), .Y(n56) );
  OR2X4 U62 ( .A(n42), .B(n94), .Y(n32) );
  NAND2X2 U63 ( .A(n42), .B(n71), .Y(n72) );
  NAND2X4 U64 ( .A(n59), .B(n58), .Y(n61) );
  OAI21X4 U65 ( .A0(n21), .A1(n61), .B0(n47), .Y(n60) );
  OAI22X4 U66 ( .A0(n45), .A1(in_17bit[1]), .B0(in_17bit[0]), .B1(in_17bit[1]), 
        .Y(n66) );
  NOR2X4 U67 ( .A(in_17bit[3]), .B(n70), .Y(n42) );
  XOR2X4 U68 ( .A(n32), .B(n71), .Y(in_17bit_b[4]) );
  XOR2X4 U69 ( .A(n73), .B(n31), .Y(in_17bit_b[5]) );
  INVX4 U70 ( .A(mul[21]), .Y(n117) );
  XOR2X4 U71 ( .A(n81), .B(n30), .Y(in_17bit_b[9]) );
  XOR2X4 U72 ( .A(n34), .B(n75), .Y(in_17bit_b[6]) );
  NOR3X2 U73 ( .A(mul[20]), .B(n12), .C(n5), .Y(n118) );
  NAND2X4 U74 ( .A(n35), .B(n75), .Y(n76) );
  OR2X4 U75 ( .A(mul[13]), .B(n103), .Y(n104) );
  XNOR2X4 U76 ( .A(mul[21]), .B(n115), .Y(out[14]) );
  XOR2X2 U77 ( .A(mul[9]), .B(n22), .Y(out[2]) );
  XNOR2X2 U78 ( .A(mul[15]), .B(n27), .Y(out[8]) );
  NAND2X2 U79 ( .A(n105), .B(n113), .Y(n27) );
  NAND2XL U80 ( .A(mul[12]), .B(n101), .Y(n15) );
  NAND2X2 U81 ( .A(n13), .B(n14), .Y(n16) );
  NAND2X4 U82 ( .A(n15), .B(n16), .Y(out[5]) );
  INVXL U83 ( .A(mul[12]), .Y(n13) );
  INVX1 U84 ( .A(n101), .Y(n14) );
  NAND2X1 U85 ( .A(n102), .B(n113), .Y(n101) );
  NAND2X4 U86 ( .A(n19), .B(n20), .Y(out[10]) );
  XOR2X4 U87 ( .A(n119), .B(mul[22]), .Y(out[15]) );
  INVX8 U88 ( .A(n51), .Y(n21) );
  XOR2X4 U89 ( .A(n57), .B(in_8bit[4]), .Y(in_8bit_b[4]) );
  NOR2X4 U90 ( .A(n8), .B(n7), .Y(n29) );
  INVXL U91 ( .A(in_17bit[8]), .Y(n79) );
  NOR2X1 U92 ( .A(n90), .B(in_17bit[13]), .Y(n37) );
  NAND2X4 U93 ( .A(n68), .B(n1), .Y(n70) );
  NOR2XL U94 ( .A(n85), .B(in_17bit[11]), .Y(n38) );
  OR2X4 U95 ( .A(n35), .B(n94), .Y(n34) );
  AND2X4 U96 ( .A(n104), .B(n113), .Y(n23) );
  XNOR2X4 U97 ( .A(mul[18]), .B(n28), .Y(out[11]) );
  XNOR2X4 U98 ( .A(n29), .B(n68), .Y(in_17bit_b[2]) );
  NAND2X2 U99 ( .A(n37), .B(n93), .Y(n95) );
  OR2X4 U100 ( .A(mul[8]), .B(out[0]), .Y(n97) );
  NAND2X4 U101 ( .A(n110), .B(n113), .Y(n28) );
  OR2X4 U102 ( .A(mul[16]), .B(n108), .Y(n109) );
  AND2X1 U103 ( .A(n98), .B(n113), .Y(n24) );
  NAND2XL U104 ( .A(n100), .B(n113), .Y(n99) );
  AND2X2 U105 ( .A(n97), .B(n113), .Y(n22) );
  INVXL U106 ( .A(in_8bit[1]), .Y(n50) );
  NAND2XL U107 ( .A(n40), .B(n83), .Y(n85) );
  NAND2X4 U108 ( .A(n65), .B(n47), .Y(n64) );
  OR2X4 U109 ( .A(mul[10]), .B(n98), .Y(n100) );
  OR2X4 U110 ( .A(mul[9]), .B(n97), .Y(n98) );
  OR2X4 U111 ( .A(mul[14]), .B(n104), .Y(n105) );
  OR2X4 U112 ( .A(mul[12]), .B(n102), .Y(n103) );
  NAND2XL U113 ( .A(out[0]), .B(n113), .Y(n96) );
  INVX4 U114 ( .A(n121), .Y(n113) );
  NAND2XL U115 ( .A(n45), .B(n80), .Y(n30) );
  AND2X4 U116 ( .A(n78), .B(n77), .Y(n41) );
  AND2X4 U117 ( .A(n74), .B(n73), .Y(n35) );
  NOR2XL U118 ( .A(n80), .B(in_17bit[9]), .Y(n40) );
  OR2X4 U119 ( .A(mul[18]), .B(n110), .Y(n116) );
  OR2X2 U120 ( .A(mul[11]), .B(n100), .Y(n102) );
  XNOR2X1 U121 ( .A(mul[8]), .B(n96), .Y(out[1]) );
  NOR2XL U122 ( .A(mul[20]), .B(n114), .Y(n122) );
  AOI21X2 U123 ( .A0(n56), .A1(n50), .B0(n48), .Y(n57) );
  INVXL U124 ( .A(in_8bit[2]), .Y(n52) );
  XNOR2X2 U125 ( .A(n87), .B(n88), .Y(in_17bit_b[12]) );
  XOR2X2 U126 ( .A(n36), .B(n79), .Y(in_17bit_b[8]) );
  NAND2XL U127 ( .A(n45), .B(n90), .Y(n89) );
  NAND2XL U128 ( .A(n45), .B(n85), .Y(n84) );
  NAND2X2 U129 ( .A(n38), .B(n88), .Y(n90) );
  NAND2X1 U130 ( .A(n41), .B(n79), .Y(n80) );
  XNOR2X2 U131 ( .A(n77), .B(n39), .Y(in_17bit_b[7]) );
  XNOR2X1 U132 ( .A(n45), .B(n47), .Y(n121) );
  NOR3X2 U133 ( .A(in_17bit[15]), .B(n95), .C(n94), .Y(in_17bit_b[16]) );
  XOR2X2 U134 ( .A(in_17bit[15]), .B(n43), .Y(in_17bit_b[15]) );
  AND2X1 U135 ( .A(n45), .B(n95), .Y(n43) );
  INVX1 U136 ( .A(in_17bit[10]), .Y(n83) );
  INVX1 U137 ( .A(in_8bit[6]), .Y(n63) );
  OAI21X4 U138 ( .A0(n114), .A1(mul[20]), .B0(n113), .Y(n115) );
  NOR2XL U139 ( .A(n37), .B(n94), .Y(n92) );
  XOR2X4 U140 ( .A(n53), .B(n52), .Y(in_8bit_b[2]) );
  XOR2X4 U141 ( .A(n64), .B(n63), .Y(in_8bit_b[6]) );
  NOR3X4 U142 ( .A(in_8bit[6]), .B(n2), .C(n48), .Y(in_8bit_b[7]) );
  XNOR2X4 U143 ( .A(in_17bit[3]), .B(n69), .Y(in_17bit_b[3]) );
  CLKINVX3 U144 ( .A(in_17bit[4]), .Y(n71) );
  CLKINVX3 U145 ( .A(in_17bit[5]), .Y(n73) );
  CLKINVX3 U146 ( .A(n72), .Y(n74) );
  CLKINVX3 U147 ( .A(in_17bit[6]), .Y(n75) );
  CLKINVX3 U148 ( .A(in_17bit[7]), .Y(n77) );
  CLKINVX3 U149 ( .A(n76), .Y(n78) );
  XNOR2X4 U150 ( .A(n82), .B(n83), .Y(in_17bit_b[10]) );
  CLKINVX3 U151 ( .A(in_17bit[11]), .Y(n86) );
  XOR2X4 U152 ( .A(n86), .B(n84), .Y(in_17bit_b[11]) );
  CLKINVX3 U153 ( .A(in_17bit[12]), .Y(n88) );
  XOR2X4 U154 ( .A(n91), .B(n89), .Y(in_17bit_b[13]) );
  CLKINVX3 U155 ( .A(in_17bit[14]), .Y(n93) );
  XNOR2X4 U156 ( .A(n92), .B(n93), .Y(in_17bit_b[14]) );
  CLKINVX3 U157 ( .A(n105), .Y(n106) );
  NAND2BX4 U158 ( .AN(mul[15]), .B(n106), .Y(n108) );
  NAND2X4 U159 ( .A(n108), .B(n113), .Y(n107) );
  XNOR2X4 U160 ( .A(mul[16]), .B(n107), .Y(out[9]) );
  NAND2BX4 U161 ( .AN(mul[17]), .B(n4), .Y(n110) );
  XOR2X4 U162 ( .A(n111), .B(n12), .Y(out[12]) );
  NAND2BX4 U163 ( .AN(mul[19]), .B(n112), .Y(n120) );
  XOR2X4 U164 ( .A(mul[23]), .B(n124), .Y(out[16]) );
endmodule


module multi16_0_DW01_add_0 ( A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, 
        A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, 
        B_20_, B_19_, B_18_, B_17_, B_16_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, 
        SUM_17_, SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, 
        SUM_9_, SUM_8_, SUM_7_, SUM_6_, SUM_5_ );
  input A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_,
         A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, B_20_, B_19_,
         B_18_, B_17_, B_16_;
  output SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, SUM_15_,
         SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, SUM_7_,
         SUM_6_, SUM_5_;
  wire   n1, n2, n3, n4, n5, n6, n8, n9, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46;

  NAND2X2 U2 ( .A(B_18_), .B(A_18_), .Y(n41) );
  CLKINVX8 U3 ( .A(n42), .Y(n27) );
  XOR2X4 U4 ( .A(n46), .B(n1), .Y(n21) );
  AND2X4 U5 ( .A(n41), .B(n23), .Y(n1) );
  INVX4 U6 ( .A(A_15_), .Y(n28) );
  BUFX8 U7 ( .A(A_6_), .Y(SUM_6_) );
  INVX3 U8 ( .A(n25), .Y(n2) );
  INVX4 U9 ( .A(n31), .Y(n4) );
  BUFX12 U10 ( .A(A_14_), .Y(SUM_14_) );
  INVX8 U11 ( .A(n28), .Y(SUM_15_) );
  BUFX12 U12 ( .A(A_11_), .Y(SUM_11_) );
  OAI21X1 U13 ( .A0(n38), .A1(n42), .B0(n2), .Y(n40) );
  NAND2X4 U14 ( .A(n3), .B(n4), .Y(n6) );
  BUFX8 U15 ( .A(A_7_), .Y(SUM_7_) );
  INVX4 U16 ( .A(n38), .Y(n26) );
  OAI21X2 U17 ( .A0(n46), .A1(n39), .B0(n41), .Y(n44) );
  AOI21X2 U18 ( .A0(n23), .A1(n40), .B0(n24), .Y(n35) );
  AOI21X2 U19 ( .A0(n31), .A1(n32), .B0(n22), .Y(n30) );
  INVX8 U20 ( .A(n21), .Y(SUM_18_) );
  OR2X4 U21 ( .A(B_20_), .B(A_20_), .Y(n32) );
  NAND2X2 U22 ( .A(n33), .B(n32), .Y(n34) );
  NAND2X4 U23 ( .A(B_20_), .B(A_20_), .Y(n33) );
  OAI21X4 U24 ( .A0(n35), .A1(n36), .B0(n37), .Y(n31) );
  NOR2BX4 U25 ( .AN(n37), .B(n36), .Y(n45) );
  NAND2X2 U26 ( .A(B_19_), .B(A_19_), .Y(n37) );
  XOR2X4 U27 ( .A(n44), .B(n45), .Y(SUM_19_) );
  NAND2X2 U28 ( .A(n34), .B(n31), .Y(n5) );
  NAND2X4 U29 ( .A(n5), .B(n6), .Y(SUM_20_) );
  CLKINVX3 U30 ( .A(n34), .Y(n3) );
  INVX8 U31 ( .A(n43), .Y(n25) );
  NOR2X2 U32 ( .A(B_19_), .B(A_19_), .Y(n36) );
  AND2X4 U33 ( .A(n9), .B(n42), .Y(SUM_16_) );
  OR2X4 U34 ( .A(A_16_), .B(B_16_), .Y(n9) );
  XOR2X4 U35 ( .A(n8), .B(n27), .Y(SUM_17_) );
  NOR2X4 U36 ( .A(n25), .B(n38), .Y(n8) );
  NAND2X4 U37 ( .A(A_17_), .B(B_17_), .Y(n43) );
  INVX2 U38 ( .A(n41), .Y(n24) );
  INVXL U39 ( .A(n33), .Y(n22) );
  BUFX4 U40 ( .A(A_9_), .Y(SUM_9_) );
  BUFX8 U41 ( .A(A_12_), .Y(SUM_12_) );
  BUFX4 U42 ( .A(A_10_), .Y(SUM_10_) );
  BUFX8 U43 ( .A(A_5_), .Y(SUM_5_) );
  BUFX4 U44 ( .A(A_8_), .Y(SUM_8_) );
  BUFX8 U45 ( .A(A_13_), .Y(SUM_13_) );
  AOI21X4 U46 ( .A0(n26), .A1(n27), .B0(n25), .Y(n46) );
  INVX4 U47 ( .A(n39), .Y(n23) );
  NOR2X4 U48 ( .A(A_18_), .B(B_18_), .Y(n39) );
  NAND2X4 U49 ( .A(A_16_), .B(B_16_), .Y(n42) );
  NOR2X4 U50 ( .A(A_17_), .B(B_17_), .Y(n38) );
  XOR2X1 U51 ( .A(n29), .B(n30), .Y(SUM_21_) );
  XNOR2X1 U52 ( .A(B_21_), .B(A_21_), .Y(n29) );
endmodule


module multi16_0_DW02_mult_0 ( A, B, PRODUCT_23_, PRODUCT_22_, PRODUCT_21_, 
        PRODUCT_20_, PRODUCT_19_, PRODUCT_18_, PRODUCT_17_, PRODUCT_16_, 
        PRODUCT_15_, PRODUCT_14_, PRODUCT_13_, PRODUCT_12_, PRODUCT_11_, 
        PRODUCT_10_, PRODUCT_9_, PRODUCT_8_, PRODUCT_7_ );
  input [16:0] A;
  input [7:0] B;
  output PRODUCT_23_, PRODUCT_22_, PRODUCT_21_, PRODUCT_20_, PRODUCT_19_,
         PRODUCT_18_, PRODUCT_17_, PRODUCT_16_, PRODUCT_15_, PRODUCT_14_,
         PRODUCT_13_, PRODUCT_12_, PRODUCT_11_, PRODUCT_10_, PRODUCT_9_,
         PRODUCT_8_, PRODUCT_7_;
  wire   ab_16__7_, ab_16__6_, ab_16__5_, ab_16__4_, ab_16__3_, ab_16__2_,
         ab_16__1_, ab_16__0_, ab_15__7_, ab_15__6_, ab_15__5_, ab_15__4_,
         ab_15__3_, ab_15__2_, ab_15__1_, ab_15__0_, ab_14__7_, ab_14__6_,
         ab_14__5_, ab_14__4_, ab_14__3_, ab_14__2_, ab_14__1_, ab_14__0_,
         ab_13__7_, ab_13__6_, ab_13__5_, ab_13__4_, ab_13__3_, ab_13__2_,
         ab_13__1_, ab_13__0_, ab_12__7_, ab_12__6_, ab_12__5_, ab_12__4_,
         ab_12__3_, ab_12__2_, ab_12__1_, ab_12__0_, ab_11__7_, ab_11__6_,
         ab_11__5_, ab_11__4_, ab_11__3_, ab_11__2_, ab_11__1_, ab_11__0_,
         ab_10__7_, ab_10__6_, ab_10__5_, ab_10__4_, ab_10__3_, ab_10__2_,
         ab_10__1_, ab_10__0_, ab_9__7_, ab_9__6_, ab_9__5_, ab_9__4_,
         ab_9__3_, ab_9__2_, ab_9__1_, ab_9__0_, ab_8__7_, ab_8__6_, ab_8__5_,
         ab_8__4_, ab_8__3_, ab_8__2_, ab_8__1_, ab_8__0_, ab_7__7_, ab_7__6_,
         ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_, ab_7__0_, ab_6__7_,
         ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_, ab_6__1_, ab_6__0_,
         ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_, ab_5__2_, ab_5__1_,
         ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_, ab_4__3_, ab_4__2_,
         ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_, ab_3__4_, ab_3__3_,
         ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_, ab_2__5_, ab_2__4_,
         ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_, ab_1__6_, ab_1__5_,
         ab_1__4_, ab_1__3_, ab_1__2_, ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_,
         ab_0__3_, ab_0__2_, CARRYB_16__6_, CARRYB_16__5_, CARRYB_16__4_,
         CARRYB_16__3_, CARRYB_16__2_, CARRYB_16__1_, CARRYB_16__0_,
         CARRYB_15__6_, CARRYB_15__5_, CARRYB_15__4_, CARRYB_15__3_,
         CARRYB_15__2_, CARRYB_15__1_, CARRYB_15__0_, CARRYB_14__6_,
         CARRYB_14__5_, CARRYB_14__4_, CARRYB_14__3_, CARRYB_14__2_,
         CARRYB_14__1_, CARRYB_14__0_, CARRYB_13__6_, CARRYB_13__5_,
         CARRYB_13__4_, CARRYB_13__3_, CARRYB_13__2_, CARRYB_13__1_,
         CARRYB_13__0_, CARRYB_12__6_, CARRYB_12__5_, CARRYB_12__4_,
         CARRYB_12__3_, CARRYB_12__2_, CARRYB_12__1_, CARRYB_12__0_,
         CARRYB_11__6_, CARRYB_11__5_, CARRYB_11__4_, CARRYB_11__3_,
         CARRYB_11__2_, CARRYB_11__1_, CARRYB_11__0_, CARRYB_10__6_,
         CARRYB_10__5_, CARRYB_10__4_, CARRYB_10__3_, CARRYB_10__2_,
         CARRYB_10__1_, CARRYB_10__0_, CARRYB_9__6_, CARRYB_9__5_,
         CARRYB_9__4_, CARRYB_9__3_, CARRYB_9__2_, CARRYB_9__1_, CARRYB_9__0_,
         CARRYB_8__6_, CARRYB_8__5_, CARRYB_8__4_, CARRYB_8__3_, CARRYB_8__2_,
         CARRYB_8__1_, CARRYB_8__0_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_,
         CARRYB_7__3_, CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_,
         CARRYB_6__5_, CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_,
         CARRYB_6__0_, CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_,
         CARRYB_5__2_, CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_,
         CARRYB_4__4_, CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_,
         CARRYB_3__6_, CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_,
         CARRYB_3__1_, CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_,
         CARRYB_2__3_, CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__2_,
         CARRYB_1__0_, SUMB_16__6_, SUMB_16__5_, SUMB_16__4_, SUMB_16__3_,
         SUMB_16__2_, SUMB_16__1_, SUMB_16__0_, SUMB_15__6_, SUMB_15__5_,
         SUMB_15__4_, SUMB_15__3_, SUMB_15__2_, SUMB_15__1_, SUMB_14__6_,
         SUMB_14__5_, SUMB_14__4_, SUMB_14__3_, SUMB_14__2_, SUMB_14__1_,
         SUMB_13__6_, SUMB_13__5_, SUMB_13__4_, SUMB_13__3_, SUMB_13__2_,
         SUMB_13__1_, SUMB_12__6_, SUMB_12__5_, SUMB_12__4_, SUMB_12__3_,
         SUMB_12__2_, SUMB_12__1_, SUMB_11__6_, SUMB_11__5_, SUMB_11__4_,
         SUMB_11__3_, SUMB_11__2_, SUMB_11__1_, SUMB_10__6_, SUMB_10__5_,
         SUMB_10__4_, SUMB_10__3_, SUMB_10__2_, SUMB_10__1_, SUMB_9__6_,
         SUMB_9__5_, SUMB_9__4_, SUMB_9__3_, SUMB_9__2_, SUMB_9__1_,
         SUMB_8__6_, SUMB_8__5_, SUMB_8__4_, SUMB_8__3_, SUMB_8__2_,
         SUMB_8__1_, SUMB_7__6_, SUMB_7__5_, SUMB_7__4_, SUMB_7__3_,
         SUMB_7__2_, SUMB_7__1_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_,
         SUMB_6__3_, SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_,
         SUMB_5__4_, SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_,
         SUMB_4__5_, SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_,
         SUMB_3__6_, SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_,
         SUMB_3__1_, SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_,
         SUMB_2__2_, SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_,
         SUMB_1__3_, SUMB_1__2_, SUMB_1__1_, PROD1_7_, A1_21_, A1_20_, A1_19_,
         A1_18_, A1_17_, A1_16_, A1_15_, A1_13_, A1_12_, A1_11_, A1_10_, A1_9_,
         A1_8_, A1_7_, A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, n3, n5, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41;

  ADDFHX2 S4_5 ( .A(ab_16__5_), .B(CARRYB_15__5_), .CI(SUMB_15__6_), .CO(
        CARRYB_16__5_), .S(SUMB_16__5_) );
  multi16_0_DW01_add_0 FS_1 ( .A_21_(A1_21_), .A_20_(A1_20_), .A_19_(A1_19_), 
        .A_18_(A1_18_), .A_17_(A1_17_), .A_16_(A1_16_), .A_15_(A1_15_), 
        .A_14_(SUMB_16__0_), .A_13_(A1_13_), .A_12_(A1_12_), .A_11_(A1_11_), 
        .A_10_(A1_10_), .A_9_(A1_9_), .A_8_(A1_8_), .A_7_(A1_7_), .A_6_(A1_6_), 
        .A_5_(PROD1_7_), .B_21_(n17), .B_20_(n16), .B_19_(n14), .B_18_(n13), 
        .B_17_(n15), .B_16_(n5), .SUM_21_(PRODUCT_23_), .SUM_20_(PRODUCT_22_), 
        .SUM_19_(PRODUCT_21_), .SUM_18_(PRODUCT_20_), .SUM_17_(PRODUCT_19_), 
        .SUM_16_(PRODUCT_18_), .SUM_15_(PRODUCT_17_), .SUM_14_(PRODUCT_16_), 
        .SUM_13_(PRODUCT_15_), .SUM_12_(PRODUCT_14_), .SUM_11_(PRODUCT_13_), 
        .SUM_10_(PRODUCT_12_), .SUM_9_(PRODUCT_11_), .SUM_8_(PRODUCT_10_), 
        .SUM_7_(PRODUCT_9_), .SUM_6_(PRODUCT_8_), .SUM_5_(PRODUCT_7_) );
  ADDFHX4 S2_14_1 ( .A(ab_14__1_), .B(CARRYB_13__1_), .CI(SUMB_13__2_), .CO(
        CARRYB_14__1_), .S(SUMB_14__1_) );
  ADDFHX4 S2_13_2 ( .A(ab_13__2_), .B(CARRYB_12__2_), .CI(SUMB_12__3_), .CO(
        CARRYB_13__2_), .S(SUMB_13__2_) );
  ADDFHX4 S2_14_2 ( .A(ab_14__2_), .B(CARRYB_13__2_), .CI(SUMB_13__3_), .CO(
        CARRYB_14__2_), .S(SUMB_14__2_) );
  ADDFHX4 S4_0 ( .A(ab_16__0_), .B(CARRYB_15__0_), .CI(SUMB_15__1_), .CO(
        CARRYB_16__0_), .S(SUMB_16__0_) );
  ADDFHX4 S2_14_4 ( .A(ab_14__4_), .B(CARRYB_13__4_), .CI(SUMB_13__5_), .CO(
        CARRYB_14__4_), .S(SUMB_14__4_) );
  ADDFHX4 S2_11_1 ( .A(ab_11__1_), .B(CARRYB_10__1_), .CI(SUMB_10__2_), .CO(
        CARRYB_11__1_), .S(SUMB_11__1_) );
  ADDFHX4 S4_2 ( .A(ab_16__2_), .B(CARRYB_15__2_), .CI(SUMB_15__3_), .CO(
        CARRYB_16__2_), .S(SUMB_16__2_) );
  ADDFHX4 S1_14_0 ( .A(ab_14__0_), .B(CARRYB_13__0_), .CI(SUMB_13__1_), .CO(
        CARRYB_14__0_), .S(A1_12_) );
  ADDFHX4 S1_15_0 ( .A(ab_15__0_), .B(CARRYB_14__0_), .CI(SUMB_14__1_), .CO(
        CARRYB_15__0_), .S(A1_13_) );
  ADDFHX4 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  ADDFHX4 S1_7_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(PROD1_7_) );
  ADDFHX4 S2_11_2 ( .A(ab_11__2_), .B(CARRYB_10__2_), .CI(SUMB_10__3_), .CO(
        CARRYB_11__2_), .S(SUMB_11__2_) );
  ADDFHX4 S2_12_2 ( .A(ab_12__2_), .B(CARRYB_11__2_), .CI(SUMB_11__3_), .CO(
        CARRYB_12__2_), .S(SUMB_12__2_) );
  ADDFHX4 S2_14_3 ( .A(ab_14__3_), .B(CARRYB_13__3_), .CI(SUMB_13__4_), .CO(
        CARRYB_14__3_), .S(SUMB_14__3_) );
  ADDFHX4 S2_15_2 ( .A(ab_15__2_), .B(CARRYB_14__2_), .CI(SUMB_14__3_), .CO(
        CARRYB_15__2_), .S(SUMB_15__2_) );
  ADDFHX4 S2_12_5 ( .A(ab_12__5_), .B(CARRYB_11__5_), .CI(SUMB_11__6_), .CO(
        CARRYB_12__5_), .S(SUMB_12__5_) );
  ADDFHX4 S2_10_1 ( .A(ab_10__1_), .B(CARRYB_9__1_), .CI(SUMB_9__2_), .CO(
        CARRYB_10__1_), .S(SUMB_10__1_) );
  ADDFHX4 S2_15_1 ( .A(ab_15__1_), .B(CARRYB_14__1_), .CI(SUMB_14__2_), .CO(
        CARRYB_15__1_), .S(SUMB_15__1_) );
  ADDFHX4 S4_1 ( .A(ab_16__1_), .B(CARRYB_15__1_), .CI(SUMB_15__2_), .CO(
        CARRYB_16__1_), .S(SUMB_16__1_) );
  ADDFHX4 S2_13_3 ( .A(ab_13__3_), .B(CARRYB_12__3_), .CI(SUMB_12__4_), .CO(
        CARRYB_13__3_), .S(SUMB_13__3_) );
  ADDFHX4 S2_11_3 ( .A(ab_11__3_), .B(CARRYB_10__3_), .CI(SUMB_10__4_), .CO(
        CARRYB_11__3_), .S(SUMB_11__3_) );
  ADDFHX4 S2_15_3 ( .A(ab_15__3_), .B(CARRYB_14__3_), .CI(SUMB_14__4_), .CO(
        CARRYB_15__3_), .S(SUMB_15__3_) );
  ADDFHX4 S2_13_4 ( .A(ab_13__4_), .B(CARRYB_12__4_), .CI(SUMB_12__5_), .CO(
        CARRYB_13__4_), .S(SUMB_13__4_) );
  ADDFHX4 S2_11_4 ( .A(ab_11__4_), .B(CARRYB_10__4_), .CI(SUMB_10__5_), .CO(
        CARRYB_11__4_), .S(SUMB_11__4_) );
  ADDFHX4 S2_12_4 ( .A(ab_12__4_), .B(CARRYB_11__4_), .CI(SUMB_11__5_), .CO(
        CARRYB_12__4_), .S(SUMB_12__4_) );
  ADDFHX4 S2_10_2 ( .A(ab_10__2_), .B(CARRYB_9__2_), .CI(SUMB_9__3_), .CO(
        CARRYB_10__2_), .S(SUMB_10__2_) );
  ADDFHX4 S2_12_3 ( .A(ab_12__3_), .B(CARRYB_11__3_), .CI(SUMB_11__4_), .CO(
        CARRYB_12__3_), .S(SUMB_12__3_) );
  ADDFHX4 S1_12_0 ( .A(ab_12__0_), .B(CARRYB_11__0_), .CI(SUMB_11__1_), .CO(
        CARRYB_12__0_), .S(A1_10_) );
  ADDFHX4 S1_13_0 ( .A(ab_13__0_), .B(CARRYB_12__0_), .CI(SUMB_12__1_), .CO(
        CARRYB_13__0_), .S(A1_11_) );
  ADDFHX4 S1_9_0 ( .A(ab_9__0_), .B(CARRYB_8__0_), .CI(SUMB_8__1_), .CO(
        CARRYB_9__0_), .S(A1_7_) );
  ADDFHX4 S1_8_0 ( .A(ab_8__0_), .B(CARRYB_7__0_), .CI(SUMB_7__1_), .CO(
        CARRYB_8__0_), .S(A1_6_) );
  ADDFHX4 S2_11_5 ( .A(ab_11__5_), .B(CARRYB_10__5_), .CI(SUMB_10__6_), .CO(
        CARRYB_11__5_), .S(SUMB_11__5_) );
  ADDFHX1 S3_15_6 ( .A(ab_15__6_), .B(CARRYB_14__6_), .CI(ab_14__7_), .CO(
        CARRYB_15__6_), .S(SUMB_15__6_) );
  ADDFX2 S5_6 ( .A(ab_16__6_), .B(CARRYB_15__6_), .CI(ab_15__7_), .CO(
        CARRYB_16__6_), .S(SUMB_16__6_) );
  ADDFHX4 S2_9_1 ( .A(ab_9__1_), .B(CARRYB_8__1_), .CI(SUMB_8__2_), .CO(
        CARRYB_9__1_), .S(SUMB_9__1_) );
  ADDFHX4 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  ADDFHX4 S4_3 ( .A(ab_16__3_), .B(CARRYB_15__3_), .CI(SUMB_15__4_), .CO(
        CARRYB_16__3_), .S(SUMB_16__3_) );
  ADDFHX4 S3_2_6 ( .A(ab_2__6_), .B(n3), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  ADDFHX4 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  ADDFHX4 S3_9_6 ( .A(ab_9__6_), .B(CARRYB_8__6_), .CI(ab_8__7_), .CO(
        CARRYB_9__6_), .S(SUMB_9__6_) );
  ADDFHX4 S3_10_6 ( .A(ab_10__6_), .B(CARRYB_9__6_), .CI(ab_9__7_), .CO(
        CARRYB_10__6_), .S(SUMB_10__6_) );
  ADDFHX4 S2_9_4 ( .A(ab_9__4_), .B(CARRYB_8__4_), .CI(SUMB_8__5_), .CO(
        CARRYB_9__4_), .S(SUMB_9__4_) );
  ADDFHX4 S2_10_4 ( .A(ab_10__4_), .B(CARRYB_9__4_), .CI(SUMB_9__5_), .CO(
        CARRYB_10__4_), .S(SUMB_10__4_) );
  ADDFHX4 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  ADDFHX4 S2_14_5 ( .A(ab_14__5_), .B(CARRYB_13__5_), .CI(SUMB_13__6_), .CO(
        CARRYB_14__5_), .S(SUMB_14__5_) );
  ADDFHX4 S2_15_5 ( .A(ab_15__5_), .B(CARRYB_14__5_), .CI(SUMB_14__6_), .CO(
        CARRYB_15__5_), .S(SUMB_15__5_) );
  ADDFHX4 S2_9_5 ( .A(ab_9__5_), .B(CARRYB_8__5_), .CI(SUMB_8__6_), .CO(
        CARRYB_9__5_), .S(SUMB_9__5_) );
  ADDFHX4 S2_10_5 ( .A(ab_10__5_), .B(CARRYB_9__5_), .CI(SUMB_9__6_), .CO(
        CARRYB_10__5_), .S(SUMB_10__5_) );
  ADDFHX4 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  ADDFHX4 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  ADDFHX4 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  ADDFHX4 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  ADDFHX4 S3_8_6 ( .A(ab_8__6_), .B(CARRYB_7__6_), .CI(ab_7__7_), .CO(
        CARRYB_8__6_), .S(SUMB_8__6_) );
  ADDFHX4 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  ADDFHX4 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  ADDFHX4 S2_7_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  ADDFHX4 S2_8_5 ( .A(ab_8__5_), .B(CARRYB_7__5_), .CI(SUMB_7__6_), .CO(
        CARRYB_8__5_), .S(SUMB_8__5_) );
  ADDFHX4 S2_13_5 ( .A(ab_13__5_), .B(CARRYB_12__5_), .CI(SUMB_12__6_), .CO(
        CARRYB_13__5_), .S(SUMB_13__5_) );
  ADDFHX4 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  ADDFHX4 S2_10_3 ( .A(ab_10__3_), .B(CARRYB_9__3_), .CI(SUMB_9__4_), .CO(
        CARRYB_10__3_), .S(SUMB_10__3_) );
  ADDFHX4 S2_2_5 ( .A(ab_2__5_), .B(n7), .CI(SUMB_1__6_), .CO(CARRYB_2__5_), 
        .S(SUMB_2__5_) );
  ADDFHX4 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  ADDFHX4 S2_9_2 ( .A(ab_9__2_), .B(CARRYB_8__2_), .CI(SUMB_8__3_), .CO(
        CARRYB_9__2_), .S(SUMB_9__2_) );
  ADDFHX4 S2_12_1 ( .A(ab_12__1_), .B(CARRYB_11__1_), .CI(SUMB_11__2_), .CO(
        CARRYB_12__1_), .S(SUMB_12__1_) );
  ADDFHX4 S2_7_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  ADDFHX4 S2_8_4 ( .A(ab_8__4_), .B(CARRYB_7__4_), .CI(SUMB_7__5_), .CO(
        CARRYB_8__4_), .S(SUMB_8__4_) );
  ADDFHX4 S2_13_1 ( .A(ab_13__1_), .B(CARRYB_12__1_), .CI(SUMB_12__2_), .CO(
        CARRYB_13__1_), .S(SUMB_13__1_) );
  ADDFHX4 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  ADDFHX4 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  ADDFHX4 S3_7_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(
        CARRYB_7__6_), .S(SUMB_7__6_) );
  ADDFHX4 S2_2_1 ( .A(ab_2__1_), .B(n8), .CI(SUMB_1__2_), .CO(CARRYB_2__1_), 
        .S(SUMB_2__1_) );
  ADDFHX4 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  ADDFHX4 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  ADDFHX4 S4_4 ( .A(ab_16__4_), .B(CARRYB_15__4_), .CI(SUMB_15__5_), .CO(
        CARRYB_16__4_), .S(SUMB_16__4_) );
  ADDFHX4 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  ADDFHX4 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  ADDFHX4 S2_7_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  ADDFHX4 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  ADDFHX4 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  ADDFHX4 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  ADDFHX4 S3_13_6 ( .A(ab_13__6_), .B(CARRYB_12__6_), .CI(ab_12__7_), .CO(
        CARRYB_13__6_), .S(SUMB_13__6_) );
  ADDFHX4 S3_14_6 ( .A(ab_14__6_), .B(CARRYB_13__6_), .CI(ab_13__7_), .CO(
        CARRYB_14__6_), .S(SUMB_14__6_) );
  ADDFHX4 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  ADDFHX4 S2_8_3 ( .A(ab_8__3_), .B(CARRYB_7__3_), .CI(SUMB_7__4_), .CO(
        CARRYB_8__3_), .S(SUMB_8__3_) );
  ADDFHX4 S2_9_3 ( .A(ab_9__3_), .B(CARRYB_8__3_), .CI(SUMB_8__4_), .CO(
        CARRYB_9__3_), .S(SUMB_9__3_) );
  ADDFHX4 S2_7_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  ADDFHX4 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  ADDFHX4 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  ADDFHX4 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  ADDFHX4 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  ADDFHX4 S2_7_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  ADDFHX4 S2_8_1 ( .A(ab_8__1_), .B(CARRYB_7__1_), .CI(SUMB_7__2_), .CO(
        CARRYB_8__1_), .S(SUMB_8__1_) );
  ADDFHX4 S3_11_6 ( .A(ab_11__6_), .B(CARRYB_10__6_), .CI(ab_10__7_), .CO(
        CARRYB_11__6_), .S(SUMB_11__6_) );
  ADDFHX4 S3_12_6 ( .A(ab_12__6_), .B(CARRYB_11__6_), .CI(ab_11__7_), .CO(
        CARRYB_12__6_), .S(SUMB_12__6_) );
  ADDFHX4 S1_11_0 ( .A(ab_11__0_), .B(CARRYB_10__0_), .CI(SUMB_10__1_), .CO(
        CARRYB_11__0_), .S(A1_9_) );
  ADDFHX4 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  ADDFHX4 S1_10_0 ( .A(ab_10__0_), .B(CARRYB_9__0_), .CI(SUMB_9__1_), .CO(
        CARRYB_10__0_), .S(A1_8_) );
  ADDFHX4 S2_2_4 ( .A(ab_2__4_), .B(n6), .CI(SUMB_1__5_), .CO(CARRYB_2__4_), 
        .S(SUMB_2__4_) );
  ADDFHX4 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  ADDFHX4 S2_2_3 ( .A(ab_2__3_), .B(n9), .CI(SUMB_1__4_), .CO(CARRYB_2__3_), 
        .S(SUMB_2__3_) );
  ADDFHX4 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  ADDFHX4 S2_8_2 ( .A(ab_8__2_), .B(CARRYB_7__2_), .CI(SUMB_7__3_), .CO(
        CARRYB_8__2_), .S(SUMB_8__2_) );
  ADDFHX4 S1_2_0 ( .A(CARRYB_1__0_), .B(ab_2__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  ADDFHX4 S2_15_4 ( .A(ab_15__4_), .B(CARRYB_14__4_), .CI(SUMB_14__5_), .CO(
        CARRYB_15__4_), .S(SUMB_15__4_) );
  XOR2X2 U2 ( .A(n41), .B(ab_0__2_), .Y(SUMB_1__1_) );
  AND2X2 U3 ( .A(CARRYB_16__2_), .B(SUMB_16__3_), .Y(n13) );
  NOR2BXL U4 ( .AN(A[0]), .B(n30), .Y(n33) );
  INVX12 U5 ( .A(A[0]), .Y(n32) );
  AND2X4 U6 ( .A(ab_0__7_), .B(ab_1__6_), .Y(n3) );
  BUFX20 U7 ( .A(A[2]), .Y(n11) );
  BUFX20 U8 ( .A(A[1]), .Y(n12) );
  NOR2BX1 U9 ( .AN(A[13]), .B(n24), .Y(ab_13__3_) );
  NOR2BX1 U10 ( .AN(A[13]), .B(n22), .Y(ab_13__4_) );
  NOR2BX1 U11 ( .AN(A[9]), .B(n22), .Y(ab_9__4_) );
  NOR2BX2 U12 ( .AN(A[8]), .B(n25), .Y(ab_8__2_) );
  NOR2BX1 U13 ( .AN(A[14]), .B(n24), .Y(ab_14__3_) );
  NOR2BX1 U14 ( .AN(A[14]), .B(n22), .Y(ab_14__4_) );
  INVX1 U15 ( .A(n25), .Y(n10) );
  NOR2BX1 U16 ( .AN(A[12]), .B(n22), .Y(ab_12__4_) );
  NOR2BX1 U17 ( .AN(A[12]), .B(n24), .Y(ab_12__3_) );
  NOR2BX1 U18 ( .AN(A[9]), .B(n26), .Y(ab_9__2_) );
  NOR2BX1 U19 ( .AN(A[12]), .B(n20), .Y(ab_12__5_) );
  NOR2BX1 U20 ( .AN(A[16]), .B(n24), .Y(ab_16__3_) );
  NOR2BX1 U21 ( .AN(A[9]), .B(n20), .Y(ab_9__5_) );
  NOR2BX1 U22 ( .AN(A[10]), .B(n24), .Y(ab_10__3_) );
  NOR2BX1 U23 ( .AN(A[10]), .B(n28), .Y(ab_10__1_) );
  NOR2BX1 U24 ( .AN(A[14]), .B(n20), .Y(ab_14__5_) );
  NOR2BX1 U25 ( .AN(A[16]), .B(n26), .Y(ab_16__2_) );
  NOR2BX1 U26 ( .AN(A[9]), .B(n40), .Y(ab_9__7_) );
  NOR2BX2 U27 ( .AN(A[3]), .B(n30), .Y(ab_3__0_) );
  AND2X4 U29 ( .A(CARRYB_16__0_), .B(SUMB_16__1_), .Y(n5) );
  AND2X4 U30 ( .A(ab_0__5_), .B(ab_1__4_), .Y(n6) );
  AND2X4 U31 ( .A(ab_0__6_), .B(ab_1__5_), .Y(n7) );
  BUFX16 U32 ( .A(n35), .Y(n19) );
  NOR2BX4 U33 ( .AN(B[5]), .B(n32), .Y(ab_0__5_) );
  NOR2BXL U34 ( .AN(A[4]), .B(n30), .Y(ab_4__0_) );
  NOR2BX2 U35 ( .AN(A[3]), .B(n23), .Y(ab_3__3_) );
  NOR2BX2 U36 ( .AN(A[3]), .B(n25), .Y(ab_3__2_) );
  NOR2BX2 U37 ( .AN(A[3]), .B(n27), .Y(ab_3__1_) );
  INVX8 U38 ( .A(n18), .Y(CARRYB_1__2_) );
  AND2X4 U39 ( .A(n41), .B(ab_0__2_), .Y(n8) );
  NOR2BX4 U40 ( .AN(n11), .B(n21), .Y(ab_2__4_) );
  NOR2BX4 U41 ( .AN(n11), .B(n23), .Y(ab_2__3_) );
  NOR2BX4 U42 ( .AN(n11), .B(n29), .Y(ab_2__6_) );
  INVX4 U43 ( .A(B[6]), .Y(n34) );
  NOR2BX4 U44 ( .AN(n11), .B(n30), .Y(ab_2__0_) );
  AND2X4 U45 ( .A(ab_1__3_), .B(ab_0__4_), .Y(n9) );
  NOR2BX4 U46 ( .AN(n11), .B(n27), .Y(ab_2__1_) );
  AND3X2 U47 ( .A(n12), .B(B[1]), .C(n33), .Y(CARRYB_1__0_) );
  AND2X4 U48 ( .A(n12), .B(n10), .Y(ab_1__2_) );
  NOR2BX4 U49 ( .AN(n11), .B(n25), .Y(ab_2__2_) );
  NOR2BX1 U50 ( .AN(n11), .B(n40), .Y(ab_2__7_) );
  NAND2X4 U51 ( .A(ab_1__2_), .B(ab_0__3_), .Y(n18) );
  XOR2X4 U52 ( .A(ab_1__2_), .B(ab_0__3_), .Y(SUMB_1__2_) );
  XOR2X4 U53 ( .A(ab_1__4_), .B(ab_0__5_), .Y(SUMB_1__4_) );
  XOR2X2 U54 ( .A(ab_1__6_), .B(ab_0__7_), .Y(SUMB_1__6_) );
  NOR2BX2 U55 ( .AN(A[4]), .B(n19), .Y(ab_4__5_) );
  NOR2BX1 U56 ( .AN(A[3]), .B(n40), .Y(ab_3__7_) );
  NOR2BX2 U57 ( .AN(A[3]), .B(n29), .Y(ab_3__6_) );
  NOR2BX2 U58 ( .AN(A[4]), .B(n25), .Y(ab_4__2_) );
  NOR2BX2 U59 ( .AN(A[4]), .B(n21), .Y(ab_4__4_) );
  BUFX20 U60 ( .A(n34), .Y(n29) );
  XOR2X4 U61 ( .A(ab_1__3_), .B(ab_0__4_), .Y(SUMB_1__3_) );
  NOR2BX4 U62 ( .AN(B[6]), .B(n32), .Y(ab_0__6_) );
  NOR2BX2 U63 ( .AN(B[4]), .B(n32), .Y(ab_0__4_) );
  NOR2BX2 U64 ( .AN(B[7]), .B(n32), .Y(ab_0__7_) );
  INVX20 U65 ( .A(B[7]), .Y(n40) );
  BUFX20 U66 ( .A(n36), .Y(n21) );
  INVX8 U67 ( .A(B[4]), .Y(n36) );
  NOR2BX2 U68 ( .AN(B[3]), .B(n32), .Y(ab_0__3_) );
  NOR2BX2 U69 ( .AN(A[3]), .B(n21), .Y(ab_3__4_) );
  NOR2BX2 U70 ( .AN(A[4]), .B(n23), .Y(ab_4__3_) );
  NOR2BX2 U71 ( .AN(A[6]), .B(n25), .Y(ab_6__2_) );
  INVX4 U72 ( .A(B[3]), .Y(n37) );
  NOR2BX1 U73 ( .AN(A[5]), .B(n29), .Y(ab_5__6_) );
  NOR2BX4 U74 ( .AN(n12), .B(n27), .Y(n41) );
  NOR2BX4 U75 ( .AN(n12), .B(n23), .Y(ab_1__3_) );
  AND2X4 U76 ( .A(n12), .B(B[6]), .Y(ab_1__6_) );
  CLKINVX8 U77 ( .A(B[0]), .Y(n30) );
  XOR2X4 U78 ( .A(ab_1__5_), .B(ab_0__6_), .Y(SUMB_1__5_) );
  XOR2X4 U79 ( .A(CARRYB_16__5_), .B(SUMB_16__6_), .Y(A1_20_) );
  NOR2BX4 U80 ( .AN(n12), .B(n21), .Y(ab_1__4_) );
  NOR2BX2 U81 ( .AN(A[3]), .B(n19), .Y(ab_3__5_) );
  BUFX12 U82 ( .A(n39), .Y(n27) );
  XOR2X4 U83 ( .A(CARRYB_16__4_), .B(SUMB_16__5_), .Y(A1_19_) );
  NOR2BX4 U84 ( .AN(n12), .B(n19), .Y(ab_1__5_) );
  XOR2X4 U85 ( .A(SUMB_16__1_), .B(CARRYB_16__0_), .Y(A1_15_) );
  NOR2BX2 U86 ( .AN(n11), .B(n19), .Y(ab_2__5_) );
  NOR2BX1 U87 ( .AN(A[14]), .B(n26), .Y(ab_14__2_) );
  AND2X4 U88 ( .A(CARRYB_16__1_), .B(SUMB_16__2_), .Y(n15) );
  NOR2BX1 U89 ( .AN(A[15]), .B(n31), .Y(ab_15__0_) );
  NOR2BX1 U90 ( .AN(A[15]), .B(n26), .Y(ab_15__2_) );
  NOR2BX1 U91 ( .AN(A[9]), .B(n28), .Y(ab_9__1_) );
  NOR2BX1 U92 ( .AN(A[12]), .B(n28), .Y(ab_12__1_) );
  NOR2BX1 U93 ( .AN(A[10]), .B(n30), .Y(ab_10__0_) );
  NOR2BX1 U94 ( .AN(A[6]), .B(n40), .Y(ab_6__7_) );
  NOR2BX2 U95 ( .AN(A[6]), .B(n29), .Y(ab_6__6_) );
  NOR2BX1 U96 ( .AN(A[6]), .B(n23), .Y(ab_6__3_) );
  NOR2BX1 U97 ( .AN(A[6]), .B(n30), .Y(ab_6__0_) );
  NOR2BX1 U98 ( .AN(A[16]), .B(n28), .Y(ab_16__1_) );
  NOR2BX1 U99 ( .AN(A[15]), .B(n22), .Y(ab_15__4_) );
  INVXL U100 ( .A(B[0]), .Y(n31) );
  BUFX8 U101 ( .A(n37), .Y(n23) );
  BUFX1 U102 ( .A(n37), .Y(n24) );
  CLKBUFXL U103 ( .A(n35), .Y(n20) );
  NOR2BX1 U104 ( .AN(A[10]), .B(n22), .Y(ab_10__4_) );
  NOR2BX1 U105 ( .AN(A[10]), .B(n20), .Y(ab_10__5_) );
  NOR2BX1 U106 ( .AN(A[13]), .B(n28), .Y(ab_13__1_) );
  NOR2BX1 U107 ( .AN(A[13]), .B(n20), .Y(ab_13__5_) );
  NOR2BX1 U108 ( .AN(A[4]), .B(n40), .Y(ab_4__7_) );
  NOR2BX1 U109 ( .AN(A[5]), .B(n27), .Y(ab_5__1_) );
  NOR2BXL U110 ( .AN(A[6]), .B(n27), .Y(ab_6__1_) );
  NOR2BXL U111 ( .AN(A[8]), .B(n27), .Y(ab_8__1_) );
  NOR2BXL U112 ( .AN(A[7]), .B(n27), .Y(ab_7__1_) );
  NOR2BX1 U113 ( .AN(A[9]), .B(n24), .Y(ab_9__3_) );
  NOR2BXL U114 ( .AN(A[12]), .B(n29), .Y(ab_12__6_) );
  NOR2BXL U115 ( .AN(A[10]), .B(n29), .Y(ab_10__6_) );
  NOR2BX1 U116 ( .AN(A[5]), .B(n25), .Y(ab_5__2_) );
  NOR2BXL U117 ( .AN(A[5]), .B(n23), .Y(ab_5__3_) );
  NOR2BXL U118 ( .AN(A[8]), .B(n21), .Y(ab_8__4_) );
  NOR2BXL U119 ( .AN(A[8]), .B(n40), .Y(ab_8__7_) );
  NOR2BXL U120 ( .AN(A[9]), .B(n29), .Y(ab_9__6_) );
  NOR2BXL U121 ( .AN(A[8]), .B(n19), .Y(ab_8__5_) );
  NOR2BXL U122 ( .AN(A[7]), .B(n25), .Y(ab_7__2_) );
  NOR2BXL U123 ( .AN(A[7]), .B(n40), .Y(ab_7__7_) );
  NOR2BXL U124 ( .AN(A[8]), .B(n29), .Y(ab_8__6_) );
  NOR2BXL U125 ( .AN(A[7]), .B(n21), .Y(ab_7__4_) );
  NOR2BXL U126 ( .AN(A[7]), .B(n29), .Y(ab_7__6_) );
  NOR2BXL U127 ( .AN(A[7]), .B(n19), .Y(ab_7__5_) );
  NOR2BXL U128 ( .AN(A[8]), .B(n23), .Y(ab_8__3_) );
  NOR2BXL U129 ( .AN(A[7]), .B(n23), .Y(ab_7__3_) );
  NOR2BX1 U130 ( .AN(A[10]), .B(n26), .Y(ab_10__2_) );
  NOR2BX1 U131 ( .AN(A[13]), .B(n26), .Y(ab_13__2_) );
  NOR2BX1 U132 ( .AN(A[12]), .B(n26), .Y(ab_12__2_) );
  NOR2BX1 U133 ( .AN(A[9]), .B(n30), .Y(ab_9__0_) );
  NOR2BXL U134 ( .AN(A[12]), .B(n30), .Y(ab_12__0_) );
  INVX4 U135 ( .A(B[1]), .Y(n39) );
  AND2X1 U136 ( .A(CARRYB_16__5_), .B(SUMB_16__6_), .Y(n17) );
  NOR2BXL U137 ( .AN(A[14]), .B(n40), .Y(ab_14__7_) );
  NOR2BX1 U138 ( .AN(A[15]), .B(n28), .Y(ab_15__1_) );
  NOR2BX1 U139 ( .AN(A[15]), .B(n24), .Y(ab_15__3_) );
  BUFX3 U140 ( .A(n36), .Y(n22) );
  BUFX12 U141 ( .A(n38), .Y(n25) );
  BUFX3 U142 ( .A(n39), .Y(n28) );
  CLKBUFXL U143 ( .A(n38), .Y(n26) );
  NOR2BXL U144 ( .AN(A[11]), .B(n30), .Y(ab_11__0_) );
  AND2X2 U145 ( .A(CARRYB_16__3_), .B(SUMB_16__4_), .Y(n14) );
  NOR2BX2 U146 ( .AN(A[14]), .B(n28), .Y(ab_14__1_) );
  NOR2BX1 U147 ( .AN(A[14]), .B(n31), .Y(ab_14__0_) );
  NOR2BX1 U148 ( .AN(A[13]), .B(n31), .Y(ab_13__0_) );
  NOR2BXL U149 ( .AN(A[7]), .B(n30), .Y(ab_7__0_) );
  NOR2BXL U150 ( .AN(A[11]), .B(n26), .Y(ab_11__2_) );
  NOR2BXL U151 ( .AN(A[11]), .B(n24), .Y(ab_11__3_) );
  NOR2BXL U152 ( .AN(A[11]), .B(n22), .Y(ab_11__4_) );
  NOR2BXL U153 ( .AN(A[8]), .B(n30), .Y(ab_8__0_) );
  NOR2BXL U154 ( .AN(A[11]), .B(n20), .Y(ab_11__5_) );
  NOR2BXL U155 ( .AN(A[11]), .B(n40), .Y(ab_11__7_) );
  NOR2BXL U156 ( .AN(A[10]), .B(n40), .Y(ab_10__7_) );
  NOR2BXL U157 ( .AN(A[11]), .B(n29), .Y(ab_11__6_) );
  NOR2BXL U158 ( .AN(A[5]), .B(n30), .Y(ab_5__0_) );
  NOR2BX1 U159 ( .AN(A[4]), .B(n27), .Y(ab_4__1_) );
  NOR2BXL U160 ( .AN(A[5]), .B(n21), .Y(ab_5__4_) );
  NOR2BXL U161 ( .AN(A[6]), .B(n21), .Y(ab_6__4_) );
  NOR2BXL U162 ( .AN(A[11]), .B(n28), .Y(ab_11__1_) );
  AND2X2 U163 ( .A(CARRYB_16__4_), .B(SUMB_16__5_), .Y(n16) );
  INVX4 U164 ( .A(B[5]), .Y(n35) );
  NOR2BX1 U165 ( .AN(A[12]), .B(n40), .Y(ab_12__7_) );
  NOR2BX1 U166 ( .AN(A[13]), .B(n29), .Y(ab_13__6_) );
  NOR2BXL U167 ( .AN(A[5]), .B(n19), .Y(ab_5__5_) );
  NOR2BXL U168 ( .AN(A[6]), .B(n19), .Y(ab_6__5_) );
  NOR2BXL U169 ( .AN(A[5]), .B(n40), .Y(ab_5__7_) );
  NOR2BX1 U170 ( .AN(A[13]), .B(n40), .Y(ab_13__7_) );
  NOR2BX1 U171 ( .AN(A[14]), .B(n29), .Y(ab_14__6_) );
  XOR2X1 U172 ( .A(CARRYB_16__6_), .B(ab_16__7_), .Y(A1_21_) );
  NOR2BX1 U173 ( .AN(A[16]), .B(n22), .Y(ab_16__4_) );
  NOR2BX1 U174 ( .AN(A[16]), .B(n20), .Y(ab_16__5_) );
  NOR2BXL U175 ( .AN(A[16]), .B(n29), .Y(ab_16__6_) );
  NOR2BXL U176 ( .AN(A[15]), .B(n40), .Y(ab_15__7_) );
  NOR2BX2 U177 ( .AN(B[2]), .B(n32), .Y(ab_0__2_) );
  NOR2BXL U178 ( .AN(A[15]), .B(n29), .Y(ab_15__6_) );
  NOR2BX1 U179 ( .AN(A[16]), .B(n31), .Y(ab_16__0_) );
  NOR2BX1 U180 ( .AN(n12), .B(n40), .Y(ab_1__7_) );
  NOR2BXL U181 ( .AN(A[15]), .B(n20), .Y(ab_15__5_) );
  NOR2BX2 U182 ( .AN(A[4]), .B(n29), .Y(ab_4__6_) );
  NOR2BXL U183 ( .AN(A[16]), .B(n40), .Y(ab_16__7_) );
  XOR2X4 U184 ( .A(SUMB_16__3_), .B(CARRYB_16__2_), .Y(A1_17_) );
  XOR2X4 U185 ( .A(CARRYB_16__3_), .B(SUMB_16__4_), .Y(A1_18_) );
  XOR2X4 U186 ( .A(SUMB_16__2_), .B(CARRYB_16__1_), .Y(A1_16_) );
  INVX8 U187 ( .A(B[2]), .Y(n38) );
endmodule


module multi16_0 ( in_17bit, in_8bit, out );
  input [16:0] in_17bit;
  input [7:0] in_8bit;
  output [16:0] out;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112;
  wire   [16:1] in_17bit_b;
  wire   [7:1] in_8bit_b;
  wire   [23:8] mul;

  multi16_0_DW02_mult_0 mult_55 ( .A({in_17bit_b, in_17bit[0]}), .B({in_8bit_b, 
        n40}), .PRODUCT_23_(mul[23]), .PRODUCT_22_(mul[22]), .PRODUCT_21_(
        mul[21]), .PRODUCT_20_(mul[20]), .PRODUCT_19_(mul[19]), .PRODUCT_18_(
        mul[18]), .PRODUCT_17_(mul[17]), .PRODUCT_16_(mul[16]), .PRODUCT_15_(
        mul[15]), .PRODUCT_14_(mul[14]), .PRODUCT_13_(mul[13]), .PRODUCT_12_(
        mul[12]), .PRODUCT_11_(mul[11]), .PRODUCT_10_(mul[10]), .PRODUCT_9_(
        mul[9]), .PRODUCT_8_(mul[8]), .PRODUCT_7_(out[0]) );
  CLKBUFX4 U2 ( .A(n39), .Y(n1) );
  BUFX12 U3 ( .A(in_17bit[16]), .Y(n39) );
  BUFX20 U4 ( .A(n1), .Y(n9) );
  DLY1X1 U5 ( .A(n101), .Y(n2) );
  NAND3X2 U6 ( .A(in_17bit[1]), .B(n39), .C(in_17bit[0]), .Y(n36) );
  NOR2XL U7 ( .A(n2), .B(mul[19]), .Y(n3) );
  AND2X2 U8 ( .A(n58), .B(n1), .Y(n32) );
  OR2X2 U9 ( .A(n26), .B(n82), .Y(n23) );
  NOR2X1 U10 ( .A(n21), .B(n82), .Y(n20) );
  BUFX8 U11 ( .A(n82), .Y(n5) );
  NAND2X4 U12 ( .A(n105), .B(n6), .Y(n103) );
  INVX8 U13 ( .A(mul[19]), .Y(n105) );
  CLKINVX4 U14 ( .A(n97), .Y(n98) );
  INVXL U15 ( .A(in_17bit[9]), .Y(n69) );
  INVX20 U16 ( .A(n109), .Y(n106) );
  NAND2X2 U17 ( .A(n31), .B(n70), .Y(n71) );
  NAND2X2 U18 ( .A(n81), .B(n80), .Y(n83) );
  BUFX4 U19 ( .A(n6), .Y(n4) );
  XOR2X4 U20 ( .A(n51), .B(in_8bit[5]), .Y(in_8bit_b[5]) );
  INVXL U21 ( .A(mul[20]), .Y(n110) );
  NOR2X2 U22 ( .A(mul[22]), .B(mul[21]), .Y(n111) );
  XNOR2X4 U23 ( .A(n102), .B(n105), .Y(out[12]) );
  NOR2X4 U24 ( .A(n8), .B(n109), .Y(n17) );
  NOR2X4 U25 ( .A(n7), .B(mul[18]), .Y(n6) );
  CLKINVX8 U26 ( .A(in_8bit[2]), .Y(n47) );
  AND2X1 U27 ( .A(n9), .B(n65), .Y(n18) );
  NOR3X2 U28 ( .A(in_17bit[15]), .B(n83), .C(n5), .Y(in_17bit_b[16]) );
  NAND2BX2 U29 ( .AN(mul[17]), .B(n98), .Y(n7) );
  NAND3BX4 U30 ( .AN(mul[20]), .B(n4), .C(n105), .Y(n107) );
  NOR2BX4 U31 ( .AN(n106), .B(n6), .Y(n102) );
  NOR2X4 U32 ( .A(n101), .B(mul[19]), .Y(n8) );
  OR2X4 U33 ( .A(mul[13]), .B(n91), .Y(n92) );
  AOI21X4 U34 ( .A0(n52), .A1(n45), .B0(n43), .Y(n51) );
  CLKINVX8 U35 ( .A(in_8bit[0]), .Y(n41) );
  OR2X4 U36 ( .A(mul[8]), .B(out[0]), .Y(n85) );
  NAND2X4 U37 ( .A(n85), .B(n106), .Y(n12) );
  XNOR2X4 U38 ( .A(mul[9]), .B(n12), .Y(out[2]) );
  NOR3X4 U39 ( .A(in_8bit[6]), .B(n56), .C(n43), .Y(in_8bit_b[7]) );
  INVX1 U40 ( .A(in_8bit[7]), .Y(n44) );
  INVX2 U41 ( .A(in_8bit[7]), .Y(n43) );
  NAND2X2 U42 ( .A(n42), .B(n48), .Y(n16) );
  NOR2X4 U43 ( .A(in_17bit[3]), .B(n58), .Y(n34) );
  NAND2X4 U44 ( .A(n97), .B(n106), .Y(n15) );
  AOI31X4 U45 ( .A0(n111), .A1(n110), .A2(n3), .B0(n109), .Y(n112) );
  NAND2X2 U46 ( .A(n91), .B(n106), .Y(n11) );
  XOR2X4 U47 ( .A(n62), .B(n60), .Y(in_17bit_b[5]) );
  NOR2X4 U48 ( .A(n65), .B(n22), .Y(n21) );
  OR2X4 U49 ( .A(n39), .B(in_17bit[1]), .Y(n38) );
  OR2X4 U50 ( .A(in_17bit[0]), .B(in_17bit[1]), .Y(n37) );
  INVX8 U51 ( .A(n50), .Y(n52) );
  CLKINVX8 U52 ( .A(in_8bit[4]), .Y(n45) );
  NAND2X4 U53 ( .A(n93), .B(n106), .Y(n14) );
  INVX8 U54 ( .A(n39), .Y(n82) );
  XNOR2X4 U55 ( .A(mul[15]), .B(n14), .Y(out[8]) );
  OAI21X4 U56 ( .A0(mul[20]), .A1(n103), .B0(n106), .Y(n104) );
  XOR2X4 U57 ( .A(in_8bit[1]), .B(n25), .Y(in_8bit_b[1]) );
  INVX8 U58 ( .A(n41), .Y(n40) );
  XOR2X2 U59 ( .A(mul[11]), .B(n10), .Y(out[4]) );
  XNOR2X4 U60 ( .A(n104), .B(mul[21]), .Y(out[14]) );
  XNOR2X2 U61 ( .A(mul[13]), .B(n11), .Y(out[6]) );
  XOR2X4 U62 ( .A(n24), .B(n59), .Y(in_17bit_b[4]) );
  OR2X4 U63 ( .A(n34), .B(n82), .Y(n24) );
  XOR2X4 U64 ( .A(n49), .B(n45), .Y(in_8bit_b[4]) );
  NAND2X4 U65 ( .A(n42), .B(n50), .Y(n49) );
  NOR2X4 U66 ( .A(n68), .B(in_17bit[9]), .Y(n31) );
  CLKINVX3 U67 ( .A(n66), .Y(n22) );
  NAND2X2 U68 ( .A(n21), .B(n67), .Y(n68) );
  NOR2X4 U69 ( .A(in_17bit[0]), .B(in_17bit[1]), .Y(n33) );
  XNOR2X2 U70 ( .A(n66), .B(n18), .Y(in_17bit_b[7]) );
  NAND2XL U71 ( .A(n27), .B(n74), .Y(n76) );
  OR2X4 U72 ( .A(mul[10]), .B(n87), .Y(n88) );
  OR2X4 U73 ( .A(mul[16]), .B(n96), .Y(n97) );
  AND2X1 U74 ( .A(n88), .B(n106), .Y(n10) );
  XNOR2X2 U75 ( .A(n20), .B(n67), .Y(in_17bit_b[8]) );
  NAND2BX4 U76 ( .AN(in_17bit[2]), .B(n33), .Y(n58) );
  OR2X4 U77 ( .A(mul[9]), .B(n85), .Y(n87) );
  OR2X4 U78 ( .A(mul[12]), .B(n90), .Y(n91) );
  OR2X4 U79 ( .A(mul[14]), .B(n92), .Y(n93) );
  OR2X4 U80 ( .A(mul[11]), .B(n88), .Y(n90) );
  XOR2X4 U81 ( .A(mul[14]), .B(n13), .Y(out[7]) );
  AND2X4 U82 ( .A(n92), .B(n106), .Y(n13) );
  XNOR2X4 U83 ( .A(n15), .B(mul[17]), .Y(out[10]) );
  XNOR2X1 U84 ( .A(in_8bit[3]), .B(n16), .Y(in_8bit_b[3]) );
  NAND2X2 U85 ( .A(n56), .B(n42), .Y(n55) );
  XOR2X4 U86 ( .A(n17), .B(mul[20]), .Y(out[13]) );
  INVX4 U87 ( .A(n44), .Y(n42) );
  XOR2X4 U88 ( .A(n23), .B(n64), .Y(in_17bit_b[6]) );
  AND2X4 U89 ( .A(n63), .B(n62), .Y(n26) );
  XOR2X2 U90 ( .A(n72), .B(n19), .Y(in_17bit_b[11]) );
  NAND2XL U91 ( .A(n9), .B(n71), .Y(n19) );
  NOR2XL U92 ( .A(n71), .B(n28), .Y(n27) );
  INVXL U93 ( .A(n72), .Y(n28) );
  XOR2X4 U94 ( .A(in_17bit[3]), .B(n32), .Y(in_17bit_b[3]) );
  OR2X4 U95 ( .A(mul[18]), .B(n7), .Y(n101) );
  XNOR2X4 U96 ( .A(n108), .B(mul[22]), .Y(out[15]) );
  XNOR2X1 U97 ( .A(mul[12]), .B(n89), .Y(out[5]) );
  NAND2X1 U98 ( .A(n90), .B(n106), .Y(n89) );
  XNOR2X1 U99 ( .A(mul[8]), .B(n84), .Y(out[1]) );
  NAND2X1 U100 ( .A(out[0]), .B(n106), .Y(n84) );
  XNOR2X2 U101 ( .A(mul[10]), .B(n86), .Y(out[3]) );
  NAND2X2 U102 ( .A(n87), .B(n106), .Y(n86) );
  INVX1 U103 ( .A(in_8bit[6]), .Y(n54) );
  OR2X4 U104 ( .A(in_8bit[3]), .B(n48), .Y(n50) );
  NAND2X2 U105 ( .A(n9), .B(n61), .Y(n60) );
  AND2X4 U106 ( .A(n40), .B(n42), .Y(n25) );
  NOR2XL U107 ( .A(n27), .B(n5), .Y(n73) );
  NAND2XL U108 ( .A(n9), .B(n76), .Y(n75) );
  NAND2BXL U109 ( .AN(n76), .B(n77), .Y(n78) );
  NOR2XL U110 ( .A(n81), .B(n5), .Y(n79) );
  XOR2X2 U111 ( .A(n29), .B(n70), .Y(in_17bit_b[10]) );
  OR2XL U112 ( .A(n31), .B(n5), .Y(n29) );
  XNOR2X2 U113 ( .A(n69), .B(n30), .Y(in_17bit_b[9]) );
  AND2X1 U114 ( .A(n9), .B(n68), .Y(n30) );
  XNOR2X1 U115 ( .A(n9), .B(n42), .Y(n109) );
  XOR2X4 U116 ( .A(n57), .B(in_17bit[2]), .Y(in_17bit_b[2]) );
  XOR2X2 U117 ( .A(in_17bit[15]), .B(n35), .Y(in_17bit_b[15]) );
  AND2X1 U118 ( .A(n9), .B(n83), .Y(n35) );
  OAI21X4 U119 ( .A0(n107), .A1(mul[21]), .B0(n106), .Y(n108) );
  AND3X4 U120 ( .A(n38), .B(n37), .C(n36), .Y(in_17bit_b[1]) );
  NOR2XL U121 ( .A(in_8bit[5]), .B(in_8bit[4]), .Y(n53) );
  OAI21X4 U122 ( .A0(n40), .A1(in_8bit[1]), .B0(n42), .Y(n46) );
  XOR2X4 U123 ( .A(n46), .B(n47), .Y(in_8bit_b[2]) );
  NAND3BX4 U124 ( .AN(in_8bit[1]), .B(n47), .C(n41), .Y(n48) );
  NAND2X4 U125 ( .A(n53), .B(n52), .Y(n56) );
  XOR2X4 U126 ( .A(n55), .B(n54), .Y(in_8bit_b[6]) );
  NOR2X4 U127 ( .A(n33), .B(n82), .Y(n57) );
  CLKINVX3 U128 ( .A(in_17bit[4]), .Y(n59) );
  CLKINVX3 U129 ( .A(in_17bit[5]), .Y(n62) );
  NAND2X4 U130 ( .A(n34), .B(n59), .Y(n61) );
  CLKINVX3 U131 ( .A(n61), .Y(n63) );
  CLKINVX3 U132 ( .A(in_17bit[6]), .Y(n64) );
  CLKINVX3 U133 ( .A(in_17bit[7]), .Y(n66) );
  NAND2X4 U134 ( .A(n26), .B(n64), .Y(n65) );
  CLKINVX3 U135 ( .A(in_17bit[8]), .Y(n67) );
  CLKINVX3 U136 ( .A(in_17bit[10]), .Y(n70) );
  CLKINVX3 U137 ( .A(in_17bit[11]), .Y(n72) );
  CLKINVX3 U138 ( .A(in_17bit[12]), .Y(n74) );
  XNOR2X4 U139 ( .A(n73), .B(n74), .Y(in_17bit_b[12]) );
  CLKINVX3 U140 ( .A(in_17bit[13]), .Y(n77) );
  XOR2X4 U141 ( .A(n77), .B(n75), .Y(in_17bit_b[13]) );
  CLKINVX3 U142 ( .A(n78), .Y(n81) );
  CLKINVX3 U143 ( .A(in_17bit[14]), .Y(n80) );
  XNOR2X4 U144 ( .A(n79), .B(n80), .Y(in_17bit_b[14]) );
  CLKINVX3 U145 ( .A(n93), .Y(n94) );
  NAND2BX4 U146 ( .AN(mul[15]), .B(n94), .Y(n96) );
  NAND2X4 U147 ( .A(n96), .B(n106), .Y(n95) );
  XNOR2X4 U148 ( .A(mul[16]), .B(n95), .Y(out[9]) );
  NAND2BX4 U149 ( .AN(mul[17]), .B(n98), .Y(n100) );
  NAND2X4 U150 ( .A(n100), .B(n106), .Y(n99) );
  XNOR2X4 U151 ( .A(mul[18]), .B(n99), .Y(out[11]) );
  XOR2X4 U152 ( .A(mul[23]), .B(n112), .Y(out[16]) );
endmodule


module butterfly_DW01_sub_25 ( A, B, DIFF );
  input [16:0] A;
  input [16:0] B;
  output [16:0] DIFF;
  wire   n166, n167, n168, n169, n170, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n26,
         n27, n28, n31, n32, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165;

  AND2X1 U3 ( .A(n26), .B(n109), .Y(n107) );
  NAND4BX1 U4 ( .AN(n40), .B(n110), .C(n1), .D(n112), .Y(n101) );
  INVX8 U5 ( .A(n151), .Y(n1) );
  AND3X2 U6 ( .A(n127), .B(n109), .C(n26), .Y(n20) );
  NAND2X1 U7 ( .A(n5), .B(n100), .Y(n97) );
  AOI21X2 U8 ( .A0(n86), .A1(n13), .B0(n88), .Y(n85) );
  NAND2X4 U9 ( .A(n112), .B(n108), .Y(n146) );
  NAND2BX2 U10 ( .AN(A[4]), .B(B[4]), .Y(n59) );
  NAND2BX2 U11 ( .AN(B[4]), .B(A[4]), .Y(n57) );
  CLKINVXL U12 ( .A(B[12]), .Y(n125) );
  AND2X4 U13 ( .A(n1), .B(n139), .Y(n2) );
  AND2X1 U14 ( .A(n5), .B(n104), .Y(n3) );
  INVX4 U15 ( .A(n6), .Y(n138) );
  NAND2X2 U16 ( .A(n142), .B(n143), .Y(n139) );
  INVX4 U17 ( .A(n143), .Y(n149) );
  BUFX4 U18 ( .A(A[10]), .Y(n15) );
  CLKBUFX8 U19 ( .A(n87), .Y(n13) );
  INVX8 U20 ( .A(n111), .Y(n151) );
  CLKINVX3 U21 ( .A(A[9]), .Y(n8) );
  INVX4 U22 ( .A(n161), .Y(n72) );
  NAND2X2 U23 ( .A(n109), .B(n26), .Y(n131) );
  NAND2X2 U24 ( .A(n77), .B(n78), .Y(n74) );
  INVX1 U25 ( .A(n7), .Y(n144) );
  INVX4 U26 ( .A(n120), .Y(n22) );
  NOR2X2 U27 ( .A(n72), .B(n77), .Y(n159) );
  INVX4 U28 ( .A(n123), .Y(n19) );
  INVX8 U29 ( .A(n110), .Y(n37) );
  AND2X2 U30 ( .A(n113), .B(n110), .Y(n10) );
  OR2X4 U31 ( .A(n55), .B(n52), .Y(n31) );
  INVX4 U32 ( .A(n118), .Y(n52) );
  CLKINVX8 U33 ( .A(n99), .Y(n4) );
  INVX8 U34 ( .A(n4), .Y(n5) );
  NAND2X4 U35 ( .A(n2), .B(n112), .Y(n109) );
  NOR2BX2 U36 ( .AN(n84), .B(n85), .Y(n83) );
  NAND3X2 U37 ( .A(n127), .B(n26), .C(n109), .Y(n137) );
  NAND2BX4 U38 ( .AN(B[12]), .B(n16), .Y(n6) );
  NAND2BX2 U39 ( .AN(A[13]), .B(B[13]), .Y(n100) );
  NAND3X4 U40 ( .A(n83), .B(n82), .C(n81), .Y(n79) );
  NOR2X4 U41 ( .A(B[9]), .B(n8), .Y(n7) );
  INVX4 U42 ( .A(A[13]), .Y(n134) );
  NAND3X2 U43 ( .A(n3), .B(n105), .C(n9), .Y(n81) );
  INVX2 U44 ( .A(n101), .Y(n95) );
  OAI21X2 U45 ( .A0(n106), .A1(n101), .B0(n107), .Y(n104) );
  CLKINVX8 U46 ( .A(n88), .Y(n9) );
  INVX4 U47 ( .A(n89), .Y(n88) );
  INVX4 U48 ( .A(n145), .Y(n39) );
  BUFX16 U49 ( .A(n169), .Y(DIFF[8]) );
  XOR2X4 U50 ( .A(n38), .B(n27), .Y(n169) );
  INVX4 U51 ( .A(A[15]), .Y(n17) );
  CLKINVX4 U52 ( .A(n17), .Y(n18) );
  NAND2X2 U53 ( .A(n67), .B(n68), .Y(n62) );
  NAND2BX4 U54 ( .AN(B[3]), .B(A[3]), .Y(n68) );
  AOI21X2 U55 ( .A0(n111), .A1(n148), .B0(n149), .Y(n147) );
  NAND2X2 U56 ( .A(n57), .B(n59), .Y(n61) );
  NAND4X4 U57 ( .A(n112), .B(n10), .C(n1), .D(n38), .Y(n127) );
  BUFX8 U58 ( .A(A[14]), .Y(n11) );
  BUFX16 U59 ( .A(n170), .Y(DIFF[5]) );
  NAND3X1 U60 ( .A(n90), .B(n100), .C(n91), .Y(n86) );
  NAND2X4 U61 ( .A(n6), .B(n126), .Y(n90) );
  OAI2BB1X4 U62 ( .A0N(n16), .A1N(n125), .B0(n93), .Y(n124) );
  XOR2X4 U63 ( .A(n14), .B(n136), .Y(n166) );
  XOR2X4 U64 ( .A(B[13]), .B(A[13]), .Y(n14) );
  AOI21X1 U65 ( .A0(n39), .A1(n110), .B0(n7), .Y(n142) );
  NAND2X4 U66 ( .A(n130), .B(n126), .Y(n128) );
  INVX2 U67 ( .A(n91), .Y(n98) );
  NAND2BX4 U68 ( .AN(B[2]), .B(A[2]), .Y(n70) );
  CLKINVX2 U69 ( .A(n58), .Y(n60) );
  INVX8 U70 ( .A(n135), .Y(n16) );
  INVX8 U71 ( .A(A[12]), .Y(n135) );
  NOR2X4 U72 ( .A(n76), .B(n72), .Y(n75) );
  NAND2BX2 U73 ( .AN(A[1]), .B(B[1]), .Y(n161) );
  XNOR2X4 U74 ( .A(B[16]), .B(A[16]), .Y(n80) );
  NAND2X2 U75 ( .A(n46), .B(n47), .Y(n41) );
  OAI21X2 U76 ( .A0(n135), .A1(B[12]), .B0(n127), .Y(n132) );
  BUFX20 U77 ( .A(n168), .Y(DIFF[10]) );
  NOR2X4 U78 ( .A(n39), .B(n40), .Y(n27) );
  NAND2X2 U79 ( .A(n43), .B(n46), .Y(n154) );
  NAND2BX4 U80 ( .AN(B[13]), .B(A[13]), .Y(n93) );
  BUFX20 U81 ( .A(n166), .Y(DIFF[13]) );
  NAND4X2 U82 ( .A(n94), .B(n95), .C(n9), .D(n96), .Y(n82) );
  BUFX12 U83 ( .A(n108), .Y(n26) );
  NAND2BX4 U84 ( .AN(B[11]), .B(A[11]), .Y(n108) );
  NOR2X2 U85 ( .A(n97), .B(n98), .Y(n96) );
  NAND2BX2 U86 ( .AN(A[8]), .B(B[8]), .Y(n113) );
  AOI2BB1X4 U87 ( .A0N(n20), .A1N(n19), .B0(n124), .Y(n121) );
  NAND2BX4 U88 ( .AN(B[10]), .B(n15), .Y(n143) );
  NOR2BX2 U89 ( .AN(n100), .B(n98), .Y(n105) );
  NAND3X4 U90 ( .A(n127), .B(n109), .C(n26), .Y(n141) );
  NAND2X4 U91 ( .A(n91), .B(n87), .Y(n129) );
  NAND2BX4 U92 ( .AN(B[15]), .B(n18), .Y(n84) );
  NOR2X4 U93 ( .A(n45), .B(n49), .Y(n48) );
  INVX4 U94 ( .A(n50), .Y(n45) );
  XOR2X4 U95 ( .A(n74), .B(n75), .Y(DIFF[1]) );
  NAND2X4 U96 ( .A(n46), .B(n156), .Y(n117) );
  NAND2BX4 U97 ( .AN(A[7]), .B(B[7]), .Y(n46) );
  XOR2X4 U98 ( .A(n148), .B(n150), .Y(n168) );
  AOI21X4 U99 ( .A0(B[13]), .A1(n134), .B0(n19), .Y(n133) );
  NAND2X4 U100 ( .A(n160), .B(n78), .Y(DIFF[0]) );
  NAND3X2 U101 ( .A(n157), .B(n50), .C(n47), .Y(n156) );
  NAND2BX4 U102 ( .AN(B[7]), .B(A[7]), .Y(n47) );
  NAND2BX4 U103 ( .AN(B[8]), .B(A[8]), .Y(n145) );
  OAI2BB1X4 U104 ( .A0N(n134), .A1N(B[13]), .B0(n91), .Y(n122) );
  NAND2BX4 U105 ( .AN(B[14]), .B(n11), .Y(n87) );
  NAND2BX4 U106 ( .AN(A[2]), .B(B[2]), .Y(n64) );
  XOR2X4 U107 ( .A(n62), .B(n63), .Y(DIFF[3]) );
  AOI21X2 U108 ( .A0(n64), .A1(n65), .B0(n66), .Y(n63) );
  INVX8 U109 ( .A(n32), .Y(DIFF[14]) );
  BUFX20 U110 ( .A(n167), .Y(DIFF[12]) );
  NAND2BX4 U111 ( .AN(B[6]), .B(A[6]), .Y(n50) );
  NAND2X2 U112 ( .A(n119), .B(n120), .Y(n23) );
  NAND2X4 U113 ( .A(n21), .B(n22), .Y(n24) );
  NAND2X4 U114 ( .A(n24), .B(n23), .Y(DIFF[15]) );
  INVX4 U115 ( .A(n119), .Y(n21) );
  NAND2BX4 U116 ( .AN(A[12]), .B(B[12]), .Y(n123) );
  NAND3X2 U117 ( .A(n118), .B(n158), .C(n43), .Y(n157) );
  INVX4 U118 ( .A(n43), .Y(n49) );
  AOI21X2 U119 ( .A0(n43), .A1(n44), .B0(n45), .Y(n42) );
  NAND2BX4 U120 ( .AN(A[6]), .B(B[6]), .Y(n43) );
  NAND2BX4 U121 ( .AN(A[10]), .B(B[10]), .Y(n111) );
  NOR2X4 U122 ( .A(n149), .B(n151), .Y(n150) );
  NAND2BX4 U123 ( .AN(A[3]), .B(B[3]), .Y(n67) );
  NAND2BX4 U124 ( .AN(A[5]), .B(B[5]), .Y(n118) );
  NAND2BX2 U125 ( .AN(B[5]), .B(A[5]), .Y(n53) );
  NAND2BX4 U126 ( .AN(A[11]), .B(B[11]), .Y(n112) );
  INVX4 U127 ( .A(n70), .Y(n66) );
  NAND2BX2 U128 ( .AN(B[1]), .B(A[1]), .Y(n73) );
  INVX4 U129 ( .A(n113), .Y(n40) );
  NAND2X4 U130 ( .A(n84), .B(n89), .Y(n120) );
  CLKINVX2 U131 ( .A(n103), .Y(n114) );
  INVXL U132 ( .A(n117), .Y(n116) );
  XOR2X4 U133 ( .A(n146), .B(n147), .Y(DIFF[11]) );
  OAI21X4 U134 ( .A0(n152), .A1(n37), .B0(n144), .Y(n148) );
  XNOR2X4 U135 ( .A(n65), .B(n28), .Y(DIFF[2]) );
  OR2X4 U136 ( .A(n66), .B(n69), .Y(n28) );
  OAI21X4 U137 ( .A0(n71), .A1(n72), .B0(n73), .Y(n65) );
  NAND2BXL U138 ( .AN(B[0]), .B(A[0]), .Y(n78) );
  NAND2BXL U139 ( .AN(A[0]), .B(B[0]), .Y(n160) );
  NAND2BX4 U140 ( .AN(n115), .B(n102), .Y(n58) );
  NAND3XL U141 ( .A(n59), .B(n118), .C(n58), .Y(n155) );
  NAND2X1 U142 ( .A(n53), .B(n57), .Y(n158) );
  XNOR2X4 U143 ( .A(n54), .B(n31), .Y(n170) );
  NAND2X1 U144 ( .A(n162), .B(n68), .Y(n115) );
  NAND3X1 U145 ( .A(n64), .B(n163), .C(n67), .Y(n162) );
  NAND3X1 U146 ( .A(n164), .B(n73), .C(n70), .Y(n163) );
  NAND2X1 U147 ( .A(n165), .B(n161), .Y(n164) );
  INVX1 U148 ( .A(n64), .Y(n69) );
  INVX1 U149 ( .A(n73), .Y(n76) );
  INVX1 U150 ( .A(n74), .Y(n71) );
  INVX1 U151 ( .A(n160), .Y(n77) );
  INVX1 U152 ( .A(n78), .Y(n165) );
  NAND4BXL U153 ( .AN(n52), .B(n59), .C(n43), .D(n46), .Y(n103) );
  NOR2XL U154 ( .A(n102), .B(n103), .Y(n94) );
  XOR2X4 U155 ( .A(n128), .B(n129), .Y(n32) );
  AOI21XL U156 ( .A0(n114), .A1(n115), .B0(n116), .Y(n106) );
  NAND3X4 U157 ( .A(n64), .B(n67), .C(n159), .Y(n102) );
  XOR2X4 U158 ( .A(n35), .B(n36), .Y(DIFF[9]) );
  NOR2X4 U159 ( .A(n7), .B(n37), .Y(n36) );
  XOR2X4 U160 ( .A(n41), .B(n42), .Y(DIFF[7]) );
  XOR2X4 U161 ( .A(n44), .B(n48), .Y(DIFF[6]) );
  OAI21X4 U162 ( .A0(n51), .A1(n52), .B0(n53), .Y(n44) );
  CLKINVX3 U163 ( .A(n54), .Y(n51) );
  CLKINVX3 U164 ( .A(n53), .Y(n55) );
  NAND2X4 U165 ( .A(n56), .B(n57), .Y(n54) );
  NAND2X4 U166 ( .A(n58), .B(n59), .Y(n56) );
  XOR2X4 U167 ( .A(n60), .B(n61), .Y(DIFF[4]) );
  XOR2X4 U168 ( .A(n79), .B(n80), .Y(DIFF[16]) );
  NAND2BX4 U169 ( .AN(A[15]), .B(B[15]), .Y(n89) );
  OAI21X4 U170 ( .A0(n121), .A1(n122), .B0(n13), .Y(n119) );
  NAND2BX4 U171 ( .AN(A[14]), .B(B[14]), .Y(n91) );
  OAI21X4 U172 ( .A0(n132), .A1(n131), .B0(n133), .Y(n130) );
  NAND2BX4 U173 ( .AN(B[13]), .B(A[13]), .Y(n126) );
  AOI21X4 U174 ( .A0(n137), .A1(n5), .B0(n138), .Y(n136) );
  XNOR2X4 U175 ( .A(n140), .B(n141), .Y(n167) );
  NAND2X4 U176 ( .A(n99), .B(n92), .Y(n140) );
  NAND2BX4 U177 ( .AN(B[12]), .B(n16), .Y(n92) );
  NAND2BX4 U178 ( .AN(A[12]), .B(B[12]), .Y(n99) );
  NAND2BX4 U179 ( .AN(A[9]), .B(B[9]), .Y(n110) );
  CLKINVX3 U180 ( .A(n35), .Y(n152) );
  NAND2X4 U181 ( .A(n153), .B(n145), .Y(n35) );
  NAND2X4 U182 ( .A(n38), .B(n113), .Y(n153) );
  OAI21X4 U183 ( .A0(n154), .A1(n155), .B0(n117), .Y(n38) );
endmodule


module butterfly_DW01_add_18 ( A, B, SUM );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  wire   n121, n1, n2, n3, n4, n5, n6, n7, n8, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120;

  XOR2X1 U2 ( .A(n99), .B(n100), .Y(SUM[12]) );
  BUFX8 U3 ( .A(n107), .Y(n1) );
  INVX1 U4 ( .A(n81), .Y(n110) );
  NAND2X2 U5 ( .A(n8), .B(n72), .Y(n105) );
  OAI21X2 U6 ( .A0(B[13]), .A1(A[13]), .B0(n89), .Y(n87) );
  NAND4X2 U7 ( .A(n11), .B(n82), .C(n81), .D(n22), .Y(n102) );
  NAND4BX1 U8 ( .AN(n25), .B(n80), .C(n81), .D(n82), .Y(n70) );
  INVXL U9 ( .A(n117), .Y(n41) );
  INVX8 U10 ( .A(n75), .Y(n117) );
  INVX3 U11 ( .A(n91), .Y(n84) );
  XOR2X2 U12 ( .A(n26), .B(n27), .Y(SUM[7]) );
  BUFX3 U13 ( .A(n121), .Y(SUM[0]) );
  XNOR2X2 U14 ( .A(n105), .B(n106), .Y(n2) );
  NOR2BX2 U15 ( .AN(n24), .B(n25), .Y(n23) );
  INVXL U16 ( .A(n83), .Y(n25) );
  NOR2BX4 U17 ( .AN(n20), .B(n21), .Y(n19) );
  XOR2X2 U18 ( .A(n18), .B(n19), .Y(SUM[9]) );
  XOR2X4 U19 ( .A(n22), .B(n23), .Y(SUM[8]) );
  NOR2BX2 U20 ( .AN(n104), .B(n110), .Y(n109) );
  XOR2X4 U21 ( .A(n109), .B(n1), .Y(SUM[10]) );
  INVX2 U22 ( .A(n33), .Y(n30) );
  XOR2X4 U23 ( .A(n94), .B(n95), .Y(SUM[14]) );
  INVX2 U24 ( .A(n3), .Y(n96) );
  INVX8 U25 ( .A(n80), .Y(n21) );
  NAND2X4 U26 ( .A(B[13]), .B(A[13]), .Y(n86) );
  AND2X4 U27 ( .A(n98), .B(n90), .Y(n3) );
  AOI21X2 U28 ( .A0(n81), .A1(n107), .B0(n108), .Y(n106) );
  NOR2X4 U29 ( .A(A[5]), .B(B[5]), .Y(n15) );
  INVX8 U30 ( .A(n2), .Y(SUM[11]) );
  XOR2X4 U31 ( .A(n33), .B(n34), .Y(SUM[6]) );
  NAND2X2 U32 ( .A(B[11]), .B(A[11]), .Y(n72) );
  NAND3X4 U33 ( .A(n65), .B(n4), .C(n64), .Y(n63) );
  OR2X4 U34 ( .A(B[15]), .B(A[15]), .Y(n4) );
  INVX3 U35 ( .A(n88), .Y(n5) );
  NOR2X4 U36 ( .A(A[14]), .B(B[14]), .Y(n88) );
  NOR2X4 U37 ( .A(A[4]), .B(B[4]), .Y(n16) );
  NAND2X4 U38 ( .A(B[15]), .B(A[15]), .Y(n92) );
  NAND2X4 U39 ( .A(A[9]), .B(B[9]), .Y(n20) );
  OR2X4 U40 ( .A(B[15]), .B(A[15]), .Y(n79) );
  NAND2X4 U41 ( .A(n99), .B(n67), .Y(n98) );
  BUFX8 U42 ( .A(A[8]), .Y(n6) );
  INVX4 U43 ( .A(n67), .Y(n101) );
  XOR2X4 U44 ( .A(n7), .B(n93), .Y(n13) );
  AND2X2 U45 ( .A(n79), .B(n92), .Y(n7) );
  OR2X4 U46 ( .A(A[11]), .B(B[11]), .Y(n8) );
  NAND4BBX2 U47 ( .AN(n15), .BN(n16), .C(n35), .D(n116), .Y(n78) );
  NOR2BX4 U48 ( .AN(n40), .B(n16), .Y(n42) );
  NAND2X2 U49 ( .A(B[12]), .B(A[12]), .Y(n90) );
  AOI21X4 U50 ( .A0(n86), .A1(n87), .B0(n88), .Y(n85) );
  NAND3X4 U51 ( .A(n8), .B(n81), .C(n103), .Y(n73) );
  NAND2X2 U52 ( .A(A[14]), .B(B[14]), .Y(n91) );
  NAND3BX2 U53 ( .AN(n15), .B(n115), .C(n35), .Y(n114) );
  NOR2BX2 U54 ( .AN(n37), .B(n15), .Y(n39) );
  OAI21X2 U55 ( .A0(n36), .A1(n15), .B0(n37), .Y(n33) );
  NOR2X4 U56 ( .A(A[13]), .B(B[13]), .Y(n14) );
  NOR2X4 U57 ( .A(n66), .B(n14), .Y(n65) );
  CLKINVX3 U58 ( .A(n90), .Y(n89) );
  NAND3X4 U59 ( .A(n102), .B(n72), .C(n73), .Y(n99) );
  OAI21X4 U60 ( .A0(n84), .A1(n85), .B0(n79), .Y(n62) );
  OAI21X4 U61 ( .A0(n111), .A1(n21), .B0(n20), .Y(n107) );
  INVX4 U62 ( .A(n18), .Y(n111) );
  NAND2X4 U63 ( .A(n67), .B(n68), .Y(n66) );
  OAI211X2 U64 ( .A0(n21), .A1(n24), .B0(n20), .C0(n104), .Y(n103) );
  INVX8 U65 ( .A(n13), .Y(SUM[15]) );
  INVX8 U66 ( .A(n17), .Y(SUM[16]) );
  NAND2X4 U67 ( .A(B[4]), .B(A[4]), .Y(n40) );
  NAND2X4 U68 ( .A(B[5]), .B(A[5]), .Y(n37) );
  OR2X4 U69 ( .A(A[1]), .B(B[1]), .Y(n54) );
  NAND2X4 U70 ( .A(B[1]), .B(A[1]), .Y(n56) );
  INVX1 U71 ( .A(n92), .Y(n61) );
  AND2X1 U72 ( .A(n83), .B(n80), .Y(n11) );
  NAND2X4 U73 ( .A(n112), .B(n24), .Y(n18) );
  NAND2X4 U74 ( .A(n22), .B(n83), .Y(n112) );
  OAI21X4 U75 ( .A0(n16), .A1(n117), .B0(n40), .Y(n38) );
  AOI21X1 U76 ( .A0(n74), .A1(n75), .B0(n76), .Y(n69) );
  NAND2X1 U77 ( .A(B[7]), .B(A[7]), .Y(n28) );
  NAND2XL U78 ( .A(B[3]), .B(A[3]), .Y(n45) );
  OAI21X4 U79 ( .A0(n117), .A1(n78), .B0(n77), .Y(n22) );
  NAND2BX4 U80 ( .AN(n29), .B(n113), .Y(n77) );
  NAND3X2 U81 ( .A(n114), .B(n32), .C(n28), .Y(n113) );
  AND2X1 U82 ( .A(n73), .B(n72), .Y(n71) );
  NOR2BX1 U83 ( .AN(n50), .B(n49), .Y(n52) );
  OAI2BB1X2 U84 ( .A0N(n54), .A1N(n55), .B0(n56), .Y(n51) );
  OAI21X2 U85 ( .A0(n69), .A1(n70), .B0(n71), .Y(n64) );
  NAND2X4 U86 ( .A(B[10]), .B(A[10]), .Y(n104) );
  OR2X4 U87 ( .A(n6), .B(B[8]), .Y(n83) );
  OR2X4 U88 ( .A(A[3]), .B(B[3]), .Y(n47) );
  OR2X4 U89 ( .A(A[2]), .B(B[2]), .Y(n53) );
  XNOR3X4 U90 ( .A(B[16]), .B(A[16]), .C(n60), .Y(n17) );
  NAND2X4 U91 ( .A(B[0]), .B(A[0]), .Y(n59) );
  NOR2BX1 U92 ( .AN(n59), .B(n12), .Y(n121) );
  NOR2XL U93 ( .A(A[0]), .B(B[0]), .Y(n12) );
  INVX1 U94 ( .A(n51), .Y(n48) );
  INVX1 U95 ( .A(n104), .Y(n108) );
  NAND2X1 U96 ( .A(n37), .B(n40), .Y(n115) );
  NOR2BX1 U97 ( .AN(n32), .B(n31), .Y(n34) );
  NOR2BXL U98 ( .AN(n28), .B(n29), .Y(n27) );
  OAI21XL U99 ( .A0(n30), .A1(n31), .B0(n32), .Y(n26) );
  INVXL U100 ( .A(n35), .Y(n31) );
  INVX1 U101 ( .A(n54), .Y(n58) );
  INVXL U102 ( .A(n78), .Y(n74) );
  INVXL U103 ( .A(n77), .Y(n76) );
  XOR2X1 U104 ( .A(n38), .B(n39), .Y(SUM[5]) );
  XOR2X1 U105 ( .A(n41), .B(n42), .Y(SUM[4]) );
  INVX1 U106 ( .A(n38), .Y(n36) );
  XOR2X1 U107 ( .A(n43), .B(n44), .Y(SUM[3]) );
  NOR2BX1 U108 ( .AN(n45), .B(n46), .Y(n44) );
  OAI21XL U109 ( .A0(n48), .A1(n49), .B0(n50), .Y(n43) );
  INVX1 U110 ( .A(n47), .Y(n46) );
  XOR2X1 U111 ( .A(n55), .B(n57), .Y(SUM[1]) );
  NOR2BX1 U112 ( .AN(n56), .B(n58), .Y(n57) );
  INVX1 U113 ( .A(n53), .Y(n49) );
  XOR2X1 U114 ( .A(n51), .B(n52), .Y(SUM[2]) );
  NAND2X1 U115 ( .A(B[6]), .B(A[6]), .Y(n32) );
  NAND2X2 U116 ( .A(n45), .B(n118), .Y(n75) );
  OAI211X1 U117 ( .A0(n119), .A1(n120), .B0(n53), .C0(n47), .Y(n118) );
  OAI21X1 U118 ( .A0(n58), .A1(n59), .B0(n56), .Y(n119) );
  CLKINVX3 U119 ( .A(n50), .Y(n120) );
  INVX1 U120 ( .A(n59), .Y(n55) );
  NAND3BX4 U121 ( .AN(n61), .B(n63), .C(n62), .Y(n60) );
  AOI21X4 U122 ( .A0(n94), .A1(n5), .B0(n84), .Y(n93) );
  NOR2BX4 U123 ( .AN(n91), .B(n88), .Y(n95) );
  OR2X4 U124 ( .A(B[14]), .B(A[14]), .Y(n68) );
  OAI21X4 U125 ( .A0(n3), .A1(n14), .B0(n86), .Y(n94) );
  XOR2X4 U126 ( .A(n96), .B(n97), .Y(SUM[13]) );
  NOR2BX4 U127 ( .AN(n86), .B(n14), .Y(n97) );
  NOR2BX4 U128 ( .AN(n90), .B(n101), .Y(n100) );
  OR2X4 U129 ( .A(A[12]), .B(B[12]), .Y(n67) );
  OR2X4 U130 ( .A(A[11]), .B(B[11]), .Y(n82) );
  OR2X4 U131 ( .A(A[10]), .B(B[10]), .Y(n81) );
  OR2X4 U132 ( .A(B[9]), .B(A[9]), .Y(n80) );
  NAND2X4 U133 ( .A(B[8]), .B(n6), .Y(n24) );
  CLKINVX3 U134 ( .A(n116), .Y(n29) );
  OR2X4 U135 ( .A(A[7]), .B(B[7]), .Y(n116) );
  OR2X4 U136 ( .A(A[6]), .B(B[6]), .Y(n35) );
  NAND2X4 U137 ( .A(B[2]), .B(A[2]), .Y(n50) );
endmodule


module butterfly_DW01_add_20 ( A, B, SUM );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  wire   n123, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122;

  CLKINVX3 U2 ( .A(n18), .Y(n10) );
  AND2X4 U3 ( .A(n85), .B(n64), .Y(n7) );
  OR2X4 U4 ( .A(A[11]), .B(B[11]), .Y(n1) );
  CLKINVX1 U5 ( .A(n103), .Y(n3) );
  INVX4 U6 ( .A(n90), .Y(n97) );
  INVX2 U7 ( .A(n92), .Y(n113) );
  NOR2BX1 U8 ( .AN(n40), .B(n19), .Y(n42) );
  AND2X2 U9 ( .A(n1), .B(n77), .Y(n2) );
  XNOR2X4 U10 ( .A(n109), .B(n2), .Y(n123) );
  NOR2BX2 U11 ( .AN(n27), .B(n28), .Y(n26) );
  OAI211X2 U12 ( .A0(n121), .A1(n122), .B0(n56), .C0(n50), .Y(n120) );
  OAI21X4 U13 ( .A0(n61), .A1(n62), .B0(n59), .Y(n121) );
  OR2X4 U14 ( .A(A[2]), .B(B[2]), .Y(n56) );
  NOR2BX4 U15 ( .AN(n108), .B(n113), .Y(n112) );
  XOR2X2 U16 ( .A(n21), .B(n22), .Y(SUM[9]) );
  XNOR2X4 U17 ( .A(n3), .B(n104), .Y(SUM[12]) );
  NAND2X4 U18 ( .A(B[11]), .B(A[11]), .Y(n77) );
  XOR2X4 U19 ( .A(n96), .B(n98), .Y(SUM[14]) );
  NAND4BX2 U20 ( .AN(n4), .B(n25), .C(n92), .D(n93), .Y(n106) );
  INVX4 U21 ( .A(n70), .Y(n105) );
  NAND2XL U22 ( .A(n94), .B(n91), .Y(n4) );
  CLKINVX2 U23 ( .A(n71), .Y(n5) );
  INVX2 U24 ( .A(n5), .Y(n6) );
  XNOR2X4 U25 ( .A(n7), .B(n95), .Y(SUM[15]) );
  NAND2X4 U26 ( .A(B[15]), .B(A[15]), .Y(n64) );
  CLKINVX3 U27 ( .A(n89), .Y(n88) );
  NAND2X4 U28 ( .A(n115), .B(n27), .Y(n21) );
  NAND2X4 U29 ( .A(n25), .B(n94), .Y(n115) );
  XOR2X4 U30 ( .A(n8), .B(n9), .Y(SUM[16]) );
  NAND3X4 U31 ( .A(n64), .B(n65), .C(n63), .Y(n8) );
  NOR2X4 U32 ( .A(A[14]), .B(B[14]), .Y(n87) );
  BUFX16 U33 ( .A(n123), .Y(SUM[11]) );
  OAI21X2 U34 ( .A0(n20), .A1(n43), .B0(n44), .Y(n41) );
  INVX4 U35 ( .A(n80), .Y(n43) );
  XOR2X4 U36 ( .A(n36), .B(n37), .Y(SUM[6]) );
  NOR2BX2 U37 ( .AN(n35), .B(n34), .Y(n37) );
  INVX8 U38 ( .A(n91), .Y(n24) );
  NOR2X4 U39 ( .A(n18), .B(n69), .Y(n68) );
  XOR2X4 U40 ( .A(B[16]), .B(A[16]), .Y(n9) );
  OAI21X2 U41 ( .A0(n72), .A1(n73), .B0(n74), .Y(n67) );
  NAND3X4 U42 ( .A(n107), .B(n92), .C(n1), .Y(n78) );
  OAI2BB1X4 U43 ( .A0N(n100), .A1N(n10), .B0(n99), .Y(n96) );
  NOR2X4 U44 ( .A(A[13]), .B(B[13]), .Y(n18) );
  AOI21X2 U45 ( .A0(n99), .A1(n86), .B0(n87), .Y(n84) );
  OAI21X4 U46 ( .A0(n39), .A1(n19), .B0(n40), .Y(n36) );
  NAND3BX2 U47 ( .AN(n19), .B(n118), .C(n38), .Y(n117) );
  NOR2X4 U48 ( .A(A[5]), .B(B[5]), .Y(n19) );
  AOI21X2 U49 ( .A0(n92), .A1(n110), .B0(n111), .Y(n109) );
  NOR2X2 U50 ( .A(A[15]), .B(B[15]), .Y(n66) );
  NAND2X4 U51 ( .A(A[13]), .B(B[13]), .Y(n99) );
  INVX4 U52 ( .A(n21), .Y(n114) );
  NAND2X4 U53 ( .A(A[14]), .B(B[14]), .Y(n90) );
  OAI211X2 U54 ( .A0(n24), .A1(n27), .B0(n23), .C0(n108), .Y(n107) );
  XOR2X4 U55 ( .A(n29), .B(n30), .Y(SUM[7]) );
  OAI21X2 U56 ( .A0(n33), .A1(n34), .B0(n35), .Y(n29) );
  NAND3X4 U57 ( .A(n106), .B(n77), .C(n78), .Y(n103) );
  OAI21X4 U58 ( .A0(n43), .A1(n83), .B0(n82), .Y(n25) );
  NAND2BX4 U59 ( .AN(n32), .B(n116), .Y(n82) );
  XOR2X2 U60 ( .A(n110), .B(n112), .Y(SUM[10]) );
  OAI21X4 U61 ( .A0(n114), .A1(n24), .B0(n23), .Y(n110) );
  NAND2X4 U62 ( .A(n71), .B(n70), .Y(n69) );
  NAND2X4 U63 ( .A(B[9]), .B(A[9]), .Y(n23) );
  OAI21X2 U64 ( .A0(B[13]), .A1(A[13]), .B0(n88), .Y(n86) );
  NAND2X1 U65 ( .A(n12), .B(n100), .Y(n13) );
  NAND2X1 U66 ( .A(n11), .B(n101), .Y(n14) );
  NAND2X4 U67 ( .A(n14), .B(n13), .Y(SUM[13]) );
  INVXL U68 ( .A(n100), .Y(n11) );
  INVX4 U69 ( .A(n101), .Y(n12) );
  NAND2X4 U70 ( .A(n102), .B(n89), .Y(n100) );
  NOR2BX4 U71 ( .AN(n99), .B(n18), .Y(n101) );
  OR2X4 U72 ( .A(n84), .B(n97), .Y(n15) );
  NAND2X4 U73 ( .A(n15), .B(n85), .Y(n63) );
  NAND2X4 U74 ( .A(n103), .B(n70), .Y(n102) );
  NAND2X4 U75 ( .A(B[5]), .B(A[5]), .Y(n40) );
  NAND2X4 U76 ( .A(B[2]), .B(A[2]), .Y(n53) );
  NAND2X4 U77 ( .A(B[4]), .B(A[4]), .Y(n44) );
  NOR2XL U78 ( .A(A[4]), .B(B[4]), .Y(n20) );
  NAND2X4 U79 ( .A(A[8]), .B(B[8]), .Y(n27) );
  OR2X4 U80 ( .A(A[1]), .B(B[1]), .Y(n57) );
  NAND2X4 U81 ( .A(B[1]), .B(A[1]), .Y(n59) );
  OR2X4 U82 ( .A(A[15]), .B(B[15]), .Y(n85) );
  OAI21X1 U83 ( .A0(n51), .A1(n52), .B0(n53), .Y(n46) );
  INVXL U84 ( .A(n50), .Y(n49) );
  NAND2X1 U85 ( .A(B[7]), .B(A[7]), .Y(n31) );
  NAND2XL U86 ( .A(B[3]), .B(A[3]), .Y(n48) );
  INVXL U87 ( .A(n78), .Y(n75) );
  INVXL U88 ( .A(n83), .Y(n79) );
  INVXL U89 ( .A(n82), .Y(n81) );
  INVX2 U90 ( .A(n41), .Y(n39) );
  OAI2BB1X2 U91 ( .A0N(n57), .A1N(n58), .B0(n59), .Y(n54) );
  NAND2X4 U92 ( .A(B[12]), .B(A[12]), .Y(n89) );
  NAND2X4 U93 ( .A(B[10]), .B(A[10]), .Y(n108) );
  OR2X4 U94 ( .A(A[7]), .B(B[7]), .Y(n119) );
  OR2X4 U95 ( .A(B[8]), .B(A[8]), .Y(n94) );
  OR2X4 U96 ( .A(A[3]), .B(B[3]), .Y(n50) );
  NAND2X4 U97 ( .A(B[0]), .B(A[0]), .Y(n62) );
  NOR2BX1 U98 ( .AN(n62), .B(n17), .Y(SUM[0]) );
  NOR2XL U99 ( .A(A[0]), .B(B[0]), .Y(n17) );
  INVX1 U100 ( .A(n54), .Y(n51) );
  AOI21X1 U101 ( .A0(n79), .A1(n80), .B0(n81), .Y(n72) );
  NAND4BXL U102 ( .AN(n28), .B(n91), .C(n92), .D(n93), .Y(n73) );
  NOR2X2 U103 ( .A(n75), .B(n76), .Y(n74) );
  NOR2BXL U104 ( .AN(n23), .B(n24), .Y(n22) );
  INVX1 U105 ( .A(n108), .Y(n111) );
  NAND4BBX2 U106 ( .AN(n19), .BN(n20), .C(n38), .D(n119), .Y(n83) );
  INVX1 U107 ( .A(n94), .Y(n28) );
  NAND3X1 U108 ( .A(n117), .B(n35), .C(n31), .Y(n116) );
  NAND2X1 U109 ( .A(n40), .B(n44), .Y(n118) );
  INVX1 U110 ( .A(n119), .Y(n32) );
  INVX1 U111 ( .A(n77), .Y(n76) );
  INVX1 U112 ( .A(n57), .Y(n61) );
  XOR2X1 U113 ( .A(n25), .B(n26), .Y(SUM[8]) );
  NAND2X2 U114 ( .A(n48), .B(n120), .Y(n80) );
  INVX1 U115 ( .A(n53), .Y(n122) );
  XOR2X1 U116 ( .A(n41), .B(n42), .Y(SUM[5]) );
  INVXL U117 ( .A(n38), .Y(n34) );
  NOR2BXL U118 ( .AN(n31), .B(n32), .Y(n30) );
  INVXL U119 ( .A(n36), .Y(n33) );
  XOR2X1 U120 ( .A(n80), .B(n45), .Y(SUM[4]) );
  NOR2BX1 U121 ( .AN(n44), .B(n20), .Y(n45) );
  INVX1 U122 ( .A(n56), .Y(n52) );
  XOR2X1 U123 ( .A(n54), .B(n55), .Y(SUM[2]) );
  NOR2BX1 U124 ( .AN(n53), .B(n52), .Y(n55) );
  XOR2X1 U125 ( .A(n46), .B(n47), .Y(SUM[3]) );
  NOR2BX1 U126 ( .AN(n48), .B(n49), .Y(n47) );
  XOR2X1 U127 ( .A(n58), .B(n60), .Y(SUM[1]) );
  NOR2BXL U128 ( .AN(n59), .B(n61), .Y(n60) );
  INVX1 U129 ( .A(n62), .Y(n58) );
  NAND2X1 U130 ( .A(B[6]), .B(A[6]), .Y(n35) );
  NAND3BX4 U131 ( .AN(n66), .B(n67), .C(n68), .Y(n65) );
  AOI21X4 U132 ( .A0(n96), .A1(n6), .B0(n97), .Y(n95) );
  NOR2BX4 U133 ( .AN(n90), .B(n87), .Y(n98) );
  OR2X4 U134 ( .A(A[14]), .B(B[14]), .Y(n71) );
  NOR2BX4 U135 ( .AN(n89), .B(n105), .Y(n104) );
  OR2X4 U136 ( .A(A[12]), .B(B[12]), .Y(n70) );
  OR2X4 U137 ( .A(A[11]), .B(B[11]), .Y(n93) );
  OR2X4 U138 ( .A(A[10]), .B(B[10]), .Y(n92) );
  OR2X4 U139 ( .A(A[9]), .B(B[9]), .Y(n91) );
  OR2X4 U140 ( .A(A[6]), .B(B[6]), .Y(n38) );
endmodule


module butterfly_DW01_add_21 ( A, B, SUM );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  wire   n122, n123, n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n13, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121;

  INVX4 U2 ( .A(n91), .Y(n114) );
  OAI2BB1X4 U3 ( .A0N(n22), .A1N(n1), .B0(n24), .Y(n111) );
  CLKINVX20 U4 ( .A(n25), .Y(n1) );
  NAND2X4 U5 ( .A(n115), .B(n28), .Y(n22) );
  OAI21X4 U6 ( .A0(n40), .A1(n19), .B0(n41), .Y(n37) );
  NAND3BX2 U7 ( .AN(n19), .B(n117), .C(n39), .Y(n116) );
  NOR2BX4 U8 ( .AN(n41), .B(n19), .Y(n43) );
  BUFX20 U9 ( .A(n122), .Y(SUM[12]) );
  XOR2X4 U10 ( .A(n101), .B(n100), .Y(SUM[13]) );
  NOR2BX4 U11 ( .AN(n89), .B(n86), .Y(n97) );
  INVX4 U12 ( .A(n89), .Y(n96) );
  INVX8 U13 ( .A(n3), .Y(n91) );
  NOR2X4 U14 ( .A(A[10]), .B(B[10]), .Y(n3) );
  INVX8 U15 ( .A(n100), .Y(n98) );
  BUFX4 U16 ( .A(n103), .Y(n4) );
  CLKINVX2 U17 ( .A(n88), .Y(n87) );
  XOR2X2 U18 ( .A(n111), .B(n113), .Y(SUM[10]) );
  CLKINVX3 U19 ( .A(n11), .Y(SUM[0]) );
  INVX1 U20 ( .A(n123), .Y(n11) );
  NOR2BX1 U21 ( .AN(n32), .B(n33), .Y(n31) );
  INVX4 U22 ( .A(n118), .Y(n33) );
  INVX2 U23 ( .A(n79), .Y(n44) );
  AOI21X4 U24 ( .A0(n91), .A1(n111), .B0(n112), .Y(n110) );
  INVX8 U25 ( .A(n15), .Y(SUM[11]) );
  NAND2X4 U26 ( .A(B[9]), .B(A[9]), .Y(n24) );
  OR2X4 U27 ( .A(A[11]), .B(B[11]), .Y(n5) );
  INVX4 U28 ( .A(n71), .Y(n105) );
  INVX3 U29 ( .A(n86), .Y(n6) );
  NOR2X4 U30 ( .A(A[14]), .B(B[14]), .Y(n86) );
  CLKINVX4 U31 ( .A(n105), .Y(n7) );
  XNOR2X4 U32 ( .A(n8), .B(n94), .Y(SUM[15]) );
  AND2X4 U33 ( .A(n84), .B(n66), .Y(n8) );
  NAND4BX4 U34 ( .AN(n109), .B(n26), .C(n91), .D(n5), .Y(n106) );
  OAI211X2 U35 ( .A0(n120), .A1(n121), .B0(n57), .C0(n51), .Y(n119) );
  INVX4 U36 ( .A(n42), .Y(n40) );
  XOR2X4 U37 ( .A(n30), .B(n31), .Y(SUM[7]) );
  OAI21X2 U38 ( .A0(n34), .A1(n35), .B0(n36), .Y(n30) );
  NAND3X4 U39 ( .A(n69), .B(n9), .C(n68), .Y(n67) );
  OR2X4 U40 ( .A(A[15]), .B(B[15]), .Y(n9) );
  NAND2X1 U41 ( .A(n93), .B(n90), .Y(n109) );
  NAND2X4 U42 ( .A(n7), .B(n72), .Y(n70) );
  NAND2X2 U43 ( .A(B[14]), .B(A[14]), .Y(n89) );
  AOI21X4 U44 ( .A0(n99), .A1(n85), .B0(n86), .Y(n83) );
  NOR2X4 U45 ( .A(n70), .B(n18), .Y(n69) );
  NAND2X2 U46 ( .A(A[11]), .B(B[11]), .Y(n76) );
  NAND3X4 U47 ( .A(n92), .B(n107), .C(n91), .Y(n77) );
  INVX8 U48 ( .A(n90), .Y(n25) );
  NAND2X2 U49 ( .A(B[15]), .B(A[15]), .Y(n66) );
  OAI21X4 U50 ( .A0(n98), .A1(n18), .B0(n99), .Y(n10) );
  NAND3X4 U51 ( .A(n67), .B(n65), .C(n66), .Y(n64) );
  OAI21X4 U52 ( .A0(n96), .A1(n83), .B0(n84), .Y(n65) );
  OAI21X2 U53 ( .A0(B[13]), .A1(A[13]), .B0(n87), .Y(n85) );
  NAND3X4 U54 ( .A(n106), .B(n77), .C(n76), .Y(n103) );
  OAI211X2 U55 ( .A0(n25), .A1(n28), .B0(n24), .C0(n108), .Y(n107) );
  NAND2X4 U56 ( .A(n71), .B(n103), .Y(n102) );
  XOR2X4 U57 ( .A(n16), .B(n110), .Y(n15) );
  XOR2X4 U58 ( .A(n22), .B(n23), .Y(SUM[9]) );
  NOR2X4 U59 ( .A(A[13]), .B(B[13]), .Y(n18) );
  NAND2X4 U60 ( .A(B[13]), .B(A[13]), .Y(n99) );
  XNOR3X4 U61 ( .A(B[16]), .B(A[16]), .C(n64), .Y(n21) );
  NAND4BBX4 U62 ( .AN(n19), .BN(n20), .C(n39), .D(n118), .Y(n82) );
  NOR2X2 U63 ( .A(A[4]), .B(B[4]), .Y(n20) );
  INVX8 U64 ( .A(n21), .Y(SUM[16]) );
  NAND2X4 U65 ( .A(B[4]), .B(A[4]), .Y(n45) );
  NAND2X1 U66 ( .A(B[1]), .B(A[1]), .Y(n60) );
  NAND2X4 U67 ( .A(B[5]), .B(A[5]), .Y(n41) );
  NAND2X4 U68 ( .A(n26), .B(n93), .Y(n115) );
  OAI21X4 U69 ( .A0(n20), .A1(n44), .B0(n45), .Y(n42) );
  OAI2BB1X1 U70 ( .A0N(n58), .A1N(n59), .B0(n60), .Y(n55) );
  NAND2X2 U71 ( .A(B[7]), .B(A[7]), .Y(n32) );
  NAND4BXL U72 ( .AN(n29), .B(n90), .C(n91), .D(n92), .Y(n74) );
  NOR2X4 U73 ( .A(A[5]), .B(B[5]), .Y(n19) );
  NAND2XL U74 ( .A(B[3]), .B(A[3]), .Y(n49) );
  OAI21X4 U75 ( .A0(n44), .A1(n82), .B0(n81), .Y(n26) );
  OAI21X2 U76 ( .A0(n73), .A1(n74), .B0(n75), .Y(n68) );
  OR2X4 U77 ( .A(n33), .B(n13), .Y(n81) );
  AND3X4 U78 ( .A(n116), .B(n36), .C(n32), .Y(n13) );
  AND2X1 U79 ( .A(n5), .B(n76), .Y(n16) );
  NAND2X4 U80 ( .A(B[12]), .B(A[12]), .Y(n88) );
  NAND2X4 U81 ( .A(B[10]), .B(A[10]), .Y(n108) );
  AND2X1 U82 ( .A(n77), .B(n76), .Y(n75) );
  OR2X4 U83 ( .A(A[8]), .B(B[8]), .Y(n93) );
  OR2X4 U84 ( .A(A[3]), .B(B[3]), .Y(n51) );
  OR2X4 U85 ( .A(A[2]), .B(B[2]), .Y(n57) );
  OR2X4 U86 ( .A(A[1]), .B(B[1]), .Y(n58) );
  NAND2X4 U87 ( .A(B[0]), .B(A[0]), .Y(n63) );
  NOR2BX1 U88 ( .AN(n63), .B(n17), .Y(n123) );
  NOR2XL U89 ( .A(A[0]), .B(B[0]), .Y(n17) );
  NOR2BX1 U90 ( .AN(n108), .B(n114), .Y(n113) );
  NOR2BXL U91 ( .AN(n24), .B(n25), .Y(n23) );
  INVX1 U92 ( .A(n93), .Y(n29) );
  NAND2X1 U93 ( .A(n41), .B(n45), .Y(n117) );
  XOR2X1 U94 ( .A(n26), .B(n27), .Y(SUM[8]) );
  NOR2BX1 U95 ( .AN(n28), .B(n29), .Y(n27) );
  XOR2X1 U96 ( .A(n37), .B(n38), .Y(SUM[6]) );
  NOR2BX1 U97 ( .AN(n36), .B(n35), .Y(n38) );
  INVX1 U98 ( .A(n37), .Y(n34) );
  INVXL U99 ( .A(n39), .Y(n35) );
  INVX1 U100 ( .A(n58), .Y(n62) );
  AOI21X1 U101 ( .A0(n78), .A1(n79), .B0(n80), .Y(n73) );
  INVXL U102 ( .A(n82), .Y(n78) );
  INVXL U103 ( .A(n81), .Y(n80) );
  XOR2X1 U104 ( .A(n42), .B(n43), .Y(SUM[5]) );
  XOR2X1 U105 ( .A(n79), .B(n46), .Y(SUM[4]) );
  NOR2BX1 U106 ( .AN(n45), .B(n20), .Y(n46) );
  XOR2X1 U107 ( .A(n59), .B(n61), .Y(SUM[1]) );
  NOR2BX1 U108 ( .AN(n60), .B(n62), .Y(n61) );
  INVX1 U109 ( .A(n57), .Y(n53) );
  XOR2X1 U110 ( .A(n55), .B(n56), .Y(SUM[2]) );
  NOR2BX1 U111 ( .AN(n54), .B(n53), .Y(n56) );
  XOR2X1 U112 ( .A(n47), .B(n48), .Y(SUM[3]) );
  OAI21XL U113 ( .A0(n52), .A1(n53), .B0(n54), .Y(n47) );
  NOR2BX1 U114 ( .AN(n49), .B(n50), .Y(n48) );
  INVX1 U115 ( .A(n55), .Y(n52) );
  INVX1 U116 ( .A(n51), .Y(n50) );
  INVXL U117 ( .A(n108), .Y(n112) );
  NAND2X1 U118 ( .A(B[6]), .B(A[6]), .Y(n36) );
  NAND2X2 U119 ( .A(n49), .B(n119), .Y(n79) );
  OAI21X1 U120 ( .A0(n62), .A1(n63), .B0(n60), .Y(n120) );
  CLKINVX3 U121 ( .A(n54), .Y(n121) );
  INVX1 U122 ( .A(n63), .Y(n59) );
  AOI21X4 U123 ( .A0(n10), .A1(n6), .B0(n96), .Y(n94) );
  OR2X4 U124 ( .A(B[15]), .B(A[15]), .Y(n84) );
  XOR2X4 U125 ( .A(n97), .B(n95), .Y(SUM[14]) );
  OR2X4 U126 ( .A(B[14]), .B(A[14]), .Y(n72) );
  OAI21X4 U127 ( .A0(n98), .A1(n18), .B0(n99), .Y(n95) );
  NOR2BX4 U128 ( .AN(n99), .B(n18), .Y(n101) );
  NAND2X4 U129 ( .A(n102), .B(n88), .Y(n100) );
  XOR2X4 U130 ( .A(n104), .B(n4), .Y(n122) );
  NOR2BX4 U131 ( .AN(n88), .B(n105), .Y(n104) );
  OR2X4 U132 ( .A(B[12]), .B(A[12]), .Y(n71) );
  OR2X4 U133 ( .A(A[11]), .B(B[11]), .Y(n92) );
  OR2X4 U134 ( .A(A[9]), .B(B[9]), .Y(n90) );
  NAND2X4 U135 ( .A(B[8]), .B(A[8]), .Y(n28) );
  OR2X4 U136 ( .A(A[7]), .B(B[7]), .Y(n118) );
  OR2X4 U137 ( .A(A[6]), .B(B[6]), .Y(n39) );
  NAND2X4 U138 ( .A(B[2]), .B(A[2]), .Y(n54) );
endmodule


module butterfly_DW01_sub_26 ( A, B, DIFF );
  input [16:0] A;
  input [16:0] B;
  output [16:0] DIFF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152;

  BUFX4 U3 ( .A(n77), .Y(n1) );
  NAND2BX2 U4 ( .AN(A[11]), .B(n8), .Y(n2) );
  INVX4 U5 ( .A(n9), .Y(n8) );
  NOR2X4 U6 ( .A(n111), .B(n107), .Y(n120) );
  BUFX1 U7 ( .A(B[15]), .Y(n5) );
  INVX2 U8 ( .A(n32), .Y(n38) );
  INVX2 U9 ( .A(n24), .Y(n22) );
  XOR2X2 U10 ( .A(n42), .B(n43), .Y(DIFF[5]) );
  CLKINVX4 U11 ( .A(n42), .Y(n39) );
  NAND2BX2 U12 ( .AN(B[3]), .B(A[3]), .Y(n55) );
  NAND2X2 U13 ( .A(n20), .B(n14), .Y(n15) );
  AOI21X2 U14 ( .A0(n96), .A1(n135), .B0(n136), .Y(n134) );
  INVX8 U15 ( .A(n18), .Y(n136) );
  NAND2X4 U16 ( .A(n110), .B(n92), .Y(n128) );
  NAND2BX4 U17 ( .AN(A[13]), .B(B[13]), .Y(n82) );
  OAI21X2 U18 ( .A0(n23), .A1(n29), .B0(n24), .Y(n130) );
  CLKINVX3 U19 ( .A(n89), .Y(n98) );
  OAI21X2 U20 ( .A0(n71), .A1(n72), .B0(n73), .Y(n69) );
  XOR2X2 U21 ( .A(n52), .B(n56), .Y(DIFF[2]) );
  NAND2X1 U22 ( .A(n35), .B(n36), .Y(n30) );
  INVX3 U23 ( .A(n148), .Y(n60) );
  NOR2X2 U24 ( .A(n64), .B(n60), .Y(n63) );
  INVXL U25 ( .A(n61), .Y(n64) );
  NAND2BX4 U26 ( .AN(B[2]), .B(A[2]), .Y(n58) );
  NAND2BX2 U27 ( .AN(A[2]), .B(B[2]), .Y(n51) );
  NAND2BX2 U28 ( .AN(A[4]), .B(B[4]), .Y(n48) );
  NAND2BX1 U29 ( .AN(B[6]), .B(A[6]), .Y(n145) );
  NOR2X2 U30 ( .A(n34), .B(n38), .Y(n37) );
  NAND2BX1 U31 ( .AN(B[4]), .B(A[4]), .Y(n46) );
  NAND2X4 U32 ( .A(n3), .B(n127), .Y(n126) );
  INVX4 U33 ( .A(n116), .Y(n3) );
  INVX4 U34 ( .A(n97), .Y(n116) );
  INVX8 U35 ( .A(n86), .Y(n85) );
  AND2X4 U36 ( .A(n114), .B(n18), .Y(n4) );
  NOR2X4 U37 ( .A(n4), .B(n116), .Y(n113) );
  INVXL U38 ( .A(A[15]), .Y(n74) );
  BUFX1 U39 ( .A(n70), .Y(n6) );
  AOI21X2 U40 ( .A0(n5), .A1(n74), .B0(n75), .Y(n73) );
  OAI21X2 U41 ( .A0(n123), .A1(n86), .B0(n76), .Y(n122) );
  NAND2X2 U42 ( .A(n82), .B(n76), .Y(n124) );
  INVX4 U43 ( .A(n70), .Y(n101) );
  INVX2 U44 ( .A(n92), .Y(n91) );
  NAND2BX4 U45 ( .AN(n116), .B(n127), .Y(n92) );
  NOR2BX2 U46 ( .AN(B[13]), .B(A[13]), .Y(n123) );
  AOI21X2 U47 ( .A0(n83), .A1(n84), .B0(n85), .Y(n79) );
  NAND2X2 U48 ( .A(n76), .B(n86), .Y(n105) );
  BUFX8 U49 ( .A(n117), .Y(n10) );
  CLKINVX4 U50 ( .A(B[11]), .Y(n9) );
  NAND2BX2 U51 ( .AN(B[7]), .B(A[7]), .Y(n36) );
  INVX4 U52 ( .A(n25), .Y(n140) );
  NAND2BX4 U53 ( .AN(B[8]), .B(A[8]), .Y(n29) );
  INVX2 U54 ( .A(n20), .Y(n139) );
  NAND2BX2 U55 ( .AN(B[14]), .B(A[14]), .Y(n77) );
  NAND2X4 U56 ( .A(n2), .B(n10), .Y(n133) );
  NAND3X4 U57 ( .A(n10), .B(n18), .C(n114), .Y(n127) );
  NAND2BX2 U58 ( .AN(B[10]), .B(A[10]), .Y(n115) );
  XOR2X4 U59 ( .A(n137), .B(n135), .Y(DIFF[10]) );
  NAND2X2 U60 ( .A(n108), .B(n77), .Y(n118) );
  INVX4 U61 ( .A(n108), .Y(n75) );
  XOR2X4 U62 ( .A(n7), .B(n100), .Y(DIFF[15]) );
  NAND2X4 U63 ( .A(n103), .B(n1), .Y(n7) );
  AOI21X4 U64 ( .A0(n121), .A1(n81), .B0(n85), .Y(n125) );
  OAI21X2 U65 ( .A0(n59), .A1(n60), .B0(n61), .Y(n52) );
  INVX2 U66 ( .A(n62), .Y(n59) );
  NAND2X4 U67 ( .A(n69), .B(n6), .Y(n67) );
  NOR2BX2 U68 ( .AN(n36), .B(n34), .Y(n141) );
  NAND2X4 U69 ( .A(n130), .B(n96), .Y(n114) );
  NOR2X4 U70 ( .A(n112), .B(n113), .Y(n109) );
  NAND2X1 U71 ( .A(n81), .B(n82), .Y(n80) );
  AOI21X2 U72 ( .A0(n109), .A1(n110), .B0(n111), .Y(n104) );
  NAND4BX4 U73 ( .AN(n131), .B(n25), .C(n96), .D(n97), .Y(n110) );
  INVX8 U74 ( .A(n132), .Y(n28) );
  NAND2XL U75 ( .A(n132), .B(n95), .Y(n131) );
  NAND2BX4 U76 ( .AN(A[8]), .B(B[8]), .Y(n132) );
  INVX3 U77 ( .A(n145), .Y(n34) );
  INVX8 U78 ( .A(n81), .Y(n111) );
  NOR2X4 U79 ( .A(n85), .B(n111), .Y(n129) );
  NAND2BX4 U80 ( .AN(A[11]), .B(n8), .Y(n97) );
  XOR2X2 U81 ( .A(n33), .B(n37), .Y(DIFF[6]) );
  NAND2X2 U82 ( .A(n9), .B(A[11]), .Y(n117) );
  XOR2X4 U83 ( .A(n133), .B(n134), .Y(DIFF[11]) );
  INVX4 U84 ( .A(n82), .Y(n107) );
  NOR2BX2 U85 ( .AN(B[15]), .B(A[15]), .Y(n102) );
  AOI21X4 U86 ( .A0(n120), .A1(n121), .B0(n122), .Y(n119) );
  XOR2X4 U87 ( .A(n124), .B(n125), .Y(DIFF[13]) );
  XOR2X4 U88 ( .A(n129), .B(n128), .Y(DIFF[12]) );
  NAND2BX4 U89 ( .AN(B[15]), .B(A[15]), .Y(n70) );
  AOI21X2 U90 ( .A0(n78), .A1(n79), .B0(n80), .Y(n71) );
  XOR2X4 U91 ( .A(n67), .B(n68), .Y(DIFF[16]) );
  OAI2BB1X4 U92 ( .A0N(n141), .A1N(n142), .B0(n35), .Y(n93) );
  NAND2BX4 U93 ( .AN(A[7]), .B(B[7]), .Y(n35) );
  NOR2X2 U94 ( .A(n88), .B(n89), .Y(n83) );
  NOR2X4 U95 ( .A(n138), .B(n136), .Y(n137) );
  NAND2BX4 U96 ( .AN(A[14]), .B(B[14]), .Y(n108) );
  NOR2X4 U97 ( .A(n27), .B(n28), .Y(n26) );
  XNOR2X4 U98 ( .A(B[16]), .B(A[16]), .Y(n68) );
  NAND2BX4 U99 ( .AN(B[13]), .B(A[13]), .Y(n76) );
  NAND2X4 U100 ( .A(n110), .B(n126), .Y(n121) );
  OR2X4 U101 ( .A(n104), .B(n105), .Y(n17) );
  NAND2BX4 U102 ( .AN(A[12]), .B(B[12]), .Y(n81) );
  NAND2BX4 U103 ( .AN(B[12]), .B(A[12]), .Y(n86) );
  NAND3X1 U104 ( .A(n51), .B(n150), .C(n54), .Y(n149) );
  NAND2BX4 U105 ( .AN(A[3]), .B(B[3]), .Y(n54) );
  INVX4 U106 ( .A(n144), .Y(n40) );
  NAND2BX4 U107 ( .AN(A[5]), .B(B[5]), .Y(n144) );
  NAND2BX4 U108 ( .AN(B[9]), .B(A[9]), .Y(n24) );
  NOR2X4 U109 ( .A(n75), .B(n107), .Y(n106) );
  OAI21X4 U110 ( .A0(n139), .A1(n23), .B0(n24), .Y(n135) );
  AOI21X2 U111 ( .A0(n32), .A1(n33), .B0(n34), .Y(n31) );
  OAI21X4 U112 ( .A0(n39), .A1(n40), .B0(n41), .Y(n33) );
  XOR2X4 U113 ( .A(n118), .B(n119), .Y(DIFF[14]) );
  NOR2X4 U114 ( .A(n102), .B(n101), .Y(n100) );
  NAND2X2 U115 ( .A(n25), .B(n11), .Y(n12) );
  NAND2X1 U116 ( .A(n140), .B(n26), .Y(n13) );
  NAND2X4 U117 ( .A(n12), .B(n13), .Y(DIFF[8]) );
  INVX2 U118 ( .A(n26), .Y(n11) );
  OAI2BB1X4 U119 ( .A0N(n98), .A1N(n47), .B0(n93), .Y(n25) );
  NAND2X2 U120 ( .A(n139), .B(n21), .Y(n16) );
  NAND2X4 U121 ( .A(n15), .B(n16), .Y(DIFF[9]) );
  INVX4 U122 ( .A(n21), .Y(n14) );
  OAI21X4 U123 ( .A0(n28), .A1(n140), .B0(n29), .Y(n20) );
  NOR2X4 U124 ( .A(n22), .B(n23), .Y(n21) );
  NAND2X4 U125 ( .A(n17), .B(n106), .Y(n103) );
  NAND4BX2 U126 ( .AN(n28), .B(n95), .C(n96), .D(n2), .Y(n88) );
  INVX4 U127 ( .A(n96), .Y(n138) );
  NAND2BX4 U128 ( .AN(A[10]), .B(B[10]), .Y(n96) );
  INVX8 U129 ( .A(n95), .Y(n23) );
  NAND2BX4 U130 ( .AN(A[9]), .B(B[9]), .Y(n95) );
  BUFX8 U131 ( .A(n115), .Y(n18) );
  NAND3X1 U132 ( .A(n51), .B(n54), .C(n146), .Y(n87) );
  NAND2XL U133 ( .A(n152), .B(n148), .Y(n151) );
  NAND3X2 U134 ( .A(n151), .B(n61), .C(n58), .Y(n150) );
  INVXL U135 ( .A(n58), .Y(n53) );
  NAND2XL U136 ( .A(n65), .B(n66), .Y(n62) );
  NAND2XL U137 ( .A(n46), .B(n48), .Y(n19) );
  NAND4BX2 U138 ( .AN(n40), .B(n48), .C(n32), .D(n35), .Y(n89) );
  NOR2X2 U139 ( .A(n60), .B(n65), .Y(n146) );
  NAND2X2 U140 ( .A(n149), .B(n55), .Y(n99) );
  NAND2X2 U141 ( .A(n47), .B(n48), .Y(n45) );
  XNOR2X1 U142 ( .A(n47), .B(n19), .Y(DIFF[4]) );
  INVXL U143 ( .A(n51), .Y(n57) );
  NAND2BX2 U144 ( .AN(A[6]), .B(B[6]), .Y(n32) );
  NAND2BXL U145 ( .AN(B[1]), .B(A[1]), .Y(n61) );
  NAND2BXL U146 ( .AN(A[1]), .B(B[1]), .Y(n148) );
  NAND2BXL U147 ( .AN(B[0]), .B(A[0]), .Y(n66) );
  NAND2BXL U148 ( .AN(A[0]), .B(B[0]), .Y(n147) );
  NAND2BX1 U149 ( .AN(n99), .B(n87), .Y(n47) );
  AOI21X1 U150 ( .A0(n93), .A1(n94), .B0(n88), .Y(n90) );
  NAND2XL U151 ( .A(n98), .B(n99), .Y(n94) );
  INVX1 U152 ( .A(n87), .Y(n84) );
  INVXL U153 ( .A(n10), .Y(n112) );
  INVX1 U154 ( .A(n29), .Y(n27) );
  XOR2X2 U155 ( .A(n30), .B(n31), .Y(DIFF[7]) );
  NOR2XL U156 ( .A(n44), .B(n40), .Y(n43) );
  INVXL U157 ( .A(n41), .Y(n44) );
  NAND3X1 U158 ( .A(n32), .B(n143), .C(n144), .Y(n142) );
  NAND2X1 U159 ( .A(n41), .B(n46), .Y(n143) );
  NAND2X2 U160 ( .A(n45), .B(n46), .Y(n42) );
  NOR2X1 U161 ( .A(n53), .B(n57), .Y(n56) );
  XOR2X1 U162 ( .A(n49), .B(n50), .Y(DIFF[3]) );
  NAND2X1 U163 ( .A(n54), .B(n55), .Y(n49) );
  AOI21XL U164 ( .A0(n51), .A1(n52), .B0(n53), .Y(n50) );
  XOR2X1 U165 ( .A(n62), .B(n63), .Y(DIFF[1]) );
  NOR2X1 U166 ( .A(n90), .B(n91), .Y(n78) );
  NAND2XL U167 ( .A(n76), .B(n77), .Y(n72) );
  INVX1 U168 ( .A(n147), .Y(n65) );
  INVX1 U169 ( .A(n66), .Y(n152) );
  NAND2X1 U170 ( .A(n147), .B(n66), .Y(DIFF[0]) );
  NAND2BX4 U171 ( .AN(B[5]), .B(A[5]), .Y(n41) );
endmodule


module butterfly_DW01_sub_31 ( A, B, DIFF );
  input [16:0] A;
  input [16:0] B;
  output [16:0] DIFF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137;

  NOR2BX4 U3 ( .AN(A[15]), .B(B[15]), .Y(n100) );
  INVX1 U4 ( .A(n73), .Y(n70) );
  OAI21X4 U5 ( .A0(n67), .A1(n68), .B0(n69), .Y(n66) );
  CLKINVX3 U6 ( .A(n75), .Y(n1) );
  CLKINVX4 U7 ( .A(n1), .Y(n2) );
  AOI21X4 U8 ( .A0(n8), .A1(n5), .B0(n104), .Y(n101) );
  CLKINVX4 U9 ( .A(n83), .Y(n5) );
  NAND3X2 U10 ( .A(n106), .B(n14), .C(n88), .Y(n8) );
  OAI2BB1X4 U11 ( .A0N(n31), .A1N(n32), .B0(n33), .Y(n26) );
  INVX2 U12 ( .A(n31), .Y(n36) );
  NAND3X1 U13 ( .A(n31), .B(n130), .C(n131), .Y(n129) );
  NAND2BX2 U14 ( .AN(B[10]), .B(A[10]), .Y(n116) );
  BUFX8 U15 ( .A(n77), .Y(n10) );
  NAND2BX4 U16 ( .AN(A[11]), .B(B[11]), .Y(n119) );
  INVX2 U17 ( .A(n33), .Y(n35) );
  NOR2X2 U18 ( .A(n82), .B(n83), .Y(n78) );
  INVX4 U19 ( .A(n24), .Y(n4) );
  AND3X4 U20 ( .A(n23), .B(n19), .C(n114), .Y(n3) );
  NAND2BXL U21 ( .AN(B[8]), .B(A[8]), .Y(n117) );
  INVX4 U22 ( .A(n40), .Y(n37) );
  NAND2X4 U23 ( .A(n43), .B(n44), .Y(n40) );
  INVX4 U24 ( .A(n117), .Y(n24) );
  XOR2X2 U25 ( .A(n32), .B(n34), .Y(DIFF[6]) );
  NAND2BX2 U26 ( .AN(A[6]), .B(B[6]), .Y(n31) );
  NAND2BX2 U27 ( .AN(B[6]), .B(A[6]), .Y(n33) );
  NAND2BX4 U28 ( .AN(B[4]), .B(A[4]), .Y(n44) );
  NAND2BX4 U29 ( .AN(A[4]), .B(B[4]), .Y(n46) );
  XNOR2X2 U30 ( .A(n23), .B(n15), .Y(DIFF[8]) );
  XOR2X4 U31 ( .A(n11), .B(n8), .Y(DIFF[12]) );
  NAND2BX4 U32 ( .AN(A[11]), .B(B[11]), .Y(n93) );
  BUFX12 U33 ( .A(n89), .Y(n14) );
  CLKINVXL U34 ( .A(B[15]), .Y(n65) );
  OAI21X2 U35 ( .A0(n74), .A1(n2), .B0(n76), .Y(n68) );
  OR2X4 U36 ( .A(A[14]), .B(n103), .Y(n9) );
  NAND4BX4 U37 ( .AN(n38), .B(n46), .C(n31), .D(n30), .Y(n82) );
  NAND2BX4 U38 ( .AN(A[7]), .B(B[7]), .Y(n30) );
  NAND2X2 U39 ( .A(n24), .B(n92), .Y(n115) );
  NAND3X1 U40 ( .A(n94), .B(n95), .C(n96), .Y(n67) );
  NAND2XL U41 ( .A(n97), .B(n77), .Y(n96) );
  XOR2X4 U42 ( .A(n6), .B(n20), .Y(DIFF[9]) );
  NOR2X4 U43 ( .A(n21), .B(n22), .Y(n6) );
  XOR2X4 U44 ( .A(n7), .B(n64), .Y(DIFF[16]) );
  XNOR2X4 U45 ( .A(B[16]), .B(A[16]), .Y(n7) );
  AND2X4 U46 ( .A(n93), .B(n89), .Y(n18) );
  NAND2XL U47 ( .A(n14), .B(n88), .Y(n87) );
  INVX4 U48 ( .A(n20), .Y(n125) );
  AOI21X2 U49 ( .A0(n114), .A1(n122), .B0(n123), .Y(n121) );
  NAND2X4 U50 ( .A(n3), .B(n119), .Y(n106) );
  AND2X2 U51 ( .A(n120), .B(n92), .Y(n19) );
  NAND2X4 U52 ( .A(n9), .B(n10), .Y(n102) );
  INVX8 U53 ( .A(n92), .Y(n22) );
  XOR2X2 U54 ( .A(n40), .B(n41), .Y(DIFF[5]) );
  NOR2X1 U55 ( .A(n42), .B(n38), .Y(n41) );
  NAND2BX4 U56 ( .AN(B[5]), .B(A[5]), .Y(n39) );
  INVX8 U57 ( .A(n72), .Y(n71) );
  NAND3BX2 U58 ( .AN(n21), .B(n115), .C(n116), .Y(n113) );
  NOR2X4 U59 ( .A(n83), .B(n97), .Y(n11) );
  BUFX3 U60 ( .A(n95), .Y(n12) );
  CLKINVX8 U61 ( .A(n103), .Y(n13) );
  INVX8 U62 ( .A(B[14]), .Y(n103) );
  NAND2BX4 U63 ( .AN(A[8]), .B(B[8]), .Y(n120) );
  NAND3X2 U64 ( .A(n10), .B(n78), .C(n79), .Y(n76) );
  NAND2X2 U65 ( .A(n94), .B(n105), .Y(n104) );
  AOI21X2 U66 ( .A0(n110), .A1(n84), .B0(n97), .Y(n112) );
  INVX8 U67 ( .A(n84), .Y(n83) );
  INVX4 U68 ( .A(n23), .Y(n126) );
  NAND2BX4 U69 ( .AN(B[11]), .B(A[11]), .Y(n89) );
  OAI2BB1X4 U70 ( .A0N(n65), .A1N(A[15]), .B0(n66), .Y(n64) );
  NAND2BX4 U71 ( .AN(B[13]), .B(A[13]), .Y(n94) );
  NAND2BX4 U72 ( .AN(A[14]), .B(n13), .Y(n73) );
  NOR2BX2 U73 ( .AN(n28), .B(n35), .Y(n128) );
  OAI2BB1X2 U74 ( .A0N(n128), .A1N(n129), .B0(n30), .Y(n91) );
  NOR2X2 U75 ( .A(n97), .B(n110), .Y(n109) );
  OAI21X4 U76 ( .A0(n101), .A1(n102), .B0(n12), .Y(n98) );
  NAND2BX4 U77 ( .AN(B[14]), .B(A[14]), .Y(n95) );
  NAND2BX4 U78 ( .AN(A[15]), .B(B[15]), .Y(n72) );
  NAND4BX2 U79 ( .AN(n25), .B(n119), .C(n114), .D(n92), .Y(n81) );
  INVX4 U80 ( .A(n114), .Y(n124) );
  NAND2BX4 U81 ( .AN(A[10]), .B(B[10]), .Y(n114) );
  NAND2X4 U82 ( .A(n84), .B(n77), .Y(n75) );
  NOR2X2 U83 ( .A(n71), .B(n70), .Y(n69) );
  NAND2BX4 U84 ( .AN(B[9]), .B(A[9]), .Y(n118) );
  INVX8 U85 ( .A(n105), .Y(n97) );
  NAND2BX4 U86 ( .AN(B[12]), .B(A[12]), .Y(n105) );
  INVX4 U87 ( .A(n116), .Y(n123) );
  INVX4 U88 ( .A(n118), .Y(n21) );
  OAI2BB1X4 U89 ( .A0N(n127), .A1N(n45), .B0(n91), .Y(n23) );
  INVX2 U90 ( .A(n82), .Y(n127) );
  OAI21X2 U91 ( .A0(n37), .A1(n38), .B0(n39), .Y(n32) );
  NAND4X1 U92 ( .A(n49), .B(n132), .C(n52), .D(n63), .Y(n80) );
  NAND2BX4 U93 ( .AN(A[9]), .B(B[9]), .Y(n92) );
  XOR2X2 U94 ( .A(n47), .B(n48), .Y(DIFF[3]) );
  AOI21X1 U95 ( .A0(n49), .A1(n50), .B0(n51), .Y(n48) );
  NAND2BX4 U96 ( .AN(A[1]), .B(B[1]), .Y(n132) );
  OAI21X2 U97 ( .A0(n56), .A1(n57), .B0(n58), .Y(n50) );
  INVX4 U98 ( .A(n132), .Y(n57) );
  NAND2BX4 U99 ( .AN(A[12]), .B(B[12]), .Y(n84) );
  NOR2BX1 U100 ( .AN(n28), .B(n29), .Y(n27) );
  NAND2X4 U101 ( .A(n90), .B(n80), .Y(n45) );
  NOR2X1 U102 ( .A(n80), .B(n81), .Y(n79) );
  INVX4 U103 ( .A(n120), .Y(n25) );
  OR2X2 U104 ( .A(n24), .B(n25), .Y(n15) );
  NAND2XL U105 ( .A(n44), .B(n46), .Y(n17) );
  NAND2BXL U106 ( .AN(B[0]), .B(A[0]), .Y(n62) );
  NAND2BXL U107 ( .AN(A[0]), .B(B[0]), .Y(n63) );
  XOR2X2 U108 ( .A(n26), .B(n27), .Y(DIFF[7]) );
  INVX4 U109 ( .A(n131), .Y(n38) );
  OAI21X2 U110 ( .A0(n134), .A1(n135), .B0(n53), .Y(n133) );
  NAND2X2 U111 ( .A(n45), .B(n46), .Y(n43) );
  XNOR2X4 U112 ( .A(n122), .B(n16), .Y(DIFF[10]) );
  OR2X4 U113 ( .A(n124), .B(n123), .Y(n16) );
  XNOR2X1 U114 ( .A(n45), .B(n17), .Y(DIFF[4]) );
  INVXL U115 ( .A(n39), .Y(n42) );
  INVXL U116 ( .A(n58), .Y(n61) );
  NAND2XL U117 ( .A(n52), .B(n53), .Y(n47) );
  INVXL U118 ( .A(n81), .Y(n85) );
  NAND2XL U119 ( .A(n39), .B(n44), .Y(n130) );
  NAND2BX2 U120 ( .AN(A[2]), .B(B[2]), .Y(n49) );
  NAND2BXL U121 ( .AN(A[3]), .B(B[3]), .Y(n52) );
  NAND2BX1 U122 ( .AN(n63), .B(n62), .Y(n59) );
  NAND2X1 U123 ( .A(n63), .B(n62), .Y(DIFF[0]) );
  XNOR2X4 U124 ( .A(n107), .B(n108), .Y(DIFF[14]) );
  AOI21X1 U125 ( .A0(n85), .A1(n86), .B0(n87), .Y(n74) );
  OAI21XL U126 ( .A0(n90), .A1(n82), .B0(n91), .Y(n86) );
  XNOR2X4 U127 ( .A(n18), .B(n121), .Y(DIFF[11]) );
  NOR2X2 U128 ( .A(n35), .B(n36), .Y(n34) );
  INVX1 U129 ( .A(n30), .Y(n29) );
  NOR2X1 U130 ( .A(n51), .B(n136), .Y(n134) );
  NAND2X1 U131 ( .A(n49), .B(n52), .Y(n135) );
  OAI21X1 U132 ( .A0(n57), .A1(n62), .B0(n58), .Y(n136) );
  INVX1 U133 ( .A(n59), .Y(n56) );
  XOR2X1 U134 ( .A(n50), .B(n54), .Y(DIFF[2]) );
  NOR2XL U135 ( .A(n51), .B(n55), .Y(n54) );
  INVX1 U136 ( .A(n49), .Y(n55) );
  XOR2X1 U137 ( .A(n59), .B(n60), .Y(DIFF[1]) );
  NOR2XL U138 ( .A(n61), .B(n57), .Y(n60) );
  NAND2BXL U139 ( .AN(A[5]), .B(B[5]), .Y(n131) );
  NAND2BXL U140 ( .AN(B[7]), .B(A[7]), .Y(n28) );
  NAND2BXL U141 ( .AN(B[2]), .B(A[2]), .Y(n137) );
  NAND2BXL U142 ( .AN(B[1]), .B(A[1]), .Y(n58) );
  NAND2BXL U143 ( .AN(B[3]), .B(A[3]), .Y(n53) );
  NAND2X2 U144 ( .A(n77), .B(n94), .Y(n111) );
  NOR2X4 U145 ( .A(n71), .B(n100), .Y(n99) );
  XOR2X4 U146 ( .A(n98), .B(n99), .Y(DIFF[15]) );
  NAND2X4 U147 ( .A(n95), .B(n73), .Y(n108) );
  OAI21X4 U148 ( .A0(n75), .A1(n109), .B0(n94), .Y(n107) );
  XOR2X4 U149 ( .A(n112), .B(n111), .Y(DIFF[13]) );
  NAND2BX4 U150 ( .AN(A[13]), .B(B[13]), .Y(n77) );
  NAND3X4 U151 ( .A(n106), .B(n14), .C(n88), .Y(n110) );
  NAND3X4 U152 ( .A(n113), .B(n93), .C(n114), .Y(n88) );
  OAI21X4 U153 ( .A0(n125), .A1(n22), .B0(n118), .Y(n122) );
  OAI21X4 U154 ( .A0(n25), .A1(n126), .B0(n4), .Y(n20) );
  CLKINVX3 U155 ( .A(n133), .Y(n90) );
  CLKINVX3 U156 ( .A(n137), .Y(n51) );
endmodule


module butterfly_DW01_add_36 ( A, B, SUM );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120;

  OAI21X1 U2 ( .A0(B[13]), .A1(n18), .B0(n97), .Y(n85) );
  AOI21X2 U3 ( .A0(n100), .A1(n65), .B0(n97), .Y(n99) );
  BUFX8 U4 ( .A(A[13]), .Y(n18) );
  CLKINVX3 U5 ( .A(n76), .Y(n86) );
  OR2X2 U6 ( .A(A[11]), .B(B[11]), .Y(n3) );
  AND2X2 U7 ( .A(n104), .B(n79), .Y(n14) );
  NOR2BX2 U8 ( .AN(n34), .B(n33), .Y(n36) );
  OAI21X1 U9 ( .A0(n32), .A1(n33), .B0(n34), .Y(n27) );
  CLKINVX8 U10 ( .A(n104), .Y(n26) );
  OR2X4 U11 ( .A(B[13]), .B(A[13]), .Y(n13) );
  NAND4BXL U12 ( .AN(n26), .B(n79), .C(n80), .D(n3), .Y(n67) );
  NAND2X2 U13 ( .A(n38), .B(n8), .Y(n9) );
  NAND2X2 U14 ( .A(n87), .B(n2), .Y(n4) );
  AND2X4 U15 ( .A(n76), .B(n77), .Y(n1) );
  INVX4 U16 ( .A(n87), .Y(n97) );
  NAND3X4 U17 ( .A(n96), .B(n69), .C(n70), .Y(n100) );
  AND2X4 U18 ( .A(n70), .B(n69), .Y(n68) );
  NAND2X4 U19 ( .A(B[9]), .B(A[9]), .Y(n21) );
  NAND2X2 U20 ( .A(B[4]), .B(A[4]), .Y(n41) );
  INVX4 U21 ( .A(n80), .Y(n108) );
  AND2X4 U22 ( .A(n81), .B(n69), .Y(n106) );
  OR2X4 U23 ( .A(A[12]), .B(B[12]), .Y(n2) );
  NAND2X4 U24 ( .A(n1), .B(n78), .Y(n63) );
  NAND2X4 U25 ( .A(B[13]), .B(n18), .Y(n84) );
  NAND3X4 U26 ( .A(n62), .B(n61), .C(n89), .Y(n59) );
  NAND2X4 U27 ( .A(B[11]), .B(A[11]), .Y(n69) );
  NAND3X2 U28 ( .A(n84), .B(n92), .C(n93), .Y(n91) );
  OAI21X4 U29 ( .A0(n113), .A1(n114), .B0(n31), .Y(n74) );
  NAND2X2 U30 ( .A(n29), .B(n34), .Y(n114) );
  NAND2X2 U31 ( .A(n91), .B(n76), .Y(n90) );
  NAND2X4 U32 ( .A(n88), .B(n90), .Y(n10) );
  NAND2BX4 U33 ( .AN(n59), .B(n60), .Y(n7) );
  XOR2X2 U34 ( .A(n54), .B(n56), .Y(SUM[1]) );
  NOR2BX1 U35 ( .AN(n55), .B(n57), .Y(n56) );
  OAI21X2 U36 ( .A0(n22), .A1(n25), .B0(n21), .Y(n102) );
  OR2X2 U37 ( .A(n18), .B(B[13]), .Y(n77) );
  NAND2X2 U38 ( .A(B[15]), .B(A[15]), .Y(n89) );
  INVX4 U39 ( .A(n23), .Y(n112) );
  OR2X4 U40 ( .A(A[6]), .B(B[6]), .Y(n115) );
  XNOR2X4 U41 ( .A(n4), .B(n100), .Y(SUM[12]) );
  NAND3BX4 U42 ( .AN(n63), .B(n64), .C(n2), .Y(n62) );
  INVX4 U43 ( .A(n60), .Y(n5) );
  OAI21X4 U44 ( .A0(n107), .A1(n108), .B0(n103), .Y(n105) );
  INVX2 U45 ( .A(n109), .Y(n107) );
  NAND2X2 U46 ( .A(B[10]), .B(A[10]), .Y(n103) );
  AOI21X2 U47 ( .A0(n84), .A1(n85), .B0(n86), .Y(n83) );
  XOR2X4 U48 ( .A(n19), .B(n20), .Y(SUM[9]) );
  AND2X4 U49 ( .A(n78), .B(n89), .Y(n11) );
  OAI21X2 U50 ( .A0(n82), .A1(n83), .B0(n78), .Y(n61) );
  NAND2X2 U51 ( .A(n84), .B(n77), .Y(n98) );
  OR2X4 U52 ( .A(A[10]), .B(B[10]), .Y(n80) );
  NAND4X2 U53 ( .A(n81), .B(n23), .C(n80), .D(n14), .Y(n96) );
  XOR2X4 U54 ( .A(n105), .B(n106), .Y(SUM[11]) );
  OAI21X4 U55 ( .A0(n112), .A1(n26), .B0(n25), .Y(n19) );
  NOR2BX4 U56 ( .AN(n25), .B(n26), .Y(n24) );
  NAND2X2 U57 ( .A(B[8]), .B(A[8]), .Y(n25) );
  NAND2X2 U58 ( .A(B[7]), .B(A[7]), .Y(n29) );
  NAND3X4 U59 ( .A(n13), .B(n65), .C(n95), .Y(n93) );
  NAND2X4 U60 ( .A(n13), .B(n97), .Y(n92) );
  NAND3X2 U61 ( .A(n96), .B(n70), .C(n69), .Y(n95) );
  OR2X4 U62 ( .A(B[14]), .B(A[14]), .Y(n76) );
  NAND2X2 U63 ( .A(A[12]), .B(B[12]), .Y(n87) );
  CLKINVX3 U64 ( .A(n75), .Y(n71) );
  NAND4BBX2 U65 ( .AN(n16), .BN(n17), .C(n115), .D(n31), .Y(n75) );
  INVX8 U66 ( .A(n79), .Y(n22) );
  NOR2BX4 U67 ( .AN(n21), .B(n22), .Y(n20) );
  XOR2X4 U68 ( .A(B[16]), .B(A[16]), .Y(n60) );
  OAI21X4 U69 ( .A0(n22), .A1(n111), .B0(n21), .Y(n109) );
  NAND2X4 U70 ( .A(n3), .B(n101), .Y(n70) );
  OAI2BB1X4 U71 ( .A0N(n80), .A1N(n102), .B0(n103), .Y(n101) );
  XOR2X4 U72 ( .A(n98), .B(n99), .Y(SUM[13]) );
  INVX2 U73 ( .A(n19), .Y(n111) );
  AOI211X4 U74 ( .A0(n37), .A1(n41), .B0(n33), .C0(n16), .Y(n113) );
  NAND2X4 U75 ( .A(B[5]), .B(A[5]), .Y(n37) );
  NOR2X4 U76 ( .A(A[5]), .B(B[5]), .Y(n16) );
  INVX8 U77 ( .A(n72), .Y(n40) );
  XOR2X4 U78 ( .A(n27), .B(n28), .Y(SUM[7]) );
  NAND2X2 U79 ( .A(n59), .B(n5), .Y(n6) );
  NAND2X4 U80 ( .A(n6), .B(n7), .Y(SUM[16]) );
  NAND2X4 U81 ( .A(n9), .B(n37), .Y(n35) );
  INVXL U82 ( .A(n16), .Y(n8) );
  XOR2X4 U83 ( .A(n35), .B(n36), .Y(SUM[6]) );
  INVX4 U84 ( .A(n35), .Y(n32) );
  XOR2X4 U85 ( .A(n109), .B(n110), .Y(SUM[10]) );
  OR2X4 U86 ( .A(A[12]), .B(B[12]), .Y(n65) );
  OAI21X4 U87 ( .A0(n17), .A1(n40), .B0(n41), .Y(n38) );
  OAI21X4 U88 ( .A0(n117), .A1(n118), .B0(n45), .Y(n72) );
  XOR2X4 U89 ( .A(n11), .B(n10), .Y(SUM[15]) );
  NAND2XL U90 ( .A(B[0]), .B(A[0]), .Y(n58) );
  INVXL U91 ( .A(n31), .Y(n30) );
  NAND2XL U92 ( .A(B[2]), .B(A[2]), .Y(n49) );
  OR2XL U93 ( .A(A[2]), .B(B[2]), .Y(n52) );
  OR2XL U94 ( .A(A[3]), .B(B[3]), .Y(n116) );
  NAND2XL U95 ( .A(B[3]), .B(A[3]), .Y(n45) );
  OR2XL U96 ( .A(A[1]), .B(B[1]), .Y(n53) );
  NAND2XL U97 ( .A(B[1]), .B(A[1]), .Y(n55) );
  NOR2BX1 U98 ( .AN(n58), .B(n12), .Y(SUM[0]) );
  NOR2XL U99 ( .A(A[0]), .B(B[0]), .Y(n12) );
  INVXL U100 ( .A(n74), .Y(n73) );
  NOR2BXL U101 ( .AN(n37), .B(n16), .Y(n39) );
  NOR2X2 U102 ( .A(n119), .B(n120), .Y(n117) );
  OAI21X2 U103 ( .A0(n57), .A1(n58), .B0(n55), .Y(n120) );
  INVX4 U104 ( .A(n115), .Y(n33) );
  OAI2BB1X2 U105 ( .A0N(n53), .A1N(n54), .B0(n55), .Y(n50) );
  XOR2X1 U106 ( .A(n50), .B(n51), .Y(SUM[2]) );
  NOR2BXL U107 ( .AN(n49), .B(n48), .Y(n51) );
  INVX1 U108 ( .A(n58), .Y(n54) );
  INVX1 U109 ( .A(n50), .Y(n47) );
  NAND2X1 U110 ( .A(n52), .B(n116), .Y(n118) );
  XOR2X1 U111 ( .A(n23), .B(n24), .Y(SUM[8]) );
  XOR2X1 U112 ( .A(n38), .B(n39), .Y(SUM[5]) );
  NOR2BX1 U113 ( .AN(n29), .B(n30), .Y(n28) );
  INVX1 U114 ( .A(n49), .Y(n119) );
  INVX1 U115 ( .A(n53), .Y(n57) );
  INVX1 U116 ( .A(n52), .Y(n48) );
  XOR2X1 U117 ( .A(n43), .B(n44), .Y(SUM[3]) );
  NOR2BX1 U118 ( .AN(n45), .B(n46), .Y(n44) );
  OAI21XL U119 ( .A0(n47), .A1(n48), .B0(n49), .Y(n43) );
  INVX1 U120 ( .A(n116), .Y(n46) );
  XOR2X1 U121 ( .A(n72), .B(n42), .Y(SUM[4]) );
  NOR2BX1 U122 ( .AN(n41), .B(n17), .Y(n42) );
  XOR2X4 U123 ( .A(n15), .B(n94), .Y(SUM[14]) );
  AND3X4 U124 ( .A(n92), .B(n84), .C(n93), .Y(n15) );
  INVXL U125 ( .A(n88), .Y(n82) );
  OAI21XL U126 ( .A0(n66), .A1(n67), .B0(n68), .Y(n64) );
  AOI21XL U127 ( .A0(n71), .A1(n72), .B0(n73), .Y(n66) );
  NOR2X2 U128 ( .A(A[4]), .B(B[4]), .Y(n17) );
  NAND2XL U129 ( .A(B[6]), .B(A[6]), .Y(n34) );
  NAND2X2 U130 ( .A(B[14]), .B(A[14]), .Y(n88) );
  OR2X4 U131 ( .A(B[15]), .B(A[15]), .Y(n78) );
  NAND2X4 U132 ( .A(n88), .B(n76), .Y(n94) );
  OR2X4 U133 ( .A(A[11]), .B(B[11]), .Y(n81) );
  NOR2BX4 U134 ( .AN(n103), .B(n108), .Y(n110) );
  OR2X4 U135 ( .A(A[8]), .B(B[8]), .Y(n104) );
  OAI21X4 U136 ( .A0(n40), .A1(n75), .B0(n74), .Y(n23) );
  OR2X4 U137 ( .A(A[7]), .B(B[7]), .Y(n31) );
  OR2X4 U138 ( .A(A[9]), .B(B[9]), .Y(n79) );
endmodule


module butterfly_DW01_add_44 ( A, B, SUM );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  wire   n133, n134, n135, n1, n2, n4, n5, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132;

  INVX2 U2 ( .A(n100), .Y(n1) );
  INVX2 U3 ( .A(n76), .Y(n100) );
  AND2X2 U4 ( .A(n11), .B(n1), .Y(n24) );
  INVX4 U5 ( .A(n77), .Y(n11) );
  NOR2X2 U6 ( .A(n13), .B(n7), .Y(n106) );
  INVX2 U7 ( .A(n73), .Y(n72) );
  INVX8 U8 ( .A(n126), .Y(n41) );
  CLKINVX2 U9 ( .A(n97), .Y(n96) );
  OAI21X4 U10 ( .A0(n124), .A1(n125), .B0(n39), .Y(n97) );
  NOR2BX1 U11 ( .AN(n42), .B(n41), .Y(n44) );
  NAND2X2 U12 ( .A(n37), .B(n42), .Y(n125) );
  XOR2X4 U13 ( .A(n105), .B(n111), .Y(SUM[12]) );
  CLKINVX8 U14 ( .A(n4), .Y(n2) );
  INVX8 U15 ( .A(n2), .Y(SUM[15]) );
  XOR2X4 U16 ( .A(n99), .B(n98), .Y(n4) );
  INVX8 U17 ( .A(n95), .Y(n127) );
  NAND2X4 U18 ( .A(B[10]), .B(A[10]), .Y(n120) );
  NOR3X4 U19 ( .A(n77), .B(n7), .C(n13), .Y(n83) );
  NOR2X2 U20 ( .A(A[4]), .B(B[4]), .Y(n26) );
  OAI21X2 U21 ( .A0(n26), .A1(n127), .B0(n49), .Y(n47) );
  NOR2BX1 U22 ( .AN(n46), .B(n25), .Y(n48) );
  INVX4 U23 ( .A(n93), .Y(n34) );
  OAI21X4 U24 ( .A0(n45), .A1(n25), .B0(n46), .Y(n43) );
  NAND2X4 U25 ( .A(B[5]), .B(A[5]), .Y(n46) );
  CLKINVX4 U26 ( .A(n27), .Y(n122) );
  XOR2X2 U27 ( .A(n27), .B(n28), .Y(SUM[9]) );
  AND2X4 U28 ( .A(n120), .B(n91), .Y(n121) );
  INVX4 U29 ( .A(n120), .Y(n119) );
  OR2X2 U30 ( .A(B[12]), .B(A[12]), .Y(n109) );
  NAND2X4 U31 ( .A(n123), .B(n33), .Y(n27) );
  NAND2X4 U32 ( .A(n31), .B(n93), .Y(n123) );
  NAND2X4 U33 ( .A(B[12]), .B(A[12]), .Y(n110) );
  XOR2X2 U34 ( .A(n31), .B(n32), .Y(SUM[8]) );
  CLKINVXL U35 ( .A(n80), .Y(n94) );
  BUFX20 U36 ( .A(n134), .Y(SUM[13]) );
  NAND2X2 U37 ( .A(B[7]), .B(A[7]), .Y(n37) );
  CLKINVX8 U38 ( .A(n133), .Y(n5) );
  INVX8 U39 ( .A(n5), .Y(SUM[14]) );
  NOR2X4 U40 ( .A(B[12]), .B(A[12]), .Y(n7) );
  NAND2X1 U41 ( .A(A[12]), .B(B[12]), .Y(n74) );
  OR2XL U42 ( .A(B[13]), .B(A[13]), .Y(n8) );
  OAI2BB1X4 U43 ( .A0N(n14), .A1N(n17), .B0(n73), .Y(n98) );
  OR2X4 U44 ( .A(B[11]), .B(A[11]), .Y(n9) );
  XOR2X4 U45 ( .A(n116), .B(n117), .Y(SUM[11]) );
  NAND2X4 U46 ( .A(n10), .B(n112), .Y(n105) );
  AND2X4 U47 ( .A(n88), .B(n89), .Y(n10) );
  INVXL U48 ( .A(A[15]), .Y(n14) );
  INVX4 U49 ( .A(n11), .Y(n12) );
  XOR2X4 U50 ( .A(n108), .B(n107), .Y(n134) );
  NAND2X2 U51 ( .A(n8), .B(n75), .Y(n107) );
  NOR2X4 U52 ( .A(B[13]), .B(A[13]), .Y(n13) );
  NAND2X4 U53 ( .A(B[13]), .B(A[13]), .Y(n75) );
  AOI21X2 U54 ( .A0(n109), .A1(n105), .B0(n104), .Y(n108) );
  CLKINVX8 U55 ( .A(n90), .Y(n30) );
  NAND2X2 U56 ( .A(B[9]), .B(A[9]), .Y(n29) );
  BUFX16 U57 ( .A(n135), .Y(SUM[10]) );
  XOR2X4 U58 ( .A(n118), .B(n121), .Y(n135) );
  NAND2X2 U59 ( .A(A[14]), .B(B[14]), .Y(n76) );
  NAND3BX2 U60 ( .AN(n81), .B(n83), .C(n82), .Y(n68) );
  XNOR2X4 U61 ( .A(n16), .B(n67), .Y(n15) );
  NAND2X4 U62 ( .A(n69), .B(n68), .Y(n16) );
  NOR2X4 U63 ( .A(n81), .B(n77), .Y(n70) );
  XOR2X2 U64 ( .A(n43), .B(n44), .Y(SUM[6]) );
  INVX4 U65 ( .A(n110), .Y(n104) );
  NOR2BX4 U66 ( .AN(n110), .B(n7), .Y(n111) );
  INVXL U67 ( .A(B[15]), .Y(n17) );
  NAND2X2 U68 ( .A(B[15]), .B(A[15]), .Y(n73) );
  NAND2X2 U69 ( .A(n102), .B(n75), .Y(n103) );
  OAI22X4 U70 ( .A0(n114), .A1(n115), .B0(A[10]), .B1(B[10]), .Y(n113) );
  OAI211X2 U71 ( .A0(n13), .A1(n74), .B0(n75), .C0(n76), .Y(n71) );
  NAND2X2 U72 ( .A(B[11]), .B(A[11]), .Y(n89) );
  NOR2X4 U73 ( .A(B[15]), .B(A[15]), .Y(n81) );
  NAND4BX2 U74 ( .AN(n22), .B(n31), .C(n91), .D(n9), .Y(n112) );
  OAI21X4 U75 ( .A0(n30), .A1(n122), .B0(n29), .Y(n118) );
  OAI21X2 U76 ( .A0(n84), .A1(n79), .B0(n85), .Y(n82) );
  NOR2X4 U77 ( .A(n30), .B(n33), .Y(n114) );
  AOI21X2 U78 ( .A0(n91), .A1(n118), .B0(n119), .Y(n117) );
  INVX2 U79 ( .A(n47), .Y(n45) );
  XOR2X4 U80 ( .A(n35), .B(n36), .Y(SUM[7]) );
  OAI21X2 U81 ( .A0(n40), .A1(n41), .B0(n42), .Y(n35) );
  AND2X4 U82 ( .A(n70), .B(n71), .Y(n18) );
  NOR2X4 U83 ( .A(n18), .B(n72), .Y(n69) );
  XOR2X4 U84 ( .A(n24), .B(n103), .Y(n133) );
  INVX8 U85 ( .A(n15), .Y(SUM[16]) );
  XOR2X4 U86 ( .A(B[16]), .B(A[16]), .Y(n67) );
  NAND4BBX2 U87 ( .AN(n25), .BN(n26), .C(n126), .D(n39), .Y(n80) );
  NAND2X4 U88 ( .A(B[2]), .B(A[2]), .Y(n57) );
  OR2XL U89 ( .A(A[2]), .B(B[2]), .Y(n60) );
  NAND2X1 U90 ( .A(B[1]), .B(A[1]), .Y(n63) );
  OAI21X4 U91 ( .A0(n127), .A1(n80), .B0(n97), .Y(n31) );
  INVXL U92 ( .A(n88), .Y(n87) );
  INVXL U93 ( .A(n89), .Y(n86) );
  INVXL U94 ( .A(n128), .Y(n54) );
  OAI2BB1X1 U95 ( .A0N(n61), .A1N(n62), .B0(n63), .Y(n58) );
  NAND2X1 U96 ( .A(B[6]), .B(A[6]), .Y(n42) );
  NAND2XL U97 ( .A(B[3]), .B(A[3]), .Y(n53) );
  NAND2XL U98 ( .A(n93), .B(n90), .Y(n22) );
  OAI21X4 U99 ( .A0(n129), .A1(n130), .B0(n53), .Y(n95) );
  NOR2X2 U100 ( .A(n131), .B(n132), .Y(n129) );
  OAI21X2 U101 ( .A0(n65), .A1(n66), .B0(n63), .Y(n132) );
  OAI21X1 U102 ( .A0(n55), .A1(n56), .B0(n57), .Y(n51) );
  OR2X4 U103 ( .A(A[8]), .B(B[8]), .Y(n93) );
  OR2X4 U104 ( .A(A[3]), .B(B[3]), .Y(n128) );
  OR2X4 U105 ( .A(A[1]), .B(B[1]), .Y(n61) );
  NAND2X4 U106 ( .A(B[0]), .B(A[0]), .Y(n66) );
  NOR2BX1 U107 ( .AN(n66), .B(n23), .Y(SUM[0]) );
  NOR2XL U108 ( .A(A[0]), .B(B[0]), .Y(n23) );
  NOR2BX1 U109 ( .AN(n29), .B(n30), .Y(n28) );
  INVX1 U110 ( .A(n58), .Y(n55) );
  AOI21X1 U111 ( .A0(n94), .A1(n95), .B0(n96), .Y(n84) );
  NAND4BXL U112 ( .AN(n34), .B(n90), .C(n91), .D(n9), .Y(n79) );
  NOR2X1 U113 ( .A(n86), .B(n87), .Y(n85) );
  NAND2XL U114 ( .A(n89), .B(n9), .Y(n116) );
  NOR2BX1 U115 ( .AN(n33), .B(n34), .Y(n32) );
  XOR2X1 U116 ( .A(n47), .B(n48), .Y(SUM[5]) );
  NOR2BX1 U117 ( .AN(n37), .B(n38), .Y(n36) );
  INVX1 U118 ( .A(n43), .Y(n40) );
  NAND2X1 U119 ( .A(n60), .B(n128), .Y(n130) );
  INVX1 U120 ( .A(n61), .Y(n65) );
  INVX1 U121 ( .A(n57), .Y(n131) );
  INVXL U122 ( .A(n39), .Y(n38) );
  XOR2X1 U123 ( .A(n51), .B(n52), .Y(SUM[3]) );
  NOR2BX1 U124 ( .AN(n53), .B(n54), .Y(n52) );
  XOR2X1 U125 ( .A(n95), .B(n50), .Y(SUM[4]) );
  NOR2BX1 U126 ( .AN(n49), .B(n26), .Y(n50) );
  INVX1 U127 ( .A(n60), .Y(n56) );
  XOR2X1 U128 ( .A(n62), .B(n64), .Y(SUM[1]) );
  NOR2BXL U129 ( .AN(n63), .B(n65), .Y(n64) );
  XOR2X1 U130 ( .A(n58), .B(n59), .Y(SUM[2]) );
  NOR2BXL U131 ( .AN(n57), .B(n56), .Y(n59) );
  INVX1 U132 ( .A(n66), .Y(n62) );
  INVX2 U133 ( .A(n29), .Y(n115) );
  NOR2X4 U134 ( .A(A[5]), .B(B[5]), .Y(n25) );
  NAND2X1 U135 ( .A(B[4]), .B(A[4]), .Y(n49) );
  INVX8 U136 ( .A(n78), .Y(n77) );
  NOR2X4 U137 ( .A(n101), .B(n100), .Y(n99) );
  AOI21X4 U138 ( .A0(n75), .A1(n102), .B0(n12), .Y(n101) );
  OAI21X4 U139 ( .A0(n104), .A1(n105), .B0(n106), .Y(n102) );
  OR2X4 U140 ( .A(B[14]), .B(A[14]), .Y(n78) );
  OAI2BB1X4 U141 ( .A0N(n113), .A1N(n120), .B0(n92), .Y(n88) );
  OR2X4 U142 ( .A(A[11]), .B(B[11]), .Y(n92) );
  OR2X4 U143 ( .A(A[10]), .B(B[10]), .Y(n91) );
  NAND2X4 U144 ( .A(B[8]), .B(A[8]), .Y(n33) );
  AOI211X2 U145 ( .A0(n46), .A1(n49), .B0(n41), .C0(n25), .Y(n124) );
  OR2X4 U146 ( .A(A[7]), .B(B[7]), .Y(n39) );
  OR2X4 U147 ( .A(A[6]), .B(B[6]), .Y(n126) );
  OR2X4 U148 ( .A(A[9]), .B(B[9]), .Y(n90) );
endmodule


module butterfly_DW01_sub_35 ( A, B, DIFF );
  input [16:0] A;
  input [16:0] B;
  output [16:0] DIFF;
  wire   n143, n144, n145, n146, n1, n2, n3, n4, n5, n6, n7, n8, n9, n11, n12,
         n13, n14, n15, n16, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142;

  NAND2X2 U3 ( .A(n75), .B(n102), .Y(n21) );
  INVX4 U4 ( .A(n102), .Y(n101) );
  INVX2 U5 ( .A(A[14]), .Y(n1) );
  CLKINVX4 U6 ( .A(n1), .Y(n2) );
  AOI21X4 U7 ( .A0(n99), .A1(n100), .B0(n101), .Y(n74) );
  NAND3X2 U8 ( .A(n103), .B(n104), .C(n90), .Y(n99) );
  XOR2X2 U9 ( .A(n31), .B(n32), .Y(DIFF[8]) );
  NOR2X2 U10 ( .A(n33), .B(n34), .Y(n32) );
  BUFX8 U11 ( .A(B[9]), .Y(n3) );
  AOI2BB1X4 U12 ( .A0N(n133), .A1N(n30), .B0(n5), .Y(n4) );
  CLKINVX12 U13 ( .A(n4), .Y(n130) );
  CLKINVX20 U14 ( .A(n125), .Y(n5) );
  XOR2X4 U15 ( .A(n130), .B(n131), .Y(DIFF[10]) );
  NAND4BBX4 U16 ( .AN(n30), .BN(n6), .C(n121), .D(n98), .Y(n115) );
  OR2X4 U17 ( .A(n126), .B(n34), .Y(n6) );
  INVX8 U18 ( .A(n106), .Y(n118) );
  INVX8 U19 ( .A(n100), .Y(n108) );
  NAND2BX4 U20 ( .AN(B[14]), .B(n2), .Y(n100) );
  NAND2BX4 U21 ( .AN(n112), .B(n113), .Y(n7) );
  NAND2BX4 U22 ( .AN(A[10]), .B(B[10]), .Y(n121) );
  INVX2 U23 ( .A(n87), .Y(n86) );
  OAI21X2 U24 ( .A0(n79), .A1(n80), .B0(n81), .Y(n78) );
  AOI21X2 U25 ( .A0(n93), .A1(B[15]), .B0(n94), .Y(n92) );
  XOR2X2 U26 ( .A(n41), .B(n43), .Y(DIFF[6]) );
  NAND2X2 U27 ( .A(n54), .B(n55), .Y(n52) );
  XOR2X2 U28 ( .A(n49), .B(n50), .Y(DIFF[5]) );
  INVX2 U29 ( .A(n49), .Y(n46) );
  XNOR2X2 U30 ( .A(n127), .B(n13), .Y(n146) );
  OAI2BB1XL U31 ( .A0N(n40), .A1N(n41), .B0(n42), .Y(n35) );
  OAI21X2 U32 ( .A0(n46), .A1(n47), .B0(n48), .Y(n41) );
  OAI21X1 U33 ( .A0(n4), .A1(n129), .B0(n123), .Y(n127) );
  NOR2X4 U34 ( .A(n132), .B(n129), .Y(n131) );
  INVX4 U35 ( .A(n121), .Y(n129) );
  XOR2X2 U36 ( .A(n27), .B(n28), .Y(DIFF[9]) );
  INVX8 U37 ( .A(n31), .Y(n126) );
  NAND4BX2 U38 ( .AN(n34), .B(n97), .C(n121), .D(n98), .Y(n80) );
  INVX2 U39 ( .A(n98), .Y(n128) );
  BUFX16 U40 ( .A(n145), .Y(DIFF[13]) );
  BUFX16 U41 ( .A(n144), .Y(DIFF[14]) );
  XNOR2X4 U42 ( .A(n116), .B(n8), .Y(n145) );
  AND2X2 U43 ( .A(n90), .B(n105), .Y(n8) );
  NAND2X4 U44 ( .A(n7), .B(n15), .Y(n22) );
  CLKINVX8 U45 ( .A(n11), .Y(n12) );
  INVX4 U46 ( .A(A[13]), .Y(n11) );
  INVX4 U47 ( .A(n93), .Y(n9) );
  INVX4 U48 ( .A(A[15]), .Y(n93) );
  XNOR2X4 U49 ( .A(n73), .B(n16), .Y(DIFF[16]) );
  OR2X4 U50 ( .A(n114), .B(n128), .Y(n13) );
  NAND3X2 U51 ( .A(n88), .B(n89), .C(n90), .Y(n14) );
  NAND2X4 U52 ( .A(n88), .B(n90), .Y(n112) );
  INVX4 U53 ( .A(n27), .Y(n133) );
  CLKINVX4 U54 ( .A(n42), .Y(n44) );
  NAND2BX4 U55 ( .AN(B[15]), .B(n9), .Y(n75) );
  NAND3BX4 U56 ( .AN(n91), .B(n92), .C(n103), .Y(n76) );
  NAND4BX2 U57 ( .AN(n80), .B(n90), .C(n84), .D(n95), .Y(n91) );
  NAND2BX4 U58 ( .AN(A[14]), .B(B[14]), .Y(n103) );
  NAND3X4 U59 ( .A(n115), .B(n82), .C(n83), .Y(n117) );
  BUFX12 U60 ( .A(n146), .Y(DIFF[11]) );
  NAND3BX4 U61 ( .AN(n14), .B(n78), .C(n102), .Y(n77) );
  NAND4BX4 U62 ( .AN(n114), .B(n115), .C(n83), .D(n106), .Y(n113) );
  INVX4 U63 ( .A(n88), .Y(n94) );
  BUFX4 U64 ( .A(n105), .Y(n15) );
  INVX4 U65 ( .A(n82), .Y(n114) );
  NAND2BX4 U66 ( .AN(B[11]), .B(A[11]), .Y(n82) );
  NAND2X4 U67 ( .A(n105), .B(n106), .Y(n104) );
  NAND2BX4 U68 ( .AN(A[9]), .B(n3), .Y(n97) );
  NOR2X4 U69 ( .A(n111), .B(n108), .Y(n23) );
  INVX12 U70 ( .A(n89), .Y(n111) );
  XOR2X4 U71 ( .A(n23), .B(n22), .Y(n144) );
  BUFX20 U72 ( .A(n143), .Y(DIFF[15]) );
  NAND2BX2 U73 ( .AN(A[8]), .B(B[8]), .Y(n134) );
  AOI21X4 U74 ( .A0(n110), .A1(n15), .B0(n111), .Y(n109) );
  NAND4BX4 U75 ( .AN(n74), .B(n76), .C(n77), .D(n75), .Y(n73) );
  XOR2X4 U76 ( .A(B[16]), .B(A[16]), .Y(n16) );
  OAI21X4 U77 ( .A0(n126), .A1(n34), .B0(n124), .Y(n27) );
  INVX4 U78 ( .A(n134), .Y(n34) );
  AND2X4 U79 ( .A(n83), .B(n82), .Y(n81) );
  XOR2X4 U80 ( .A(n35), .B(n36), .Y(DIFF[7]) );
  OAI2BB1X4 U81 ( .A0N(n84), .A1N(n54), .B0(n87), .Y(n31) );
  NAND3X4 U82 ( .A(n120), .B(n121), .C(n98), .Y(n83) );
  NAND3BX2 U83 ( .AN(n29), .B(n122), .C(n123), .Y(n120) );
  XOR2X4 U84 ( .A(n107), .B(n21), .Y(n143) );
  NAND2BX4 U85 ( .AN(A[15]), .B(B[15]), .Y(n102) );
  AOI21X2 U86 ( .A0(n117), .A1(n88), .B0(n118), .Y(n116) );
  NOR2BX2 U87 ( .AN(n37), .B(n44), .Y(n135) );
  NAND2BX4 U88 ( .AN(A[13]), .B(B[13]), .Y(n90) );
  NAND2BX2 U89 ( .AN(B[7]), .B(A[7]), .Y(n37) );
  NAND2BX4 U90 ( .AN(B[8]), .B(A[8]), .Y(n124) );
  NAND2BX2 U91 ( .AN(B[5]), .B(A[5]), .Y(n48) );
  NAND2BX1 U92 ( .AN(B[1]), .B(A[1]), .Y(n67) );
  NAND2BX2 U93 ( .AN(B[2]), .B(A[2]), .Y(n141) );
  INVX4 U94 ( .A(n97), .Y(n30) );
  NAND2BX4 U95 ( .AN(n85), .B(n96), .Y(n54) );
  AOI21XL U96 ( .A0(n58), .A1(n59), .B0(n60), .Y(n57) );
  NAND2XL U97 ( .A(n61), .B(n62), .Y(n56) );
  AND2X2 U98 ( .A(n58), .B(n61), .Y(n26) );
  OR2X2 U99 ( .A(n60), .B(n140), .Y(n25) );
  NAND2BX2 U100 ( .AN(A[1]), .B(B[1]), .Y(n139) );
  NAND2BX1 U101 ( .AN(B[3]), .B(A[3]), .Y(n62) );
  NAND4BX2 U102 ( .AN(n47), .B(n55), .C(n40), .D(n39), .Y(n142) );
  NAND2XL U103 ( .A(n52), .B(n53), .Y(n49) );
  XNOR2X1 U104 ( .A(n54), .B(n24), .Y(DIFF[4]) );
  NAND2XL U105 ( .A(n53), .B(n55), .Y(n24) );
  OAI21XL U106 ( .A0(n65), .A1(n66), .B0(n67), .Y(n59) );
  INVX2 U107 ( .A(n68), .Y(n65) );
  INVXL U108 ( .A(n96), .Y(n95) );
  NOR2XL U109 ( .A(n60), .B(n64), .Y(n63) );
  NAND2BX4 U110 ( .AN(B[6]), .B(A[6]), .Y(n42) );
  NAND2BX4 U111 ( .AN(A[5]), .B(B[5]), .Y(n138) );
  NAND2BX4 U112 ( .AN(A[2]), .B(B[2]), .Y(n58) );
  NAND2BX4 U113 ( .AN(A[3]), .B(B[3]), .Y(n61) );
  OAI2BB1X4 U114 ( .A0N(n25), .A1N(n26), .B0(n62), .Y(n85) );
  NAND2BX4 U115 ( .AN(B[0]), .B(A[0]), .Y(n71) );
  NAND2BXL U116 ( .AN(A[0]), .B(B[0]), .Y(n72) );
  NOR2X1 U117 ( .A(n29), .B(n30), .Y(n28) );
  INVX1 U118 ( .A(n123), .Y(n132) );
  INVX1 U119 ( .A(n138), .Y(n47) );
  INVX1 U120 ( .A(n124), .Y(n33) );
  OAI2BB1X2 U121 ( .A0N(n135), .A1N(n136), .B0(n39), .Y(n87) );
  NAND3X1 U122 ( .A(n40), .B(n137), .C(n138), .Y(n136) );
  NAND2X1 U123 ( .A(n48), .B(n53), .Y(n137) );
  AOI21XL U124 ( .A0(n84), .A1(n85), .B0(n86), .Y(n79) );
  NOR2XL U125 ( .A(n44), .B(n45), .Y(n43) );
  INVXL U126 ( .A(n40), .Y(n45) );
  NOR2XL U127 ( .A(n51), .B(n47), .Y(n50) );
  INVX1 U128 ( .A(n48), .Y(n51) );
  NOR2BX1 U129 ( .AN(n37), .B(n38), .Y(n36) );
  INVXL U130 ( .A(n39), .Y(n38) );
  INVX1 U131 ( .A(n139), .Y(n66) );
  XOR2X1 U132 ( .A(n59), .B(n63), .Y(DIFF[2]) );
  INVX1 U133 ( .A(n58), .Y(n64) );
  XOR2X1 U134 ( .A(n56), .B(n57), .Y(DIFF[3]) );
  XOR2X1 U135 ( .A(n68), .B(n69), .Y(DIFF[1]) );
  NOR2XL U136 ( .A(n70), .B(n66), .Y(n69) );
  INVX1 U137 ( .A(n67), .Y(n70) );
  NAND2X1 U138 ( .A(n33), .B(n97), .Y(n122) );
  OAI21X1 U139 ( .A0(n66), .A1(n71), .B0(n67), .Y(n140) );
  NAND2BX2 U140 ( .AN(A[4]), .B(B[4]), .Y(n55) );
  NAND2BX2 U141 ( .AN(B[4]), .B(A[4]), .Y(n53) );
  NAND4X1 U142 ( .A(n58), .B(n139), .C(n61), .D(n72), .Y(n96) );
  NAND2BX1 U143 ( .AN(n72), .B(n71), .Y(n68) );
  NAND2X1 U144 ( .A(n72), .B(n71), .Y(DIFF[0]) );
  NAND2BX4 U145 ( .AN(B[13]), .B(n12), .Y(n105) );
  NOR2X4 U146 ( .A(n109), .B(n108), .Y(n107) );
  NAND2BX4 U147 ( .AN(A[14]), .B(B[14]), .Y(n89) );
  NAND2BX4 U148 ( .AN(n112), .B(n113), .Y(n110) );
  XOR2X4 U149 ( .A(n117), .B(n119), .Y(DIFF[12]) );
  NOR2X4 U150 ( .A(n118), .B(n94), .Y(n119) );
  NAND2BX4 U151 ( .AN(A[12]), .B(B[12]), .Y(n88) );
  NAND2BX4 U152 ( .AN(B[12]), .B(A[12]), .Y(n106) );
  CLKINVX3 U153 ( .A(n125), .Y(n29) );
  NAND2BX4 U154 ( .AN(A[11]), .B(B[11]), .Y(n98) );
  NAND2BX4 U155 ( .AN(B[10]), .B(A[10]), .Y(n123) );
  NAND2BX4 U156 ( .AN(B[9]), .B(A[9]), .Y(n125) );
  CLKINVX3 U157 ( .A(n141), .Y(n60) );
  CLKINVX3 U158 ( .A(n142), .Y(n84) );
  NAND2BX4 U159 ( .AN(A[7]), .B(B[7]), .Y(n39) );
  NAND2BX4 U160 ( .AN(A[6]), .B(B[6]), .Y(n40) );
endmodule


module butterfly_DW01_add_49 ( A, B, SUM );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  wire   n144, n145, n146, n147, n148, n149, n1, n2, n3, n5, n6, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n34, n35, n36, n37, n38, n39, n40, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143;

  NAND4X4 U2 ( .A(n1), .B(n2), .C(n3), .D(n112), .Y(n120) );
  CLKINVX20 U3 ( .A(n34), .Y(n1) );
  CLKINVX20 U4 ( .A(n9), .Y(n2) );
  AND2X2 U5 ( .A(n103), .B(n100), .Y(n23) );
  INVX2 U6 ( .A(n119), .Y(n105) );
  CLKINVX1 U7 ( .A(n123), .Y(n6) );
  BUFX8 U8 ( .A(n111), .Y(n3) );
  OAI2BB1X2 U9 ( .A0N(B[12]), .A1N(A[12]), .B0(n119), .Y(n118) );
  NAND4BXL U10 ( .AN(n51), .B(n110), .C(n3), .D(n112), .Y(n91) );
  NAND4X2 U11 ( .A(n16), .B(n101), .C(n6), .D(n103), .Y(n88) );
  OAI21X2 U12 ( .A0(n108), .A1(n8), .B0(n109), .Y(n106) );
  OR2X4 U13 ( .A(A[12]), .B(B[12]), .Y(n103) );
  CLKINVX4 U14 ( .A(n20), .Y(n101) );
  BUFX12 U15 ( .A(n149), .Y(SUM[6]) );
  BUFX8 U16 ( .A(n93), .Y(n5) );
  AND3X4 U17 ( .A(n94), .B(n120), .C(n5), .Y(n18) );
  AND2X2 U18 ( .A(n94), .B(n5), .Y(n92) );
  NAND2X2 U19 ( .A(n111), .B(n135), .Y(n11) );
  OR2X4 U20 ( .A(B[11]), .B(A[11]), .Y(n112) );
  NAND2X2 U21 ( .A(B[9]), .B(A[9]), .Y(n46) );
  NOR2X4 U22 ( .A(n10), .B(n20), .Y(n115) );
  NAND2BX4 U23 ( .AN(n88), .B(n89), .Y(n87) );
  INVX8 U24 ( .A(n102), .Y(n123) );
  OAI2BB1X2 U25 ( .A0N(n80), .A1N(n81), .B0(n82), .Y(n77) );
  OAI21X2 U26 ( .A0(n74), .A1(n75), .B0(n76), .Y(n69) );
  NAND2X2 U27 ( .A(n120), .B(n126), .Y(n125) );
  INVX2 U28 ( .A(n52), .Y(n27) );
  INVXL U29 ( .A(n48), .Y(n9) );
  OAI21X1 U30 ( .A0(n90), .A1(n91), .B0(n92), .Y(n89) );
  BUFX12 U31 ( .A(n148), .Y(SUM[7]) );
  INVXL U32 ( .A(n130), .Y(n8) );
  INVX4 U33 ( .A(n100), .Y(n108) );
  AND2X2 U34 ( .A(B[15]), .B(A[15]), .Y(n10) );
  NAND3X4 U35 ( .A(n17), .B(n3), .C(n131), .Y(n94) );
  AND2X4 U36 ( .A(n11), .B(n132), .Y(n134) );
  NAND2X4 U37 ( .A(n132), .B(n111), .Y(n12) );
  NAND2X4 U38 ( .A(B[10]), .B(A[10]), .Y(n132) );
  INVX4 U39 ( .A(n140), .Y(n55) );
  XNOR2X4 U40 ( .A(n135), .B(n12), .Y(n147) );
  XOR2X4 U41 ( .A(n86), .B(n14), .Y(n13) );
  CLKINVX20 U42 ( .A(n13), .Y(SUM[16]) );
  XNOR2X4 U43 ( .A(B[16]), .B(A[16]), .Y(n14) );
  NAND2X1 U44 ( .A(n5), .B(n94), .Y(n124) );
  NAND2X1 U45 ( .A(A[14]), .B(B[14]), .Y(n109) );
  NAND2X2 U46 ( .A(n16), .B(n102), .Y(n117) );
  NOR2BX4 U47 ( .AN(n82), .B(n84), .Y(n83) );
  INVX4 U48 ( .A(n80), .Y(n84) );
  OR2X4 U49 ( .A(B[12]), .B(A[12]), .Y(n15) );
  NAND2X2 U50 ( .A(B[4]), .B(A[4]), .Y(n67) );
  CLKINVX8 U51 ( .A(n108), .Y(n16) );
  OR2X4 U52 ( .A(B[11]), .B(A[11]), .Y(n17) );
  XOR2X4 U53 ( .A(n21), .B(n18), .Y(n145) );
  NAND2X2 U54 ( .A(n17), .B(n93), .Y(n133) );
  NAND2BX4 U55 ( .AN(n55), .B(n137), .Y(n98) );
  NAND2X4 U56 ( .A(A[12]), .B(B[12]), .Y(n126) );
  BUFX20 U57 ( .A(n146), .Y(SUM[11]) );
  NAND2X4 U58 ( .A(n52), .B(n28), .Y(n29) );
  INVX4 U59 ( .A(n53), .Y(n28) );
  XNOR2X4 U60 ( .A(n115), .B(n114), .Y(n19) );
  NOR2BX4 U61 ( .AN(n71), .B(n72), .Y(n70) );
  NAND2X2 U62 ( .A(B[3]), .B(A[3]), .Y(n71) );
  INVX8 U63 ( .A(n110), .Y(n47) );
  INVX4 U64 ( .A(n64), .Y(n62) );
  NAND2X4 U65 ( .A(B[2]), .B(A[2]), .Y(n76) );
  INVXL U66 ( .A(A[14]), .Y(n25) );
  AOI21X4 U67 ( .A0(n129), .A1(n15), .B0(n130), .Y(n128) );
  NOR2X4 U68 ( .A(A[15]), .B(B[15]), .Y(n20) );
  AND2X4 U69 ( .A(n104), .B(n37), .Y(n40) );
  OAI21X2 U70 ( .A0(n105), .A1(n106), .B0(n107), .Y(n104) );
  BUFX20 U71 ( .A(n147), .Y(SUM[10]) );
  NAND2X4 U72 ( .A(B[13]), .B(A[13]), .Y(n119) );
  OAI21X4 U73 ( .A0(n117), .A1(n116), .B0(n109), .Y(n114) );
  AOI21X2 U74 ( .A0(n103), .A1(n129), .B0(n118), .Y(n116) );
  NAND2X2 U75 ( .A(B[7]), .B(A[7]), .Y(n54) );
  NAND2X4 U76 ( .A(n15), .B(n126), .Y(n21) );
  OAI2BB1X4 U77 ( .A0N(n22), .A1N(n23), .B0(n119), .Y(n121) );
  OR2X4 U78 ( .A(n124), .B(n125), .Y(n22) );
  INVX4 U79 ( .A(n126), .Y(n130) );
  INVXL U80 ( .A(B[14]), .Y(n24) );
  AOI2BB1X4 U81 ( .A0N(n24), .A1N(n25), .B0(n123), .Y(n122) );
  NOR2X2 U82 ( .A(n20), .B(n123), .Y(n107) );
  NAND2X4 U83 ( .A(B[6]), .B(A[6]), .Y(n58) );
  BUFX8 U84 ( .A(B[5]), .Y(n26) );
  NAND4BBX2 U85 ( .AN(n38), .BN(n39), .C(n61), .D(n140), .Y(n99) );
  OR2X4 U86 ( .A(A[7]), .B(B[7]), .Y(n140) );
  NAND3X4 U87 ( .A(n120), .B(n93), .C(n94), .Y(n129) );
  BUFX20 U88 ( .A(n144), .Y(SUM[13]) );
  BUFX20 U89 ( .A(n145), .Y(SUM[12]) );
  XOR2X4 U90 ( .A(n48), .B(n49), .Y(SUM[8]) );
  NAND2X2 U91 ( .A(B[8]), .B(A[8]), .Y(n50) );
  NOR2BX4 U92 ( .AN(n85), .B(n36), .Y(SUM[0]) );
  NAND2X4 U93 ( .A(B[0]), .B(A[0]), .Y(n85) );
  NAND2X2 U94 ( .A(n71), .B(n141), .Y(n96) );
  OAI211X2 U95 ( .A0(n142), .A1(n143), .B0(n79), .C0(n73), .Y(n141) );
  INVX8 U96 ( .A(n96), .Y(n66) );
  XOR2X4 U97 ( .A(n96), .B(n68), .Y(SUM[4]) );
  NOR2BX4 U98 ( .AN(n67), .B(n39), .Y(n68) );
  NOR2X2 U99 ( .A(A[4]), .B(B[4]), .Y(n39) );
  BUFX20 U100 ( .A(n35), .Y(SUM[14]) );
  INVX4 U101 ( .A(n61), .Y(n57) );
  OR2X4 U102 ( .A(A[6]), .B(B[6]), .Y(n61) );
  XOR2X4 U103 ( .A(n77), .B(n78), .Y(SUM[2]) );
  NOR2BX4 U104 ( .AN(n76), .B(n75), .Y(n78) );
  INVX4 U105 ( .A(n113), .Y(n51) );
  OR2X4 U106 ( .A(A[8]), .B(B[8]), .Y(n113) );
  NAND2X4 U107 ( .A(n26), .B(A[5]), .Y(n63) );
  NOR2X4 U108 ( .A(A[5]), .B(n26), .Y(n38) );
  NAND2X4 U109 ( .A(n27), .B(n53), .Y(n30) );
  NAND2X4 U110 ( .A(n29), .B(n30), .Y(n148) );
  NOR2BX4 U111 ( .AN(n54), .B(n55), .Y(n53) );
  NAND2X2 U112 ( .A(n100), .B(n119), .Y(n127) );
  OR2X4 U113 ( .A(B[13]), .B(A[13]), .Y(n100) );
  INVX8 U114 ( .A(n19), .Y(SUM[15]) );
  OR2X4 U115 ( .A(A[10]), .B(B[10]), .Y(n111) );
  OAI21X4 U116 ( .A0(n136), .A1(n47), .B0(n46), .Y(n135) );
  NAND2X4 U117 ( .A(B[11]), .B(A[11]), .Y(n93) );
  INVX4 U118 ( .A(n59), .Y(n56) );
  OAI21X4 U119 ( .A0(n66), .A1(n99), .B0(n98), .Y(n48) );
  XOR2X4 U120 ( .A(n69), .B(n70), .Y(SUM[3]) );
  INVXL U121 ( .A(n98), .Y(n97) );
  INVX4 U122 ( .A(n79), .Y(n75) );
  NAND2XL U123 ( .A(n113), .B(n110), .Y(n34) );
  OAI211X4 U124 ( .A0(n47), .A1(n50), .B0(n46), .C0(n132), .Y(n131) );
  XOR2X4 U125 ( .A(n127), .B(n128), .Y(n144) );
  OR2X4 U126 ( .A(A[3]), .B(B[3]), .Y(n73) );
  XOR2X4 U127 ( .A(n121), .B(n122), .Y(n35) );
  NOR2XL U128 ( .A(A[0]), .B(B[0]), .Y(n36) );
  NAND2XL U129 ( .A(B[15]), .B(A[15]), .Y(n37) );
  INVX1 U130 ( .A(n99), .Y(n95) );
  OAI21XL U131 ( .A0(n84), .A1(n85), .B0(n82), .Y(n142) );
  INVX1 U132 ( .A(n76), .Y(n143) );
  NAND3X1 U133 ( .A(n138), .B(n58), .C(n54), .Y(n137) );
  NAND3BX1 U134 ( .AN(n38), .B(n139), .C(n61), .Y(n138) );
  NAND2X1 U135 ( .A(n63), .B(n67), .Y(n139) );
  INVX1 U136 ( .A(n77), .Y(n74) );
  INVX1 U137 ( .A(n73), .Y(n72) );
  INVX1 U138 ( .A(n85), .Y(n81) );
  AOI21XL U139 ( .A0(n95), .A1(n96), .B0(n97), .Y(n90) );
  NAND2X1 U140 ( .A(B[1]), .B(A[1]), .Y(n82) );
  OR2X2 U141 ( .A(A[2]), .B(B[2]), .Y(n79) );
  OR2X2 U142 ( .A(A[1]), .B(B[1]), .Y(n80) );
  XOR2X4 U143 ( .A(n44), .B(n45), .Y(SUM[9]) );
  NOR2BX4 U144 ( .AN(n46), .B(n47), .Y(n45) );
  NOR2BX4 U145 ( .AN(n50), .B(n51), .Y(n49) );
  OAI21X4 U146 ( .A0(n56), .A1(n57), .B0(n58), .Y(n52) );
  XOR2X4 U147 ( .A(n59), .B(n60), .Y(n149) );
  NOR2BX4 U148 ( .AN(n58), .B(n57), .Y(n60) );
  OAI21X4 U149 ( .A0(n62), .A1(n38), .B0(n63), .Y(n59) );
  XOR2X4 U150 ( .A(n64), .B(n65), .Y(SUM[5]) );
  NOR2BX4 U151 ( .AN(n63), .B(n38), .Y(n65) );
  OAI21X4 U152 ( .A0(n39), .A1(n66), .B0(n67), .Y(n64) );
  XOR2X4 U153 ( .A(n81), .B(n83), .Y(SUM[1]) );
  NAND2X4 U154 ( .A(n40), .B(n87), .Y(n86) );
  OR2X4 U155 ( .A(B[14]), .B(A[14]), .Y(n102) );
  XOR2X4 U156 ( .A(n133), .B(n134), .Y(n146) );
  OR2X4 U157 ( .A(A[9]), .B(B[9]), .Y(n110) );
  CLKINVX3 U158 ( .A(n44), .Y(n136) );
  OAI2BB1X4 U159 ( .A0N(n113), .A1N(n48), .B0(n50), .Y(n44) );
endmodule


module butterfly_DW01_add_48 ( A, B, SUM );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  wire   n128, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127;

  INVX8 U2 ( .A(n6), .Y(n7) );
  OAI2BB1X1 U3 ( .A0N(A[12]), .A1N(B[12]), .B0(n101), .Y(n100) );
  INVX1 U4 ( .A(n81), .Y(n10) );
  AND2X2 U5 ( .A(n77), .B(n107), .Y(n4) );
  BUFX3 U6 ( .A(n107), .Y(n12) );
  OAI2BB1X1 U7 ( .A0N(n75), .A1N(n76), .B0(n4), .Y(n3) );
  INVX4 U8 ( .A(n124), .Y(n41) );
  AND2X4 U9 ( .A(n102), .B(n78), .Y(n1) );
  NAND2X4 U10 ( .A(n1), .B(n8), .Y(n105) );
  NOR2X2 U11 ( .A(B[12]), .B(A[12]), .Y(n15) );
  OAI21X2 U12 ( .A0(n59), .A1(n60), .B0(n61), .Y(n54) );
  INVX4 U13 ( .A(n65), .Y(n69) );
  INVX2 U14 ( .A(n91), .Y(n33) );
  OAI21X2 U15 ( .A0(n69), .A1(n70), .B0(n67), .Y(n126) );
  CLKINVX3 U16 ( .A(n61), .Y(n127) );
  NAND3X2 U17 ( .A(n122), .B(n44), .C(n40), .Y(n121) );
  AOI21X2 U18 ( .A0(n92), .A1(n116), .B0(n117), .Y(n115) );
  XOR2X4 U19 ( .A(n2), .B(n17), .Y(n29) );
  NAND2X2 U20 ( .A(n93), .B(n87), .Y(n2) );
  INVX2 U21 ( .A(n87), .Y(n6) );
  NAND3X4 U22 ( .A(n7), .B(n88), .C(n102), .Y(n99) );
  BUFX8 U23 ( .A(A[14]), .Y(n5) );
  NAND3X4 U24 ( .A(n102), .B(n88), .C(n7), .Y(n110) );
  AND2X4 U25 ( .A(n32), .B(n91), .Y(n31) );
  NOR2X2 U26 ( .A(n15), .B(n13), .Y(n104) );
  INVX4 U27 ( .A(n92), .Y(n119) );
  NAND2X2 U28 ( .A(A[10]), .B(B[10]), .Y(n114) );
  NAND2X2 U29 ( .A(B[11]), .B(A[11]), .Y(n87) );
  INVX8 U30 ( .A(n78), .Y(n111) );
  NOR2X4 U31 ( .A(n111), .B(n15), .Y(n112) );
  INVX4 U32 ( .A(n10), .Y(n11) );
  AND2X2 U33 ( .A(n7), .B(n88), .Y(n8) );
  DLY1X1 U34 ( .A(n88), .Y(n9) );
  AND2X4 U35 ( .A(n77), .B(n74), .Y(n96) );
  OAI211X4 U36 ( .A0(n33), .A1(n36), .B0(n32), .C0(n114), .Y(n113) );
  INVX4 U37 ( .A(n115), .Y(n17) );
  NOR2X2 U38 ( .A(A[13]), .B(B[13]), .Y(n13) );
  OAI21XL U39 ( .A0(n13), .A1(n78), .B0(n101), .Y(n75) );
  BUFX8 U40 ( .A(B[14]), .Y(n14) );
  INVX8 U41 ( .A(n90), .Y(n51) );
  NOR2BX4 U42 ( .AN(n67), .B(n69), .Y(n68) );
  NAND2X2 U43 ( .A(B[15]), .B(A[15]), .Y(n77) );
  NAND2X4 U44 ( .A(n76), .B(n107), .Y(n21) );
  NAND2X4 U45 ( .A(n14), .B(n5), .Y(n107) );
  NAND2X2 U46 ( .A(B[7]), .B(A[7]), .Y(n40) );
  AOI21X1 U47 ( .A0(n82), .A1(n110), .B0(n100), .Y(n97) );
  NOR2BX4 U48 ( .AN(n36), .B(n37), .Y(n35) );
  NAND2X4 U49 ( .A(B[8]), .B(A[8]), .Y(n36) );
  NOR2BX4 U50 ( .AN(n61), .B(n60), .Y(n63) );
  INVX8 U51 ( .A(n64), .Y(n60) );
  NAND2X4 U52 ( .A(A[12]), .B(B[12]), .Y(n78) );
  OR2X4 U53 ( .A(A[11]), .B(B[11]), .Y(n16) );
  INVX4 U54 ( .A(n94), .Y(n37) );
  NAND2X4 U55 ( .A(n81), .B(n101), .Y(n108) );
  NAND4X4 U56 ( .A(n93), .B(n34), .C(n92), .D(n22), .Y(n102) );
  NAND2X4 U57 ( .A(B[6]), .B(A[6]), .Y(n44) );
  NOR2BX2 U58 ( .AN(n70), .B(n20), .Y(SUM[0]) );
  NAND2X4 U59 ( .A(B[0]), .B(A[0]), .Y(n70) );
  INVX8 U60 ( .A(n29), .Y(SUM[11]) );
  NOR2X4 U61 ( .A(A[4]), .B(B[4]), .Y(n26) );
  INVX8 U62 ( .A(n18), .Y(SUM[4]) );
  NAND3X4 U63 ( .A(n16), .B(n113), .C(n92), .Y(n88) );
  NAND2X4 U64 ( .A(B[5]), .B(A[5]), .Y(n48) );
  NAND4BBX2 U65 ( .AN(n25), .BN(n26), .C(n47), .D(n124), .Y(n80) );
  NAND2X4 U66 ( .A(B[4]), .B(A[4]), .Y(n52) );
  OAI21X2 U67 ( .A0(n42), .A1(n43), .B0(n44), .Y(n38) );
  NOR2BX4 U68 ( .AN(n40), .B(n41), .Y(n39) );
  NOR2BX4 U69 ( .AN(n56), .B(n57), .Y(n55) );
  NAND2X2 U70 ( .A(B[9]), .B(A[9]), .Y(n32) );
  CLKINVX4 U71 ( .A(n25), .Y(n23) );
  NAND3BX1 U72 ( .AN(n25), .B(n123), .C(n47), .Y(n122) );
  NAND2X2 U73 ( .A(n48), .B(n52), .Y(n123) );
  INVX4 U74 ( .A(n45), .Y(n42) );
  INVX1 U75 ( .A(n101), .Y(n106) );
  CLKINVX2 U76 ( .A(n53), .Y(n19) );
  XOR2X2 U77 ( .A(n90), .B(n19), .Y(n18) );
  INVX2 U78 ( .A(n62), .Y(n59) );
  OAI21X4 U79 ( .A0(n120), .A1(n33), .B0(n32), .Y(n116) );
  NOR2XL U80 ( .A(A[0]), .B(B[0]), .Y(n20) );
  INVX2 U81 ( .A(n79), .Y(n85) );
  NAND2X1 U82 ( .A(B[3]), .B(A[3]), .Y(n56) );
  NAND2X2 U83 ( .A(B[1]), .B(A[1]), .Y(n67) );
  XNOR2X4 U84 ( .A(n21), .B(n103), .Y(n27) );
  INVX1 U85 ( .A(n70), .Y(n66) );
  AND2X1 U86 ( .A(n94), .B(n91), .Y(n22) );
  OAI2BB1X4 U87 ( .A0N(n49), .A1N(n23), .B0(n48), .Y(n45) );
  XNOR2X4 U88 ( .A(n109), .B(n108), .Y(n24) );
  INVX8 U89 ( .A(n24), .Y(SUM[13]) );
  NOR2BX1 U90 ( .AN(n52), .B(n26), .Y(n53) );
  INVX1 U91 ( .A(n114), .Y(n117) );
  INVXL U92 ( .A(n58), .Y(n57) );
  OAI2BB1X1 U93 ( .A0N(n65), .A1N(n66), .B0(n67), .Y(n62) );
  NOR2X4 U94 ( .A(A[5]), .B(B[5]), .Y(n25) );
  NOR2X2 U95 ( .A(n84), .B(n83), .Y(n73) );
  AOI21X2 U96 ( .A0(n85), .A1(n34), .B0(n86), .Y(n83) );
  INVX8 U97 ( .A(n27), .Y(SUM[14]) );
  BUFX20 U98 ( .A(n128), .Y(SUM[15]) );
  NAND2XL U99 ( .A(n7), .B(n9), .Y(n86) );
  NAND4BXL U100 ( .AN(n37), .B(n91), .C(n92), .D(n16), .Y(n79) );
  NAND3XL U101 ( .A(n11), .B(n76), .C(n82), .Y(n84) );
  NAND2X2 U102 ( .A(n76), .B(n11), .Y(n98) );
  XOR2X4 U103 ( .A(n30), .B(n31), .Y(SUM[9]) );
  XOR2X4 U104 ( .A(n34), .B(n35), .Y(SUM[8]) );
  XOR2X4 U105 ( .A(n38), .B(n39), .Y(SUM[7]) );
  XOR2X4 U106 ( .A(n45), .B(n46), .Y(SUM[6]) );
  NOR2BX4 U107 ( .AN(n44), .B(n43), .Y(n46) );
  CLKINVX3 U108 ( .A(n47), .Y(n43) );
  XOR2X4 U109 ( .A(n49), .B(n50), .Y(SUM[5]) );
  NOR2BX4 U110 ( .AN(n48), .B(n25), .Y(n50) );
  OAI21X4 U111 ( .A0(n26), .A1(n51), .B0(n52), .Y(n49) );
  XOR2X4 U112 ( .A(n54), .B(n55), .Y(SUM[3]) );
  XOR2X4 U113 ( .A(n62), .B(n63), .Y(SUM[2]) );
  XOR2X4 U114 ( .A(n66), .B(n68), .Y(SUM[1]) );
  XOR2X4 U115 ( .A(n72), .B(n71), .Y(SUM[16]) );
  XNOR2X4 U116 ( .A(B[16]), .B(A[16]), .Y(n72) );
  OAI21X4 U117 ( .A0(n73), .A1(n3), .B0(n74), .Y(n71) );
  XOR2X4 U118 ( .A(n95), .B(n96), .Y(n128) );
  OR2X4 U119 ( .A(B[15]), .B(A[15]), .Y(n74) );
  OAI21X4 U120 ( .A0(n98), .A1(n97), .B0(n12), .Y(n95) );
  NAND2X4 U121 ( .A(A[13]), .B(B[13]), .Y(n101) );
  AOI21X4 U122 ( .A0(n104), .A1(n105), .B0(n106), .Y(n103) );
  OR2X4 U123 ( .A(A[14]), .B(B[14]), .Y(n76) );
  AOI21X4 U124 ( .A0(n82), .A1(n99), .B0(n111), .Y(n109) );
  OR2X4 U125 ( .A(A[13]), .B(B[13]), .Y(n81) );
  XOR2X4 U126 ( .A(n112), .B(n110), .Y(SUM[12]) );
  OR2X4 U127 ( .A(A[12]), .B(B[12]), .Y(n82) );
  OR2X4 U128 ( .A(B[11]), .B(A[11]), .Y(n93) );
  XOR2X4 U129 ( .A(n118), .B(n116), .Y(SUM[10]) );
  NOR2BX4 U130 ( .AN(n114), .B(n119), .Y(n118) );
  OR2X4 U131 ( .A(A[10]), .B(B[10]), .Y(n92) );
  OR2X4 U132 ( .A(A[9]), .B(B[9]), .Y(n91) );
  CLKINVX3 U133 ( .A(n30), .Y(n120) );
  OAI2BB1X4 U134 ( .A0N(n94), .A1N(n34), .B0(n36), .Y(n30) );
  OAI21X4 U135 ( .A0(n51), .A1(n80), .B0(n89), .Y(n34) );
  NAND2BX4 U136 ( .AN(n41), .B(n121), .Y(n89) );
  OR2X4 U137 ( .A(A[7]), .B(B[7]), .Y(n124) );
  OR2X4 U138 ( .A(A[6]), .B(B[6]), .Y(n47) );
  NAND2X4 U139 ( .A(n56), .B(n125), .Y(n90) );
  OAI211X2 U140 ( .A0(n126), .A1(n127), .B0(n64), .C0(n58), .Y(n125) );
  OR2X4 U141 ( .A(A[3]), .B(B[3]), .Y(n58) );
  OR2X4 U142 ( .A(A[2]), .B(B[2]), .Y(n64) );
  NAND2X4 U143 ( .A(B[2]), .B(A[2]), .Y(n61) );
  OR2X4 U144 ( .A(A[1]), .B(B[1]), .Y(n65) );
  OR2X4 U145 ( .A(A[8]), .B(B[8]), .Y(n94) );
endmodule


module butterfly_DW01_add_50 ( A, B, SUM );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  wire   n138, n139, n140, n141, n142, n143, n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n13, n14, n15, n16, n19, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137;

  NAND2X2 U2 ( .A(n11), .B(n99), .Y(n97) );
  OR2X4 U3 ( .A(A[11]), .B(B[11]), .Y(n1) );
  CLKBUFX8 U4 ( .A(n113), .Y(n4) );
  NAND2X2 U5 ( .A(n24), .B(n78), .Y(n77) );
  INVX3 U6 ( .A(n119), .Y(n2) );
  CLKINVX4 U7 ( .A(n2), .Y(n3) );
  NOR3X4 U8 ( .A(n112), .B(n4), .C(n105), .Y(n109) );
  AND2X4 U9 ( .A(n83), .B(n5), .Y(n81) );
  BUFX8 U10 ( .A(n82), .Y(n5) );
  INVX2 U11 ( .A(n85), .Y(n55) );
  BUFX20 U12 ( .A(n142), .Y(SUM[9]) );
  INVX3 U13 ( .A(n103), .Y(n120) );
  XOR2X4 U14 ( .A(n6), .B(n118), .Y(n139) );
  NAND2X2 U15 ( .A(n89), .B(n102), .Y(n6) );
  OR2X4 U16 ( .A(A[12]), .B(B[12]), .Y(n7) );
  INVX2 U17 ( .A(B[15]), .Y(n8) );
  CLKINVX4 U18 ( .A(n8), .Y(n9) );
  CLKINVX3 U19 ( .A(n104), .Y(n15) );
  INVX2 U20 ( .A(n102), .Y(n116) );
  INVX8 U21 ( .A(n91), .Y(n104) );
  CLKINVX4 U22 ( .A(n33), .Y(n130) );
  NAND4BBX2 U23 ( .AN(n29), .BN(n30), .C(n50), .D(n134), .Y(n88) );
  NOR2BX4 U24 ( .AN(n43), .B(n44), .Y(n42) );
  BUFX20 U25 ( .A(n143), .Y(SUM[7]) );
  BUFX8 U26 ( .A(n110), .Y(n10) );
  XOR2X4 U27 ( .A(A[16]), .B(B[16]), .Y(n75) );
  INVX8 U28 ( .A(n98), .Y(n11) );
  NOR2X2 U29 ( .A(B[14]), .B(A[14]), .Y(n112) );
  INVX4 U30 ( .A(n106), .Y(n98) );
  INVXL U31 ( .A(n105), .Y(n16) );
  INVX1 U32 ( .A(n123), .Y(n127) );
  BUFX20 U33 ( .A(n139), .Y(SUM[13]) );
  BUFX12 U34 ( .A(n94), .Y(n13) );
  NOR2X2 U35 ( .A(n112), .B(n105), .Y(n100) );
  OR2X4 U36 ( .A(A[6]), .B(B[6]), .Y(n50) );
  NAND2X4 U37 ( .A(B[12]), .B(A[12]), .Y(n103) );
  INVX3 U38 ( .A(n57), .Y(n22) );
  NAND2X2 U39 ( .A(B[4]), .B(A[4]), .Y(n56) );
  INVX8 U40 ( .A(n89), .Y(n105) );
  XOR2X4 U41 ( .A(n14), .B(n75), .Y(SUM[16]) );
  NAND2X4 U42 ( .A(n76), .B(n77), .Y(n14) );
  NAND2X2 U43 ( .A(B[6]), .B(A[6]), .Y(n47) );
  BUFX20 U44 ( .A(n141), .Y(SUM[10]) );
  NAND2X4 U45 ( .A(n5), .B(n1), .Y(n124) );
  XOR2X4 U46 ( .A(n58), .B(n59), .Y(SUM[3]) );
  OAI21X1 U47 ( .A0(n63), .A1(n64), .B0(n65), .Y(n58) );
  NAND2X2 U48 ( .A(n106), .B(n91), .Y(n23) );
  INVX4 U49 ( .A(n134), .Y(n44) );
  NAND2X2 U50 ( .A(B[7]), .B(A[7]), .Y(n43) );
  INVX8 U51 ( .A(n93), .Y(n36) );
  BUFX20 U52 ( .A(n138), .Y(SUM[14]) );
  NAND2X2 U53 ( .A(B[11]), .B(A[11]), .Y(n82) );
  OAI2BB1X4 U54 ( .A0N(A[15]), .A1N(n9), .B0(n90), .Y(n107) );
  AND4X2 U55 ( .A(n16), .B(n90), .C(n15), .D(n7), .Y(n24) );
  NOR2BX4 U56 ( .AN(n71), .B(n73), .Y(n72) );
  INVX2 U57 ( .A(n69), .Y(n73) );
  AOI21X4 U58 ( .A0(n13), .A1(n126), .B0(n127), .Y(n125) );
  AND2X1 U59 ( .A(n9), .B(A[15]), .Y(n26) );
  NOR2X2 U60 ( .A(A[4]), .B(B[4]), .Y(n30) );
  NAND2X2 U61 ( .A(B[1]), .B(A[1]), .Y(n71) );
  OAI211X4 U62 ( .A0(n36), .A1(n39), .B0(n35), .C0(n123), .Y(n122) );
  NAND2X4 U63 ( .A(A[13]), .B(B[13]), .Y(n102) );
  NOR2BX4 U64 ( .AN(n74), .B(n25), .Y(SUM[0]) );
  NAND2X4 U65 ( .A(B[0]), .B(A[0]), .Y(n74) );
  NAND2BX2 U66 ( .AN(n44), .B(n131), .Y(n87) );
  XOR2X4 U67 ( .A(n66), .B(n67), .Y(SUM[2]) );
  NOR2BX4 U68 ( .AN(n65), .B(n64), .Y(n67) );
  NAND2X2 U69 ( .A(B[10]), .B(A[10]), .Y(n123) );
  NAND4BX4 U70 ( .AN(n21), .B(n95), .C(n13), .D(n37), .Y(n117) );
  INVX8 U71 ( .A(n92), .Y(n113) );
  NAND2X4 U72 ( .A(B[9]), .B(A[9]), .Y(n35) );
  NOR2BX2 U73 ( .AN(n60), .B(n61), .Y(n59) );
  INVX8 U74 ( .A(n28), .Y(SUM[15]) );
  NAND2X2 U75 ( .A(n100), .B(n101), .Y(n99) );
  OR2X4 U76 ( .A(A[8]), .B(B[8]), .Y(n96) );
  NAND2X4 U77 ( .A(B[8]), .B(A[8]), .Y(n39) );
  AND2X4 U78 ( .A(n97), .B(n90), .Y(n19) );
  NOR2X4 U79 ( .A(n19), .B(n26), .Y(n76) );
  OR2X4 U80 ( .A(A[10]), .B(B[10]), .Y(n94) );
  BUFX20 U81 ( .A(n140), .Y(SUM[12]) );
  CLKINVX2 U82 ( .A(n65), .Y(n137) );
  OAI21X1 U83 ( .A0(n73), .A1(n74), .B0(n71), .Y(n136) );
  NAND3XL U84 ( .A(n132), .B(n47), .C(n43), .Y(n131) );
  NAND3BXL U85 ( .AN(n29), .B(n133), .C(n50), .Y(n132) );
  XNOR2X4 U86 ( .A(n85), .B(n22), .Y(SUM[4]) );
  OAI2BB1X2 U87 ( .A0N(n69), .A1N(n70), .B0(n71), .Y(n66) );
  INVX2 U88 ( .A(n62), .Y(n61) );
  XOR2X4 U89 ( .A(n126), .B(n128), .Y(n141) );
  INVX4 U90 ( .A(n96), .Y(n40) );
  INVX4 U91 ( .A(n50), .Y(n46) );
  NOR2X4 U92 ( .A(A[5]), .B(B[5]), .Y(n29) );
  NAND2X1 U93 ( .A(B[3]), .B(A[3]), .Y(n60) );
  NAND2X2 U94 ( .A(B[5]), .B(A[5]), .Y(n52) );
  NAND2X1 U95 ( .A(B[2]), .B(A[2]), .Y(n65) );
  INVXL U96 ( .A(n88), .Y(n84) );
  NOR2BX4 U97 ( .AN(n123), .B(n129), .Y(n128) );
  INVX4 U98 ( .A(n94), .Y(n129) );
  NAND2XL U99 ( .A(n96), .B(n93), .Y(n21) );
  NAND2XL U100 ( .A(n52), .B(n56), .Y(n133) );
  OAI21X4 U101 ( .A0(n130), .A1(n36), .B0(n35), .Y(n126) );
  XOR2X4 U102 ( .A(n114), .B(n23), .Y(n138) );
  OR2X4 U103 ( .A(A[2]), .B(B[2]), .Y(n68) );
  NOR2XL U104 ( .A(A[0]), .B(B[0]), .Y(n25) );
  OR2X4 U105 ( .A(A[12]), .B(B[12]), .Y(n92) );
  INVXL U106 ( .A(n87), .Y(n86) );
  XNOR2X4 U107 ( .A(n124), .B(n125), .Y(n27) );
  INVX8 U108 ( .A(n27), .Y(SUM[11]) );
  NAND4BXL U109 ( .AN(n40), .B(n93), .C(n13), .D(n1), .Y(n80) );
  INVX1 U110 ( .A(n66), .Y(n63) );
  NOR2BX1 U111 ( .AN(n56), .B(n30), .Y(n57) );
  INVX1 U112 ( .A(n68), .Y(n64) );
  INVX1 U113 ( .A(n74), .Y(n70) );
  XNOR2X4 U114 ( .A(n107), .B(n108), .Y(n28) );
  NAND2XL U115 ( .A(n102), .B(n103), .Y(n101) );
  OAI21XL U116 ( .A0(n79), .A1(n80), .B0(n81), .Y(n78) );
  AOI21XL U117 ( .A0(n84), .A1(n85), .B0(n86), .Y(n79) );
  OR2X2 U118 ( .A(A[1]), .B(B[1]), .Y(n69) );
  NAND3X4 U119 ( .A(n81), .B(n117), .C(n103), .Y(n110) );
  NAND2X2 U120 ( .A(B[14]), .B(A[14]), .Y(n106) );
  XOR2X4 U121 ( .A(n33), .B(n34), .Y(n142) );
  NOR2BX4 U122 ( .AN(n35), .B(n36), .Y(n34) );
  XOR2X4 U123 ( .A(n37), .B(n38), .Y(SUM[8]) );
  NOR2BX4 U124 ( .AN(n39), .B(n40), .Y(n38) );
  XOR2X4 U125 ( .A(n41), .B(n42), .Y(n143) );
  OAI21X4 U126 ( .A0(n45), .A1(n46), .B0(n47), .Y(n41) );
  CLKINVX3 U127 ( .A(n48), .Y(n45) );
  XOR2X4 U128 ( .A(n48), .B(n49), .Y(SUM[6]) );
  NOR2BX4 U129 ( .AN(n47), .B(n46), .Y(n49) );
  OAI21X4 U130 ( .A0(n51), .A1(n29), .B0(n52), .Y(n48) );
  CLKINVX3 U131 ( .A(n53), .Y(n51) );
  XOR2X4 U132 ( .A(n53), .B(n54), .Y(SUM[5]) );
  NOR2BX4 U133 ( .AN(n52), .B(n29), .Y(n54) );
  OAI21X4 U134 ( .A0(n30), .A1(n55), .B0(n56), .Y(n53) );
  XOR2X4 U135 ( .A(n70), .B(n72), .Y(SUM[1]) );
  AOI21X4 U136 ( .A0(n10), .A1(n109), .B0(n111), .Y(n108) );
  OAI21X4 U137 ( .A0(n104), .A1(n102), .B0(n11), .Y(n111) );
  OR2X4 U138 ( .A(B[15]), .B(A[15]), .Y(n90) );
  AOI21X4 U139 ( .A0(n115), .A1(n110), .B0(n116), .Y(n114) );
  NOR2X4 U140 ( .A(n105), .B(n4), .Y(n115) );
  OR2X4 U141 ( .A(B[14]), .B(A[14]), .Y(n91) );
  AOI21X4 U142 ( .A0(n119), .A1(n7), .B0(n120), .Y(n118) );
  OR2X4 U143 ( .A(B[13]), .B(A[13]), .Y(n89) );
  XOR2X4 U144 ( .A(n3), .B(n121), .Y(n140) );
  NOR2BX4 U145 ( .AN(n103), .B(n113), .Y(n121) );
  NAND3X4 U146 ( .A(n117), .B(n5), .C(n83), .Y(n119) );
  NAND3X4 U147 ( .A(n122), .B(n95), .C(n13), .Y(n83) );
  OR2X4 U148 ( .A(A[11]), .B(B[11]), .Y(n95) );
  OR2X4 U149 ( .A(A[9]), .B(B[9]), .Y(n93) );
  OAI2BB1X4 U150 ( .A0N(n96), .A1N(n37), .B0(n39), .Y(n33) );
  OAI21X4 U151 ( .A0(n55), .A1(n88), .B0(n87), .Y(n37) );
  OR2X4 U152 ( .A(A[7]), .B(B[7]), .Y(n134) );
  NAND2X4 U153 ( .A(n60), .B(n135), .Y(n85) );
  OAI211X2 U154 ( .A0(n136), .A1(n137), .B0(n68), .C0(n62), .Y(n135) );
  OR2X4 U155 ( .A(A[3]), .B(B[3]), .Y(n62) );
endmodule


module butterfly_DW01_add_61 ( A, B, SUM );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130;

  NAND3X1 U2 ( .A(n77), .B(n84), .C(n78), .Y(n81) );
  NAND2X2 U3 ( .A(B[10]), .B(A[10]), .Y(n117) );
  NAND2X4 U4 ( .A(B[4]), .B(A[4]), .Y(n42) );
  NOR2X2 U5 ( .A(A[4]), .B(B[4]), .Y(n18) );
  INVX4 U6 ( .A(n98), .Y(n100) );
  XOR2X4 U7 ( .A(n106), .B(n1), .Y(SUM[12]) );
  AND2X4 U8 ( .A(n5), .B(n85), .Y(n1) );
  INVX8 U9 ( .A(n117), .Y(n116) );
  NAND2X2 U10 ( .A(B[12]), .B(A[12]), .Y(n85) );
  OR2X2 U11 ( .A(A[12]), .B(B[12]), .Y(n5) );
  NOR2BX2 U12 ( .AN(n35), .B(n34), .Y(n37) );
  NAND2X2 U13 ( .A(n78), .B(n77), .Y(n88) );
  INVX1 U14 ( .A(A[15]), .Y(n3) );
  OAI21X2 U15 ( .A0(n18), .A1(n125), .B0(n42), .Y(n40) );
  NAND3X1 U16 ( .A(n77), .B(n78), .C(n79), .Y(n66) );
  OR2X4 U17 ( .A(A[5]), .B(B[5]), .Y(n2) );
  XOR2X2 U18 ( .A(n36), .B(n37), .Y(SUM[6]) );
  CLKINVX8 U19 ( .A(n70), .Y(n80) );
  NOR2BX4 U20 ( .AN(n21), .B(n22), .Y(n20) );
  OAI21X4 U21 ( .A0(n33), .A1(n34), .B0(n35), .Y(n28) );
  NAND2X2 U22 ( .A(B[6]), .B(A[6]), .Y(n35) );
  NAND3X4 U23 ( .A(n23), .B(n80), .C(n5), .Y(n90) );
  NAND2X4 U24 ( .A(n23), .B(n27), .Y(n121) );
  OAI2BB1X4 U25 ( .A0N(n23), .A1N(n80), .B0(n71), .Y(n106) );
  OR2X2 U26 ( .A(A[12]), .B(B[12]), .Y(n4) );
  INVX4 U27 ( .A(n96), .Y(n105) );
  NAND2X2 U28 ( .A(n4), .B(n96), .Y(n95) );
  NAND2BX4 U29 ( .AN(n105), .B(n107), .Y(n71) );
  AND2X2 U30 ( .A(B[11]), .B(A[11]), .Y(n14) );
  INVX2 U31 ( .A(n79), .Y(n83) );
  INVX2 U32 ( .A(n112), .Y(n119) );
  AOI21X2 U33 ( .A0(n81), .A1(n82), .B0(n83), .Y(n63) );
  NOR3BX4 U34 ( .AN(n90), .B(n91), .C(n92), .Y(n89) );
  OR2X4 U35 ( .A(A[12]), .B(B[12]), .Y(n68) );
  NAND2BX4 U36 ( .AN(B[15]), .B(n3), .Y(n79) );
  NAND3BX4 U37 ( .AN(n63), .B(n65), .C(n64), .Y(n61) );
  INVX4 U38 ( .A(n86), .Y(n6) );
  XOR2X2 U39 ( .A(n23), .B(n24), .Y(SUM[8]) );
  NOR2BX2 U40 ( .AN(n25), .B(n26), .Y(n24) );
  NAND2X4 U41 ( .A(B[8]), .B(A[8]), .Y(n25) );
  OR2X4 U42 ( .A(A[3]), .B(B[3]), .Y(n126) );
  XOR2X2 U43 ( .A(n40), .B(n41), .Y(SUM[5]) );
  NAND2X2 U44 ( .A(n94), .B(n15), .Y(n107) );
  XOR2X2 U45 ( .A(B[16]), .B(A[16]), .Y(n62) );
  INVX8 U46 ( .A(n111), .Y(n22) );
  NAND2X4 U47 ( .A(B[9]), .B(A[9]), .Y(n21) );
  NAND3BX4 U48 ( .AN(n66), .B(n67), .C(n11), .Y(n65) );
  NAND2X4 U49 ( .A(n121), .B(n25), .Y(n19) );
  AOI21X2 U50 ( .A0(n21), .A1(n25), .B0(n22), .Y(n108) );
  NAND2X2 U51 ( .A(n94), .B(n15), .Y(n103) );
  NAND2X2 U52 ( .A(n93), .B(n12), .Y(n92) );
  INVX4 U53 ( .A(n93), .Y(n99) );
  AND2X4 U54 ( .A(n93), .B(n78), .Y(n16) );
  NAND2X4 U55 ( .A(B[13]), .B(A[13]), .Y(n93) );
  NAND2X2 U56 ( .A(n87), .B(n86), .Y(n8) );
  NAND2X4 U57 ( .A(n7), .B(n6), .Y(n9) );
  NAND2X4 U58 ( .A(n8), .B(n9), .Y(SUM[15]) );
  INVX4 U59 ( .A(n87), .Y(n7) );
  OAI21X4 U60 ( .A0(n88), .A1(n89), .B0(n82), .Y(n86) );
  NAND2X4 U61 ( .A(n64), .B(n79), .Y(n87) );
  OAI21X2 U62 ( .A0(A[11]), .A1(B[11]), .B0(n112), .Y(n109) );
  INVX8 U63 ( .A(n2), .Y(n10) );
  BUFX2 U64 ( .A(n4), .Y(n11) );
  INVX4 U65 ( .A(n104), .Y(n12) );
  CLKINVX8 U66 ( .A(n85), .Y(n104) );
  OR2X4 U67 ( .A(A[9]), .B(B[9]), .Y(n111) );
  XOR2X4 U68 ( .A(n19), .B(n20), .Y(SUM[9]) );
  NOR2BX4 U69 ( .AN(n117), .B(n119), .Y(n118) );
  XOR2X4 U70 ( .A(n118), .B(n115), .Y(SUM[10]) );
  XOR2X4 U71 ( .A(n97), .B(n13), .Y(SUM[14]) );
  NAND2X4 U72 ( .A(n82), .B(n77), .Y(n13) );
  AOI21X4 U73 ( .A0(n112), .A1(n115), .B0(n116), .Y(n114) );
  NAND2X2 U74 ( .A(B[14]), .B(A[14]), .Y(n82) );
  NOR2X2 U75 ( .A(n129), .B(n130), .Y(n127) );
  OAI21X1 U76 ( .A0(n59), .A1(n60), .B0(n57), .Y(n130) );
  INVX2 U77 ( .A(n36), .Y(n33) );
  NAND2X2 U78 ( .A(n96), .B(n15), .Y(n113) );
  NOR2BX4 U79 ( .AN(n68), .B(n105), .Y(n102) );
  OR2X4 U80 ( .A(B[13]), .B(A[13]), .Y(n78) );
  NAND2X2 U81 ( .A(B[5]), .B(A[5]), .Y(n39) );
  OR2X2 U82 ( .A(A[11]), .B(B[11]), .Y(n96) );
  XOR2X4 U83 ( .A(n113), .B(n114), .Y(SUM[11]) );
  XOR2X4 U84 ( .A(n28), .B(n29), .Y(SUM[7]) );
  AOI21X2 U85 ( .A0(n94), .A1(n15), .B0(n95), .Y(n91) );
  AOI21X4 U86 ( .A0(n102), .A1(n103), .B0(n104), .Y(n101) );
  OAI21X4 U87 ( .A0(n122), .A1(n123), .B0(n32), .Y(n75) );
  NAND2X1 U88 ( .A(B[7]), .B(A[7]), .Y(n30) );
  XOR2X4 U89 ( .A(n61), .B(n62), .Y(SUM[16]) );
  AOI211X2 U90 ( .A0(n39), .A1(n42), .B0(n34), .C0(n10), .Y(n122) );
  OR2X4 U91 ( .A(A[10]), .B(B[10]), .Y(n112) );
  OAI21X4 U92 ( .A0(n116), .A1(n108), .B0(n112), .Y(n94) );
  NAND4BBX2 U93 ( .AN(n10), .BN(n18), .C(n124), .D(n32), .Y(n76) );
  NAND2X2 U94 ( .A(B[15]), .B(A[15]), .Y(n64) );
  INVX4 U95 ( .A(n14), .Y(n15) );
  OR2X4 U96 ( .A(A[14]), .B(B[14]), .Y(n77) );
  OAI21X4 U97 ( .A0(n38), .A1(n10), .B0(n39), .Y(n36) );
  INVX4 U98 ( .A(n40), .Y(n38) );
  NOR2BX2 U99 ( .AN(n39), .B(n10), .Y(n41) );
  INVX2 U100 ( .A(n19), .Y(n120) );
  NAND2XL U101 ( .A(B[3]), .B(A[3]), .Y(n47) );
  NAND2XL U102 ( .A(B[1]), .B(A[1]), .Y(n57) );
  OR2XL U103 ( .A(A[1]), .B(B[1]), .Y(n55) );
  NAND2XL U104 ( .A(B[0]), .B(A[0]), .Y(n60) );
  OAI21X4 U105 ( .A0(n125), .A1(n76), .B0(n75), .Y(n23) );
  XNOR2X4 U106 ( .A(n100), .B(n16), .Y(SUM[13]) );
  OAI21X4 U107 ( .A0(n120), .A1(n22), .B0(n21), .Y(n115) );
  OAI21X4 U108 ( .A0(n127), .A1(n128), .B0(n47), .Y(n73) );
  NAND2X2 U109 ( .A(n30), .B(n35), .Y(n123) );
  INVX4 U110 ( .A(n124), .Y(n34) );
  AOI21XL U111 ( .A0(n72), .A1(n73), .B0(n74), .Y(n69) );
  CLKINVX3 U112 ( .A(n51), .Y(n129) );
  XOR2X1 U113 ( .A(n45), .B(n46), .Y(SUM[3]) );
  OAI21XL U114 ( .A0(n49), .A1(n50), .B0(n51), .Y(n45) );
  NOR2BX2 U115 ( .AN(n47), .B(n48), .Y(n46) );
  OAI2BB1X2 U116 ( .A0N(n55), .A1N(n56), .B0(n57), .Y(n52) );
  NOR2BX1 U117 ( .AN(n51), .B(n50), .Y(n53) );
  XOR2X1 U118 ( .A(n56), .B(n58), .Y(SUM[1]) );
  OR2XL U119 ( .A(A[2]), .B(B[2]), .Y(n54) );
  NOR2BX1 U120 ( .AN(n60), .B(n17), .Y(SUM[0]) );
  NOR2XL U121 ( .A(A[0]), .B(B[0]), .Y(n17) );
  INVX1 U122 ( .A(n125), .Y(n43) );
  INVX1 U123 ( .A(n73), .Y(n125) );
  NAND2X1 U124 ( .A(n12), .B(n93), .Y(n84) );
  INVX1 U125 ( .A(n27), .Y(n26) );
  NOR2BX2 U126 ( .AN(n30), .B(n31), .Y(n29) );
  INVXL U127 ( .A(n32), .Y(n31) );
  OAI21XL U128 ( .A0(n69), .A1(n70), .B0(n71), .Y(n67) );
  INVXL U129 ( .A(n76), .Y(n72) );
  INVXL U130 ( .A(n75), .Y(n74) );
  NAND2X1 U131 ( .A(n54), .B(n126), .Y(n128) );
  INVX1 U132 ( .A(n55), .Y(n59) );
  INVX1 U133 ( .A(n54), .Y(n50) );
  INVX1 U134 ( .A(n52), .Y(n49) );
  XOR2X1 U135 ( .A(n43), .B(n44), .Y(SUM[4]) );
  NOR2BX1 U136 ( .AN(n42), .B(n18), .Y(n44) );
  XOR2X2 U137 ( .A(n52), .B(n53), .Y(SUM[2]) );
  INVX1 U138 ( .A(n126), .Y(n48) );
  NOR2BXL U139 ( .AN(n57), .B(n59), .Y(n58) );
  INVX1 U140 ( .A(n60), .Y(n56) );
  NAND2XL U141 ( .A(n111), .B(n27), .Y(n110) );
  NAND2X2 U142 ( .A(B[2]), .B(A[2]), .Y(n51) );
  AOI21X4 U143 ( .A0(n98), .A1(n78), .B0(n99), .Y(n97) );
  NAND2X4 U144 ( .A(n101), .B(n90), .Y(n98) );
  OR2X4 U145 ( .A(n109), .B(n110), .Y(n70) );
  OR2X4 U146 ( .A(A[8]), .B(B[8]), .Y(n27) );
  OR2X4 U147 ( .A(A[7]), .B(B[7]), .Y(n32) );
  OR2X4 U148 ( .A(A[6]), .B(B[6]), .Y(n124) );
endmodule


module butterfly_DW01_sub_57 ( A, B, DIFF );
  input [16:0] A;
  input [16:0] B;
  output [16:0] DIFF;
  wire   n153, n1, n2, n3, n4, n5, n6, n8, n9, n10, n11, n12, n13, n14, n16,
         n17, n18, n19, n20, n21, n22, n23, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152;

  BUFX2 U3 ( .A(n101), .Y(n5) );
  INVX3 U4 ( .A(n101), .Y(n114) );
  CLKINVX8 U5 ( .A(n2), .Y(n1) );
  INVX8 U6 ( .A(n94), .Y(n2) );
  INVX8 U7 ( .A(n2), .Y(n3) );
  CLKINVX4 U8 ( .A(n100), .Y(n110) );
  INVX1 U9 ( .A(n104), .Y(n23) );
  INVX8 U10 ( .A(n106), .Y(n18) );
  NAND2X4 U11 ( .A(n97), .B(n21), .Y(n84) );
  INVX8 U12 ( .A(A[15]), .Y(n97) );
  CLKINVX3 U13 ( .A(n135), .Y(n13) );
  INVX4 U14 ( .A(n146), .Y(n50) );
  NAND2BX4 U15 ( .AN(A[5]), .B(B[5]), .Y(n146) );
  XNOR2X4 U16 ( .A(n4), .B(n122), .Y(DIFF[12]) );
  NAND2X2 U17 ( .A(n116), .B(n120), .Y(n4) );
  XOR2X4 U18 ( .A(n8), .B(n113), .Y(n6) );
  BUFX16 U19 ( .A(n153), .Y(DIFF[13]) );
  XOR2X2 U20 ( .A(n26), .B(n118), .Y(n153) );
  BUFX12 U21 ( .A(B[15]), .Y(n21) );
  NOR2X4 U22 ( .A(n9), .B(n17), .Y(n8) );
  AND3X4 U23 ( .A(n116), .B(n3), .C(n117), .Y(n9) );
  INVX4 U24 ( .A(n112), .Y(n10) );
  INVX8 U25 ( .A(n93), .Y(n112) );
  NAND2BX4 U26 ( .AN(A[10]), .B(B[10]), .Y(n128) );
  NAND2X2 U27 ( .A(n11), .B(n1), .Y(n115) );
  INVX2 U28 ( .A(n131), .Y(n129) );
  AND2X4 U29 ( .A(A[12]), .B(n105), .Y(n11) );
  NOR2BX4 U30 ( .AN(A[10]), .B(B[10]), .Y(n130) );
  NAND2BX4 U31 ( .AN(B[10]), .B(A[10]), .Y(n139) );
  INVX2 U32 ( .A(n128), .Y(n138) );
  INVX2 U33 ( .A(n139), .Y(n141) );
  NOR2BX2 U34 ( .AN(B[10]), .B(A[10]), .Y(n132) );
  XNOR2X4 U35 ( .A(n143), .B(n35), .Y(DIFF[8]) );
  INVX4 U36 ( .A(n127), .Y(n32) );
  OAI21X4 U37 ( .A0(n142), .A1(n32), .B0(n33), .Y(n140) );
  NOR2X2 U38 ( .A(n36), .B(n37), .Y(n35) );
  INVX2 U39 ( .A(n140), .Y(n137) );
  NOR2X2 U40 ( .A(n31), .B(n32), .Y(n30) );
  OAI21X2 U41 ( .A0(n49), .A1(n50), .B0(n51), .Y(n42) );
  INVX4 U42 ( .A(n92), .Y(n98) );
  XNOR2X4 U43 ( .A(n140), .B(n12), .Y(DIFF[10]) );
  OR2X4 U44 ( .A(n138), .B(n141), .Y(n12) );
  XNOR2X4 U45 ( .A(n134), .B(n13), .Y(DIFF[11]) );
  XOR2X2 U46 ( .A(n42), .B(n46), .Y(DIFF[6]) );
  CLKINVX3 U47 ( .A(n136), .Y(n14) );
  INVX2 U48 ( .A(n125), .Y(n136) );
  INVX8 U49 ( .A(n6), .Y(DIFF[14]) );
  NAND4BBX1 U50 ( .AN(n99), .BN(n86), .C(n88), .D(n94), .Y(n95) );
  BUFX4 U51 ( .A(A[13]), .Y(n16) );
  NAND2X4 U52 ( .A(n115), .B(n18), .Y(n17) );
  AOI21X2 U53 ( .A0(n117), .A1(n92), .B0(n119), .Y(n118) );
  NAND2BX4 U54 ( .AN(A[12]), .B(n22), .Y(n116) );
  AOI21X4 U55 ( .A0(A[12]), .A1(n105), .B0(n106), .Y(n102) );
  INVX8 U56 ( .A(n107), .Y(n106) );
  XOR2X4 U57 ( .A(n78), .B(n20), .Y(n19) );
  XOR2X4 U58 ( .A(B[16]), .B(A[16]), .Y(n20) );
  AND3X4 U59 ( .A(n116), .B(n93), .C(n3), .Y(n28) );
  OAI2BB1X4 U60 ( .A0N(n104), .A1N(B[14]), .B0(n1), .Y(n103) );
  NAND2BX4 U61 ( .AN(B[14]), .B(n23), .Y(n101) );
  XOR2X2 U62 ( .A(n39), .B(n40), .Y(DIFF[7]) );
  NAND2XL U63 ( .A(n3), .B(n18), .Y(n26) );
  CLKINVX8 U64 ( .A(B[12]), .Y(n105) );
  INVX4 U65 ( .A(n133), .Y(n37) );
  NAND2X4 U66 ( .A(n33), .B(n38), .Y(n126) );
  OR2X4 U67 ( .A(n103), .B(n102), .Y(n25) );
  AOI21X4 U68 ( .A0(n97), .A1(n21), .B0(n98), .Y(n96) );
  OAI21X2 U69 ( .A0(n85), .A1(n86), .B0(n87), .Y(n83) );
  NAND4BX4 U70 ( .AN(n132), .B(n133), .C(n125), .D(n127), .Y(n86) );
  INVX8 U71 ( .A(n105), .Y(n22) );
  NAND3BX4 U72 ( .AN(n95), .B(n96), .C(n10), .Y(n81) );
  INVX4 U73 ( .A(A[14]), .Y(n104) );
  NAND2X2 U74 ( .A(n121), .B(n87), .Y(n122) );
  OAI2BB1X4 U75 ( .A0N(n123), .A1N(n124), .B0(n14), .Y(n87) );
  NAND3X4 U76 ( .A(n28), .B(n83), .C(n84), .Y(n82) );
  NAND4BX4 U77 ( .AN(n79), .B(n80), .C(n81), .D(n82), .Y(n78) );
  OAI21X4 U78 ( .A0(n143), .A1(n37), .B0(n38), .Y(n29) );
  OAI21X2 U79 ( .A0(n137), .A1(n138), .B0(n139), .Y(n134) );
  NAND2X4 U80 ( .A(n121), .B(n87), .Y(n117) );
  NAND2BX4 U81 ( .AN(A[14]), .B(B[14]), .Y(n93) );
  OAI2BB1X4 U82 ( .A0N(n101), .A1N(n25), .B0(n100), .Y(n80) );
  INVX4 U83 ( .A(n111), .Y(n79) );
  NAND2BX4 U84 ( .AN(A[15]), .B(n21), .Y(n100) );
  INVX8 U85 ( .A(n19), .Y(DIFF[16]) );
  NAND2BX4 U86 ( .AN(B[5]), .B(A[5]), .Y(n51) );
  NAND2BX4 U87 ( .AN(A[9]), .B(B[9]), .Y(n127) );
  NAND2BX2 U88 ( .AN(B[12]), .B(A[12]), .Y(n120) );
  NAND2BX4 U89 ( .AN(A[8]), .B(B[8]), .Y(n133) );
  NAND2BX4 U90 ( .AN(B[13]), .B(n16), .Y(n107) );
  INVX4 U91 ( .A(n29), .Y(n142) );
  NAND2BX2 U92 ( .AN(B[7]), .B(A[7]), .Y(n45) );
  NAND2BX4 U93 ( .AN(A[1]), .B(B[1]), .Y(n75) );
  OAI2BB1X4 U94 ( .A0N(n88), .A1N(n57), .B0(n91), .Y(n34) );
  NAND3X1 U95 ( .A(n126), .B(n127), .C(n128), .Y(n124) );
  INVX4 U96 ( .A(n34), .Y(n143) );
  NAND3X1 U97 ( .A(n146), .B(n147), .C(n41), .Y(n145) );
  NOR2X2 U98 ( .A(n129), .B(n130), .Y(n123) );
  NAND2BX4 U99 ( .AN(n86), .B(n34), .Y(n121) );
  NAND2X4 U100 ( .A(n44), .B(n144), .Y(n91) );
  NAND3X2 U101 ( .A(n145), .B(n48), .C(n45), .Y(n144) );
  NAND4BX2 U102 ( .AN(n50), .B(n58), .C(n41), .D(n44), .Y(n152) );
  NAND2BX4 U103 ( .AN(n89), .B(n99), .Y(n57) );
  INVXL U104 ( .A(n48), .Y(n43) );
  XNOR2X1 U105 ( .A(n57), .B(n27), .Y(DIFF[4]) );
  NAND2XL U106 ( .A(n56), .B(n58), .Y(n27) );
  NAND2XL U107 ( .A(n64), .B(n65), .Y(n59) );
  NOR2XL U108 ( .A(n74), .B(n70), .Y(n73) );
  INVXL U109 ( .A(n71), .Y(n74) );
  NAND2BX4 U110 ( .AN(B[11]), .B(A[11]), .Y(n131) );
  NAND2BX2 U111 ( .AN(B[15]), .B(A[15]), .Y(n111) );
  NAND2BX4 U112 ( .AN(B[4]), .B(A[4]), .Y(n56) );
  NAND2BX4 U113 ( .AN(B[2]), .B(A[2]), .Y(n68) );
  NAND2BX4 U114 ( .AN(B[0]), .B(A[0]), .Y(n76) );
  NAND2BXL U115 ( .AN(A[0]), .B(B[0]), .Y(n77) );
  AOI21XL U116 ( .A0(n88), .A1(n89), .B0(n90), .Y(n85) );
  INVX1 U117 ( .A(n91), .Y(n90) );
  XOR2X1 U118 ( .A(n29), .B(n30), .Y(DIFF[9]) );
  INVXL U119 ( .A(n33), .Y(n31) );
  NOR2BX1 U120 ( .AN(n131), .B(n136), .Y(n135) );
  NAND2X1 U121 ( .A(n51), .B(n56), .Y(n147) );
  NOR2X1 U122 ( .A(n43), .B(n47), .Y(n46) );
  INVXL U123 ( .A(n41), .Y(n47) );
  INVXL U124 ( .A(n38), .Y(n36) );
  NAND2X2 U125 ( .A(n148), .B(n65), .Y(n89) );
  NAND3X1 U126 ( .A(n61), .B(n149), .C(n64), .Y(n148) );
  NAND3X1 U127 ( .A(n150), .B(n71), .C(n68), .Y(n149) );
  NAND2X1 U128 ( .A(n151), .B(n75), .Y(n150) );
  XOR2X1 U129 ( .A(n52), .B(n53), .Y(DIFF[5]) );
  NOR2XL U130 ( .A(n54), .B(n50), .Y(n53) );
  INVX1 U131 ( .A(n51), .Y(n54) );
  NAND2XL U132 ( .A(n44), .B(n45), .Y(n39) );
  AOI21XL U133 ( .A0(n41), .A1(n42), .B0(n43), .Y(n40) );
  INVX1 U134 ( .A(n52), .Y(n49) );
  NAND2X1 U135 ( .A(n55), .B(n56), .Y(n52) );
  NAND2XL U136 ( .A(n57), .B(n58), .Y(n55) );
  XOR2X1 U137 ( .A(n62), .B(n66), .Y(DIFF[2]) );
  NOR2X1 U138 ( .A(n63), .B(n67), .Y(n66) );
  INVXL U139 ( .A(n61), .Y(n67) );
  XOR2X1 U140 ( .A(n72), .B(n73), .Y(DIFF[1]) );
  XOR2X1 U141 ( .A(n59), .B(n60), .Y(DIFF[3]) );
  AOI21XL U142 ( .A0(n61), .A1(n62), .B0(n63), .Y(n60) );
  OAI21XL U143 ( .A0(n69), .A1(n70), .B0(n71), .Y(n62) );
  INVX1 U144 ( .A(n72), .Y(n69) );
  INVX1 U145 ( .A(n75), .Y(n70) );
  INVX1 U146 ( .A(n68), .Y(n63) );
  NAND2BX2 U147 ( .AN(A[3]), .B(B[3]), .Y(n64) );
  NAND4X1 U148 ( .A(n77), .B(n75), .C(n61), .D(n64), .Y(n99) );
  NAND2BX1 U149 ( .AN(B[6]), .B(A[6]), .Y(n48) );
  NAND2BX2 U150 ( .AN(B[1]), .B(A[1]), .Y(n71) );
  NAND2BX1 U151 ( .AN(B[3]), .B(A[3]), .Y(n65) );
  INVX1 U152 ( .A(n76), .Y(n151) );
  NAND2X1 U153 ( .A(n77), .B(n76), .Y(DIFF[0]) );
  NAND2BX1 U154 ( .AN(n77), .B(n76), .Y(n72) );
  XOR2X4 U155 ( .A(n108), .B(n109), .Y(DIFF[15]) );
  NOR2X4 U156 ( .A(n110), .B(n79), .Y(n109) );
  OAI21X4 U157 ( .A0(n8), .A1(n112), .B0(n5), .Y(n108) );
  NOR2X4 U158 ( .A(n112), .B(n114), .Y(n113) );
  CLKINVX3 U159 ( .A(n120), .Y(n119) );
  NAND2BX4 U160 ( .AN(A[13]), .B(B[13]), .Y(n94) );
  NAND2BX4 U161 ( .AN(A[12]), .B(n22), .Y(n92) );
  NAND2BX4 U162 ( .AN(A[11]), .B(B[11]), .Y(n125) );
  NAND2BX4 U163 ( .AN(B[9]), .B(A[9]), .Y(n33) );
  NAND2BX4 U164 ( .AN(B[8]), .B(A[8]), .Y(n38) );
  NAND2BX4 U165 ( .AN(A[2]), .B(B[2]), .Y(n61) );
  CLKINVX3 U166 ( .A(n152), .Y(n88) );
  NAND2BX4 U167 ( .AN(A[7]), .B(B[7]), .Y(n44) );
  NAND2BX4 U168 ( .AN(A[6]), .B(B[6]), .Y(n41) );
  NAND2BX4 U169 ( .AN(A[4]), .B(B[4]), .Y(n58) );
endmodule


module butterfly_DW01_add_77 ( A, B, SUM );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127;

  AND2X2 U2 ( .A(n67), .B(n75), .Y(n4) );
  INVX4 U3 ( .A(n64), .Y(n63) );
  NAND2X4 U4 ( .A(B[15]), .B(A[15]), .Y(n64) );
  BUFX4 U5 ( .A(n67), .Y(n1) );
  NAND2X2 U6 ( .A(B[14]), .B(A[14]), .Y(n67) );
  OAI2BB1X1 U7 ( .A0N(n19), .A1N(n97), .B0(n77), .Y(n106) );
  NOR2X2 U8 ( .A(A[4]), .B(B[4]), .Y(n14) );
  NAND2X4 U9 ( .A(n121), .B(n21), .Y(n15) );
  NOR2BX4 U10 ( .AN(n21), .B(n22), .Y(n20) );
  NAND2X4 U11 ( .A(B[8]), .B(A[8]), .Y(n21) );
  OAI21X2 U12 ( .A0(A[10]), .A1(B[10]), .B0(n109), .Y(n92) );
  NAND3X4 U13 ( .A(n92), .B(n91), .C(n5), .Y(n108) );
  NAND2X4 U14 ( .A(n82), .B(n1), .Y(n6) );
  INVX1 U15 ( .A(A[15]), .Y(n3) );
  NAND3X1 U16 ( .A(n91), .B(n5), .C(n92), .Y(n90) );
  AOI21X2 U17 ( .A0(n61), .A1(n62), .B0(n63), .Y(n60) );
  OAI211X1 U18 ( .A0(n86), .A1(n65), .B0(n66), .C0(n67), .Y(n62) );
  INVX2 U19 ( .A(n23), .Y(n22) );
  NOR2BX2 U20 ( .AN(n39), .B(n14), .Y(n40) );
  INVX4 U21 ( .A(n68), .Y(n86) );
  AND2X4 U22 ( .A(B[11]), .B(A[11]), .Y(n2) );
  XOR2X4 U23 ( .A(n116), .B(n118), .Y(SUM[10]) );
  XOR2X4 U24 ( .A(n15), .B(n16), .Y(SUM[9]) );
  NOR2BX2 U25 ( .AN(n17), .B(n18), .Y(n16) );
  AOI211X2 U26 ( .A0(n35), .A1(n39), .B0(n30), .C0(n13), .Y(n122) );
  NAND2X4 U27 ( .A(B[4]), .B(A[4]), .Y(n39) );
  XOR2X4 U28 ( .A(n114), .B(n115), .Y(SUM[11]) );
  NOR2BX4 U29 ( .AN(n91), .B(n119), .Y(n118) );
  INVX4 U30 ( .A(n91), .Y(n117) );
  OR2X4 U31 ( .A(A[8]), .B(B[8]), .Y(n23) );
  INVX1 U32 ( .A(n113), .Y(n119) );
  NAND2X2 U33 ( .A(B[10]), .B(A[10]), .Y(n91) );
  NAND2X4 U34 ( .A(n104), .B(n65), .Y(n102) );
  NAND2X2 U35 ( .A(n89), .B(n5), .Y(n114) );
  CLKINVX8 U36 ( .A(n2), .Y(n5) );
  NAND3BX2 U37 ( .AN(n72), .B(n73), .C(n74), .Y(n59) );
  NAND2BX4 U38 ( .AN(B[15]), .B(n3), .Y(n69) );
  NAND3BX2 U39 ( .AN(n11), .B(n89), .C(n90), .Y(n88) );
  NOR2XL U40 ( .A(A[15]), .B(B[15]), .Y(n72) );
  XOR2X4 U41 ( .A(n8), .B(n4), .Y(SUM[14]) );
  CLKINVX8 U42 ( .A(n70), .Y(n97) );
  NAND2X4 U43 ( .A(n66), .B(n65), .Y(n94) );
  NOR2X4 U44 ( .A(B[12]), .B(A[12]), .Y(n11) );
  NOR2X2 U45 ( .A(A[12]), .B(B[12]), .Y(n95) );
  NAND3BX2 U46 ( .AN(n11), .B(n19), .C(n97), .Y(n103) );
  OAI21X2 U47 ( .A0(A[11]), .A1(B[11]), .B0(n113), .Y(n110) );
  NOR2BX2 U48 ( .AN(n69), .B(n85), .Y(n61) );
  OAI21X4 U49 ( .A0(A[12]), .A1(B[12]), .B0(n89), .Y(n105) );
  INVX8 U50 ( .A(n75), .Y(n85) );
  NAND2X4 U51 ( .A(n59), .B(n60), .Y(n57) );
  NAND2X4 U52 ( .A(B[12]), .B(A[12]), .Y(n65) );
  XOR2X2 U53 ( .A(n79), .B(n40), .Y(SUM[4]) );
  NAND2X2 U54 ( .A(n19), .B(n97), .Y(n96) );
  XOR2X4 U55 ( .A(n106), .B(n107), .Y(SUM[12]) );
  NAND2X4 U56 ( .A(n87), .B(n88), .Y(n83) );
  NOR2X4 U57 ( .A(n93), .B(n94), .Y(n87) );
  NOR2X4 U58 ( .A(n95), .B(n96), .Y(n93) );
  OR2X4 U59 ( .A(A[6]), .B(B[6]), .Y(n124) );
  NOR3X2 U60 ( .A(n85), .B(n11), .C(n86), .Y(n74) );
  NAND2X4 U61 ( .A(n83), .B(n84), .Y(n82) );
  NAND2X2 U62 ( .A(B[9]), .B(A[9]), .Y(n17) );
  INVX2 U63 ( .A(n99), .Y(n100) );
  NAND2X4 U64 ( .A(B[5]), .B(A[5]), .Y(n35) );
  OAI21X4 U65 ( .A0(n34), .A1(n13), .B0(n35), .Y(n32) );
  NOR2BX4 U66 ( .AN(n35), .B(n13), .Y(n37) );
  XOR2X2 U67 ( .A(B[16]), .B(A[16]), .Y(n58) );
  NAND2X4 U68 ( .A(B[13]), .B(A[13]), .Y(n66) );
  NAND2X2 U69 ( .A(n66), .B(n68), .Y(n101) );
  OR2X4 U70 ( .A(A[13]), .B(B[13]), .Y(n68) );
  NAND2BX4 U71 ( .AN(n105), .B(n108), .Y(n104) );
  NOR2BX2 U72 ( .AN(n65), .B(n95), .Y(n107) );
  NOR2BX4 U73 ( .AN(n26), .B(n27), .Y(n25) );
  NAND2X2 U74 ( .A(B[7]), .B(A[7]), .Y(n26) );
  NOR2X4 U75 ( .A(n85), .B(n86), .Y(n84) );
  OR2X4 U76 ( .A(A[10]), .B(B[10]), .Y(n113) );
  AOI21X2 U77 ( .A0(n17), .A1(n21), .B0(n18), .Y(n109) );
  XOR2X2 U78 ( .A(n32), .B(n33), .Y(SUM[6]) );
  NOR2BX2 U79 ( .AN(n31), .B(n30), .Y(n33) );
  OAI21X2 U80 ( .A0(n29), .A1(n30), .B0(n31), .Y(n24) );
  INVX2 U81 ( .A(n32), .Y(n29) );
  XOR2X4 U82 ( .A(n24), .B(n25), .Y(SUM[7]) );
  NAND4BBX2 U83 ( .AN(n13), .BN(n14), .C(n124), .D(n28), .Y(n71) );
  OAI21X4 U84 ( .A0(n122), .A1(n123), .B0(n28), .Y(n81) );
  AOI21X2 U85 ( .A0(n113), .A1(n116), .B0(n117), .Y(n115) );
  NOR2X4 U86 ( .A(A[5]), .B(B[5]), .Y(n13) );
  NAND2X2 U87 ( .A(n19), .B(n23), .Y(n121) );
  XOR2X4 U88 ( .A(n58), .B(n57), .Y(SUM[16]) );
  NAND2X1 U89 ( .A(B[1]), .B(A[1]), .Y(n53) );
  XOR2X4 U90 ( .A(n100), .B(n101), .Y(SUM[13]) );
  INVX4 U91 ( .A(n124), .Y(n30) );
  INVX4 U92 ( .A(n15), .Y(n120) );
  OR2X4 U93 ( .A(A[1]), .B(B[1]), .Y(n51) );
  OAI21X4 U94 ( .A0(n120), .A1(n18), .B0(n17), .Y(n116) );
  XOR2X2 U95 ( .A(n19), .B(n20), .Y(SUM[8]) );
  OAI2BB1X4 U96 ( .A0N(n9), .A1N(n10), .B0(n43), .Y(n79) );
  OR2X4 U97 ( .A(A[7]), .B(B[7]), .Y(n28) );
  NAND2XL U98 ( .A(n112), .B(n23), .Y(n111) );
  INVX4 U99 ( .A(n79), .Y(n38) );
  XOR2X4 U100 ( .A(n6), .B(n7), .Y(SUM[15]) );
  AND2X4 U101 ( .A(n64), .B(n69), .Y(n7) );
  NAND2X2 U102 ( .A(n89), .B(n108), .Y(n77) );
  NAND2X4 U103 ( .A(n98), .B(n66), .Y(n8) );
  OR2X2 U104 ( .A(n126), .B(n127), .Y(n9) );
  AND2X2 U105 ( .A(n50), .B(n125), .Y(n10) );
  NAND2X2 U106 ( .A(n26), .B(n31), .Y(n123) );
  OAI21X4 U107 ( .A0(n14), .A1(n38), .B0(n39), .Y(n36) );
  CLKINVX3 U108 ( .A(n47), .Y(n126) );
  INVX2 U109 ( .A(n36), .Y(n34) );
  INVX4 U110 ( .A(n112), .Y(n18) );
  OAI21XL U111 ( .A0(n45), .A1(n46), .B0(n47), .Y(n41) );
  XOR2X1 U112 ( .A(n48), .B(n49), .Y(SUM[2]) );
  OAI2BB1X2 U113 ( .A0N(n51), .A1N(n52), .B0(n53), .Y(n48) );
  XOR2X1 U114 ( .A(n52), .B(n54), .Y(SUM[1]) );
  OR2X4 U115 ( .A(B[14]), .B(A[14]), .Y(n75) );
  OR2XL U116 ( .A(A[2]), .B(B[2]), .Y(n50) );
  OR2XL U117 ( .A(A[3]), .B(B[3]), .Y(n125) );
  NAND2X1 U118 ( .A(B[0]), .B(A[0]), .Y(n56) );
  NOR2BX1 U119 ( .AN(n56), .B(n12), .Y(SUM[0]) );
  NOR2XL U120 ( .A(A[0]), .B(B[0]), .Y(n12) );
  AOI21X1 U121 ( .A0(n78), .A1(n79), .B0(n80), .Y(n76) );
  INVX1 U122 ( .A(n71), .Y(n78) );
  INVX1 U123 ( .A(n81), .Y(n80) );
  OAI21XL U124 ( .A0(n76), .A1(n70), .B0(n77), .Y(n73) );
  OAI21XL U125 ( .A0(n55), .A1(n56), .B0(n53), .Y(n127) );
  XOR2X1 U126 ( .A(n36), .B(n37), .Y(SUM[5]) );
  INVX1 U127 ( .A(n28), .Y(n27) );
  INVX1 U128 ( .A(n51), .Y(n55) );
  INVX1 U129 ( .A(n50), .Y(n46) );
  XOR2X2 U130 ( .A(n41), .B(n42), .Y(SUM[3]) );
  NOR2BX1 U131 ( .AN(n43), .B(n44), .Y(n42) );
  INVX1 U132 ( .A(n48), .Y(n45) );
  NOR2BX1 U133 ( .AN(n47), .B(n46), .Y(n49) );
  NOR2BXL U134 ( .AN(n53), .B(n55), .Y(n54) );
  INVX1 U135 ( .A(n125), .Y(n44) );
  INVX1 U136 ( .A(n56), .Y(n52) );
  NAND2XL U137 ( .A(B[6]), .B(A[6]), .Y(n31) );
  NAND2X2 U138 ( .A(B[2]), .B(A[2]), .Y(n47) );
  NAND2XL U139 ( .A(B[3]), .B(A[3]), .Y(n43) );
  NAND2X2 U140 ( .A(n68), .B(n99), .Y(n98) );
  NAND2BX4 U141 ( .AN(n102), .B(n103), .Y(n99) );
  OR2X4 U142 ( .A(n111), .B(n110), .Y(n70) );
  OR2X4 U143 ( .A(A[11]), .B(B[11]), .Y(n89) );
  OR2X4 U144 ( .A(A[9]), .B(B[9]), .Y(n112) );
  OAI21X4 U145 ( .A0(n38), .A1(n71), .B0(n81), .Y(n19) );
endmodule


module butterfly_DW01_add_73 ( A, B, SUM );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  wire   n1, n2, n3, n4, n5, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135;

  INVX4 U2 ( .A(n11), .Y(n1) );
  NOR2BX2 U3 ( .AN(n99), .B(n103), .Y(n102) );
  BUFX1 U4 ( .A(n99), .Y(n9) );
  NOR2X2 U5 ( .A(B[15]), .B(A[15]), .Y(n2) );
  NAND2X4 U6 ( .A(n126), .B(n41), .Y(n35) );
  NAND2X4 U7 ( .A(n39), .B(n118), .Y(n126) );
  BUFX8 U8 ( .A(B[12]), .Y(n19) );
  CLKINVX4 U9 ( .A(n107), .Y(n25) );
  INVX4 U10 ( .A(n79), .Y(n112) );
  NAND2X4 U11 ( .A(n16), .B(n25), .Y(n26) );
  INVX2 U12 ( .A(n24), .Y(n16) );
  NAND2X1 U13 ( .A(n107), .B(n24), .Y(n27) );
  XOR2X4 U14 ( .A(n100), .B(n4), .Y(n3) );
  OR2X4 U15 ( .A(n5), .B(n1), .Y(n4) );
  XOR2X4 U16 ( .A(n110), .B(n111), .Y(SUM[12]) );
  AND2X2 U17 ( .A(A[15]), .B(B[15]), .Y(n5) );
  INVX8 U18 ( .A(n3), .Y(SUM[15]) );
  OAI21X2 U19 ( .A0(n53), .A1(n33), .B0(n54), .Y(n51) );
  XOR2X2 U20 ( .A(n51), .B(n52), .Y(SUM[6]) );
  AND2X2 U21 ( .A(n79), .B(n78), .Y(n7) );
  XOR2X4 U22 ( .A(n43), .B(n44), .Y(SUM[7]) );
  NAND2BX2 U23 ( .AN(n119), .B(n120), .Y(n23) );
  BUFX4 U24 ( .A(n83), .Y(n8) );
  NAND2XL U25 ( .A(B[11]), .B(A[11]), .Y(n83) );
  NOR2BX2 U26 ( .AN(n115), .B(n124), .Y(n123) );
  INVX2 U27 ( .A(n120), .Y(n21) );
  NAND2X2 U28 ( .A(n28), .B(n91), .Y(n98) );
  NOR2X4 U29 ( .A(n117), .B(n42), .Y(n116) );
  INVX4 U30 ( .A(n118), .Y(n42) );
  INVX3 U31 ( .A(n39), .Y(n117) );
  AOI211X2 U32 ( .A0(n54), .A1(n57), .B0(n49), .C0(n33), .Y(n127) );
  INVXL U33 ( .A(n88), .Y(n87) );
  AND2X2 U34 ( .A(n84), .B(n8), .Y(n82) );
  NAND2X4 U35 ( .A(n19), .B(A[12]), .Y(n109) );
  OR2X4 U36 ( .A(A[2]), .B(B[2]), .Y(n69) );
  NAND2BX4 U37 ( .AN(n10), .B(n114), .Y(n84) );
  NAND2X4 U38 ( .A(n95), .B(n94), .Y(n10) );
  INVX4 U39 ( .A(n2), .Y(n11) );
  NOR2X4 U40 ( .A(A[5]), .B(B[5]), .Y(n33) );
  INVX8 U41 ( .A(n91), .Y(n104) );
  OAI211X2 U42 ( .A0(n38), .A1(n41), .B0(n37), .C0(n115), .Y(n114) );
  INVX8 U43 ( .A(n93), .Y(n38) );
  NAND2X4 U44 ( .A(B[9]), .B(A[9]), .Y(n37) );
  NAND2X4 U45 ( .A(n7), .B(n30), .Y(n77) );
  INVX4 U46 ( .A(B[16]), .Y(n12) );
  NAND2X2 U47 ( .A(A[16]), .B(B[16]), .Y(n14) );
  NAND2X4 U48 ( .A(n13), .B(n12), .Y(n15) );
  NAND2X4 U49 ( .A(n14), .B(n15), .Y(n18) );
  INVX4 U50 ( .A(A[16]), .Y(n13) );
  NAND2X2 U51 ( .A(A[14]), .B(B[14]), .Y(n99) );
  INVX2 U52 ( .A(n90), .Y(n103) );
  OAI21X4 U53 ( .A0(n130), .A1(n89), .B0(n88), .Y(n39) );
  INVX8 U54 ( .A(n106), .Y(n24) );
  NAND2X4 U55 ( .A(B[6]), .B(A[6]), .Y(n50) );
  CLKINVX2 U56 ( .A(n89), .Y(n85) );
  NAND4BBX2 U57 ( .AN(n33), .BN(n34), .C(n129), .D(n47), .Y(n89) );
  XOR2X2 U58 ( .A(n35), .B(n36), .Y(SUM[9]) );
  XOR2X4 U59 ( .A(n32), .B(n18), .Y(n17) );
  AOI22X2 U60 ( .A0(n19), .A1(A[12]), .B0(B[13]), .B1(A[13]), .Y(n97) );
  OAI21X2 U61 ( .A0(n80), .A1(n81), .B0(n82), .Y(n78) );
  NAND2X2 U62 ( .A(B[13]), .B(A[13]), .Y(n105) );
  OAI21X4 U63 ( .A0(n24), .A1(n104), .B0(n105), .Y(n20) );
  OAI21X2 U64 ( .A0(n24), .A1(n104), .B0(n105), .Y(n101) );
  OAI21X2 U65 ( .A0(n34), .A1(n130), .B0(n57), .Y(n55) );
  NOR2X4 U66 ( .A(A[4]), .B(B[4]), .Y(n34) );
  OAI21X4 U67 ( .A0(n97), .A1(n98), .B0(n99), .Y(n96) );
  NAND2X4 U68 ( .A(n110), .B(n79), .Y(n108) );
  NAND3X4 U69 ( .A(n84), .B(n8), .C(n113), .Y(n110) );
  OR2X4 U70 ( .A(A[14]), .B(B[14]), .Y(n28) );
  XOR2X4 U71 ( .A(n121), .B(n123), .Y(SUM[10]) );
  NAND4X2 U72 ( .A(n116), .B(n93), .C(n94), .D(n95), .Y(n113) );
  NAND2X2 U73 ( .A(n119), .B(n21), .Y(n22) );
  NAND2X4 U74 ( .A(n22), .B(n23), .Y(SUM[11]) );
  AOI21X2 U75 ( .A0(n94), .A1(n121), .B0(n122), .Y(n120) );
  NAND2X4 U76 ( .A(n26), .B(n27), .Y(SUM[13]) );
  NAND2X4 U77 ( .A(n108), .B(n109), .Y(n106) );
  NAND2X4 U78 ( .A(B[8]), .B(A[8]), .Y(n41) );
  NOR2BX2 U79 ( .AN(n37), .B(n38), .Y(n36) );
  INVX8 U80 ( .A(n17), .Y(SUM[16]) );
  NAND2X4 U81 ( .A(n76), .B(n77), .Y(n32) );
  OAI21X4 U82 ( .A0(n132), .A1(n133), .B0(n62), .Y(n86) );
  OAI21X4 U83 ( .A0(n125), .A1(n38), .B0(n37), .Y(n121) );
  NAND2X4 U84 ( .A(B[4]), .B(A[4]), .Y(n57) );
  NAND2X4 U85 ( .A(B[2]), .B(A[2]), .Y(n66) );
  NAND2X1 U86 ( .A(B[7]), .B(A[7]), .Y(n45) );
  INVX4 U87 ( .A(n35), .Y(n125) );
  NAND2X2 U88 ( .A(B[5]), .B(A[5]), .Y(n54) );
  NAND2X1 U89 ( .A(B[1]), .B(A[1]), .Y(n72) );
  AND3X4 U90 ( .A(n92), .B(n91), .C(n90), .Y(n30) );
  INVXL U91 ( .A(n131), .Y(n63) );
  OAI2BB1X1 U92 ( .A0N(n70), .A1N(n71), .B0(n72), .Y(n67) );
  NAND2XL U93 ( .A(B[3]), .B(A[3]), .Y(n62) );
  NOR2BX4 U94 ( .AN(n105), .B(n104), .Y(n107) );
  OAI21X2 U95 ( .A0(n127), .A1(n128), .B0(n47), .Y(n88) );
  NAND2X2 U96 ( .A(n45), .B(n50), .Y(n128) );
  INVX4 U97 ( .A(n129), .Y(n49) );
  INVX2 U98 ( .A(n55), .Y(n53) );
  NOR2X2 U99 ( .A(n134), .B(n135), .Y(n132) );
  OAI21X2 U100 ( .A0(n74), .A1(n75), .B0(n72), .Y(n135) );
  OAI21X1 U101 ( .A0(n64), .A1(n65), .B0(n66), .Y(n60) );
  NAND2X2 U102 ( .A(B[10]), .B(A[10]), .Y(n115) );
  OR2X4 U103 ( .A(A[3]), .B(B[3]), .Y(n131) );
  OR2X4 U104 ( .A(A[1]), .B(B[1]), .Y(n70) );
  NAND2X4 U105 ( .A(B[0]), .B(A[0]), .Y(n75) );
  NOR2BX1 U106 ( .AN(n75), .B(n31), .Y(SUM[0]) );
  NOR2XL U107 ( .A(A[0]), .B(B[0]), .Y(n31) );
  INVX1 U108 ( .A(n130), .Y(n58) );
  INVX1 U109 ( .A(n86), .Y(n130) );
  INVX1 U110 ( .A(n51), .Y(n48) );
  INVX1 U111 ( .A(n67), .Y(n64) );
  NAND4BXL U112 ( .AN(n42), .B(n95), .C(n94), .D(n93), .Y(n81) );
  AOI21X1 U113 ( .A0(n85), .A1(n86), .B0(n87), .Y(n80) );
  INVXL U114 ( .A(n94), .Y(n124) );
  NAND2XL U115 ( .A(n8), .B(n95), .Y(n119) );
  INVX1 U116 ( .A(n115), .Y(n122) );
  XOR2X1 U117 ( .A(n39), .B(n40), .Y(SUM[8]) );
  NOR2BXL U118 ( .AN(n41), .B(n42), .Y(n40) );
  NAND2X1 U119 ( .A(n69), .B(n131), .Y(n133) );
  INVX1 U120 ( .A(n70), .Y(n74) );
  INVX1 U121 ( .A(n66), .Y(n134) );
  NOR2BXL U122 ( .AN(n50), .B(n49), .Y(n52) );
  XOR2X1 U123 ( .A(n55), .B(n56), .Y(SUM[5]) );
  NOR2BX1 U124 ( .AN(n54), .B(n33), .Y(n56) );
  NOR2BX1 U125 ( .AN(n45), .B(n46), .Y(n44) );
  OAI21XL U126 ( .A0(n48), .A1(n49), .B0(n50), .Y(n43) );
  INVXL U127 ( .A(n47), .Y(n46) );
  XOR2X1 U128 ( .A(n60), .B(n61), .Y(SUM[3]) );
  NOR2BX1 U129 ( .AN(n62), .B(n63), .Y(n61) );
  XOR2X1 U130 ( .A(n58), .B(n59), .Y(SUM[4]) );
  NOR2BX1 U131 ( .AN(n57), .B(n34), .Y(n59) );
  INVX1 U132 ( .A(n69), .Y(n65) );
  XOR2X1 U133 ( .A(n67), .B(n68), .Y(SUM[2]) );
  NOR2BXL U134 ( .AN(n66), .B(n65), .Y(n68) );
  XOR2X1 U135 ( .A(n71), .B(n73), .Y(SUM[1]) );
  NOR2BXL U136 ( .AN(n72), .B(n74), .Y(n73) );
  INVX1 U137 ( .A(n75), .Y(n71) );
  XOR2X4 U138 ( .A(n101), .B(n102), .Y(SUM[14]) );
  AOI21X4 U139 ( .A0(n96), .A1(n11), .B0(n5), .Y(n76) );
  OR2X4 U140 ( .A(B[15]), .B(A[15]), .Y(n92) );
  OAI2BB1X4 U141 ( .A0N(n90), .A1N(n20), .B0(n9), .Y(n100) );
  OR2X4 U142 ( .A(A[14]), .B(B[14]), .Y(n90) );
  OR2X4 U143 ( .A(A[13]), .B(B[13]), .Y(n91) );
  NOR2BX4 U144 ( .AN(n109), .B(n112), .Y(n111) );
  OR2X4 U145 ( .A(A[12]), .B(B[12]), .Y(n79) );
  OR2X4 U146 ( .A(B[11]), .B(A[11]), .Y(n95) );
  OR2X4 U147 ( .A(B[10]), .B(A[10]), .Y(n94) );
  OR2X4 U148 ( .A(A[9]), .B(B[9]), .Y(n93) );
  OR2X4 U149 ( .A(A[8]), .B(B[8]), .Y(n118) );
  OR2X4 U150 ( .A(A[7]), .B(B[7]), .Y(n47) );
  OR2X4 U151 ( .A(A[6]), .B(B[6]), .Y(n129) );
endmodule


module butterfly_DW01_sub_64 ( A, B, DIFF );
  input [16:0] A;
  input [16:0] B;
  output [16:0] DIFF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142;

  INVX4 U3 ( .A(n109), .Y(n1) );
  CLKINVX8 U4 ( .A(n74), .Y(n109) );
  INVX1 U5 ( .A(B[13]), .Y(n9) );
  NAND2X4 U6 ( .A(n4), .B(B[15]), .Y(n77) );
  INVX20 U7 ( .A(A[15]), .Y(n4) );
  AOI2BB1X4 U8 ( .A0N(n3), .A1N(n2), .B0(n79), .Y(n65) );
  CLKINVX20 U9 ( .A(n78), .Y(n2) );
  OR2X4 U10 ( .A(n87), .B(n88), .Y(n3) );
  OAI2BB1X2 U11 ( .A0N(n11), .A1N(n10), .B0(n76), .Y(n101) );
  OAI21X2 U12 ( .A0(n90), .A1(n91), .B0(n92), .Y(n87) );
  NAND4BX2 U13 ( .AN(n25), .B(n95), .C(n96), .D(n97), .Y(n94) );
  NAND2X2 U14 ( .A(n93), .B(n83), .Y(n91) );
  NAND2BX4 U15 ( .AN(n5), .B(n70), .Y(n68) );
  NAND2X4 U16 ( .A(n74), .B(n7), .Y(n5) );
  NOR2X2 U17 ( .A(n80), .B(n110), .Y(n67) );
  INVX8 U18 ( .A(n77), .Y(n80) );
  INVX8 U19 ( .A(n102), .Y(n115) );
  NAND2BX4 U20 ( .AN(A[12]), .B(n18), .Y(n82) );
  CLKINVX2 U21 ( .A(n113), .Y(n7) );
  INVX3 U22 ( .A(n10), .Y(n71) );
  NAND3X2 U23 ( .A(n48), .B(n51), .C(n136), .Y(n90) );
  INVX1 U24 ( .A(A[14]), .Y(n8) );
  XOR2X2 U25 ( .A(n46), .B(n47), .Y(DIFF[3]) );
  NAND2X1 U26 ( .A(n43), .B(n45), .Y(n13) );
  INVX2 U27 ( .A(n96), .Y(n130) );
  NAND2X2 U28 ( .A(n83), .B(n84), .Y(n78) );
  INVXL U29 ( .A(n58), .Y(n60) );
  NOR2X2 U30 ( .A(n50), .B(n54), .Y(n53) );
  AND2X4 U31 ( .A(n139), .B(n52), .Y(n6) );
  INVX1 U32 ( .A(A[13]), .Y(n11) );
  NAND2BX4 U33 ( .AN(n18), .B(A[12]), .Y(n73) );
  NOR2BX2 U34 ( .AN(n18), .B(A[12]), .Y(n116) );
  BUFX8 U35 ( .A(B[12]), .Y(n18) );
  AND2X4 U36 ( .A(n97), .B(n92), .Y(n17) );
  NAND2BX4 U37 ( .AN(A[5]), .B(B[5]), .Y(n134) );
  NAND2BX4 U38 ( .AN(B[5]), .B(A[5]), .Y(n38) );
  XOR2X2 U39 ( .A(n39), .B(n40), .Y(DIFF[5]) );
  NAND2BX1 U40 ( .AN(A[8]), .B(B[8]), .Y(n142) );
  NAND2BX2 U41 ( .AN(A[3]), .B(B[3]), .Y(n51) );
  NAND2BX4 U42 ( .AN(B[3]), .B(A[3]), .Y(n52) );
  NAND2X2 U43 ( .A(n38), .B(n43), .Y(n135) );
  NAND2X2 U44 ( .A(n42), .B(n43), .Y(n39) );
  NAND2BX1 U45 ( .AN(B[4]), .B(A[4]), .Y(n43) );
  INVX2 U46 ( .A(n73), .Y(n72) );
  INVX4 U47 ( .A(n75), .Y(n113) );
  INVX4 U48 ( .A(n9), .Y(n10) );
  NAND2BX4 U49 ( .AN(A[7]), .B(B[7]), .Y(n31) );
  NAND2BX4 U50 ( .AN(A[14]), .B(B[14]), .Y(n76) );
  XOR2X4 U51 ( .A(n26), .B(n27), .Y(DIFF[7]) );
  INVX1 U52 ( .A(A[12]), .Y(n118) );
  NAND2BX4 U53 ( .AN(n18), .B(A[12]), .Y(n103) );
  NAND2BX4 U54 ( .AN(B[9]), .B(A[9]), .Y(n124) );
  NAND2BX4 U55 ( .AN(B[7]), .B(A[7]), .Y(n32) );
  NAND3X2 U56 ( .A(n133), .B(n35), .C(n32), .Y(n132) );
  NAND4BX4 U57 ( .AN(n80), .B(n81), .C(n76), .D(n82), .Y(n79) );
  NAND2BX1 U58 ( .AN(A[13]), .B(n10), .Y(n81) );
  AOI21X4 U59 ( .A0(n82), .A1(n102), .B0(n108), .Y(n106) );
  OR2X4 U60 ( .A(B[14]), .B(n8), .Y(n74) );
  AND2X1 U61 ( .A(B[13]), .B(n11), .Y(n114) );
  NAND2BX4 U62 ( .AN(B[13]), .B(A[13]), .Y(n75) );
  NOR2X4 U63 ( .A(n80), .B(n99), .Y(n14) );
  NOR2BX2 U64 ( .AN(A[15]), .B(B[15]), .Y(n99) );
  NAND2X4 U65 ( .A(n103), .B(n75), .Y(n108) );
  NAND3BX2 U66 ( .AN(n20), .B(n121), .C(n122), .Y(n120) );
  NAND2BX4 U67 ( .AN(B[10]), .B(A[10]), .Y(n122) );
  NOR2X4 U68 ( .A(n20), .B(n21), .Y(n12) );
  NAND2BX4 U69 ( .AN(B[11]), .B(A[11]), .Y(n92) );
  NOR2X4 U70 ( .A(n106), .B(n107), .Y(n105) );
  NAND3X4 U71 ( .A(n120), .B(n96), .C(n97), .Y(n89) );
  AOI21X2 U72 ( .A0(n96), .A1(n127), .B0(n128), .Y(n126) );
  NAND2BX4 U73 ( .AN(A[10]), .B(B[10]), .Y(n96) );
  AOI21X2 U74 ( .A0(n82), .A1(n102), .B0(n108), .Y(n100) );
  INVX4 U75 ( .A(n76), .Y(n110) );
  NAND3X4 U76 ( .A(n119), .B(n92), .C(n89), .Y(n102) );
  NAND4BX2 U77 ( .AN(n16), .B(n95), .C(n96), .D(n97), .Y(n119) );
  INVX4 U78 ( .A(n122), .Y(n128) );
  NAND2X4 U79 ( .A(n31), .B(n132), .Y(n86) );
  OAI2BB1X2 U80 ( .A0N(n93), .A1N(n44), .B0(n86), .Y(n22) );
  XOR2X4 U81 ( .A(n19), .B(n12), .Y(DIFF[9]) );
  NAND2BX4 U82 ( .AN(B[6]), .B(A[6]), .Y(n35) );
  NAND2BX4 U83 ( .AN(A[9]), .B(B[9]), .Y(n95) );
  CLKINVX4 U84 ( .A(n95), .Y(n21) );
  XOR2X2 U85 ( .A(n22), .B(n23), .Y(DIFF[8]) );
  NAND2BX4 U86 ( .AN(B[8]), .B(A[8]), .Y(n123) );
  NOR2X2 U87 ( .A(n30), .B(n34), .Y(n33) );
  INVX2 U88 ( .A(n28), .Y(n34) );
  INVX2 U89 ( .A(n138), .Y(n57) );
  XNOR2X2 U90 ( .A(n44), .B(n13), .Y(DIFF[4]) );
  AOI21X4 U91 ( .A0(n28), .A1(n29), .B0(n30), .Y(n27) );
  NAND2X2 U92 ( .A(n31), .B(n32), .Y(n26) );
  OAI21X2 U93 ( .A0(n36), .A1(n37), .B0(n38), .Y(n29) );
  CLKINVX3 U94 ( .A(n137), .Y(n61) );
  AOI21X1 U95 ( .A0(n48), .A1(n49), .B0(n50), .Y(n47) );
  NAND2BX1 U96 ( .AN(A[4]), .B(B[4]), .Y(n45) );
  NAND2X4 U97 ( .A(n44), .B(n45), .Y(n42) );
  NOR2X2 U98 ( .A(n24), .B(n25), .Y(n23) );
  INVX4 U99 ( .A(n35), .Y(n30) );
  NAND3X2 U100 ( .A(n48), .B(n140), .C(n51), .Y(n139) );
  NAND3X2 U101 ( .A(n141), .B(n58), .C(n55), .Y(n140) );
  XOR2X4 U102 ( .A(n98), .B(n14), .Y(DIFF[15]) );
  INVXL U103 ( .A(n55), .Y(n50) );
  INVX4 U104 ( .A(n124), .Y(n20) );
  XOR2X1 U105 ( .A(n59), .B(n15), .Y(DIFF[1]) );
  NOR2XL U106 ( .A(n60), .B(n57), .Y(n15) );
  NAND2XL U107 ( .A(n24), .B(n95), .Y(n121) );
  NAND2XL U108 ( .A(n51), .B(n52), .Y(n46) );
  NAND2XL U109 ( .A(n61), .B(n62), .Y(n59) );
  NAND2XL U110 ( .A(n137), .B(n62), .Y(DIFF[0]) );
  NAND2BXL U111 ( .AN(A[2]), .B(B[2]), .Y(n48) );
  NAND2BXL U112 ( .AN(B[0]), .B(A[0]), .Y(n62) );
  OAI21XL U113 ( .A0(n6), .A1(n85), .B0(n86), .Y(n84) );
  OR2XL U114 ( .A(n125), .B(n25), .Y(n16) );
  XNOR2X4 U115 ( .A(n17), .B(n126), .Y(DIFF[11]) );
  INVX1 U116 ( .A(n134), .Y(n37) );
  INVX1 U117 ( .A(n123), .Y(n24) );
  INVXL U118 ( .A(n89), .Y(n88) );
  INVX1 U119 ( .A(n48), .Y(n54) );
  NOR2XL U120 ( .A(n41), .B(n37), .Y(n40) );
  INVX1 U121 ( .A(n38), .Y(n41) );
  NAND2BX1 U122 ( .AN(n62), .B(n138), .Y(n141) );
  OAI21XL U123 ( .A0(n56), .A1(n57), .B0(n58), .Y(n49) );
  INVX1 U124 ( .A(n59), .Y(n56) );
  NAND2BXL U125 ( .AN(B[1]), .B(A[1]), .Y(n58) );
  NAND2BXL U126 ( .AN(B[2]), .B(A[2]), .Y(n55) );
  NAND2BXL U127 ( .AN(A[1]), .B(B[1]), .Y(n138) );
  NAND2BXL U128 ( .AN(A[0]), .B(B[0]), .Y(n137) );
  NAND2BX1 U129 ( .AN(B[15]), .B(A[15]), .Y(n69) );
  NOR2BX1 U130 ( .AN(B[13]), .B(A[13]), .Y(n107) );
  XOR2X4 U131 ( .A(n29), .B(n33), .Y(DIFF[6]) );
  CLKINVX3 U132 ( .A(n39), .Y(n36) );
  XOR2X4 U133 ( .A(n49), .B(n53), .Y(DIFF[2]) );
  XOR2X4 U134 ( .A(n63), .B(n64), .Y(DIFF[16]) );
  XOR2X4 U135 ( .A(B[16]), .B(A[16]), .Y(n64) );
  NOR2X4 U136 ( .A(n66), .B(n65), .Y(n63) );
  OAI2BB1X4 U137 ( .A0N(n67), .A1N(n68), .B0(n69), .Y(n66) );
  OAI21X4 U138 ( .A0(n71), .A1(A[13]), .B0(n72), .Y(n70) );
  CLKINVX3 U139 ( .A(n94), .Y(n83) );
  OAI21X4 U140 ( .A0(n101), .A1(n100), .B0(n1), .Y(n98) );
  XOR2X4 U141 ( .A(n104), .B(n105), .Y(DIFF[14]) );
  NOR2X4 U142 ( .A(n109), .B(n110), .Y(n104) );
  XOR2X4 U143 ( .A(n111), .B(n112), .Y(DIFF[13]) );
  NOR2X4 U144 ( .A(n113), .B(n114), .Y(n112) );
  OAI21X4 U145 ( .A0(n115), .A1(n116), .B0(n73), .Y(n111) );
  XOR2X4 U146 ( .A(n117), .B(n115), .Y(DIFF[12]) );
  OAI2BB1X4 U147 ( .A0N(n18), .A1N(n118), .B0(n73), .Y(n117) );
  NAND2BX4 U148 ( .AN(A[11]), .B(B[11]), .Y(n97) );
  XOR2X4 U149 ( .A(n127), .B(n129), .Y(DIFF[10]) );
  NOR2X4 U150 ( .A(n128), .B(n130), .Y(n129) );
  OAI21X4 U151 ( .A0(n131), .A1(n21), .B0(n124), .Y(n127) );
  CLKINVX3 U152 ( .A(n19), .Y(n131) );
  OAI21X4 U153 ( .A0(n25), .A1(n125), .B0(n123), .Y(n19) );
  CLKINVX3 U154 ( .A(n22), .Y(n125) );
  NAND3X4 U155 ( .A(n134), .B(n135), .C(n28), .Y(n133) );
  NAND2X4 U156 ( .A(n6), .B(n90), .Y(n44) );
  NOR2X4 U157 ( .A(n57), .B(n61), .Y(n136) );
  CLKINVX3 U158 ( .A(n85), .Y(n93) );
  NAND4BX4 U159 ( .AN(n37), .B(n45), .C(n28), .D(n31), .Y(n85) );
  NAND2BX4 U160 ( .AN(A[6]), .B(B[6]), .Y(n28) );
  CLKINVX3 U161 ( .A(n142), .Y(n25) );
endmodule


module butterfly_DW01_add_85 ( A, B, SUM );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137;

  OAI21X2 U2 ( .A0(n105), .A1(n106), .B0(n13), .Y(n1) );
  AOI21X4 U3 ( .A0(n24), .A1(n107), .B0(n108), .Y(n105) );
  OR2X4 U4 ( .A(n98), .B(n104), .Y(n2) );
  INVX8 U5 ( .A(n89), .Y(n104) );
  NAND2X2 U6 ( .A(A[11]), .B(B[11]), .Y(n81) );
  BUFX3 U7 ( .A(n90), .Y(n16) );
  NOR2X4 U8 ( .A(n98), .B(n104), .Y(n103) );
  INVX8 U9 ( .A(n99), .Y(n98) );
  CLKBUFX4 U10 ( .A(n100), .Y(n13) );
  NAND3X2 U11 ( .A(n15), .B(n13), .C(n101), .Y(n97) );
  NAND2BX4 U12 ( .AN(B[13]), .B(n3), .Y(n88) );
  CLKINVX20 U13 ( .A(A[13]), .Y(n3) );
  NAND2BX2 U14 ( .AN(n74), .B(n75), .Y(n73) );
  NAND4X2 U15 ( .A(n89), .B(n12), .C(n16), .D(n91), .Y(n74) );
  INVX4 U16 ( .A(n45), .Y(n41) );
  CLKINVX8 U17 ( .A(n80), .Y(n4) );
  INVX8 U18 ( .A(n81), .Y(n80) );
  NAND2XL U19 ( .A(B[4]), .B(A[4]), .Y(n5) );
  NAND2XL U20 ( .A(B[4]), .B(A[4]), .Y(n6) );
  XOR2X2 U21 ( .A(n48), .B(n49), .Y(SUM[5]) );
  OAI21X4 U22 ( .A0(n26), .A1(n50), .B0(n51), .Y(n48) );
  NAND2BX4 U23 ( .AN(B[11]), .B(n7), .Y(n94) );
  CLKINVX20 U24 ( .A(A[11]), .Y(n7) );
  AND2X2 U25 ( .A(A[12]), .B(n27), .Y(n8) );
  NAND2BX4 U26 ( .AN(B[14]), .B(n9), .Y(n90) );
  CLKINVX20 U27 ( .A(A[14]), .Y(n9) );
  NAND2X2 U28 ( .A(n103), .B(n18), .Y(n20) );
  NAND2X2 U29 ( .A(n88), .B(n15), .Y(n115) );
  INVX4 U30 ( .A(n84), .Y(n50) );
  CLKINVX3 U31 ( .A(n87), .Y(n83) );
  OAI2BB1X2 U32 ( .A0N(n27), .A1N(A[12]), .B0(n15), .Y(n108) );
  AND2X2 U33 ( .A(n32), .B(n14), .Y(n10) );
  AND2X4 U34 ( .A(B[13]), .B(A[13]), .Y(n11) );
  NAND2X1 U35 ( .A(B[8]), .B(A[8]), .Y(n34) );
  OR2X4 U36 ( .A(A[8]), .B(B[8]), .Y(n95) );
  XOR2X2 U37 ( .A(n32), .B(n33), .Y(SUM[8]) );
  OR2X4 U38 ( .A(A[3]), .B(B[3]), .Y(n57) );
  NAND2X1 U39 ( .A(B[3]), .B(A[3]), .Y(n55) );
  INVX4 U40 ( .A(n48), .Y(n46) );
  NAND2X2 U41 ( .A(n130), .B(n34), .Y(n28) );
  NOR2BX4 U42 ( .AN(n38), .B(n39), .Y(n37) );
  INVX4 U43 ( .A(n134), .Y(n39) );
  OAI211X2 U44 ( .A0(n31), .A1(n34), .B0(n30), .C0(n122), .Y(n121) );
  NAND3X2 U45 ( .A(n109), .B(n4), .C(n82), .Y(n117) );
  NAND2X4 U46 ( .A(n72), .B(n73), .Y(n70) );
  NAND3XL U47 ( .A(A[12]), .B(n88), .C(n27), .Y(n101) );
  OR2X1 U48 ( .A(A[12]), .B(n27), .Y(n22) );
  BUFX8 U49 ( .A(n88), .Y(n12) );
  NAND3X4 U50 ( .A(n109), .B(n4), .C(n82), .Y(n107) );
  AND2X2 U51 ( .A(n89), .B(n16), .Y(n96) );
  NAND2X4 U52 ( .A(n27), .B(A[12]), .Y(n119) );
  BUFX16 U53 ( .A(B[12]), .Y(n27) );
  NAND3X4 U54 ( .A(n10), .B(n94), .C(n93), .Y(n109) );
  NAND3X1 U55 ( .A(n4), .B(n82), .C(n109), .Y(n113) );
  AND2X1 U56 ( .A(n95), .B(n92), .Y(n14) );
  INVX8 U57 ( .A(n11), .Y(n15) );
  OR2X4 U58 ( .A(A[12]), .B(n27), .Y(n23) );
  INVX4 U59 ( .A(n93), .Y(n128) );
  NAND4BBX4 U60 ( .AN(n25), .BN(n26), .C(n45), .D(n134), .Y(n87) );
  NAND2BX4 U61 ( .AN(n39), .B(n131), .Y(n86) );
  OAI21X4 U62 ( .A0(n129), .A1(n31), .B0(n30), .Y(n125) );
  INVX4 U63 ( .A(n28), .Y(n129) );
  NAND2X4 U64 ( .A(B[9]), .B(A[9]), .Y(n30) );
  NAND2X2 U65 ( .A(B[7]), .B(A[7]), .Y(n38) );
  AND2X4 U66 ( .A(n114), .B(n15), .Y(n111) );
  NAND2X2 U67 ( .A(B[15]), .B(A[15]), .Y(n99) );
  NAND2X4 U68 ( .A(n8), .B(n88), .Y(n114) );
  NAND3X2 U69 ( .A(n88), .B(n22), .C(n113), .Y(n112) );
  NAND2X4 U70 ( .A(n32), .B(n95), .Y(n130) );
  NAND3X2 U71 ( .A(n132), .B(n42), .C(n38), .Y(n131) );
  NAND2X4 U72 ( .A(n2), .B(n1), .Y(n19) );
  XOR2X4 U73 ( .A(n110), .B(n17), .Y(SUM[14]) );
  AND2X4 U74 ( .A(n90), .B(n100), .Y(n17) );
  XOR2X2 U75 ( .A(n28), .B(n29), .Y(SUM[9]) );
  NOR2BX2 U76 ( .AN(n30), .B(n31), .Y(n29) );
  INVX4 U77 ( .A(n92), .Y(n31) );
  OR2X4 U78 ( .A(A[12]), .B(n27), .Y(n91) );
  AOI21X4 U79 ( .A0(n96), .A1(n97), .B0(n98), .Y(n72) );
  NAND2X2 U80 ( .A(n90), .B(n12), .Y(n106) );
  NAND2X4 U81 ( .A(n111), .B(n112), .Y(n110) );
  NOR2BX2 U82 ( .AN(n34), .B(n35), .Y(n33) );
  NOR2X2 U83 ( .A(A[5]), .B(B[5]), .Y(n25) );
  NAND2X2 U84 ( .A(B[5]), .B(A[5]), .Y(n47) );
  NOR2BX2 U85 ( .AN(n47), .B(n25), .Y(n49) );
  NAND2X2 U86 ( .A(n94), .B(n81), .Y(n123) );
  OAI21X4 U87 ( .A0(n105), .A1(n106), .B0(n13), .Y(n102) );
  NAND2X2 U88 ( .A(B[14]), .B(A[14]), .Y(n100) );
  OR2X4 U89 ( .A(B[15]), .B(A[15]), .Y(n89) );
  XOR2X2 U90 ( .A(n43), .B(n44), .Y(SUM[6]) );
  OAI21X2 U91 ( .A0(n46), .A1(n25), .B0(n47), .Y(n43) );
  XOR2X2 U92 ( .A(B[16]), .B(A[16]), .Y(n71) );
  CLKINVX4 U93 ( .A(n102), .Y(n18) );
  XOR2X4 U94 ( .A(n70), .B(n71), .Y(SUM[16]) );
  INVX4 U95 ( .A(n119), .Y(n118) );
  XOR2X4 U96 ( .A(n123), .B(n124), .Y(SUM[11]) );
  AOI21X2 U97 ( .A0(n93), .A1(n125), .B0(n126), .Y(n124) );
  NAND3BX4 U98 ( .AN(n25), .B(n133), .C(n45), .Y(n132) );
  XNOR2X4 U99 ( .A(n107), .B(n120), .Y(SUM[12]) );
  NAND2X4 U100 ( .A(n119), .B(n91), .Y(n120) );
  AOI21X4 U101 ( .A0(n117), .A1(n23), .B0(n118), .Y(n116) );
  NAND3X4 U102 ( .A(n94), .B(n93), .C(n121), .Y(n82) );
  XOR2X4 U103 ( .A(n115), .B(n116), .Y(SUM[13]) );
  NAND2X4 U104 ( .A(B[10]), .B(A[10]), .Y(n122) );
  INVX2 U105 ( .A(n43), .Y(n40) );
  NOR2X4 U106 ( .A(A[4]), .B(B[4]), .Y(n26) );
  NAND2X4 U107 ( .A(n19), .B(n20), .Y(SUM[15]) );
  INVX4 U108 ( .A(n64), .Y(n68) );
  OAI21X4 U109 ( .A0(n50), .A1(n87), .B0(n86), .Y(n32) );
  INVXL U110 ( .A(n86), .Y(n85) );
  NOR2BX1 U111 ( .AN(n42), .B(n41), .Y(n44) );
  OAI211X2 U112 ( .A0(n136), .A1(n137), .B0(n63), .C0(n57), .Y(n135) );
  OAI21X2 U113 ( .A0(n68), .A1(n69), .B0(n66), .Y(n136) );
  CLKINVX4 U114 ( .A(n60), .Y(n137) );
  OAI21XL U115 ( .A0(n58), .A1(n59), .B0(n60), .Y(n53) );
  INVX2 U116 ( .A(n61), .Y(n58) );
  XOR2X1 U117 ( .A(n61), .B(n62), .Y(SUM[2]) );
  INVXL U118 ( .A(n57), .Y(n56) );
  XOR2X1 U119 ( .A(n65), .B(n67), .Y(SUM[1]) );
  NAND2XL U120 ( .A(B[4]), .B(A[4]), .Y(n51) );
  NAND2XL U121 ( .A(B[1]), .B(A[1]), .Y(n66) );
  OR2X4 U122 ( .A(A[9]), .B(B[9]), .Y(n92) );
  OR2XL U123 ( .A(A[2]), .B(B[2]), .Y(n63) );
  NAND2X1 U124 ( .A(B[0]), .B(A[0]), .Y(n69) );
  NOR2BX1 U125 ( .AN(n69), .B(n21), .Y(SUM[0]) );
  NOR2XL U126 ( .A(A[0]), .B(B[0]), .Y(n21) );
  INVX1 U127 ( .A(n122), .Y(n126) );
  NAND2X1 U128 ( .A(n47), .B(n5), .Y(n133) );
  XOR2X2 U129 ( .A(n36), .B(n37), .Y(SUM[7]) );
  OAI21X1 U130 ( .A0(n40), .A1(n41), .B0(n42), .Y(n36) );
  INVXL U131 ( .A(n95), .Y(n35) );
  NAND2X2 U132 ( .A(n55), .B(n135), .Y(n84) );
  OAI21X1 U133 ( .A0(n76), .A1(n77), .B0(n78), .Y(n75) );
  AOI21XL U134 ( .A0(n83), .A1(n84), .B0(n85), .Y(n76) );
  NAND4BXL U135 ( .AN(n35), .B(n92), .C(n93), .D(n94), .Y(n77) );
  NOR2X1 U136 ( .A(n79), .B(n80), .Y(n78) );
  INVX1 U137 ( .A(n63), .Y(n59) );
  XOR2X2 U138 ( .A(n53), .B(n54), .Y(SUM[3]) );
  NOR2BX1 U139 ( .AN(n55), .B(n56), .Y(n54) );
  XOR2X1 U140 ( .A(n84), .B(n52), .Y(SUM[4]) );
  NOR2BX1 U141 ( .AN(n6), .B(n26), .Y(n52) );
  NOR2BX1 U142 ( .AN(n60), .B(n59), .Y(n62) );
  NOR2BXL U143 ( .AN(n66), .B(n68), .Y(n67) );
  OAI2BB1X1 U144 ( .A0N(n64), .A1N(n65), .B0(n66), .Y(n61) );
  INVX1 U145 ( .A(n69), .Y(n65) );
  OR2X2 U146 ( .A(A[7]), .B(B[7]), .Y(n134) );
  OR2XL U147 ( .A(A[12]), .B(n27), .Y(n24) );
  NAND2X1 U148 ( .A(B[6]), .B(A[6]), .Y(n42) );
  NAND2X2 U149 ( .A(B[2]), .B(A[2]), .Y(n60) );
  OR2X2 U150 ( .A(A[1]), .B(B[1]), .Y(n64) );
  INVXL U151 ( .A(n82), .Y(n79) );
  XOR2X4 U152 ( .A(n125), .B(n127), .Y(SUM[10]) );
  NOR2BX4 U153 ( .AN(n122), .B(n128), .Y(n127) );
  OR2X4 U154 ( .A(A[10]), .B(B[10]), .Y(n93) );
  OR2X4 U155 ( .A(A[6]), .B(B[6]), .Y(n45) );
endmodule


module butterfly_DW01_sub_69 ( A, B, DIFF );
  input [16:0] A;
  input [16:0] B;
  output [16:0] DIFF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145;

  CLKINVX8 U3 ( .A(B[12]), .Y(n20) );
  CLKINVX8 U4 ( .A(n20), .Y(n19) );
  CLKINVX8 U5 ( .A(n20), .Y(n18) );
  OR2X4 U6 ( .A(B[15]), .B(n1), .Y(n97) );
  CLKINVX20 U7 ( .A(A[15]), .Y(n1) );
  NAND3X2 U8 ( .A(n12), .B(n118), .C(n101), .Y(n98) );
  NAND2BX1 U9 ( .AN(A[13]), .B(B[13]), .Y(n118) );
  OAI21X2 U10 ( .A0(n107), .A1(n115), .B0(n102), .Y(n114) );
  NAND2X2 U11 ( .A(n2), .B(B[14]), .Y(n87) );
  CLKINVX20 U12 ( .A(A[14]), .Y(n2) );
  OAI21X2 U13 ( .A0(n105), .A1(n106), .B0(n12), .Y(n104) );
  XNOR2X4 U14 ( .A(B[16]), .B(A[16]), .Y(n68) );
  NAND3BX4 U15 ( .AN(n72), .B(n73), .C(n74), .Y(n71) );
  CLKINVX8 U16 ( .A(n26), .Y(n126) );
  OAI2BB1X4 U17 ( .A0N(n82), .A1N(n46), .B0(n85), .Y(n26) );
  CLKINVX4 U18 ( .A(n90), .Y(n82) );
  NOR2X1 U19 ( .A(n76), .B(n90), .Y(n89) );
  NAND2X2 U20 ( .A(n86), .B(n123), .Y(n122) );
  INVX8 U21 ( .A(n97), .Y(n96) );
  OAI2BB1X4 U22 ( .A0N(n3), .A1N(n18), .B0(n116), .Y(n110) );
  CLKINVX20 U23 ( .A(A[12]), .Y(n3) );
  NOR2X2 U24 ( .A(n9), .B(n110), .Y(n105) );
  NAND2BX4 U25 ( .AN(B[14]), .B(A[14]), .Y(n99) );
  INVX4 U26 ( .A(n81), .Y(n78) );
  NOR2BX4 U27 ( .AN(n80), .B(n78), .Y(n117) );
  NAND2BX4 U28 ( .AN(n19), .B(A[12]), .Y(n108) );
  NAND2BX4 U29 ( .AN(n19), .B(A[12]), .Y(n115) );
  NAND2BX4 U30 ( .AN(A[15]), .B(B[15]), .Y(n74) );
  NAND2BX4 U31 ( .AN(A[13]), .B(B[13]), .Y(n116) );
  OR2X4 U32 ( .A(B[13]), .B(n4), .Y(n102) );
  CLKINVX20 U33 ( .A(A[13]), .Y(n4) );
  INVX2 U34 ( .A(n5), .Y(n29) );
  INVX1 U35 ( .A(n109), .Y(n8) );
  INVX1 U36 ( .A(A[8]), .Y(n6) );
  INVX4 U37 ( .A(n91), .Y(n24) );
  NAND2X2 U38 ( .A(n35), .B(n36), .Y(n30) );
  INVX1 U39 ( .A(n32), .Y(n37) );
  NOR2X2 U40 ( .A(B[8]), .B(n6), .Y(n5) );
  NOR2X4 U41 ( .A(n135), .B(n133), .Y(n134) );
  NAND2BX2 U42 ( .AN(A[8]), .B(B[8]), .Y(n145) );
  NAND2BX4 U43 ( .AN(B[5]), .B(A[5]), .Y(n41) );
  NAND2BX2 U44 ( .AN(A[5]), .B(B[5]), .Y(n139) );
  NAND2BX2 U45 ( .AN(A[3]), .B(B[3]), .Y(n53) );
  NAND2BX2 U46 ( .AN(B[3]), .B(A[3]), .Y(n54) );
  NAND3X1 U47 ( .A(n50), .B(n142), .C(n53), .Y(n141) );
  NAND4X2 U48 ( .A(n66), .B(n64), .C(n50), .D(n53), .Y(n94) );
  NAND2X1 U49 ( .A(n53), .B(n54), .Y(n48) );
  NAND2BX4 U50 ( .AN(B[6]), .B(A[6]), .Y(n38) );
  NAND3X2 U51 ( .A(n138), .B(n38), .C(n36), .Y(n137) );
  INVX4 U52 ( .A(n38), .Y(n34) );
  XNOR2X4 U53 ( .A(n123), .B(n124), .Y(DIFF[12]) );
  NOR2X4 U54 ( .A(n7), .B(n8), .Y(n9) );
  INVX4 U55 ( .A(n117), .Y(n7) );
  XOR2X4 U56 ( .A(n130), .B(n131), .Y(DIFF[11]) );
  NOR2X4 U57 ( .A(n95), .B(n96), .Y(n69) );
  AOI21X4 U58 ( .A0(n98), .A1(n11), .B0(n100), .Y(n95) );
  NAND3X1 U59 ( .A(n116), .B(n86), .C(n12), .Y(n72) );
  BUFX12 U60 ( .A(n87), .Y(n12) );
  INVX8 U61 ( .A(n10), .Y(n11) );
  NAND3X4 U62 ( .A(n129), .B(n91), .C(n92), .Y(n127) );
  NAND2X4 U63 ( .A(n11), .B(n12), .Y(n111) );
  NAND4BX4 U64 ( .AN(n24), .B(n125), .C(n92), .D(n93), .Y(n109) );
  INVX4 U65 ( .A(n74), .Y(n100) );
  NAND2BX4 U66 ( .AN(A[1]), .B(B[1]), .Y(n64) );
  OAI21X2 U67 ( .A0(n58), .A1(n59), .B0(n60), .Y(n51) );
  INVX4 U68 ( .A(n64), .Y(n59) );
  NAND2BX4 U69 ( .AN(B[1]), .B(A[1]), .Y(n60) );
  INVX4 U70 ( .A(n21), .Y(n136) );
  NAND3X4 U71 ( .A(n69), .B(n70), .C(n71), .Y(n67) );
  NAND4X2 U72 ( .A(n16), .B(n88), .C(n116), .D(n89), .Y(n70) );
  NAND2X1 U73 ( .A(n115), .B(n102), .Y(n101) );
  NAND2X2 U74 ( .A(n104), .B(n11), .Y(n103) );
  NOR2X1 U75 ( .A(n5), .B(n28), .Y(n27) );
  CLKINVX4 U76 ( .A(n145), .Y(n28) );
  XOR2X2 U77 ( .A(n21), .B(n22), .Y(DIFF[9]) );
  XOR2X2 U78 ( .A(n26), .B(n27), .Y(DIFF[8]) );
  OAI21X2 U79 ( .A0(n107), .A1(n108), .B0(n102), .Y(n106) );
  CLKINVX8 U80 ( .A(n99), .Y(n10) );
  XNOR2X4 U81 ( .A(n120), .B(n121), .Y(DIFF[13]) );
  NAND2BX4 U82 ( .AN(B[7]), .B(A[7]), .Y(n36) );
  NOR2X1 U83 ( .A(n126), .B(n28), .Y(n125) );
  INVX3 U84 ( .A(n116), .Y(n107) );
  NAND2X2 U85 ( .A(n25), .B(n29), .Y(n129) );
  OAI21X4 U86 ( .A0(n28), .A1(n126), .B0(n29), .Y(n21) );
  AND3X2 U87 ( .A(n74), .B(n86), .C(n12), .Y(n16) );
  INVX4 U88 ( .A(n25), .Y(n23) );
  OAI21X4 U89 ( .A0(n136), .A1(n24), .B0(n25), .Y(n132) );
  NAND2BX4 U90 ( .AN(B[9]), .B(A[9]), .Y(n25) );
  INVX8 U91 ( .A(n128), .Y(n133) );
  NAND2BX4 U92 ( .AN(B[10]), .B(A[10]), .Y(n128) );
  NAND2X2 U93 ( .A(n118), .B(n102), .Y(n121) );
  NOR2X4 U94 ( .A(n113), .B(n114), .Y(n112) );
  NAND2BX4 U95 ( .AN(n83), .B(n94), .Y(n46) );
  XOR2X2 U96 ( .A(n30), .B(n31), .Y(DIFF[7]) );
  AOI21X2 U97 ( .A0(n32), .A1(n33), .B0(n34), .Y(n31) );
  OAI21X2 U98 ( .A0(n39), .A1(n40), .B0(n41), .Y(n33) );
  INVX2 U99 ( .A(n42), .Y(n39) );
  NAND2BX4 U100 ( .AN(A[2]), .B(B[2]), .Y(n50) );
  NAND2X4 U101 ( .A(n127), .B(n128), .Y(n119) );
  NAND2BX4 U102 ( .AN(A[9]), .B(B[9]), .Y(n91) );
  NAND3X2 U103 ( .A(n81), .B(n80), .C(n109), .Y(n123) );
  NAND2BX4 U104 ( .AN(B[11]), .B(A[11]), .Y(n80) );
  NAND2X4 U105 ( .A(n93), .B(n119), .Y(n81) );
  XNOR2X4 U106 ( .A(n103), .B(n13), .Y(DIFF[15]) );
  XOR2X4 U107 ( .A(n111), .B(n112), .Y(DIFF[14]) );
  XOR2X4 U108 ( .A(n67), .B(n68), .Y(DIFF[16]) );
  NAND4BX1 U109 ( .AN(n28), .B(n91), .C(n92), .D(n93), .Y(n76) );
  INVX4 U110 ( .A(n92), .Y(n135) );
  NAND2BX4 U111 ( .AN(A[10]), .B(B[10]), .Y(n92) );
  AOI21X2 U112 ( .A0(n92), .A1(n132), .B0(n133), .Y(n131) );
  NOR2X1 U113 ( .A(n34), .B(n37), .Y(n15) );
  NAND2X2 U114 ( .A(n46), .B(n47), .Y(n44) );
  NAND2X2 U115 ( .A(n93), .B(n80), .Y(n130) );
  NOR2XL U116 ( .A(n43), .B(n40), .Y(n14) );
  NAND2X1 U117 ( .A(n144), .B(n64), .Y(n143) );
  NAND3X1 U118 ( .A(n139), .B(n140), .C(n32), .Y(n138) );
  XOR2X1 U119 ( .A(n33), .B(n15), .Y(DIFF[6]) );
  NOR2X1 U120 ( .A(n52), .B(n56), .Y(n55) );
  XOR2X1 U121 ( .A(n46), .B(n17), .Y(DIFF[4]) );
  OR2X4 U122 ( .A(n100), .B(n96), .Y(n13) );
  XOR2X1 U123 ( .A(n42), .B(n14), .Y(DIFF[5]) );
  NAND2X2 U124 ( .A(n35), .B(n137), .Y(n85) );
  NAND4BX2 U125 ( .AN(n40), .B(n47), .C(n32), .D(n35), .Y(n90) );
  NAND2X2 U126 ( .A(n141), .B(n54), .Y(n83) );
  INVXL U127 ( .A(n57), .Y(n52) );
  XOR2X1 U128 ( .A(n51), .B(n55), .Y(DIFF[2]) );
  XOR2X1 U129 ( .A(n48), .B(n49), .Y(DIFF[3]) );
  NAND2XL U130 ( .A(n66), .B(n65), .Y(DIFF[0]) );
  NAND2BXL U131 ( .AN(A[4]), .B(B[4]), .Y(n47) );
  NAND2BXL U132 ( .AN(B[4]), .B(A[4]), .Y(n45) );
  NAND2BXL U133 ( .AN(B[0]), .B(A[0]), .Y(n65) );
  OAI21XL U134 ( .A0(n75), .A1(n76), .B0(n77), .Y(n73) );
  AOI21XL U135 ( .A0(n82), .A1(n83), .B0(n84), .Y(n75) );
  NOR2X1 U136 ( .A(n78), .B(n79), .Y(n77) );
  INVX1 U137 ( .A(n85), .Y(n84) );
  XOR2X2 U138 ( .A(n132), .B(n134), .Y(DIFF[10]) );
  NOR2X2 U139 ( .A(n23), .B(n24), .Y(n22) );
  INVX1 U140 ( .A(n94), .Y(n88) );
  INVX1 U141 ( .A(n139), .Y(n40) );
  NAND2X1 U142 ( .A(n41), .B(n45), .Y(n140) );
  INVX1 U143 ( .A(n80), .Y(n79) );
  INVX1 U144 ( .A(n50), .Y(n56) );
  AOI21X1 U145 ( .A0(n50), .A1(n51), .B0(n52), .Y(n49) );
  XOR2X1 U146 ( .A(n61), .B(n62), .Y(DIFF[1]) );
  NOR2X1 U147 ( .A(n63), .B(n59), .Y(n62) );
  INVX1 U148 ( .A(n60), .Y(n63) );
  AND2X2 U149 ( .A(n45), .B(n47), .Y(n17) );
  NAND2X2 U150 ( .A(n44), .B(n45), .Y(n42) );
  NAND3X1 U151 ( .A(n143), .B(n60), .C(n57), .Y(n142) );
  INVX1 U152 ( .A(n61), .Y(n58) );
  NAND2BX1 U153 ( .AN(n66), .B(n65), .Y(n61) );
  INVX1 U154 ( .A(n65), .Y(n144) );
  NAND2BXL U155 ( .AN(B[2]), .B(A[2]), .Y(n57) );
  NAND2BXL U156 ( .AN(A[0]), .B(B[0]), .Y(n66) );
  NAND2X2 U157 ( .A(n122), .B(n115), .Y(n120) );
  AOI21X2 U158 ( .A0(n117), .A1(n109), .B0(n110), .Y(n113) );
  CLKINVX3 U159 ( .A(n41), .Y(n43) );
  NAND2X4 U160 ( .A(n108), .B(n86), .Y(n124) );
  NAND2BX4 U161 ( .AN(A[12]), .B(n18), .Y(n86) );
  NAND2BX4 U162 ( .AN(A[11]), .B(B[11]), .Y(n93) );
  NAND2BX4 U163 ( .AN(A[7]), .B(B[7]), .Y(n35) );
  NAND2BX4 U164 ( .AN(A[6]), .B(B[6]), .Y(n32) );
endmodule


module butterfly_DW01_sub_71 ( A, B, DIFF );
  input [16:0] A;
  input [16:0] B;
  output [16:0] DIFF;
  wire   n161, n162, n163, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n33, n34, n35, n36, n37, n38, n39, n40, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160;

  INVX2 U3 ( .A(n101), .Y(n23) );
  INVX3 U4 ( .A(A[13]), .Y(n22) );
  CLKINVX3 U5 ( .A(n128), .Y(n8) );
  XNOR2X4 U6 ( .A(n119), .B(n1), .Y(n161) );
  NAND2X4 U7 ( .A(n92), .B(n109), .Y(n1) );
  CLKINVX4 U8 ( .A(n16), .Y(n144) );
  BUFX4 U9 ( .A(A[11]), .Y(n7) );
  BUFX20 U10 ( .A(n163), .Y(DIFF[7]) );
  INVX3 U11 ( .A(n133), .Y(n2) );
  BUFX8 U12 ( .A(B[10]), .Y(n3) );
  NOR2BX4 U13 ( .AN(n9), .B(n122), .Y(n121) );
  OAI21X2 U14 ( .A0(n145), .A1(n146), .B0(n138), .Y(n142) );
  OAI21X1 U15 ( .A0(n93), .A1(n2), .B0(n95), .Y(n90) );
  NOR2X2 U16 ( .A(n100), .B(n101), .Y(n89) );
  NAND3X2 U17 ( .A(n153), .B(n154), .C(n52), .Y(n152) );
  INVX4 U18 ( .A(n108), .Y(n135) );
  INVX2 U19 ( .A(n109), .Y(n100) );
  NOR2X2 U20 ( .A(n80), .B(n84), .Y(n155) );
  XNOR2X2 U21 ( .A(n47), .B(n26), .Y(n25) );
  XOR2X4 U22 ( .A(n69), .B(n70), .Y(DIFF[3]) );
  NAND2BX2 U23 ( .AN(A[11]), .B(B[11]), .Y(n115) );
  NAND2BX4 U24 ( .AN(A[10]), .B(n3), .Y(n114) );
  BUFX8 U25 ( .A(B[9]), .Y(n4) );
  NAND2BX4 U26 ( .AN(n18), .B(n115), .Y(n129) );
  BUFX8 U27 ( .A(A[15]), .Y(n19) );
  NOR2X4 U28 ( .A(n101), .B(n123), .Y(n122) );
  NAND4BX4 U29 ( .AN(n101), .B(n14), .C(n12), .D(n125), .Y(n120) );
  NAND2BX4 U30 ( .AN(A[12]), .B(n6), .Y(n124) );
  INVX4 U31 ( .A(n138), .Y(n148) );
  XNOR2X2 U32 ( .A(n43), .B(n44), .Y(n5) );
  CLKINVX20 U33 ( .A(n5), .Y(DIFF[9]) );
  BUFX8 U34 ( .A(B[12]), .Y(n6) );
  BUFX12 U35 ( .A(B[13]), .Y(n24) );
  INVX2 U36 ( .A(n9), .Y(n97) );
  NAND2BX4 U37 ( .AN(B[14]), .B(n11), .Y(n9) );
  INVX8 U38 ( .A(n113), .Y(n46) );
  AND2X4 U39 ( .A(n10), .B(n124), .Y(n127) );
  NAND2X4 U40 ( .A(n24), .B(n22), .Y(n10) );
  BUFX8 U41 ( .A(A[14]), .Y(n11) );
  INVX4 U42 ( .A(n52), .Y(n58) );
  INVXL U43 ( .A(n135), .Y(n12) );
  AOI21X2 U44 ( .A0(n89), .A1(n90), .B0(n91), .Y(n88) );
  INVX8 U45 ( .A(n111), .Y(n128) );
  CLKINVX4 U46 ( .A(n93), .Y(n14) );
  INVX3 U47 ( .A(n99), .Y(n93) );
  AND4X4 U48 ( .A(n109), .B(n23), .C(n124), .D(n14), .Y(n15) );
  NAND3X4 U49 ( .A(n71), .B(n74), .C(n155), .Y(n104) );
  NAND2BX4 U50 ( .AN(A[11]), .B(B[11]), .Y(n16) );
  NAND2BX4 U51 ( .AN(A[1]), .B(B[1]), .Y(n157) );
  NAND2BX4 U52 ( .AN(B[1]), .B(A[1]), .Y(n81) );
  INVX4 U53 ( .A(n140), .Y(n45) );
  INVX8 U54 ( .A(n94), .Y(n133) );
  NAND2BX4 U55 ( .AN(A[10]), .B(n3), .Y(n17) );
  INVX3 U56 ( .A(n123), .Y(n96) );
  INVX8 U57 ( .A(n141), .Y(n49) );
  NAND3X2 U58 ( .A(n47), .B(n17), .C(n28), .Y(n18) );
  NAND4BX4 U59 ( .AN(n128), .B(n94), .C(n110), .D(n129), .Y(n125) );
  NAND3X4 U60 ( .A(n136), .B(n16), .C(n17), .Y(n110) );
  NAND2X4 U61 ( .A(n156), .B(n85), .Y(DIFF[0]) );
  NAND2BX4 U62 ( .AN(B[0]), .B(A[0]), .Y(n85) );
  XNOR2X4 U63 ( .A(B[16]), .B(A[16]), .Y(n21) );
  XNOR2X4 U64 ( .A(n147), .B(n29), .Y(n33) );
  INVX4 U65 ( .A(n47), .Y(n150) );
  NAND2BX4 U66 ( .AN(B[14]), .B(n11), .Y(n98) );
  AOI21X4 U67 ( .A0(n132), .A1(n124), .B0(n133), .Y(n131) );
  BUFX20 U68 ( .A(n162), .Y(DIFF[13]) );
  INVX4 U69 ( .A(n43), .Y(n149) );
  INVX4 U70 ( .A(n147), .Y(n145) );
  INVX4 U71 ( .A(n114), .Y(n146) );
  NOR2X2 U72 ( .A(n96), .B(n97), .Y(n95) );
  NAND2BX4 U73 ( .AN(B[15]), .B(n19), .Y(n92) );
  NAND3X4 U74 ( .A(n129), .B(n8), .C(n110), .Y(n132) );
  NAND4BX4 U75 ( .AN(n104), .B(n36), .C(n102), .D(n15), .Y(n87) );
  XOR2X4 U76 ( .A(n20), .B(n21), .Y(DIFF[16]) );
  NAND3X4 U77 ( .A(n86), .B(n87), .C(n88), .Y(n20) );
  INVX8 U78 ( .A(n25), .Y(DIFF[8]) );
  BUFX20 U79 ( .A(n161), .Y(DIFF[15]) );
  NAND2BX4 U80 ( .AN(A[4]), .B(B[4]), .Y(n68) );
  XOR2X4 U81 ( .A(n130), .B(n131), .Y(n162) );
  NAND2BX4 U82 ( .AN(A[5]), .B(B[5]), .Y(n153) );
  NAND2BX4 U83 ( .AN(B[3]), .B(A[3]), .Y(n75) );
  AOI21X1 U84 ( .A0(n71), .A1(n72), .B0(n73), .Y(n70) );
  INVX8 U85 ( .A(n33), .Y(DIFF[10]) );
  XOR2X4 U86 ( .A(n72), .B(n76), .Y(DIFF[2]) );
  OAI21X2 U87 ( .A0(n105), .A1(n106), .B0(n15), .Y(n86) );
  NAND2X4 U88 ( .A(n55), .B(n151), .Y(n118) );
  NAND3X4 U89 ( .A(n152), .B(n59), .C(n56), .Y(n151) );
  NAND2BX4 U90 ( .AN(B[5]), .B(A[5]), .Y(n62) );
  XNOR2X4 U91 ( .A(n82), .B(n27), .Y(DIFF[1]) );
  NAND2BX4 U92 ( .AN(A[3]), .B(B[3]), .Y(n74) );
  NAND2BX4 U93 ( .AN(B[4]), .B(A[4]), .Y(n66) );
  NAND2X2 U94 ( .A(n55), .B(n56), .Y(n50) );
  AOI21X2 U95 ( .A0(n52), .A1(n53), .B0(n54), .Y(n51) );
  OAI21X4 U96 ( .A0(n79), .A1(n80), .B0(n81), .Y(n72) );
  OR2X4 U97 ( .A(n83), .B(n80), .Y(n27) );
  NAND2XL U98 ( .A(n62), .B(n66), .Y(n154) );
  NAND2BX4 U99 ( .AN(B[9]), .B(A[9]), .Y(n140) );
  NOR2X4 U100 ( .A(n48), .B(n49), .Y(n26) );
  INVX4 U101 ( .A(n153), .Y(n61) );
  INVX8 U102 ( .A(n34), .Y(DIFF[11]) );
  NAND2X4 U103 ( .A(n99), .B(n123), .Y(n130) );
  NAND2BXL U104 ( .AN(A[0]), .B(B[0]), .Y(n156) );
  OAI2BB1X4 U105 ( .A0N(n36), .A1N(n67), .B0(n118), .Y(n47) );
  INVXL U106 ( .A(n118), .Y(n117) );
  INVX4 U107 ( .A(n157), .Y(n80) );
  AND2X1 U108 ( .A(n141), .B(n113), .Y(n28) );
  INVX4 U109 ( .A(n78), .Y(n73) );
  OR2X4 U110 ( .A(n64), .B(n61), .Y(n39) );
  NAND2X4 U111 ( .A(n84), .B(n85), .Y(n82) );
  NAND2X4 U112 ( .A(n67), .B(n68), .Y(n65) );
  INVXL U113 ( .A(n61), .Y(n37) );
  INVX4 U114 ( .A(n142), .Y(n35) );
  NOR2X4 U115 ( .A(n148), .B(n146), .Y(n29) );
  NAND3BXL U116 ( .AN(n30), .B(n81), .C(n78), .Y(n159) );
  AND2X1 U117 ( .A(n160), .B(n157), .Y(n30) );
  XNOR2X4 U118 ( .A(n126), .B(n31), .Y(n40) );
  NAND2X2 U119 ( .A(n107), .B(n98), .Y(n31) );
  XOR2X4 U120 ( .A(n134), .B(n132), .Y(DIFF[12]) );
  NAND2BX4 U121 ( .AN(B[10]), .B(A[10]), .Y(n138) );
  NAND2BX4 U122 ( .AN(B[7]), .B(A[7]), .Y(n56) );
  NAND2BX4 U123 ( .AN(n116), .B(n104), .Y(n67) );
  XOR2X4 U124 ( .A(n143), .B(n35), .Y(n34) );
  AND4X4 U125 ( .A(n37), .B(n68), .C(n52), .D(n55), .Y(n36) );
  NAND2XL U126 ( .A(n110), .B(n111), .Y(n106) );
  NOR2XL U127 ( .A(n112), .B(n103), .Y(n105) );
  AOI21XL U128 ( .A0(n36), .A1(n116), .B0(n117), .Y(n112) );
  INVXL U129 ( .A(n71), .Y(n77) );
  XOR2X4 U130 ( .A(n67), .B(n38), .Y(DIFF[4]) );
  AND2X2 U131 ( .A(n66), .B(n68), .Y(n38) );
  NAND2X1 U132 ( .A(n74), .B(n75), .Y(n69) );
  XNOR2X4 U133 ( .A(n63), .B(n39), .Y(DIFF[5]) );
  INVX1 U134 ( .A(n81), .Y(n83) );
  INVX1 U135 ( .A(n82), .Y(n79) );
  INVX1 U136 ( .A(n156), .Y(n84) );
  INVX1 U137 ( .A(n85), .Y(n160) );
  NAND3BX2 U138 ( .AN(n45), .B(n137), .C(n138), .Y(n136) );
  NAND2XL U139 ( .A(n48), .B(n113), .Y(n137) );
  INVX8 U140 ( .A(n40), .Y(DIFF[14]) );
  INVX1 U141 ( .A(n92), .Y(n91) );
  NAND2BX4 U142 ( .AN(B[12]), .B(A[12]), .Y(n94) );
  NAND4BXL U143 ( .AN(n49), .B(n113), .C(n17), .D(n115), .Y(n103) );
  NAND2BX4 U144 ( .AN(A[12]), .B(n6), .Y(n108) );
  INVX8 U145 ( .A(n107), .Y(n101) );
  NOR2X4 U146 ( .A(n45), .B(n46), .Y(n44) );
  XOR2X4 U147 ( .A(n50), .B(n51), .Y(n163) );
  XOR2X4 U148 ( .A(n53), .B(n57), .Y(DIFF[6]) );
  NOR2X4 U149 ( .A(n54), .B(n58), .Y(n57) );
  CLKINVX3 U150 ( .A(n59), .Y(n54) );
  OAI21X4 U151 ( .A0(n60), .A1(n61), .B0(n62), .Y(n53) );
  CLKINVX3 U152 ( .A(n63), .Y(n60) );
  CLKINVX3 U153 ( .A(n62), .Y(n64) );
  NAND2X4 U154 ( .A(n65), .B(n66), .Y(n63) );
  NOR2X4 U155 ( .A(n73), .B(n77), .Y(n76) );
  CLKINVX3 U156 ( .A(n103), .Y(n102) );
  NAND2BX4 U157 ( .AN(A[15]), .B(B[15]), .Y(n109) );
  NAND2X4 U158 ( .A(n120), .B(n121), .Y(n119) );
  AOI21X4 U159 ( .A0(n127), .A1(n125), .B0(n96), .Y(n126) );
  NAND2BX4 U160 ( .AN(A[14]), .B(B[14]), .Y(n107) );
  NAND2BX4 U161 ( .AN(B[13]), .B(A[13]), .Y(n123) );
  NAND2BX4 U162 ( .AN(A[13]), .B(n24), .Y(n99) );
  NOR2X4 U163 ( .A(n133), .B(n135), .Y(n134) );
  CLKINVX3 U164 ( .A(n139), .Y(n48) );
  NOR2X4 U165 ( .A(n128), .B(n144), .Y(n143) );
  NAND2BX4 U166 ( .AN(B[11]), .B(n7), .Y(n111) );
  OAI21X4 U167 ( .A0(n149), .A1(n46), .B0(n140), .Y(n147) );
  NAND2BX4 U168 ( .AN(A[9]), .B(n4), .Y(n113) );
  OAI21X4 U169 ( .A0(n150), .A1(n49), .B0(n139), .Y(n43) );
  NAND2BX4 U170 ( .AN(B[8]), .B(A[8]), .Y(n139) );
  NAND2BX4 U171 ( .AN(A[8]), .B(B[8]), .Y(n141) );
  NAND2BX4 U172 ( .AN(B[6]), .B(A[6]), .Y(n59) );
  NAND2X4 U173 ( .A(n158), .B(n75), .Y(n116) );
  NAND3X4 U174 ( .A(n71), .B(n159), .C(n74), .Y(n158) );
  NAND2BX4 U175 ( .AN(B[2]), .B(A[2]), .Y(n78) );
  NAND2BX4 U176 ( .AN(A[2]), .B(B[2]), .Y(n71) );
  NAND2BX4 U177 ( .AN(A[7]), .B(B[7]), .Y(n55) );
  NAND2BX4 U178 ( .AN(A[6]), .B(B[6]), .Y(n52) );
endmodule


module butterfly_DW01_add_90 ( A, B, SUM );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132;

  CLKBUFX4 U2 ( .A(A[12]), .Y(n24) );
  BUFX1 U3 ( .A(n86), .Y(n1) );
  NAND2X2 U4 ( .A(n15), .B(n9), .Y(n2) );
  INVX4 U5 ( .A(n14), .Y(n15) );
  INVX4 U6 ( .A(n8), .Y(n9) );
  OAI21XL U7 ( .A0(A[12]), .A1(B[12]), .B0(n90), .Y(n104) );
  NAND2X2 U8 ( .A(B[12]), .B(A[12]), .Y(n114) );
  NAND2X2 U9 ( .A(B[11]), .B(A[11]), .Y(n77) );
  AND2X2 U10 ( .A(n84), .B(n87), .Y(n6) );
  NAND2X2 U11 ( .A(n84), .B(n101), .Y(n113) );
  NAND3X1 U12 ( .A(n3), .B(n24), .C(n84), .Y(n95) );
  INVX2 U13 ( .A(B[14]), .Y(n8) );
  XOR2X2 U14 ( .A(n80), .B(n49), .Y(SUM[4]) );
  BUFX12 U15 ( .A(B[12]), .Y(n3) );
  XOR2X2 U16 ( .A(n45), .B(n46), .Y(SUM[5]) );
  NAND2X4 U17 ( .A(n114), .B(n115), .Y(n112) );
  BUFX8 U18 ( .A(n122), .Y(n4) );
  AND2X2 U19 ( .A(A[15]), .B(B[15]), .Y(n5) );
  NAND2X2 U20 ( .A(B[13]), .B(A[13]), .Y(n101) );
  INVX2 U21 ( .A(n129), .Y(n36) );
  INVX2 U22 ( .A(n45), .Y(n43) );
  XOR2X2 U23 ( .A(n50), .B(n51), .Y(SUM[3]) );
  INVX4 U24 ( .A(n30), .Y(n17) );
  NAND2X2 U25 ( .A(n16), .B(n30), .Y(n19) );
  NOR2BX4 U26 ( .AN(n31), .B(n32), .Y(n30) );
  XOR2X2 U27 ( .A(n33), .B(n34), .Y(SUM[7]) );
  NAND2X1 U28 ( .A(B[6]), .B(A[6]), .Y(n39) );
  NAND3X2 U29 ( .A(n24), .B(n3), .C(n84), .Y(n109) );
  NAND3X2 U30 ( .A(n101), .B(n109), .C(n110), .Y(n12) );
  XOR2X4 U31 ( .A(n25), .B(n26), .Y(SUM[9]) );
  AND2X4 U32 ( .A(n86), .B(n84), .Y(n100) );
  NOR2XL U33 ( .A(A[11]), .B(B[11]), .Y(n118) );
  NAND3X2 U34 ( .A(n90), .B(n89), .C(n107), .Y(n78) );
  AND3X2 U35 ( .A(n1), .B(n85), .C(n6), .Y(n11) );
  NAND2X2 U36 ( .A(B[7]), .B(A[7]), .Y(n35) );
  OAI21X2 U37 ( .A0(n92), .A1(n91), .B0(n85), .Y(n69) );
  NAND2X4 U38 ( .A(n13), .B(n85), .Y(n10) );
  NAND2X4 U39 ( .A(n11), .B(n71), .Y(n70) );
  XNOR2X4 U40 ( .A(n7), .B(n121), .Y(SUM[11]) );
  AND2X4 U41 ( .A(n90), .B(n77), .Y(n7) );
  XNOR2X4 U42 ( .A(n96), .B(n10), .Y(SUM[15]) );
  NAND2X4 U43 ( .A(n2), .B(n97), .Y(n96) );
  NAND2X2 U44 ( .A(B[1]), .B(A[1]), .Y(n63) );
  NAND2X2 U45 ( .A(n111), .B(n87), .Y(n115) );
  NAND2X4 U46 ( .A(n114), .B(n87), .Y(n20) );
  AOI2BB1X1 U47 ( .A0N(n15), .A1N(n9), .B0(n95), .Y(n91) );
  XNOR2X4 U48 ( .A(n12), .B(n108), .Y(SUM[14]) );
  NAND4BX2 U49 ( .AN(n118), .B(n29), .C(n89), .D(n119), .Y(n116) );
  INVX4 U50 ( .A(n5), .Y(n13) );
  NAND2X4 U51 ( .A(n15), .B(n9), .Y(n94) );
  NOR2BX4 U52 ( .AN(n117), .B(n106), .Y(n124) );
  INVX4 U53 ( .A(n89), .Y(n106) );
  CLKINVX2 U54 ( .A(A[14]), .Y(n14) );
  NAND3X1 U55 ( .A(n86), .B(B[13]), .C(A[13]), .Y(n93) );
  OAI211X2 U56 ( .A0(n131), .A1(n132), .B0(n60), .C0(n54), .Y(n130) );
  OR2X4 U57 ( .A(A[3]), .B(B[3]), .Y(n54) );
  OAI21X2 U58 ( .A0(n37), .A1(n38), .B0(n39), .Y(n33) );
  OR2X4 U59 ( .A(A[7]), .B(B[7]), .Y(n129) );
  NAND3X4 U60 ( .A(n70), .B(n13), .C(n69), .Y(n67) );
  XOR2X2 U61 ( .A(B[16]), .B(A[16]), .Y(n68) );
  XOR2X4 U62 ( .A(n4), .B(n124), .Y(SUM[10]) );
  CLKINVX2 U63 ( .A(n29), .Y(n16) );
  NAND2X2 U64 ( .A(n29), .B(n17), .Y(n18) );
  OAI2BB1X4 U65 ( .A0N(n120), .A1N(n29), .B0(n31), .Y(n25) );
  NOR2X2 U66 ( .A(n28), .B(n106), .Y(n105) );
  NAND2X4 U67 ( .A(B[5]), .B(A[5]), .Y(n44) );
  OAI21X4 U68 ( .A0(n125), .A1(n28), .B0(n27), .Y(n122) );
  NAND2X2 U69 ( .A(B[9]), .B(A[9]), .Y(n27) );
  NAND2X2 U70 ( .A(n44), .B(n48), .Y(n128) );
  NAND2X2 U71 ( .A(n2), .B(n93), .Y(n92) );
  OAI21X4 U72 ( .A0(n98), .A1(n99), .B0(n100), .Y(n97) );
  AOI31X4 U73 ( .A0(n102), .A1(n103), .A2(n77), .B0(n104), .Y(n98) );
  XOR2X2 U74 ( .A(n40), .B(n41), .Y(SUM[6]) );
  OR2X4 U75 ( .A(A[13]), .B(B[13]), .Y(n84) );
  NAND3X2 U76 ( .A(n84), .B(n87), .C(n111), .Y(n110) );
  XNOR2X4 U77 ( .A(n111), .B(n20), .Y(SUM[12]) );
  NAND2X4 U78 ( .A(n94), .B(n86), .Y(n108) );
  NAND2X4 U79 ( .A(B[10]), .B(A[10]), .Y(n117) );
  OAI211X2 U80 ( .A0(n28), .A1(n31), .B0(n27), .C0(n117), .Y(n107) );
  INVX8 U81 ( .A(n88), .Y(n28) );
  NAND2X4 U82 ( .A(B[8]), .B(A[8]), .Y(n31) );
  OAI21X2 U83 ( .A0(n55), .A1(n56), .B0(n57), .Y(n50) );
  INVX4 U84 ( .A(n25), .Y(n125) );
  AOI21X2 U85 ( .A0(n89), .A1(n122), .B0(n123), .Y(n121) );
  OR2X4 U86 ( .A(A[15]), .B(B[15]), .Y(n85) );
  OR2X4 U87 ( .A(A[14]), .B(B[14]), .Y(n86) );
  NAND2X4 U88 ( .A(B[2]), .B(A[2]), .Y(n57) );
  OAI21X2 U89 ( .A0(n43), .A1(n22), .B0(n44), .Y(n40) );
  XNOR2X4 U90 ( .A(n112), .B(n113), .Y(SUM[13]) );
  NOR2X1 U91 ( .A(n28), .B(n32), .Y(n119) );
  INVX4 U92 ( .A(n120), .Y(n32) );
  OR2X4 U93 ( .A(A[8]), .B(B[8]), .Y(n120) );
  NOR2X4 U94 ( .A(A[5]), .B(B[5]), .Y(n22) );
  NAND2X4 U95 ( .A(n18), .B(n19), .Y(SUM[8]) );
  INVX4 U96 ( .A(n80), .Y(n47) );
  INVXL U97 ( .A(n66), .Y(n62) );
  OAI21X2 U98 ( .A0(n23), .A1(n47), .B0(n48), .Y(n45) );
  OAI2BB1X1 U99 ( .A0N(n3), .A1N(n24), .B0(n101), .Y(n99) );
  NOR2XL U100 ( .A(A[0]), .B(B[0]), .Y(n21) );
  OAI21X4 U101 ( .A0(n47), .A1(n83), .B0(n82), .Y(n29) );
  INVXL U102 ( .A(n83), .Y(n79) );
  INVXL U103 ( .A(n82), .Y(n81) );
  INVX2 U104 ( .A(n40), .Y(n37) );
  NAND2X2 U105 ( .A(n52), .B(n130), .Y(n80) );
  OAI21X2 U106 ( .A0(n65), .A1(n66), .B0(n63), .Y(n131) );
  INVX4 U107 ( .A(n61), .Y(n65) );
  XOR2X1 U108 ( .A(n58), .B(n59), .Y(SUM[2]) );
  NOR2BXL U109 ( .AN(n57), .B(n56), .Y(n59) );
  NAND2XL U110 ( .A(B[4]), .B(A[4]), .Y(n48) );
  NAND2XL U111 ( .A(B[3]), .B(A[3]), .Y(n52) );
  NOR2XL U112 ( .A(A[4]), .B(B[4]), .Y(n23) );
  OR2X4 U113 ( .A(A[12]), .B(B[12]), .Y(n87) );
  OR2XL U114 ( .A(A[2]), .B(B[2]), .Y(n60) );
  NOR2BX1 U115 ( .AN(n66), .B(n21), .Y(SUM[0]) );
  INVX1 U116 ( .A(n78), .Y(n75) );
  NAND4BBX2 U117 ( .AN(n22), .BN(n23), .C(n42), .D(n129), .Y(n83) );
  INVX1 U118 ( .A(n117), .Y(n123) );
  NAND2BX2 U119 ( .AN(n36), .B(n126), .Y(n82) );
  NAND3X1 U120 ( .A(n127), .B(n39), .C(n35), .Y(n126) );
  NAND3BX1 U121 ( .AN(n22), .B(n128), .C(n42), .Y(n127) );
  INVXL U122 ( .A(n42), .Y(n38) );
  NOR2BX2 U123 ( .AN(n39), .B(n38), .Y(n41) );
  NOR2BX1 U124 ( .AN(n44), .B(n22), .Y(n46) );
  NOR2BXL U125 ( .AN(n35), .B(n36), .Y(n34) );
  OAI21XL U126 ( .A0(n72), .A1(n73), .B0(n74), .Y(n71) );
  AOI21X1 U127 ( .A0(n79), .A1(n80), .B0(n81), .Y(n72) );
  NAND4BXL U128 ( .AN(n32), .B(n88), .C(n89), .D(n90), .Y(n73) );
  NOR2X1 U129 ( .A(n75), .B(n76), .Y(n74) );
  INVX1 U130 ( .A(n57), .Y(n132) );
  INVX1 U131 ( .A(n77), .Y(n76) );
  INVX1 U132 ( .A(n60), .Y(n56) );
  NOR2BX1 U133 ( .AN(n52), .B(n53), .Y(n51) );
  INVX1 U134 ( .A(n58), .Y(n55) );
  NOR2BX1 U135 ( .AN(n48), .B(n23), .Y(n49) );
  XOR2X1 U136 ( .A(n62), .B(n64), .Y(SUM[1]) );
  NOR2BXL U137 ( .AN(n63), .B(n65), .Y(n64) );
  INVX1 U138 ( .A(n54), .Y(n53) );
  OAI2BB1X1 U139 ( .A0N(n61), .A1N(n62), .B0(n63), .Y(n58) );
  NAND2XL U140 ( .A(n107), .B(n89), .Y(n102) );
  NAND3BXL U141 ( .AN(n32), .B(n29), .C(n105), .Y(n103) );
  OR2X2 U142 ( .A(A[1]), .B(B[1]), .Y(n61) );
  NAND2X1 U143 ( .A(B[0]), .B(A[0]), .Y(n66) );
  NOR2BX4 U144 ( .AN(n27), .B(n28), .Y(n26) );
  XOR2X4 U145 ( .A(n67), .B(n68), .Y(SUM[16]) );
  NAND3X4 U146 ( .A(n116), .B(n77), .C(n78), .Y(n111) );
  OR2X4 U147 ( .A(A[11]), .B(B[11]), .Y(n90) );
  OR2X4 U148 ( .A(A[10]), .B(B[10]), .Y(n89) );
  OR2X4 U149 ( .A(B[9]), .B(A[9]), .Y(n88) );
  OR2X4 U150 ( .A(A[6]), .B(B[6]), .Y(n42) );
endmodule


module butterfly_DW01_sub_70 ( A, B, DIFF );
  input [16:0] A;
  input [16:0] B;
  output [16:0] DIFF;
  wire   n147, n1, n2, n3, n4, n5, n6, n7, n8, n9, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146;

  NAND2X1 U3 ( .A(n1), .B(B[15]), .Y(n79) );
  CLKINVX20 U4 ( .A(A[15]), .Y(n1) );
  INVX4 U5 ( .A(n11), .Y(n85) );
  NOR2X4 U6 ( .A(n112), .B(n14), .Y(n116) );
  CLKINVX2 U7 ( .A(n80), .Y(n2) );
  NAND2X2 U8 ( .A(n74), .B(n11), .Y(n123) );
  NAND2X2 U9 ( .A(n3), .B(B[14]), .Y(n83) );
  CLKINVX20 U10 ( .A(A[14]), .Y(n3) );
  XOR2X4 U11 ( .A(n4), .B(n115), .Y(DIFF[14]) );
  NAND2X2 U12 ( .A(n83), .B(n78), .Y(n4) );
  OR2X2 U13 ( .A(B[15]), .B(n13), .Y(n72) );
  XOR2X4 U14 ( .A(n5), .B(n6), .Y(DIFF[16]) );
  NAND3X4 U15 ( .A(n67), .B(n66), .C(n68), .Y(n5) );
  XNOR2X4 U16 ( .A(B[16]), .B(A[16]), .Y(n6) );
  NOR2X4 U17 ( .A(n20), .B(n21), .Y(n19) );
  INVX4 U18 ( .A(n22), .Y(n20) );
  NAND2X4 U19 ( .A(n119), .B(n99), .Y(n95) );
  INVXL U20 ( .A(n99), .Y(n8) );
  OR2X4 U21 ( .A(B[13]), .B(n7), .Y(n110) );
  CLKINVX20 U22 ( .A(A[13]), .Y(n7) );
  NAND2X1 U23 ( .A(n110), .B(n74), .Y(n109) );
  OAI21X4 U24 ( .A0(n104), .A1(n105), .B0(n9), .Y(n103) );
  AOI2BB1X4 U25 ( .A0N(n114), .A1N(n8), .B0(n124), .Y(n122) );
  NOR2BX4 U26 ( .AN(n30), .B(n31), .Y(n29) );
  NAND2BX2 U27 ( .AN(B[7]), .B(A[7]), .Y(n30) );
  BUFX4 U28 ( .A(n78), .Y(n9) );
  AOI21X2 U29 ( .A0(n107), .A1(n108), .B0(n109), .Y(n104) );
  INVX3 U30 ( .A(n99), .Y(n112) );
  NOR2BX2 U31 ( .AN(n79), .B(n80), .Y(n69) );
  INVX1 U32 ( .A(A[15]), .Y(n13) );
  NAND2BX1 U33 ( .AN(n15), .B(A[1]), .Y(n60) );
  BUFX4 U34 ( .A(n147), .Y(DIFF[8]) );
  XOR2X2 U35 ( .A(n52), .B(n56), .Y(DIFF[2]) );
  OAI21X2 U36 ( .A0(n58), .A1(n59), .B0(n60), .Y(n52) );
  INVX4 U37 ( .A(n140), .Y(n59) );
  XOR2X4 U38 ( .A(n132), .B(n130), .Y(DIFF[10]) );
  NOR2X4 U39 ( .A(n25), .B(n26), .Y(n24) );
  BUFX8 U40 ( .A(n120), .Y(n11) );
  NAND2BX1 U41 ( .AN(A[3]), .B(B[3]), .Y(n54) );
  INVX4 U42 ( .A(n18), .Y(n134) );
  INVX8 U43 ( .A(n126), .Y(n131) );
  AND2X1 U44 ( .A(n96), .B(n95), .Y(n94) );
  NAND3XL U45 ( .A(n96), .B(n113), .C(n114), .Y(n117) );
  OAI21X2 U46 ( .A0(n73), .A1(n74), .B0(n75), .Y(n70) );
  NAND2X2 U47 ( .A(n22), .B(n27), .Y(n127) );
  NAND3X4 U48 ( .A(n127), .B(n97), .C(n98), .Y(n125) );
  NAND2X4 U49 ( .A(n99), .B(n96), .Y(n128) );
  NAND2BX4 U50 ( .AN(A[9]), .B(B[9]), .Y(n97) );
  AND2X2 U51 ( .A(B[15]), .B(n13), .Y(n90) );
  OR2X4 U52 ( .A(n111), .B(B[12]), .Y(n74) );
  NOR2X4 U53 ( .A(n133), .B(n131), .Y(n132) );
  INVX2 U54 ( .A(n98), .Y(n133) );
  INVX8 U55 ( .A(n82), .Y(n73) );
  XOR2X4 U56 ( .A(n18), .B(n19), .Y(DIFF[9]) );
  XNOR2X4 U57 ( .A(n121), .B(n12), .Y(DIFF[13]) );
  OR2X4 U58 ( .A(n76), .B(n73), .Y(n12) );
  NAND4BX1 U59 ( .AN(n81), .B(n82), .C(n84), .D(n2), .Y(n67) );
  INVX8 U60 ( .A(n97), .Y(n21) );
  NAND2X2 U61 ( .A(n82), .B(n11), .Y(n14) );
  INVX4 U62 ( .A(n78), .Y(n77) );
  NAND4BX1 U63 ( .AN(n40), .B(n48), .C(n33), .D(n32), .Y(n145) );
  NAND2BX4 U64 ( .AN(A[6]), .B(B[6]), .Y(n33) );
  INVX4 U65 ( .A(n139), .Y(n40) );
  NAND2BX4 U66 ( .AN(A[5]), .B(B[5]), .Y(n139) );
  OR2X4 U67 ( .A(B[14]), .B(n106), .Y(n78) );
  NAND3XL U68 ( .A(n114), .B(n113), .C(n96), .Y(n107) );
  CLKINVX4 U69 ( .A(n119), .Y(n113) );
  NAND4BX2 U70 ( .AN(n26), .B(n23), .C(n97), .D(n98), .Y(n114) );
  NAND4BX1 U71 ( .AN(n26), .B(n97), .C(n98), .D(n99), .Y(n86) );
  NAND2X4 U72 ( .A(n125), .B(n126), .Y(n119) );
  NOR2X4 U73 ( .A(n85), .B(n90), .Y(n84) );
  INVX8 U74 ( .A(n110), .Y(n76) );
  AOI21XL U75 ( .A0(B[12]), .A1(n111), .B0(n112), .Y(n108) );
  NAND2BX4 U76 ( .AN(B[5]), .B(A[5]), .Y(n41) );
  NAND2BX4 U77 ( .AN(A[11]), .B(B[11]), .Y(n99) );
  AOI21X4 U78 ( .A0(n69), .A1(n70), .B0(n71), .Y(n68) );
  OAI21X4 U79 ( .A0(n122), .A1(n85), .B0(n74), .Y(n121) );
  OAI21X2 U80 ( .A0(n73), .A1(n74), .B0(n110), .Y(n118) );
  NOR2X4 U81 ( .A(n76), .B(n77), .Y(n75) );
  NAND2BX1 U82 ( .AN(B[6]), .B(A[6]), .Y(n35) );
  BUFX8 U83 ( .A(B[1]), .Y(n15) );
  XOR2X4 U84 ( .A(n128), .B(n129), .Y(DIFF[11]) );
  NAND2XL U85 ( .A(n46), .B(n48), .Y(n17) );
  NAND2BX2 U86 ( .AN(A[7]), .B(B[7]), .Y(n32) );
  XOR2X4 U87 ( .A(n103), .B(n16), .Y(DIFF[15]) );
  AND2X4 U88 ( .A(n79), .B(n72), .Y(n16) );
  NAND2BX2 U89 ( .AN(A[12]), .B(B[12]), .Y(n120) );
  INVX4 U90 ( .A(n83), .Y(n80) );
  INVX3 U91 ( .A(n145), .Y(n87) );
  CLKINVX1 U92 ( .A(n32), .Y(n31) );
  OAI2BB1X2 U93 ( .A0N(n136), .A1N(n137), .B0(n32), .Y(n102) );
  NAND2BX4 U94 ( .AN(B[9]), .B(A[9]), .Y(n22) );
  AOI21X4 U95 ( .A0(n116), .A1(n117), .B0(n118), .Y(n115) );
  NAND2BX4 U96 ( .AN(A[10]), .B(B[10]), .Y(n98) );
  CLKINVX3 U97 ( .A(n23), .Y(n135) );
  OAI2BB1X4 U98 ( .A0N(n87), .A1N(n47), .B0(n102), .Y(n23) );
  NAND2X2 U99 ( .A(n41), .B(n46), .Y(n138) );
  NAND2BX4 U100 ( .AN(A[13]), .B(B[13]), .Y(n82) );
  NOR3X2 U101 ( .A(n80), .B(n85), .C(n73), .Y(n92) );
  OAI21X4 U102 ( .A0(n26), .A1(n135), .B0(n27), .Y(n18) );
  OAI21X4 U103 ( .A0(n134), .A1(n21), .B0(n22), .Y(n130) );
  NAND2BX4 U104 ( .AN(B[4]), .B(A[4]), .Y(n46) );
  NAND2BX4 U105 ( .AN(B[10]), .B(A[10]), .Y(n126) );
  XOR2X4 U106 ( .A(n123), .B(n122), .Y(DIFF[12]) );
  NAND2BX1 U107 ( .AN(A[2]), .B(B[2]), .Y(n51) );
  NAND2BX4 U108 ( .AN(B[8]), .B(A[8]), .Y(n27) );
  NAND2BX4 U109 ( .AN(B[11]), .B(A[11]), .Y(n96) );
  AOI21X2 U110 ( .A0(n98), .A1(n130), .B0(n131), .Y(n129) );
  OAI21X2 U111 ( .A0(n39), .A1(n40), .B0(n41), .Y(n34) );
  INVX1 U112 ( .A(n27), .Y(n25) );
  NAND2BX4 U113 ( .AN(n100), .B(n89), .Y(n47) );
  INVXL U114 ( .A(n89), .Y(n88) );
  INVX2 U115 ( .A(n42), .Y(n39) );
  INVX4 U116 ( .A(n35), .Y(n37) );
  NOR2X2 U117 ( .A(n53), .B(n143), .Y(n141) );
  OAI21X2 U118 ( .A0(n59), .A1(n64), .B0(n60), .Y(n143) );
  NAND2X2 U119 ( .A(n47), .B(n48), .Y(n45) );
  XOR2X1 U120 ( .A(n42), .B(n43), .Y(DIFF[5]) );
  NOR2X1 U121 ( .A(n44), .B(n40), .Y(n43) );
  NAND2X2 U122 ( .A(n96), .B(n95), .Y(n124) );
  NOR2BX2 U123 ( .AN(n30), .B(n37), .Y(n136) );
  XNOR2X1 U124 ( .A(n47), .B(n17), .Y(DIFF[4]) );
  NAND2BXL U125 ( .AN(B[3]), .B(A[3]), .Y(n55) );
  NAND2BXL U126 ( .AN(A[4]), .B(B[4]), .Y(n48) );
  NAND2BXL U127 ( .AN(A[1]), .B(n15), .Y(n140) );
  OAI21XL U128 ( .A0(n93), .A1(n86), .B0(n94), .Y(n91) );
  NAND2BXL U129 ( .AN(B[2]), .B(A[2]), .Y(n144) );
  NAND2BXL U130 ( .AN(A[0]), .B(B[0]), .Y(n65) );
  NAND2BXL U131 ( .AN(B[0]), .B(A[0]), .Y(n64) );
  NAND3BXL U132 ( .AN(n86), .B(n87), .C(n88), .Y(n81) );
  AOI21XL U133 ( .A0(n87), .A1(n100), .B0(n101), .Y(n93) );
  INVX1 U134 ( .A(n102), .Y(n101) );
  INVX1 U135 ( .A(n72), .Y(n71) );
  OAI21X2 U136 ( .A0(n141), .A1(n142), .B0(n55), .Y(n100) );
  NAND2X1 U137 ( .A(n51), .B(n54), .Y(n142) );
  XOR2X2 U138 ( .A(n34), .B(n36), .Y(DIFF[6]) );
  NOR2X2 U139 ( .A(n37), .B(n38), .Y(n36) );
  INVX1 U140 ( .A(n33), .Y(n38) );
  XOR2X1 U141 ( .A(n23), .B(n24), .Y(n147) );
  INVX1 U142 ( .A(n41), .Y(n44) );
  XOR2X2 U143 ( .A(n28), .B(n29), .Y(DIFF[7]) );
  OAI2BB1X1 U144 ( .A0N(n33), .A1N(n34), .B0(n35), .Y(n28) );
  NAND2X2 U145 ( .A(n45), .B(n46), .Y(n42) );
  NAND3X1 U146 ( .A(n33), .B(n138), .C(n139), .Y(n137) );
  INVX1 U147 ( .A(n61), .Y(n58) );
  NAND4X1 U148 ( .A(n51), .B(n140), .C(n54), .D(n65), .Y(n89) );
  NOR2XL U149 ( .A(n53), .B(n57), .Y(n56) );
  INVX1 U150 ( .A(n51), .Y(n57) );
  XOR2X1 U151 ( .A(n49), .B(n50), .Y(DIFF[3]) );
  NAND2X1 U152 ( .A(n54), .B(n55), .Y(n49) );
  AOI21XL U153 ( .A0(n51), .A1(n52), .B0(n53), .Y(n50) );
  XOR2X1 U154 ( .A(n61), .B(n62), .Y(DIFF[1]) );
  NOR2XL U155 ( .A(n63), .B(n59), .Y(n62) );
  INVX1 U156 ( .A(n60), .Y(n63) );
  NAND2BX1 U157 ( .AN(n65), .B(n64), .Y(n61) );
  NAND2X1 U158 ( .A(n65), .B(n64), .Y(DIFF[0]) );
  OAI2BB1X1 U159 ( .A0N(n106), .A1N(B[14]), .B0(n82), .Y(n105) );
  INVX1 U160 ( .A(A[14]), .Y(n106) );
  NAND3BX1 U161 ( .AN(n90), .B(n91), .C(n92), .Y(n66) );
  NAND2BXL U162 ( .AN(A[8]), .B(B[8]), .Y(n146) );
  INVX1 U163 ( .A(A[12]), .Y(n111) );
  CLKINVX3 U164 ( .A(n144), .Y(n53) );
  CLKINVX3 U165 ( .A(n146), .Y(n26) );
endmodule


module butterfly_DW01_add_91 ( A, B, SUM );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139;

  NAND2X2 U2 ( .A(n90), .B(n104), .Y(n124) );
  CLKBUFX4 U3 ( .A(A[12]), .Y(n1) );
  INVX3 U4 ( .A(n70), .Y(n69) );
  NAND2X2 U5 ( .A(B[15]), .B(A[15]), .Y(n70) );
  NOR2X4 U6 ( .A(n101), .B(n120), .Y(n97) );
  NAND2X4 U7 ( .A(n4), .B(n87), .Y(n95) );
  AOI21X4 U8 ( .A0(n67), .A1(n68), .B0(n69), .Y(n66) );
  NOR2X4 U9 ( .A(n74), .B(n75), .Y(n67) );
  NAND2X2 U10 ( .A(B[12]), .B(A[12]), .Y(n99) );
  NAND2X2 U11 ( .A(B[11]), .B(A[11]), .Y(n104) );
  XOR2X4 U12 ( .A(n28), .B(n29), .Y(SUM[8]) );
  NOR2BX4 U13 ( .AN(n30), .B(n31), .Y(n29) );
  XOR2X4 U14 ( .A(n24), .B(n25), .Y(SUM[9]) );
  XOR2X4 U15 ( .A(n126), .B(n128), .Y(SUM[10]) );
  INVX2 U16 ( .A(n124), .Y(n14) );
  NOR2BX2 U17 ( .AN(n34), .B(n35), .Y(n33) );
  INVX4 U18 ( .A(n90), .Y(n101) );
  NAND4BX1 U19 ( .AN(n31), .B(n88), .C(n5), .D(n90), .Y(n79) );
  BUFX4 U20 ( .A(n118), .Y(n2) );
  NAND2X4 U21 ( .A(B[9]), .B(A[9]), .Y(n26) );
  NOR2BX4 U22 ( .AN(n104), .B(n81), .Y(n80) );
  NOR3X4 U23 ( .A(n81), .B(n112), .C(n113), .Y(n108) );
  INVX4 U24 ( .A(n115), .Y(n81) );
  OAI21X1 U25 ( .A0(n78), .A1(n79), .B0(n80), .Y(n77) );
  NAND2X4 U26 ( .A(B[13]), .B(A[13]), .Y(n100) );
  NAND2XL U27 ( .A(n99), .B(n100), .Y(n98) );
  AOI21X2 U28 ( .A0(n96), .A1(n97), .B0(n98), .Y(n94) );
  NAND2X2 U29 ( .A(n6), .B(n73), .Y(n109) );
  INVX4 U30 ( .A(n20), .Y(n9) );
  INVX1 U31 ( .A(n87), .Y(n75) );
  NOR2BX2 U32 ( .AN(n39), .B(n38), .Y(n41) );
  INVX4 U33 ( .A(n134), .Y(n38) );
  XOR2X2 U34 ( .A(n40), .B(n41), .Y(SUM[6]) );
  NAND2X1 U35 ( .A(B[6]), .B(A[6]), .Y(n39) );
  NAND2X2 U36 ( .A(B[5]), .B(A[5]), .Y(n43) );
  NAND2X2 U37 ( .A(B[4]), .B(A[4]), .Y(n47) );
  NAND2X2 U38 ( .A(B[14]), .B(A[14]), .Y(n72) );
  NAND2X2 U39 ( .A(n70), .B(n76), .Y(n93) );
  NAND3X2 U40 ( .A(n71), .B(n72), .C(n100), .Y(n68) );
  AND2X4 U41 ( .A(n72), .B(n87), .Y(n107) );
  INVX1 U42 ( .A(n105), .Y(n103) );
  NAND2X4 U43 ( .A(n3), .B(n77), .Y(n65) );
  AND4X2 U44 ( .A(n4), .B(n76), .C(n87), .D(n6), .Y(n3) );
  BUFX8 U45 ( .A(n73), .Y(n4) );
  CLKINVX3 U46 ( .A(n129), .Y(n5) );
  INVX2 U47 ( .A(n89), .Y(n129) );
  NAND2X2 U48 ( .A(B[10]), .B(A[10]), .Y(n122) );
  NAND2X2 U49 ( .A(n118), .B(n19), .Y(n117) );
  OAI21X4 U50 ( .A0(n94), .A1(n95), .B0(n72), .Y(n92) );
  INVX4 U51 ( .A(n91), .Y(n31) );
  CLKINVX8 U52 ( .A(n120), .Y(n6) );
  INVX8 U53 ( .A(n19), .Y(n120) );
  XOR2X4 U54 ( .A(n7), .B(n8), .Y(SUM[16]) );
  NAND2X4 U55 ( .A(n65), .B(n66), .Y(n7) );
  XOR2X4 U56 ( .A(A[16]), .B(B[16]), .Y(n8) );
  AOI21X2 U57 ( .A0(n89), .A1(n126), .B0(n127), .Y(n125) );
  OAI21X4 U58 ( .A0(n130), .A1(n27), .B0(n26), .Y(n126) );
  INVX2 U59 ( .A(n122), .Y(n127) );
  INVX2 U60 ( .A(n104), .Y(n112) );
  NAND2X4 U61 ( .A(n9), .B(n116), .Y(n12) );
  NAND2X4 U62 ( .A(n100), .B(n73), .Y(n116) );
  CLKINVX3 U63 ( .A(n76), .Y(n74) );
  NAND3XL U64 ( .A(n102), .B(n103), .C(n104), .Y(n96) );
  NAND2X4 U65 ( .A(n121), .B(n122), .Y(n105) );
  NAND2BX4 U66 ( .AN(n102), .B(n90), .Y(n114) );
  OR2X4 U67 ( .A(A[11]), .B(B[11]), .Y(n90) );
  INVX4 U68 ( .A(n114), .Y(n113) );
  NAND2X4 U69 ( .A(n105), .B(n90), .Y(n115) );
  INVX2 U70 ( .A(n100), .Y(n111) );
  INVX4 U71 ( .A(n116), .Y(n10) );
  NOR2BX4 U72 ( .AN(n26), .B(n27), .Y(n25) );
  INVX4 U73 ( .A(n88), .Y(n27) );
  NAND3X4 U74 ( .A(n114), .B(n104), .C(n115), .Y(n118) );
  NAND4X2 U75 ( .A(n28), .B(n89), .C(n91), .D(n88), .Y(n102) );
  OR2X4 U76 ( .A(A[12]), .B(B[12]), .Y(n19) );
  NAND2X2 U77 ( .A(n20), .B(n10), .Y(n11) );
  NAND3X2 U78 ( .A(n88), .B(n123), .C(n89), .Y(n121) );
  NAND2XL U79 ( .A(n26), .B(n30), .Y(n123) );
  OR2X4 U80 ( .A(A[13]), .B(B[13]), .Y(n73) );
  OAI21X4 U81 ( .A0(n23), .A1(n46), .B0(n47), .Y(n44) );
  INVX4 U82 ( .A(n83), .Y(n46) );
  NOR2X4 U83 ( .A(A[4]), .B(B[4]), .Y(n23) );
  AOI21X2 U84 ( .A0(n73), .A1(n21), .B0(n111), .Y(n110) );
  OAI21X4 U85 ( .A0(n46), .A1(n86), .B0(n85), .Y(n28) );
  OAI21X4 U86 ( .A0(n132), .A1(n133), .B0(n36), .Y(n85) );
  AOI211X2 U87 ( .A0(n43), .A1(n47), .B0(n38), .C0(n22), .Y(n132) );
  NAND2X2 U88 ( .A(n131), .B(n30), .Y(n24) );
  NAND2X4 U89 ( .A(B[8]), .B(A[8]), .Y(n30) );
  XOR2X4 U90 ( .A(n2), .B(n119), .Y(SUM[12]) );
  NOR2BX4 U91 ( .AN(n99), .B(n120), .Y(n119) );
  OR2X4 U92 ( .A(A[2]), .B(B[2]), .Y(n58) );
  XOR2X2 U93 ( .A(n32), .B(n33), .Y(SUM[7]) );
  OAI21X1 U94 ( .A0(n37), .A1(n38), .B0(n39), .Y(n32) );
  OR2X2 U95 ( .A(A[8]), .B(B[8]), .Y(n91) );
  OR2X4 U96 ( .A(A[14]), .B(B[14]), .Y(n87) );
  OR2X4 U97 ( .A(A[9]), .B(B[9]), .Y(n88) );
  NOR2BX2 U98 ( .AN(n122), .B(n129), .Y(n128) );
  NAND2X4 U99 ( .A(n11), .B(n12), .Y(SUM[13]) );
  AND2X4 U100 ( .A(n99), .B(n117), .Y(n20) );
  OR2X4 U101 ( .A(n108), .B(n109), .Y(n13) );
  NAND2X4 U102 ( .A(n13), .B(n110), .Y(n106) );
  XOR2X4 U103 ( .A(n106), .B(n107), .Y(SUM[14]) );
  NAND2X2 U104 ( .A(n124), .B(n15), .Y(n16) );
  NAND2X2 U105 ( .A(n14), .B(n125), .Y(n17) );
  NAND2X4 U106 ( .A(n16), .B(n17), .Y(SUM[11]) );
  INVX2 U107 ( .A(n125), .Y(n15) );
  XNOR2X4 U108 ( .A(n93), .B(n92), .Y(SUM[15]) );
  OAI21X4 U109 ( .A0(n42), .A1(n22), .B0(n43), .Y(n40) );
  NAND4BBX2 U110 ( .AN(n22), .BN(n23), .C(n134), .D(n36), .Y(n86) );
  NOR2BX4 U111 ( .AN(n43), .B(n22), .Y(n45) );
  NOR2X4 U112 ( .A(A[5]), .B(B[5]), .Y(n22) );
  CLKINVX3 U113 ( .A(n24), .Y(n130) );
  OAI21X4 U114 ( .A0(n136), .A1(n137), .B0(n51), .Y(n83) );
  NAND2X1 U115 ( .A(B[1]), .B(A[1]), .Y(n61) );
  NAND2X2 U116 ( .A(B[2]), .B(A[2]), .Y(n55) );
  NAND2X2 U117 ( .A(n28), .B(n91), .Y(n131) );
  OR2X4 U118 ( .A(A[7]), .B(B[7]), .Y(n36) );
  NAND2X4 U119 ( .A(B[0]), .B(A[0]), .Y(n64) );
  NOR2BX2 U120 ( .AN(n55), .B(n54), .Y(n57) );
  OR2X4 U121 ( .A(A[3]), .B(B[3]), .Y(n135) );
  OR2X4 U122 ( .A(A[1]), .B(B[1]), .Y(n59) );
  NOR2BX1 U123 ( .AN(n64), .B(n18), .Y(SUM[0]) );
  NOR2XL U124 ( .A(A[0]), .B(B[0]), .Y(n18) );
  NAND2X2 U125 ( .A(n34), .B(n39), .Y(n133) );
  NOR2X2 U126 ( .A(n138), .B(n139), .Y(n136) );
  OAI21X2 U127 ( .A0(n63), .A1(n64), .B0(n61), .Y(n139) );
  INVX2 U128 ( .A(n40), .Y(n37) );
  OAI2BB1X2 U129 ( .A0N(n59), .A1N(n60), .B0(n61), .Y(n56) );
  OR2X2 U130 ( .A(A[6]), .B(B[6]), .Y(n134) );
  OR2X4 U131 ( .A(A[15]), .B(B[15]), .Y(n76) );
  INVX1 U132 ( .A(n64), .Y(n60) );
  INVX1 U133 ( .A(n86), .Y(n82) );
  INVX1 U134 ( .A(n85), .Y(n84) );
  INVX1 U135 ( .A(n56), .Y(n53) );
  INVX1 U136 ( .A(n44), .Y(n42) );
  NAND2X1 U137 ( .A(n58), .B(n135), .Y(n137) );
  XOR2X1 U138 ( .A(n44), .B(n45), .Y(SUM[5]) );
  AOI21XL U139 ( .A0(n82), .A1(n83), .B0(n84), .Y(n78) );
  INVX1 U140 ( .A(n36), .Y(n35) );
  INVX1 U141 ( .A(n59), .Y(n63) );
  INVX1 U142 ( .A(n58), .Y(n54) );
  XOR2X1 U143 ( .A(n83), .B(n48), .Y(SUM[4]) );
  NOR2BX1 U144 ( .AN(n47), .B(n23), .Y(n48) );
  XOR2X1 U145 ( .A(n56), .B(n57), .Y(SUM[2]) );
  INVX1 U146 ( .A(n55), .Y(n138) );
  XOR2X1 U147 ( .A(n49), .B(n50), .Y(SUM[3]) );
  NOR2BX1 U148 ( .AN(n51), .B(n52), .Y(n50) );
  OAI21XL U149 ( .A0(n53), .A1(n54), .B0(n55), .Y(n49) );
  INVX1 U150 ( .A(n135), .Y(n52) );
  XOR2X1 U151 ( .A(n60), .B(n62), .Y(SUM[1]) );
  NOR2BXL U152 ( .AN(n61), .B(n63), .Y(n62) );
  AND2X1 U153 ( .A(n1), .B(B[12]), .Y(n21) );
  NAND2XL U154 ( .A(B[7]), .B(A[7]), .Y(n34) );
  NAND2XL U155 ( .A(B[3]), .B(A[3]), .Y(n51) );
  NAND3XL U156 ( .A(n1), .B(B[12]), .C(n73), .Y(n71) );
  OR2X4 U157 ( .A(A[10]), .B(B[10]), .Y(n89) );
endmodule


module butterfly_DW01_add_98 ( A, B, SUM );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126;

  DLY1X1 U2 ( .A(B[14]), .Y(n14) );
  AND2X4 U3 ( .A(B[15]), .B(A[15]), .Y(n1) );
  CLKBUFX4 U4 ( .A(n86), .Y(n12) );
  AND3X4 U5 ( .A(n78), .B(n110), .C(n77), .Y(n2) );
  NAND2X4 U6 ( .A(n3), .B(n71), .Y(n70) );
  AND4X2 U7 ( .A(n84), .B(n85), .C(n12), .D(n13), .Y(n3) );
  NAND2BX4 U8 ( .AN(n1), .B(n85), .Y(n9) );
  NAND2X2 U9 ( .A(B[10]), .B(A[10]), .Y(n112) );
  INVX8 U10 ( .A(n11), .Y(n24) );
  AND2X4 U11 ( .A(A[14]), .B(B[14]), .Y(n11) );
  NAND2X2 U12 ( .A(B[4]), .B(A[4]), .Y(n48) );
  NOR2BX4 U13 ( .AN(n39), .B(n38), .Y(n41) );
  INVX1 U14 ( .A(n42), .Y(n38) );
  OAI21X1 U15 ( .A0(n37), .A1(n38), .B0(n39), .Y(n33) );
  NAND3X2 U16 ( .A(n121), .B(n39), .C(n35), .Y(n120) );
  OR2X1 U17 ( .A(B[10]), .B(A[10]), .Y(n4) );
  AND2X4 U18 ( .A(n86), .B(n24), .Y(n5) );
  INVXL U19 ( .A(n29), .Y(n6) );
  NAND4BBX4 U20 ( .AN(n7), .BN(n6), .C(n89), .D(n90), .Y(n110) );
  NAND2XL U21 ( .A(n91), .B(n88), .Y(n7) );
  OAI21X1 U22 ( .A0(n65), .A1(n66), .B0(n63), .Y(n125) );
  CLKINVX2 U23 ( .A(n83), .Y(n79) );
  NOR2BX1 U24 ( .AN(n44), .B(n22), .Y(n46) );
  NOR2X2 U25 ( .A(n92), .B(n1), .Y(n69) );
  AND2X4 U26 ( .A(B[13]), .B(A[13]), .Y(n8) );
  NAND2X4 U27 ( .A(B[8]), .B(A[8]), .Y(n31) );
  OR2X4 U28 ( .A(A[8]), .B(B[8]), .Y(n91) );
  OAI21X4 U29 ( .A0(n23), .A1(n47), .B0(n48), .Y(n45) );
  NOR2BX2 U30 ( .AN(n48), .B(n23), .Y(n49) );
  NOR2X2 U31 ( .A(A[4]), .B(B[4]), .Y(n23) );
  XOR2X2 U32 ( .A(n40), .B(n41), .Y(SUM[6]) );
  NAND2X2 U33 ( .A(B[9]), .B(A[9]), .Y(n27) );
  OR2X4 U34 ( .A(A[9]), .B(B[9]), .Y(n88) );
  INVX4 U35 ( .A(n80), .Y(n47) );
  XOR2X4 U36 ( .A(n117), .B(n115), .Y(SUM[10]) );
  AOI21X2 U37 ( .A0(n89), .A1(n115), .B0(n116), .Y(n114) );
  XNOR2X4 U38 ( .A(n97), .B(n9), .Y(SUM[15]) );
  NAND2X4 U39 ( .A(n17), .B(n96), .Y(n101) );
  AOI21X4 U40 ( .A0(n13), .A1(n10), .B0(n101), .Y(n98) );
  NAND2X4 U41 ( .A(n10), .B(n18), .Y(n19) );
  INVX4 U42 ( .A(n2), .Y(n10) );
  OAI21X4 U43 ( .A0(n103), .A1(n104), .B0(n17), .Y(n102) );
  AOI21X2 U44 ( .A0(A[14]), .A1(n14), .B0(n95), .Y(n93) );
  NAND2X2 U45 ( .A(n12), .B(n85), .Y(n94) );
  NOR2BX2 U46 ( .AN(n84), .B(n96), .Y(n95) );
  NAND2X4 U47 ( .A(n84), .B(n17), .Y(n106) );
  NAND2X4 U48 ( .A(B[12]), .B(A[12]), .Y(n96) );
  XOR2X4 U49 ( .A(n102), .B(n5), .Y(SUM[14]) );
  XOR2X4 U50 ( .A(n25), .B(n26), .Y(SUM[9]) );
  NAND2X2 U51 ( .A(n90), .B(n77), .Y(n113) );
  CLKINVX8 U52 ( .A(n87), .Y(n109) );
  OR2X4 U53 ( .A(A[12]), .B(B[12]), .Y(n87) );
  NAND2X2 U54 ( .A(n84), .B(n86), .Y(n99) );
  NAND2X2 U55 ( .A(B[7]), .B(A[7]), .Y(n35) );
  NAND2X4 U56 ( .A(n69), .B(n70), .Y(n67) );
  NAND2X2 U57 ( .A(B[11]), .B(A[11]), .Y(n77) );
  AOI21X2 U58 ( .A0(n93), .A1(n17), .B0(n94), .Y(n92) );
  NAND2X2 U59 ( .A(n87), .B(n84), .Y(n104) );
  INVX4 U60 ( .A(n89), .Y(n118) );
  OR2X4 U61 ( .A(B[10]), .B(A[10]), .Y(n89) );
  NAND4BBX2 U62 ( .AN(n22), .BN(n23), .C(n42), .D(n123), .Y(n83) );
  OAI2BB1X4 U63 ( .A0N(n91), .A1N(n29), .B0(n31), .Y(n25) );
  XOR2X2 U64 ( .A(n29), .B(n30), .Y(SUM[8]) );
  INVX4 U65 ( .A(n109), .Y(n13) );
  NOR2X4 U66 ( .A(A[5]), .B(B[5]), .Y(n22) );
  OR2X4 U67 ( .A(A[7]), .B(B[7]), .Y(n123) );
  NAND2BX4 U68 ( .AN(n36), .B(n120), .Y(n82) );
  INVX2 U69 ( .A(n108), .Y(n18) );
  NAND2X2 U70 ( .A(n2), .B(n108), .Y(n20) );
  NOR2BX4 U71 ( .AN(n96), .B(n109), .Y(n108) );
  NAND2X4 U72 ( .A(n15), .B(n24), .Y(n97) );
  NOR2X1 U73 ( .A(n105), .B(n100), .Y(n103) );
  INVX4 U74 ( .A(n91), .Y(n32) );
  AND2X4 U75 ( .A(n100), .B(n87), .Y(n16) );
  OAI21X4 U76 ( .A0(n43), .A1(n22), .B0(n44), .Y(n40) );
  NAND2X1 U77 ( .A(n44), .B(n48), .Y(n122) );
  NAND2X4 U78 ( .A(B[5]), .B(A[5]), .Y(n44) );
  XOR2X2 U79 ( .A(B[16]), .B(A[16]), .Y(n68) );
  OAI211X2 U80 ( .A0(n28), .A1(n31), .B0(n27), .C0(n112), .Y(n111) );
  NAND3X4 U81 ( .A(n90), .B(n4), .C(n111), .Y(n78) );
  OR2X4 U82 ( .A(B[13]), .B(A[13]), .Y(n84) );
  INVX2 U83 ( .A(n45), .Y(n43) );
  NOR2BX2 U84 ( .AN(n27), .B(n28), .Y(n26) );
  NOR2BX4 U85 ( .AN(n112), .B(n118), .Y(n117) );
  XOR2X4 U86 ( .A(n113), .B(n114), .Y(SUM[11]) );
  INVX4 U87 ( .A(n88), .Y(n28) );
  OR2X4 U88 ( .A(A[14]), .B(B[14]), .Y(n86) );
  INVX4 U89 ( .A(n96), .Y(n105) );
  OR2X4 U90 ( .A(n99), .B(n98), .Y(n15) );
  NOR2X4 U91 ( .A(n16), .B(n105), .Y(n107) );
  XOR2X4 U92 ( .A(n107), .B(n106), .Y(SUM[13]) );
  OR2X4 U93 ( .A(B[15]), .B(A[15]), .Y(n85) );
  NAND2X4 U94 ( .A(n19), .B(n20), .Y(SUM[12]) );
  XOR2X4 U95 ( .A(n67), .B(n68), .Y(SUM[16]) );
  INVX8 U96 ( .A(n8), .Y(n17) );
  NAND3X4 U97 ( .A(n78), .B(n110), .C(n77), .Y(n100) );
  OR2X2 U98 ( .A(A[1]), .B(B[1]), .Y(n61) );
  NAND3BX1 U99 ( .AN(n22), .B(n122), .C(n42), .Y(n121) );
  NOR2BXL U100 ( .AN(n63), .B(n65), .Y(n64) );
  NAND2XL U101 ( .A(B[1]), .B(A[1]), .Y(n63) );
  OAI21X4 U102 ( .A0(n47), .A1(n83), .B0(n82), .Y(n29) );
  INVXL U103 ( .A(n112), .Y(n116) );
  INVXL U104 ( .A(n78), .Y(n75) );
  OAI21X4 U105 ( .A0(n119), .A1(n28), .B0(n27), .Y(n115) );
  INVX4 U106 ( .A(n25), .Y(n119) );
  XOR2X2 U107 ( .A(n33), .B(n34), .Y(SUM[7]) );
  INVX2 U108 ( .A(n40), .Y(n37) );
  INVXL U109 ( .A(n77), .Y(n76) );
  INVXL U110 ( .A(n60), .Y(n56) );
  INVXL U111 ( .A(n54), .Y(n53) );
  CLKINVX3 U112 ( .A(n57), .Y(n126) );
  INVXL U113 ( .A(n66), .Y(n62) );
  NOR2BX1 U114 ( .AN(n66), .B(n21), .Y(SUM[0]) );
  NOR2XL U115 ( .A(A[0]), .B(B[0]), .Y(n21) );
  INVX1 U116 ( .A(n82), .Y(n81) );
  NOR2BX1 U117 ( .AN(n31), .B(n32), .Y(n30) );
  XOR2X1 U118 ( .A(n45), .B(n46), .Y(SUM[5]) );
  NOR2BX1 U119 ( .AN(n35), .B(n36), .Y(n34) );
  OAI21XL U120 ( .A0(n72), .A1(n73), .B0(n74), .Y(n71) );
  AOI21X1 U121 ( .A0(n79), .A1(n80), .B0(n81), .Y(n72) );
  NAND4BXL U122 ( .AN(n32), .B(n88), .C(n89), .D(n90), .Y(n73) );
  NOR2X1 U123 ( .A(n75), .B(n76), .Y(n74) );
  INVX1 U124 ( .A(n123), .Y(n36) );
  INVX1 U125 ( .A(n61), .Y(n65) );
  XOR2X1 U126 ( .A(n80), .B(n49), .Y(SUM[4]) );
  XOR2X1 U127 ( .A(n62), .B(n64), .Y(SUM[1]) );
  XOR2X1 U128 ( .A(n58), .B(n59), .Y(SUM[2]) );
  NOR2BX1 U129 ( .AN(n57), .B(n56), .Y(n59) );
  XOR2X1 U130 ( .A(n50), .B(n51), .Y(SUM[3]) );
  OAI21XL U131 ( .A0(n55), .A1(n56), .B0(n57), .Y(n50) );
  NOR2BX1 U132 ( .AN(n52), .B(n53), .Y(n51) );
  INVX1 U133 ( .A(n58), .Y(n55) );
  OAI2BB1X1 U134 ( .A0N(n61), .A1N(n62), .B0(n63), .Y(n58) );
  NAND2XL U135 ( .A(B[6]), .B(A[6]), .Y(n39) );
  OR2X2 U136 ( .A(A[6]), .B(B[6]), .Y(n42) );
  NAND2X2 U137 ( .A(n52), .B(n124), .Y(n80) );
  OAI211X1 U138 ( .A0(n125), .A1(n126), .B0(n60), .C0(n54), .Y(n124) );
  OR2X2 U139 ( .A(A[3]), .B(B[3]), .Y(n54) );
  NAND2X1 U140 ( .A(B[2]), .B(A[2]), .Y(n57) );
  NAND2X1 U141 ( .A(B[3]), .B(A[3]), .Y(n52) );
  OR2X2 U142 ( .A(A[2]), .B(B[2]), .Y(n60) );
  NAND2X2 U143 ( .A(B[0]), .B(A[0]), .Y(n66) );
  OR2X4 U144 ( .A(B[11]), .B(A[11]), .Y(n90) );
endmodule


module butterfly_DW01_sub_77 ( A, B, DIFF );
  input [16:0] A;
  input [16:0] B;
  output [16:0] DIFF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161;

  NAND3X2 U3 ( .A(n97), .B(n5), .C(n96), .Y(n83) );
  NAND2BX2 U4 ( .AN(B[11]), .B(A[11]), .Y(n135) );
  AND4X4 U5 ( .A(n108), .B(n16), .C(n124), .D(n93), .Y(n120) );
  NOR2BX4 U6 ( .AN(n85), .B(n86), .Y(n84) );
  NAND2BX4 U7 ( .AN(B[15]), .B(n1), .Y(n85) );
  CLKINVX20 U8 ( .A(n2), .Y(n1) );
  CLKINVX20 U9 ( .A(A[15]), .Y(n2) );
  AND2X2 U10 ( .A(B[14]), .B(n14), .Y(n3) );
  INVX4 U11 ( .A(n129), .Y(n110) );
  INVX3 U12 ( .A(n113), .Y(n145) );
  NAND2BX4 U13 ( .AN(B[3]), .B(A[3]), .Y(n70) );
  NAND2BX4 U14 ( .AN(A[3]), .B(B[3]), .Y(n69) );
  NAND4X4 U15 ( .A(n6), .B(n33), .C(n112), .D(n113), .Y(n124) );
  OR2X4 U16 ( .A(B[14]), .B(n14), .Y(n4) );
  INVX2 U17 ( .A(n100), .Y(n99) );
  NOR2X4 U18 ( .A(n109), .B(n110), .Y(n108) );
  INVX8 U19 ( .A(n39), .Y(n20) );
  AOI21X4 U20 ( .A0(n4), .A1(n87), .B0(n89), .Y(n86) );
  NAND3X2 U21 ( .A(n153), .B(n154), .C(n47), .Y(n152) );
  NAND2X2 U22 ( .A(n57), .B(n61), .Y(n154) );
  NAND3X2 U23 ( .A(n66), .B(n69), .C(n155), .Y(n103) );
  INVXL U24 ( .A(n41), .Y(n6) );
  INVX1 U25 ( .A(A[15]), .Y(n10) );
  CLKINVX3 U26 ( .A(n31), .Y(n21) );
  INVX2 U27 ( .A(B[16]), .Y(n24) );
  NAND2X1 U28 ( .A(n69), .B(n70), .Y(n64) );
  INVX1 U29 ( .A(A[12]), .Y(n17) );
  INVX1 U30 ( .A(A[14]), .Y(n14) );
  AND2X4 U31 ( .A(n94), .B(n95), .Y(n5) );
  OR2X4 U32 ( .A(n43), .B(n44), .Y(n32) );
  INVX4 U33 ( .A(n150), .Y(n44) );
  OAI21X1 U34 ( .A0(n74), .A1(n75), .B0(n76), .Y(n67) );
  INVX3 U35 ( .A(n157), .Y(n75) );
  INVX4 U36 ( .A(n140), .Y(n149) );
  OAI21X2 U37 ( .A0(n146), .A1(n138), .B0(n140), .Y(n143) );
  NAND2X4 U38 ( .A(n133), .B(n100), .Y(n34) );
  INVX4 U39 ( .A(n133), .Y(n132) );
  XOR2X2 U40 ( .A(n45), .B(n46), .Y(DIFF[7]) );
  NAND2BX1 U41 ( .AN(B[2]), .B(A[2]), .Y(n73) );
  NAND4BX2 U42 ( .AN(n56), .B(n63), .C(n47), .D(n50), .Y(n102) );
  XNOR2X4 U43 ( .A(n42), .B(n32), .Y(DIFF[8]) );
  OR2X4 U44 ( .A(n40), .B(n41), .Y(n31) );
  INVX8 U45 ( .A(n141), .Y(n40) );
  AND2X4 U46 ( .A(n108), .B(n124), .Y(n7) );
  NOR2X4 U47 ( .A(n7), .B(n128), .Y(n126) );
  OAI21X4 U48 ( .A0(n138), .A1(n139), .B0(n140), .Y(n137) );
  INVX4 U49 ( .A(n42), .Y(n136) );
  NAND2BX4 U50 ( .AN(B[7]), .B(A[7]), .Y(n51) );
  XOR2X4 U51 ( .A(n8), .B(n125), .Y(DIFF[14]) );
  NAND2X4 U52 ( .A(n88), .B(n9), .Y(n8) );
  NAND2X4 U53 ( .A(B[14]), .B(n14), .Y(n9) );
  OR2X4 U54 ( .A(B[14]), .B(n14), .Y(n88) );
  NAND2X4 U55 ( .A(B[15]), .B(n10), .Y(n106) );
  OR2X4 U56 ( .A(B[12]), .B(n17), .Y(n93) );
  INVX4 U57 ( .A(n147), .Y(n146) );
  CLKINVX8 U58 ( .A(n90), .Y(n98) );
  OAI2BB1X4 U59 ( .A0N(n17), .A1N(B[12]), .B0(n18), .Y(n128) );
  NOR3X4 U60 ( .A(n89), .B(n98), .C(n3), .Y(n105) );
  OR2X4 U61 ( .A(B[13]), .B(n19), .Y(n15) );
  NAND3X2 U62 ( .A(n18), .B(n91), .C(n9), .Y(n87) );
  INVX4 U63 ( .A(n135), .Y(n109) );
  CLKINVXL U64 ( .A(B[12]), .Y(n11) );
  INVX2 U65 ( .A(n11), .Y(n12) );
  XNOR2X4 U66 ( .A(n130), .B(n13), .Y(DIFF[13]) );
  AND2X4 U67 ( .A(n18), .B(n15), .Y(n13) );
  INVXL U68 ( .A(n101), .Y(n95) );
  AND2X4 U69 ( .A(n92), .B(n90), .Y(n123) );
  NAND2X4 U70 ( .A(n17), .B(B[12]), .Y(n100) );
  NAND2X4 U71 ( .A(B[14]), .B(n14), .Y(n92) );
  NAND2BX4 U72 ( .AN(n81), .B(n28), .Y(n30) );
  NAND2X4 U73 ( .A(n85), .B(n106), .Y(n119) );
  OR2X4 U74 ( .A(B[13]), .B(n19), .Y(n16) );
  INVX3 U75 ( .A(n131), .Y(n134) );
  NAND3X4 U76 ( .A(n129), .B(n135), .C(n124), .Y(n131) );
  INVXL U77 ( .A(A[13]), .Y(n19) );
  OR2X4 U78 ( .A(B[12]), .B(n17), .Y(n133) );
  NAND2BX4 U79 ( .AN(A[13]), .B(B[13]), .Y(n18) );
  INVX8 U80 ( .A(n106), .Y(n89) );
  XOR2X4 U81 ( .A(n147), .B(n148), .Y(DIFF[10]) );
  NAND2X2 U82 ( .A(n93), .B(n16), .Y(n91) );
  OAI21X4 U83 ( .A0(n98), .A1(n93), .B0(n16), .Y(n127) );
  NAND2X4 U84 ( .A(n122), .B(n123), .Y(n121) );
  XNOR2X4 U85 ( .A(n118), .B(n119), .Y(DIFF[15]) );
  NAND2BX2 U86 ( .AN(A[8]), .B(B[8]), .Y(n150) );
  OAI21X4 U87 ( .A0(n20), .A1(n41), .B0(n141), .Y(n147) );
  NAND2BX4 U88 ( .AN(A[10]), .B(B[10]), .Y(n112) );
  NAND2X4 U89 ( .A(n24), .B(A[16]), .Y(n27) );
  NAND2X1 U90 ( .A(B[16]), .B(n25), .Y(n26) );
  INVX4 U91 ( .A(n38), .Y(n28) );
  NAND3BX2 U92 ( .AN(A[12]), .B(n12), .C(n15), .Y(n122) );
  NAND3X4 U93 ( .A(n152), .B(n54), .C(n51), .Y(n151) );
  INVX4 U94 ( .A(n54), .Y(n49) );
  NAND2BX4 U95 ( .AN(B[6]), .B(A[6]), .Y(n54) );
  INVX8 U96 ( .A(n142), .Y(n43) );
  NAND2BX4 U97 ( .AN(B[8]), .B(A[8]), .Y(n142) );
  XOR2X4 U98 ( .A(n143), .B(n144), .Y(DIFF[11]) );
  NAND2BX2 U99 ( .AN(A[7]), .B(B[7]), .Y(n50) );
  CLKINVX8 U100 ( .A(n111), .Y(n41) );
  AOI21X2 U101 ( .A0(n43), .A1(n111), .B0(n40), .Y(n139) );
  NAND4BX2 U102 ( .AN(n44), .B(n111), .C(n112), .D(n113), .Y(n101) );
  NAND2BX4 U103 ( .AN(A[9]), .B(B[9]), .Y(n111) );
  NAND3X4 U104 ( .A(n82), .B(n83), .C(n84), .Y(n81) );
  NAND3X2 U105 ( .A(n104), .B(n100), .C(n105), .Y(n82) );
  NOR2X4 U106 ( .A(n149), .B(n138), .Y(n148) );
  INVX8 U107 ( .A(n112), .Y(n138) );
  NAND2BX4 U108 ( .AN(B[10]), .B(A[10]), .Y(n140) );
  NAND2BX4 U109 ( .AN(A[5]), .B(B[5]), .Y(n153) );
  OAI21X2 U110 ( .A0(n55), .A1(n56), .B0(n57), .Y(n48) );
  INVX4 U111 ( .A(n153), .Y(n56) );
  NAND2BX4 U112 ( .AN(B[5]), .B(A[5]), .Y(n57) );
  NAND2BX4 U113 ( .AN(A[11]), .B(B[11]), .Y(n113) );
  NAND2BX4 U114 ( .AN(B[9]), .B(A[9]), .Y(n141) );
  NAND2X2 U115 ( .A(n39), .B(n31), .Y(n22) );
  NAND2X4 U116 ( .A(n20), .B(n21), .Y(n23) );
  NAND2X4 U117 ( .A(n22), .B(n23), .Y(DIFF[9]) );
  NAND2X4 U118 ( .A(n26), .B(n27), .Y(n38) );
  INVX1 U119 ( .A(A[16]), .Y(n25) );
  NAND2X2 U120 ( .A(n81), .B(n38), .Y(n29) );
  NAND2X4 U121 ( .A(n30), .B(n29), .Y(DIFF[16]) );
  NOR2X2 U122 ( .A(n89), .B(n3), .Y(n97) );
  NOR2XL U123 ( .A(n136), .B(n44), .Y(n33) );
  AOI21X1 U124 ( .A0(n47), .A1(n48), .B0(n49), .Y(n46) );
  NAND2BXL U125 ( .AN(A[1]), .B(B[1]), .Y(n157) );
  NAND2X4 U126 ( .A(n50), .B(n151), .Y(n117) );
  NAND2XL U127 ( .A(n50), .B(n51), .Y(n45) );
  NAND2BXL U128 ( .AN(B[0]), .B(A[0]), .Y(n80) );
  INVXL U129 ( .A(n117), .Y(n116) );
  NAND2X2 U130 ( .A(n60), .B(n61), .Y(n58) );
  NAND2X2 U131 ( .A(n62), .B(n63), .Y(n60) );
  OAI21X1 U132 ( .A0(n107), .A1(n101), .B0(n108), .Y(n104) );
  NAND2X2 U133 ( .A(n158), .B(n70), .Y(n115) );
  NAND3X2 U134 ( .A(n66), .B(n159), .C(n69), .Y(n158) );
  NAND3X2 U135 ( .A(n160), .B(n76), .C(n73), .Y(n159) );
  NAND2X2 U136 ( .A(n161), .B(n157), .Y(n160) );
  XOR2X1 U137 ( .A(n48), .B(n52), .Y(DIFF[6]) );
  NOR2XL U138 ( .A(n49), .B(n53), .Y(n52) );
  INVX2 U139 ( .A(n47), .Y(n53) );
  XOR2X4 U140 ( .A(n134), .B(n34), .Y(DIFF[12]) );
  XOR2X1 U141 ( .A(n58), .B(n35), .Y(DIFF[5]) );
  NOR2XL U142 ( .A(n59), .B(n56), .Y(n35) );
  XNOR2X1 U143 ( .A(n62), .B(n36), .Y(DIFF[4]) );
  NAND2XL U144 ( .A(n61), .B(n63), .Y(n36) );
  XOR2X1 U145 ( .A(n77), .B(n37), .Y(DIFF[1]) );
  NOR2XL U146 ( .A(n78), .B(n75), .Y(n37) );
  INVXL U147 ( .A(n73), .Y(n68) );
  INVXL U148 ( .A(n66), .Y(n72) );
  XOR2X1 U149 ( .A(n64), .B(n65), .Y(DIFF[3]) );
  AOI21XL U150 ( .A0(n66), .A1(n67), .B0(n68), .Y(n65) );
  CLKINVX3 U151 ( .A(n156), .Y(n79) );
  NAND2XL U152 ( .A(n156), .B(n80), .Y(DIFF[0]) );
  NOR2XL U153 ( .A(n102), .B(n103), .Y(n94) );
  NOR2XL U154 ( .A(n98), .B(n99), .Y(n96) );
  NAND2BX4 U155 ( .AN(n115), .B(n103), .Y(n62) );
  AOI21XL U156 ( .A0(n114), .A1(n115), .B0(n116), .Y(n107) );
  INVX1 U157 ( .A(n58), .Y(n55) );
  INVX1 U158 ( .A(n77), .Y(n74) );
  XOR2X2 U159 ( .A(n67), .B(n71), .Y(DIFF[2]) );
  NOR2X1 U160 ( .A(n68), .B(n72), .Y(n71) );
  INVX1 U161 ( .A(n80), .Y(n161) );
  NAND2XL U162 ( .A(n79), .B(n80), .Y(n77) );
  NAND2BX1 U163 ( .AN(A[2]), .B(B[2]), .Y(n66) );
  NAND2BX2 U164 ( .AN(A[4]), .B(B[4]), .Y(n63) );
  NAND2BX1 U165 ( .AN(B[1]), .B(A[1]), .Y(n76) );
  NAND2BXL U166 ( .AN(A[0]), .B(B[0]), .Y(n156) );
  CLKINVX3 U167 ( .A(n57), .Y(n59) );
  CLKINVX3 U168 ( .A(n76), .Y(n78) );
  OAI21X4 U169 ( .A0(n120), .A1(n121), .B0(n4), .Y(n118) );
  NOR2X4 U170 ( .A(n126), .B(n127), .Y(n125) );
  AOI21X4 U171 ( .A0(n131), .A1(n100), .B0(n132), .Y(n130) );
  NAND2BX4 U172 ( .AN(A[13]), .B(B[13]), .Y(n90) );
  NAND2X4 U173 ( .A(n137), .B(n113), .Y(n129) );
  NOR2X4 U174 ( .A(n145), .B(n109), .Y(n144) );
  OAI21X4 U175 ( .A0(n136), .A1(n44), .B0(n142), .Y(n39) );
  OAI2BB1X4 U176 ( .A0N(n114), .A1N(n62), .B0(n117), .Y(n42) );
  NAND2BX4 U177 ( .AN(B[4]), .B(A[4]), .Y(n61) );
  NOR2X4 U178 ( .A(n75), .B(n79), .Y(n155) );
  CLKINVX3 U179 ( .A(n102), .Y(n114) );
  NAND2BX4 U180 ( .AN(A[6]), .B(B[6]), .Y(n47) );
endmodule


module butterfly_DW01_add_100 ( A, B, SUM );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  wire   n128, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127;

  BUFX4 U2 ( .A(n92), .Y(n1) );
  INVX1 U3 ( .A(n111), .Y(n2) );
  INVX3 U4 ( .A(n112), .Y(n111) );
  NAND4BX2 U5 ( .AN(n2), .B(n87), .C(n88), .D(n89), .Y(n74) );
  OR2X4 U6 ( .A(A[3]), .B(B[3]), .Y(n53) );
  BUFX4 U7 ( .A(B[10]), .Y(n11) );
  AND2X2 U8 ( .A(B[11]), .B(A[11]), .Y(n3) );
  INVX20 U9 ( .A(n3), .Y(n76) );
  NOR2BX4 U10 ( .AN(n117), .B(n10), .Y(n118) );
  NAND2XL U11 ( .A(B[7]), .B(A[7]), .Y(n34) );
  NOR2X4 U12 ( .A(B[11]), .B(A[11]), .Y(n112) );
  NAND3X4 U13 ( .A(n83), .B(n103), .C(n104), .Y(n102) );
  NAND2X1 U14 ( .A(n91), .B(n92), .Y(n90) );
  INVX1 U15 ( .A(A[12]), .Y(n9) );
  AND2X2 U16 ( .A(n96), .B(n84), .Y(n20) );
  INVX1 U17 ( .A(A[11]), .Y(n7) );
  INVX2 U18 ( .A(n96), .Y(n68) );
  CLKINVX4 U19 ( .A(n24), .Y(n119) );
  OR2X1 U20 ( .A(A[2]), .B(B[2]), .Y(n59) );
  NAND2X1 U21 ( .A(B[2]), .B(A[2]), .Y(n56) );
  NOR2X2 U22 ( .A(A[4]), .B(B[4]), .Y(n23) );
  OAI21X4 U23 ( .A0(n23), .A1(n124), .B0(n46), .Y(n44) );
  XOR2X2 U24 ( .A(n39), .B(n40), .Y(SUM[6]) );
  AOI21X4 U25 ( .A0(n104), .A1(n103), .B0(n107), .Y(n106) );
  INVXL U26 ( .A(B[11]), .Y(n6) );
  NAND2X4 U27 ( .A(B[12]), .B(A[12]), .Y(n95) );
  NAND2X4 U28 ( .A(n15), .B(n20), .Y(n17) );
  CLKINVX4 U29 ( .A(n19), .Y(n15) );
  NAND2X1 U30 ( .A(n96), .B(n84), .Y(n4) );
  AND2X4 U31 ( .A(n77), .B(n76), .Y(n75) );
  NAND2X2 U32 ( .A(n19), .B(n4), .Y(n16) );
  OR2X4 U33 ( .A(A[15]), .B(B[15]), .Y(n84) );
  XNOR2X4 U34 ( .A(n5), .B(n104), .Y(SUM[12]) );
  NAND2X4 U35 ( .A(n95), .B(n86), .Y(n5) );
  OAI2BB1X4 U36 ( .A0N(n6), .A1N(n7), .B0(n76), .Y(n114) );
  NAND3BX2 U37 ( .AN(n9), .B(n8), .C(B[12]), .Y(n101) );
  NAND2X1 U38 ( .A(n94), .B(n95), .Y(n93) );
  NAND2X2 U39 ( .A(B[14]), .B(A[14]), .Y(n92) );
  NAND2XL U40 ( .A(n84), .B(n90), .Y(n69) );
  OR2X4 U41 ( .A(A[13]), .B(B[13]), .Y(n8) );
  NAND4XL U42 ( .A(n8), .B(n84), .C(n85), .D(n86), .Y(n71) );
  AOI21X4 U43 ( .A0(n87), .A1(n116), .B0(n109), .Y(n115) );
  OAI21X4 U44 ( .A0(n119), .A1(n27), .B0(n26), .Y(n116) );
  NAND2X4 U45 ( .A(B[6]), .B(A[6]), .Y(n38) );
  OR2X4 U46 ( .A(A[12]), .B(B[12]), .Y(n86) );
  XOR2X4 U47 ( .A(n116), .B(n118), .Y(SUM[10]) );
  NAND2X2 U48 ( .A(n24), .B(n12), .Y(n13) );
  NAND2X2 U49 ( .A(B[9]), .B(A[9]), .Y(n26) );
  OAI2BB1X4 U50 ( .A0N(n89), .A1N(n28), .B0(n30), .Y(n24) );
  NAND2X4 U51 ( .A(B[8]), .B(A[8]), .Y(n30) );
  NAND3BX4 U52 ( .AN(n68), .B(n70), .C(n69), .Y(n66) );
  NAND2BX4 U53 ( .AN(n71), .B(n72), .Y(n70) );
  OR2X4 U54 ( .A(B[12]), .B(A[12]), .Y(n103) );
  XOR2X4 U55 ( .A(B[16]), .B(A[16]), .Y(n67) );
  NOR2X2 U56 ( .A(A[5]), .B(B[5]), .Y(n22) );
  NAND2X2 U57 ( .A(n83), .B(n94), .Y(n105) );
  NAND3X1 U58 ( .A(n85), .B(n93), .C(n83), .Y(n91) );
  NAND2X4 U59 ( .A(n85), .B(n98), .Y(n97) );
  XOR2X4 U60 ( .A(n114), .B(n115), .Y(SUM[11]) );
  NAND2X2 U61 ( .A(B[4]), .B(A[4]), .Y(n46) );
  NAND2X2 U62 ( .A(n43), .B(n46), .Y(n122) );
  NOR2X4 U63 ( .A(B[10]), .B(A[10]), .Y(n10) );
  INVX2 U64 ( .A(n39), .Y(n36) );
  OAI21X2 U65 ( .A0(n42), .A1(n22), .B0(n43), .Y(n39) );
  NOR2BX4 U66 ( .AN(n26), .B(n27), .Y(n25) );
  INVX8 U67 ( .A(n88), .Y(n27) );
  INVX2 U68 ( .A(n95), .Y(n107) );
  XNOR2X4 U69 ( .A(n98), .B(n99), .Y(SUM[14]) );
  NAND2X4 U70 ( .A(n92), .B(n85), .Y(n99) );
  NAND2X4 U71 ( .A(n97), .B(n1), .Y(n19) );
  XOR2X4 U72 ( .A(n66), .B(n67), .Y(SUM[16]) );
  NAND2X2 U73 ( .A(B[15]), .B(A[15]), .Y(n96) );
  INVX8 U74 ( .A(n117), .Y(n109) );
  NAND2X4 U75 ( .A(n11), .B(A[10]), .Y(n117) );
  NAND4BBX2 U76 ( .AN(n22), .BN(n23), .C(n41), .D(n123), .Y(n82) );
  INVX4 U77 ( .A(n41), .Y(n37) );
  NAND3BX2 U78 ( .AN(n22), .B(n122), .C(n41), .Y(n121) );
  OR2X4 U79 ( .A(A[6]), .B(B[6]), .Y(n41) );
  INVX2 U80 ( .A(n44), .Y(n42) );
  OR2X4 U81 ( .A(A[7]), .B(B[7]), .Y(n123) );
  NOR2BX2 U82 ( .AN(n30), .B(n31), .Y(n29) );
  INVX4 U83 ( .A(n89), .Y(n31) );
  OR2X4 U84 ( .A(A[8]), .B(B[8]), .Y(n89) );
  NAND4BX2 U85 ( .AN(n112), .B(n28), .C(n87), .D(n113), .Y(n108) );
  NOR2X2 U86 ( .A(n27), .B(n31), .Y(n113) );
  NAND2X2 U87 ( .A(B[13]), .B(A[13]), .Y(n94) );
  NAND2X2 U88 ( .A(n119), .B(n25), .Y(n14) );
  NAND2X4 U89 ( .A(n13), .B(n14), .Y(SUM[9]) );
  INVX2 U90 ( .A(n25), .Y(n12) );
  NAND2X4 U91 ( .A(n16), .B(n17), .Y(SUM[15]) );
  CLKINVX3 U92 ( .A(n94), .Y(n100) );
  BUFX4 U93 ( .A(n128), .Y(SUM[8]) );
  NAND3BX4 U94 ( .AN(n100), .B(n101), .C(n102), .Y(n98) );
  NAND3X4 U95 ( .A(n108), .B(n76), .C(n77), .Y(n104) );
  OAI21X4 U96 ( .A0(n109), .A1(n110), .B0(n111), .Y(n77) );
  OAI21X2 U97 ( .A0(n36), .A1(n37), .B0(n38), .Y(n32) );
  XOR2X2 U98 ( .A(n32), .B(n33), .Y(SUM[7]) );
  OAI21X2 U99 ( .A0(n64), .A1(n65), .B0(n62), .Y(n126) );
  CLKINVX3 U100 ( .A(n56), .Y(n127) );
  OAI211X2 U101 ( .A0(n126), .A1(n127), .B0(n59), .C0(n53), .Y(n125) );
  NOR2BX1 U102 ( .AN(n56), .B(n55), .Y(n58) );
  NOR2BX1 U103 ( .AN(n38), .B(n37), .Y(n40) );
  NOR2BXL U104 ( .AN(n43), .B(n22), .Y(n45) );
  NAND2BX4 U105 ( .AN(n35), .B(n120), .Y(n81) );
  OR2XL U106 ( .A(A[1]), .B(B[1]), .Y(n60) );
  OAI21X4 U107 ( .A0(n124), .A1(n82), .B0(n81), .Y(n28) );
  CLKINVX3 U108 ( .A(n124), .Y(n47) );
  INVX2 U109 ( .A(n79), .Y(n124) );
  XOR2X2 U110 ( .A(n44), .B(n45), .Y(SUM[5]) );
  NAND3X2 U111 ( .A(n121), .B(n38), .C(n34), .Y(n120) );
  XOR2X1 U112 ( .A(n28), .B(n29), .Y(n128) );
  INVXL U113 ( .A(n53), .Y(n52) );
  OAI2BB1X2 U114 ( .A0N(n60), .A1N(n61), .B0(n62), .Y(n57) );
  XOR2X1 U115 ( .A(n61), .B(n63), .Y(SUM[1]) );
  AOI211X2 U116 ( .A0(n26), .A1(n30), .B0(n10), .C0(n27), .Y(n110) );
  NAND2XL U117 ( .A(B[3]), .B(A[3]), .Y(n51) );
  OR2X4 U118 ( .A(B[13]), .B(A[13]), .Y(n83) );
  NAND2XL U119 ( .A(B[1]), .B(A[1]), .Y(n62) );
  NAND2XL U120 ( .A(B[0]), .B(A[0]), .Y(n65) );
  NOR2BX1 U121 ( .AN(n65), .B(n21), .Y(SUM[0]) );
  NOR2XL U122 ( .A(A[0]), .B(B[0]), .Y(n21) );
  INVX1 U123 ( .A(n81), .Y(n80) );
  INVX1 U124 ( .A(n82), .Y(n78) );
  OAI21XL U125 ( .A0(n73), .A1(n74), .B0(n75), .Y(n72) );
  AOI21X1 U126 ( .A0(n78), .A1(n79), .B0(n80), .Y(n73) );
  NOR2BX1 U127 ( .AN(n34), .B(n35), .Y(n33) );
  INVX1 U128 ( .A(n123), .Y(n35) );
  INVX1 U129 ( .A(n60), .Y(n64) );
  XOR2X1 U130 ( .A(n49), .B(n50), .Y(SUM[3]) );
  OAI21XL U131 ( .A0(n54), .A1(n55), .B0(n56), .Y(n49) );
  NOR2BX1 U132 ( .AN(n51), .B(n52), .Y(n50) );
  INVX1 U133 ( .A(n57), .Y(n54) );
  XOR2X1 U134 ( .A(n47), .B(n48), .Y(SUM[4]) );
  NOR2BX1 U135 ( .AN(n46), .B(n23), .Y(n48) );
  NAND2X2 U136 ( .A(n51), .B(n125), .Y(n79) );
  INVX1 U137 ( .A(n59), .Y(n55) );
  XOR2X2 U138 ( .A(n57), .B(n58), .Y(SUM[2]) );
  NOR2BXL U139 ( .AN(n62), .B(n64), .Y(n63) );
  INVX1 U140 ( .A(n65), .Y(n61) );
  NAND2XL U141 ( .A(B[5]), .B(A[5]), .Y(n43) );
  OR2X4 U142 ( .A(B[14]), .B(A[14]), .Y(n85) );
  XOR2X4 U143 ( .A(n105), .B(n106), .Y(SUM[13]) );
  OR2X4 U144 ( .A(B[10]), .B(A[10]), .Y(n87) );
  OR2X4 U145 ( .A(B[9]), .B(A[9]), .Y(n88) );
endmodule


module butterfly_DW01_sub_90 ( A, B, DIFF );
  input [16:0] A;
  input [16:0] B;
  output [16:0] DIFF;
  wire   n163, n164, n165, n166, n167, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n18, n20, n21, n22, n23, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162;

  BUFX8 U3 ( .A(n113), .Y(n1) );
  BUFX12 U4 ( .A(n111), .Y(n9) );
  CLKBUFX8 U5 ( .A(n100), .Y(n16) );
  BUFX4 U6 ( .A(n119), .Y(n2) );
  BUFX8 U7 ( .A(n99), .Y(n6) );
  BUFX4 U8 ( .A(A[11]), .Y(n11) );
  NAND2BX2 U9 ( .AN(B[11]), .B(n11), .Y(n3) );
  NAND2BX2 U10 ( .AN(B[11]), .B(n11), .Y(n4) );
  BUFX8 U11 ( .A(A[14]), .Y(n10) );
  NAND2BXL U12 ( .AN(n9), .B(n119), .Y(n110) );
  BUFX8 U13 ( .A(n139), .Y(n5) );
  INVX3 U14 ( .A(n89), .Y(n88) );
  NOR2BX4 U15 ( .AN(B[15]), .B(A[15]), .Y(n14) );
  INVX8 U16 ( .A(n116), .Y(n109) );
  NAND2X2 U17 ( .A(n134), .B(n18), .Y(n119) );
  BUFX20 U18 ( .A(n104), .Y(n8) );
  NOR2BX1 U19 ( .AN(n6), .B(n14), .Y(n107) );
  CLKINVX4 U20 ( .A(n106), .Y(n95) );
  INVX4 U21 ( .A(n155), .Y(n58) );
  NOR2X2 U22 ( .A(n77), .B(n81), .Y(n157) );
  NAND4BX2 U23 ( .AN(n58), .B(n65), .C(n49), .D(n52), .Y(n106) );
  NAND2BX4 U24 ( .AN(B[1]), .B(A[1]), .Y(n78) );
  NAND2X2 U25 ( .A(n72), .B(n73), .Y(n21) );
  NAND2BX2 U26 ( .AN(B[3]), .B(A[3]), .Y(n73) );
  AOI21X2 U27 ( .A0(n69), .A1(n70), .B0(n71), .Y(n68) );
  NAND3X2 U28 ( .A(n144), .B(n102), .C(n103), .Y(n142) );
  NAND4X2 U29 ( .A(n102), .B(n145), .C(n43), .D(n103), .Y(n123) );
  INVX4 U30 ( .A(n103), .Y(n150) );
  NAND2X4 U31 ( .A(n97), .B(n98), .Y(n84) );
  INVX8 U32 ( .A(n150), .Y(n7) );
  NAND2X4 U33 ( .A(n52), .B(n53), .Y(n47) );
  OAI21X4 U34 ( .A0(n86), .A1(n87), .B0(n88), .Y(n85) );
  AOI21X2 U35 ( .A0(n15), .A1(n125), .B0(n126), .Y(n124) );
  BUFX12 U36 ( .A(B[13]), .Y(n18) );
  XOR2X4 U37 ( .A(B[16]), .B(A[16]), .Y(n28) );
  INVX1 U38 ( .A(n133), .Y(n12) );
  NOR2X4 U39 ( .A(n94), .B(n89), .Y(n98) );
  INVX8 U40 ( .A(n102), .Y(n41) );
  NAND2X2 U41 ( .A(n158), .B(n82), .Y(DIFF[0]) );
  NAND2BX4 U42 ( .AN(B[0]), .B(A[0]), .Y(n82) );
  AND2X2 U43 ( .A(n12), .B(n113), .Y(n26) );
  AOI21X4 U44 ( .A0(n18), .A1(n134), .B0(n9), .Y(n132) );
  INVX8 U45 ( .A(n122), .Y(n15) );
  INVX8 U46 ( .A(n8), .Y(n122) );
  NAND2X2 U47 ( .A(n101), .B(n100), .Y(n130) );
  XNOR2X4 U48 ( .A(n127), .B(n128), .Y(n165) );
  NAND2X4 U49 ( .A(n139), .B(n100), .Y(n138) );
  INVX2 U50 ( .A(n4), .Y(n126) );
  NAND2X2 U51 ( .A(n112), .B(n9), .Y(n121) );
  NAND2X4 U52 ( .A(n18), .B(n134), .Y(n101) );
  INVX8 U53 ( .A(A[13]), .Y(n134) );
  OR2X4 U54 ( .A(n80), .B(n77), .Y(n35) );
  INVX4 U55 ( .A(n159), .Y(n77) );
  NOR2X4 U56 ( .A(n132), .B(n133), .Y(n131) );
  AOI21X2 U57 ( .A0(n92), .A1(n93), .B0(n94), .Y(n86) );
  NAND4BX2 U58 ( .AN(n45), .B(n102), .C(n7), .D(n15), .Y(n94) );
  NAND2BX4 U59 ( .AN(B[5]), .B(A[5]), .Y(n59) );
  NAND4BX4 U60 ( .AN(n14), .B(n6), .C(n2), .D(n16), .Y(n89) );
  INVX8 U61 ( .A(n145), .Y(n45) );
  XNOR2X4 U62 ( .A(n148), .B(n25), .Y(n13) );
  NAND2BX4 U63 ( .AN(n123), .B(n8), .Y(n141) );
  NAND2X2 U64 ( .A(n136), .B(n91), .Y(n135) );
  NAND2X4 U65 ( .A(n8), .B(n125), .Y(n90) );
  OAI21X2 U66 ( .A0(n122), .A1(n123), .B0(n124), .Y(n120) );
  INVX8 U67 ( .A(n13), .Y(DIFF[10]) );
  AOI21X2 U68 ( .A0(n107), .A1(n108), .B0(n109), .Y(n83) );
  AOI2BB1X2 U69 ( .A0N(n122), .A1N(n123), .B0(n135), .Y(n129) );
  INVX4 U70 ( .A(n112), .Y(n133) );
  NAND2X2 U71 ( .A(n15), .B(n125), .Y(n136) );
  AOI21X2 U72 ( .A0(n7), .A1(n148), .B0(n149), .Y(n147) );
  AOI21X4 U73 ( .A0(n120), .A1(n16), .B0(n121), .Y(n117) );
  BUFX20 U74 ( .A(n167), .Y(DIFF[11]) );
  NAND2BX4 U75 ( .AN(B[15]), .B(A[15]), .Y(n116) );
  NAND2X4 U76 ( .A(n8), .B(n91), .Y(n146) );
  NAND2BX4 U77 ( .AN(B[4]), .B(A[4]), .Y(n63) );
  NAND2BX4 U78 ( .AN(A[4]), .B(B[4]), .Y(n65) );
  AND2X4 U79 ( .A(n138), .B(n111), .Y(n34) );
  XNOR2X4 U80 ( .A(n79), .B(n35), .Y(DIFF[1]) );
  INVX4 U81 ( .A(n143), .Y(n149) );
  NAND2X4 U82 ( .A(n63), .B(n65), .Y(n67) );
  NAND2X2 U83 ( .A(n64), .B(n65), .Y(n62) );
  NAND2BX4 U84 ( .AN(B[12]), .B(A[12]), .Y(n111) );
  BUFX20 U85 ( .A(n163), .Y(DIFF[16]) );
  NAND2X4 U86 ( .A(n142), .B(n143), .Y(n125) );
  NAND2X4 U87 ( .A(n119), .B(n99), .Y(n118) );
  BUFX20 U88 ( .A(n165), .Y(DIFF[14]) );
  NOR2X4 U89 ( .A(n109), .B(n14), .Y(n115) );
  BUFX20 U90 ( .A(n166), .Y(DIFF[13]) );
  BUFX20 U91 ( .A(n164), .Y(DIFF[15]) );
  OAI21X4 U92 ( .A0(n118), .A1(n117), .B0(n1), .Y(n114) );
  NAND2BX4 U93 ( .AN(A[5]), .B(B[5]), .Y(n155) );
  OAI21X4 U94 ( .A0(n45), .A1(n152), .B0(n46), .Y(n39) );
  INVX4 U95 ( .A(n43), .Y(n152) );
  OAI21X1 U96 ( .A0(n76), .A1(n77), .B0(n78), .Y(n70) );
  INVX2 U97 ( .A(n64), .Y(n66) );
  NAND2BX4 U98 ( .AN(A[3]), .B(B[3]), .Y(n72) );
  NAND3X2 U99 ( .A(n154), .B(n56), .C(n53), .Y(n153) );
  NAND2BX4 U100 ( .AN(B[7]), .B(A[7]), .Y(n53) );
  NAND3X1 U101 ( .A(n155), .B(n156), .C(n49), .Y(n154) );
  OAI21X4 U102 ( .A0(n151), .A1(n41), .B0(n42), .Y(n148) );
  INVX2 U103 ( .A(n39), .Y(n151) );
  INVX8 U104 ( .A(n32), .Y(DIFF[8]) );
  XOR2X4 U105 ( .A(n43), .B(n33), .Y(n32) );
  NAND2BX4 U106 ( .AN(B[8]), .B(A[8]), .Y(n46) );
  INVX4 U107 ( .A(n56), .Y(n51) );
  NAND2BX4 U108 ( .AN(A[2]), .B(B[2]), .Y(n69) );
  NAND2X2 U109 ( .A(n26), .B(n110), .Y(n108) );
  INVX2 U110 ( .A(n46), .Y(n44) );
  INVX8 U111 ( .A(n30), .Y(DIFF[9]) );
  AOI21X4 U112 ( .A0(n49), .A1(n50), .B0(n51), .Y(n48) );
  INVX4 U113 ( .A(n49), .Y(n55) );
  NAND2BX4 U114 ( .AN(A[6]), .B(B[6]), .Y(n49) );
  XOR2X4 U115 ( .A(n39), .B(n31), .Y(n30) );
  NAND2XL U116 ( .A(n59), .B(n63), .Y(n156) );
  OR2X4 U117 ( .A(n40), .B(n41), .Y(n31) );
  XOR2X4 U118 ( .A(n34), .B(n137), .Y(n166) );
  XOR2X4 U119 ( .A(n5), .B(n140), .Y(n29) );
  INVX8 U120 ( .A(n29), .Y(DIFF[12]) );
  NAND2BXL U121 ( .AN(A[0]), .B(B[0]), .Y(n158) );
  NAND2X2 U122 ( .A(n52), .B(n153), .Y(n92) );
  NAND2X4 U123 ( .A(n81), .B(n82), .Y(n79) );
  XOR2X4 U124 ( .A(n60), .B(n20), .Y(DIFF[5]) );
  NOR2X4 U125 ( .A(n61), .B(n58), .Y(n20) );
  XOR2X4 U126 ( .A(n21), .B(n68), .Y(DIFF[3]) );
  XOR2X4 U127 ( .A(n70), .B(n22), .Y(DIFF[2]) );
  NOR2X4 U128 ( .A(n71), .B(n74), .Y(n22) );
  NAND3XL U129 ( .A(n23), .B(n78), .C(n75), .Y(n161) );
  NAND2XL U130 ( .A(n162), .B(n159), .Y(n23) );
  NOR2X4 U131 ( .A(n150), .B(n149), .Y(n25) );
  XOR2X4 U132 ( .A(n27), .B(n28), .Y(n163) );
  AND3X4 U133 ( .A(n83), .B(n84), .C(n85), .Y(n27) );
  INVX1 U134 ( .A(n158), .Y(n81) );
  INVX1 U135 ( .A(n82), .Y(n162) );
  NAND2BX4 U136 ( .AN(n96), .B(n105), .Y(n64) );
  NAND2XL U137 ( .A(n95), .B(n96), .Y(n93) );
  OR2X4 U138 ( .A(n44), .B(n45), .Y(n33) );
  NOR2XL U139 ( .A(n105), .B(n106), .Y(n97) );
  NAND2XL U140 ( .A(n3), .B(n90), .Y(n87) );
  NAND2XL U141 ( .A(n42), .B(n46), .Y(n144) );
  INVX1 U142 ( .A(n79), .Y(n76) );
  NAND3X4 U143 ( .A(n69), .B(n72), .C(n157), .Y(n105) );
  CLKINVX3 U144 ( .A(n42), .Y(n40) );
  XOR2X4 U145 ( .A(n47), .B(n48), .Y(DIFF[7]) );
  XOR2X4 U146 ( .A(n50), .B(n54), .Y(DIFF[6]) );
  NOR2X4 U147 ( .A(n51), .B(n55), .Y(n54) );
  OAI21X4 U148 ( .A0(n57), .A1(n58), .B0(n59), .Y(n50) );
  CLKINVX3 U149 ( .A(n60), .Y(n57) );
  CLKINVX3 U150 ( .A(n59), .Y(n61) );
  NAND2X4 U151 ( .A(n62), .B(n63), .Y(n60) );
  XOR2X4 U152 ( .A(n66), .B(n67), .Y(DIFF[4]) );
  CLKINVX3 U153 ( .A(n69), .Y(n74) );
  CLKINVX3 U154 ( .A(n75), .Y(n71) );
  CLKINVX3 U155 ( .A(n78), .Y(n80) );
  XOR2X4 U156 ( .A(n114), .B(n115), .Y(n164) );
  NAND2X4 U157 ( .A(n113), .B(n99), .Y(n128) );
  NAND2BX4 U158 ( .AN(B[14]), .B(n10), .Y(n113) );
  NAND2BX4 U159 ( .AN(A[14]), .B(B[14]), .Y(n99) );
  OAI21X4 U160 ( .A0(n130), .A1(n129), .B0(n131), .Y(n127) );
  NAND2X4 U161 ( .A(n101), .B(n112), .Y(n137) );
  NAND2BX4 U162 ( .AN(B[13]), .B(A[13]), .Y(n112) );
  NAND2X4 U163 ( .A(n111), .B(n100), .Y(n140) );
  NAND2BX4 U164 ( .AN(A[12]), .B(B[12]), .Y(n100) );
  NAND3X4 U165 ( .A(n141), .B(n90), .C(n3), .Y(n139) );
  XOR2X4 U166 ( .A(n146), .B(n147), .Y(n167) );
  NAND2BX4 U167 ( .AN(B[11]), .B(n11), .Y(n91) );
  NAND2BX4 U168 ( .AN(A[11]), .B(B[11]), .Y(n104) );
  NAND2BX4 U169 ( .AN(B[10]), .B(A[10]), .Y(n143) );
  NAND2BX4 U170 ( .AN(A[10]), .B(B[10]), .Y(n103) );
  NAND2BX4 U171 ( .AN(B[9]), .B(A[9]), .Y(n42) );
  NAND2BX4 U172 ( .AN(A[9]), .B(B[9]), .Y(n102) );
  OAI2BB1X4 U173 ( .A0N(n95), .A1N(n64), .B0(n92), .Y(n43) );
  NAND2BX4 U174 ( .AN(B[6]), .B(A[6]), .Y(n56) );
  NAND2X4 U175 ( .A(n160), .B(n73), .Y(n96) );
  NAND3X4 U176 ( .A(n69), .B(n161), .C(n72), .Y(n160) );
  NAND2BX4 U177 ( .AN(B[2]), .B(A[2]), .Y(n75) );
  NAND2BX4 U178 ( .AN(A[1]), .B(B[1]), .Y(n159) );
  NAND2BX4 U179 ( .AN(A[7]), .B(B[7]), .Y(n52) );
  NAND2BX4 U180 ( .AN(A[8]), .B(B[8]), .Y(n145) );
endmodule


module butterfly_DW01_sub_81 ( A, B, DIFF );
  input [16:0] A;
  input [16:0] B;
  output [16:0] DIFF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148;

  NAND2BX1 U3 ( .AN(B[11]), .B(A[11]), .Y(n79) );
  NAND2BX2 U4 ( .AN(A[14]), .B(B[14]), .Y(n1) );
  NAND2BX2 U5 ( .AN(A[14]), .B(B[14]), .Y(n86) );
  INVX4 U6 ( .A(n86), .Y(n2) );
  CLKINVX8 U7 ( .A(n2), .Y(n3) );
  NAND3X4 U8 ( .A(n4), .B(n72), .C(n73), .Y(n71) );
  AND3X4 U9 ( .A(n85), .B(n3), .C(n117), .Y(n4) );
  CLKINVX2 U10 ( .A(B[13]), .Y(n108) );
  NAND2BX2 U11 ( .AN(B[13]), .B(A[13]), .Y(n101) );
  NAND2BX4 U12 ( .AN(A[3]), .B(B[3]), .Y(n53) );
  NAND3X1 U13 ( .A(n117), .B(n73), .C(n112), .Y(n116) );
  OAI21X2 U14 ( .A0(A[13]), .A1(n108), .B0(n101), .Y(n120) );
  INVX8 U15 ( .A(n132), .Y(n26) );
  NAND2BX4 U16 ( .AN(A[8]), .B(B[8]), .Y(n132) );
  CLKINVX4 U17 ( .A(B[15]), .Y(n5) );
  INVX4 U18 ( .A(n5), .Y(n6) );
  CLKINVX2 U19 ( .A(A[13]), .Y(n118) );
  NAND2BX4 U20 ( .AN(A[13]), .B(B[13]), .Y(n73) );
  NAND2BX4 U21 ( .AN(A[12]), .B(B[12]), .Y(n122) );
  NAND2BX2 U22 ( .AN(A[12]), .B(B[12]), .Y(n117) );
  INVX1 U23 ( .A(n68), .Y(n10) );
  INVX2 U24 ( .A(n122), .Y(n12) );
  NOR2X2 U25 ( .A(n43), .B(n39), .Y(n42) );
  CLKINVX3 U26 ( .A(n143), .Y(n64) );
  INVX2 U27 ( .A(n3), .Y(n98) );
  BUFX8 U28 ( .A(n79), .Y(n15) );
  INVX1 U29 ( .A(n12), .Y(n11) );
  AND3X4 U30 ( .A(n124), .B(n15), .C(n80), .Y(n7) );
  NAND3XL U31 ( .A(n147), .B(n60), .C(n57), .Y(n146) );
  OAI21X1 U32 ( .A0(n58), .A1(n59), .B0(n60), .Y(n51) );
  NAND2X4 U33 ( .A(n122), .B(n100), .Y(n18) );
  NAND2BX4 U34 ( .AN(B[12]), .B(A[12]), .Y(n100) );
  NAND2BX2 U35 ( .AN(B[4]), .B(A[4]), .Y(n45) );
  NAND3X2 U36 ( .A(n140), .B(n141), .C(n30), .Y(n139) );
  INVX4 U37 ( .A(n140), .Y(n39) );
  BUFX3 U38 ( .A(n30), .Y(n8) );
  INVX4 U39 ( .A(n37), .Y(n32) );
  NAND2BX1 U40 ( .AN(B[6]), .B(A[6]), .Y(n37) );
  XOR2X4 U41 ( .A(n31), .B(n35), .Y(DIFF[6]) );
  NOR2X2 U42 ( .A(n32), .B(n36), .Y(n35) );
  NOR2X4 U43 ( .A(n22), .B(n23), .Y(n21) );
  INVX8 U44 ( .A(n130), .Y(n22) );
  XOR2X2 U45 ( .A(n41), .B(n42), .Y(DIFF[5]) );
  NAND2X1 U46 ( .A(n46), .B(n47), .Y(n44) );
  XNOR2X4 U47 ( .A(n46), .B(n17), .Y(DIFF[4]) );
  NAND2BX4 U48 ( .AN(n82), .B(n90), .Y(n46) );
  XOR2X4 U49 ( .A(n28), .B(n29), .Y(DIFF[7]) );
  AOI21X2 U50 ( .A0(n8), .A1(n31), .B0(n32), .Y(n29) );
  XOR2X4 U51 ( .A(n7), .B(n18), .Y(DIFF[12]) );
  NAND2X4 U52 ( .A(n15), .B(n93), .Y(n133) );
  XNOR2X4 U53 ( .A(n9), .B(n133), .Y(DIFF[11]) );
  NAND2X2 U54 ( .A(n14), .B(n134), .Y(n9) );
  NAND4BX4 U55 ( .AN(n131), .B(n24), .C(n126), .D(n93), .Y(n124) );
  NAND2X4 U56 ( .A(n14), .B(n126), .Y(n16) );
  NAND4BX2 U57 ( .AN(n26), .B(n92), .C(n126), .D(n93), .Y(n75) );
  NAND2BX4 U58 ( .AN(A[10]), .B(B[10]), .Y(n126) );
  NAND4X4 U59 ( .A(n70), .B(n71), .C(n69), .D(n10), .Y(n66) );
  XNOR2X4 U60 ( .A(n135), .B(n16), .Y(DIFF[10]) );
  NAND3X4 U61 ( .A(n11), .B(n87), .C(n88), .Y(n70) );
  NOR2X4 U62 ( .A(n97), .B(n98), .Y(n96) );
  AOI21X2 U63 ( .A0(n112), .A1(n122), .B0(n123), .Y(n121) );
  NAND2BX4 U64 ( .AN(B[9]), .B(A[9]), .Y(n130) );
  INVX4 U65 ( .A(n102), .Y(n94) );
  NAND2BX4 U66 ( .AN(B[14]), .B(A[14]), .Y(n102) );
  OAI21X2 U67 ( .A0(A[13]), .A1(n108), .B0(n1), .Y(n107) );
  OAI2BB1X2 U68 ( .A0N(B[13]), .A1N(n118), .B0(n119), .Y(n115) );
  XNOR2X2 U69 ( .A(B[16]), .B(A[16]), .Y(n67) );
  NAND2BX1 U70 ( .AN(B[15]), .B(A[15]), .Y(n105) );
  NAND2BX4 U71 ( .AN(B[7]), .B(A[7]), .Y(n34) );
  OAI2BB1X1 U72 ( .A0N(A[12]), .A1N(n113), .B0(n101), .Y(n109) );
  INVX4 U73 ( .A(n85), .Y(n97) );
  OAI21X4 U74 ( .A0(n94), .A1(n95), .B0(n96), .Y(n69) );
  NAND2X4 U75 ( .A(n3), .B(n85), .Y(n89) );
  NAND2XL U76 ( .A(n40), .B(n45), .Y(n141) );
  INVXL U77 ( .A(B[12]), .Y(n113) );
  NAND2BX4 U78 ( .AN(B[8]), .B(A[8]), .Y(n129) );
  XOR2X2 U79 ( .A(n24), .B(n25), .Y(DIFF[8]) );
  NOR2X2 U80 ( .A(n26), .B(n27), .Y(n25) );
  NOR2X4 U81 ( .A(n13), .B(n89), .Y(n88) );
  NAND2BX2 U82 ( .AN(B[10]), .B(A[10]), .Y(n128) );
  INVX4 U83 ( .A(n92), .Y(n23) );
  NOR2X2 U84 ( .A(n109), .B(n110), .Y(n106) );
  NOR2BXL U85 ( .AN(B[13]), .B(A[13]), .Y(n99) );
  OAI21X4 U86 ( .A0(n38), .A1(n39), .B0(n40), .Y(n31) );
  NAND2X2 U87 ( .A(n126), .B(n135), .Y(n134) );
  NAND3BX4 U88 ( .AN(n22), .B(n127), .C(n14), .Y(n125) );
  AOI21X2 U89 ( .A0(n111), .A1(B[12]), .B0(n7), .Y(n110) );
  NOR2BX1 U90 ( .AN(A[12]), .B(B[12]), .Y(n119) );
  INVX4 U91 ( .A(n24), .Y(n137) );
  NOR2X4 U92 ( .A(n97), .B(n68), .Y(n104) );
  INVX4 U93 ( .A(n105), .Y(n68) );
  NAND2X4 U94 ( .A(n1), .B(n102), .Y(n114) );
  INVX4 U95 ( .A(n20), .Y(n136) );
  AOI21X1 U96 ( .A0(n81), .A1(n82), .B0(n83), .Y(n74) );
  CLKINVX4 U97 ( .A(n91), .Y(n81) );
  NAND2BX2 U98 ( .AN(A[5]), .B(B[5]), .Y(n140) );
  NAND2BX4 U99 ( .AN(B[5]), .B(A[5]), .Y(n40) );
  BUFX8 U100 ( .A(n128), .Y(n14) );
  XOR2X4 U101 ( .A(n120), .B(n121), .Y(DIFF[13]) );
  NAND3X4 U102 ( .A(n93), .B(n126), .C(n125), .Y(n80) );
  OAI21X4 U103 ( .A0(n106), .A1(n107), .B0(n102), .Y(n103) );
  INVX2 U104 ( .A(n100), .Y(n123) );
  XOR2X4 U105 ( .A(n103), .B(n104), .Y(DIFF[15]) );
  NAND2BX4 U106 ( .AN(A[15]), .B(n6), .Y(n85) );
  XOR2X4 U107 ( .A(n66), .B(n67), .Y(DIFF[16]) );
  AND3X4 U108 ( .A(n101), .B(n115), .C(n116), .Y(n19) );
  XOR2X4 U109 ( .A(n19), .B(n114), .Y(DIFF[14]) );
  NAND2BX4 U110 ( .AN(A[9]), .B(B[9]), .Y(n92) );
  INVX4 U111 ( .A(n129), .Y(n27) );
  OAI21X4 U112 ( .A0(n26), .A1(n137), .B0(n129), .Y(n20) );
  XOR2X2 U113 ( .A(n51), .B(n55), .Y(DIFF[2]) );
  INVX2 U114 ( .A(n61), .Y(n58) );
  INVX2 U115 ( .A(n144), .Y(n59) );
  NAND2BX4 U116 ( .AN(A[2]), .B(B[2]), .Y(n50) );
  NAND2BX4 U117 ( .AN(A[7]), .B(B[7]), .Y(n33) );
  OAI21X4 U118 ( .A0(n23), .A1(n136), .B0(n130), .Y(n135) );
  AND2X1 U119 ( .A(n118), .B(B[13]), .Y(n13) );
  OAI2BB1X4 U120 ( .A0N(n81), .A1N(n46), .B0(n84), .Y(n24) );
  NAND2BX2 U121 ( .AN(A[6]), .B(B[6]), .Y(n30) );
  INVX2 U122 ( .A(n41), .Y(n38) );
  NAND3X1 U123 ( .A(n50), .B(n53), .C(n142), .Y(n90) );
  NAND2XL U124 ( .A(n64), .B(n65), .Y(n61) );
  NAND2X4 U125 ( .A(n33), .B(n138), .Y(n84) );
  INVX1 U126 ( .A(n65), .Y(n148) );
  XOR2X2 U127 ( .A(n20), .B(n21), .Y(DIFF[9]) );
  NAND3X4 U128 ( .A(n124), .B(n15), .C(n80), .Y(n112) );
  NAND4BX2 U129 ( .AN(n39), .B(n47), .C(n30), .D(n33), .Y(n91) );
  NOR2X2 U130 ( .A(n59), .B(n64), .Y(n142) );
  NAND2X2 U131 ( .A(n145), .B(n54), .Y(n82) );
  NAND3X2 U132 ( .A(n50), .B(n146), .C(n53), .Y(n145) );
  NAND2XL U133 ( .A(n148), .B(n144), .Y(n147) );
  NAND3X2 U134 ( .A(n139), .B(n37), .C(n34), .Y(n138) );
  INVXL U135 ( .A(n80), .Y(n77) );
  NAND2XL U136 ( .A(n45), .B(n47), .Y(n17) );
  INVXL U137 ( .A(n50), .Y(n56) );
  NAND2XL U138 ( .A(n53), .B(n54), .Y(n48) );
  INVXL U139 ( .A(n57), .Y(n52) );
  NAND2BXL U140 ( .AN(B[1]), .B(A[1]), .Y(n60) );
  NAND2XL U141 ( .A(n143), .B(n65), .Y(DIFF[0]) );
  OAI21XL U142 ( .A0(n74), .A1(n75), .B0(n76), .Y(n72) );
  NOR2X1 U143 ( .A(n77), .B(n78), .Y(n76) );
  INVX1 U144 ( .A(n84), .Y(n83) );
  NAND2X1 U145 ( .A(n132), .B(n92), .Y(n131) );
  INVX1 U146 ( .A(n30), .Y(n36) );
  NAND2X1 U147 ( .A(n33), .B(n34), .Y(n28) );
  INVX1 U148 ( .A(n40), .Y(n43) );
  INVX1 U149 ( .A(n15), .Y(n78) );
  NOR2X1 U150 ( .A(n52), .B(n56), .Y(n55) );
  XOR2X1 U151 ( .A(n48), .B(n49), .Y(DIFF[3]) );
  AOI21XL U152 ( .A0(n50), .A1(n51), .B0(n52), .Y(n49) );
  XOR2X1 U153 ( .A(n61), .B(n62), .Y(DIFF[1]) );
  NOR2XL U154 ( .A(n63), .B(n59), .Y(n62) );
  INVX1 U155 ( .A(n60), .Y(n63) );
  NAND2X2 U156 ( .A(n44), .B(n45), .Y(n41) );
  NAND2XL U157 ( .A(n27), .B(n92), .Y(n127) );
  OAI21XL U158 ( .A0(n99), .A1(n100), .B0(n101), .Y(n95) );
  NAND2BX1 U159 ( .AN(A[4]), .B(B[4]), .Y(n47) );
  NAND2BX1 U160 ( .AN(B[3]), .B(A[3]), .Y(n54) );
  NAND2BXL U161 ( .AN(A[1]), .B(B[1]), .Y(n144) );
  NAND2BX1 U162 ( .AN(B[2]), .B(A[2]), .Y(n57) );
  NOR3XL U163 ( .A(n90), .B(n75), .C(n91), .Y(n87) );
  NAND2BX1 U164 ( .AN(B[0]), .B(A[0]), .Y(n65) );
  NAND2BX1 U165 ( .AN(A[0]), .B(B[0]), .Y(n143) );
  INVXL U166 ( .A(A[12]), .Y(n111) );
  NAND2BX4 U167 ( .AN(A[11]), .B(B[11]), .Y(n93) );
endmodule


module butterfly_DW01_add_104 ( A, B, SUM );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  wire   n126, n127, n1, n3, n5, n6, n7, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125;

  INVX16 U2 ( .A(n73), .Y(n93) );
  OR2X4 U3 ( .A(A[15]), .B(B[15]), .Y(n1) );
  NAND2X4 U4 ( .A(n81), .B(n82), .Y(n80) );
  BUFX20 U5 ( .A(n127), .Y(SUM[13]) );
  XOR2X4 U6 ( .A(n97), .B(n98), .Y(n127) );
  NAND2X2 U7 ( .A(n74), .B(n82), .Y(n97) );
  INVX2 U8 ( .A(n85), .Y(n114) );
  INVX3 U9 ( .A(n78), .Y(n15) );
  AOI21X1 U10 ( .A0(n68), .A1(n69), .B0(n70), .Y(n65) );
  INVX2 U11 ( .A(n6), .Y(n7) );
  INVX1 U12 ( .A(n23), .Y(n10) );
  NOR2BX2 U13 ( .AN(n43), .B(n17), .Y(n44) );
  XNOR2X4 U14 ( .A(n92), .B(n90), .Y(n3) );
  XOR2X2 U15 ( .A(n23), .B(n24), .Y(SUM[8]) );
  XOR2X2 U16 ( .A(n34), .B(n35), .Y(SUM[6]) );
  XOR2X4 U17 ( .A(n27), .B(n28), .Y(SUM[7]) );
  NAND4BBX4 U18 ( .AN(n38), .BN(n17), .C(n36), .D(n120), .Y(n72) );
  OAI21X4 U19 ( .A0(n17), .A1(n42), .B0(n43), .Y(n40) );
  NOR2X2 U20 ( .A(A[4]), .B(B[4]), .Y(n17) );
  AOI21X2 U21 ( .A0(B[11]), .A1(A[11]), .B0(n106), .Y(n105) );
  INVX8 U22 ( .A(n84), .Y(n22) );
  NOR2BX2 U23 ( .AN(n107), .B(n114), .Y(n113) );
  NOR2BX4 U24 ( .AN(n83), .B(n96), .Y(n98) );
  INVX8 U25 ( .A(n3), .Y(SUM[14]) );
  OR2XL U26 ( .A(A[14]), .B(B[14]), .Y(n5) );
  NAND2X4 U27 ( .A(B[14]), .B(A[14]), .Y(n81) );
  NAND2X4 U28 ( .A(n116), .B(n25), .Y(n19) );
  NAND2X4 U29 ( .A(n23), .B(n87), .Y(n116) );
  XNOR2X4 U30 ( .A(n108), .B(n109), .Y(SUM[11]) );
  NAND2X2 U31 ( .A(n107), .B(n111), .Y(n108) );
  NOR2BX4 U32 ( .AN(n81), .B(n93), .Y(n92) );
  NAND2X4 U33 ( .A(n1), .B(n73), .Y(n77) );
  NAND2X1 U34 ( .A(n78), .B(n75), .Y(n88) );
  NAND2X1 U35 ( .A(n64), .B(n63), .Y(n6) );
  NAND2X4 U36 ( .A(n16), .B(n7), .Y(n62) );
  OAI21X2 U37 ( .A0(n65), .A1(n66), .B0(n67), .Y(n63) );
  OR2X4 U38 ( .A(B[12]), .B(A[12]), .Y(n64) );
  XOR2X4 U39 ( .A(n19), .B(n20), .Y(SUM[9]) );
  NOR2BX2 U40 ( .AN(n21), .B(n22), .Y(n20) );
  BUFX20 U41 ( .A(n126), .Y(SUM[15]) );
  NAND2X4 U42 ( .A(n86), .B(n101), .Y(n100) );
  NAND2X2 U43 ( .A(n83), .B(n64), .Y(n102) );
  NAND2X2 U44 ( .A(B[13]), .B(A[13]), .Y(n82) );
  NAND2X1 U45 ( .A(A[15]), .B(B[15]), .Y(n78) );
  NOR2X4 U46 ( .A(n79), .B(n80), .Y(n76) );
  OR2X4 U47 ( .A(B[11]), .B(A[11]), .Y(n9) );
  NAND4BBX4 U48 ( .AN(n11), .BN(n10), .C(n85), .D(n86), .Y(n99) );
  NAND2XL U49 ( .A(n87), .B(n84), .Y(n11) );
  NAND4BX1 U50 ( .AN(n26), .B(n84), .C(n85), .D(n9), .Y(n66) );
  NAND2X2 U51 ( .A(n9), .B(n110), .Y(n109) );
  OAI2BB1X4 U52 ( .A0N(n85), .A1N(n104), .B0(n105), .Y(n101) );
  NAND2X4 U53 ( .A(B[9]), .B(A[9]), .Y(n21) );
  NOR2BX4 U54 ( .AN(n74), .B(n83), .Y(n79) );
  OAI21X1 U55 ( .A0(n31), .A1(n32), .B0(n33), .Y(n27) );
  OAI21X2 U56 ( .A0(n22), .A1(n25), .B0(n21), .Y(n104) );
  OAI21X4 U57 ( .A0(n42), .A1(n72), .B0(n71), .Y(n23) );
  XOR2X4 U58 ( .A(n112), .B(n113), .Y(SUM[10]) );
  OAI21X4 U59 ( .A0(n22), .A1(n115), .B0(n21), .Y(n112) );
  NAND2X2 U60 ( .A(n99), .B(n67), .Y(n103) );
  NAND2X2 U61 ( .A(n9), .B(n101), .Y(n67) );
  AOI2BB2X4 U62 ( .B0(n99), .B1(n100), .A0N(B[12]), .A1N(A[12]), .Y(n96) );
  INVX2 U63 ( .A(n19), .Y(n115) );
  NAND2X4 U64 ( .A(B[4]), .B(A[4]), .Y(n43) );
  OAI21X4 U65 ( .A0(n95), .A1(n96), .B0(n74), .Y(n94) );
  INVX4 U66 ( .A(n83), .Y(n95) );
  NAND2X4 U67 ( .A(B[10]), .B(A[10]), .Y(n107) );
  XNOR2X4 U68 ( .A(n102), .B(n103), .Y(SUM[12]) );
  INVXL U69 ( .A(n81), .Y(n91) );
  AND3X4 U70 ( .A(n73), .B(n75), .C(n74), .Y(n16) );
  AOI2BB1X4 U71 ( .A0N(n76), .A1N(n77), .B0(n15), .Y(n14) );
  INVX4 U72 ( .A(n69), .Y(n42) );
  NAND2BX4 U73 ( .AN(n30), .B(n12), .Y(n71) );
  NAND3X2 U74 ( .A(n117), .B(n33), .C(n29), .Y(n12) );
  OAI2BB1XL U75 ( .A0N(n55), .A1N(n56), .B0(n57), .Y(n52) );
  XOR2X4 U76 ( .A(n88), .B(n89), .Y(n126) );
  NAND2X1 U77 ( .A(B[6]), .B(A[6]), .Y(n33) );
  NAND2X1 U78 ( .A(B[3]), .B(A[3]), .Y(n47) );
  NOR2BX1 U79 ( .AN(n60), .B(n13), .Y(SUM[0]) );
  NOR2XL U80 ( .A(A[0]), .B(B[0]), .Y(n13) );
  INVX1 U81 ( .A(n72), .Y(n68) );
  INVX1 U82 ( .A(n71), .Y(n70) );
  INVX1 U83 ( .A(n52), .Y(n49) );
  INVXL U84 ( .A(n87), .Y(n26) );
  NAND2XL U85 ( .A(n85), .B(n112), .Y(n111) );
  NOR2BXL U86 ( .AN(n29), .B(n30), .Y(n28) );
  INVX1 U87 ( .A(n34), .Y(n31) );
  NOR2BX1 U88 ( .AN(n25), .B(n26), .Y(n24) );
  XOR2X1 U89 ( .A(n40), .B(n41), .Y(SUM[5]) );
  NOR2BXL U90 ( .AN(n39), .B(n38), .Y(n41) );
  OAI21XL U91 ( .A0(n37), .A1(n38), .B0(n39), .Y(n34) );
  INVX1 U92 ( .A(n40), .Y(n37) );
  INVXL U93 ( .A(n36), .Y(n32) );
  NOR2BXL U94 ( .AN(n33), .B(n32), .Y(n35) );
  XOR2X1 U95 ( .A(n45), .B(n46), .Y(SUM[3]) );
  NOR2BX1 U96 ( .AN(n47), .B(n48), .Y(n46) );
  OAI21XL U97 ( .A0(n49), .A1(n50), .B0(n51), .Y(n45) );
  INVXL U98 ( .A(n121), .Y(n48) );
  XOR2X1 U99 ( .A(n69), .B(n44), .Y(SUM[4]) );
  INVXL U100 ( .A(n54), .Y(n50) );
  XOR2X1 U101 ( .A(n56), .B(n58), .Y(SUM[1]) );
  NOR2BXL U102 ( .AN(n57), .B(n59), .Y(n58) );
  XOR2X1 U103 ( .A(n52), .B(n53), .Y(SUM[2]) );
  NOR2BX1 U104 ( .AN(n51), .B(n50), .Y(n53) );
  INVXL U105 ( .A(n60), .Y(n56) );
  INVX2 U106 ( .A(n107), .Y(n106) );
  NAND2XL U107 ( .A(A[11]), .B(B[11]), .Y(n110) );
  NAND2X1 U108 ( .A(B[7]), .B(A[7]), .Y(n29) );
  NAND2X2 U109 ( .A(B[5]), .B(A[5]), .Y(n39) );
  NAND2X1 U110 ( .A(B[1]), .B(A[1]), .Y(n57) );
  XNOR2X4 U111 ( .A(n61), .B(n18), .Y(SUM[16]) );
  XNOR2X4 U112 ( .A(B[16]), .B(A[16]), .Y(n18) );
  AOI21X4 U113 ( .A0(n90), .A1(n5), .B0(n91), .Y(n89) );
  NAND2X4 U114 ( .A(n14), .B(n62), .Y(n61) );
  OR2X4 U115 ( .A(A[15]), .B(B[15]), .Y(n75) );
  OR2X4 U116 ( .A(B[14]), .B(A[14]), .Y(n73) );
  NAND2X4 U117 ( .A(n82), .B(n94), .Y(n90) );
  OR2X4 U118 ( .A(A[13]), .B(B[13]), .Y(n74) );
  NAND2X4 U119 ( .A(B[12]), .B(A[12]), .Y(n83) );
  OR2X4 U120 ( .A(B[11]), .B(A[11]), .Y(n86) );
  OR2X4 U121 ( .A(A[10]), .B(B[10]), .Y(n85) );
  NAND2X4 U122 ( .A(B[8]), .B(A[8]), .Y(n25) );
  OR2X4 U123 ( .A(B[8]), .B(A[8]), .Y(n87) );
  NAND3X4 U124 ( .A(n118), .B(n36), .C(n119), .Y(n117) );
  NAND2X4 U125 ( .A(n39), .B(n43), .Y(n119) );
  CLKINVX3 U126 ( .A(n120), .Y(n30) );
  OR2X4 U127 ( .A(A[7]), .B(B[7]), .Y(n120) );
  OR2X4 U128 ( .A(A[6]), .B(B[6]), .Y(n36) );
  CLKINVX3 U129 ( .A(n118), .Y(n38) );
  OR2X4 U130 ( .A(A[5]), .B(B[5]), .Y(n118) );
  OAI21X4 U131 ( .A0(n122), .A1(n123), .B0(n47), .Y(n69) );
  NAND2X4 U132 ( .A(n54), .B(n121), .Y(n123) );
  OR2X4 U133 ( .A(A[3]), .B(B[3]), .Y(n121) );
  OR2X4 U134 ( .A(A[2]), .B(B[2]), .Y(n54) );
  NOR2X4 U135 ( .A(n124), .B(n125), .Y(n122) );
  OAI21X4 U136 ( .A0(n59), .A1(n60), .B0(n57), .Y(n125) );
  CLKINVX3 U137 ( .A(n55), .Y(n59) );
  OR2X4 U138 ( .A(A[1]), .B(B[1]), .Y(n55) );
  CLKINVX3 U139 ( .A(n51), .Y(n124) );
  NAND2X4 U140 ( .A(B[2]), .B(A[2]), .Y(n51) );
  OR2X4 U141 ( .A(A[9]), .B(B[9]), .Y(n84) );
  NAND2X4 U142 ( .A(B[0]), .B(A[0]), .Y(n60) );
endmodule


module butterfly_DW01_sub_91 ( A, B, DIFF );
  input [16:0] A;
  input [16:0] B;
  output [16:0] DIFF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136;

  INVX8 U3 ( .A(n103), .Y(n5) );
  INVX8 U4 ( .A(n86), .Y(n92) );
  INVX2 U5 ( .A(A[14]), .Y(n108) );
  INVX8 U6 ( .A(n20), .Y(n1) );
  BUFX20 U7 ( .A(n85), .Y(n20) );
  INVX2 U8 ( .A(n20), .Y(n95) );
  NAND2BX2 U9 ( .AN(B[10]), .B(A[10]), .Y(n117) );
  NAND3X4 U10 ( .A(n103), .B(n20), .C(n8), .Y(n70) );
  NAND2BX2 U11 ( .AN(A[4]), .B(B[4]), .Y(n48) );
  BUFX4 U12 ( .A(A[8]), .Y(n2) );
  INVX4 U13 ( .A(n42), .Y(n39) );
  NAND2BX2 U14 ( .AN(B[6]), .B(A[6]), .Y(n38) );
  INVX4 U15 ( .A(n118), .Y(n125) );
  NAND4BX1 U16 ( .AN(n29), .B(n99), .C(n118), .D(n119), .Y(n74) );
  BUFX8 U17 ( .A(A[15]), .Y(n3) );
  NAND2BX4 U18 ( .AN(A[11]), .B(B[11]), .Y(n119) );
  NAND3X4 U19 ( .A(n6), .B(n99), .C(n118), .Y(n116) );
  CLKBUFX2 U20 ( .A(n106), .Y(n4) );
  NAND2X2 U21 ( .A(n20), .B(n94), .Y(n113) );
  NAND3X1 U22 ( .A(n129), .B(n130), .C(n36), .Y(n128) );
  NAND2X4 U23 ( .A(n105), .B(n96), .Y(n16) );
  XOR2X2 U24 ( .A(n52), .B(n56), .Y(DIFF[2]) );
  NOR2X1 U25 ( .A(n53), .B(n57), .Y(n56) );
  INVX4 U26 ( .A(n99), .Y(n24) );
  NAND2X2 U27 ( .A(n120), .B(n99), .Y(n15) );
  AND2X4 U28 ( .A(n93), .B(n84), .Y(n110) );
  NAND2BX1 U29 ( .AN(B[7]), .B(A[7]), .Y(n33) );
  CLKINVX4 U30 ( .A(n136), .Y(n80) );
  NAND4BX2 U31 ( .AN(n40), .B(n48), .C(n36), .D(n35), .Y(n136) );
  BUFX12 U32 ( .A(B[14]), .Y(n7) );
  NAND2BX4 U33 ( .AN(A[14]), .B(n7), .Y(n103) );
  XOR2X4 U34 ( .A(n4), .B(n114), .Y(DIFF[12]) );
  NAND2BX4 U35 ( .AN(A[7]), .B(B[7]), .Y(n35) );
  AND3X4 U36 ( .A(n103), .B(n8), .C(n20), .Y(n11) );
  NOR2BX4 U37 ( .AN(n72), .B(n112), .Y(n114) );
  XOR2X2 U38 ( .A(n26), .B(n27), .Y(DIFF[8]) );
  AOI21X2 U39 ( .A0(n118), .A1(n122), .B0(n123), .Y(n121) );
  NAND2X1 U40 ( .A(n25), .B(n30), .Y(n6) );
  NAND2BX4 U41 ( .AN(A[15]), .B(B[15]), .Y(n86) );
  NAND2BX4 U42 ( .AN(A[13]), .B(B[13]), .Y(n85) );
  AOI21X4 U43 ( .A0(n108), .A1(n7), .B0(n94), .Y(n107) );
  NAND2BX4 U44 ( .AN(A[15]), .B(B[15]), .Y(n8) );
  BUFX3 U45 ( .A(n94), .Y(n9) );
  NAND2BX4 U46 ( .AN(B[12]), .B(A[12]), .Y(n96) );
  NAND3X4 U47 ( .A(n20), .B(n84), .C(n104), .Y(n102) );
  CLKINVX3 U48 ( .A(n87), .Y(n10) );
  OR2X4 U49 ( .A(n1), .B(n96), .Y(n12) );
  NAND2BX4 U50 ( .AN(A[12]), .B(B[12]), .Y(n72) );
  NAND3BX4 U51 ( .AN(n70), .B(n71), .C(n72), .Y(n69) );
  NAND2BX4 U52 ( .AN(B[11]), .B(A[11]), .Y(n78) );
  AOI21X4 U53 ( .A0(n11), .A1(n10), .B0(n88), .Y(n68) );
  NAND4BX2 U54 ( .AN(n15), .B(n26), .C(n118), .D(n119), .Y(n115) );
  AND2X4 U55 ( .A(n93), .B(n94), .Y(n13) );
  NAND2BX4 U56 ( .AN(B[13]), .B(A[13]), .Y(n94) );
  NAND2X4 U57 ( .A(n89), .B(n90), .Y(n88) );
  NOR2BX4 U58 ( .AN(n93), .B(n107), .Y(n101) );
  NAND2BX4 U59 ( .AN(B[15]), .B(n3), .Y(n90) );
  OAI2BB1X4 U60 ( .A0N(n21), .A1N(n99), .B0(n25), .Y(n122) );
  INVX4 U61 ( .A(n117), .Y(n123) );
  NAND2BX2 U62 ( .AN(B[5]), .B(A[5]), .Y(n41) );
  XNOR2X4 U63 ( .A(B[16]), .B(A[16]), .Y(n67) );
  OAI2BB1X4 U64 ( .A0N(n12), .A1N(n13), .B0(n91), .Y(n89) );
  NAND2X4 U65 ( .A(n101), .B(n102), .Y(n17) );
  OAI21X4 U66 ( .A0(n95), .A1(n111), .B0(n9), .Y(n109) );
  INVX1 U67 ( .A(n41), .Y(n44) );
  NAND2X1 U68 ( .A(n41), .B(n46), .Y(n130) );
  NAND2X4 U69 ( .A(n105), .B(n96), .Y(n104) );
  NAND2X4 U70 ( .A(n106), .B(n72), .Y(n105) );
  NAND2BX4 U71 ( .AN(B[8]), .B(n2), .Y(n30) );
  NAND2X4 U72 ( .A(n90), .B(n8), .Y(n100) );
  NAND2BX4 U73 ( .AN(A[9]), .B(B[9]), .Y(n99) );
  XOR2X4 U74 ( .A(n66), .B(n67), .Y(DIFF[16]) );
  NAND2X4 U75 ( .A(n68), .B(n69), .Y(n66) );
  NAND2X4 U76 ( .A(n35), .B(n127), .Y(n83) );
  NAND3X2 U77 ( .A(n128), .B(n38), .C(n33), .Y(n127) );
  NAND2BX4 U78 ( .AN(A[0]), .B(B[0]), .Y(n65) );
  AOI21X2 U79 ( .A0(n51), .A1(n52), .B0(n53), .Y(n50) );
  OAI21X4 U80 ( .A0(n58), .A1(n59), .B0(n60), .Y(n52) );
  INVXL U81 ( .A(n61), .Y(n58) );
  NAND2BX4 U82 ( .AN(B[1]), .B(A[1]), .Y(n60) );
  XNOR2X4 U83 ( .A(n17), .B(n100), .Y(DIFF[15]) );
  AOI21X2 U84 ( .A0(n106), .A1(n72), .B0(n112), .Y(n111) );
  NAND2BX4 U85 ( .AN(A[10]), .B(B[10]), .Y(n118) );
  OAI21X2 U86 ( .A0(n39), .A1(n40), .B0(n41), .Y(n37) );
  NOR2X4 U87 ( .A(n92), .B(n5), .Y(n91) );
  NAND2BX4 U88 ( .AN(B[9]), .B(A[9]), .Y(n25) );
  NAND2BX4 U89 ( .AN(B[14]), .B(A[14]), .Y(n93) );
  NAND2BX4 U90 ( .AN(A[14]), .B(n7), .Y(n84) );
  INVX4 U91 ( .A(n96), .Y(n112) );
  XNOR2X4 U92 ( .A(n113), .B(n16), .Y(DIFF[13]) );
  XOR2X2 U93 ( .A(n42), .B(n43), .Y(DIFF[5]) );
  INVX4 U94 ( .A(n35), .Y(n34) );
  NAND2X4 U95 ( .A(n45), .B(n46), .Y(n42) );
  NAND2X4 U96 ( .A(n47), .B(n48), .Y(n45) );
  NOR2X4 U97 ( .A(n28), .B(n29), .Y(n27) );
  XOR2X2 U98 ( .A(n37), .B(n19), .Y(DIFF[6]) );
  AND2X2 U99 ( .A(n38), .B(n36), .Y(n19) );
  OAI2BB1X2 U100 ( .A0N(n36), .A1N(n37), .B0(n38), .Y(n31) );
  INVX4 U101 ( .A(n30), .Y(n28) );
  NOR2X2 U102 ( .A(n44), .B(n40), .Y(n43) );
  XNOR2X1 U103 ( .A(n47), .B(n14), .Y(DIFF[4]) );
  NAND2XL U104 ( .A(n46), .B(n48), .Y(n14) );
  XOR2X1 U105 ( .A(n61), .B(n62), .Y(DIFF[1]) );
  INVXL U106 ( .A(n60), .Y(n63) );
  INVXL U107 ( .A(n51), .Y(n57) );
  NAND2XL U108 ( .A(n54), .B(n55), .Y(n49) );
  NAND4X2 U109 ( .A(n51), .B(n131), .C(n54), .D(n65), .Y(n98) );
  INVXL U110 ( .A(n79), .Y(n76) );
  XNOR2X4 U111 ( .A(n18), .B(n121), .Y(DIFF[11]) );
  AND2X2 U112 ( .A(n119), .B(n78), .Y(n18) );
  XOR2X2 U113 ( .A(n31), .B(n32), .Y(DIFF[7]) );
  OAI21XL U114 ( .A0(n73), .A1(n74), .B0(n75), .Y(n71) );
  AOI21XL U115 ( .A0(n80), .A1(n81), .B0(n82), .Y(n73) );
  NOR2X1 U116 ( .A(n76), .B(n77), .Y(n75) );
  INVX1 U117 ( .A(n83), .Y(n82) );
  INVXL U118 ( .A(n78), .Y(n77) );
  NAND2BX4 U119 ( .AN(n81), .B(n98), .Y(n47) );
  NOR2XL U120 ( .A(n63), .B(n59), .Y(n62) );
  INVX1 U121 ( .A(n98), .Y(n97) );
  NAND2BX1 U122 ( .AN(A[2]), .B(B[2]), .Y(n51) );
  INVX1 U123 ( .A(n135), .Y(n53) );
  NAND2BX1 U124 ( .AN(B[2]), .B(A[2]), .Y(n135) );
  NAND2BX1 U125 ( .AN(A[3]), .B(B[3]), .Y(n54) );
  NAND2BX1 U126 ( .AN(B[3]), .B(A[3]), .Y(n55) );
  NAND2BXL U127 ( .AN(n65), .B(n64), .Y(n61) );
  NAND2XL U128 ( .A(n65), .B(n64), .Y(DIFF[0]) );
  NAND4BXL U129 ( .AN(n74), .B(n97), .C(n80), .D(n72), .Y(n87) );
  XOR2X4 U130 ( .A(n21), .B(n22), .Y(DIFF[9]) );
  NOR2X4 U131 ( .A(n23), .B(n24), .Y(n22) );
  CLKINVX3 U132 ( .A(n25), .Y(n23) );
  NOR2BX4 U133 ( .AN(n33), .B(n34), .Y(n32) );
  XOR2X4 U134 ( .A(n49), .B(n50), .Y(DIFF[3]) );
  XOR2X4 U135 ( .A(n109), .B(n110), .Y(DIFF[14]) );
  NAND3X4 U136 ( .A(n115), .B(n78), .C(n79), .Y(n106) );
  OAI2BB1X4 U137 ( .A0N(n117), .A1N(n116), .B0(n119), .Y(n79) );
  XOR2X4 U138 ( .A(n122), .B(n124), .Y(DIFF[10]) );
  NOR2X4 U139 ( .A(n125), .B(n123), .Y(n124) );
  OAI21X4 U140 ( .A0(n29), .A1(n126), .B0(n30), .Y(n21) );
  CLKINVX3 U141 ( .A(n26), .Y(n126) );
  OAI2BB1X4 U142 ( .A0N(n80), .A1N(n47), .B0(n83), .Y(n26) );
  NAND2BX4 U143 ( .AN(B[4]), .B(A[4]), .Y(n46) );
  OAI21X4 U144 ( .A0(n132), .A1(n133), .B0(n55), .Y(n81) );
  NAND2X4 U145 ( .A(n51), .B(n54), .Y(n133) );
  NOR2X4 U146 ( .A(n53), .B(n134), .Y(n132) );
  OAI21X4 U147 ( .A0(n59), .A1(n64), .B0(n60), .Y(n134) );
  CLKINVX3 U148 ( .A(n131), .Y(n59) );
  NAND2BX4 U149 ( .AN(A[1]), .B(B[1]), .Y(n131) );
  NAND2BX4 U150 ( .AN(A[6]), .B(B[6]), .Y(n36) );
  CLKINVX3 U151 ( .A(n129), .Y(n40) );
  NAND2BX4 U152 ( .AN(A[5]), .B(B[5]), .Y(n129) );
  CLKINVX3 U153 ( .A(n120), .Y(n29) );
  NAND2BX4 U154 ( .AN(A[8]), .B(B[8]), .Y(n120) );
  NAND2BX4 U155 ( .AN(B[0]), .B(A[0]), .Y(n64) );
endmodule


module butterfly ( calc_in, rotation, calc_out );
  input [135:0] calc_in;
  input [2:0] rotation;
  output [135:0] calc_out;
  wire   n128, n129, n130, n131, n132, n133, n134, N9, N42, n7, n13, N306,
         N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295,
         N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284,
         N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273,
         N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228,
         N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217,
         N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206,
         N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195,
         N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184,
         N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173,
         N172, N171, N136, N135, N134, N133, N132, N131, N130, N129, N128,
         N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117,
         N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106,
         N105, N104, N103, N340, N339, N338, N337, N336, N335, N334, N333,
         N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322,
         N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311,
         N310, N309, N308, N307, N272, N271, N270, N269, N268, N267, N266,
         N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255,
         N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244,
         N243, N242, N241, N240, N239, N170, N169, N168, N167, N166, N165,
         N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154,
         N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143,
         N142, N141, N140, N139, N138, N137, N99, N98, N97, N96, N95, N94, N93,
         N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79,
         N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N102, N101, N100,
         n8, n9, n10, n12, n14, n15, n16, n17, n18, n20, n21, n22, n23, n24,
         n25, n28, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103;
  wire   [16:0] temp_2_1_real;
  wire   [16:0] temp_2_2_real;
  wire   [16:0] temp_2_1_imag;
  wire   [16:0] temp_2_2_imag;
  wire   [16:0] temp_3_1_real;
  wire   [16:0] temp_3_2_real;
  wire   [16:0] temp_3_1_imag;
  wire   [16:0] temp_3_2_imag;
  wire   [16:0] temp_4_1_real;
  wire   [16:0] temp_4_2_real;
  wire   [16:0] temp_4_1_imag;
  wire   [16:0] temp_4_2_imag;
  wire   [16:0] temp_1_real;
  wire   [16:0] temp_1_imag;
  wire   [16:0] temp_2_real;
  wire   [16:0] temp_2_imag;
  wire   [16:0] temp_3_real;
  wire   [16:0] temp_3_imag;

  multi16_11 multiBRR ( .in_17bit({calc_in[67:53], n49, n66}), .in_8bit({1'b0, 
        n36, n82, 1'b1, n80, n73, n76, n38}), .out(temp_2_1_real) );
  multi16_10 multiBII ( .in_17bit({calc_in[50:38], n33, calc_in[36:34]}), 
        .in_8bit({n91, n52, n37, 1'b0, n8, n79, n91, n103}), .out(
        temp_2_2_real) );
  multi16_9 multiBRI ( .in_17bit({calc_in[67:53], n49, n66}), .in_8bit({n91, 
        n53, n100, 1'b0, n98, n95, n91, n52}), .out(temp_2_1_imag) );
  multi16_8 multiBIR ( .in_17bit({calc_in[50:38], n33, calc_in[36:34]}), 
        .in_8bit({1'b0, n36, n82, 1'b1, n34, n73, n76, n93}), .out(
        temp_2_2_imag) );
  multi16_7 multiCRR ( .in_17bit(calc_in[101:85]), .in_8bit({n101, n74, n39, 
        n75, n75, n39, n63, N42}), .out(temp_3_1_real) );
  multi16_6 multiCII ( .in_17bit({calc_in[84:71], n54, n44, n60}), .in_8bit({
        n91, 1'b0, n98, 1'b0, 1'b0, n8, n98, n100}), .out(temp_3_2_real) );
  multi16_5 multiCRI ( .in_17bit(calc_in[101:85]), .in_8bit({n91, 1'b0, n8, 
        1'b0, 1'b0, n8, n98, n37}), .out(temp_3_1_imag) );
  multi16_4 multiCIR ( .in_17bit({calc_in[84:70], n44, n60}), .in_8bit({n101, 
        n75, n93, n73, n74, n38, n63, N42}), .out(temp_3_2_imag) );
  multi16_3 multiDRR ( .in_17bit({calc_in[135:123], n50, calc_in[121:119]}), 
        .in_8bit({n90, N42, n36, n74, n39, n35, n83, n74}), .out(temp_4_1_real) );
  multi16_2 multiDII ( .in_17bit({calc_in[118:106], n42, calc_in[104], n65, 
        n71}), .in_8bit({n95, 1'b0, n90, n101, n53, n100, n95, n102}), .out(
        temp_4_2_real) );
  multi16_1 multiDRI ( .in_17bit({calc_in[135:123], n50, calc_in[121:119]}), 
        .in_8bit({n94, 1'b0, n90, n101, n103, n37, n95, n9}), .out(
        temp_4_1_imag) );
  multi16_0 multiDIR ( .in_17bit({calc_in[118:106], n42, calc_in[104], n65, 
        n71}), .in_8bit({n89, N42, n76, n75, n93, n35, n83, n73}), .out(
        temp_4_2_imag) );
  butterfly_DW01_sub_25 sub_278 ( .A(temp_3_1_real), .B({temp_3_2_real[16:14], 
        n55, n62, temp_3_2_real[11:0]}), .DIFF(temp_2_real) );
  butterfly_DW01_add_18 add_0_root_add_0_root_add_292_3 ( .A({N102, N101, N100, 
        N99, N98, N97, N96, N95, N94, N93, N92, N91, n22, N89, N88, N87, N86}), 
        .B({N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, 
        N72, N71, N70, N69}), .SUM({calc_out[33:31], n131, calc_out[29:17]})
         );
  butterfly_DW01_add_20 add_0_root_sub_0_root_sub_296_2 ( .A({N204, N203, N202, 
        N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, 
        N189, N188}), .B({N187, N186, N185, N184, N183, N182, N181, N180, N179, 
        N178, N177, N176, N175, N174, N173, N172, N171}), .SUM(calc_out[84:68]) );
  butterfly_DW01_add_21 add_0_root_add_0_root_add_293_3 ( .A({N136, N135, N134, 
        N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, 
        N121, N120}), .B({N119, N118, N117, N116, N115, N114, N113, N112, N111, 
        N110, N109, N108, N107, N106, N105, N104, N103}), .SUM({calc_out[16], 
        n132, n133, n134, calc_out[12:0]}) );
  butterfly_DW01_sub_26 sub_1_root_sub_0_root_add_301 ( .A({n67, 
        temp_3_real[15:13], n72, temp_3_real[11:5], n18, temp_3_real[3:0]}), 
        .B({n68, temp_2_imag[15:9], n58, temp_2_imag[7:0]}), .DIFF({N323, N322, 
        N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, 
        N309, N308, N307}) );
  butterfly_DW01_sub_31 sub_1_root_sub_0_root_sub_299_2 ( .A(temp_1_real), .B(
        {n67, temp_3_real[15:13], n72, n46, temp_3_real[10:5], n18, 
        temp_3_real[3:0]}), .DIFF({N255, N254, N253, N252, N251, N250, N249, 
        N248, N247, N246, N245, N244, N243, N242, N241, N240, N239}) );
  butterfly_DW01_add_36 add_1_root_add_0_root_add_292_3 ( .A(temp_1_real), .B(
        {n67, temp_3_real[15:13], n72, temp_3_real[11:5], n18, 
        temp_3_real[3:0]}), .SUM({N85, N84, N83, N82, N81, N80, N79, N78, N77, 
        N76, N75, N74, N73, N72, N71, N70, N69}) );
  butterfly_DW01_add_44 add_0_root_sub_0_root_sub_299_2 ( .A({N272, N271, N270, 
        N269, N268, N267, N266, N265, N264, N263, n15, N261, N260, N259, N258, 
        N257, N256}), .B({N255, N254, N253, N252, N251, N250, N249, N248, N247, 
        N246, n28, N244, N243, N242, N241, N240, N239}), .SUM({
        calc_out[118:115], n128, calc_out[113:102]}) );
  butterfly_DW01_sub_35 sub_0_root_sub_0_root_sub_295_2 ( .A({N170, N169, N168, 
        N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, 
        N155, N154}), .B({N153, N152, N151, N150, N149, N148, N147, N146, N145, 
        N144, N143, N142, N141, N140, N139, N138, N137}), .DIFF({
        calc_out[101:96], n129, calc_out[94:85]}) );
  butterfly_DW01_add_49 add_282 ( .A(temp_4_1_imag), .B(temp_4_2_imag), .SUM(
        temp_3_imag) );
  butterfly_DW01_add_48 add_276 ( .A(temp_2_1_imag), .B(temp_2_2_imag), .SUM(
        temp_1_imag) );
  butterfly_DW01_add_50 add_279 ( .A(temp_3_1_imag), .B(temp_3_2_imag), .SUM(
        temp_2_imag) );
  butterfly_DW01_add_61 add_2_root_add_0_root_add_292_3 ( .A(calc_in[33:17]), 
        .B({n64, n69, temp_2_real[14:12], n43, temp_2_real[10:8], n51, n31, 
        temp_2_real[5:0]}), .SUM({N102, N101, N100, N99, N98, N97, N96, N95, 
        N94, N93, N92, N91, N90, N89, N88, N87, N86}) );
  butterfly_DW01_sub_57 sub_0_root_sub_0_root_sub_300_2 ( .A({N306, N305, N304, 
        N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, 
        N291, N290}), .B({N289, N288, N287, N286, N285, N284, n70, N282, N281, 
        N280, N279, N278, N277, N276, N275, N274, N273}), .DIFF({
        calc_out[67:61], n130, calc_out[59:51]}) );
  butterfly_DW01_add_77 add_2_root_sub_0_root_sub_295_2 ( .A(calc_in[33:17]), 
        .B({n64, n69, temp_2_real[14:12], n43, temp_2_real[10:8], n51, n31, 
        temp_2_real[5:0]}), .SUM({N170, N169, N168, N167, N166, N165, N164, 
        N163, N162, N161, N160, N159, N158, N157, N156, N155, N154}) );
  butterfly_DW01_add_73 add_0_root_sub_0_root_add_301 ( .A({N340, N339, N338, 
        N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, 
        N325, N324}), .B({N323, N322, N321, N320, N319, N318, N317, N316, N315, 
        N314, N313, N312, N311, N310, N309, N308, N307}), .SUM(calc_out[50:34]) );
  butterfly_DW01_sub_64 sub_2_root_sub_0_root_add_298 ( .A(calc_in[33:17]), 
        .B({n41, temp_1_imag[15:13], n92, temp_1_imag[11], n61, n24, n23, 
        temp_1_imag[7], n20, temp_1_imag[5:4], n16, temp_1_imag[2:0]}), .DIFF(
        {N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, 
        N227, N226, N225, N224, N223, N222}) );
  butterfly_DW01_add_85 add_2_root_sub_0_root_sub_300_2 ( .A(calc_in[33:17]), 
        .B({n41, temp_1_imag[15:13], n92, temp_1_imag[11], n61, temp_1_imag[9], 
        n23, temp_1_imag[7], n20, temp_1_imag[5:4], n16, temp_1_imag[2:0]}), 
        .SUM({N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, 
        N295, N294, N293, N292, N291, N290}) );
  butterfly_DW01_sub_69 sub_2_root_sub_0_root_sub_296_2 ( .A(calc_in[16:0]), 
        .B({n14, temp_1_imag[15:13], n92, temp_1_imag[11], n61, temp_1_imag[9], 
        n23, temp_1_imag[7], n20, temp_1_imag[5:4], n16, temp_1_imag[2:0]}), 
        .DIFF({N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, 
        N194, N193, N192, N191, N190, N189, N188}) );
  butterfly_DW01_sub_71 sub_281 ( .A({n48, temp_4_1_real[15:0]}), .B(
        temp_4_2_real), .DIFF(temp_3_real) );
  butterfly_DW01_add_90 add_1_root_add_0_root_add_293_3 ( .A({n41, 
        temp_1_imag[15:13], n92, temp_1_imag[11], n61, n24, n23, 
        temp_1_imag[7], n20, temp_1_imag[5:4], n16, temp_1_imag[2:0]}), .B({
        temp_3_imag[16:10], n17, temp_3_imag[8:6], n21, temp_3_imag[4:0]}), 
        .SUM({N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, 
        N108, N107, N106, N105, N104, N103}) );
  butterfly_DW01_sub_70 sub_2_root_sub_0_root_add_301 ( .A(calc_in[16:0]), .B(
        temp_1_real), .DIFF({N340, N339, N338, N337, N336, N335, N334, N333, 
        N332, N331, N330, N329, N328, N327, N326, N325, N324}) );
  butterfly_DW01_add_91 add_1_root_sub_0_root_sub_295_2 ( .A(temp_1_real), .B(
        {n67, temp_3_real[15:13], n72, temp_3_real[11:5], n18, 
        temp_3_real[3:0]}), .SUM({N153, N152, N151, N150, N149, N148, N147, 
        N146, N145, N144, N143, N142, N141, N140, N139, N138, N137}) );
  butterfly_DW01_add_98 add_1_root_sub_0_root_sub_300_2 ( .A({
        temp_3_imag[16:10], n17, temp_3_imag[8:6], n21, temp_3_imag[4:0]}), 
        .B({n64, n69, temp_2_real[14:12], n43, temp_2_real[10:8], n51, n31, 
        temp_2_real[5:0]}), .SUM({N289, N288, N287, N286, N285, N284, N283, 
        N282, N281, N280, N279, N278, N277, N276, N275, N274, N273}) );
  butterfly_DW01_sub_77 sub_2_root_sub_0_root_sub_299_2 ( .A(calc_in[16:0]), 
        .B({temp_2_imag[16:9], n58, temp_2_imag[7:0]}), .DIFF({N272, N271, 
        N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, 
        N258, N257, N256}) );
  butterfly_DW01_add_100 add_2_root_add_0_root_add_293_3 ( .A(calc_in[16:0]), 
        .B({n68, temp_2_imag[15:9], n58, temp_2_imag[7:0]}), .SUM({N136, N135, 
        N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, 
        N122, N121, N120}) );
  butterfly_DW01_sub_90 sub_275 ( .A(temp_2_1_real), .B(temp_2_2_real), .DIFF(
        temp_1_real) );
  butterfly_DW01_sub_81 sub_1_root_sub_0_root_sub_296_2 ( .A({n68, 
        temp_2_imag[15:9], n58, temp_2_imag[7:0]}), .B({temp_3_imag[16:10], 
        n17, temp_3_imag[8:6], n21, temp_3_imag[4:0]}), .DIFF({N187, N186, 
        N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, 
        N173, N172, N171}) );
  butterfly_DW01_add_104 add_0_root_sub_0_root_add_298 ( .A({N238, N237, N236, 
        N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, 
        N223, N222}), .B({N221, N220, N219, N218, N217, N216, N215, N214, N213, 
        N212, N211, N210, N209, N208, N207, N206, N205}), .SUM(
        calc_out[135:119]) );
  butterfly_DW01_sub_91 sub_1_root_sub_0_root_add_298 ( .A({temp_3_imag[16:10], 
        n17, temp_3_imag[8:6], n21, temp_3_imag[4:0]}), .B({n64, n69, 
        temp_2_real[14:12], n43, temp_2_real[10:8], n51, n31, temp_2_real[5:0]}), .DIFF({N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, 
        N210, N209, N208, N207, N206, N205}) );
  BUFX20 U9 ( .A(temp_1_imag[16]), .Y(n41) );
  BUFX20 U10 ( .A(temp_2_imag[16]), .Y(n68) );
  INVX20 U11 ( .A(n80), .Y(n8) );
  INVX2 U12 ( .A(temp_1_imag[16]), .Y(n12) );
  BUFX20 U13 ( .A(n102), .Y(n9) );
  CLKINVX8 U14 ( .A(n96), .Y(n102) );
  CLKINVX12 U15 ( .A(n97), .Y(n101) );
  AOI21X2 U16 ( .A0(n85), .A1(n86), .B0(n87), .Y(n10) );
  CLKBUFX8 U17 ( .A(calc_in[70]), .Y(n54) );
  BUFX12 U18 ( .A(n132), .Y(calc_out[15]) );
  INVX1 U19 ( .A(n78), .Y(n34) );
  INVX3 U20 ( .A(n78), .Y(n35) );
  INVX4 U21 ( .A(n12), .Y(n14) );
  BUFX4 U22 ( .A(N262), .Y(n15) );
  BUFX12 U23 ( .A(temp_1_imag[3]), .Y(n16) );
  BUFX20 U24 ( .A(n128), .Y(calc_out[114]) );
  BUFX16 U25 ( .A(temp_3_imag[9]), .Y(n17) );
  BUFX16 U26 ( .A(temp_3_real[4]), .Y(n18) );
  BUFX20 U27 ( .A(n133), .Y(calc_out[14]) );
  BUFX16 U28 ( .A(temp_1_imag[6]), .Y(n20) );
  BUFX20 U29 ( .A(N283), .Y(n70) );
  BUFX16 U30 ( .A(temp_3_imag[5]), .Y(n21) );
  BUFX8 U31 ( .A(N90), .Y(n22) );
  BUFX16 U32 ( .A(temp_1_imag[8]), .Y(n23) );
  BUFX8 U33 ( .A(temp_1_imag[9]), .Y(n24) );
  CLKINVX4 U34 ( .A(n130), .Y(n25) );
  INVX4 U35 ( .A(n25), .Y(calc_out[60]) );
  INVX8 U36 ( .A(n56), .Y(calc_out[95]) );
  BUFX8 U37 ( .A(N245), .Y(n28) );
  BUFX20 U38 ( .A(n134), .Y(calc_out[13]) );
  BUFX20 U39 ( .A(n131), .Y(calc_out[30]) );
  BUFX12 U40 ( .A(temp_2_real[6]), .Y(n31) );
  BUFX20 U41 ( .A(temp_2_imag[8]), .Y(n58) );
  CLKINVX8 U42 ( .A(n87), .Y(n32) );
  INVX8 U43 ( .A(rotation[2]), .Y(n87) );
  BUFX20 U44 ( .A(temp_3_2_real[12]), .Y(n62) );
  BUFX16 U45 ( .A(n97), .Y(n76) );
  BUFX20 U46 ( .A(temp_2_real[11]), .Y(n43) );
  BUFX12 U47 ( .A(calc_in[37]), .Y(n33) );
  CLKBUFX12 U48 ( .A(n84), .Y(n91) );
  INVX8 U49 ( .A(n7), .Y(n81) );
  INVX8 U50 ( .A(n81), .Y(n82) );
  INVX8 U51 ( .A(rotation[1]), .Y(n86) );
  INVX8 U52 ( .A(n78), .Y(n80) );
  OR2X2 U53 ( .A(n77), .B(n87), .Y(n47) );
  BUFX4 U54 ( .A(n97), .Y(n36) );
  INVX8 U55 ( .A(n82), .Y(n37) );
  INVX8 U56 ( .A(n94), .Y(n38) );
  INVX8 U57 ( .A(n94), .Y(n39) );
  BUFX16 U58 ( .A(calc_in[105]), .Y(n42) );
  BUFX20 U59 ( .A(calc_in[69]), .Y(n44) );
  AND2X4 U60 ( .A(rotation[0]), .B(rotation[2]), .Y(n40) );
  INVX8 U61 ( .A(n45), .Y(n46) );
  BUFX16 U62 ( .A(n13), .Y(n83) );
  INVX8 U63 ( .A(N9), .Y(n94) );
  BUFX20 U64 ( .A(calc_in[122]), .Y(n50) );
  BUFX20 U65 ( .A(temp_3_2_real[13]), .Y(n55) );
  NAND3X2 U66 ( .A(rotation[0]), .B(n59), .C(n32), .Y(n96) );
  BUFX8 U67 ( .A(temp_4_1_real[16]), .Y(n48) );
  BUFX20 U68 ( .A(temp_1_imag[10]), .Y(n61) );
  INVX8 U69 ( .A(temp_3_real[11]), .Y(n45) );
  INVX20 U70 ( .A(n47), .Y(n95) );
  INVX4 U71 ( .A(n86), .Y(n59) );
  INVX20 U72 ( .A(n10), .Y(N42) );
  CLKINVX4 U73 ( .A(n38), .Y(n79) );
  INVX12 U74 ( .A(n99), .Y(n90) );
  BUFX20 U75 ( .A(temp_2_real[7]), .Y(n51) );
  BUFX20 U76 ( .A(calc_in[51]), .Y(n66) );
  BUFX20 U77 ( .A(temp_3_real[16]), .Y(n67) );
  BUFX20 U78 ( .A(calc_in[52]), .Y(n49) );
  INVX3 U79 ( .A(rotation[0]), .Y(n85) );
  BUFX16 U80 ( .A(temp_2_real[16]), .Y(n64) );
  BUFX20 U81 ( .A(calc_in[103]), .Y(n65) );
  BUFX20 U82 ( .A(calc_in[68]), .Y(n60) );
  BUFX20 U83 ( .A(temp_2_real[15]), .Y(n69) );
  NAND3BX4 U84 ( .AN(rotation[0]), .B(rotation[1]), .C(rotation[2]), .Y(n7) );
  INVX8 U85 ( .A(n83), .Y(n52) );
  INVX8 U86 ( .A(n83), .Y(n53) );
  BUFX20 U87 ( .A(temp_3_real[12]), .Y(n72) );
  CLKINVX4 U88 ( .A(n129), .Y(n56) );
  BUFX20 U89 ( .A(n88), .Y(n74) );
  INVX8 U90 ( .A(n81), .Y(n63) );
  AND2X4 U91 ( .A(rotation[0]), .B(rotation[2]), .Y(n78) );
  BUFX20 U92 ( .A(calc_in[102]), .Y(n71) );
  BUFX20 U93 ( .A(temp_1_imag[12]), .Y(n92) );
  INVX20 U94 ( .A(n80), .Y(n98) );
  INVX8 U95 ( .A(n83), .Y(n103) );
  NAND3BX2 U96 ( .AN(rotation[1]), .B(rotation[2]), .C(rotation[0]), .Y(n13)
         );
  NAND2X4 U97 ( .A(n40), .B(n59), .Y(n97) );
  BUFX20 U98 ( .A(n88), .Y(n73) );
  INVX8 U99 ( .A(n82), .Y(n100) );
  NAND2BX4 U100 ( .AN(n77), .B(n32), .Y(N9) );
  NAND2X4 U101 ( .A(rotation[1]), .B(rotation[2]), .Y(n99) );
  INVX8 U102 ( .A(n94), .Y(n93) );
  CLKBUFX20 U103 ( .A(n88), .Y(n75) );
  INVX8 U104 ( .A(n89), .Y(n88) );
  XNOR2X4 U105 ( .A(rotation[0]), .B(rotation[1]), .Y(n77) );
  AOI21X4 U106 ( .A0(n85), .A1(n86), .B0(n87), .Y(n84) );
  CLKINVX8 U107 ( .A(n99), .Y(n89) );
endmodule


module reg1 ( clk, rst_n, data_in_2, reg_datain_flag, data_out_2 );
  input [135:0] data_in_2;
  output [135:0] data_out_2;
  input clk, rst_n, reg_datain_flag;
  wire   reg_flag_mux, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62,
         N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76,
         N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90,
         N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, N124, N125,
         N126, N127, N128, N129, N130, N131, N132, N133, N134, N135, N136,
         N137, N138, N139, N140, N141, N142, N143, N144, N145, N146, N147,
         N148, N149, N150, N151, N152, N153, N154, N155, N156, N157, N158,
         N159, N160, N161, N162, N163, N164, N165, N166, N167, N168, N169,
         N170, N171, N172, N173, N174, N175, N176, N177, N178, N179, N180,
         N181, N182, N183, N184, N185, N186, N187, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n961, n962, n963, n964, n965, n966, n968,
         n969, n971, n973, n974, n975, n976, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n7, n8, n9, n10, n45, n245, n317, n318, n614, n616,
         n618, n620, n622, n624, n626, n628, n630, n632, n634, n636, n638,
         n640, n642, n644, n646, n648, n650, n652, n654, n656, n658, n660,
         n662, n664, n666, n668, n670, n672, n674, n676, n678, n680, n682,
         n684, n958, n960, n970, n977, n1118, n1120, n1122, n1124, n1126,
         n1128, n1130, n1132, n1134, n1136, n1138, n1140, n1142, n1144, n1146,
         n1148, n1150, n1152, n1154, n1156, n1158, n1160, n1162, n1164, n1166,
         n1168, n1170, n1172, n1174, n1176, n1178, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250;
  wire   [1:0] counter1;
  wire   [33:0] R0;
  wire   [33:0] R1;
  wire   [33:0] R4;
  wire   [33:0] R5;
  wire   [33:0] R8;
  wire   [33:0] R9;
  wire   [33:0] R12;
  wire   [33:0] R13;
  wire   [1:0] counter2;

  EDFFX4 data_out_2_reg_130_ ( .D(N182), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[130]) );
  EDFFX4 data_out_2_reg_129_ ( .D(N181), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[129]) );
  EDFFX4 data_out_2_reg_128_ ( .D(N180), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[128]) );
  EDFFX4 data_out_2_reg_127_ ( .D(N179), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[127]) );
  EDFFX4 data_out_2_reg_126_ ( .D(N178), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[126]) );
  EDFFX4 data_out_2_reg_125_ ( .D(N177), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[125]) );
  EDFFX4 data_out_2_reg_120_ ( .D(N172), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[120]) );
  EDFFX4 data_out_2_reg_119_ ( .D(N171), .E(n1243), .CK(clk), .Q(
        data_out_2[119]) );
  EDFFX4 data_out_2_reg_118_ ( .D(N170), .E(n1243), .CK(clk), .Q(
        data_out_2[118]) );
  EDFFX4 data_out_2_reg_113_ ( .D(N165), .E(n1243), .CK(clk), .Q(
        data_out_2[113]) );
  EDFFX4 data_out_2_reg_111_ ( .D(N163), .E(n1244), .CK(clk), .Q(
        data_out_2[111]) );
  EDFFX4 data_out_2_reg_110_ ( .D(N162), .E(n1243), .CK(clk), .Q(
        data_out_2[110]) );
  EDFFX4 data_out_2_reg_109_ ( .D(N161), .E(n1244), .CK(clk), .Q(
        data_out_2[109]) );
  EDFFX4 data_out_2_reg_101_ ( .D(N153), .E(n1244), .CK(clk), .Q(
        data_out_2[101]) );
  EDFFX4 data_out_2_reg_84_ ( .D(N136), .E(n1243), .CK(clk), .Q(data_out_2[84]) );
  EDFFX4 data_out_2_reg_69_ ( .D(N121), .E(n1244), .CK(clk), .Q(data_out_2[69]) );
  EDFFX4 data_out_2_reg_68_ ( .D(N120), .E(n1243), .CK(clk), .Q(data_out_2[68]) );
  EDFFX4 data_out_2_reg_67_ ( .D(N119), .E(n1243), .CK(clk), .Q(data_out_2[67]) );
  EDFFX4 data_out_2_reg_63_ ( .D(N115), .E(n1244), .CK(clk), .Q(data_out_2[63]) );
  EDFFX4 data_out_2_reg_50_ ( .D(N102), .E(n1244), .CK(clk), .Q(data_out_2[50]) );
  CLKINVX4 U302 ( .A(rst_n), .Y(n961) );
  DFFXL R13_reg_30_ ( .D(n1180), .CK(clk), .Q(R13[30]) );
  DFFXL R9_reg_30_ ( .D(n1178), .CK(clk), .Q(R9[30]) );
  DFFXL R5_reg_30_ ( .D(n1176), .CK(clk), .Q(R5[30]) );
  DFFXL R1_reg_30_ ( .D(n1174), .CK(clk), .Q(R1[30]) );
  DFFXL R12_reg_12_ ( .D(n1172), .CK(clk), .Q(R12[12]) );
  DFFXL R8_reg_12_ ( .D(n1170), .CK(clk), .Q(R8[12]) );
  DFFXL R4_reg_12_ ( .D(n1168), .CK(clk), .Q(R4[12]) );
  DFFXL R0_reg_12_ ( .D(n1166), .CK(clk), .Q(R0[12]) );
  DFFXL R13_reg_12_ ( .D(n1164), .CK(clk), .Q(R13[12]) );
  DFFXL R9_reg_12_ ( .D(n1162), .CK(clk), .Q(R9[12]) );
  DFFXL R5_reg_12_ ( .D(n1160), .CK(clk), .Q(R5[12]) );
  DFFXL R1_reg_12_ ( .D(n1158), .CK(clk), .Q(R1[12]) );
  DFFXL R12_reg_13_ ( .D(n1156), .CK(clk), .Q(R12[13]) );
  DFFXL R8_reg_13_ ( .D(n1154), .CK(clk), .Q(R8[13]) );
  DFFXL R4_reg_13_ ( .D(n1152), .CK(clk), .Q(R4[13]) );
  DFFXL R0_reg_13_ ( .D(n1150), .CK(clk), .Q(R0[13]) );
  DFFXL R13_reg_13_ ( .D(n1148), .CK(clk), .Q(R13[13]) );
  DFFXL R9_reg_13_ ( .D(n1146), .CK(clk), .Q(R9[13]) );
  DFFXL R5_reg_13_ ( .D(n1144), .CK(clk), .Q(R5[13]) );
  DFFXL R1_reg_13_ ( .D(n1142), .CK(clk), .Q(R1[13]) );
  DFFXL R13_reg_31_ ( .D(n1140), .CK(clk), .Q(R13[31]) );
  DFFXL R9_reg_31_ ( .D(n1138), .CK(clk), .Q(R9[31]) );
  DFFXL R5_reg_31_ ( .D(n1136), .CK(clk), .Q(R5[31]) );
  DFFXL R1_reg_31_ ( .D(n1134), .CK(clk), .Q(R1[31]) );
  DFFXL R13_reg_14_ ( .D(n1132), .CK(clk), .Q(R13[14]) );
  DFFXL R9_reg_14_ ( .D(n1130), .CK(clk), .Q(R9[14]) );
  DFFXL R5_reg_14_ ( .D(n1128), .CK(clk), .Q(R5[14]) );
  DFFXL R1_reg_14_ ( .D(n1126), .CK(clk), .Q(R1[14]) );
  DFFXL R12_reg_30_ ( .D(n1124), .CK(clk), .Q(R12[30]) );
  DFFXL R8_reg_30_ ( .D(n1122), .CK(clk), .Q(R8[30]) );
  DFFXL R4_reg_30_ ( .D(n1120), .CK(clk), .Q(R4[30]) );
  DFFXL R0_reg_30_ ( .D(n1118), .CK(clk), .Q(R0[30]) );
  DFFXL R12_reg_16_ ( .D(n977), .CK(clk), .Q(R12[16]) );
  DFFXL R8_reg_16_ ( .D(n970), .CK(clk), .Q(R8[16]) );
  DFFXL R4_reg_16_ ( .D(n960), .CK(clk), .Q(R4[16]) );
  DFFXL R0_reg_16_ ( .D(n958), .CK(clk), .Q(R0[16]) );
  DFFXL R12_reg_31_ ( .D(n684), .CK(clk), .Q(R12[31]) );
  DFFXL R8_reg_31_ ( .D(n682), .CK(clk), .Q(R8[31]) );
  DFFXL R4_reg_31_ ( .D(n680), .CK(clk), .Q(R4[31]) );
  DFFXL R0_reg_31_ ( .D(n678), .CK(clk), .Q(R0[31]) );
  DFFXL R13_reg_16_ ( .D(n676), .CK(clk), .Q(R13[16]) );
  DFFXL R9_reg_16_ ( .D(n674), .CK(clk), .Q(R9[16]) );
  DFFXL R5_reg_16_ ( .D(n672), .CK(clk), .Q(R5[16]) );
  DFFXL R1_reg_16_ ( .D(n670), .CK(clk), .Q(R1[16]) );
  MX2X1 R12_reg_32__U3 ( .A(R12[32]), .B(data_in_2[32]), .S0(n1208), .Y(n668)
         );
  DFFXL R12_reg_32_ ( .D(n668), .CK(clk), .Q(R12[32]) );
  MX2X1 R8_reg_32__U3 ( .A(R8[32]), .B(data_in_2[32]), .S0(n1191), .Y(n666) );
  DFFXL R8_reg_32_ ( .D(n666), .CK(clk), .Q(R8[32]) );
  MX2X1 R4_reg_32__U3 ( .A(R4[32]), .B(data_in_2[32]), .S0(n1214), .Y(n664) );
  DFFXL R4_reg_32_ ( .D(n664), .CK(clk), .Q(R4[32]) );
  MX2X1 R0_reg_32__U3 ( .A(R0[32]), .B(data_in_2[32]), .S0(n1194), .Y(n662) );
  DFFXL R0_reg_32_ ( .D(n662), .CK(clk), .Q(R0[32]) );
  DFFXL R12_reg_33_ ( .D(n660), .CK(clk), .Q(R12[33]) );
  DFFXL R8_reg_33_ ( .D(n658), .CK(clk), .Q(R8[33]) );
  DFFXL R4_reg_33_ ( .D(n656), .CK(clk), .Q(R4[33]) );
  DFFXL R0_reg_33_ ( .D(n654), .CK(clk), .Q(R0[33]) );
  DFFXL R13_reg_32_ ( .D(n652), .CK(clk), .Q(R13[32]) );
  DFFXL R9_reg_32_ ( .D(n650), .CK(clk), .Q(R9[32]) );
  DFFXL R5_reg_32_ ( .D(n648), .CK(clk), .Q(R5[32]) );
  DFFXL R1_reg_32_ ( .D(n646), .CK(clk), .Q(R1[32]) );
  DFFXL R12_reg_14_ ( .D(n644), .CK(clk), .Q(R12[14]) );
  DFFXL R8_reg_14_ ( .D(n642), .CK(clk), .Q(R8[14]) );
  DFFXL R4_reg_14_ ( .D(n640), .CK(clk), .Q(R4[14]) );
  DFFXL R0_reg_14_ ( .D(n638), .CK(clk), .Q(R0[14]) );
  DFFXL R13_reg_33_ ( .D(n636), .CK(clk), .Q(R13[33]) );
  DFFXL R9_reg_33_ ( .D(n634), .CK(clk), .Q(R9[33]) );
  DFFXL R5_reg_33_ ( .D(n632), .CK(clk), .Q(R5[33]) );
  DFFXL R1_reg_33_ ( .D(n630), .CK(clk), .Q(R1[33]) );
  MX2X1 R12_reg_15__U3 ( .A(R12[15]), .B(data_in_2[15]), .S0(n1207), .Y(n628)
         );
  DFFXL R12_reg_15_ ( .D(n628), .CK(clk), .Q(R12[15]) );
  MX2X1 R8_reg_15__U3 ( .A(R8[15]), .B(data_in_2[15]), .S0(n1189), .Y(n626) );
  DFFXL R8_reg_15_ ( .D(n626), .CK(clk), .Q(R8[15]) );
  MX2X1 R4_reg_15__U3 ( .A(R4[15]), .B(data_in_2[15]), .S0(n1214), .Y(n624) );
  DFFXL R4_reg_15_ ( .D(n624), .CK(clk), .Q(R4[15]) );
  MX2X1 R0_reg_15__U3 ( .A(R0[15]), .B(data_in_2[15]), .S0(n1194), .Y(n622) );
  DFFXL R0_reg_15_ ( .D(n622), .CK(clk), .Q(R0[15]) );
  DFFXL R13_reg_15_ ( .D(n620), .CK(clk), .Q(R13[15]) );
  DFFXL R9_reg_15_ ( .D(n618), .CK(clk), .Q(R9[15]) );
  DFFXL R5_reg_15_ ( .D(n616), .CK(clk), .Q(R5[15]) );
  DFFXL R1_reg_15_ ( .D(n614), .CK(clk), .Q(R1[15]) );
  EDFFX1 R10_reg_24_ ( .D(data_in_2[92]), .E(n1186), .CK(clk), .QN(n729) );
  EDFFX1 R10_reg_23_ ( .D(data_in_2[91]), .E(n1191), .CK(clk), .QN(n730) );
  EDFFX1 R10_reg_22_ ( .D(data_in_2[90]), .E(n1189), .CK(clk), .QN(n731) );
  EDFFX1 R10_reg_21_ ( .D(data_in_2[89]), .E(n1187), .CK(clk), .QN(n732) );
  EDFFX1 R10_reg_20_ ( .D(data_in_2[88]), .E(n1191), .CK(clk), .QN(n733) );
  EDFFX1 R10_reg_19_ ( .D(data_in_2[87]), .E(n1188), .CK(clk), .QN(n734) );
  EDFFX1 R10_reg_7_ ( .D(data_in_2[75]), .E(n1187), .CK(clk), .QN(n746) );
  EDFFX1 R10_reg_6_ ( .D(data_in_2[74]), .E(n1187), .CK(clk), .QN(n747) );
  EDFFX1 R10_reg_5_ ( .D(data_in_2[73]), .E(n1187), .CK(clk), .QN(n748) );
  EDFFX1 R10_reg_4_ ( .D(data_in_2[72]), .E(n1187), .CK(clk), .QN(n749) );
  EDFFX1 R10_reg_3_ ( .D(data_in_2[71]), .E(n1187), .CK(clk), .QN(n750) );
  EDFFX1 R10_reg_2_ ( .D(data_in_2[70]), .E(n1187), .CK(clk), .QN(n751) );
  EDFFX1 R10_reg_1_ ( .D(data_in_2[69]), .E(n1186), .CK(clk), .QN(n752) );
  EDFFX1 R14_reg_24_ ( .D(data_in_2[92]), .E(n971), .CK(clk), .QN(n763) );
  EDFFX1 R14_reg_23_ ( .D(data_in_2[91]), .E(n971), .CK(clk), .QN(n764) );
  EDFFX1 R14_reg_22_ ( .D(data_in_2[90]), .E(n971), .CK(clk), .QN(n765) );
  EDFFX1 R14_reg_21_ ( .D(data_in_2[89]), .E(n971), .CK(clk), .QN(n766) );
  EDFFX1 R14_reg_20_ ( .D(data_in_2[88]), .E(n971), .CK(clk), .QN(n767) );
  EDFFX1 R14_reg_7_ ( .D(data_in_2[75]), .E(n1211), .CK(clk), .QN(n780) );
  EDFFX1 R14_reg_6_ ( .D(data_in_2[74]), .E(n1206), .CK(clk), .QN(n781) );
  EDFFX1 R14_reg_5_ ( .D(data_in_2[73]), .E(n1207), .CK(clk), .QN(n782) );
  EDFFX1 R14_reg_4_ ( .D(data_in_2[72]), .E(n1208), .CK(clk), .QN(n783) );
  EDFFX1 R14_reg_3_ ( .D(data_in_2[71]), .E(n1207), .CK(clk), .QN(n784) );
  EDFFX1 R14_reg_2_ ( .D(data_in_2[70]), .E(n1206), .CK(clk), .QN(n785) );
  EDFFX1 R14_reg_1_ ( .D(data_in_2[69]), .E(n971), .CK(clk), .QN(n786) );
  EDFFX1 R2_reg_24_ ( .D(data_in_2[92]), .E(n1196), .CK(clk), .QN(n831) );
  EDFFX1 R2_reg_23_ ( .D(data_in_2[91]), .E(n1196), .CK(clk), .QN(n832) );
  EDFFX1 R2_reg_22_ ( .D(data_in_2[90]), .E(n1196), .CK(clk), .QN(n833) );
  EDFFX1 R2_reg_21_ ( .D(data_in_2[89]), .E(n1196), .CK(clk), .QN(n834) );
  EDFFX1 R2_reg_20_ ( .D(data_in_2[88]), .E(n1196), .CK(clk), .QN(n835) );
  EDFFX1 R2_reg_19_ ( .D(data_in_2[87]), .E(n1196), .CK(clk), .QN(n836) );
  EDFFX1 R2_reg_7_ ( .D(data_in_2[75]), .E(n1195), .CK(clk), .QN(n848) );
  EDFFX1 R2_reg_6_ ( .D(data_in_2[74]), .E(n1195), .CK(clk), .QN(n849) );
  EDFFX1 R2_reg_5_ ( .D(data_in_2[73]), .E(n1195), .CK(clk), .QN(n850) );
  EDFFX1 R2_reg_4_ ( .D(data_in_2[72]), .E(n1194), .CK(clk), .QN(n851) );
  EDFFX1 R2_reg_3_ ( .D(data_in_2[71]), .E(n1194), .CK(clk), .QN(n852) );
  EDFFX1 R2_reg_2_ ( .D(data_in_2[70]), .E(n1195), .CK(clk), .QN(n853) );
  EDFFX1 R2_reg_1_ ( .D(data_in_2[69]), .E(n1194), .CK(clk), .QN(n854) );
  EDFFXL R6_reg_28_ ( .D(data_in_2[96]), .E(n1216), .CK(clk), .QN(n895) );
  EDFFXL R6_reg_27_ ( .D(data_in_2[95]), .E(n969), .CK(clk), .QN(n896) );
  EDFFXL R6_reg_26_ ( .D(data_in_2[94]), .E(n1214), .CK(clk), .QN(n897) );
  EDFFXL R6_reg_25_ ( .D(data_in_2[93]), .E(n1216), .CK(clk), .QN(n898) );
  EDFFXL R6_reg_24_ ( .D(data_in_2[92]), .E(n969), .CK(clk), .QN(n899) );
  EDFFXL R6_reg_23_ ( .D(data_in_2[91]), .E(n1214), .CK(clk), .QN(n900) );
  EDFFXL R6_reg_22_ ( .D(data_in_2[90]), .E(n1214), .CK(clk), .QN(n901) );
  EDFFXL R6_reg_21_ ( .D(data_in_2[89]), .E(n1216), .CK(clk), .QN(n902) );
  EDFFXL R6_reg_20_ ( .D(data_in_2[88]), .E(n1216), .CK(clk), .QN(n903) );
  EDFFXL R6_reg_19_ ( .D(data_in_2[87]), .E(n1214), .CK(clk), .QN(n904) );
  EDFFXL R6_reg_18_ ( .D(data_in_2[86]), .E(n969), .CK(clk), .QN(n905) );
  EDFFXL R6_reg_11_ ( .D(data_in_2[79]), .E(n969), .CK(clk), .QN(n912) );
  EDFFXL R6_reg_10_ ( .D(data_in_2[78]), .E(n1216), .CK(clk), .QN(n913) );
  EDFFXL R6_reg_9_ ( .D(data_in_2[77]), .E(n969), .CK(clk), .QN(n914) );
  EDFFXL R6_reg_8_ ( .D(data_in_2[76]), .E(n1215), .CK(clk), .QN(n915) );
  EDFFXL R6_reg_7_ ( .D(data_in_2[75]), .E(n1216), .CK(clk), .QN(n916) );
  EDFFXL R6_reg_6_ ( .D(data_in_2[74]), .E(n969), .CK(clk), .QN(n917) );
  EDFFXL R6_reg_5_ ( .D(data_in_2[73]), .E(n969), .CK(clk), .QN(n918) );
  EDFFXL R6_reg_4_ ( .D(data_in_2[72]), .E(n1215), .CK(clk), .QN(n919) );
  EDFFXL R6_reg_3_ ( .D(data_in_2[71]), .E(n1216), .CK(clk), .QN(n920) );
  EDFFXL R6_reg_2_ ( .D(data_in_2[70]), .E(n969), .CK(clk), .QN(n921) );
  EDFFXL R6_reg_1_ ( .D(data_in_2[69]), .E(n969), .CK(clk), .QN(n922) );
  EDFFX1 R11_reg_26_ ( .D(data_in_2[128]), .E(n1188), .CK(clk), .QN(n693) );
  EDFFX1 R11_reg_23_ ( .D(data_in_2[125]), .E(n1188), .CK(clk), .QN(n696) );
  EDFFX1 R11_reg_22_ ( .D(data_in_2[124]), .E(n1188), .CK(clk), .QN(n697) );
  EDFFX1 R11_reg_21_ ( .D(data_in_2[123]), .E(n1188), .CK(clk), .QN(n698) );
  EDFFX1 R11_reg_20_ ( .D(data_in_2[122]), .E(n1188), .CK(clk), .QN(n699) );
  EDFFX1 R11_reg_19_ ( .D(data_in_2[121]), .E(n1188), .CK(clk), .QN(n700) );
  EDFFX1 R11_reg_7_ ( .D(data_in_2[109]), .E(n317), .CK(clk), .QN(n712) );
  EDFFX1 R11_reg_6_ ( .D(data_in_2[108]), .E(n1187), .CK(clk), .QN(n713) );
  EDFFX1 R11_reg_5_ ( .D(data_in_2[107]), .E(n1188), .CK(clk), .QN(n714) );
  EDFFX1 R11_reg_4_ ( .D(data_in_2[106]), .E(n1191), .CK(clk), .QN(n715) );
  EDFFX1 R11_reg_3_ ( .D(data_in_2[105]), .E(n1191), .CK(clk), .QN(n716) );
  EDFFX1 R11_reg_2_ ( .D(data_in_2[104]), .E(n1191), .CK(clk), .QN(n717) );
  EDFFX1 R15_reg_26_ ( .D(data_in_2[128]), .E(n1211), .CK(clk), .QN(n795) );
  EDFFX1 R15_reg_23_ ( .D(data_in_2[125]), .E(n1211), .CK(clk), .QN(n798) );
  EDFFX1 R15_reg_22_ ( .D(data_in_2[124]), .E(n1206), .CK(clk), .QN(n799) );
  EDFFX1 R15_reg_21_ ( .D(data_in_2[123]), .E(n1206), .CK(clk), .QN(n800) );
  EDFFX1 R15_reg_20_ ( .D(data_in_2[122]), .E(n1211), .CK(clk), .QN(n801) );
  EDFFX1 R15_reg_19_ ( .D(data_in_2[121]), .E(n1211), .CK(clk), .QN(n802) );
  EDFFX1 R15_reg_7_ ( .D(data_in_2[109]), .E(n1206), .CK(clk), .QN(n814) );
  EDFFX1 R15_reg_6_ ( .D(data_in_2[108]), .E(n1206), .CK(clk), .QN(n815) );
  EDFFX1 R15_reg_5_ ( .D(data_in_2[107]), .E(n1206), .CK(clk), .QN(n816) );
  EDFFX1 R15_reg_4_ ( .D(data_in_2[106]), .E(n1206), .CK(clk), .QN(n817) );
  EDFFX1 R15_reg_3_ ( .D(data_in_2[105]), .E(n1206), .CK(clk), .QN(n818) );
  EDFFX1 R15_reg_2_ ( .D(data_in_2[104]), .E(n1206), .CK(clk), .QN(n819) );
  EDFFX1 R3_reg_26_ ( .D(data_in_2[128]), .E(n1194), .CK(clk), .QN(n863) );
  EDFFX1 R3_reg_23_ ( .D(data_in_2[125]), .E(n1195), .CK(clk), .QN(n866) );
  EDFFX1 R3_reg_22_ ( .D(data_in_2[124]), .E(n1195), .CK(clk), .QN(n867) );
  EDFFX1 R3_reg_21_ ( .D(data_in_2[123]), .E(n1194), .CK(clk), .QN(n868) );
  EDFFX1 R3_reg_20_ ( .D(data_in_2[122]), .E(n1194), .CK(clk), .QN(n869) );
  EDFFX1 R3_reg_19_ ( .D(data_in_2[121]), .E(n1195), .CK(clk), .QN(n870) );
  EDFFX1 R3_reg_7_ ( .D(data_in_2[109]), .E(n1194), .CK(clk), .QN(n882) );
  EDFFX1 R3_reg_6_ ( .D(data_in_2[108]), .E(n1195), .CK(clk), .QN(n883) );
  EDFFX1 R3_reg_5_ ( .D(data_in_2[107]), .E(n1194), .CK(clk), .QN(n884) );
  EDFFX1 R3_reg_4_ ( .D(data_in_2[106]), .E(n1196), .CK(clk), .QN(n885) );
  EDFFX1 R3_reg_3_ ( .D(data_in_2[105]), .E(n1194), .CK(clk), .QN(n886) );
  EDFFX1 R3_reg_2_ ( .D(data_in_2[104]), .E(n1194), .CK(clk), .QN(n887) );
  EDFFXL R7_reg_29_ ( .D(data_in_2[131]), .E(n1216), .CK(clk), .QN(n928) );
  EDFFXL R7_reg_28_ ( .D(data_in_2[130]), .E(n1214), .CK(clk), .QN(n929) );
  EDFFXL R7_reg_27_ ( .D(data_in_2[129]), .E(n1215), .CK(clk), .QN(n930) );
  EDFFXL R7_reg_26_ ( .D(data_in_2[128]), .E(n1216), .CK(clk), .QN(n931) );
  EDFFXL R7_reg_25_ ( .D(data_in_2[127]), .E(n1214), .CK(clk), .QN(n932) );
  EDFFXL R7_reg_24_ ( .D(data_in_2[126]), .E(n1215), .CK(clk), .QN(n933) );
  EDFFXL R7_reg_23_ ( .D(data_in_2[125]), .E(n1216), .CK(clk), .QN(n934) );
  EDFFXL R7_reg_22_ ( .D(data_in_2[124]), .E(n969), .CK(clk), .QN(n935) );
  EDFFXL R7_reg_21_ ( .D(data_in_2[123]), .E(n969), .CK(clk), .QN(n936) );
  EDFFXL R7_reg_20_ ( .D(data_in_2[122]), .E(n969), .CK(clk), .QN(n937) );
  EDFFXL R7_reg_19_ ( .D(data_in_2[121]), .E(n969), .CK(clk), .QN(n938) );
  EDFFXL R7_reg_18_ ( .D(data_in_2[120]), .E(n969), .CK(clk), .QN(n939) );
  EDFFXL R7_reg_11_ ( .D(data_in_2[113]), .E(n969), .CK(clk), .QN(n946) );
  EDFFXL R7_reg_10_ ( .D(data_in_2[112]), .E(n1215), .CK(clk), .QN(n947) );
  EDFFXL R7_reg_9_ ( .D(data_in_2[111]), .E(n1216), .CK(clk), .QN(n948) );
  EDFFXL R7_reg_8_ ( .D(data_in_2[110]), .E(n1215), .CK(clk), .QN(n949) );
  EDFFXL R7_reg_7_ ( .D(data_in_2[109]), .E(n1216), .CK(clk), .QN(n950) );
  EDFFXL R7_reg_6_ ( .D(data_in_2[108]), .E(n1216), .CK(clk), .QN(n951) );
  EDFFXL R7_reg_5_ ( .D(data_in_2[107]), .E(n1215), .CK(clk), .QN(n952) );
  EDFFXL R7_reg_4_ ( .D(data_in_2[106]), .E(n1216), .CK(clk), .QN(n953) );
  EDFFXL R7_reg_3_ ( .D(data_in_2[105]), .E(n1215), .CK(clk), .QN(n954) );
  EDFFXL R7_reg_2_ ( .D(data_in_2[104]), .E(n1215), .CK(clk), .QN(n955) );
  EDFFXL R7_reg_1_ ( .D(data_in_2[103]), .E(n1215), .CK(clk), .QN(n956) );
  EDFFX1 R8_reg_22_ ( .D(data_in_2[22]), .E(n1190), .CK(clk), .Q(R8[22]) );
  EDFFX1 R8_reg_21_ ( .D(data_in_2[21]), .E(n1190), .CK(clk), .Q(R8[21]) );
  EDFFX1 R8_reg_20_ ( .D(data_in_2[20]), .E(n1190), .CK(clk), .Q(R8[20]) );
  EDFFX1 R8_reg_19_ ( .D(data_in_2[19]), .E(n1190), .CK(clk), .Q(R8[19]) );
  EDFFX1 R8_reg_18_ ( .D(data_in_2[18]), .E(n1190), .CK(clk), .Q(R8[18]) );
  EDFFX1 R8_reg_7_ ( .D(data_in_2[7]), .E(n1189), .CK(clk), .Q(R8[7]) );
  EDFFX1 R8_reg_6_ ( .D(data_in_2[6]), .E(n1189), .CK(clk), .Q(R8[6]) );
  EDFFX1 R8_reg_4_ ( .D(data_in_2[4]), .E(n1187), .CK(clk), .Q(R8[4]) );
  EDFFX1 R8_reg_3_ ( .D(data_in_2[3]), .E(n1188), .CK(clk), .Q(R8[3]) );
  EDFFX1 R8_reg_2_ ( .D(data_in_2[2]), .E(n1186), .CK(clk), .Q(R8[2]) );
  EDFFX1 R8_reg_1_ ( .D(data_in_2[1]), .E(n1188), .CK(clk), .Q(R8[1]) );
  EDFFX1 R8_reg_0_ ( .D(data_in_2[0]), .E(n1191), .CK(clk), .Q(R8[0]) );
  EDFFX1 R12_reg_22_ ( .D(data_in_2[22]), .E(n1209), .CK(clk), .Q(R12[22]) );
  EDFFX1 R12_reg_21_ ( .D(data_in_2[21]), .E(n1208), .CK(clk), .Q(R12[21]) );
  EDFFX1 R12_reg_20_ ( .D(data_in_2[20]), .E(n1211), .CK(clk), .Q(R12[20]) );
  EDFFX1 R12_reg_19_ ( .D(data_in_2[19]), .E(n1209), .CK(clk), .Q(R12[19]) );
  EDFFX1 R12_reg_18_ ( .D(data_in_2[18]), .E(n1208), .CK(clk), .Q(R12[18]) );
  EDFFX1 R12_reg_7_ ( .D(data_in_2[7]), .E(n1207), .CK(clk), .Q(R12[7]) );
  EDFFX1 R12_reg_6_ ( .D(data_in_2[6]), .E(n1207), .CK(clk), .Q(R12[6]) );
  EDFFX1 R12_reg_4_ ( .D(data_in_2[4]), .E(n1207), .CK(clk), .Q(R12[4]) );
  EDFFX1 R12_reg_3_ ( .D(data_in_2[3]), .E(n1207), .CK(clk), .Q(R12[3]) );
  EDFFX1 R12_reg_2_ ( .D(data_in_2[2]), .E(n1211), .CK(clk), .Q(R12[2]) );
  EDFFX1 R12_reg_1_ ( .D(data_in_2[1]), .E(n1211), .CK(clk), .Q(R12[1]) );
  EDFFX1 R12_reg_0_ ( .D(data_in_2[0]), .E(n1208), .CK(clk), .Q(R12[0]) );
  EDFFX1 R0_reg_22_ ( .D(data_in_2[22]), .E(n1194), .CK(clk), .Q(R0[22]) );
  EDFFX1 R0_reg_21_ ( .D(data_in_2[21]), .E(n1194), .CK(clk), .Q(R0[21]) );
  EDFFX1 R0_reg_20_ ( .D(data_in_2[20]), .E(n1194), .CK(clk), .Q(R0[20]) );
  EDFFX1 R0_reg_19_ ( .D(data_in_2[19]), .E(n1194), .CK(clk), .Q(R0[19]) );
  EDFFX1 R0_reg_18_ ( .D(data_in_2[18]), .E(n1194), .CK(clk), .Q(R0[18]) );
  EDFFX1 R0_reg_7_ ( .D(data_in_2[7]), .E(n1194), .CK(clk), .Q(R0[7]) );
  EDFFX1 R0_reg_6_ ( .D(data_in_2[6]), .E(n1195), .CK(clk), .Q(R0[6]) );
  EDFFX1 R0_reg_4_ ( .D(data_in_2[4]), .E(n1195), .CK(clk), .Q(R0[4]) );
  EDFFX1 R0_reg_3_ ( .D(data_in_2[3]), .E(n1194), .CK(clk), .Q(R0[3]) );
  EDFFX1 R0_reg_2_ ( .D(data_in_2[2]), .E(n1195), .CK(clk), .Q(R0[2]) );
  EDFFX1 R0_reg_1_ ( .D(data_in_2[1]), .E(n1195), .CK(clk), .Q(R0[1]) );
  EDFFX1 R0_reg_0_ ( .D(data_in_2[0]), .E(n1195), .CK(clk), .Q(R0[0]) );
  EDFFXL R4_reg_28_ ( .D(data_in_2[28]), .E(n1214), .CK(clk), .Q(R4[28]) );
  EDFFXL R4_reg_27_ ( .D(data_in_2[27]), .E(n1214), .CK(clk), .Q(R4[27]) );
  EDFFXL R4_reg_26_ ( .D(data_in_2[26]), .E(n1214), .CK(clk), .Q(R4[26]) );
  EDFFXL R4_reg_25_ ( .D(data_in_2[25]), .E(n1214), .CK(clk), .Q(R4[25]) );
  EDFFXL R4_reg_24_ ( .D(data_in_2[24]), .E(n1214), .CK(clk), .Q(R4[24]) );
  EDFFXL R4_reg_23_ ( .D(data_in_2[23]), .E(n1214), .CK(clk), .Q(R4[23]) );
  EDFFXL R4_reg_22_ ( .D(data_in_2[22]), .E(n1214), .CK(clk), .Q(R4[22]) );
  EDFFXL R4_reg_21_ ( .D(data_in_2[21]), .E(n1214), .CK(clk), .Q(R4[21]) );
  EDFFXL R4_reg_20_ ( .D(data_in_2[20]), .E(n1214), .CK(clk), .Q(R4[20]) );
  EDFFXL R4_reg_19_ ( .D(data_in_2[19]), .E(n1214), .CK(clk), .Q(R4[19]) );
  EDFFXL R4_reg_18_ ( .D(data_in_2[18]), .E(n1214), .CK(clk), .Q(R4[18]) );
  EDFFXL R4_reg_11_ ( .D(data_in_2[11]), .E(n1215), .CK(clk), .Q(R4[11]) );
  EDFFXL R4_reg_10_ ( .D(data_in_2[10]), .E(n1215), .CK(clk), .Q(R4[10]) );
  EDFFXL R4_reg_9_ ( .D(data_in_2[9]), .E(n1215), .CK(clk), .Q(R4[9]) );
  EDFFXL R4_reg_8_ ( .D(data_in_2[8]), .E(n1215), .CK(clk), .Q(R4[8]) );
  EDFFXL R4_reg_7_ ( .D(data_in_2[7]), .E(n1215), .CK(clk), .Q(R4[7]) );
  EDFFXL R4_reg_5_ ( .D(data_in_2[5]), .E(n1215), .CK(clk), .Q(R4[5]) );
  EDFFXL R4_reg_4_ ( .D(data_in_2[4]), .E(n1215), .CK(clk), .Q(R4[4]) );
  EDFFXL R4_reg_3_ ( .D(data_in_2[3]), .E(n1215), .CK(clk), .Q(R4[3]) );
  EDFFXL R4_reg_2_ ( .D(data_in_2[2]), .E(n1215), .CK(clk), .Q(R4[2]) );
  EDFFXL R4_reg_1_ ( .D(data_in_2[1]), .E(n1215), .CK(clk), .Q(R4[1]) );
  EDFFX1 R4_reg_0_ ( .D(data_in_2[0]), .E(n1215), .CK(clk), .Q(R4[0]) );
  EDFFXL R13_reg_29_ ( .D(data_in_2[63]), .E(n1210), .CK(clk), .Q(R13[29]) );
  EDFFXL R13_reg_28_ ( .D(data_in_2[62]), .E(n1210), .CK(clk), .Q(R13[28]) );
  EDFFXL R13_reg_27_ ( .D(data_in_2[61]), .E(n1210), .CK(clk), .Q(R13[27]) );
  EDFFXL R13_reg_26_ ( .D(data_in_2[60]), .E(n1210), .CK(clk), .Q(R13[26]) );
  EDFFXL R13_reg_25_ ( .D(data_in_2[59]), .E(n1210), .CK(clk), .Q(R13[25]) );
  EDFFXL R13_reg_24_ ( .D(data_in_2[58]), .E(n1210), .CK(clk), .Q(R13[24]) );
  EDFFXL R13_reg_23_ ( .D(data_in_2[57]), .E(n1210), .CK(clk), .Q(R13[23]) );
  EDFFXL R13_reg_22_ ( .D(data_in_2[56]), .E(n1210), .CK(clk), .Q(R13[22]) );
  EDFFXL R13_reg_21_ ( .D(data_in_2[55]), .E(n1210), .CK(clk), .Q(R13[21]) );
  EDFFXL R13_reg_20_ ( .D(data_in_2[54]), .E(n1210), .CK(clk), .Q(R13[20]) );
  EDFFXL R13_reg_11_ ( .D(data_in_2[45]), .E(n1209), .CK(clk), .Q(R13[11]) );
  EDFFXL R13_reg_10_ ( .D(data_in_2[44]), .E(n1209), .CK(clk), .Q(R13[10]) );
  EDFFXL R13_reg_9_ ( .D(data_in_2[43]), .E(n1209), .CK(clk), .Q(R13[9]) );
  EDFFXL R13_reg_8_ ( .D(data_in_2[42]), .E(n1209), .CK(clk), .Q(R13[8]) );
  EDFFXL R13_reg_7_ ( .D(data_in_2[41]), .E(n1209), .CK(clk), .Q(R13[7]) );
  EDFFXL R13_reg_6_ ( .D(data_in_2[40]), .E(n1209), .CK(clk), .Q(R13[6]) );
  EDFFXL R13_reg_5_ ( .D(data_in_2[39]), .E(n1208), .CK(clk), .Q(R13[5]) );
  EDFFXL R13_reg_4_ ( .D(data_in_2[38]), .E(n1208), .CK(clk), .Q(R13[4]) );
  EDFFXL R13_reg_3_ ( .D(data_in_2[37]), .E(n1208), .CK(clk), .Q(R13[3]) );
  EDFFXL R13_reg_2_ ( .D(data_in_2[36]), .E(n1208), .CK(clk), .Q(R13[2]) );
  EDFFXL R9_reg_29_ ( .D(data_in_2[63]), .E(n1186), .CK(clk), .Q(R9[29]) );
  EDFFXL R9_reg_28_ ( .D(data_in_2[62]), .E(n1186), .CK(clk), .Q(R9[28]) );
  EDFFXL R9_reg_27_ ( .D(data_in_2[61]), .E(n1186), .CK(clk), .Q(R9[27]) );
  EDFFXL R9_reg_26_ ( .D(data_in_2[60]), .E(n1186), .CK(clk), .Q(R9[26]) );
  EDFFXL R9_reg_25_ ( .D(data_in_2[59]), .E(n1186), .CK(clk), .Q(R9[25]) );
  EDFFXL R9_reg_24_ ( .D(data_in_2[58]), .E(n1186), .CK(clk), .Q(R9[24]) );
  EDFFXL R9_reg_23_ ( .D(data_in_2[57]), .E(n317), .CK(clk), .Q(R9[23]) );
  EDFFXL R9_reg_22_ ( .D(data_in_2[56]), .E(n317), .CK(clk), .Q(R9[22]) );
  EDFFXL R9_reg_21_ ( .D(data_in_2[55]), .E(n317), .CK(clk), .Q(R9[21]) );
  EDFFXL R9_reg_20_ ( .D(data_in_2[54]), .E(n317), .CK(clk), .Q(R9[20]) );
  EDFFXL R9_reg_11_ ( .D(data_in_2[45]), .E(n1185), .CK(clk), .Q(R9[11]) );
  EDFFXL R9_reg_10_ ( .D(data_in_2[44]), .E(n1185), .CK(clk), .Q(R9[10]) );
  EDFFXL R9_reg_9_ ( .D(data_in_2[43]), .E(n1185), .CK(clk), .Q(R9[9]) );
  EDFFXL R9_reg_8_ ( .D(data_in_2[42]), .E(n1185), .CK(clk), .Q(R9[8]) );
  EDFFXL R9_reg_7_ ( .D(data_in_2[41]), .E(n1185), .CK(clk), .Q(R9[7]) );
  EDFFXL R9_reg_6_ ( .D(data_in_2[40]), .E(n1185), .CK(clk), .Q(R9[6]) );
  EDFFXL R9_reg_5_ ( .D(data_in_2[39]), .E(n1185), .CK(clk), .Q(R9[5]) );
  EDFFXL R9_reg_4_ ( .D(data_in_2[38]), .E(n1185), .CK(clk), .Q(R9[4]) );
  EDFFXL R9_reg_3_ ( .D(data_in_2[37]), .E(n1185), .CK(clk), .Q(R9[3]) );
  EDFFXL R9_reg_2_ ( .D(data_in_2[36]), .E(n1185), .CK(clk), .Q(R9[2]) );
  EDFFXL R1_reg_29_ ( .D(data_in_2[63]), .E(n1195), .CK(clk), .Q(R1[29]) );
  EDFFXL R1_reg_28_ ( .D(data_in_2[62]), .E(n1194), .CK(clk), .Q(R1[28]) );
  EDFFXL R1_reg_27_ ( .D(data_in_2[61]), .E(n1194), .CK(clk), .Q(R1[27]) );
  EDFFXL R1_reg_26_ ( .D(data_in_2[60]), .E(n1195), .CK(clk), .Q(R1[26]) );
  EDFFXL R1_reg_25_ ( .D(data_in_2[59]), .E(n1195), .CK(clk), .Q(R1[25]) );
  EDFFXL R1_reg_24_ ( .D(data_in_2[58]), .E(n1195), .CK(clk), .Q(R1[24]) );
  EDFFXL R1_reg_23_ ( .D(data_in_2[57]), .E(n1195), .CK(clk), .Q(R1[23]) );
  EDFFXL R1_reg_22_ ( .D(data_in_2[56]), .E(n1195), .CK(clk), .Q(R1[22]) );
  EDFFXL R1_reg_21_ ( .D(data_in_2[55]), .E(n1195), .CK(clk), .Q(R1[21]) );
  EDFFXL R1_reg_20_ ( .D(data_in_2[54]), .E(n1195), .CK(clk), .Q(R1[20]) );
  EDFFXL R1_reg_11_ ( .D(data_in_2[45]), .E(n1195), .CK(clk), .Q(R1[11]) );
  EDFFXL R1_reg_10_ ( .D(data_in_2[44]), .E(n1195), .CK(clk), .Q(R1[10]) );
  EDFFXL R1_reg_9_ ( .D(data_in_2[43]), .E(n1195), .CK(clk), .Q(R1[9]) );
  EDFFXL R1_reg_8_ ( .D(data_in_2[42]), .E(n1195), .CK(clk), .Q(R1[8]) );
  EDFFXL R1_reg_7_ ( .D(data_in_2[41]), .E(n1195), .CK(clk), .Q(R1[7]) );
  EDFFXL R1_reg_6_ ( .D(data_in_2[40]), .E(n1195), .CK(clk), .Q(R1[6]) );
  EDFFXL R1_reg_5_ ( .D(data_in_2[39]), .E(n1195), .CK(clk), .Q(R1[5]) );
  EDFFXL R1_reg_4_ ( .D(data_in_2[38]), .E(n1195), .CK(clk), .Q(R1[4]) );
  EDFFXL R1_reg_3_ ( .D(data_in_2[37]), .E(n1196), .CK(clk), .Q(R1[3]) );
  EDFFXL R1_reg_2_ ( .D(data_in_2[36]), .E(n1196), .CK(clk), .Q(R1[2]) );
  EDFFXL R5_reg_29_ ( .D(data_in_2[63]), .E(n1215), .CK(clk), .Q(R5[29]) );
  EDFFXL R5_reg_28_ ( .D(data_in_2[62]), .E(n1215), .CK(clk), .Q(R5[28]) );
  EDFFXL R5_reg_27_ ( .D(data_in_2[61]), .E(n1215), .CK(clk), .Q(R5[27]) );
  EDFFXL R5_reg_26_ ( .D(data_in_2[60]), .E(n1216), .CK(clk), .Q(R5[26]) );
  EDFFXL R5_reg_25_ ( .D(data_in_2[59]), .E(n1216), .CK(clk), .Q(R5[25]) );
  EDFFXL R5_reg_24_ ( .D(data_in_2[58]), .E(n1216), .CK(clk), .Q(R5[24]) );
  EDFFXL R5_reg_23_ ( .D(data_in_2[57]), .E(n1216), .CK(clk), .Q(R5[23]) );
  EDFFXL R5_reg_22_ ( .D(data_in_2[56]), .E(n1216), .CK(clk), .Q(R5[22]) );
  EDFFXL R5_reg_21_ ( .D(data_in_2[55]), .E(n1216), .CK(clk), .Q(R5[21]) );
  EDFFXL R5_reg_20_ ( .D(data_in_2[54]), .E(n1216), .CK(clk), .Q(R5[20]) );
  EDFFXL R5_reg_11_ ( .D(data_in_2[45]), .E(n1216), .CK(clk), .Q(R5[11]) );
  EDFFXL R5_reg_10_ ( .D(data_in_2[44]), .E(n1216), .CK(clk), .Q(R5[10]) );
  EDFFXL R5_reg_9_ ( .D(data_in_2[43]), .E(n1216), .CK(clk), .Q(R5[9]) );
  EDFFXL R5_reg_8_ ( .D(data_in_2[42]), .E(n1216), .CK(clk), .Q(R5[8]) );
  EDFFXL R5_reg_7_ ( .D(data_in_2[41]), .E(n1216), .CK(clk), .Q(R5[7]) );
  EDFFXL R5_reg_6_ ( .D(data_in_2[40]), .E(n1216), .CK(clk), .Q(R5[6]) );
  EDFFXL R5_reg_5_ ( .D(data_in_2[39]), .E(n1216), .CK(clk), .Q(R5[5]) );
  EDFFXL R5_reg_4_ ( .D(data_in_2[38]), .E(n1214), .CK(clk), .Q(R5[4]) );
  EDFFXL R5_reg_3_ ( .D(data_in_2[37]), .E(n1215), .CK(clk), .Q(R5[3]) );
  EDFFXL R5_reg_2_ ( .D(data_in_2[36]), .E(n1216), .CK(clk), .Q(R5[2]) );
  DFFHQX1 counter1_reg_0_ ( .D(n1116), .CK(clk), .Q(counter1[0]) );
  DFFHQX1 counter1_reg_1_ ( .D(n1115), .CK(clk), .Q(counter1[1]) );
  DFFHQX1 counter2_reg_0_ ( .D(n1114), .CK(clk), .Q(counter2[0]) );
  DFFHQX1 counter2_reg_1_ ( .D(n1113), .CK(clk), .Q(counter2[1]) );
  EDFFX1 data_out_2_reg_81_ ( .D(N133), .E(n1243), .CK(clk), .Q(data_out_2[81]) );
  EDFFX1 data_out_2_reg_80_ ( .D(N132), .E(n1243), .CK(clk), .Q(data_out_2[80]) );
  EDFFX1 data_out_2_reg_79_ ( .D(N131), .E(n1243), .CK(clk), .Q(data_out_2[79]) );
  EDFFX1 data_out_2_reg_97_ ( .D(N149), .E(n1243), .CK(clk), .Q(data_out_2[97]) );
  EDFFX1 data_out_2_reg_98_ ( .D(N150), .E(n1243), .CK(clk), .Q(data_out_2[98]) );
  EDFFX1 data_out_2_reg_115_ ( .D(N167), .E(n1243), .CK(clk), .Q(
        data_out_2[115]) );
  EDFFX1 data_out_2_reg_46_ ( .D(N98), .E(n1244), .CK(clk), .Q(data_out_2[46])
         );
  EDFFX1 data_out_2_reg_96_ ( .D(N148), .E(n1243), .CK(clk), .Q(data_out_2[96]) );
  EDFFX1 data_out_2_reg_95_ ( .D(N147), .E(n1243), .CK(clk), .Q(data_out_2[95]) );
  EDFFX1 data_out_2_reg_47_ ( .D(N99), .E(n1244), .CK(clk), .Q(data_out_2[47])
         );
  EDFFX1 data_out_2_reg_78_ ( .D(N130), .E(n1244), .CK(clk), .Q(data_out_2[78]) );
  EDFFX1 data_out_2_reg_77_ ( .D(N129), .E(n1243), .CK(clk), .Q(data_out_2[77]) );
  EDFFX1 data_out_2_reg_93_ ( .D(N145), .E(n1243), .CK(clk), .Q(data_out_2[93]) );
  EDFFX1 data_out_2_reg_94_ ( .D(N146), .E(n1243), .CK(clk), .Q(data_out_2[94]) );
  EDFFX1 data_out_2_reg_75_ ( .D(N127), .E(n1243), .CK(clk), .Q(data_out_2[75]) );
  EDFFX1 data_out_2_reg_74_ ( .D(N126), .E(n1244), .CK(clk), .Q(data_out_2[74]) );
  EDFFX1 data_out_2_reg_90_ ( .D(N142), .E(n1243), .CK(clk), .Q(data_out_2[90]) );
  EDFFX1 data_out_2_reg_92_ ( .D(N144), .E(n1243), .CK(clk), .Q(data_out_2[92]) );
  EDFFX1 data_out_2_reg_36_ ( .D(N88), .E(n1244), .CK(clk), .Q(data_out_2[36])
         );
  EDFFX1 data_out_2_reg_72_ ( .D(N124), .E(n1243), .CK(clk), .Q(data_out_2[72]) );
  EDFFX1 data_out_2_reg_89_ ( .D(N141), .E(n1243), .CK(clk), .Q(data_out_2[89]) );
  EDFFX1 data_out_2_reg_37_ ( .D(N89), .E(n1244), .CK(clk), .Q(data_out_2[37])
         );
  EDFFX1 data_out_2_reg_55_ ( .D(N107), .E(n1244), .CK(clk), .Q(data_out_2[55]) );
  EDFFX1 data_out_2_reg_106_ ( .D(N158), .E(n1244), .CK(clk), .Q(
        data_out_2[106]) );
  EDFFX1 data_out_2_reg_38_ ( .D(N90), .E(n1244), .CK(clk), .Q(data_out_2[38])
         );
  EDFFX1 data_out_2_reg_123_ ( .D(N175), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[123]) );
  EDFFX1 data_out_2_reg_104_ ( .D(N156), .E(n1243), .CK(clk), .Q(
        data_out_2[104]) );
  EDFFX1 data_out_2_reg_52_ ( .D(N104), .E(n1244), .CK(clk), .Q(data_out_2[52]) );
  EDFFX1 data_out_2_reg_86_ ( .D(N138), .E(n1243), .CK(clk), .Q(data_out_2[86]) );
  EDFFX1 data_out_2_reg_103_ ( .D(N155), .E(n1243), .CK(clk), .Q(
        data_out_2[103]) );
  EDFFX1 data_out_2_reg_85_ ( .D(N137), .E(n1243), .CK(clk), .Q(data_out_2[85]) );
  EDFFX1 data_out_2_reg_35_ ( .D(N87), .E(n1244), .CK(clk), .Q(data_out_2[35])
         );
  EDFFX1 data_out_2_reg_87_ ( .D(N139), .E(n1243), .CK(clk), .Q(data_out_2[87]) );
  EDFFX1 data_out_2_reg_70_ ( .D(N122), .E(n1244), .CK(clk), .Q(data_out_2[70]) );
  EDFFX1 data_out_2_reg_53_ ( .D(N105), .E(n1244), .CK(clk), .Q(data_out_2[53]) );
  EDFFX1 data_out_2_reg_121_ ( .D(N173), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[121]) );
  EDFFX1 data_out_2_reg_135_ ( .D(N187), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[135]) );
  EDFFX1 data_out_2_reg_114_ ( .D(N166), .E(n1244), .CK(clk), .Q(
        data_out_2[114]) );
  EDFFX1 data_out_2_reg_45_ ( .D(N97), .E(n1244), .CK(clk), .Q(data_out_2[45])
         );
  EDFFX1 data_out_2_reg_60_ ( .D(N112), .E(n1244), .CK(clk), .Q(data_out_2[60]) );
  EDFFX1 data_out_2_reg_107_ ( .D(N159), .E(n1243), .CK(clk), .Q(
        data_out_2[107]) );
  EDFFX1 data_out_2_reg_39_ ( .D(N91), .E(n1243), .CK(clk), .Q(data_out_2[39])
         );
  EDFFX1 data_out_2_reg_56_ ( .D(N108), .E(n1244), .CK(clk), .Q(data_out_2[56]) );
  EDFFX2 data_out_2_reg_122_ ( .D(N174), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[122]) );
  EDFFX2 data_out_2_reg_54_ ( .D(N106), .E(n1244), .CK(clk), .Q(data_out_2[54]) );
  EDFFX2 data_out_2_reg_91_ ( .D(N143), .E(n1243), .CK(clk), .Q(data_out_2[91]) );
  EDFFX2 data_out_2_reg_71_ ( .D(N123), .E(n1244), .CK(clk), .Q(data_out_2[71]) );
  EDFFX2 data_out_2_reg_51_ ( .D(N103), .E(n1244), .CK(clk), .Q(data_out_2[51]) );
  EDFFX2 data_out_2_reg_34_ ( .D(N86), .E(n1244), .CK(clk), .Q(data_out_2[34])
         );
  EDFFX2 data_out_2_reg_102_ ( .D(N154), .E(n1243), .CK(clk), .Q(
        data_out_2[102]) );
  EDFFX2 data_out_2_reg_88_ ( .D(N140), .E(n1243), .CK(clk), .Q(data_out_2[88]) );
  EDFFX1 data_out_2_reg_132_ ( .D(N184), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[132]) );
  EDFFX1 data_out_2_reg_58_ ( .D(N110), .E(n1244), .CK(clk), .Q(data_out_2[58]) );
  EDFFX1 data_out_2_reg_73_ ( .D(N125), .E(n1243), .CK(clk), .Q(data_out_2[73]) );
  EDFFX1 data_out_2_reg_57_ ( .D(N109), .E(n1244), .CK(clk), .Q(data_out_2[57]) );
  EDFFX1 data_out_2_reg_65_ ( .D(N117), .E(n1244), .CK(clk), .Q(data_out_2[65]) );
  EDFFX1 data_out_2_reg_64_ ( .D(N116), .E(n1243), .CK(clk), .Q(data_out_2[64]) );
  EDFFX1 data_out_2_reg_44_ ( .D(N96), .E(n1244), .CK(clk), .Q(data_out_2[44])
         );
  EDFFX1 data_out_2_reg_43_ ( .D(N95), .E(n1244), .CK(clk), .Q(data_out_2[43])
         );
  EDFFX1 data_out_2_reg_42_ ( .D(N94), .E(n1244), .CK(clk), .Q(data_out_2[42])
         );
  EDFFX1 data_out_2_reg_59_ ( .D(N111), .E(n1244), .CK(clk), .Q(data_out_2[59]) );
  EDFFX1 data_out_2_reg_124_ ( .D(N176), .E(n1244), .CK(clk), .Q(
        data_out_2[124]) );
  EDFFX1 data_out_2_reg_108_ ( .D(N160), .E(n1244), .CK(clk), .Q(
        data_out_2[108]) );
  EDFFX1 data_out_2_reg_40_ ( .D(N92), .E(n1244), .CK(clk), .Q(data_out_2[40])
         );
  EDFFX1 data_out_2_reg_105_ ( .D(N157), .E(n1243), .CK(clk), .Q(
        data_out_2[105]) );
  EDFFXL R8_reg_25_ ( .D(data_in_2[25]), .E(n1190), .CK(clk), .Q(R8[25]) );
  EDFFXL R12_reg_25_ ( .D(data_in_2[25]), .E(n971), .CK(clk), .Q(R12[25]) );
  EDFFXL R0_reg_25_ ( .D(data_in_2[25]), .E(n1194), .CK(clk), .Q(R0[25]) );
  EDFFXL R8_reg_26_ ( .D(data_in_2[26]), .E(n1190), .CK(clk), .Q(R8[26]) );
  EDFFXL R12_reg_26_ ( .D(data_in_2[26]), .E(n1209), .CK(clk), .Q(R12[26]) );
  EDFFXL R0_reg_26_ ( .D(data_in_2[26]), .E(n1194), .CK(clk), .Q(R0[26]) );
  EDFFXL R8_reg_28_ ( .D(data_in_2[28]), .E(n1190), .CK(clk), .Q(R8[28]) );
  EDFFXL R12_reg_28_ ( .D(data_in_2[28]), .E(n1208), .CK(clk), .Q(R12[28]) );
  EDFFXL R0_reg_28_ ( .D(data_in_2[28]), .E(n1194), .CK(clk), .Q(R0[28]) );
  EDFFXL R10_reg_9_ ( .D(data_in_2[77]), .E(n1187), .CK(clk), .QN(n744) );
  EDFFXL R14_reg_9_ ( .D(data_in_2[77]), .E(n1209), .CK(clk), .QN(n778) );
  EDFFXL R2_reg_9_ ( .D(data_in_2[77]), .E(n1194), .CK(clk), .QN(n846) );
  EDFFXL R2_reg_27_ ( .D(data_in_2[95]), .E(n1196), .CK(clk), .QN(n828) );
  EDFFXL R14_reg_27_ ( .D(data_in_2[95]), .E(n1210), .CK(clk), .QN(n760) );
  EDFFXL R10_reg_27_ ( .D(data_in_2[95]), .E(n1191), .CK(clk), .QN(n726) );
  EDFFXL R10_reg_8_ ( .D(data_in_2[76]), .E(n1187), .CK(clk), .QN(n745) );
  EDFFXL R14_reg_8_ ( .D(data_in_2[76]), .E(n1210), .CK(clk), .QN(n779) );
  EDFFXL R2_reg_8_ ( .D(data_in_2[76]), .E(n1195), .CK(clk), .QN(n847) );
  EDFFXL R11_reg_11_ ( .D(data_in_2[113]), .E(n317), .CK(clk), .QN(n708) );
  EDFFXL R15_reg_11_ ( .D(data_in_2[113]), .E(n1206), .CK(clk), .QN(n810) );
  EDFFXL R3_reg_11_ ( .D(data_in_2[113]), .E(n1196), .CK(clk), .QN(n878) );
  EDFFXL R8_reg_8_ ( .D(data_in_2[8]), .E(n1189), .CK(clk), .Q(R8[8]) );
  EDFFXL R12_reg_8_ ( .D(data_in_2[8]), .E(n1207), .CK(clk), .Q(R12[8]) );
  EDFFXL R0_reg_8_ ( .D(data_in_2[8]), .E(n318), .CK(clk), .Q(R0[8]) );
  EDFFXL R8_reg_24_ ( .D(data_in_2[24]), .E(n1190), .CK(clk), .Q(R8[24]) );
  EDFFXL R12_reg_24_ ( .D(data_in_2[24]), .E(n1208), .CK(clk), .Q(R12[24]) );
  EDFFXL R0_reg_24_ ( .D(data_in_2[24]), .E(n1194), .CK(clk), .Q(R0[24]) );
  EDFFX1 R4_reg_6_ ( .D(data_in_2[6]), .E(n1215), .CK(clk), .Q(R4[6]) );
  EDFFXL R8_reg_11_ ( .D(data_in_2[11]), .E(n1189), .CK(clk), .Q(R8[11]) );
  EDFFXL R12_reg_11_ ( .D(data_in_2[11]), .E(n1207), .CK(clk), .Q(R12[11]) );
  EDFFXL R0_reg_11_ ( .D(data_in_2[11]), .E(n1194), .CK(clk), .Q(R0[11]) );
  EDFFXL R11_reg_8_ ( .D(data_in_2[110]), .E(n317), .CK(clk), .QN(n711) );
  EDFFXL R15_reg_8_ ( .D(data_in_2[110]), .E(n1206), .CK(clk), .QN(n813) );
  EDFFXL R3_reg_8_ ( .D(data_in_2[110]), .E(n1195), .CK(clk), .QN(n881) );
  EDFFXL R8_reg_27_ ( .D(data_in_2[27]), .E(n1190), .CK(clk), .Q(R8[27]) );
  EDFFXL R12_reg_27_ ( .D(data_in_2[27]), .E(n1211), .CK(clk), .Q(R12[27]) );
  EDFFXL R0_reg_27_ ( .D(data_in_2[27]), .E(n1194), .CK(clk), .Q(R0[27]) );
  EDFFXL R14_reg_26_ ( .D(data_in_2[94]), .E(n1210), .CK(clk), .QN(n761) );
  EDFFXL R2_reg_26_ ( .D(data_in_2[94]), .E(n1196), .CK(clk), .QN(n829) );
  EDFFXL R10_reg_26_ ( .D(data_in_2[94]), .E(n1185), .CK(clk), .QN(n727) );
  EDFFXL R11_reg_9_ ( .D(data_in_2[111]), .E(n317), .CK(clk), .QN(n710) );
  EDFFXL R15_reg_9_ ( .D(data_in_2[111]), .E(n1206), .CK(clk), .QN(n812) );
  EDFFXL R3_reg_9_ ( .D(data_in_2[111]), .E(n1194), .CK(clk), .QN(n880) );
  EDFFXL R8_reg_23_ ( .D(data_in_2[23]), .E(n1190), .CK(clk), .Q(R8[23]) );
  EDFFXL R12_reg_23_ ( .D(data_in_2[23]), .E(n1210), .CK(clk), .Q(R12[23]) );
  EDFFXL R0_reg_23_ ( .D(data_in_2[23]), .E(n1194), .CK(clk), .Q(R0[23]) );
  EDFFXL data_out_2_reg_49_ ( .D(N101), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[49]) );
  EDFFXL data_out_2_reg_48_ ( .D(N100), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[48]) );
  EDFFXL data_out_2_reg_134_ ( .D(N186), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[134]) );
  EDFFXL data_out_2_reg_133_ ( .D(N185), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[133]) );
  EDFFXL data_out_2_reg_117_ ( .D(N169), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[117]) );
  EDFFXL data_out_2_reg_116_ ( .D(N168), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[116]) );
  EDFFXL data_out_2_reg_100_ ( .D(N152), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[100]) );
  EDFFXL data_out_2_reg_99_ ( .D(N151), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[99]) );
  EDFFXL data_out_2_reg_83_ ( .D(N135), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[83]) );
  EDFFXL data_out_2_reg_82_ ( .D(N134), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[82]) );
  EDFFXL data_out_2_reg_33_ ( .D(N85), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[33]) );
  EDFFXL data_out_2_reg_32_ ( .D(N84), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[32]) );
  EDFFXL data_out_2_reg_31_ ( .D(N83), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[31]) );
  EDFFXL data_out_2_reg_30_ ( .D(N82), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[30]) );
  EDFFXL data_out_2_reg_29_ ( .D(N81), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[29]) );
  EDFFXL data_out_2_reg_28_ ( .D(N80), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[28]) );
  EDFFXL data_out_2_reg_27_ ( .D(N79), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[27]) );
  EDFFXL data_out_2_reg_26_ ( .D(N78), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[26]) );
  EDFFXL data_out_2_reg_25_ ( .D(N77), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[25]) );
  EDFFXL data_out_2_reg_24_ ( .D(N76), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[24]) );
  EDFFXL data_out_2_reg_23_ ( .D(N75), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[23]) );
  EDFFXL data_out_2_reg_22_ ( .D(N74), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[22]) );
  EDFFXL data_out_2_reg_21_ ( .D(N73), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[21]) );
  EDFFXL data_out_2_reg_20_ ( .D(N72), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[20]) );
  EDFFXL data_out_2_reg_19_ ( .D(N71), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[19]) );
  EDFFXL data_out_2_reg_18_ ( .D(N70), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[18]) );
  EDFFXL data_out_2_reg_17_ ( .D(N69), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[17]) );
  EDFFXL data_out_2_reg_16_ ( .D(N68), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[16]) );
  EDFFXL data_out_2_reg_15_ ( .D(N67), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[15]) );
  EDFFXL data_out_2_reg_14_ ( .D(N66), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[14]) );
  EDFFXL data_out_2_reg_13_ ( .D(N65), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[13]) );
  EDFFXL data_out_2_reg_12_ ( .D(N64), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[12]) );
  EDFFXL data_out_2_reg_11_ ( .D(N63), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[11]) );
  EDFFXL data_out_2_reg_10_ ( .D(N62), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[10]) );
  EDFFXL data_out_2_reg_9_ ( .D(N61), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[9]) );
  EDFFXL data_out_2_reg_8_ ( .D(N60), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[8]) );
  EDFFXL data_out_2_reg_7_ ( .D(N59), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[7]) );
  EDFFXL data_out_2_reg_6_ ( .D(N58), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[6]) );
  EDFFXL data_out_2_reg_5_ ( .D(N57), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[5]) );
  EDFFXL data_out_2_reg_4_ ( .D(N56), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[4]) );
  EDFFXL data_out_2_reg_3_ ( .D(N55), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[3]) );
  EDFFXL data_out_2_reg_2_ ( .D(N54), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[2]) );
  EDFFXL data_out_2_reg_1_ ( .D(N53), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[1]) );
  EDFFXL data_out_2_reg_0_ ( .D(N52), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[0]) );
  EDFFXL data_out_2_reg_66_ ( .D(N118), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[66]) );
  EDFFXL R13_reg_17_ ( .D(data_in_2[51]), .E(n971), .CK(clk), .Q(R13[17]) );
  EDFFXL R9_reg_17_ ( .D(data_in_2[51]), .E(n317), .CK(clk), .Q(R9[17]) );
  EDFFXL R5_reg_17_ ( .D(data_in_2[51]), .E(n969), .CK(clk), .Q(R5[17]) );
  EDFFXL R1_reg_17_ ( .D(data_in_2[51]), .E(n318), .CK(clk), .Q(R1[17]) );
  EDFFXL R12_reg_17_ ( .D(data_in_2[17]), .E(n971), .CK(clk), .Q(R12[17]) );
  EDFFXL R8_reg_17_ ( .D(data_in_2[17]), .E(n317), .CK(clk), .Q(R8[17]) );
  EDFFXL R4_reg_17_ ( .D(data_in_2[17]), .E(n969), .CK(clk), .Q(R4[17]) );
  EDFFXL R0_reg_17_ ( .D(data_in_2[17]), .E(n318), .CK(clk), .Q(R0[17]) );
  EDFFXL R13_reg_0_ ( .D(data_in_2[34]), .E(n971), .CK(clk), .Q(R13[0]) );
  EDFFXL R9_reg_0_ ( .D(data_in_2[34]), .E(n317), .CK(clk), .Q(R9[0]) );
  EDFFXL R5_reg_0_ ( .D(data_in_2[34]), .E(n969), .CK(clk), .Q(R5[0]) );
  EDFFXL R1_reg_0_ ( .D(data_in_2[34]), .E(n318), .CK(clk), .Q(R1[0]) );
  EDFFXL data_out_2_reg_41_ ( .D(N93), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[41]) );
  EDFFXL data_out_2_reg_61_ ( .D(N113), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[61]) );
  EDFFXL data_out_2_reg_76_ ( .D(N128), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[76]) );
  EDFFXL data_out_2_reg_131_ ( .D(N183), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[131]) );
  EDFFXL data_out_2_reg_112_ ( .D(N164), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[112]) );
  EDFFXL data_out_2_reg_62_ ( .D(N114), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[62]) );
  EDFFXL R13_reg_1_ ( .D(data_in_2[35]), .E(n971), .CK(clk), .Q(R13[1]) );
  EDFFXL R9_reg_1_ ( .D(data_in_2[35]), .E(n317), .CK(clk), .Q(R9[1]) );
  EDFFXL R5_reg_1_ ( .D(data_in_2[35]), .E(n969), .CK(clk), .Q(R5[1]) );
  EDFFXL R1_reg_1_ ( .D(data_in_2[35]), .E(n318), .CK(clk), .Q(R1[1]) );
  EDFFXL R13_reg_18_ ( .D(data_in_2[52]), .E(n971), .CK(clk), .Q(R13[18]) );
  EDFFXL R9_reg_18_ ( .D(data_in_2[52]), .E(n317), .CK(clk), .Q(R9[18]) );
  EDFFXL R5_reg_18_ ( .D(data_in_2[52]), .E(n969), .CK(clk), .Q(R5[18]) );
  EDFFXL R1_reg_18_ ( .D(data_in_2[52]), .E(n318), .CK(clk), .Q(R1[18]) );
  EDFFXL R13_reg_19_ ( .D(data_in_2[53]), .E(n971), .CK(clk), .Q(R13[19]) );
  EDFFXL R9_reg_19_ ( .D(data_in_2[53]), .E(n317), .CK(clk), .Q(R9[19]) );
  EDFFXL R5_reg_19_ ( .D(data_in_2[53]), .E(n969), .CK(clk), .Q(R5[19]) );
  EDFFXL R1_reg_19_ ( .D(data_in_2[53]), .E(n318), .CK(clk), .Q(R1[19]) );
  EDFFXL R15_reg_17_ ( .D(data_in_2[119]), .E(n971), .CK(clk), .QN(n804) );
  EDFFXL R11_reg_17_ ( .D(data_in_2[119]), .E(n317), .CK(clk), .QN(n702) );
  EDFFXL R7_reg_17_ ( .D(data_in_2[119]), .E(n969), .CK(clk), .QN(n940) );
  EDFFXL R3_reg_17_ ( .D(data_in_2[119]), .E(n318), .CK(clk), .QN(n872) );
  EDFFXL R14_reg_0_ ( .D(data_in_2[68]), .E(n971), .CK(clk), .QN(n787) );
  EDFFXL R10_reg_0_ ( .D(data_in_2[68]), .E(n317), .CK(clk), .QN(n753) );
  EDFFXL R6_reg_0_ ( .D(data_in_2[68]), .E(n969), .CK(clk), .QN(n923) );
  EDFFXL R2_reg_0_ ( .D(data_in_2[68]), .E(n318), .CK(clk), .QN(n855) );
  EDFFXL R14_reg_17_ ( .D(data_in_2[85]), .E(n971), .CK(clk), .QN(n770) );
  EDFFXL R10_reg_17_ ( .D(data_in_2[85]), .E(n317), .CK(clk), .QN(n736) );
  EDFFXL R6_reg_17_ ( .D(data_in_2[85]), .E(n969), .CK(clk), .QN(n906) );
  EDFFXL R2_reg_17_ ( .D(data_in_2[85]), .E(n318), .CK(clk), .QN(n838) );
  EDFFXL R15_reg_0_ ( .D(data_in_2[102]), .E(n971), .CK(clk), .QN(n821) );
  EDFFXL R11_reg_0_ ( .D(data_in_2[102]), .E(n317), .CK(clk), .QN(n719) );
  EDFFXL R7_reg_0_ ( .D(data_in_2[102]), .E(n969), .CK(clk), .QN(n957) );
  EDFFXL R3_reg_0_ ( .D(data_in_2[102]), .E(n318), .CK(clk), .QN(n889) );
  EDFFXL R14_reg_18_ ( .D(data_in_2[86]), .E(n971), .CK(clk), .QN(n769) );
  EDFFXL R10_reg_18_ ( .D(data_in_2[86]), .E(n317), .CK(clk), .QN(n735) );
  EDFFXL R2_reg_18_ ( .D(data_in_2[86]), .E(n318), .CK(clk), .QN(n837) );
  EDFFXL R15_reg_1_ ( .D(data_in_2[103]), .E(n971), .CK(clk), .QN(n820) );
  EDFFXL R11_reg_1_ ( .D(data_in_2[103]), .E(n317), .CK(clk), .QN(n718) );
  EDFFXL R3_reg_1_ ( .D(data_in_2[103]), .E(n318), .CK(clk), .QN(n888) );
  EDFFXL R15_reg_18_ ( .D(data_in_2[120]), .E(n971), .CK(clk), .QN(n803) );
  EDFFXL R11_reg_18_ ( .D(data_in_2[120]), .E(n317), .CK(clk), .QN(n701) );
  EDFFXL R3_reg_18_ ( .D(data_in_2[120]), .E(n318), .CK(clk), .QN(n871) );
  EDFFXL R14_reg_19_ ( .D(data_in_2[87]), .E(n1206), .CK(clk), .QN(n768) );
  DFFHQXL R0_reg_29_ ( .D(n1181), .CK(clk), .Q(R0[29]) );
  DFFHQXL R4_reg_29_ ( .D(n1182), .CK(clk), .Q(R4[29]) );
  DFFHQXL R8_reg_29_ ( .D(n1183), .CK(clk), .Q(R8[29]) );
  DFFHQXL R12_reg_29_ ( .D(n1184), .CK(clk), .Q(R12[29]) );
  EDFFXL R7_reg_12_ ( .D(data_in_2[114]), .E(n969), .CK(clk), .QN(n945) );
  EDFFXL R3_reg_12_ ( .D(data_in_2[114]), .E(n318), .CK(clk), .QN(n877) );
  EDFFXL R15_reg_12_ ( .D(data_in_2[114]), .E(n971), .CK(clk), .QN(n809) );
  EDFFXL R11_reg_12_ ( .D(data_in_2[114]), .E(n317), .CK(clk), .QN(n707) );
  EDFFXL R7_reg_30_ ( .D(data_in_2[132]), .E(n969), .CK(clk), .QN(n927) );
  EDFFXL R3_reg_30_ ( .D(data_in_2[132]), .E(n318), .CK(clk), .QN(n859) );
  EDFFXL R15_reg_30_ ( .D(data_in_2[132]), .E(n971), .CK(clk), .QN(n791) );
  EDFFXL R11_reg_30_ ( .D(data_in_2[132]), .E(n317), .CK(clk), .QN(n689) );
  EDFFXL R6_reg_29_ ( .D(data_in_2[97]), .E(n969), .CK(clk), .QN(n894) );
  EDFFXL R2_reg_29_ ( .D(data_in_2[97]), .E(n318), .CK(clk), .QN(n826) );
  EDFFXL R14_reg_29_ ( .D(data_in_2[97]), .E(n971), .CK(clk), .QN(n758) );
  EDFFXL R10_reg_29_ ( .D(data_in_2[97]), .E(n317), .CK(clk), .QN(n724) );
  EDFFXL R6_reg_13_ ( .D(data_in_2[81]), .E(n969), .CK(clk), .QN(n910) );
  EDFFXL R2_reg_13_ ( .D(data_in_2[81]), .E(n318), .CK(clk), .QN(n842) );
  EDFFXL R14_reg_13_ ( .D(data_in_2[81]), .E(n971), .CK(clk), .QN(n774) );
  EDFFXL R10_reg_13_ ( .D(data_in_2[81]), .E(n317), .CK(clk), .QN(n740) );
  EDFFXL R6_reg_12_ ( .D(data_in_2[80]), .E(n969), .CK(clk), .QN(n911) );
  EDFFXL R2_reg_12_ ( .D(data_in_2[80]), .E(n318), .CK(clk), .QN(n843) );
  EDFFXL R7_reg_13_ ( .D(data_in_2[115]), .E(n969), .CK(clk), .QN(n944) );
  EDFFXL R3_reg_13_ ( .D(data_in_2[115]), .E(n318), .CK(clk), .QN(n876) );
  EDFFXL R14_reg_12_ ( .D(data_in_2[80]), .E(n971), .CK(clk), .QN(n775) );
  EDFFXL R10_reg_12_ ( .D(data_in_2[80]), .E(n317), .CK(clk), .QN(n741) );
  EDFFXL R15_reg_13_ ( .D(data_in_2[115]), .E(n971), .CK(clk), .QN(n808) );
  EDFFXL R11_reg_13_ ( .D(data_in_2[115]), .E(n317), .CK(clk), .QN(n706) );
  EDFFXL R7_reg_31_ ( .D(data_in_2[133]), .E(n969), .CK(clk), .QN(n926) );
  EDFFXL R3_reg_31_ ( .D(data_in_2[133]), .E(n318), .CK(clk), .QN(n858) );
  EDFFXL R15_reg_31_ ( .D(data_in_2[133]), .E(n971), .CK(clk), .QN(n790) );
  EDFFXL R11_reg_31_ ( .D(data_in_2[133]), .E(n317), .CK(clk), .QN(n688) );
  EDFFXL R15_reg_32_ ( .D(data_in_2[134]), .E(n971), .CK(clk), .QN(n789) );
  EDFFXL R6_reg_30_ ( .D(data_in_2[98]), .E(n969), .CK(clk), .QN(n893) );
  EDFFXL R2_reg_30_ ( .D(data_in_2[98]), .E(n318), .CK(clk), .QN(n825) );
  EDFFXL R14_reg_30_ ( .D(data_in_2[98]), .E(n971), .CK(clk), .QN(n757) );
  EDFFXL R10_reg_30_ ( .D(data_in_2[98]), .E(n317), .CK(clk), .QN(n723) );
  EDFFXL R7_reg_14_ ( .D(data_in_2[116]), .E(n969), .CK(clk), .QN(n943) );
  EDFFXL R3_reg_14_ ( .D(data_in_2[116]), .E(n318), .CK(clk), .QN(n875) );
  EDFFXL R15_reg_14_ ( .D(data_in_2[116]), .E(n971), .CK(clk), .QN(n807) );
  EDFFXL R11_reg_14_ ( .D(data_in_2[116]), .E(n317), .CK(clk), .QN(n705) );
  EDFFXL R6_reg_31_ ( .D(data_in_2[99]), .E(n969), .CK(clk), .QN(n892) );
  EDFFXL R2_reg_31_ ( .D(data_in_2[99]), .E(n318), .CK(clk), .QN(n824) );
  EDFFXL R14_reg_31_ ( .D(data_in_2[99]), .E(n971), .CK(clk), .QN(n756) );
  EDFFXL R10_reg_31_ ( .D(data_in_2[99]), .E(n317), .CK(clk), .QN(n722) );
  EDFFXL R7_reg_32_ ( .D(data_in_2[134]), .E(n969), .CK(clk), .QN(n925) );
  EDFFXL R3_reg_32_ ( .D(data_in_2[134]), .E(n318), .CK(clk), .QN(n857) );
  EDFFXL R11_reg_32_ ( .D(data_in_2[134]), .E(n317), .CK(clk), .QN(n687) );
  EDFFXL R7_reg_33_ ( .D(data_in_2[135]), .E(n969), .CK(clk), .QN(n924) );
  EDFFXL R11_reg_33_ ( .D(data_in_2[135]), .E(n317), .CK(clk), .QN(n686) );
  EDFFXL R7_reg_15_ ( .D(data_in_2[117]), .E(n969), .CK(clk), .QN(n942) );
  EDFFXL R3_reg_15_ ( .D(data_in_2[117]), .E(n318), .CK(clk), .QN(n874) );
  EDFFXL R7_reg_16_ ( .D(data_in_2[118]), .E(n969), .CK(clk), .QN(n941) );
  EDFFXL R3_reg_16_ ( .D(data_in_2[118]), .E(n318), .CK(clk), .QN(n873) );
  EDFFXL R15_reg_15_ ( .D(data_in_2[117]), .E(n971), .CK(clk), .QN(n806) );
  EDFFXL R11_reg_15_ ( .D(data_in_2[117]), .E(n317), .CK(clk), .QN(n704) );
  EDFFXL R11_reg_16_ ( .D(data_in_2[118]), .E(n317), .CK(clk), .QN(n703) );
  EDFFXL R15_reg_16_ ( .D(data_in_2[118]), .E(n971), .CK(clk), .QN(n805) );
  EDFFXL R6_reg_32_ ( .D(data_in_2[100]), .E(n969), .CK(clk), .QN(n891) );
  EDFFXL R2_reg_32_ ( .D(data_in_2[100]), .E(n318), .CK(clk), .QN(n823) );
  EDFFXL R14_reg_32_ ( .D(data_in_2[100]), .E(n971), .CK(clk), .QN(n755) );
  EDFFXL R10_reg_32_ ( .D(data_in_2[100]), .E(n317), .CK(clk), .QN(n721) );
  EDFFXL R6_reg_15_ ( .D(data_in_2[83]), .E(n969), .CK(clk), .QN(n908) );
  EDFFXL R2_reg_15_ ( .D(data_in_2[83]), .E(n318), .CK(clk), .QN(n840) );
  EDFFXL R14_reg_15_ ( .D(data_in_2[83]), .E(n971), .CK(clk), .QN(n772) );
  EDFFXL R10_reg_15_ ( .D(data_in_2[83]), .E(n317), .CK(clk), .QN(n738) );
  EDFFXL R3_reg_33_ ( .D(data_in_2[135]), .E(n318), .CK(clk), .QN(n856) );
  EDFFXL R15_reg_33_ ( .D(data_in_2[135]), .E(n971), .CK(clk), .QN(n788) );
  EDFFXL R6_reg_16_ ( .D(data_in_2[84]), .E(n969), .CK(clk), .QN(n907) );
  EDFFXL R2_reg_16_ ( .D(data_in_2[84]), .E(n318), .CK(clk), .QN(n839) );
  EDFFXL R6_reg_33_ ( .D(data_in_2[101]), .E(n969), .CK(clk), .QN(n890) );
  EDFFXL R2_reg_33_ ( .D(data_in_2[101]), .E(n318), .CK(clk), .QN(n822) );
  EDFFXL R14_reg_16_ ( .D(data_in_2[84]), .E(n971), .CK(clk), .QN(n771) );
  EDFFXL R10_reg_16_ ( .D(data_in_2[84]), .E(n317), .CK(clk), .QN(n737) );
  EDFFXL R14_reg_33_ ( .D(data_in_2[101]), .E(n971), .CK(clk), .QN(n754) );
  EDFFXL R10_reg_33_ ( .D(data_in_2[101]), .E(n317), .CK(clk), .QN(n720) );
  DFFHQX4 reg_flag_mux_reg ( .D(n1246), .CK(clk), .Q(reg_flag_mux) );
  EDFFXL R2_reg_25_ ( .D(data_in_2[93]), .E(n1196), .CK(clk), .QN(n830) );
  EDFFXL R14_reg_25_ ( .D(data_in_2[93]), .E(n971), .CK(clk), .QN(n762) );
  EDFFXL R10_reg_25_ ( .D(data_in_2[93]), .E(n1185), .CK(clk), .QN(n728) );
  EDFFXL R10_reg_10_ ( .D(data_in_2[78]), .E(n1187), .CK(clk), .QN(n743) );
  EDFFXL R14_reg_10_ ( .D(data_in_2[78]), .E(n971), .CK(clk), .QN(n777) );
  EDFFXL R2_reg_10_ ( .D(data_in_2[78]), .E(n1195), .CK(clk), .QN(n845) );
  EDFFXL R11_reg_25_ ( .D(data_in_2[127]), .E(n1188), .CK(clk), .QN(n694) );
  EDFFXL R15_reg_25_ ( .D(data_in_2[127]), .E(n971), .CK(clk), .QN(n796) );
  EDFFXL R3_reg_25_ ( .D(data_in_2[127]), .E(n1195), .CK(clk), .QN(n864) );
  EDFFXL R0_reg_10_ ( .D(data_in_2[10]), .E(n1195), .CK(clk), .Q(R0[10]) );
  EDFFXL R8_reg_10_ ( .D(data_in_2[10]), .E(n1189), .CK(clk), .Q(R8[10]) );
  EDFFXL R12_reg_10_ ( .D(data_in_2[10]), .E(n1207), .CK(clk), .Q(R12[10]) );
  EDFFX2 R10_reg_14_ ( .D(data_in_2[82]), .E(n317), .CK(clk), .QN(n739) );
  EDFFX2 R14_reg_14_ ( .D(data_in_2[82]), .E(n971), .CK(clk), .QN(n773) );
  EDFFX2 R2_reg_14_ ( .D(data_in_2[82]), .E(n318), .CK(clk), .QN(n841) );
  EDFFX2 R6_reg_14_ ( .D(data_in_2[82]), .E(n969), .CK(clk), .QN(n909) );
  EDFFXL R11_reg_29_ ( .D(data_in_2[131]), .E(n1185), .CK(clk), .QN(n690) );
  EDFFXL R15_reg_29_ ( .D(data_in_2[131]), .E(n1210), .CK(clk), .QN(n792) );
  EDFFXL R3_reg_29_ ( .D(data_in_2[131]), .E(n1196), .CK(clk), .QN(n860) );
  EDFFXL R11_reg_10_ ( .D(data_in_2[112]), .E(n317), .CK(clk), .QN(n709) );
  EDFFXL R15_reg_10_ ( .D(data_in_2[112]), .E(n1206), .CK(clk), .QN(n811) );
  EDFFXL R3_reg_10_ ( .D(data_in_2[112]), .E(n1194), .CK(clk), .QN(n879) );
  EDFFXL R15_reg_28_ ( .D(data_in_2[130]), .E(n1211), .CK(clk), .QN(n793) );
  EDFFXL R11_reg_28_ ( .D(data_in_2[130]), .E(n1186), .CK(clk), .QN(n691) );
  EDFFXL R3_reg_28_ ( .D(data_in_2[130]), .E(n1195), .CK(clk), .QN(n861) );
  EDFFXL R10_reg_11_ ( .D(data_in_2[79]), .E(n1187), .CK(clk), .QN(n742) );
  EDFFXL R14_reg_11_ ( .D(data_in_2[79]), .E(n1206), .CK(clk), .QN(n776) );
  EDFFXL R2_reg_11_ ( .D(data_in_2[79]), .E(n1195), .CK(clk), .QN(n844) );
  EDFFXL R3_reg_24_ ( .D(data_in_2[126]), .E(n1195), .CK(clk), .QN(n865) );
  EDFFXL R15_reg_24_ ( .D(data_in_2[126]), .E(n1210), .CK(clk), .QN(n797) );
  EDFFXL R11_reg_24_ ( .D(data_in_2[126]), .E(n1188), .CK(clk), .QN(n695) );
  EDFFXL R0_reg_9_ ( .D(data_in_2[9]), .E(n1194), .CK(clk), .Q(R0[9]) );
  EDFFXL R8_reg_9_ ( .D(data_in_2[9]), .E(n1189), .CK(clk), .Q(R8[9]) );
  EDFFXL R12_reg_9_ ( .D(data_in_2[9]), .E(n1207), .CK(clk), .Q(R12[9]) );
  EDFFXL R0_reg_5_ ( .D(data_in_2[5]), .E(n1194), .CK(clk), .Q(R0[5]) );
  EDFFXL R8_reg_5_ ( .D(data_in_2[5]), .E(n1185), .CK(clk), .Q(R8[5]) );
  EDFFXL R12_reg_5_ ( .D(data_in_2[5]), .E(n1207), .CK(clk), .Q(R12[5]) );
  EDFFXL R10_reg_28_ ( .D(data_in_2[96]), .E(n1191), .CK(clk), .QN(n725) );
  EDFFXL R2_reg_28_ ( .D(data_in_2[96]), .E(n1196), .CK(clk), .QN(n827) );
  EDFFXL R14_reg_28_ ( .D(data_in_2[96]), .E(n1211), .CK(clk), .QN(n759) );
  EDFFXL R11_reg_27_ ( .D(data_in_2[129]), .E(n1188), .CK(clk), .QN(n692) );
  EDFFXL R15_reg_27_ ( .D(data_in_2[129]), .E(n1211), .CK(clk), .QN(n794) );
  EDFFXL R3_reg_27_ ( .D(data_in_2[129]), .E(n1194), .CK(clk), .QN(n862) );
  MX2X2 U3 ( .A(R0[33]), .B(data_in_2[33]), .S0(n1194), .Y(n654) );
  MX2X2 U4 ( .A(R12[33]), .B(data_in_2[33]), .S0(n1208), .Y(n660) );
  MX2X2 U5 ( .A(R8[33]), .B(data_in_2[33]), .S0(n1191), .Y(n658) );
  MX2X2 U6 ( .A(R4[33]), .B(data_in_2[33]), .S0(n1214), .Y(n656) );
  MX2X2 U7 ( .A(R0[12]), .B(data_in_2[12]), .S0(n1194), .Y(n1166) );
  MX2X2 U8 ( .A(R12[12]), .B(data_in_2[12]), .S0(n1207), .Y(n1172) );
  MX2X2 U9 ( .A(R8[12]), .B(data_in_2[12]), .S0(n1189), .Y(n1170) );
  MX2X2 U10 ( .A(R4[12]), .B(data_in_2[12]), .S0(n1215), .Y(n1168) );
  MX2X2 U11 ( .A(R0[13]), .B(data_in_2[13]), .S0(n1195), .Y(n1150) );
  MX2X2 U12 ( .A(R12[13]), .B(data_in_2[13]), .S0(n1207), .Y(n1156) );
  MX2X2 U13 ( .A(R8[13]), .B(data_in_2[13]), .S0(n1189), .Y(n1154) );
  MX2X2 U14 ( .A(R4[13]), .B(data_in_2[13]), .S0(n1215), .Y(n1152) );
  MX2X2 U15 ( .A(R0[14]), .B(data_in_2[14]), .S0(n1194), .Y(n638) );
  MX2X2 U16 ( .A(R12[14]), .B(data_in_2[14]), .S0(n1207), .Y(n644) );
  MX2X2 U17 ( .A(R8[14]), .B(data_in_2[14]), .S0(n1189), .Y(n642) );
  MX2X2 U18 ( .A(R4[14]), .B(data_in_2[14]), .S0(n1214), .Y(n640) );
  MX2X2 U19 ( .A(R0[31]), .B(data_in_2[31]), .S0(n1194), .Y(n678) );
  MX2X2 U20 ( .A(R12[31]), .B(data_in_2[31]), .S0(n1208), .Y(n684) );
  MX2X2 U21 ( .A(R4[31]), .B(data_in_2[31]), .S0(n1214), .Y(n680) );
  MX2X2 U22 ( .A(R8[31]), .B(data_in_2[31]), .S0(n1191), .Y(n682) );
  MX2X2 U23 ( .A(data_in_2[64]), .B(R9[30]), .S0(n1193), .Y(n1178) );
  MX2X2 U24 ( .A(R5[30]), .B(data_in_2[64]), .S0(n1215), .Y(n1176) );
  MX2X2 U25 ( .A(R1[30]), .B(data_in_2[64]), .S0(n1194), .Y(n1174) );
  MX2X2 U26 ( .A(R13[30]), .B(data_in_2[64]), .S0(n1211), .Y(n1180) );
  MX2X2 U27 ( .A(R1[15]), .B(data_in_2[49]), .S0(n1195), .Y(n614) );
  MX2X2 U28 ( .A(R13[15]), .B(data_in_2[49]), .S0(n1209), .Y(n620) );
  MX2X2 U29 ( .A(R5[15]), .B(data_in_2[49]), .S0(n1216), .Y(n616) );
  MX2X2 U30 ( .A(R9[15]), .B(data_in_2[49]), .S0(n317), .Y(n618) );
  MX2X2 U31 ( .A(data_in_2[65]), .B(R1[31]), .S0(n7), .Y(n1134) );
  CLKINVX20 U32 ( .A(n1194), .Y(n7) );
  MX2X2 U33 ( .A(R13[31]), .B(data_in_2[65]), .S0(n1211), .Y(n1140) );
  MX2X2 U34 ( .A(R5[31]), .B(data_in_2[65]), .S0(n1215), .Y(n1136) );
  MX2X2 U35 ( .A(data_in_2[50]), .B(R1[16]), .S0(n8), .Y(n670) );
  CLKINVX20 U36 ( .A(n1195), .Y(n8) );
  INVXL U37 ( .A(n971), .Y(n1212) );
  OR2X2 U38 ( .A(counter2[0]), .B(counter2[1]), .Y(n9) );
  OR2X2 U39 ( .A(n1249), .B(counter2[1]), .Y(n10) );
  AND3X2 U40 ( .A(counter1[0]), .B(n1248), .C(reg_datain_flag), .Y(n318) );
  INVX1 U41 ( .A(n1214), .Y(n245) );
  INVX1 U42 ( .A(n1197), .Y(n1196) );
  MX2X2 U43 ( .A(R4[29]), .B(data_in_2[29]), .S0(n1214), .Y(n1182) );
  MX2X2 U44 ( .A(R0[29]), .B(data_in_2[29]), .S0(n1194), .Y(n1181) );
  MX2X2 U45 ( .A(R12[29]), .B(data_in_2[29]), .S0(n1208), .Y(n1184) );
  MX2X2 U46 ( .A(R8[29]), .B(data_in_2[29]), .S0(n1190), .Y(n1183) );
  MX2X4 U47 ( .A(data_in_2[30]), .B(R12[30]), .S0(n1213), .Y(n1124) );
  MX2X2 U48 ( .A(R13[12]), .B(n45), .S0(n1209), .Y(n1164) );
  MX2X2 U49 ( .A(R5[12]), .B(n45), .S0(n1216), .Y(n1160) );
  MX2X2 U50 ( .A(R1[12]), .B(n45), .S0(n1195), .Y(n1158) );
  MX2X2 U51 ( .A(R9[12]), .B(n45), .S0(n317), .Y(n1162) );
  BUFX8 U52 ( .A(data_in_2[46]), .Y(n45) );
  MX2X2 U53 ( .A(R13[14]), .B(data_in_2[48]), .S0(n1209), .Y(n1132) );
  MX2X2 U54 ( .A(R9[14]), .B(data_in_2[48]), .S0(n317), .Y(n1130) );
  MX2X2 U55 ( .A(R1[14]), .B(data_in_2[48]), .S0(n1195), .Y(n1126) );
  MX2X2 U56 ( .A(R5[14]), .B(data_in_2[48]), .S0(n1216), .Y(n1128) );
  MX2X2 U57 ( .A(R8[16]), .B(data_in_2[16]), .S0(n1189), .Y(n970) );
  MX2X2 U58 ( .A(R12[16]), .B(data_in_2[16]), .S0(n971), .Y(n977) );
  MX2X2 U59 ( .A(R4[16]), .B(data_in_2[16]), .S0(n1214), .Y(n960) );
  MX2X2 U60 ( .A(R0[16]), .B(data_in_2[16]), .S0(n1194), .Y(n958) );
  MX2X2 U61 ( .A(R13[32]), .B(data_in_2[66]), .S0(n1211), .Y(n652) );
  MX2X2 U62 ( .A(R5[32]), .B(data_in_2[66]), .S0(n1215), .Y(n648) );
  MX2X2 U63 ( .A(data_in_2[50]), .B(R13[16]), .S0(n1212), .Y(n676) );
  MX2X2 U64 ( .A(data_in_2[50]), .B(R9[16]), .S0(n1193), .Y(n674) );
  MX2X2 U65 ( .A(data_in_2[67]), .B(R13[33]), .S0(n1212), .Y(n636) );
  MX2X2 U66 ( .A(R1[32]), .B(data_in_2[66]), .S0(n1195), .Y(n646) );
  MX2X2 U67 ( .A(R9[32]), .B(data_in_2[66]), .S0(n1186), .Y(n650) );
  MX2X4 U68 ( .A(R9[31]), .B(data_in_2[65]), .S0(n1186), .Y(n1138) );
  MX2X2 U69 ( .A(data_in_2[67]), .B(R5[33]), .S0(n245), .Y(n632) );
  MX2X2 U70 ( .A(data_in_2[67]), .B(R1[33]), .S0(n1197), .Y(n630) );
  MX2X2 U71 ( .A(data_in_2[67]), .B(R9[33]), .S0(n1192), .Y(n634) );
  MX2X2 U72 ( .A(R5[16]), .B(data_in_2[50]), .S0(n1216), .Y(n672) );
  AND2X4 U73 ( .A(reg_datain_flag), .B(n964), .Y(n317) );
  NOR2X4 U74 ( .A(n973), .B(n1248), .Y(n969) );
  NAND2X1 U75 ( .A(reg_datain_flag), .B(n1247), .Y(n973) );
  NOR2X4 U76 ( .A(n973), .B(counter1[1]), .Y(n971) );
  MX2X2 U77 ( .A(R0[30]), .B(data_in_2[30]), .S0(n1194), .Y(n1118) );
  MX2X2 U78 ( .A(R8[30]), .B(data_in_2[30]), .S0(n1191), .Y(n1122) );
  MX2X2 U79 ( .A(data_in_2[30]), .B(R4[30]), .S0(n245), .Y(n1120) );
  MX2X2 U80 ( .A(R13[13]), .B(data_in_2[47]), .S0(n1209), .Y(n1148) );
  MX2X2 U81 ( .A(R9[13]), .B(data_in_2[47]), .S0(n317), .Y(n1146) );
  MX2X2 U82 ( .A(R5[13]), .B(data_in_2[47]), .S0(n1216), .Y(n1144) );
  MX2X2 U83 ( .A(R1[13]), .B(data_in_2[47]), .S0(n1195), .Y(n1142) );
  CLKINVX3 U84 ( .A(n1217), .Y(n1216) );
  CLKINVX3 U85 ( .A(n1217), .Y(n1215) );
  INVX1 U86 ( .A(n1213), .Y(n1206) );
  INVX1 U87 ( .A(n1212), .Y(n1210) );
  INVX1 U88 ( .A(n1213), .Y(n1207) );
  INVX1 U89 ( .A(n1213), .Y(n1208) );
  INVX1 U90 ( .A(n1213), .Y(n1209) );
  INVX1 U91 ( .A(n969), .Y(n1217) );
  CLKINVX3 U92 ( .A(n1217), .Y(n1214) );
  INVX1 U93 ( .A(n10), .Y(n1232) );
  INVX1 U94 ( .A(n10), .Y(n1233) );
  INVX1 U95 ( .A(n10), .Y(n1234) );
  INVX1 U96 ( .A(n10), .Y(n1227) );
  INVX1 U97 ( .A(n10), .Y(n1228) );
  INVX1 U98 ( .A(n10), .Y(n1229) );
  INVX1 U99 ( .A(n10), .Y(n1230) );
  INVX1 U100 ( .A(n10), .Y(n1231) );
  CLKINVX3 U101 ( .A(n1197), .Y(n1195) );
  INVX1 U102 ( .A(n9), .Y(n1203) );
  INVX1 U103 ( .A(n9), .Y(n1204) );
  INVX1 U104 ( .A(n9), .Y(n1205) );
  INVX1 U105 ( .A(n9), .Y(n1198) );
  INVX1 U106 ( .A(n9), .Y(n1199) );
  INVX1 U107 ( .A(n9), .Y(n1200) );
  INVX1 U108 ( .A(n9), .Y(n1201) );
  INVX1 U109 ( .A(n9), .Y(n1202) );
  INVX1 U110 ( .A(n1242), .Y(n1237) );
  INVX1 U111 ( .A(n1242), .Y(n1236) );
  INVX1 U112 ( .A(n1242), .Y(n1241) );
  INVX1 U113 ( .A(n1242), .Y(n1240) );
  INVX1 U114 ( .A(n1242), .Y(n1239) );
  INVX1 U115 ( .A(n1242), .Y(n1238) );
  INVX1 U116 ( .A(n1225), .Y(n1222) );
  INVX1 U117 ( .A(n1225), .Y(n1223) );
  INVX1 U118 ( .A(n1225), .Y(n1224) );
  INVX1 U119 ( .A(n1225), .Y(n1218) );
  INVX1 U120 ( .A(n1225), .Y(n1219) );
  INVX1 U121 ( .A(n1225), .Y(n1220) );
  INVX1 U122 ( .A(n1225), .Y(n1221) );
  INVX1 U123 ( .A(n1193), .Y(n1185) );
  INVX1 U124 ( .A(n1192), .Y(n1188) );
  INVX1 U125 ( .A(n1192), .Y(n1190) );
  INVX1 U126 ( .A(n1192), .Y(n1187) );
  INVX1 U127 ( .A(n1192), .Y(n1186) );
  INVX1 U128 ( .A(n1193), .Y(n1189) );
  INVX1 U129 ( .A(n1193), .Y(n1191) );
  INVX1 U130 ( .A(n1212), .Y(n1211) );
  INVX1 U131 ( .A(n966), .Y(n1250) );
  INVX1 U132 ( .A(n971), .Y(n1213) );
  NOR2X1 U133 ( .A(n1248), .B(n1247), .Y(n964) );
  INVX1 U134 ( .A(n10), .Y(n1226) );
  CLKINVX3 U135 ( .A(n1197), .Y(n1194) );
  INVX1 U136 ( .A(n318), .Y(n1197) );
  CLKINVX3 U137 ( .A(n1245), .Y(n1244) );
  CLKINVX3 U138 ( .A(n1245), .Y(n1243) );
  INVX1 U139 ( .A(n1242), .Y(n1235) );
  INVX1 U140 ( .A(n968), .Y(n1225) );
  INVX1 U141 ( .A(n317), .Y(n1193) );
  INVX1 U142 ( .A(n317), .Y(n1192) );
  INVX1 U143 ( .A(n963), .Y(n1242) );
  OAI32X1 U144 ( .A0(n961), .A1(counter2[0]), .A2(n966), .B0(n1249), .B1(n1250), .Y(n1114) );
  NOR2X1 U145 ( .A(n961), .B(reg_flag_mux), .Y(n966) );
  OAI22X1 U146 ( .A0(n1247), .A1(n974), .B0(n961), .B1(n973), .Y(n1116) );
  NAND2BX1 U147 ( .AN(reg_datain_flag), .B(rst_n), .Y(n974) );
  OAI21XL U148 ( .A0(n1248), .A1(n974), .B0(n975), .Y(n1115) );
  OAI21XL U149 ( .A0(n1194), .A1(n1214), .B0(rst_n), .Y(n975) );
  OAI2BB2X1 U150 ( .B0(n965), .B1(n961), .A0N(counter2[1]), .A1N(n966), .Y(
        n1113) );
  AOI21X1 U151 ( .A0(n1230), .A1(n1250), .B0(n1225), .Y(n965) );
  INVX1 U152 ( .A(n962), .Y(n1246) );
  AOI32X1 U153 ( .A0(n1243), .A1(n1235), .A2(rst_n), .B0(n964), .B1(rst_n), 
        .Y(n962) );
  AOI22X1 U154 ( .A0(R13[28]), .A1(n1231), .B0(n1200), .B1(R12[28]), .Y(n1030)
         );
  NAND2X1 U155 ( .A(counter2[1]), .B(n1249), .Y(n968) );
  NAND2X1 U156 ( .A(counter2[1]), .B(counter2[0]), .Y(n963) );
  OAI221XL U157 ( .A0(n877), .A1(n1237), .B0(n843), .B1(n1222), .C0(n1012), 
        .Y(N64) );
  AOI22X1 U158 ( .A0(R1[12]), .A1(n1232), .B0(n1203), .B1(R0[12]), .Y(n1012)
         );
  OAI221XL U159 ( .A0(n876), .A1(n1237), .B0(n842), .B1(n1222), .C0(n1011), 
        .Y(N65) );
  AOI22X1 U160 ( .A0(R1[13]), .A1(n1232), .B0(n1203), .B1(R0[13]), .Y(n1011)
         );
  OAI221XL U161 ( .A0(n875), .A1(n1237), .B0(n841), .B1(n1222), .C0(n1010), 
        .Y(N66) );
  AOI22X1 U162 ( .A0(R1[14]), .A1(n1232), .B0(n1203), .B1(R0[14]), .Y(n1010)
         );
  OAI221XL U163 ( .A0(n874), .A1(n1237), .B0(n840), .B1(n1222), .C0(n1009), 
        .Y(N67) );
  AOI22X1 U164 ( .A0(R1[15]), .A1(n1232), .B0(n1203), .B1(R0[15]), .Y(n1009)
         );
  OAI221XL U165 ( .A0(n873), .A1(n1237), .B0(n839), .B1(n1222), .C0(n1008), 
        .Y(N68) );
  AOI22X1 U166 ( .A0(R1[16]), .A1(n1233), .B0(n1203), .B1(R0[16]), .Y(n1008)
         );
  OAI221XL U167 ( .A0(n860), .A1(n1236), .B0(n826), .B1(n1223), .C0(n995), .Y(
        N81) );
  AOI22X1 U168 ( .A0(R1[29]), .A1(n1234), .B0(n1204), .B1(R0[29]), .Y(n995) );
  OAI221XL U169 ( .A0(n859), .A1(n1236), .B0(n825), .B1(n1223), .C0(n994), .Y(
        N82) );
  AOI22X1 U170 ( .A0(R1[30]), .A1(n1234), .B0(n1204), .B1(R0[30]), .Y(n994) );
  OAI221XL U171 ( .A0(n858), .A1(n1236), .B0(n824), .B1(n1223), .C0(n993), .Y(
        N83) );
  AOI22X1 U172 ( .A0(R1[31]), .A1(n1234), .B0(n1204), .B1(R0[31]), .Y(n993) );
  OAI221XL U173 ( .A0(n857), .A1(n1236), .B0(n823), .B1(n1224), .C0(n992), .Y(
        N84) );
  AOI22X1 U174 ( .A0(R1[32]), .A1(n1234), .B0(n1205), .B1(R0[32]), .Y(n992) );
  OAI221XL U175 ( .A0(n856), .A1(n1236), .B0(n822), .B1(n1224), .C0(n991), .Y(
        N85) );
  AOI22X1 U176 ( .A0(R1[33]), .A1(n1234), .B0(n1205), .B1(R0[33]), .Y(n991) );
  OAI221XL U177 ( .A0(n945), .A1(n1235), .B0(n911), .B1(n1223), .C0(n978), .Y(
        N98) );
  AOI22X1 U178 ( .A0(R5[12]), .A1(n1233), .B0(n1205), .B1(R4[12]), .Y(n978) );
  OAI221XL U179 ( .A0(n944), .A1(n1235), .B0(n910), .B1(n1222), .C0(n976), .Y(
        N99) );
  AOI22X1 U180 ( .A0(R5[13]), .A1(n1232), .B0(n1205), .B1(R4[13]), .Y(n976) );
  OAI221XL U181 ( .A0(n943), .A1(n1235), .B0(n909), .B1(n1218), .C0(n1112), 
        .Y(N100) );
  AOI22X1 U182 ( .A0(R5[14]), .A1(n1226), .B0(n1198), .B1(R4[14]), .Y(n1112)
         );
  OAI221XL U183 ( .A0(n942), .A1(n963), .B0(n908), .B1(n1218), .C0(n1111), .Y(
        N101) );
  AOI22X1 U184 ( .A0(R5[15]), .A1(n1226), .B0(n1198), .B1(R4[15]), .Y(n1111)
         );
  OAI221XL U185 ( .A0(n941), .A1(n963), .B0(n907), .B1(n1218), .C0(n1110), .Y(
        N102) );
  AOI22X1 U186 ( .A0(R5[16]), .A1(n1226), .B0(n1198), .B1(R4[16]), .Y(n1110)
         );
  OAI221XL U187 ( .A0(n928), .A1(n963), .B0(n894), .B1(n1219), .C0(n1097), .Y(
        N115) );
  AOI22X1 U188 ( .A0(R5[29]), .A1(n1227), .B0(n1199), .B1(R4[29]), .Y(n1097)
         );
  OAI221XL U189 ( .A0(n927), .A1(n1238), .B0(n893), .B1(n1219), .C0(n1096), 
        .Y(N116) );
  AOI22X1 U190 ( .A0(R5[30]), .A1(n1227), .B0(n1199), .B1(R4[30]), .Y(n1096)
         );
  OAI221XL U191 ( .A0(n926), .A1(n1241), .B0(n892), .B1(n1219), .C0(n1095), 
        .Y(N117) );
  AOI22X1 U192 ( .A0(R5[31]), .A1(n1227), .B0(n1199), .B1(R4[31]), .Y(n1095)
         );
  OAI221XL U193 ( .A0(n925), .A1(n963), .B0(n891), .B1(n1219), .C0(n1094), .Y(
        N118) );
  AOI22X1 U194 ( .A0(R5[32]), .A1(n1227), .B0(n1199), .B1(R4[32]), .Y(n1094)
         );
  OAI221XL U195 ( .A0(n924), .A1(n963), .B0(n890), .B1(n1219), .C0(n1093), .Y(
        N119) );
  AOI22X1 U196 ( .A0(R5[33]), .A1(n1227), .B0(n1199), .B1(R4[33]), .Y(n1093)
         );
  OAI221XL U197 ( .A0(n707), .A1(n1241), .B0(n741), .B1(n1220), .C0(n1080), 
        .Y(N132) );
  AOI22X1 U198 ( .A0(R9[12]), .A1(n1228), .B0(n1200), .B1(R8[12]), .Y(n1080)
         );
  OAI221XL U199 ( .A0(n706), .A1(n1240), .B0(n740), .B1(n1220), .C0(n1079), 
        .Y(N133) );
  AOI22X1 U200 ( .A0(R9[13]), .A1(n1228), .B0(n1200), .B1(R8[13]), .Y(n1079)
         );
  OAI221XL U201 ( .A0(n705), .A1(n1240), .B0(n739), .B1(n1220), .C0(n1078), 
        .Y(N134) );
  AOI22X1 U202 ( .A0(R9[14]), .A1(n1228), .B0(n1200), .B1(R8[14]), .Y(n1078)
         );
  OAI221XL U203 ( .A0(n704), .A1(n1240), .B0(n738), .B1(n1220), .C0(n1077), 
        .Y(N135) );
  AOI22X1 U204 ( .A0(R9[15]), .A1(n1228), .B0(n1200), .B1(R8[15]), .Y(n1077)
         );
  OAI221XL U205 ( .A0(n703), .A1(n1240), .B0(n737), .B1(n968), .C0(n1076), .Y(
        N136) );
  AOI22X1 U206 ( .A0(R9[16]), .A1(n1228), .B0(n1201), .B1(R8[16]), .Y(n1076)
         );
  OAI221XL U207 ( .A0(n690), .A1(n1239), .B0(n724), .B1(n1223), .C0(n1063), 
        .Y(N149) );
  AOI22X1 U208 ( .A0(R9[29]), .A1(n1231), .B0(n1201), .B1(R8[29]), .Y(n1063)
         );
  OAI221XL U209 ( .A0(n689), .A1(n1239), .B0(n723), .B1(n1222), .C0(n1062), 
        .Y(N150) );
  AOI22X1 U210 ( .A0(R9[30]), .A1(n1227), .B0(n1201), .B1(R8[30]), .Y(n1062)
         );
  OAI221XL U211 ( .A0(n688), .A1(n1239), .B0(n722), .B1(n968), .C0(n1061), .Y(
        N151) );
  AOI22X1 U212 ( .A0(R9[31]), .A1(n1227), .B0(n1201), .B1(R8[31]), .Y(n1061)
         );
  OAI221XL U213 ( .A0(n687), .A1(n1239), .B0(n721), .B1(n968), .C0(n1060), .Y(
        N152) );
  AOI22X1 U214 ( .A0(R9[32]), .A1(n1229), .B0(n1201), .B1(R8[32]), .Y(n1060)
         );
  OAI221XL U215 ( .A0(n686), .A1(n1239), .B0(n720), .B1(n968), .C0(n1059), .Y(
        N153) );
  AOI22X1 U216 ( .A0(R9[33]), .A1(n1229), .B0(n1201), .B1(R8[33]), .Y(n1059)
         );
  OAI221XL U217 ( .A0(n809), .A1(n1241), .B0(n775), .B1(n1221), .C0(n1046), 
        .Y(N166) );
  AOI22X1 U218 ( .A0(R13[12]), .A1(n1230), .B0(n1201), .B1(R12[12]), .Y(n1046)
         );
  OAI221XL U219 ( .A0(n808), .A1(n1240), .B0(n774), .B1(n1219), .C0(n1045), 
        .Y(N167) );
  AOI22X1 U220 ( .A0(R13[13]), .A1(n1230), .B0(n1203), .B1(R12[13]), .Y(n1045)
         );
  OAI221XL U221 ( .A0(n807), .A1(n1236), .B0(n773), .B1(n968), .C0(n1044), .Y(
        N168) );
  AOI22X1 U222 ( .A0(R13[14]), .A1(n1230), .B0(n1199), .B1(R12[14]), .Y(n1044)
         );
  OAI221XL U223 ( .A0(n806), .A1(n1238), .B0(n772), .B1(n968), .C0(n1043), .Y(
        N169) );
  AOI22X1 U224 ( .A0(R13[15]), .A1(n1230), .B0(n1204), .B1(R12[15]), .Y(n1043)
         );
  OAI221XL U225 ( .A0(n805), .A1(n1236), .B0(n771), .B1(n1223), .C0(n1042), 
        .Y(N170) );
  AOI22X1 U226 ( .A0(R13[16]), .A1(n1230), .B0(n1202), .B1(R12[16]), .Y(n1042)
         );
  OAI221XL U227 ( .A0(n792), .A1(n963), .B0(n758), .B1(n1224), .C0(n1029), .Y(
        N183) );
  AOI22X1 U228 ( .A0(R13[29]), .A1(n1231), .B0(n1203), .B1(R12[29]), .Y(n1029)
         );
  OAI221XL U229 ( .A0(n791), .A1(n1236), .B0(n757), .B1(n1221), .C0(n1028), 
        .Y(N184) );
  AOI22X1 U230 ( .A0(R13[30]), .A1(n1231), .B0(n1202), .B1(R12[30]), .Y(n1028)
         );
  OAI221XL U231 ( .A0(n790), .A1(n1238), .B0(n756), .B1(n1221), .C0(n1027), 
        .Y(N185) );
  AOI22X1 U232 ( .A0(R13[31]), .A1(n1231), .B0(n1202), .B1(R12[31]), .Y(n1027)
         );
  OAI221XL U233 ( .A0(n789), .A1(n1238), .B0(n755), .B1(n1221), .C0(n1026), 
        .Y(N186) );
  AOI22X1 U234 ( .A0(R13[32]), .A1(n1231), .B0(n1202), .B1(R12[32]), .Y(n1026)
         );
  OAI221XL U235 ( .A0(n788), .A1(n1238), .B0(n754), .B1(n1221), .C0(n1025), 
        .Y(N187) );
  AOI22X1 U236 ( .A0(R13[33]), .A1(n1231), .B0(n1202), .B1(R12[33]), .Y(n1025)
         );
  OAI221XL U237 ( .A0(n889), .A1(n1238), .B0(n855), .B1(n1221), .C0(n1024), 
        .Y(N52) );
  AOI22X1 U238 ( .A0(R1[0]), .A1(n1231), .B0(n1202), .B1(R0[0]), .Y(n1024) );
  OAI221XL U239 ( .A0(n888), .A1(n1238), .B0(n854), .B1(n1221), .C0(n1023), 
        .Y(N53) );
  AOI22X1 U240 ( .A0(R1[1]), .A1(n1231), .B0(n1202), .B1(R0[1]), .Y(n1023) );
  OAI221XL U241 ( .A0(n887), .A1(n1238), .B0(n853), .B1(n1221), .C0(n1022), 
        .Y(N54) );
  AOI22X1 U242 ( .A0(R1[2]), .A1(n1231), .B0(n1202), .B1(R0[2]), .Y(n1022) );
  OAI221XL U243 ( .A0(n886), .A1(n1238), .B0(n852), .B1(n1221), .C0(n1021), 
        .Y(N55) );
  AOI22X1 U244 ( .A0(R1[3]), .A1(n1232), .B0(n1202), .B1(R0[3]), .Y(n1021) );
  OAI221XL U245 ( .A0(n885), .A1(n1238), .B0(n851), .B1(n1221), .C0(n1020), 
        .Y(N56) );
  AOI22X1 U246 ( .A0(R1[4]), .A1(n1232), .B0(n1202), .B1(R0[4]), .Y(n1020) );
  OAI221XL U247 ( .A0(n884), .A1(n1238), .B0(n850), .B1(n1221), .C0(n1019), 
        .Y(N57) );
  AOI22X1 U248 ( .A0(R1[5]), .A1(n1232), .B0(n1202), .B1(R0[5]), .Y(n1019) );
  OAI221XL U249 ( .A0(n883), .A1(n1238), .B0(n849), .B1(n1221), .C0(n1018), 
        .Y(N58) );
  AOI22X1 U250 ( .A0(R1[6]), .A1(n1232), .B0(n1202), .B1(R0[6]), .Y(n1018) );
  OAI221XL U251 ( .A0(n882), .A1(n1238), .B0(n848), .B1(n1221), .C0(n1017), 
        .Y(N59) );
  AOI22X1 U252 ( .A0(R1[7]), .A1(n1232), .B0(n1202), .B1(R0[7]), .Y(n1017) );
  OAI221XL U253 ( .A0(n881), .A1(n1238), .B0(n847), .B1(n1222), .C0(n1016), 
        .Y(N60) );
  AOI22X1 U254 ( .A0(R1[8]), .A1(n1232), .B0(n1203), .B1(R0[8]), .Y(n1016) );
  OAI221XL U255 ( .A0(n880), .A1(n1238), .B0(n846), .B1(n1222), .C0(n1015), 
        .Y(N61) );
  AOI22X1 U256 ( .A0(R1[9]), .A1(n1232), .B0(n1203), .B1(R0[9]), .Y(n1015) );
  OAI221XL U257 ( .A0(n879), .A1(n1237), .B0(n845), .B1(n1222), .C0(n1014), 
        .Y(N62) );
  AOI22X1 U258 ( .A0(R1[10]), .A1(n1232), .B0(n1203), .B1(R0[10]), .Y(n1014)
         );
  OAI221XL U259 ( .A0(n878), .A1(n1237), .B0(n844), .B1(n1222), .C0(n1013), 
        .Y(N63) );
  AOI22X1 U260 ( .A0(R1[11]), .A1(n1232), .B0(n1203), .B1(R0[11]), .Y(n1013)
         );
  OAI221XL U261 ( .A0(n872), .A1(n1237), .B0(n838), .B1(n1222), .C0(n1007), 
        .Y(N69) );
  AOI22X1 U262 ( .A0(R1[17]), .A1(n1233), .B0(n1203), .B1(R0[17]), .Y(n1007)
         );
  OAI221XL U263 ( .A0(n871), .A1(n1237), .B0(n837), .B1(n1222), .C0(n1006), 
        .Y(N70) );
  AOI22X1 U264 ( .A0(R1[18]), .A1(n1233), .B0(n1203), .B1(R0[18]), .Y(n1006)
         );
  OAI221XL U265 ( .A0(n870), .A1(n1237), .B0(n836), .B1(n1222), .C0(n1005), 
        .Y(N71) );
  AOI22X1 U266 ( .A0(R1[19]), .A1(n1233), .B0(n1203), .B1(R0[19]), .Y(n1005)
         );
  OAI221XL U267 ( .A0(n869), .A1(n1237), .B0(n835), .B1(n1223), .C0(n1004), 
        .Y(N72) );
  AOI22X1 U268 ( .A0(R1[20]), .A1(n1233), .B0(n1204), .B1(R0[20]), .Y(n1004)
         );
  OAI221XL U269 ( .A0(n868), .A1(n1237), .B0(n834), .B1(n1223), .C0(n1003), 
        .Y(N73) );
  AOI22X1 U270 ( .A0(R1[21]), .A1(n1233), .B0(n1204), .B1(R0[21]), .Y(n1003)
         );
  OAI221XL U271 ( .A0(n867), .A1(n1237), .B0(n833), .B1(n1223), .C0(n1002), 
        .Y(N74) );
  AOI22X1 U272 ( .A0(R1[22]), .A1(n1233), .B0(n1204), .B1(R0[22]), .Y(n1002)
         );
  OAI221XL U273 ( .A0(n866), .A1(n1236), .B0(n832), .B1(n1223), .C0(n1001), 
        .Y(N75) );
  AOI22X1 U274 ( .A0(R1[23]), .A1(n1233), .B0(n1204), .B1(R0[23]), .Y(n1001)
         );
  OAI221XL U275 ( .A0(n865), .A1(n1236), .B0(n831), .B1(n1223), .C0(n1000), 
        .Y(N76) );
  AOI22X1 U276 ( .A0(R1[24]), .A1(n1233), .B0(n1204), .B1(R0[24]), .Y(n1000)
         );
  OAI221XL U277 ( .A0(n864), .A1(n1236), .B0(n830), .B1(n1223), .C0(n999), .Y(
        N77) );
  AOI22X1 U278 ( .A0(R1[25]), .A1(n1233), .B0(n1204), .B1(R0[25]), .Y(n999) );
  OAI221XL U279 ( .A0(n863), .A1(n1236), .B0(n829), .B1(n1223), .C0(n998), .Y(
        N78) );
  AOI22X1 U280 ( .A0(R1[26]), .A1(n1233), .B0(n1204), .B1(R0[26]), .Y(n998) );
  OAI221XL U281 ( .A0(n862), .A1(n1236), .B0(n828), .B1(n1223), .C0(n997), .Y(
        N79) );
  AOI22X1 U282 ( .A0(R1[27]), .A1(n1233), .B0(n1204), .B1(R0[27]), .Y(n997) );
  OAI221XL U283 ( .A0(n861), .A1(n1236), .B0(n827), .B1(n1223), .C0(n996), .Y(
        N80) );
  AOI22X1 U284 ( .A0(R1[28]), .A1(n1233), .B0(n1204), .B1(R0[28]), .Y(n996) );
  OAI221XL U285 ( .A0(n957), .A1(n1236), .B0(n923), .B1(n1224), .C0(n990), .Y(
        N86) );
  AOI22X1 U286 ( .A0(R5[0]), .A1(n1234), .B0(n1205), .B1(R4[0]), .Y(n990) );
  OAI221XL U287 ( .A0(n956), .A1(n1236), .B0(n922), .B1(n1224), .C0(n989), .Y(
        N87) );
  AOI22X1 U288 ( .A0(R5[1]), .A1(n1234), .B0(n1205), .B1(R4[1]), .Y(n989) );
  OAI221XL U289 ( .A0(n955), .A1(n1235), .B0(n921), .B1(n1224), .C0(n988), .Y(
        N88) );
  AOI22X1 U290 ( .A0(R5[2]), .A1(n1234), .B0(n1205), .B1(R4[2]), .Y(n988) );
  OAI221XL U291 ( .A0(n954), .A1(n1235), .B0(n920), .B1(n1224), .C0(n987), .Y(
        N89) );
  AOI22X1 U292 ( .A0(R5[3]), .A1(n1234), .B0(n1205), .B1(R4[3]), .Y(n987) );
  OAI221XL U293 ( .A0(n953), .A1(n1235), .B0(n919), .B1(n1224), .C0(n986), .Y(
        N90) );
  AOI22X1 U294 ( .A0(R5[4]), .A1(n1234), .B0(n1205), .B1(R4[4]), .Y(n986) );
  OAI221XL U295 ( .A0(n952), .A1(n1235), .B0(n918), .B1(n1224), .C0(n985), .Y(
        N91) );
  AOI22X1 U296 ( .A0(R5[5]), .A1(n1234), .B0(n1205), .B1(R4[5]), .Y(n985) );
  OAI221XL U297 ( .A0(n951), .A1(n1235), .B0(n917), .B1(n1224), .C0(n984), .Y(
        N92) );
  AOI22X1 U298 ( .A0(R5[6]), .A1(n1234), .B0(n1205), .B1(R4[6]), .Y(n984) );
  OAI221XL U299 ( .A0(n950), .A1(n1235), .B0(n916), .B1(n1224), .C0(n983), .Y(
        N93) );
  AOI22X1 U300 ( .A0(R5[7]), .A1(n1234), .B0(n1205), .B1(R4[7]), .Y(n983) );
  OAI221XL U301 ( .A0(n949), .A1(n1235), .B0(n915), .B1(n1224), .C0(n982), .Y(
        N94) );
  AOI22X1 U303 ( .A0(R5[8]), .A1(n1233), .B0(n1205), .B1(R4[8]), .Y(n982) );
  OAI221XL U304 ( .A0(n948), .A1(n1235), .B0(n914), .B1(n1224), .C0(n981), .Y(
        N95) );
  AOI22X1 U305 ( .A0(R5[9]), .A1(n1232), .B0(n1205), .B1(R4[9]), .Y(n981) );
  OAI221XL U306 ( .A0(n947), .A1(n1235), .B0(n913), .B1(n1219), .C0(n980), .Y(
        N96) );
  AOI22X1 U307 ( .A0(R5[10]), .A1(n1228), .B0(n1203), .B1(R4[10]), .Y(n980) );
  OAI221XL U308 ( .A0(n946), .A1(n1235), .B0(n912), .B1(n1219), .C0(n979), .Y(
        N97) );
  AOI22X1 U309 ( .A0(R5[11]), .A1(n1229), .B0(n1204), .B1(R4[11]), .Y(n979) );
  OAI221XL U310 ( .A0(n940), .A1(n1237), .B0(n906), .B1(n1218), .C0(n1109), 
        .Y(N103) );
  AOI22X1 U311 ( .A0(R5[17]), .A1(n1226), .B0(n1198), .B1(R4[17]), .Y(n1109)
         );
  OAI221XL U312 ( .A0(n939), .A1(n1239), .B0(n905), .B1(n1218), .C0(n1108), 
        .Y(N104) );
  AOI22X1 U313 ( .A0(R5[18]), .A1(n1226), .B0(n1198), .B1(R4[18]), .Y(n1108)
         );
  OAI221XL U314 ( .A0(n938), .A1(n1235), .B0(n904), .B1(n1218), .C0(n1107), 
        .Y(N105) );
  AOI22X1 U315 ( .A0(R5[19]), .A1(n1226), .B0(n1198), .B1(R4[19]), .Y(n1107)
         );
  OAI221XL U316 ( .A0(n937), .A1(n1237), .B0(n903), .B1(n1218), .C0(n1106), 
        .Y(N106) );
  AOI22X1 U317 ( .A0(R5[20]), .A1(n1226), .B0(n1198), .B1(R4[20]), .Y(n1106)
         );
  OAI221XL U318 ( .A0(n936), .A1(n1240), .B0(n902), .B1(n1218), .C0(n1105), 
        .Y(N107) );
  AOI22X1 U319 ( .A0(R5[21]), .A1(n1226), .B0(n1198), .B1(R4[21]), .Y(n1105)
         );
  OAI221XL U320 ( .A0(n935), .A1(n1235), .B0(n901), .B1(n1218), .C0(n1104), 
        .Y(N108) );
  AOI22X1 U321 ( .A0(R5[22]), .A1(n1226), .B0(n1198), .B1(R4[22]), .Y(n1104)
         );
  OAI221XL U322 ( .A0(n934), .A1(n963), .B0(n900), .B1(n1218), .C0(n1103), .Y(
        N109) );
  AOI22X1 U323 ( .A0(R5[23]), .A1(n1226), .B0(n1198), .B1(R4[23]), .Y(n1103)
         );
  OAI221XL U324 ( .A0(n933), .A1(n963), .B0(n899), .B1(n1218), .C0(n1102), .Y(
        N110) );
  AOI22X1 U325 ( .A0(R5[24]), .A1(n1226), .B0(n1198), .B1(R4[24]), .Y(n1102)
         );
  OAI221XL U326 ( .A0(n932), .A1(n963), .B0(n898), .B1(n1218), .C0(n1101), .Y(
        N111) );
  AOI22X1 U327 ( .A0(R5[25]), .A1(n1226), .B0(n1198), .B1(R4[25]), .Y(n1101)
         );
  OAI221XL U328 ( .A0(n931), .A1(n963), .B0(n897), .B1(n1219), .C0(n1100), .Y(
        N112) );
  AOI22X1 U329 ( .A0(R5[26]), .A1(n1226), .B0(n1199), .B1(R4[26]), .Y(n1100)
         );
  OAI221XL U330 ( .A0(n930), .A1(n963), .B0(n896), .B1(n1219), .C0(n1099), .Y(
        N113) );
  AOI22X1 U331 ( .A0(R5[27]), .A1(n1227), .B0(n1199), .B1(R4[27]), .Y(n1099)
         );
  OAI221XL U332 ( .A0(n929), .A1(n1237), .B0(n895), .B1(n1219), .C0(n1098), 
        .Y(N114) );
  AOI22X1 U333 ( .A0(R5[28]), .A1(n1227), .B0(n1199), .B1(R4[28]), .Y(n1098)
         );
  OAI221XL U334 ( .A0(n719), .A1(n1241), .B0(n753), .B1(n1219), .C0(n1092), 
        .Y(N120) );
  AOI22X1 U335 ( .A0(R9[0]), .A1(n1227), .B0(n1199), .B1(R8[0]), .Y(n1092) );
  OAI221XL U336 ( .A0(n718), .A1(n1241), .B0(n752), .B1(n1219), .C0(n1091), 
        .Y(N121) );
  AOI22X1 U337 ( .A0(R9[1]), .A1(n1227), .B0(n1199), .B1(R8[1]), .Y(n1091) );
  OAI221XL U338 ( .A0(n717), .A1(n1241), .B0(n751), .B1(n1219), .C0(n1090), 
        .Y(N122) );
  AOI22X1 U339 ( .A0(R9[2]), .A1(n1227), .B0(n1199), .B1(R8[2]), .Y(n1090) );
  OAI221XL U340 ( .A0(n716), .A1(n1241), .B0(n750), .B1(n1219), .C0(n1089), 
        .Y(N123) );
  AOI22X1 U341 ( .A0(R9[3]), .A1(n1227), .B0(n1199), .B1(R8[3]), .Y(n1089) );
  OAI221XL U342 ( .A0(n715), .A1(n1241), .B0(n749), .B1(n1220), .C0(n1088), 
        .Y(N124) );
  AOI22X1 U343 ( .A0(R9[4]), .A1(n1227), .B0(n1200), .B1(R8[4]), .Y(n1088) );
  OAI221XL U344 ( .A0(n714), .A1(n1241), .B0(n748), .B1(n1220), .C0(n1087), 
        .Y(N125) );
  AOI22X1 U345 ( .A0(R9[5]), .A1(n1227), .B0(n1200), .B1(R8[5]), .Y(n1087) );
  OAI221XL U346 ( .A0(n713), .A1(n1241), .B0(n747), .B1(n1220), .C0(n1086), 
        .Y(N126) );
  AOI22X1 U347 ( .A0(R9[6]), .A1(n1228), .B0(n1200), .B1(R8[6]), .Y(n1086) );
  OAI221XL U348 ( .A0(n712), .A1(n1241), .B0(n746), .B1(n1220), .C0(n1085), 
        .Y(N127) );
  AOI22X1 U349 ( .A0(R9[7]), .A1(n1228), .B0(n1200), .B1(R8[7]), .Y(n1085) );
  OAI221XL U350 ( .A0(n711), .A1(n1241), .B0(n745), .B1(n1220), .C0(n1084), 
        .Y(N128) );
  AOI22X1 U351 ( .A0(R9[8]), .A1(n1228), .B0(n1200), .B1(R8[8]), .Y(n1084) );
  OAI221XL U352 ( .A0(n710), .A1(n1241), .B0(n744), .B1(n1220), .C0(n1083), 
        .Y(N129) );
  AOI22X1 U353 ( .A0(R9[9]), .A1(n1228), .B0(n1200), .B1(R8[9]), .Y(n1083) );
  OAI221XL U354 ( .A0(n709), .A1(n1241), .B0(n743), .B1(n1220), .C0(n1082), 
        .Y(N130) );
  AOI22X1 U355 ( .A0(R9[10]), .A1(n1228), .B0(n1200), .B1(R8[10]), .Y(n1082)
         );
  OAI221XL U356 ( .A0(n708), .A1(n1241), .B0(n742), .B1(n1220), .C0(n1081), 
        .Y(N131) );
  AOI22X1 U357 ( .A0(R9[11]), .A1(n1228), .B0(n1200), .B1(R8[11]), .Y(n1081)
         );
  OAI221XL U358 ( .A0(n702), .A1(n1240), .B0(n736), .B1(n1223), .C0(n1075), 
        .Y(N137) );
  AOI22X1 U359 ( .A0(R9[17]), .A1(n1228), .B0(n1204), .B1(R8[17]), .Y(n1075)
         );
  OAI221XL U360 ( .A0(n701), .A1(n1240), .B0(n735), .B1(n1222), .C0(n1074), 
        .Y(N138) );
  AOI22X1 U361 ( .A0(R9[18]), .A1(n1228), .B0(n1204), .B1(R8[18]), .Y(n1074)
         );
  OAI221XL U362 ( .A0(n700), .A1(n1240), .B0(n734), .B1(n1219), .C0(n1073), 
        .Y(N139) );
  AOI22X1 U363 ( .A0(R9[19]), .A1(n1234), .B0(n1200), .B1(R8[19]), .Y(n1073)
         );
  OAI221XL U364 ( .A0(n699), .A1(n1240), .B0(n733), .B1(n1224), .C0(n1072), 
        .Y(N140) );
  AOI22X1 U365 ( .A0(R9[20]), .A1(n1228), .B0(n1202), .B1(R8[20]), .Y(n1072)
         );
  OAI221XL U366 ( .A0(n698), .A1(n1240), .B0(n732), .B1(n1223), .C0(n1071), 
        .Y(N141) );
  AOI22X1 U367 ( .A0(R9[21]), .A1(n1226), .B0(n1203), .B1(R8[21]), .Y(n1071)
         );
  OAI221XL U368 ( .A0(n697), .A1(n1240), .B0(n731), .B1(n1222), .C0(n1070), 
        .Y(N142) );
  AOI22X1 U369 ( .A0(R9[22]), .A1(n1231), .B0(n1200), .B1(R8[22]), .Y(n1070)
         );
  OAI221XL U370 ( .A0(n696), .A1(n1240), .B0(n730), .B1(n1218), .C0(n1069), 
        .Y(N143) );
  AOI22X1 U371 ( .A0(R9[23]), .A1(n1231), .B0(n1199), .B1(R8[23]), .Y(n1069)
         );
  OAI221XL U372 ( .A0(n695), .A1(n1240), .B0(n729), .B1(n1220), .C0(n1068), 
        .Y(N144) );
  AOI22X1 U373 ( .A0(R9[24]), .A1(n1227), .B0(n1203), .B1(R8[24]), .Y(n1068)
         );
  OAI221XL U374 ( .A0(n694), .A1(n1240), .B0(n728), .B1(n1221), .C0(n1067), 
        .Y(N145) );
  AOI22X1 U375 ( .A0(R9[25]), .A1(n1234), .B0(n1205), .B1(R8[25]), .Y(n1067)
         );
  OAI221XL U376 ( .A0(n693), .A1(n1239), .B0(n727), .B1(n1221), .C0(n1066), 
        .Y(N146) );
  AOI22X1 U377 ( .A0(R9[26]), .A1(n1226), .B0(n1198), .B1(R8[26]), .Y(n1066)
         );
  OAI221XL U378 ( .A0(n692), .A1(n1239), .B0(n726), .B1(n1220), .C0(n1065), 
        .Y(N147) );
  AOI22X1 U379 ( .A0(R9[27]), .A1(n1230), .B0(n1205), .B1(R8[27]), .Y(n1065)
         );
  OAI221XL U380 ( .A0(n691), .A1(n1239), .B0(n725), .B1(n1219), .C0(n1064), 
        .Y(N148) );
  AOI22X1 U381 ( .A0(R9[28]), .A1(n1229), .B0(n1201), .B1(R8[28]), .Y(n1064)
         );
  OAI221XL U382 ( .A0(n821), .A1(n1239), .B0(n787), .B1(n968), .C0(n1058), .Y(
        N154) );
  AOI22X1 U383 ( .A0(R13[0]), .A1(n1229), .B0(n1201), .B1(R12[0]), .Y(n1058)
         );
  OAI221XL U384 ( .A0(n820), .A1(n1239), .B0(n786), .B1(n1218), .C0(n1057), 
        .Y(N155) );
  AOI22X1 U385 ( .A0(R13[1]), .A1(n1229), .B0(n1201), .B1(R12[1]), .Y(n1057)
         );
  OAI221XL U386 ( .A0(n819), .A1(n1239), .B0(n785), .B1(n968), .C0(n1056), .Y(
        N156) );
  AOI22X1 U387 ( .A0(R13[2]), .A1(n1229), .B0(n1201), .B1(R12[2]), .Y(n1056)
         );
  OAI221XL U388 ( .A0(n818), .A1(n1239), .B0(n784), .B1(n968), .C0(n1055), .Y(
        N157) );
  AOI22X1 U389 ( .A0(R13[3]), .A1(n1229), .B0(n1201), .B1(R12[3]), .Y(n1055)
         );
  OAI221XL U390 ( .A0(n817), .A1(n1239), .B0(n783), .B1(n968), .C0(n1054), .Y(
        N158) );
  AOI22X1 U391 ( .A0(R13[4]), .A1(n1229), .B0(n1201), .B1(R12[4]), .Y(n1054)
         );
  OAI221XL U392 ( .A0(n816), .A1(n1236), .B0(n782), .B1(n968), .C0(n1053), .Y(
        N159) );
  AOI22X1 U393 ( .A0(R13[5]), .A1(n1229), .B0(n1201), .B1(R12[5]), .Y(n1053)
         );
  OAI221XL U394 ( .A0(n815), .A1(n1239), .B0(n781), .B1(n1224), .C0(n1052), 
        .Y(N160) );
  AOI22X1 U395 ( .A0(R13[6]), .A1(n1229), .B0(n1200), .B1(R12[6]), .Y(n1052)
         );
  OAI221XL U396 ( .A0(n814), .A1(n1238), .B0(n780), .B1(n1222), .C0(n1051), 
        .Y(N161) );
  AOI22X1 U397 ( .A0(R13[7]), .A1(n1229), .B0(n1199), .B1(R12[7]), .Y(n1051)
         );
  OAI221XL U398 ( .A0(n813), .A1(n1241), .B0(n779), .B1(n968), .C0(n1050), .Y(
        N162) );
  AOI22X1 U399 ( .A0(R13[8]), .A1(n1229), .B0(n1205), .B1(R12[8]), .Y(n1050)
         );
  OAI221XL U400 ( .A0(n812), .A1(n1240), .B0(n778), .B1(n968), .C0(n1049), .Y(
        N163) );
  AOI22X1 U401 ( .A0(R13[9]), .A1(n1229), .B0(n1200), .B1(R12[9]), .Y(n1049)
         );
  OAI221XL U402 ( .A0(n811), .A1(n1237), .B0(n777), .B1(n968), .C0(n1048), .Y(
        N164) );
  AOI22X1 U403 ( .A0(R13[10]), .A1(n1229), .B0(n1198), .B1(R12[10]), .Y(n1048)
         );
  OAI221XL U404 ( .A0(n810), .A1(n1237), .B0(n776), .B1(n1218), .C0(n1047), 
        .Y(N165) );
  AOI22X1 U405 ( .A0(R13[11]), .A1(n1230), .B0(n1198), .B1(R12[11]), .Y(n1047)
         );
  OAI221XL U406 ( .A0(n804), .A1(n1239), .B0(n770), .B1(n968), .C0(n1041), .Y(
        N171) );
  AOI22X1 U407 ( .A0(R13[17]), .A1(n1230), .B0(n1201), .B1(R12[17]), .Y(n1041)
         );
  OAI221XL U408 ( .A0(n803), .A1(n1235), .B0(n769), .B1(n1218), .C0(n1040), 
        .Y(N172) );
  AOI22X1 U409 ( .A0(R13[18]), .A1(n1230), .B0(n1202), .B1(R12[18]), .Y(n1040)
         );
  OAI221XL U410 ( .A0(n802), .A1(n1239), .B0(n768), .B1(n1224), .C0(n1039), 
        .Y(N173) );
  AOI22X1 U411 ( .A0(R13[19]), .A1(n1230), .B0(n1198), .B1(R12[19]), .Y(n1039)
         );
  OAI221XL U412 ( .A0(n801), .A1(n1240), .B0(n767), .B1(n1221), .C0(n1038), 
        .Y(N174) );
  AOI22X1 U413 ( .A0(R13[20]), .A1(n1230), .B0(n1199), .B1(R12[20]), .Y(n1038)
         );
  OAI221XL U414 ( .A0(n800), .A1(n1238), .B0(n766), .B1(n1220), .C0(n1037), 
        .Y(N175) );
  AOI22X1 U415 ( .A0(R13[21]), .A1(n1230), .B0(n1201), .B1(R12[21]), .Y(n1037)
         );
  OAI221XL U416 ( .A0(n799), .A1(n1241), .B0(n765), .B1(n1220), .C0(n1036), 
        .Y(N176) );
  AOI22X1 U417 ( .A0(R13[22]), .A1(n1230), .B0(n1202), .B1(R12[22]), .Y(n1036)
         );
  OAI221XL U418 ( .A0(n798), .A1(n963), .B0(n764), .B1(n1224), .C0(n1035), .Y(
        N177) );
  AOI22X1 U419 ( .A0(R13[23]), .A1(n1230), .B0(n1204), .B1(R12[23]), .Y(n1035)
         );
  OAI221XL U420 ( .A0(n797), .A1(n963), .B0(n763), .B1(n968), .C0(n1034), .Y(
        N178) );
  AOI22X1 U421 ( .A0(R13[24]), .A1(n1231), .B0(n1199), .B1(R12[24]), .Y(n1034)
         );
  OAI221XL U422 ( .A0(n796), .A1(n963), .B0(n762), .B1(n968), .C0(n1033), .Y(
        N179) );
  AOI22X1 U423 ( .A0(R13[25]), .A1(n1231), .B0(n1202), .B1(R12[25]), .Y(n1033)
         );
  OAI221XL U424 ( .A0(n795), .A1(n963), .B0(n761), .B1(n1220), .C0(n1032), .Y(
        N180) );
  AOI22X1 U425 ( .A0(R13[26]), .A1(n1231), .B0(n1198), .B1(R12[26]), .Y(n1032)
         );
  OAI221XL U426 ( .A0(n794), .A1(n963), .B0(n760), .B1(n1221), .C0(n1031), .Y(
        N181) );
  AOI22X1 U427 ( .A0(R13[27]), .A1(n1231), .B0(n1201), .B1(R12[27]), .Y(n1031)
         );
  INVX1 U428 ( .A(counter1[1]), .Y(n1248) );
  INVX1 U429 ( .A(counter1[0]), .Y(n1247) );
  INVX1 U430 ( .A(counter2[0]), .Y(n1249) );
  INVX1 U431 ( .A(reg_flag_mux), .Y(n1245) );
  OAI221XL U432 ( .A0(n793), .A1(n963), .B0(n759), .B1(n1218), .C0(n1030), .Y(
        N182) );
endmodule


module p_s ( clk, rst_n, data_in_3, p_s_flag_in, data_out_3 );
  input [135:0] data_in_3;
  output [33:0] data_out_3;
  input clk, rst_n, p_s_flag_in;
  wire   N26, N50, N52, N119, N120, N121, N122, N123, N124, N125, N126, N127,
         N128, N129, N130, N131, N132, N133, N134, N135, N136, N137, N138,
         N139, N140, N141, N142, N143, N144, N145, N146, N147, N148, N149,
         N150, N151, N152, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n862, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n883, n884, n885, n887, n888, n889, n890,
         n893, n895, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1, n3, n4, n6, n7, n10, n11, n12, n13, n14, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n59, n60, n186, n188, n190,
         n192, n194, n196, n198, n200, n202, n204, n206, n208, n249, n250,
         n251, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n583, n584, n858, n859, n860, n861, n863, n864, n865,
         n866, n867, n881, n882, n886, n891, n892, n894, n896, n1166, n1167,
         n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
         n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
         n1188, n1189, n1190, n1191, n1192, n1194, n1196, n1198, n1200, n1202,
         n1204, n1206, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
         n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
         n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
         n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
         n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
         n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
         n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
         n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283;
  wire   [1:0] counter_1;
  wire   [32:0] R0;
  wire   [33:0] R12;
  wire   [31:0] R1;
  wire   [33:0] R13;
  wire   [33:0] R2;
  wire   [33:0] R14;
  wire   [33:0] R3;
  wire   [32:0] R15;
  wire   [3:0] counter_2;

  AND2X2 U321 ( .A(n1158), .B(n870), .Y(n887) );
  AND2X2 U324 ( .A(counter_2[3]), .B(n862), .Y(n1158) );
  AND2X2 U326 ( .A(counter_2[3]), .B(counter_2[0]), .Y(n1159) );
  DFFXL R15_reg_13_ ( .D(n1208), .CK(clk), .Q(R15[13]) );
  DFFXL R14_reg_13_ ( .D(n1206), .CK(clk), .Q(R14[13]) );
  DFFXL R13_reg_13_ ( .D(n1204), .CK(clk), .Q(R13[13]) );
  DFFXL R12_reg_13_ ( .D(n1202), .CK(clk), .Q(R12[13]) );
  DFFXL R3_reg_29_ ( .D(n1200), .CK(clk), .Q(R3[29]) );
  DFFXL R2_reg_29_ ( .D(n1198), .CK(clk), .Q(R2[29]) );
  DFFXL R1_reg_29_ ( .D(n1196), .CK(clk), .Q(R1[29]) );
  DFFXL R0_reg_29_ ( .D(n1194), .CK(clk), .Q(R0[29]) );
  EDFFX1 R7_reg_22_ ( .D(data_in_3[56]), .E(n1265), .CK(clk), .QN(n597) );
  EDFFX1 R7_reg_21_ ( .D(data_in_3[55]), .E(n1265), .CK(clk), .QN(n598) );
  EDFFX1 R7_reg_20_ ( .D(data_in_3[54]), .E(n1265), .CK(clk), .QN(n599) );
  EDFFX1 R7_reg_19_ ( .D(data_in_3[53]), .E(n1265), .CK(clk), .QN(n600) );
  EDFFX1 R7_reg_18_ ( .D(data_in_3[52]), .E(n1265), .CK(clk), .QN(n601) );
  EDFFX1 R7_reg_10_ ( .D(data_in_3[44]), .E(n1264), .CK(clk), .QN(n609) );
  EDFFX1 R7_reg_9_ ( .D(data_in_3[43]), .E(n1264), .CK(clk), .QN(n610) );
  EDFFX1 R7_reg_6_ ( .D(data_in_3[40]), .E(n1264), .CK(clk), .QN(n613) );
  EDFFX1 R7_reg_5_ ( .D(data_in_3[39]), .E(n1261), .CK(clk), .QN(n614) );
  EDFFX1 R7_reg_4_ ( .D(data_in_3[38]), .E(n1261), .CK(clk), .QN(n615) );
  EDFFX1 R7_reg_3_ ( .D(data_in_3[37]), .E(n1260), .CK(clk), .QN(n616) );
  EDFFX1 R7_reg_2_ ( .D(data_in_3[36]), .E(n1261), .CK(clk), .QN(n617) );
  EDFFX1 R6_reg_22_ ( .D(data_in_3[56]), .E(n1276), .CK(clk), .QN(n665) );
  EDFFX1 R6_reg_21_ ( .D(data_in_3[55]), .E(n1276), .CK(clk), .QN(n666) );
  EDFFX1 R6_reg_20_ ( .D(data_in_3[54]), .E(n1276), .CK(clk), .QN(n667) );
  EDFFX1 R6_reg_19_ ( .D(data_in_3[53]), .E(n1276), .CK(clk), .QN(n668) );
  EDFFX1 R6_reg_18_ ( .D(data_in_3[52]), .E(n1276), .CK(clk), .QN(n669) );
  EDFFX1 R6_reg_10_ ( .D(data_in_3[44]), .E(n1269), .CK(clk), .QN(n677) );
  EDFFX1 R6_reg_9_ ( .D(data_in_3[43]), .E(n1276), .CK(clk), .QN(n678) );
  EDFFX1 R6_reg_6_ ( .D(data_in_3[40]), .E(n1269), .CK(clk), .QN(n681) );
  EDFFX1 R6_reg_5_ ( .D(data_in_3[39]), .E(n1273), .CK(clk), .QN(n682) );
  EDFFX1 R6_reg_4_ ( .D(data_in_3[38]), .E(n1275), .CK(clk), .QN(n683) );
  EDFFX1 R6_reg_3_ ( .D(data_in_3[37]), .E(n1276), .CK(clk), .QN(n684) );
  EDFFX1 R6_reg_2_ ( .D(data_in_3[36]), .E(n1272), .CK(clk), .QN(n685) );
  EDFFX1 R4_reg_22_ ( .D(data_in_3[56]), .E(n1213), .CK(clk), .QN(n733) );
  EDFFX1 R4_reg_21_ ( .D(data_in_3[55]), .E(n1213), .CK(clk), .QN(n734) );
  EDFFX1 R4_reg_20_ ( .D(data_in_3[54]), .E(n1213), .CK(clk), .QN(n735) );
  EDFFX1 R4_reg_19_ ( .D(data_in_3[53]), .E(n1213), .CK(clk), .QN(n736) );
  EDFFX1 R4_reg_18_ ( .D(data_in_3[52]), .E(n1213), .CK(clk), .QN(n737) );
  EDFFX1 R4_reg_10_ ( .D(data_in_3[44]), .E(n1212), .CK(clk), .QN(n745) );
  EDFFX1 R4_reg_9_ ( .D(data_in_3[43]), .E(n1210), .CK(clk), .QN(n746) );
  EDFFX1 R4_reg_6_ ( .D(data_in_3[40]), .E(n1212), .CK(clk), .QN(n749) );
  EDFFX1 R4_reg_5_ ( .D(data_in_3[39]), .E(n1215), .CK(clk), .QN(n750) );
  EDFFX1 R4_reg_4_ ( .D(data_in_3[38]), .E(n1213), .CK(clk), .QN(n751) );
  EDFFX1 R4_reg_3_ ( .D(data_in_3[37]), .E(n1213), .CK(clk), .QN(n752) );
  EDFFX1 R4_reg_2_ ( .D(data_in_3[36]), .E(n1212), .CK(clk), .QN(n753) );
  EDFFXL R5_reg_29_ ( .D(data_in_3[63]), .E(n1221), .CK(clk), .QN(n794) );
  EDFFXL R5_reg_28_ ( .D(data_in_3[62]), .E(n1220), .CK(clk), .QN(n795) );
  EDFFXL R5_reg_27_ ( .D(data_in_3[61]), .E(n1221), .CK(clk), .QN(n796) );
  EDFFXL R5_reg_26_ ( .D(data_in_3[60]), .E(n1221), .CK(clk), .QN(n797) );
  EDFFXL R5_reg_25_ ( .D(data_in_3[59]), .E(n1221), .CK(clk), .QN(n798) );
  EDFFXL R5_reg_24_ ( .D(data_in_3[58]), .E(n1221), .CK(clk), .QN(n799) );
  EDFFXL R5_reg_23_ ( .D(data_in_3[57]), .E(n1221), .CK(clk), .QN(n800) );
  EDFFXL R5_reg_22_ ( .D(data_in_3[56]), .E(n1221), .CK(clk), .QN(n801) );
  EDFFXL R5_reg_21_ ( .D(data_in_3[55]), .E(n1221), .CK(clk), .QN(n802) );
  EDFFXL R5_reg_20_ ( .D(data_in_3[54]), .E(n1221), .CK(clk), .QN(n803) );
  EDFFXL R5_reg_19_ ( .D(data_in_3[53]), .E(n1221), .CK(clk), .QN(n804) );
  EDFFXL R5_reg_18_ ( .D(data_in_3[52]), .E(n1221), .CK(clk), .QN(n805) );
  EDFFXL R5_reg_11_ ( .D(data_in_3[45]), .E(n1220), .CK(clk), .QN(n812) );
  EDFFXL R5_reg_10_ ( .D(data_in_3[44]), .E(n1220), .CK(clk), .QN(n813) );
  EDFFXL R5_reg_9_ ( .D(data_in_3[43]), .E(n1220), .CK(clk), .QN(n814) );
  EDFFXL R5_reg_8_ ( .D(data_in_3[42]), .E(n1220), .CK(clk), .QN(n815) );
  EDFFXL R5_reg_7_ ( .D(data_in_3[41]), .E(n1220), .CK(clk), .QN(n816) );
  EDFFXL R5_reg_6_ ( .D(data_in_3[40]), .E(n1220), .CK(clk), .QN(n817) );
  EDFFXL R5_reg_5_ ( .D(data_in_3[39]), .E(n1220), .CK(clk), .QN(n818) );
  EDFFXL R5_reg_4_ ( .D(data_in_3[38]), .E(n1220), .CK(clk), .QN(n819) );
  EDFFXL R5_reg_3_ ( .D(data_in_3[37]), .E(n1223), .CK(clk), .QN(n820) );
  EDFFXL R5_reg_2_ ( .D(data_in_3[36]), .E(n1223), .CK(clk), .QN(n821) );
  EDFFXL R5_reg_1_ ( .D(data_in_3[35]), .E(n1223), .CK(clk), .QN(n822) );
  EDFFXL R10_reg_28_ ( .D(data_in_3[96]), .E(n1270), .CK(clk), .QN(n625) );
  EDFFXL R10_reg_27_ ( .D(data_in_3[95]), .E(n1270), .CK(clk), .QN(n626) );
  EDFFXL R10_reg_26_ ( .D(data_in_3[94]), .E(n1270), .CK(clk), .QN(n627) );
  EDFFXL R10_reg_25_ ( .D(data_in_3[93]), .E(n1270), .CK(clk), .QN(n628) );
  EDFFXL R10_reg_24_ ( .D(data_in_3[92]), .E(n1270), .CK(clk), .QN(n629) );
  EDFFXL R10_reg_23_ ( .D(data_in_3[91]), .E(n1270), .CK(clk), .QN(n630) );
  EDFFXL R10_reg_22_ ( .D(data_in_3[90]), .E(n1270), .CK(clk), .QN(n631) );
  EDFFXL R10_reg_21_ ( .D(data_in_3[89]), .E(n1270), .CK(clk), .QN(n632) );
  EDFFXL R10_reg_20_ ( .D(data_in_3[88]), .E(n1270), .CK(clk), .QN(n633) );
  EDFFXL R10_reg_19_ ( .D(data_in_3[87]), .E(n1270), .CK(clk), .QN(n634) );
  EDFFXL R10_reg_18_ ( .D(data_in_3[86]), .E(n1270), .CK(clk), .QN(n635) );
  EDFFXL R10_reg_11_ ( .D(data_in_3[79]), .E(n1269), .CK(clk), .QN(n642) );
  EDFFXL R10_reg_10_ ( .D(data_in_3[78]), .E(n1269), .CK(clk), .QN(n643) );
  EDFFXL R10_reg_8_ ( .D(data_in_3[76]), .E(n1269), .CK(clk), .QN(n645) );
  EDFFXL R10_reg_7_ ( .D(data_in_3[75]), .E(n1269), .CK(clk), .QN(n646) );
  EDFFXL R10_reg_6_ ( .D(data_in_3[74]), .E(n1269), .CK(clk), .QN(n647) );
  EDFFXL R10_reg_5_ ( .D(data_in_3[73]), .E(n1269), .CK(clk), .QN(n648) );
  EDFFXL R10_reg_4_ ( .D(data_in_3[72]), .E(n1269), .CK(clk), .QN(n649) );
  EDFFXL R10_reg_3_ ( .D(data_in_3[71]), .E(n1269), .CK(clk), .QN(n650) );
  EDFFXL R10_reg_2_ ( .D(data_in_3[70]), .E(n1269), .CK(clk), .QN(n651) );
  EDFFXL R10_reg_1_ ( .D(data_in_3[69]), .E(n1272), .CK(clk), .QN(n652) );
  EDFFXL R11_reg_28_ ( .D(data_in_3[96]), .E(n1261), .CK(clk), .QN(n693) );
  EDFFXL R11_reg_27_ ( .D(data_in_3[95]), .E(n1261), .CK(clk), .QN(n694) );
  EDFFXL R11_reg_26_ ( .D(data_in_3[94]), .E(n1261), .CK(clk), .QN(n695) );
  EDFFXL R11_reg_25_ ( .D(data_in_3[93]), .E(n1260), .CK(clk), .QN(n696) );
  EDFFXL R11_reg_24_ ( .D(data_in_3[92]), .E(n1258), .CK(clk), .QN(n697) );
  EDFFXL R11_reg_23_ ( .D(data_in_3[91]), .E(n1264), .CK(clk), .QN(n698) );
  EDFFXL R11_reg_22_ ( .D(data_in_3[90]), .E(n1260), .CK(clk), .QN(n699) );
  EDFFXL R11_reg_21_ ( .D(data_in_3[89]), .E(n1264), .CK(clk), .QN(n700) );
  EDFFXL R11_reg_20_ ( .D(data_in_3[88]), .E(n1259), .CK(clk), .QN(n701) );
  EDFFXL R11_reg_19_ ( .D(data_in_3[87]), .E(n1264), .CK(clk), .QN(n702) );
  EDFFXL R11_reg_18_ ( .D(data_in_3[86]), .E(n1260), .CK(clk), .QN(n703) );
  EDFFXL R11_reg_11_ ( .D(data_in_3[79]), .E(n1259), .CK(clk), .QN(n710) );
  EDFFXL R11_reg_10_ ( .D(data_in_3[78]), .E(n1261), .CK(clk), .QN(n711) );
  EDFFXL R11_reg_8_ ( .D(data_in_3[76]), .E(n1258), .CK(clk), .QN(n713) );
  EDFFXL R11_reg_7_ ( .D(data_in_3[75]), .E(n1259), .CK(clk), .QN(n714) );
  EDFFXL R11_reg_6_ ( .D(data_in_3[74]), .E(n1264), .CK(clk), .QN(n715) );
  EDFFXL R11_reg_5_ ( .D(data_in_3[73]), .E(n1258), .CK(clk), .QN(n716) );
  EDFFXL R11_reg_4_ ( .D(data_in_3[72]), .E(n1264), .CK(clk), .QN(n717) );
  EDFFXL R11_reg_3_ ( .D(data_in_3[71]), .E(n1264), .CK(clk), .QN(n718) );
  EDFFXL R11_reg_2_ ( .D(data_in_3[70]), .E(n1264), .CK(clk), .QN(n719) );
  EDFFXL R11_reg_1_ ( .D(data_in_3[69]), .E(n1260), .CK(clk), .QN(n720) );
  EDFFXL R8_reg_28_ ( .D(data_in_3[96]), .E(n1213), .CK(clk), .QN(n761) );
  EDFFXL R8_reg_27_ ( .D(data_in_3[95]), .E(n1212), .CK(clk), .QN(n762) );
  EDFFXL R8_reg_26_ ( .D(data_in_3[94]), .E(n1213), .CK(clk), .QN(n763) );
  EDFFXL R8_reg_25_ ( .D(data_in_3[93]), .E(n1212), .CK(clk), .QN(n764) );
  EDFFXL R8_reg_24_ ( .D(data_in_3[92]), .E(n1212), .CK(clk), .QN(n765) );
  EDFFXL R8_reg_23_ ( .D(data_in_3[91]), .E(n1212), .CK(clk), .QN(n766) );
  EDFFXL R8_reg_22_ ( .D(data_in_3[90]), .E(n1212), .CK(clk), .QN(n767) );
  EDFFXL R8_reg_21_ ( .D(data_in_3[89]), .E(n1212), .CK(clk), .QN(n768) );
  EDFFXL R8_reg_20_ ( .D(data_in_3[88]), .E(n1212), .CK(clk), .QN(n769) );
  EDFFXL R8_reg_19_ ( .D(data_in_3[87]), .E(n1212), .CK(clk), .QN(n770) );
  EDFFXL R8_reg_18_ ( .D(data_in_3[86]), .E(n1212), .CK(clk), .QN(n771) );
  EDFFXL R8_reg_11_ ( .D(data_in_3[79]), .E(n1211), .CK(clk), .QN(n778) );
  EDFFXL R8_reg_10_ ( .D(data_in_3[78]), .E(n1210), .CK(clk), .QN(n779) );
  EDFFXL R8_reg_8_ ( .D(data_in_3[76]), .E(n1212), .CK(clk), .QN(n781) );
  EDFFXL R8_reg_7_ ( .D(data_in_3[75]), .E(n1214), .CK(clk), .QN(n782) );
  EDFFXL R8_reg_6_ ( .D(data_in_3[74]), .E(n1209), .CK(clk), .QN(n783) );
  EDFFXL R8_reg_5_ ( .D(data_in_3[73]), .E(n1215), .CK(clk), .QN(n784) );
  EDFFXL R8_reg_4_ ( .D(data_in_3[72]), .E(n1209), .CK(clk), .QN(n785) );
  EDFFXL R8_reg_3_ ( .D(data_in_3[71]), .E(n1211), .CK(clk), .QN(n786) );
  EDFFXL R8_reg_2_ ( .D(data_in_3[70]), .E(n1215), .CK(clk), .QN(n787) );
  EDFFXL R8_reg_1_ ( .D(data_in_3[69]), .E(n1211), .CK(clk), .QN(n788) );
  EDFFXL R9_reg_28_ ( .D(data_in_3[96]), .E(n1220), .CK(clk), .QN(n829) );
  EDFFXL R9_reg_27_ ( .D(data_in_3[95]), .E(n1223), .CK(clk), .QN(n830) );
  EDFFXL R9_reg_26_ ( .D(data_in_3[94]), .E(n1223), .CK(clk), .QN(n831) );
  EDFFXL R9_reg_25_ ( .D(data_in_3[93]), .E(n249), .CK(clk), .QN(n832) );
  EDFFXL R9_reg_24_ ( .D(data_in_3[92]), .E(n249), .CK(clk), .QN(n833) );
  EDFFXL R9_reg_23_ ( .D(data_in_3[91]), .E(n1219), .CK(clk), .QN(n834) );
  EDFFXL R9_reg_22_ ( .D(data_in_3[90]), .E(n1223), .CK(clk), .QN(n835) );
  EDFFXL R9_reg_21_ ( .D(data_in_3[89]), .E(n1217), .CK(clk), .QN(n836) );
  EDFFXL R9_reg_20_ ( .D(data_in_3[88]), .E(n1221), .CK(clk), .QN(n837) );
  EDFFXL R9_reg_19_ ( .D(data_in_3[87]), .E(n249), .CK(clk), .QN(n838) );
  EDFFXL R9_reg_18_ ( .D(data_in_3[86]), .E(n1222), .CK(clk), .QN(n839) );
  EDFFXL R9_reg_11_ ( .D(data_in_3[79]), .E(n1223), .CK(clk), .QN(n846) );
  EDFFXL R9_reg_10_ ( .D(data_in_3[78]), .E(n1217), .CK(clk), .QN(n847) );
  EDFFXL R9_reg_8_ ( .D(data_in_3[76]), .E(n1222), .CK(clk), .QN(n849) );
  EDFFXL R9_reg_7_ ( .D(data_in_3[75]), .E(n1220), .CK(clk), .QN(n850) );
  EDFFXL R9_reg_6_ ( .D(data_in_3[74]), .E(n1223), .CK(clk), .QN(n851) );
  EDFFXL R9_reg_5_ ( .D(data_in_3[73]), .E(n1221), .CK(clk), .QN(n852) );
  EDFFXL R9_reg_4_ ( .D(data_in_3[72]), .E(n1217), .CK(clk), .QN(n853) );
  EDFFXL R9_reg_3_ ( .D(data_in_3[71]), .E(n1221), .CK(clk), .QN(n854) );
  EDFFXL R9_reg_2_ ( .D(data_in_3[70]), .E(n1220), .CK(clk), .QN(n855) );
  EDFFXL R9_reg_1_ ( .D(data_in_3[69]), .E(n1219), .CK(clk), .QN(n856) );
  EDFFXL R15_reg_29_ ( .D(data_in_3[131]), .E(n1260), .CK(clk), .Q(R15[29]) );
  EDFFXL R15_reg_28_ ( .D(data_in_3[130]), .E(n1260), .CK(clk), .Q(R15[28]) );
  EDFFXL R15_reg_27_ ( .D(data_in_3[129]), .E(n1260), .CK(clk), .Q(R15[27]) );
  EDFFXL R15_reg_26_ ( .D(data_in_3[128]), .E(n1260), .CK(clk), .Q(R15[26]) );
  EDFFXL R15_reg_25_ ( .D(data_in_3[127]), .E(n1260), .CK(clk), .Q(R15[25]) );
  EDFFXL R15_reg_24_ ( .D(data_in_3[126]), .E(n1260), .CK(clk), .Q(R15[24]) );
  EDFFXL R15_reg_23_ ( .D(data_in_3[125]), .E(n1259), .CK(clk), .Q(R15[23]) );
  EDFFXL R15_reg_22_ ( .D(data_in_3[124]), .E(n1259), .CK(clk), .Q(R15[22]) );
  EDFFXL R15_reg_21_ ( .D(data_in_3[123]), .E(n1259), .CK(clk), .Q(R15[21]) );
  EDFFXL R15_reg_20_ ( .D(data_in_3[122]), .E(n1259), .CK(clk), .Q(R15[20]) );
  EDFFXL R15_reg_19_ ( .D(data_in_3[121]), .E(n1259), .CK(clk), .Q(R15[19]) );
  EDFFXL R15_reg_11_ ( .D(data_in_3[113]), .E(n1258), .CK(clk), .Q(R15[11]) );
  EDFFXL R15_reg_10_ ( .D(data_in_3[112]), .E(n1258), .CK(clk), .Q(R15[10]) );
  EDFFXL R15_reg_9_ ( .D(data_in_3[111]), .E(n1258), .CK(clk), .Q(R15[9]) );
  EDFFXL R15_reg_8_ ( .D(data_in_3[110]), .E(n1258), .CK(clk), .Q(R15[8]) );
  EDFFXL R15_reg_7_ ( .D(data_in_3[109]), .E(n1258), .CK(clk), .Q(R15[7]) );
  EDFFXL R15_reg_6_ ( .D(data_in_3[108]), .E(n1258), .CK(clk), .Q(R15[6]) );
  EDFFXL R15_reg_5_ ( .D(data_in_3[107]), .E(n1258), .CK(clk), .Q(R15[5]) );
  EDFFXL R15_reg_4_ ( .D(data_in_3[106]), .E(n1258), .CK(clk), .Q(R15[4]) );
  EDFFXL R15_reg_3_ ( .D(data_in_3[105]), .E(n1258), .CK(clk), .Q(R15[3]) );
  EDFFXL R15_reg_2_ ( .D(data_in_3[104]), .E(n1258), .CK(clk), .Q(R15[2]) );
  EDFFXL R12_reg_29_ ( .D(data_in_3[131]), .E(n1211), .CK(clk), .Q(R12[29]) );
  EDFFXL R12_reg_28_ ( .D(data_in_3[130]), .E(n1211), .CK(clk), .Q(R12[28]) );
  EDFFXL R12_reg_27_ ( .D(data_in_3[129]), .E(n1211), .CK(clk), .Q(R12[27]) );
  EDFFXL R12_reg_26_ ( .D(data_in_3[128]), .E(n1211), .CK(clk), .Q(R12[26]) );
  EDFFXL R12_reg_25_ ( .D(data_in_3[127]), .E(n1211), .CK(clk), .Q(R12[25]) );
  EDFFXL R12_reg_24_ ( .D(data_in_3[126]), .E(n1211), .CK(clk), .Q(R12[24]) );
  EDFFXL R12_reg_23_ ( .D(data_in_3[125]), .E(n1210), .CK(clk), .Q(R12[23]) );
  EDFFXL R12_reg_22_ ( .D(data_in_3[124]), .E(n1210), .CK(clk), .Q(R12[22]) );
  EDFFXL R12_reg_21_ ( .D(data_in_3[123]), .E(n1210), .CK(clk), .Q(R12[21]) );
  EDFFXL R12_reg_20_ ( .D(data_in_3[122]), .E(n1210), .CK(clk), .Q(R12[20]) );
  EDFFXL R12_reg_19_ ( .D(data_in_3[121]), .E(n1210), .CK(clk), .Q(R12[19]) );
  EDFFXL R12_reg_11_ ( .D(data_in_3[113]), .E(n1209), .CK(clk), .Q(R12[11]) );
  EDFFXL R12_reg_10_ ( .D(data_in_3[112]), .E(n1209), .CK(clk), .Q(R12[10]) );
  EDFFXL R12_reg_9_ ( .D(data_in_3[111]), .E(n1209), .CK(clk), .Q(R12[9]) );
  EDFFXL R12_reg_8_ ( .D(data_in_3[110]), .E(n1209), .CK(clk), .Q(R12[8]) );
  EDFFXL R12_reg_7_ ( .D(data_in_3[109]), .E(n1209), .CK(clk), .Q(R12[7]) );
  EDFFXL R12_reg_6_ ( .D(data_in_3[108]), .E(n1209), .CK(clk), .Q(R12[6]) );
  EDFFXL R12_reg_5_ ( .D(data_in_3[107]), .E(n1209), .CK(clk), .Q(R12[5]) );
  EDFFXL R12_reg_4_ ( .D(data_in_3[106]), .E(n1209), .CK(clk), .Q(R12[4]) );
  EDFFXL R12_reg_3_ ( .D(data_in_3[105]), .E(n1209), .CK(clk), .Q(R12[3]) );
  EDFFXL R12_reg_2_ ( .D(data_in_3[104]), .E(n1209), .CK(clk), .Q(R12[2]) );
  EDFFXL R3_reg_28_ ( .D(data_in_3[28]), .E(n1264), .CK(clk), .Q(R3[28]) );
  EDFFXL R3_reg_27_ ( .D(data_in_3[27]), .E(n1263), .CK(clk), .Q(R3[27]) );
  EDFFXL R3_reg_24_ ( .D(data_in_3[24]), .E(n1263), .CK(clk), .Q(R3[24]) );
  EDFFXL R3_reg_23_ ( .D(data_in_3[23]), .E(n1263), .CK(clk), .Q(R3[23]) );
  EDFFXL R3_reg_22_ ( .D(data_in_3[22]), .E(n1263), .CK(clk), .Q(R3[22]) );
  EDFFXL R3_reg_21_ ( .D(data_in_3[21]), .E(n1263), .CK(clk), .Q(R3[21]) );
  EDFFXL R3_reg_20_ ( .D(data_in_3[20]), .E(n1263), .CK(clk), .Q(R3[20]) );
  EDFFXL R3_reg_19_ ( .D(data_in_3[19]), .E(n1263), .CK(clk), .Q(R3[19]) );
  EDFFXL R3_reg_18_ ( .D(data_in_3[18]), .E(n1263), .CK(clk), .Q(R3[18]) );
  EDFFXL R3_reg_11_ ( .D(data_in_3[11]), .E(n1262), .CK(clk), .Q(R3[11]) );
  EDFFXL R3_reg_10_ ( .D(data_in_3[10]), .E(n1262), .CK(clk), .Q(R3[10]) );
  EDFFXL R3_reg_9_ ( .D(data_in_3[9]), .E(n1262), .CK(clk), .Q(R3[9]) );
  EDFFXL R3_reg_8_ ( .D(data_in_3[8]), .E(n1262), .CK(clk), .Q(R3[8]) );
  EDFFXL R3_reg_7_ ( .D(data_in_3[7]), .E(n1262), .CK(clk), .Q(R3[7]) );
  EDFFXL R3_reg_5_ ( .D(data_in_3[5]), .E(n1262), .CK(clk), .Q(R3[5]) );
  EDFFXL R3_reg_4_ ( .D(data_in_3[4]), .E(n1262), .CK(clk), .Q(R3[4]) );
  EDFFXL R3_reg_3_ ( .D(data_in_3[3]), .E(n1261), .CK(clk), .Q(R3[3]) );
  EDFFXL R3_reg_2_ ( .D(data_in_3[2]), .E(n1261), .CK(clk), .Q(R3[2]) );
  EDFFXL R3_reg_1_ ( .D(data_in_3[1]), .E(n1261), .CK(clk), .Q(R3[1]) );
  EDFFX1 R3_reg_0_ ( .D(data_in_3[0]), .E(n1261), .CK(clk), .Q(R3[0]) );
  EDFFXL R0_reg_28_ ( .D(data_in_3[28]), .E(n250), .CK(clk), .Q(R0[28]) );
  EDFFXL R0_reg_27_ ( .D(data_in_3[27]), .E(n250), .CK(clk), .Q(R0[27]) );
  EDFFXL R0_reg_24_ ( .D(data_in_3[24]), .E(n250), .CK(clk), .Q(R0[24]) );
  EDFFXL R0_reg_23_ ( .D(data_in_3[23]), .E(n250), .CK(clk), .Q(R0[23]) );
  EDFFXL R0_reg_22_ ( .D(data_in_3[22]), .E(n1213), .CK(clk), .Q(R0[22]) );
  EDFFXL R0_reg_21_ ( .D(data_in_3[21]), .E(n1210), .CK(clk), .Q(R0[21]) );
  EDFFXL R0_reg_20_ ( .D(data_in_3[20]), .E(n1214), .CK(clk), .Q(R0[20]) );
  EDFFXL R0_reg_19_ ( .D(data_in_3[19]), .E(n1215), .CK(clk), .Q(R0[19]) );
  EDFFXL R0_reg_18_ ( .D(data_in_3[18]), .E(n1212), .CK(clk), .Q(R0[18]) );
  EDFFXL R0_reg_11_ ( .D(data_in_3[11]), .E(n1214), .CK(clk), .Q(R0[11]) );
  EDFFXL R0_reg_10_ ( .D(data_in_3[10]), .E(n1214), .CK(clk), .Q(R0[10]) );
  EDFFXL R0_reg_9_ ( .D(data_in_3[9]), .E(n1214), .CK(clk), .Q(R0[9]) );
  EDFFXL R0_reg_8_ ( .D(data_in_3[8]), .E(n1214), .CK(clk), .Q(R0[8]) );
  EDFFXL R0_reg_7_ ( .D(data_in_3[7]), .E(n1214), .CK(clk), .Q(R0[7]) );
  EDFFXL R0_reg_5_ ( .D(data_in_3[5]), .E(n1215), .CK(clk), .Q(R0[5]) );
  EDFFXL R0_reg_4_ ( .D(data_in_3[4]), .E(n1211), .CK(clk), .Q(R0[4]) );
  EDFFXL R0_reg_3_ ( .D(data_in_3[3]), .E(n1215), .CK(clk), .Q(R0[3]) );
  EDFFXL R0_reg_2_ ( .D(data_in_3[2]), .E(n1215), .CK(clk), .Q(R0[2]) );
  EDFFXL R0_reg_1_ ( .D(data_in_3[1]), .E(n1209), .CK(clk), .Q(R0[1]) );
  EDFFX1 R0_reg_0_ ( .D(data_in_3[0]), .E(n1215), .CK(clk), .Q(R0[0]) );
  EDFFXL R1_reg_28_ ( .D(data_in_3[28]), .E(n1222), .CK(clk), .Q(R1[28]) );
  EDFFXL R1_reg_27_ ( .D(data_in_3[27]), .E(n1223), .CK(clk), .Q(R1[27]) );
  EDFFXL R1_reg_24_ ( .D(data_in_3[24]), .E(n1218), .CK(clk), .Q(R1[24]) );
  EDFFXL R1_reg_23_ ( .D(data_in_3[23]), .E(n1219), .CK(clk), .Q(R1[23]) );
  EDFFXL R1_reg_22_ ( .D(data_in_3[22]), .E(n1222), .CK(clk), .Q(R1[22]) );
  EDFFXL R1_reg_21_ ( .D(data_in_3[21]), .E(n1223), .CK(clk), .Q(R1[21]) );
  EDFFXL R1_reg_20_ ( .D(data_in_3[20]), .E(n249), .CK(clk), .Q(R1[20]) );
  EDFFXL R1_reg_19_ ( .D(data_in_3[19]), .E(n249), .CK(clk), .Q(R1[19]) );
  EDFFXL R1_reg_18_ ( .D(data_in_3[18]), .E(n1220), .CK(clk), .Q(R1[18]) );
  EDFFXL R1_reg_11_ ( .D(data_in_3[11]), .E(n1222), .CK(clk), .Q(R1[11]) );
  EDFFXL R1_reg_10_ ( .D(data_in_3[10]), .E(n1222), .CK(clk), .Q(R1[10]) );
  EDFFXL R1_reg_9_ ( .D(data_in_3[9]), .E(n1222), .CK(clk), .Q(R1[9]) );
  EDFFXL R1_reg_8_ ( .D(data_in_3[8]), .E(n1222), .CK(clk), .Q(R1[8]) );
  EDFFXL R1_reg_7_ ( .D(data_in_3[7]), .E(n1222), .CK(clk), .Q(R1[7]) );
  EDFFXL R1_reg_5_ ( .D(data_in_3[5]), .E(n1220), .CK(clk), .Q(R1[5]) );
  EDFFXL R1_reg_4_ ( .D(data_in_3[4]), .E(n1220), .CK(clk), .Q(R1[4]) );
  EDFFXL R1_reg_3_ ( .D(data_in_3[3]), .E(n1217), .CK(clk), .Q(R1[3]) );
  EDFFXL R1_reg_2_ ( .D(data_in_3[2]), .E(n1221), .CK(clk), .Q(R1[2]) );
  EDFFXL R1_reg_1_ ( .D(data_in_3[1]), .E(n1220), .CK(clk), .Q(R1[1]) );
  EDFFX1 R1_reg_0_ ( .D(data_in_3[0]), .E(n1218), .CK(clk), .Q(R1[0]) );
  EDFFXL R14_reg_29_ ( .D(data_in_3[131]), .E(n1273), .CK(clk), .Q(R14[29]) );
  EDFFXL R14_reg_28_ ( .D(data_in_3[130]), .E(n1273), .CK(clk), .Q(R14[28]) );
  EDFFXL R14_reg_27_ ( .D(data_in_3[129]), .E(n1272), .CK(clk), .Q(R14[27]) );
  EDFFXL R14_reg_26_ ( .D(data_in_3[128]), .E(n1272), .CK(clk), .Q(R14[26]) );
  EDFFXL R14_reg_25_ ( .D(data_in_3[127]), .E(n1272), .CK(clk), .Q(R14[25]) );
  EDFFXL R14_reg_24_ ( .D(data_in_3[126]), .E(n1272), .CK(clk), .Q(R14[24]) );
  EDFFXL R14_reg_23_ ( .D(data_in_3[125]), .E(n1272), .CK(clk), .Q(R14[23]) );
  EDFFXL R14_reg_22_ ( .D(data_in_3[124]), .E(n1272), .CK(clk), .Q(R14[22]) );
  EDFFXL R14_reg_21_ ( .D(data_in_3[123]), .E(n1272), .CK(clk), .Q(R14[21]) );
  EDFFXL R14_reg_20_ ( .D(data_in_3[122]), .E(n1272), .CK(clk), .Q(R14[20]) );
  EDFFXL R14_reg_19_ ( .D(data_in_3[121]), .E(n1272), .CK(clk), .Q(R14[19]) );
  EDFFXL R14_reg_11_ ( .D(data_in_3[113]), .E(n1271), .CK(clk), .Q(R14[11]) );
  EDFFXL R14_reg_10_ ( .D(data_in_3[112]), .E(n1271), .CK(clk), .Q(R14[10]) );
  EDFFXL R14_reg_9_ ( .D(data_in_3[111]), .E(n1271), .CK(clk), .Q(R14[9]) );
  EDFFXL R14_reg_8_ ( .D(data_in_3[110]), .E(n1271), .CK(clk), .Q(R14[8]) );
  EDFFXL R14_reg_7_ ( .D(data_in_3[109]), .E(n1271), .CK(clk), .Q(R14[7]) );
  EDFFXL R14_reg_6_ ( .D(data_in_3[108]), .E(n1271), .CK(clk), .Q(R14[6]) );
  EDFFXL R14_reg_5_ ( .D(data_in_3[107]), .E(n1271), .CK(clk), .Q(R14[5]) );
  EDFFXL R14_reg_4_ ( .D(data_in_3[106]), .E(n1271), .CK(clk), .Q(R14[4]) );
  EDFFXL R14_reg_3_ ( .D(data_in_3[105]), .E(n1270), .CK(clk), .Q(R14[3]) );
  EDFFXL R14_reg_2_ ( .D(data_in_3[104]), .E(n1270), .CK(clk), .Q(R14[2]) );
  EDFFXL R13_reg_29_ ( .D(data_in_3[131]), .E(n1219), .CK(clk), .Q(R13[29]) );
  EDFFXL R13_reg_28_ ( .D(data_in_3[130]), .E(n1219), .CK(clk), .Q(R13[28]) );
  EDFFXL R13_reg_27_ ( .D(data_in_3[129]), .E(n1219), .CK(clk), .Q(R13[27]) );
  EDFFXL R13_reg_26_ ( .D(data_in_3[128]), .E(n1219), .CK(clk), .Q(R13[26]) );
  EDFFXL R13_reg_25_ ( .D(data_in_3[127]), .E(n1219), .CK(clk), .Q(R13[25]) );
  EDFFXL R13_reg_24_ ( .D(data_in_3[126]), .E(n1219), .CK(clk), .Q(R13[24]) );
  EDFFXL R13_reg_23_ ( .D(data_in_3[125]), .E(n1218), .CK(clk), .Q(R13[23]) );
  EDFFXL R13_reg_22_ ( .D(data_in_3[124]), .E(n1218), .CK(clk), .Q(R13[22]) );
  EDFFXL R13_reg_21_ ( .D(data_in_3[123]), .E(n1218), .CK(clk), .Q(R13[21]) );
  EDFFXL R13_reg_20_ ( .D(data_in_3[122]), .E(n1218), .CK(clk), .Q(R13[20]) );
  EDFFXL R13_reg_19_ ( .D(data_in_3[121]), .E(n1218), .CK(clk), .Q(R13[19]) );
  EDFFXL R13_reg_11_ ( .D(data_in_3[113]), .E(n1217), .CK(clk), .Q(R13[11]) );
  EDFFXL R13_reg_10_ ( .D(data_in_3[112]), .E(n1217), .CK(clk), .Q(R13[10]) );
  EDFFXL R13_reg_9_ ( .D(data_in_3[111]), .E(n1217), .CK(clk), .Q(R13[9]) );
  EDFFXL R13_reg_8_ ( .D(data_in_3[110]), .E(n1217), .CK(clk), .Q(R13[8]) );
  EDFFXL R13_reg_7_ ( .D(data_in_3[109]), .E(n1217), .CK(clk), .Q(R13[7]) );
  EDFFXL R13_reg_6_ ( .D(data_in_3[108]), .E(n1217), .CK(clk), .Q(R13[6]) );
  EDFFXL R13_reg_5_ ( .D(data_in_3[107]), .E(n1217), .CK(clk), .Q(R13[5]) );
  EDFFXL R13_reg_4_ ( .D(data_in_3[106]), .E(n1217), .CK(clk), .Q(R13[4]) );
  EDFFXL R13_reg_3_ ( .D(data_in_3[105]), .E(n1217), .CK(clk), .Q(R13[3]) );
  EDFFXL R13_reg_2_ ( .D(data_in_3[104]), .E(n1217), .CK(clk), .Q(R13[2]) );
  EDFFXL R2_reg_28_ ( .D(data_in_3[28]), .E(n1275), .CK(clk), .Q(R2[28]) );
  EDFFXL R2_reg_27_ ( .D(data_in_3[27]), .E(n1275), .CK(clk), .Q(R2[27]) );
  EDFFXL R2_reg_24_ ( .D(data_in_3[24]), .E(n1275), .CK(clk), .Q(R2[24]) );
  EDFFXL R2_reg_23_ ( .D(data_in_3[23]), .E(n1275), .CK(clk), .Q(R2[23]) );
  EDFFXL R2_reg_22_ ( .D(data_in_3[22]), .E(n1275), .CK(clk), .Q(R2[22]) );
  EDFFXL R2_reg_21_ ( .D(data_in_3[21]), .E(n1275), .CK(clk), .Q(R2[21]) );
  EDFFXL R2_reg_20_ ( .D(data_in_3[20]), .E(n1275), .CK(clk), .Q(R2[20]) );
  EDFFXL R2_reg_19_ ( .D(data_in_3[19]), .E(n1275), .CK(clk), .Q(R2[19]) );
  EDFFXL R2_reg_18_ ( .D(data_in_3[18]), .E(n1275), .CK(clk), .Q(R2[18]) );
  EDFFXL R2_reg_11_ ( .D(data_in_3[11]), .E(n1274), .CK(clk), .Q(R2[11]) );
  EDFFXL R2_reg_10_ ( .D(data_in_3[10]), .E(n1274), .CK(clk), .Q(R2[10]) );
  EDFFXL R2_reg_9_ ( .D(data_in_3[9]), .E(n1274), .CK(clk), .Q(R2[9]) );
  EDFFXL R2_reg_8_ ( .D(data_in_3[8]), .E(n1274), .CK(clk), .Q(R2[8]) );
  EDFFXL R2_reg_7_ ( .D(data_in_3[7]), .E(n1274), .CK(clk), .Q(R2[7]) );
  EDFFXL R2_reg_5_ ( .D(data_in_3[5]), .E(n1273), .CK(clk), .Q(R2[5]) );
  EDFFXL R2_reg_4_ ( .D(data_in_3[4]), .E(n1273), .CK(clk), .Q(R2[4]) );
  EDFFXL R2_reg_3_ ( .D(data_in_3[3]), .E(n1273), .CK(clk), .Q(R2[3]) );
  EDFFXL R2_reg_2_ ( .D(data_in_3[2]), .E(n1273), .CK(clk), .Q(R2[2]) );
  EDFFXL R2_reg_1_ ( .D(data_in_3[1]), .E(n1273), .CK(clk), .Q(R2[1]) );
  EDFFX1 R2_reg_0_ ( .D(data_in_3[0]), .E(n1273), .CK(clk), .Q(R2[0]) );
  JKFFRXL counter_1_reg_0_ ( .J(1'b1), .K(1'b1), .CK(clk), .RN(rst_n), .Q(
        counter_1[0]), .QN(n585) );
  DFFRHQX1 counter_1_reg_1_ ( .D(N26), .CK(clk), .RN(rst_n), .Q(counter_1[1])
         );
  JKFFRXL counter_2_reg_0_ ( .J(1'b1), .K(1'b1), .CK(clk), .RN(rst_n), .Q(
        counter_2[0]), .QN(n862) );
  DFFRHQX1 counter_2_reg_1_ ( .D(N50), .CK(clk), .RN(rst_n), .Q(counter_2[1])
         );
  DFFRHQX1 counter_2_reg_2_ ( .D(n1280), .CK(clk), .RN(rst_n), .Q(counter_2[2]) );
  DFFRHQX1 counter_2_reg_3_ ( .D(N52), .CK(clk), .RN(rst_n), .Q(counter_2[3])
         );
  EDFFX1 data_out_3_reg_23_ ( .D(N142), .E(n1279), .CK(clk), .Q(data_out_3[23]) );
  EDFFX1 data_out_3_reg_22_ ( .D(N141), .E(n1279), .CK(clk), .Q(data_out_3[22]) );
  EDFFX1 data_out_3_reg_21_ ( .D(N140), .E(n1279), .CK(clk), .Q(data_out_3[21]) );
  EDFFX1 data_out_3_reg_20_ ( .D(N139), .E(n1279), .CK(clk), .Q(data_out_3[20]) );
  EDFFX1 data_out_3_reg_19_ ( .D(N138), .E(n1279), .CK(clk), .Q(data_out_3[19]) );
  EDFFX1 data_out_3_reg_18_ ( .D(N137), .E(n1279), .CK(clk), .Q(data_out_3[18]) );
  EDFFX1 data_out_3_reg_17_ ( .D(N136), .E(n1279), .CK(clk), .Q(data_out_3[17]) );
  EDFFX1 data_out_3_reg_16_ ( .D(N135), .E(n1279), .CK(clk), .Q(data_out_3[16]) );
  EDFFX1 data_out_3_reg_15_ ( .D(N134), .E(n1279), .CK(clk), .Q(data_out_3[15]) );
  EDFFX1 data_out_3_reg_14_ ( .D(N133), .E(n1279), .CK(clk), .Q(data_out_3[14]) );
  EDFFX1 data_out_3_reg_13_ ( .D(N132), .E(n1279), .CK(clk), .Q(data_out_3[13]) );
  EDFFX1 data_out_3_reg_12_ ( .D(N131), .E(n1279), .CK(clk), .Q(data_out_3[12]) );
  EDFFX1 data_out_3_reg_11_ ( .D(N130), .E(n1279), .CK(clk), .Q(data_out_3[11]) );
  EDFFX1 data_out_3_reg_10_ ( .D(N129), .E(n1279), .CK(clk), .Q(data_out_3[10]) );
  EDFFXL R4_reg_11_ ( .D(data_in_3[45]), .E(n1212), .CK(clk), .QN(n744) );
  EDFFXL R6_reg_11_ ( .D(data_in_3[45]), .E(n1273), .CK(clk), .QN(n676) );
  EDFFXL R7_reg_11_ ( .D(data_in_3[45]), .E(n1264), .CK(clk), .QN(n608) );
  EDFFXL R7_reg_27_ ( .D(data_in_3[61]), .E(n1265), .CK(clk), .QN(n592) );
  EDFFXL R6_reg_27_ ( .D(data_in_3[61]), .E(n1270), .CK(clk), .QN(n660) );
  EDFFXL R4_reg_27_ ( .D(data_in_3[61]), .E(n1213), .CK(clk), .QN(n728) );
  EDFFXL R6_reg_26_ ( .D(data_in_3[60]), .E(n1274), .CK(clk), .QN(n661) );
  EDFFXL R4_reg_26_ ( .D(data_in_3[60]), .E(n1213), .CK(clk), .QN(n729) );
  EDFFXL R7_reg_26_ ( .D(data_in_3[60]), .E(n1265), .CK(clk), .QN(n593) );
  EDFFXL R7_reg_25_ ( .D(data_in_3[59]), .E(n1265), .CK(clk), .QN(n594) );
  EDFFXL R6_reg_25_ ( .D(data_in_3[59]), .E(n1271), .CK(clk), .QN(n662) );
  EDFFXL R4_reg_25_ ( .D(data_in_3[59]), .E(n1213), .CK(clk), .QN(n730) );
  EDFFXL R7_reg_7_ ( .D(data_in_3[41]), .E(n1264), .CK(clk), .QN(n612) );
  EDFFXL R6_reg_7_ ( .D(data_in_3[41]), .E(n1275), .CK(clk), .QN(n680) );
  EDFFXL R4_reg_7_ ( .D(data_in_3[41]), .E(n1215), .CK(clk), .QN(n748) );
  EDFFX1 R2_reg_6_ ( .D(data_in_3[6]), .E(n1274), .CK(clk), .Q(R2[6]) );
  EDFFX1 R1_reg_6_ ( .D(data_in_3[6]), .E(n1222), .CK(clk), .Q(R1[6]) );
  EDFFX1 R0_reg_6_ ( .D(data_in_3[6]), .E(n1214), .CK(clk), .Q(R0[6]) );
  EDFFX1 R3_reg_6_ ( .D(data_in_3[6]), .E(n1262), .CK(clk), .Q(R3[6]) );
  EDFFXL R7_reg_28_ ( .D(data_in_3[62]), .E(n1265), .CK(clk), .QN(n591) );
  EDFFXL R6_reg_28_ ( .D(data_in_3[62]), .E(n1269), .CK(clk), .QN(n659) );
  EDFFXL R4_reg_28_ ( .D(data_in_3[62]), .E(n1209), .CK(clk), .QN(n727) );
  EDFFXL R7_reg_8_ ( .D(data_in_3[42]), .E(n1264), .CK(clk), .QN(n611) );
  EDFFXL R6_reg_8_ ( .D(data_in_3[42]), .E(n1272), .CK(clk), .QN(n679) );
  EDFFXL R4_reg_8_ ( .D(data_in_3[42]), .E(n1210), .CK(clk), .QN(n747) );
  DFFXL R1_reg_16_ ( .D(n1168), .CK(clk), .Q(n208) );
  DFFXL R0_reg_16_ ( .D(n1167), .CK(clk), .Q(n206) );
  DFFXL R13_reg_15_ ( .D(n865), .CK(clk), .Q(n204) );
  DFFXL R12_reg_15_ ( .D(n864), .CK(clk), .Q(n202) );
  DFFXL R14_reg_15_ ( .D(n866), .CK(clk), .Q(n200) );
  DFFXL R12_reg_16_ ( .D(n567), .CK(clk), .Q(n198) );
  DFFXL R1_reg_33_ ( .D(n583), .CK(clk), .Q(n196) );
  DFFXL R0_reg_33_ ( .D(n581), .CK(clk), .Q(n194) );
  DFFXL R2_reg_32_ ( .D(n861), .CK(clk), .Q(n192) );
  DFFXL R1_reg_32_ ( .D(n860), .CK(clk), .Q(n190) );
  DFFXL R2_reg_16_ ( .D(n1169), .CK(clk), .Q(n188) );
  DFFXL R13_reg_16_ ( .D(n568), .CK(clk), .Q(n186) );
  EDFFXL data_out_3_reg_7_ ( .D(N126), .E(n1279), .CK(clk), .Q(data_out_3[7])
         );
  EDFFXL data_out_3_reg_6_ ( .D(N125), .E(n1279), .CK(clk), .Q(data_out_3[6])
         );
  EDFFXL data_out_3_reg_5_ ( .D(N124), .E(n1279), .CK(clk), .Q(data_out_3[5])
         );
  EDFFXL data_out_3_reg_4_ ( .D(N123), .E(n1279), .CK(clk), .Q(data_out_3[4])
         );
  EDFFXL data_out_3_reg_3_ ( .D(N122), .E(n1279), .CK(clk), .Q(data_out_3[3])
         );
  EDFFXL data_out_3_reg_2_ ( .D(N121), .E(n1279), .CK(clk), .Q(data_out_3[2])
         );
  EDFFXL data_out_3_reg_1_ ( .D(N120), .E(n1279), .CK(clk), .Q(data_out_3[1])
         );
  EDFFXL data_out_3_reg_0_ ( .D(N119), .E(n1279), .CK(clk), .Q(data_out_3[0])
         );
  EDFFXL data_out_3_reg_9_ ( .D(N128), .E(n1279), .CK(clk), .Q(data_out_3[9])
         );
  EDFFXL data_out_3_reg_8_ ( .D(N127), .E(n1279), .CK(clk), .Q(data_out_3[8])
         );
  EDFFXL data_out_3_reg_32_ ( .D(N151), .E(n1279), .CK(clk), .Q(data_out_3[32]) );
  EDFFXL data_out_3_reg_31_ ( .D(N150), .E(n1279), .CK(clk), .Q(data_out_3[31]) );
  EDFFXL data_out_3_reg_30_ ( .D(N149), .E(n1279), .CK(clk), .Q(data_out_3[30]) );
  EDFFXL data_out_3_reg_29_ ( .D(N148), .E(n1279), .CK(clk), .Q(data_out_3[29]) );
  EDFFXL data_out_3_reg_28_ ( .D(N147), .E(n1279), .CK(clk), .Q(data_out_3[28]) );
  EDFFXL data_out_3_reg_27_ ( .D(N146), .E(n1279), .CK(clk), .Q(data_out_3[27]) );
  EDFFXL data_out_3_reg_26_ ( .D(N145), .E(n1279), .CK(clk), .Q(data_out_3[26]) );
  EDFFXL data_out_3_reg_25_ ( .D(N144), .E(n1279), .CK(clk), .Q(data_out_3[25]) );
  EDFFXL data_out_3_reg_24_ ( .D(N143), .E(n1279), .CK(clk), .Q(data_out_3[24]) );
  EDFFXL R15_reg_17_ ( .D(data_in_3[119]), .E(n1263), .CK(clk), .Q(R15[17]) );
  EDFFXL R14_reg_17_ ( .D(data_in_3[119]), .E(n20), .CK(clk), .Q(R14[17]) );
  EDFFXL R13_reg_17_ ( .D(data_in_3[119]), .E(n249), .CK(clk), .Q(R13[17]) );
  EDFFXL R12_reg_17_ ( .D(data_in_3[119]), .E(n250), .CK(clk), .Q(R12[17]) );
  EDFFXL R3_reg_17_ ( .D(data_in_3[17]), .E(n1257), .CK(clk), .Q(R3[17]) );
  EDFFXL R2_reg_17_ ( .D(data_in_3[17]), .E(n20), .CK(clk), .Q(R2[17]) );
  EDFFXL R1_reg_17_ ( .D(data_in_3[17]), .E(n249), .CK(clk), .Q(R1[17]) );
  EDFFXL R0_reg_17_ ( .D(data_in_3[17]), .E(n250), .CK(clk), .Q(R0[17]) );
  EDFFXL R15_reg_0_ ( .D(data_in_3[102]), .E(n1262), .CK(clk), .Q(R15[0]) );
  EDFFXL R13_reg_0_ ( .D(data_in_3[102]), .E(n249), .CK(clk), .Q(R13[0]) );
  EDFFXL R12_reg_0_ ( .D(data_in_3[102]), .E(n250), .CK(clk), .Q(R12[0]) );
  EDFFXL R15_reg_1_ ( .D(data_in_3[103]), .E(n1257), .CK(clk), .Q(R15[1]) );
  EDFFXL R14_reg_1_ ( .D(data_in_3[103]), .E(n20), .CK(clk), .Q(R14[1]) );
  EDFFXL R13_reg_1_ ( .D(data_in_3[103]), .E(n249), .CK(clk), .Q(R13[1]) );
  EDFFXL R12_reg_1_ ( .D(data_in_3[103]), .E(n250), .CK(clk), .Q(R12[1]) );
  EDFFXL R15_reg_18_ ( .D(data_in_3[120]), .E(n1265), .CK(clk), .Q(R15[18]) );
  EDFFXL R14_reg_18_ ( .D(data_in_3[120]), .E(n20), .CK(clk), .Q(R14[18]) );
  EDFFXL R13_reg_18_ ( .D(data_in_3[120]), .E(n249), .CK(clk), .Q(R13[18]) );
  EDFFXL R12_reg_18_ ( .D(data_in_3[120]), .E(n250), .CK(clk), .Q(R12[18]) );
  EDFFXL R11_reg_0_ ( .D(data_in_3[68]), .E(n1263), .CK(clk), .QN(n721) );
  EDFFXL R9_reg_0_ ( .D(data_in_3[68]), .E(n249), .CK(clk), .QN(n857) );
  EDFFXL R8_reg_0_ ( .D(data_in_3[68]), .E(n250), .CK(clk), .QN(n789) );
  EDFFXL R7_reg_17_ ( .D(data_in_3[51]), .E(n1257), .CK(clk), .QN(n602) );
  EDFFXL R6_reg_17_ ( .D(data_in_3[51]), .E(n1273), .CK(clk), .QN(n670) );
  EDFFXL R5_reg_17_ ( .D(data_in_3[51]), .E(n249), .CK(clk), .QN(n806) );
  EDFFXL R4_reg_17_ ( .D(data_in_3[51]), .E(n250), .CK(clk), .QN(n738) );
  EDFFXL R11_reg_17_ ( .D(data_in_3[85]), .E(n1262), .CK(clk), .QN(n704) );
  EDFFXL R10_reg_17_ ( .D(data_in_3[85]), .E(n20), .CK(clk), .QN(n636) );
  EDFFXL R9_reg_17_ ( .D(data_in_3[85]), .E(n249), .CK(clk), .QN(n840) );
  EDFFXL R8_reg_17_ ( .D(data_in_3[85]), .E(n250), .CK(clk), .QN(n772) );
  EDFFXL R7_reg_0_ ( .D(data_in_3[34]), .E(n1257), .CK(clk), .QN(n619) );
  EDFFXL R5_reg_0_ ( .D(data_in_3[34]), .E(n249), .CK(clk), .QN(n823) );
  EDFFXL R4_reg_0_ ( .D(data_in_3[34]), .E(n250), .CK(clk), .QN(n755) );
  EDFFXL R7_reg_1_ ( .D(data_in_3[35]), .E(n1257), .CK(clk), .QN(n618) );
  EDFFXL R6_reg_1_ ( .D(data_in_3[35]), .E(n20), .CK(clk), .QN(n686) );
  EDFFXL R4_reg_1_ ( .D(data_in_3[35]), .E(n250), .CK(clk), .QN(n754) );
  DFFHQXL R15_reg_12_ ( .D(n1180), .CK(clk), .Q(R15[12]) );
  DFFHQXL R12_reg_12_ ( .D(n1177), .CK(clk), .Q(R12[12]) );
  DFFHQXL R14_reg_12_ ( .D(n1179), .CK(clk), .Q(R14[12]) );
  DFFHQXL R13_reg_12_ ( .D(n1178), .CK(clk), .Q(R13[12]) );
  DFFHQXL R1_reg_12_ ( .D(n1190), .CK(clk), .Q(R1[12]) );
  DFFHQXL R0_reg_12_ ( .D(n1189), .CK(clk), .Q(R0[12]) );
  DFFHQXL R3_reg_12_ ( .D(n1192), .CK(clk), .Q(R3[12]) );
  DFFHQXL R2_reg_12_ ( .D(n1191), .CK(clk), .Q(R2[12]) );
  DFFHQXL R15_reg_30_ ( .D(n1188), .CK(clk), .Q(R15[30]) );
  DFFHQXL R14_reg_30_ ( .D(n1187), .CK(clk), .Q(R14[30]) );
  DFFHQXL R13_reg_30_ ( .D(n1186), .CK(clk), .Q(R13[30]) );
  DFFHQXL R12_reg_30_ ( .D(n1185), .CK(clk), .Q(R12[30]) );
  DFFHQXL R1_reg_13_ ( .D(n1182), .CK(clk), .Q(R1[13]) );
  DFFHQXL R0_reg_13_ ( .D(n1181), .CK(clk), .Q(R0[13]) );
  DFFHQXL R3_reg_13_ ( .D(n1184), .CK(clk), .Q(R3[13]) );
  DFFHQXL R2_reg_13_ ( .D(n1183), .CK(clk), .Q(R2[13]) );
  DFFHQXL R2_reg_30_ ( .D(n1173), .CK(clk), .Q(R2[30]) );
  DFFHQXL R1_reg_30_ ( .D(n1172), .CK(clk), .Q(R1[30]) );
  DFFHQXL R0_reg_30_ ( .D(n1171), .CK(clk), .Q(R0[30]) );
  DFFHQXL R3_reg_30_ ( .D(n1174), .CK(clk), .Q(R3[30]) );
  DFFHQXL R2_reg_31_ ( .D(n896), .CK(clk), .Q(R2[31]) );
  DFFHQXL R1_reg_31_ ( .D(n894), .CK(clk), .Q(R1[31]) );
  DFFHQXL R0_reg_31_ ( .D(n892), .CK(clk), .Q(R0[31]) );
  DFFHQXL R3_reg_31_ ( .D(n1166), .CK(clk), .Q(R3[31]) );
  DFFHQXL R15_reg_14_ ( .D(n891), .CK(clk), .Q(R15[14]) );
  DFFHQXL R12_reg_14_ ( .D(n881), .CK(clk), .Q(R12[14]) );
  DFFHQXL R14_reg_14_ ( .D(n886), .CK(clk), .Q(R14[14]) );
  DFFHQXL R13_reg_14_ ( .D(n882), .CK(clk), .Q(R13[14]) );
  DFFHQXL R15_reg_31_ ( .D(n578), .CK(clk), .Q(R15[31]) );
  DFFHQXL R14_reg_31_ ( .D(n577), .CK(clk), .Q(R14[31]) );
  DFFHQXL R13_reg_31_ ( .D(n576), .CK(clk), .Q(R13[31]) );
  DFFHQXL R12_reg_31_ ( .D(n575), .CK(clk), .Q(R12[31]) );
  DFFHQXL R1_reg_14_ ( .D(n572), .CK(clk), .Q(R1[14]) );
  DFFHQXL R0_reg_14_ ( .D(n571), .CK(clk), .Q(R0[14]) );
  DFFHQXL R3_reg_14_ ( .D(n574), .CK(clk), .Q(R3[14]) );
  DFFHQXL R2_reg_14_ ( .D(n573), .CK(clk), .Q(R2[14]) );
  DFFHQXL R15_reg_32_ ( .D(n580), .CK(clk), .Q(R15[32]) );
  DFFHQXL R14_reg_32_ ( .D(n579), .CK(clk), .Q(R14[32]) );
  DFFHQXL R13_reg_32_ ( .D(n1176), .CK(clk), .Q(R13[32]) );
  DFFHQXL R12_reg_32_ ( .D(n1175), .CK(clk), .Q(R12[32]) );
  DFFHQXL R3_reg_32_ ( .D(n863), .CK(clk), .Q(R3[32]) );
  DFFHQXL R15_reg_15_ ( .D(n867), .CK(clk), .Q(R15[15]) );
  DFFHQXL R0_reg_32_ ( .D(n859), .CK(clk), .Q(R0[32]) );
  DFFHQXL R2_reg_33_ ( .D(n584), .CK(clk), .Q(R2[33]) );
  DFFHQXL R1_reg_15_ ( .D(n564), .CK(clk), .Q(R1[15]) );
  DFFHQXL R0_reg_15_ ( .D(n563), .CK(clk), .Q(R0[15]) );
  DFFHQXL R3_reg_15_ ( .D(n566), .CK(clk), .Q(R3[15]) );
  DFFHQXL R3_reg_33_ ( .D(n858), .CK(clk), .Q(R3[33]) );
  DFFHQXL R2_reg_15_ ( .D(n565), .CK(clk), .Q(R2[15]) );
  DFFHQXL R14_reg_33_ ( .D(n561), .CK(clk), .Q(R14[33]) );
  DFFHQXL R13_reg_33_ ( .D(n560), .CK(clk), .Q(R13[33]) );
  DFFHQXL R12_reg_33_ ( .D(n559), .CK(clk), .Q(R12[33]) );
  EDFFXL R11_reg_29_ ( .D(data_in_3[97]), .E(n1264), .CK(clk), .QN(n692) );
  EDFFXL R10_reg_29_ ( .D(data_in_3[97]), .E(n1276), .CK(clk), .QN(n624) );
  EDFFXL R9_reg_29_ ( .D(data_in_3[97]), .E(n249), .CK(clk), .QN(n828) );
  EDFFXL R11_reg_13_ ( .D(data_in_3[81]), .E(n1265), .CK(clk), .QN(n708) );
  EDFFXL R10_reg_13_ ( .D(data_in_3[81]), .E(n20), .CK(clk), .QN(n640) );
  EDFFXL R9_reg_13_ ( .D(data_in_3[81]), .E(n249), .CK(clk), .QN(n844) );
  EDFFXL R8_reg_13_ ( .D(data_in_3[81]), .E(n250), .CK(clk), .QN(n776) );
  EDFFXL R11_reg_12_ ( .D(data_in_3[80]), .E(n1263), .CK(clk), .QN(n709) );
  EDFFXL R10_reg_12_ ( .D(data_in_3[80]), .E(n20), .CK(clk), .QN(n641) );
  EDFFXL R9_reg_12_ ( .D(data_in_3[80]), .E(n249), .CK(clk), .QN(n845) );
  EDFFXL R6_reg_13_ ( .D(data_in_3[47]), .E(n1269), .CK(clk), .QN(n674) );
  EDFFXL R4_reg_13_ ( .D(data_in_3[47]), .E(n250), .CK(clk), .QN(n742) );
  EDFFXL R7_reg_13_ ( .D(data_in_3[47]), .E(n1257), .CK(clk), .QN(n606) );
  EDFFXL R5_reg_13_ ( .D(data_in_3[47]), .E(n249), .CK(clk), .QN(n810) );
  EDFFXL R11_reg_30_ ( .D(data_in_3[98]), .E(n1262), .CK(clk), .QN(n691) );
  EDFFXL R10_reg_30_ ( .D(data_in_3[98]), .E(n20), .CK(clk), .QN(n623) );
  EDFFXL R9_reg_30_ ( .D(data_in_3[98]), .E(n249), .CK(clk), .QN(n827) );
  EDFFXL R11_reg_31_ ( .D(data_in_3[99]), .E(n1258), .CK(clk), .QN(n690) );
  EDFFXL R8_reg_31_ ( .D(data_in_3[99]), .E(n250), .CK(clk), .QN(n758) );
  EDFFXL R10_reg_31_ ( .D(data_in_3[99]), .E(n20), .CK(clk), .QN(n622) );
  EDFFXL R9_reg_31_ ( .D(data_in_3[99]), .E(n249), .CK(clk), .QN(n826) );
  EDFFXL R7_reg_31_ ( .D(data_in_3[65]), .E(n1257), .CK(clk), .QN(n588) );
  EDFFXL R6_reg_31_ ( .D(data_in_3[65]), .E(n20), .CK(clk), .QN(n656) );
  EDFFXL R4_reg_31_ ( .D(data_in_3[65]), .E(n250), .CK(clk), .QN(n724) );
  EDFFXL R5_reg_31_ ( .D(data_in_3[65]), .E(n249), .CK(clk), .QN(n792) );
  EDFFXL R6_reg_14_ ( .D(data_in_3[48]), .E(n1276), .CK(clk), .QN(n673) );
  EDFFXL R4_reg_14_ ( .D(data_in_3[48]), .E(n250), .CK(clk), .QN(n741) );
  EDFFXL R7_reg_14_ ( .D(data_in_3[48]), .E(n1257), .CK(clk), .QN(n605) );
  EDFFXL R5_reg_14_ ( .D(data_in_3[48]), .E(n249), .CK(clk), .QN(n809) );
  EDFFXL R10_reg_15_ ( .D(data_in_3[83]), .E(n20), .CK(clk), .QN(n638) );
  EDFFXL R6_reg_12_ ( .D(data_in_3[46]), .E(n20), .CK(clk), .QN(n675) );
  EDFFXL R7_reg_12_ ( .D(data_in_3[46]), .E(n1257), .CK(clk), .QN(n607) );
  EDFFXL R5_reg_12_ ( .D(data_in_3[46]), .E(n249), .CK(clk), .QN(n811) );
  EDFFXL R8_reg_30_ ( .D(data_in_3[98]), .E(n250), .CK(clk), .QN(n759) );
  EDFFXL R11_reg_32_ ( .D(data_in_3[100]), .E(n1265), .CK(clk), .QN(n689) );
  EDFFXL R8_reg_32_ ( .D(data_in_3[100]), .E(n250), .CK(clk), .QN(n757) );
  EDFFXL R10_reg_32_ ( .D(data_in_3[100]), .E(n20), .CK(clk), .QN(n621) );
  EDFFXL R9_reg_32_ ( .D(data_in_3[100]), .E(n249), .CK(clk), .QN(n825) );
  EDFFXL R10_reg_16_ ( .D(data_in_3[84]), .E(n1274), .CK(clk), .QN(n637) );
  EDFFXL R8_reg_33_ ( .D(data_in_3[101]), .E(n250), .CK(clk), .QN(n756) );
  EDFFXL R11_reg_33_ ( .D(data_in_3[101]), .E(n1263), .CK(clk), .QN(n688) );
  EDFFXL R11_reg_15_ ( .D(data_in_3[83]), .E(n1258), .CK(clk), .QN(n706) );
  EDFFXL R9_reg_15_ ( .D(data_in_3[83]), .E(n249), .CK(clk), .QN(n842) );
  EDFFXL R8_reg_15_ ( .D(data_in_3[83]), .E(n250), .CK(clk), .QN(n774) );
  EDFFXL R7_reg_32_ ( .D(data_in_3[66]), .E(n1257), .CK(clk), .QN(n587) );
  EDFFXL R7_reg_33_ ( .D(data_in_3[67]), .E(n1257), .CK(clk), .QN(n586) );
  EDFFXL R6_reg_15_ ( .D(data_in_3[49]), .E(n1270), .CK(clk), .QN(n672) );
  EDFFXL R4_reg_15_ ( .D(data_in_3[49]), .E(n250), .CK(clk), .QN(n740) );
  EDFFXL R7_reg_15_ ( .D(data_in_3[49]), .E(n1257), .CK(clk), .QN(n604) );
  EDFFXL R5_reg_15_ ( .D(data_in_3[49]), .E(n249), .CK(clk), .QN(n808) );
  EDFFXL R6_reg_32_ ( .D(data_in_3[66]), .E(n1275), .CK(clk), .QN(n655) );
  EDFFXL R4_reg_32_ ( .D(data_in_3[66]), .E(n250), .CK(clk), .QN(n723) );
  EDFFXL R5_reg_32_ ( .D(data_in_3[66]), .E(n249), .CK(clk), .QN(n791) );
  EDFFXL R11_reg_16_ ( .D(data_in_3[84]), .E(n1263), .CK(clk), .QN(n705) );
  EDFFXL R9_reg_16_ ( .D(data_in_3[84]), .E(n249), .CK(clk), .QN(n841) );
  EDFFXL R8_reg_16_ ( .D(data_in_3[84]), .E(n250), .CK(clk), .QN(n773) );
  EDFFXL R6_reg_33_ ( .D(data_in_3[67]), .E(n20), .CK(clk), .QN(n654) );
  EDFFXL R4_reg_33_ ( .D(data_in_3[67]), .E(n250), .CK(clk), .QN(n722) );
  EDFFXL R5_reg_33_ ( .D(data_in_3[67]), .E(n249), .CK(clk), .QN(n790) );
  EDFFXL R4_reg_16_ ( .D(data_in_3[50]), .E(n250), .CK(clk), .QN(n739) );
  EDFFXL R10_reg_33_ ( .D(data_in_3[101]), .E(n1272), .CK(clk), .QN(n620) );
  EDFFXL R9_reg_33_ ( .D(data_in_3[101]), .E(n249), .CK(clk), .QN(n824) );
  EDFFXL R6_reg_16_ ( .D(data_in_3[50]), .E(n1271), .CK(clk), .QN(n671) );
  EDFFXL R5_reg_16_ ( .D(data_in_3[50]), .E(n249), .CK(clk), .QN(n807) );
  EDFFXL R7_reg_16_ ( .D(data_in_3[50]), .E(n1257), .CK(clk), .QN(n603) );
  JKFFRX2 p_s_flag_out_reg ( .J(n1283), .K(1'b0), .CK(clk), .RN(rst_n), .Q(
        n1279) );
  EDFFX1 data_out_3_reg_33_ ( .D(N152), .E(n1279), .CK(clk), .Q(data_out_3[33]) );
  EDFFX1 R14_reg_0_ ( .D(data_in_3[102]), .E(n1276), .CK(clk), .Q(R14[0]) );
  EDFFX1 R6_reg_0_ ( .D(data_in_3[34]), .E(n1273), .CK(clk), .QN(n687) );
  EDFFX1 R10_reg_0_ ( .D(data_in_3[68]), .E(n1276), .CK(clk), .QN(n653) );
  EDFFX2 R4_reg_12_ ( .D(data_in_3[46]), .E(n250), .CK(clk), .QN(n743) );
  EDFFXL R7_reg_29_ ( .D(data_in_3[63]), .E(n1265), .CK(clk), .QN(n590) );
  EDFFXL R6_reg_29_ ( .D(data_in_3[63]), .E(n1270), .CK(clk), .QN(n658) );
  EDFFXL R4_reg_29_ ( .D(data_in_3[63]), .E(n1215), .CK(clk), .QN(n726) );
  EDFFXL R7_reg_24_ ( .D(data_in_3[58]), .E(n1265), .CK(clk), .QN(n595) );
  EDFFXL R6_reg_24_ ( .D(data_in_3[58]), .E(n1272), .CK(clk), .QN(n663) );
  EDFFXL R4_reg_24_ ( .D(data_in_3[58]), .E(n1213), .CK(clk), .QN(n731) );
  EDFFX2 R4_reg_30_ ( .D(data_in_3[64]), .E(n250), .CK(clk), .QN(n725) );
  EDFFX2 R8_reg_14_ ( .D(data_in_3[82]), .E(n250), .CK(clk), .QN(n775) );
  EDFFX2 R9_reg_14_ ( .D(data_in_3[82]), .E(n249), .CK(clk), .QN(n843) );
  EDFFX2 R10_reg_14_ ( .D(data_in_3[82]), .E(n1274), .CK(clk), .QN(n639) );
  EDFFX2 R11_reg_14_ ( .D(data_in_3[82]), .E(n1263), .CK(clk), .QN(n707) );
  EDFFX2 R5_reg_30_ ( .D(data_in_3[64]), .E(n249), .CK(clk), .QN(n793) );
  EDFFX2 R8_reg_29_ ( .D(data_in_3[97]), .E(n250), .CK(clk), .QN(n760) );
  EDFFX2 R8_reg_12_ ( .D(data_in_3[80]), .E(n250), .CK(clk), .QN(n777) );
  EDFFXL R10_reg_9_ ( .D(data_in_3[77]), .E(n1269), .CK(clk), .QN(n644) );
  EDFFXL R11_reg_9_ ( .D(data_in_3[77]), .E(n1264), .CK(clk), .QN(n712) );
  EDFFXL R8_reg_9_ ( .D(data_in_3[77]), .E(n1209), .CK(clk), .QN(n780) );
  EDFFXL R9_reg_9_ ( .D(data_in_3[77]), .E(n1217), .CK(clk), .QN(n848) );
  EDFFXL R3_reg_26_ ( .D(data_in_3[26]), .E(n1263), .CK(clk), .Q(R3[26]) );
  EDFFXL R0_reg_26_ ( .D(data_in_3[26]), .E(n1213), .CK(clk), .Q(R0[26]) );
  EDFFXL R1_reg_26_ ( .D(data_in_3[26]), .E(n1217), .CK(clk), .Q(R1[26]) );
  EDFFXL R2_reg_26_ ( .D(data_in_3[26]), .E(n1275), .CK(clk), .Q(R2[26]) );
  EDFFXL R7_reg_23_ ( .D(data_in_3[57]), .E(n1265), .CK(clk), .QN(n596) );
  EDFFXL R6_reg_23_ ( .D(data_in_3[57]), .E(n1276), .CK(clk), .QN(n664) );
  EDFFXL R4_reg_23_ ( .D(data_in_3[57]), .E(n1213), .CK(clk), .QN(n732) );
  EDFFXL R3_reg_25_ ( .D(data_in_3[25]), .E(n1263), .CK(clk), .Q(R3[25]) );
  EDFFXL R0_reg_25_ ( .D(data_in_3[25]), .E(n1209), .CK(clk), .Q(R0[25]) );
  EDFFXL R1_reg_25_ ( .D(data_in_3[25]), .E(n1221), .CK(clk), .Q(R1[25]) );
  EDFFXL R2_reg_25_ ( .D(data_in_3[25]), .E(n1275), .CK(clk), .Q(R2[25]) );
  EDFFXL R7_reg_30_ ( .D(data_in_3[64]), .E(n1257), .CK(clk), .QN(n589) );
  EDFFXL R6_reg_30_ ( .D(data_in_3[64]), .E(n1269), .CK(clk), .QN(n657) );
  DFFXL R14_reg_16_ ( .D(n569), .CK(clk), .Q(n7) );
  DFFXL R15_reg_33_ ( .D(n562), .CK(clk), .Q(n6) );
  DFFXL R15_reg_16_ ( .D(n570), .CK(clk), .Q(n4) );
  DFFXL R3_reg_16_ ( .D(n1170), .CK(clk), .Q(n1) );
  MX2X1 U3 ( .A(n6), .B(data_in_3[135]), .S0(n1260), .Y(n562) );
  MX2X1 U6 ( .A(data_in_3[118]), .B(n186), .S0(n3), .Y(n568) );
  CLKINVX20 U7 ( .A(n1218), .Y(n3) );
  MX2X1 U8 ( .A(data_in_3[118]), .B(n198), .S0(n13), .Y(n567) );
  INVX20 U9 ( .A(n1210), .Y(n13) );
  NAND2X4 U10 ( .A(data_in_3[33]), .B(n17), .Y(n18) );
  NAND2X4 U11 ( .A(data_in_3[33]), .B(n10), .Y(n11) );
  MX2X2 U12 ( .A(n194), .B(data_in_3[33]), .S0(n1215), .Y(n581) );
  MX2X2 U13 ( .A(n196), .B(data_in_3[33]), .S0(n1223), .Y(n583) );
  MX2X4 U14 ( .A(data_in_3[118]), .B(n7), .S0(n1277), .Y(n569) );
  MX2X4 U15 ( .A(data_in_3[118]), .B(n4), .S0(n1268), .Y(n570) );
  NAND2X4 U16 ( .A(n60), .B(n59), .Y(n1170) );
  NAND2X4 U17 ( .A(R3[33]), .B(n1267), .Y(n12) );
  NAND2X2 U18 ( .A(n11), .B(n12), .Y(n858) );
  INVX12 U19 ( .A(n1267), .Y(n10) );
  INVX2 U20 ( .A(n1257), .Y(n1267) );
  MX2X4 U21 ( .A(data_in_3[12]), .B(R1[12]), .S0(n1224), .Y(n1190) );
  MX2X2 U22 ( .A(R15[12]), .B(data_in_3[114]), .S0(n1259), .Y(n1180) );
  MX2X2 U23 ( .A(R3[29]), .B(data_in_3[29]), .S0(n1262), .Y(n1200) );
  MX2X2 U24 ( .A(R0[29]), .B(data_in_3[29]), .S0(n1214), .Y(n1194) );
  MX2X2 U25 ( .A(R2[29]), .B(data_in_3[29]), .S0(n1275), .Y(n1198) );
  MX2X2 U26 ( .A(R1[29]), .B(data_in_3[29]), .S0(n1218), .Y(n1196) );
  MX2X4 U27 ( .A(data_in_3[13]), .B(R3[13]), .S0(n1266), .Y(n1184) );
  MX2X4 U28 ( .A(data_in_3[115]), .B(R12[13]), .S0(n13), .Y(n1202) );
  MX2X2 U29 ( .A(R13[12]), .B(data_in_3[114]), .S0(n1218), .Y(n1178) );
  MX2X4 U30 ( .A(data_in_3[114]), .B(R12[12]), .S0(n14), .Y(n1177) );
  CLKINVX20 U31 ( .A(n1210), .Y(n14) );
  NAND2X4 U32 ( .A(R2[33]), .B(n1277), .Y(n19) );
  NAND2X2 U33 ( .A(n18), .B(n19), .Y(n584) );
  INVX12 U34 ( .A(n1277), .Y(n17) );
  INVX1 U35 ( .A(n20), .Y(n1277) );
  NAND2X2 U36 ( .A(n1), .B(n1267), .Y(n60) );
  MX2X2 U37 ( .A(R14[12]), .B(data_in_3[114]), .S0(n1271), .Y(n1179) );
  NOR3X2 U38 ( .A(counter_1[1]), .B(p_s_flag_in), .C(counter_1[0]), .Y(n20) );
  AND2X2 U39 ( .A(n1163), .B(n873), .Y(n21) );
  NAND2X1 U40 ( .A(n1159), .B(n872), .Y(n22) );
  NAND2X1 U41 ( .A(n1159), .B(n870), .Y(n23) );
  NAND2X1 U42 ( .A(n872), .B(n1164), .Y(n24) );
  NAND2X1 U43 ( .A(n1158), .B(n872), .Y(n25) );
  NAND2X1 U44 ( .A(n1163), .B(n872), .Y(n26) );
  NAND2X1 U45 ( .A(n1163), .B(n870), .Y(n27) );
  INVXL U46 ( .A(n250), .Y(n1216) );
  MX2X2 U47 ( .A(R14[13]), .B(data_in_3[115]), .S0(n1271), .Y(n1206) );
  MX2X2 U48 ( .A(R13[13]), .B(data_in_3[115]), .S0(n1218), .Y(n1204) );
  MX2X2 U49 ( .A(R15[13]), .B(data_in_3[115]), .S0(n1259), .Y(n1208) );
  MX2X2 U50 ( .A(R0[12]), .B(data_in_3[12]), .S0(n1214), .Y(n1189) );
  MX2X2 U51 ( .A(R2[12]), .B(data_in_3[12]), .S0(n1274), .Y(n1191) );
  MX2X2 U52 ( .A(R3[12]), .B(data_in_3[12]), .S0(n1262), .Y(n1192) );
  MX2X2 U53 ( .A(R12[30]), .B(data_in_3[132]), .S0(n1211), .Y(n1185) );
  MX2X2 U54 ( .A(R13[30]), .B(data_in_3[132]), .S0(n1219), .Y(n1186) );
  MX2X2 U55 ( .A(R14[30]), .B(data_in_3[132]), .S0(n1273), .Y(n1187) );
  MX2X2 U56 ( .A(R15[30]), .B(data_in_3[132]), .S0(n1260), .Y(n1188) );
  MX2X2 U57 ( .A(data_in_3[133]), .B(R15[31]), .S0(n1267), .Y(n578) );
  MX2X2 U58 ( .A(R13[31]), .B(data_in_3[133]), .S0(n1219), .Y(n576) );
  MX2X2 U59 ( .A(R0[13]), .B(data_in_3[13]), .S0(n1214), .Y(n1181) );
  MX2X2 U60 ( .A(R1[13]), .B(data_in_3[13]), .S0(n1222), .Y(n1182) );
  MX2X2 U61 ( .A(R2[13]), .B(data_in_3[13]), .S0(n1274), .Y(n1183) );
  MX2X2 U62 ( .A(R14[31]), .B(data_in_3[133]), .S0(n1273), .Y(n577) );
  MX2X2 U63 ( .A(R12[31]), .B(data_in_3[133]), .S0(n1211), .Y(n575) );
  MX2X4 U64 ( .A(data_in_3[134]), .B(R14[32]), .S0(n1278), .Y(n579) );
  MX2X2 U65 ( .A(n188), .B(data_in_3[16]), .S0(n1274), .Y(n1169) );
  MX2X2 U66 ( .A(n206), .B(data_in_3[16]), .S0(n1214), .Y(n1167) );
  MX2X2 U67 ( .A(n208), .B(data_in_3[16]), .S0(n1222), .Y(n1168) );
  NAND2X4 U68 ( .A(data_in_3[16]), .B(n1261), .Y(n59) );
  MX2X1 U69 ( .A(n190), .B(data_in_3[32]), .S0(n1223), .Y(n860) );
  MX2X1 U71 ( .A(n192), .B(data_in_3[32]), .S0(n1276), .Y(n861) );
  MX2X4 U72 ( .A(data_in_3[117]), .B(R15[15]), .S0(n1268), .Y(n867) );
  MX2X2 U73 ( .A(R3[30]), .B(data_in_3[30]), .S0(n1260), .Y(n1174) );
  MX2X2 U74 ( .A(R0[30]), .B(data_in_3[30]), .S0(n1215), .Y(n1171) );
  MX2X2 U75 ( .A(R1[30]), .B(data_in_3[30]), .S0(n1223), .Y(n1172) );
  MX2X2 U76 ( .A(R2[30]), .B(data_in_3[30]), .S0(n1276), .Y(n1173) );
  MX2X2 U77 ( .A(R0[14]), .B(data_in_3[14]), .S0(n1214), .Y(n571) );
  MX2X2 U78 ( .A(R1[14]), .B(data_in_3[14]), .S0(n1222), .Y(n572) );
  MX2X2 U79 ( .A(R2[14]), .B(data_in_3[14]), .S0(n1274), .Y(n573) );
  MX2X2 U80 ( .A(R3[14]), .B(data_in_3[14]), .S0(n1262), .Y(n574) );
  MX2X2 U81 ( .A(R3[31]), .B(data_in_3[31]), .S0(n1265), .Y(n1166) );
  MX2X2 U82 ( .A(R0[31]), .B(data_in_3[31]), .S0(n1215), .Y(n892) );
  MX2X2 U83 ( .A(R1[31]), .B(data_in_3[31]), .S0(n1223), .Y(n894) );
  MX2X2 U84 ( .A(R2[31]), .B(data_in_3[31]), .S0(n1276), .Y(n896) );
  MX2X2 U85 ( .A(data_in_3[32]), .B(R3[32]), .S0(n251), .Y(n863) );
  MX2X2 U86 ( .A(n202), .B(data_in_3[117]), .S0(n1210), .Y(n864) );
  MX2X2 U87 ( .A(n204), .B(data_in_3[117]), .S0(n1218), .Y(n865) );
  MX2X2 U88 ( .A(n200), .B(data_in_3[117]), .S0(n1271), .Y(n866) );
  MX2X2 U89 ( .A(R0[15]), .B(data_in_3[15]), .S0(n1214), .Y(n563) );
  MX2X2 U90 ( .A(R1[15]), .B(data_in_3[15]), .S0(n1222), .Y(n564) );
  MX2X2 U91 ( .A(R2[15]), .B(data_in_3[15]), .S0(n1274), .Y(n565) );
  MX2X2 U92 ( .A(R3[15]), .B(data_in_3[15]), .S0(n1262), .Y(n566) );
  MX2X2 U93 ( .A(R15[32]), .B(data_in_3[134]), .S0(n1260), .Y(n580) );
  MX2X2 U94 ( .A(R12[32]), .B(data_in_3[134]), .S0(n1211), .Y(n1175) );
  MX2X2 U95 ( .A(R13[32]), .B(data_in_3[134]), .S0(n1219), .Y(n1176) );
  MX2X2 U96 ( .A(R12[33]), .B(data_in_3[135]), .S0(n1211), .Y(n559) );
  MX2X2 U97 ( .A(R13[33]), .B(data_in_3[135]), .S0(n1219), .Y(n560) );
  MX2X2 U98 ( .A(R14[33]), .B(data_in_3[135]), .S0(n1273), .Y(n561) );
  MX2X2 U99 ( .A(R12[14]), .B(data_in_3[116]), .S0(n1210), .Y(n881) );
  MX2X2 U100 ( .A(R13[14]), .B(data_in_3[116]), .S0(n1218), .Y(n882) );
  MX2X2 U101 ( .A(R15[14]), .B(data_in_3[116]), .S0(n1259), .Y(n891) );
  MX2X2 U102 ( .A(R14[14]), .B(data_in_3[116]), .S0(n1271), .Y(n886) );
  MX2X2 U103 ( .A(R0[32]), .B(data_in_3[32]), .S0(n1215), .Y(n859) );
  INVX1 U104 ( .A(n868), .Y(n1225) );
  INVX1 U105 ( .A(n868), .Y(n1226) );
  INVX1 U106 ( .A(n23), .Y(n1244) );
  INVX1 U107 ( .A(n25), .Y(n1250) );
  INVX1 U108 ( .A(n1242), .Y(n1241) );
  INVX1 U109 ( .A(n26), .Y(n1234) );
  INVX1 U110 ( .A(n27), .Y(n1228) );
  INVX1 U111 ( .A(n22), .Y(n1252) );
  INVX1 U112 ( .A(n24), .Y(n1236) );
  INVX1 U113 ( .A(n1256), .Y(n1255) );
  INVX1 U114 ( .A(n1248), .Y(n1247) );
  INVX1 U115 ( .A(n1240), .Y(n1239) );
  INVX1 U116 ( .A(n1232), .Y(n1231) );
  INVX1 U117 ( .A(n21), .Y(n1230) );
  INVX1 U118 ( .A(n1254), .Y(n1253) );
  INVX1 U119 ( .A(n1246), .Y(n1245) );
  INVX1 U120 ( .A(n1238), .Y(n1237) );
  INVX1 U121 ( .A(n1277), .Y(n1272) );
  INVX1 U122 ( .A(n1266), .Y(n1263) );
  INVX1 U123 ( .A(n1267), .Y(n1260) );
  INVX1 U124 ( .A(n1278), .Y(n1271) );
  INVX1 U125 ( .A(n1266), .Y(n1262) );
  INVX1 U126 ( .A(n1278), .Y(n1273) );
  INVX1 U127 ( .A(n1268), .Y(n1259) );
  INVX1 U128 ( .A(n1278), .Y(n1274) );
  INVX1 U129 ( .A(n1268), .Y(n1258) );
  INVX1 U130 ( .A(n1266), .Y(n1265) );
  INVX1 U131 ( .A(n1277), .Y(n1275) );
  INVX1 U132 ( .A(n1277), .Y(n1269) );
  INVX1 U133 ( .A(n1278), .Y(n1270) );
  INVX1 U134 ( .A(n1268), .Y(n1261) );
  INVX1 U135 ( .A(n251), .Y(n1264) );
  INVX1 U136 ( .A(n1277), .Y(n1276) );
  INVX1 U137 ( .A(n22), .Y(n1251) );
  INVX1 U138 ( .A(n23), .Y(n1243) );
  INVX1 U139 ( .A(n24), .Y(n1235) );
  INVX1 U140 ( .A(n25), .Y(n1249) );
  INVX1 U141 ( .A(n27), .Y(n1227) );
  INVX1 U142 ( .A(n888), .Y(n1240) );
  INVX1 U143 ( .A(n893), .Y(n1232) );
  INVX1 U144 ( .A(n21), .Y(n1229) );
  INVX1 U145 ( .A(n1224), .Y(n1221) );
  INVX1 U146 ( .A(n1216), .Y(n1213) );
  INVX1 U147 ( .A(n1216), .Y(n1212) );
  INVX1 U148 ( .A(n1224), .Y(n1219) );
  INVX1 U149 ( .A(n1224), .Y(n1220) );
  INVX1 U150 ( .A(n1216), .Y(n1211) );
  INVX1 U151 ( .A(n1224), .Y(n1218) );
  INVX1 U152 ( .A(n1224), .Y(n1222) );
  INVX1 U153 ( .A(n1216), .Y(n1210) );
  INVX1 U154 ( .A(n1216), .Y(n1214) );
  INVX1 U155 ( .A(n1216), .Y(n1215) );
  INVX1 U156 ( .A(n1224), .Y(n1223) );
  INVX1 U157 ( .A(n1264), .Y(n1268) );
  INVX1 U158 ( .A(n1257), .Y(n1266) );
  INVX1 U159 ( .A(n20), .Y(n1278) );
  INVX1 U160 ( .A(n883), .Y(n1248) );
  INVX1 U161 ( .A(n884), .Y(n1246) );
  INVX1 U162 ( .A(n878), .Y(n1256) );
  INVX1 U163 ( .A(n879), .Y(n1254) );
  INVX1 U164 ( .A(n887), .Y(n1242) );
  INVX1 U165 ( .A(n889), .Y(n1238) );
  INVX1 U166 ( .A(n26), .Y(n1233) );
  INVX1 U167 ( .A(n1224), .Y(n1217) );
  INVX1 U168 ( .A(n1216), .Y(n1209) );
  NOR2X1 U169 ( .A(n1282), .B(n1281), .Y(n870) );
  NAND2X1 U170 ( .A(n1164), .B(n870), .Y(n868) );
  NAND2X1 U171 ( .A(n1160), .B(n1159), .Y(n878) );
  NAND2X1 U172 ( .A(n873), .B(n1159), .Y(n883) );
  NAND2X1 U173 ( .A(n1160), .B(n1158), .Y(n879) );
  NAND2X1 U174 ( .A(n873), .B(n1158), .Y(n884) );
  NAND2X1 U175 ( .A(n873), .B(n1164), .Y(n893) );
  NAND2X1 U176 ( .A(n1160), .B(n1164), .Y(n888) );
  NAND2X1 U177 ( .A(n1163), .B(n1160), .Y(n889) );
  INVX1 U178 ( .A(n251), .Y(n1257) );
  INVX1 U179 ( .A(n249), .Y(n1224) );
  NOR2X1 U180 ( .A(n1282), .B(counter_2[1]), .Y(n873) );
  NOR2X1 U181 ( .A(counter_2[2]), .B(counter_2[1]), .Y(n1160) );
  NOR2X1 U182 ( .A(n862), .B(counter_2[3]), .Y(n1164) );
  OAI221XL U183 ( .A0(n857), .A1(n878), .B0(n823), .B1(n1253), .C0(n1157), .Y(
        n1156) );
  AOI22X1 U184 ( .A0(n1251), .A1(R2[0]), .B0(n1249), .B1(R13[0]), .Y(n1157) );
  OAI221XL U185 ( .A0(n856), .A1(n1255), .B0(n822), .B1(n1253), .C0(n1149), 
        .Y(n1148) );
  AOI22X1 U186 ( .A0(n1251), .A1(R2[1]), .B0(n1249), .B1(R13[1]), .Y(n1149) );
  OAI221XL U187 ( .A0(n855), .A1(n878), .B0(n821), .B1(n1253), .C0(n1141), .Y(
        n1140) );
  AOI22X1 U188 ( .A0(n1251), .A1(R2[2]), .B0(n1249), .B1(R13[2]), .Y(n1141) );
  OAI221XL U189 ( .A0(n854), .A1(n878), .B0(n820), .B1(n1253), .C0(n1133), .Y(
        n1132) );
  AOI22X1 U190 ( .A0(n1251), .A1(R2[3]), .B0(n1249), .B1(R13[3]), .Y(n1133) );
  OAI221XL U191 ( .A0(n853), .A1(n878), .B0(n819), .B1(n1253), .C0(n1125), .Y(
        n1124) );
  AOI22X1 U192 ( .A0(n1251), .A1(R2[4]), .B0(n1249), .B1(R13[4]), .Y(n1125) );
  OAI221XL U193 ( .A0(n852), .A1(n878), .B0(n818), .B1(n1253), .C0(n1117), .Y(
        n1116) );
  AOI22X1 U194 ( .A0(n1251), .A1(R2[5]), .B0(n1249), .B1(R13[5]), .Y(n1117) );
  OAI221XL U195 ( .A0(n851), .A1(n878), .B0(n817), .B1(n1253), .C0(n1109), .Y(
        n1108) );
  AOI22X1 U196 ( .A0(n1251), .A1(R2[6]), .B0(n1249), .B1(R13[6]), .Y(n1109) );
  OAI221XL U197 ( .A0(n850), .A1(n878), .B0(n816), .B1(n1253), .C0(n1101), .Y(
        n1100) );
  AOI22X1 U198 ( .A0(n1251), .A1(R2[7]), .B0(n1249), .B1(R13[7]), .Y(n1101) );
  OAI221XL U199 ( .A0(n849), .A1(n1255), .B0(n815), .B1(n1253), .C0(n1093), 
        .Y(n1092) );
  AOI22X1 U200 ( .A0(n1251), .A1(R2[8]), .B0(n1249), .B1(R13[8]), .Y(n1093) );
  OAI221XL U201 ( .A0(n848), .A1(n1255), .B0(n814), .B1(n1253), .C0(n1085), 
        .Y(n1084) );
  AOI22X1 U202 ( .A0(n1251), .A1(R2[9]), .B0(n1249), .B1(R13[9]), .Y(n1085) );
  OAI221XL U203 ( .A0(n847), .A1(n1255), .B0(n813), .B1(n879), .C0(n1077), .Y(
        n1076) );
  AOI22X1 U204 ( .A0(n1251), .A1(R2[10]), .B0(n1249), .B1(R13[10]), .Y(n1077)
         );
  OAI221XL U205 ( .A0(n846), .A1(n1255), .B0(n812), .B1(n879), .C0(n1069), .Y(
        n1068) );
  AOI22X1 U206 ( .A0(n1251), .A1(R2[11]), .B0(n1249), .B1(R13[11]), .Y(n1069)
         );
  OAI221XL U207 ( .A0(n840), .A1(n1255), .B0(n806), .B1(n879), .C0(n1021), .Y(
        n1020) );
  AOI22X1 U208 ( .A0(n1252), .A1(R2[17]), .B0(n1250), .B1(R13[17]), .Y(n1021)
         );
  OAI221XL U209 ( .A0(n839), .A1(n1255), .B0(n805), .B1(n879), .C0(n1013), .Y(
        n1012) );
  AOI22X1 U210 ( .A0(n1251), .A1(R2[18]), .B0(n1250), .B1(R13[18]), .Y(n1013)
         );
  OAI221XL U211 ( .A0(n838), .A1(n1255), .B0(n804), .B1(n879), .C0(n1005), .Y(
        n1004) );
  AOI22X1 U212 ( .A0(n1252), .A1(R2[19]), .B0(n1250), .B1(R13[19]), .Y(n1005)
         );
  OAI221XL U213 ( .A0(n837), .A1(n1255), .B0(n803), .B1(n879), .C0(n997), .Y(
        n996) );
  AOI22X1 U214 ( .A0(n1251), .A1(R2[20]), .B0(n1250), .B1(R13[20]), .Y(n997)
         );
  OAI221XL U215 ( .A0(n836), .A1(n878), .B0(n802), .B1(n879), .C0(n989), .Y(
        n988) );
  AOI22X1 U216 ( .A0(n1252), .A1(R2[21]), .B0(n1250), .B1(R13[21]), .Y(n989)
         );
  OAI221XL U217 ( .A0(n835), .A1(n878), .B0(n801), .B1(n1253), .C0(n981), .Y(
        n980) );
  AOI22X1 U218 ( .A0(n1252), .A1(R2[22]), .B0(n1250), .B1(R13[22]), .Y(n981)
         );
  OAI221XL U219 ( .A0(n834), .A1(n878), .B0(n800), .B1(n1253), .C0(n973), .Y(
        n972) );
  AOI22X1 U220 ( .A0(n1251), .A1(R2[23]), .B0(n1250), .B1(R13[23]), .Y(n973)
         );
  OAI221XL U221 ( .A0(n833), .A1(n878), .B0(n799), .B1(n1253), .C0(n965), .Y(
        n964) );
  AOI22X1 U222 ( .A0(n1252), .A1(R2[24]), .B0(n1250), .B1(R13[24]), .Y(n965)
         );
  OAI221XL U223 ( .A0(n832), .A1(n878), .B0(n798), .B1(n879), .C0(n957), .Y(
        n956) );
  AOI22X1 U224 ( .A0(n1252), .A1(R2[25]), .B0(n1249), .B1(R13[25]), .Y(n957)
         );
  OAI221XL U225 ( .A0(n831), .A1(n878), .B0(n797), .B1(n879), .C0(n949), .Y(
        n948) );
  AOI22X1 U226 ( .A0(n1252), .A1(R2[26]), .B0(n1250), .B1(R13[26]), .Y(n949)
         );
  OAI221XL U227 ( .A0(n830), .A1(n878), .B0(n796), .B1(n879), .C0(n941), .Y(
        n940) );
  AOI22X1 U228 ( .A0(n1252), .A1(R2[27]), .B0(n1249), .B1(R13[27]), .Y(n941)
         );
  OAI221XL U229 ( .A0(n829), .A1(n878), .B0(n795), .B1(n879), .C0(n933), .Y(
        n932) );
  AOI22X1 U230 ( .A0(n1252), .A1(R2[28]), .B0(n1250), .B1(R13[28]), .Y(n933)
         );
  OAI221XL U231 ( .A0(n828), .A1(n878), .B0(n794), .B1(n879), .C0(n925), .Y(
        n924) );
  AOI22X1 U232 ( .A0(n1252), .A1(R2[29]), .B0(n1249), .B1(R13[29]), .Y(n925)
         );
  NOR2X1 U233 ( .A(counter_2[3]), .B(counter_2[0]), .Y(n1163) );
  NOR2X1 U234 ( .A(n1281), .B(counter_2[2]), .Y(n872) );
  AND3X2 U235 ( .A(counter_1[0]), .B(n1283), .C(counter_1[1]), .Y(n249) );
  AND3X2 U236 ( .A(n585), .B(n1283), .C(counter_1[1]), .Y(n250) );
  INVX1 U237 ( .A(p_s_flag_in), .Y(n1283) );
  INVX1 U238 ( .A(counter_2[1]), .Y(n1281) );
  AOI22X1 U239 ( .A0(n1244), .A1(R3[12]), .B0(n1241), .B1(R14[12]), .Y(n1062)
         );
  AOI22X1 U240 ( .A0(n1236), .A1(R0[12]), .B0(n1234), .B1(R15[12]), .Y(n1063)
         );
  AOI22X1 U241 ( .A0(n1225), .A1(R1[12]), .B0(n1228), .B1(R12[12]), .Y(n1064)
         );
  AOI22X1 U242 ( .A0(n1244), .A1(R3[13]), .B0(n1241), .B1(R14[13]), .Y(n1054)
         );
  AOI22X1 U243 ( .A0(n1236), .A1(R0[13]), .B0(n1234), .B1(R15[13]), .Y(n1055)
         );
  AOI22X1 U244 ( .A0(n1225), .A1(R1[13]), .B0(n1228), .B1(R12[13]), .Y(n1056)
         );
  AOI22X1 U245 ( .A0(n1244), .A1(R3[14]), .B0(n1241), .B1(R14[14]), .Y(n1046)
         );
  AOI22X1 U246 ( .A0(n1235), .A1(R0[14]), .B0(n1234), .B1(R15[14]), .Y(n1047)
         );
  AOI22X1 U247 ( .A0(n1225), .A1(R1[14]), .B0(n1228), .B1(R12[14]), .Y(n1048)
         );
  AOI22X1 U248 ( .A0(n1244), .A1(R3[15]), .B0(n1241), .B1(n200), .Y(n1038) );
  AOI22X1 U249 ( .A0(n1236), .A1(R0[15]), .B0(n1234), .B1(R15[15]), .Y(n1039)
         );
  AOI22X1 U250 ( .A0(n1225), .A1(R1[15]), .B0(n1228), .B1(n202), .Y(n1040) );
  AOI22X1 U251 ( .A0(n1244), .A1(n1), .B0(n1241), .B1(n7), .Y(n1030) );
  AOI22X1 U252 ( .A0(n1235), .A1(n206), .B0(n1234), .B1(n4), .Y(n1031) );
  AOI22X1 U253 ( .A0(n1225), .A1(n208), .B0(n1228), .B1(n198), .Y(n1032) );
  AOI22X1 U254 ( .A0(n1244), .A1(R3[30]), .B0(n887), .B1(R14[30]), .Y(n918) );
  AOI22X1 U255 ( .A0(n1236), .A1(R0[30]), .B0(n1233), .B1(R15[30]), .Y(n919)
         );
  AOI22X1 U256 ( .A0(n1225), .A1(R1[30]), .B0(n1227), .B1(R12[30]), .Y(n920)
         );
  AOI22X1 U257 ( .A0(n1243), .A1(R3[31]), .B0(n887), .B1(R14[31]), .Y(n910) );
  AOI22X1 U258 ( .A0(n1236), .A1(R0[31]), .B0(n1234), .B1(R15[31]), .Y(n911)
         );
  AOI22X1 U259 ( .A0(n1226), .A1(R1[31]), .B0(n1228), .B1(R12[31]), .Y(n912)
         );
  AOI22X1 U260 ( .A0(n1244), .A1(R3[32]), .B0(n887), .B1(R14[32]), .Y(n902) );
  AOI22X1 U261 ( .A0(n1236), .A1(R0[32]), .B0(n1233), .B1(R15[32]), .Y(n903)
         );
  AOI22X1 U262 ( .A0(n1225), .A1(n190), .B0(n1227), .B1(R12[32]), .Y(n904) );
  AOI22X1 U263 ( .A0(n1243), .A1(R3[33]), .B0(n887), .B1(R14[33]), .Y(n885) );
  AOI22X1 U264 ( .A0(n1236), .A1(n194), .B0(n1234), .B1(n6), .Y(n890) );
  AOI22X1 U265 ( .A0(n1226), .A1(n196), .B0(n1228), .B1(R12[33]), .Y(n895) );
  OAI221XL U266 ( .A0(n845), .A1(n1255), .B0(n811), .B1(n879), .C0(n1061), .Y(
        n1060) );
  AOI22X1 U267 ( .A0(n1252), .A1(R2[12]), .B0(n1250), .B1(R13[12]), .Y(n1061)
         );
  OAI221XL U268 ( .A0(n844), .A1(n1255), .B0(n810), .B1(n1253), .C0(n1053), 
        .Y(n1052) );
  AOI22X1 U269 ( .A0(n1251), .A1(R2[13]), .B0(n1250), .B1(R13[13]), .Y(n1053)
         );
  OAI221XL U270 ( .A0(n843), .A1(n1255), .B0(n809), .B1(n1253), .C0(n1045), 
        .Y(n1044) );
  AOI22X1 U271 ( .A0(n1252), .A1(R2[14]), .B0(n1250), .B1(R13[14]), .Y(n1045)
         );
  OAI221XL U272 ( .A0(n842), .A1(n1255), .B0(n808), .B1(n1253), .C0(n1037), 
        .Y(n1036) );
  AOI22X1 U273 ( .A0(n1251), .A1(R2[15]), .B0(n1250), .B1(n204), .Y(n1037) );
  OAI221XL U274 ( .A0(n841), .A1(n1255), .B0(n807), .B1(n1253), .C0(n1029), 
        .Y(n1028) );
  AOI22X1 U275 ( .A0(n1252), .A1(n188), .B0(n1250), .B1(n186), .Y(n1029) );
  OAI221XL U276 ( .A0(n827), .A1(n1255), .B0(n793), .B1(n879), .C0(n917), .Y(
        n916) );
  AOI22X1 U277 ( .A0(n1252), .A1(R2[30]), .B0(n1250), .B1(R13[30]), .Y(n917)
         );
  OAI221XL U278 ( .A0(n826), .A1(n1255), .B0(n792), .B1(n879), .C0(n909), .Y(
        n908) );
  AOI22X1 U279 ( .A0(n1252), .A1(R2[31]), .B0(n1249), .B1(R13[31]), .Y(n909)
         );
  OAI221XL U280 ( .A0(n825), .A1(n1255), .B0(n791), .B1(n879), .C0(n901), .Y(
        n900) );
  AOI22X1 U281 ( .A0(n1252), .A1(n192), .B0(n1250), .B1(R13[32]), .Y(n901) );
  OAI221XL U282 ( .A0(n824), .A1(n878), .B0(n790), .B1(n879), .C0(n880), .Y(
        n877) );
  AOI22X1 U283 ( .A0(n1252), .A1(R2[33]), .B0(n1249), .B1(R13[33]), .Y(n880)
         );
  AOI22X1 U284 ( .A0(n1243), .A1(R3[29]), .B0(n887), .B1(R14[29]), .Y(n926) );
  AOI22X1 U285 ( .A0(n1236), .A1(R0[29]), .B0(n1233), .B1(R15[29]), .Y(n927)
         );
  AOI22X1 U286 ( .A0(n1226), .A1(R1[29]), .B0(n1228), .B1(R12[29]), .Y(n928)
         );
  INVX1 U287 ( .A(counter_2[2]), .Y(n1282) );
  AOI22X1 U288 ( .A0(n1243), .A1(R3[0]), .B0(n887), .B1(R14[0]), .Y(n1161) );
  AOI22X1 U289 ( .A0(n1235), .A1(R0[0]), .B0(n1233), .B1(R15[0]), .Y(n1162) );
  AOI22X1 U290 ( .A0(n1226), .A1(R1[0]), .B0(n1227), .B1(R12[0]), .Y(n1165) );
  AOI22X1 U291 ( .A0(n1243), .A1(R3[1]), .B0(n887), .B1(R14[1]), .Y(n1150) );
  AOI22X1 U292 ( .A0(n1235), .A1(R0[1]), .B0(n1233), .B1(R15[1]), .Y(n1151) );
  AOI22X1 U293 ( .A0(n1226), .A1(R1[1]), .B0(n1227), .B1(R12[1]), .Y(n1152) );
  AOI22X1 U294 ( .A0(n1243), .A1(R3[2]), .B0(n887), .B1(R14[2]), .Y(n1142) );
  AOI22X1 U295 ( .A0(n1235), .A1(R0[2]), .B0(n1233), .B1(R15[2]), .Y(n1143) );
  AOI22X1 U296 ( .A0(n1226), .A1(R1[2]), .B0(n1227), .B1(R12[2]), .Y(n1144) );
  AOI22X1 U297 ( .A0(n1243), .A1(R3[3]), .B0(n887), .B1(R14[3]), .Y(n1134) );
  AOI22X1 U298 ( .A0(n1235), .A1(R0[3]), .B0(n1233), .B1(R15[3]), .Y(n1135) );
  AOI22X1 U299 ( .A0(n1226), .A1(R1[3]), .B0(n1227), .B1(R12[3]), .Y(n1136) );
  AOI22X1 U300 ( .A0(n1243), .A1(R3[4]), .B0(n887), .B1(R14[4]), .Y(n1126) );
  AOI22X1 U301 ( .A0(n1235), .A1(R0[4]), .B0(n1233), .B1(R15[4]), .Y(n1127) );
  AOI22X1 U302 ( .A0(n1226), .A1(R1[4]), .B0(n1227), .B1(R12[4]), .Y(n1128) );
  AOI22X1 U303 ( .A0(n1243), .A1(R3[5]), .B0(n887), .B1(R14[5]), .Y(n1118) );
  AOI22X1 U304 ( .A0(n1235), .A1(R0[5]), .B0(n1233), .B1(R15[5]), .Y(n1119) );
  AOI22X1 U305 ( .A0(n1226), .A1(R1[5]), .B0(n1227), .B1(R12[5]), .Y(n1120) );
  AOI22X1 U306 ( .A0(n1243), .A1(R3[6]), .B0(n887), .B1(R14[6]), .Y(n1110) );
  AOI22X1 U307 ( .A0(n1235), .A1(R0[6]), .B0(n1233), .B1(R15[6]), .Y(n1111) );
  AOI22X1 U308 ( .A0(n1226), .A1(R1[6]), .B0(n1227), .B1(R12[6]), .Y(n1112) );
  AOI22X1 U309 ( .A0(n1243), .A1(R3[7]), .B0(n887), .B1(R14[7]), .Y(n1102) );
  AOI22X1 U310 ( .A0(n1235), .A1(R0[7]), .B0(n1233), .B1(R15[7]), .Y(n1103) );
  AOI22X1 U311 ( .A0(n1226), .A1(R1[7]), .B0(n1227), .B1(R12[7]), .Y(n1104) );
  AOI22X1 U312 ( .A0(n1243), .A1(R3[8]), .B0(n887), .B1(R14[8]), .Y(n1094) );
  AOI22X1 U313 ( .A0(n1235), .A1(R0[8]), .B0(n1233), .B1(R15[8]), .Y(n1095) );
  AOI22X1 U314 ( .A0(n1226), .A1(R1[8]), .B0(n1227), .B1(R12[8]), .Y(n1096) );
  AOI22X1 U315 ( .A0(n1243), .A1(R3[9]), .B0(n887), .B1(R14[9]), .Y(n1086) );
  AOI22X1 U316 ( .A0(n1235), .A1(R0[9]), .B0(n1233), .B1(R15[9]), .Y(n1087) );
  AOI22X1 U317 ( .A0(n1226), .A1(R1[9]), .B0(n1227), .B1(R12[9]), .Y(n1088) );
  AOI22X1 U318 ( .A0(n1243), .A1(R3[10]), .B0(n887), .B1(R14[10]), .Y(n1078)
         );
  AOI22X1 U319 ( .A0(n1235), .A1(R0[10]), .B0(n1233), .B1(R15[10]), .Y(n1079)
         );
  AOI22X1 U320 ( .A0(n1225), .A1(R1[10]), .B0(n1227), .B1(R12[10]), .Y(n1080)
         );
  AOI22X1 U322 ( .A0(n1243), .A1(R3[11]), .B0(n887), .B1(R14[11]), .Y(n1070)
         );
  AOI22X1 U323 ( .A0(n1235), .A1(R0[11]), .B0(n1233), .B1(R15[11]), .Y(n1071)
         );
  AOI22X1 U325 ( .A0(n1225), .A1(R1[11]), .B0(n1227), .B1(R12[11]), .Y(n1072)
         );
  AOI22X1 U327 ( .A0(n1244), .A1(R3[17]), .B0(n1241), .B1(R14[17]), .Y(n1022)
         );
  AOI22X1 U328 ( .A0(n1236), .A1(R0[17]), .B0(n1234), .B1(R15[17]), .Y(n1023)
         );
  AOI22X1 U329 ( .A0(n1225), .A1(R1[17]), .B0(n1228), .B1(R12[17]), .Y(n1024)
         );
  AOI22X1 U330 ( .A0(n1244), .A1(R3[18]), .B0(n1241), .B1(R14[18]), .Y(n1014)
         );
  AOI22X1 U331 ( .A0(n1236), .A1(R0[18]), .B0(n1234), .B1(R15[18]), .Y(n1015)
         );
  AOI22X1 U332 ( .A0(n1225), .A1(R1[18]), .B0(n1228), .B1(R12[18]), .Y(n1016)
         );
  AOI22X1 U333 ( .A0(n1244), .A1(R3[19]), .B0(n1241), .B1(R14[19]), .Y(n1006)
         );
  AOI22X1 U334 ( .A0(n1235), .A1(R0[19]), .B0(n1234), .B1(R15[19]), .Y(n1007)
         );
  AOI22X1 U335 ( .A0(n1225), .A1(R1[19]), .B0(n1228), .B1(R12[19]), .Y(n1008)
         );
  AOI22X1 U336 ( .A0(n1244), .A1(R3[20]), .B0(n1241), .B1(R14[20]), .Y(n998)
         );
  AOI22X1 U337 ( .A0(n1236), .A1(R0[20]), .B0(n1234), .B1(R15[20]), .Y(n999)
         );
  AOI22X1 U338 ( .A0(n1225), .A1(R1[20]), .B0(n1228), .B1(R12[20]), .Y(n1000)
         );
  AOI22X1 U339 ( .A0(n1244), .A1(R3[21]), .B0(n1241), .B1(R14[21]), .Y(n990)
         );
  AOI22X1 U340 ( .A0(n1235), .A1(R0[21]), .B0(n1234), .B1(R15[21]), .Y(n991)
         );
  AOI22X1 U341 ( .A0(n1225), .A1(R1[21]), .B0(n1228), .B1(R12[21]), .Y(n992)
         );
  AOI22X1 U342 ( .A0(n1244), .A1(R3[22]), .B0(n1241), .B1(R14[22]), .Y(n982)
         );
  AOI22X1 U343 ( .A0(n1236), .A1(R0[22]), .B0(n1234), .B1(R15[22]), .Y(n983)
         );
  AOI22X1 U344 ( .A0(n1226), .A1(R1[22]), .B0(n1228), .B1(R12[22]), .Y(n984)
         );
  AOI22X1 U345 ( .A0(n1244), .A1(R3[23]), .B0(n1241), .B1(R14[23]), .Y(n974)
         );
  AOI22X1 U346 ( .A0(n1235), .A1(R0[23]), .B0(n1234), .B1(R15[23]), .Y(n975)
         );
  AOI22X1 U347 ( .A0(n1226), .A1(R1[23]), .B0(n1228), .B1(R12[23]), .Y(n976)
         );
  AOI22X1 U348 ( .A0(n1244), .A1(R3[24]), .B0(n887), .B1(R14[24]), .Y(n966) );
  AOI22X1 U349 ( .A0(n1236), .A1(R0[24]), .B0(n1234), .B1(R15[24]), .Y(n967)
         );
  AOI22X1 U350 ( .A0(n1226), .A1(R1[24]), .B0(n1227), .B1(R12[24]), .Y(n968)
         );
  AOI22X1 U351 ( .A0(n1243), .A1(R3[25]), .B0(n887), .B1(R14[25]), .Y(n958) );
  AOI22X1 U352 ( .A0(n1236), .A1(R0[25]), .B0(n1233), .B1(R15[25]), .Y(n959)
         );
  AOI22X1 U353 ( .A0(n1225), .A1(R1[25]), .B0(n1228), .B1(R12[25]), .Y(n960)
         );
  AOI22X1 U354 ( .A0(n1244), .A1(R3[26]), .B0(n887), .B1(R14[26]), .Y(n950) );
  AOI22X1 U355 ( .A0(n1236), .A1(R0[26]), .B0(n1234), .B1(R15[26]), .Y(n951)
         );
  AOI22X1 U356 ( .A0(n1226), .A1(R1[26]), .B0(n1227), .B1(R12[26]), .Y(n952)
         );
  AOI22X1 U357 ( .A0(n1243), .A1(R3[27]), .B0(n887), .B1(R14[27]), .Y(n942) );
  AOI22X1 U358 ( .A0(n1236), .A1(R0[27]), .B0(n1233), .B1(R15[27]), .Y(n943)
         );
  AOI22X1 U359 ( .A0(n1225), .A1(R1[27]), .B0(n1228), .B1(R12[27]), .Y(n944)
         );
  AOI22X1 U360 ( .A0(n1244), .A1(R3[28]), .B0(n887), .B1(R14[28]), .Y(n934) );
  AOI22X1 U361 ( .A0(n1236), .A1(R0[28]), .B0(n1234), .B1(R15[28]), .Y(n935)
         );
  AOI22X1 U362 ( .A0(n1225), .A1(R1[28]), .B0(n1227), .B1(R12[28]), .Y(n936)
         );
  OR4X2 U363 ( .A(n1057), .B(n1058), .C(n1059), .D(n1060), .Y(N131) );
  OAI221XL U364 ( .A0(n777), .A1(n1231), .B0(n743), .B1(n1230), .C0(n1064), 
        .Y(n1057) );
  OAI221XL U365 ( .A0(n709), .A1(n1239), .B0(n607), .B1(n889), .C0(n1063), .Y(
        n1058) );
  OAI221XL U366 ( .A0(n641), .A1(n1247), .B0(n675), .B1(n884), .C0(n1062), .Y(
        n1059) );
  OR4X2 U367 ( .A(n1049), .B(n1050), .C(n1051), .D(n1052), .Y(N132) );
  OAI221XL U368 ( .A0(n776), .A1(n1231), .B0(n742), .B1(n1230), .C0(n1056), 
        .Y(n1049) );
  OAI221XL U369 ( .A0(n708), .A1(n1239), .B0(n606), .B1(n889), .C0(n1055), .Y(
        n1050) );
  OAI221XL U370 ( .A0(n640), .A1(n1247), .B0(n674), .B1(n884), .C0(n1054), .Y(
        n1051) );
  OR4X2 U371 ( .A(n1041), .B(n1042), .C(n1043), .D(n1044), .Y(N133) );
  OAI221XL U372 ( .A0(n775), .A1(n1231), .B0(n741), .B1(n1230), .C0(n1048), 
        .Y(n1041) );
  OAI221XL U373 ( .A0(n707), .A1(n1239), .B0(n605), .B1(n889), .C0(n1047), .Y(
        n1042) );
  OAI221XL U374 ( .A0(n639), .A1(n1247), .B0(n673), .B1(n884), .C0(n1046), .Y(
        n1043) );
  OR4X2 U375 ( .A(n1033), .B(n1034), .C(n1035), .D(n1036), .Y(N134) );
  OAI221XL U376 ( .A0(n774), .A1(n1231), .B0(n740), .B1(n1230), .C0(n1040), 
        .Y(n1033) );
  OAI221XL U377 ( .A0(n706), .A1(n1239), .B0(n604), .B1(n889), .C0(n1039), .Y(
        n1034) );
  OAI221XL U378 ( .A0(n638), .A1(n1247), .B0(n672), .B1(n884), .C0(n1038), .Y(
        n1035) );
  OR4X2 U379 ( .A(n1025), .B(n1026), .C(n1027), .D(n1028), .Y(N135) );
  OAI221XL U380 ( .A0(n773), .A1(n1231), .B0(n739), .B1(n1230), .C0(n1032), 
        .Y(n1025) );
  OAI221XL U381 ( .A0(n705), .A1(n1239), .B0(n603), .B1(n889), .C0(n1031), .Y(
        n1026) );
  OAI221XL U382 ( .A0(n637), .A1(n1247), .B0(n671), .B1(n884), .C0(n1030), .Y(
        n1027) );
  OR4X2 U383 ( .A(n921), .B(n922), .C(n923), .D(n924), .Y(N148) );
  OAI221XL U384 ( .A0(n760), .A1(n1231), .B0(n726), .B1(n1229), .C0(n928), .Y(
        n921) );
  OAI221XL U385 ( .A0(n692), .A1(n1239), .B0(n590), .B1(n1237), .C0(n927), .Y(
        n922) );
  OAI221XL U386 ( .A0(n624), .A1(n883), .B0(n658), .B1(n1245), .C0(n926), .Y(
        n923) );
  OR4X2 U387 ( .A(n913), .B(n914), .C(n915), .D(n916), .Y(N149) );
  OAI221XL U388 ( .A0(n759), .A1(n893), .B0(n725), .B1(n1229), .C0(n920), .Y(
        n913) );
  OAI221XL U389 ( .A0(n691), .A1(n888), .B0(n589), .B1(n889), .C0(n919), .Y(
        n914) );
  OAI221XL U390 ( .A0(n623), .A1(n883), .B0(n657), .B1(n1245), .C0(n918), .Y(
        n915) );
  OR4X2 U391 ( .A(n905), .B(n906), .C(n907), .D(n908), .Y(N150) );
  OAI221XL U392 ( .A0(n758), .A1(n893), .B0(n724), .B1(n1229), .C0(n912), .Y(
        n905) );
  OAI221XL U393 ( .A0(n690), .A1(n888), .B0(n588), .B1(n889), .C0(n911), .Y(
        n906) );
  OAI221XL U394 ( .A0(n622), .A1(n883), .B0(n656), .B1(n1245), .C0(n910), .Y(
        n907) );
  OR4X2 U395 ( .A(n897), .B(n898), .C(n899), .D(n900), .Y(N151) );
  OAI221XL U396 ( .A0(n757), .A1(n893), .B0(n723), .B1(n1229), .C0(n904), .Y(
        n897) );
  OAI221XL U397 ( .A0(n689), .A1(n888), .B0(n587), .B1(n889), .C0(n903), .Y(
        n898) );
  OAI221XL U398 ( .A0(n621), .A1(n883), .B0(n655), .B1(n884), .C0(n902), .Y(
        n899) );
  OR4X2 U399 ( .A(n874), .B(n875), .C(n876), .D(n877), .Y(N152) );
  OAI221XL U400 ( .A0(n756), .A1(n893), .B0(n722), .B1(n1229), .C0(n895), .Y(
        n874) );
  OAI221XL U401 ( .A0(n688), .A1(n888), .B0(n586), .B1(n1237), .C0(n890), .Y(
        n875) );
  OAI221XL U402 ( .A0(n620), .A1(n883), .B0(n654), .B1(n1245), .C0(n885), .Y(
        n876) );
  OR4X2 U403 ( .A(n1153), .B(n1154), .C(n1155), .D(n1156), .Y(N119) );
  OAI221XL U404 ( .A0(n789), .A1(n1231), .B0(n755), .B1(n1230), .C0(n1165), 
        .Y(n1153) );
  OAI221XL U405 ( .A0(n721), .A1(n1239), .B0(n619), .B1(n1237), .C0(n1162), 
        .Y(n1154) );
  OAI221XL U406 ( .A0(n653), .A1(n883), .B0(n687), .B1(n1245), .C0(n1161), .Y(
        n1155) );
  OR4X2 U407 ( .A(n1145), .B(n1146), .C(n1147), .D(n1148), .Y(N120) );
  OAI221XL U408 ( .A0(n788), .A1(n1231), .B0(n754), .B1(n1229), .C0(n1152), 
        .Y(n1145) );
  OAI221XL U409 ( .A0(n720), .A1(n1239), .B0(n618), .B1(n1237), .C0(n1151), 
        .Y(n1146) );
  OAI221XL U410 ( .A0(n652), .A1(n1247), .B0(n686), .B1(n1245), .C0(n1150), 
        .Y(n1147) );
  OR4X2 U411 ( .A(n1137), .B(n1138), .C(n1139), .D(n1140), .Y(N121) );
  OAI221XL U412 ( .A0(n787), .A1(n893), .B0(n753), .B1(n1230), .C0(n1144), .Y(
        n1137) );
  OAI221XL U413 ( .A0(n719), .A1(n888), .B0(n617), .B1(n1237), .C0(n1143), .Y(
        n1138) );
  OAI221XL U414 ( .A0(n651), .A1(n883), .B0(n685), .B1(n1245), .C0(n1142), .Y(
        n1139) );
  OR4X2 U415 ( .A(n1129), .B(n1130), .C(n1131), .D(n1132), .Y(N122) );
  OAI221XL U416 ( .A0(n786), .A1(n893), .B0(n752), .B1(n1229), .C0(n1136), .Y(
        n1129) );
  OAI221XL U417 ( .A0(n718), .A1(n888), .B0(n616), .B1(n1237), .C0(n1135), .Y(
        n1130) );
  OAI221XL U418 ( .A0(n650), .A1(n883), .B0(n684), .B1(n1245), .C0(n1134), .Y(
        n1131) );
  OR4X2 U419 ( .A(n1121), .B(n1122), .C(n1123), .D(n1124), .Y(N123) );
  OAI221XL U420 ( .A0(n785), .A1(n893), .B0(n751), .B1(n1230), .C0(n1128), .Y(
        n1121) );
  OAI221XL U421 ( .A0(n717), .A1(n888), .B0(n615), .B1(n1237), .C0(n1127), .Y(
        n1122) );
  OAI221XL U422 ( .A0(n649), .A1(n883), .B0(n683), .B1(n1245), .C0(n1126), .Y(
        n1123) );
  OR4X2 U423 ( .A(n1113), .B(n1114), .C(n1115), .D(n1116), .Y(N124) );
  OAI221XL U424 ( .A0(n784), .A1(n893), .B0(n750), .B1(n1229), .C0(n1120), .Y(
        n1113) );
  OAI221XL U425 ( .A0(n716), .A1(n888), .B0(n614), .B1(n1237), .C0(n1119), .Y(
        n1114) );
  OAI221XL U426 ( .A0(n648), .A1(n883), .B0(n682), .B1(n1245), .C0(n1118), .Y(
        n1115) );
  OR4X2 U427 ( .A(n1105), .B(n1106), .C(n1107), .D(n1108), .Y(N125) );
  OAI221XL U428 ( .A0(n783), .A1(n893), .B0(n749), .B1(n1230), .C0(n1112), .Y(
        n1105) );
  OAI221XL U429 ( .A0(n715), .A1(n888), .B0(n613), .B1(n1237), .C0(n1111), .Y(
        n1106) );
  OAI221XL U430 ( .A0(n647), .A1(n883), .B0(n681), .B1(n1245), .C0(n1110), .Y(
        n1107) );
  OR4X2 U431 ( .A(n1097), .B(n1098), .C(n1099), .D(n1100), .Y(N126) );
  OAI221XL U432 ( .A0(n782), .A1(n893), .B0(n748), .B1(n1229), .C0(n1104), .Y(
        n1097) );
  OAI221XL U433 ( .A0(n714), .A1(n888), .B0(n612), .B1(n1237), .C0(n1103), .Y(
        n1098) );
  OAI221XL U434 ( .A0(n646), .A1(n883), .B0(n680), .B1(n1245), .C0(n1102), .Y(
        n1099) );
  OR4X2 U435 ( .A(n1089), .B(n1090), .C(n1091), .D(n1092), .Y(N127) );
  OAI221XL U436 ( .A0(n781), .A1(n1231), .B0(n747), .B1(n1230), .C0(n1096), 
        .Y(n1089) );
  OAI221XL U437 ( .A0(n713), .A1(n1239), .B0(n611), .B1(n1237), .C0(n1095), 
        .Y(n1090) );
  OAI221XL U438 ( .A0(n645), .A1(n1247), .B0(n679), .B1(n1245), .C0(n1094), 
        .Y(n1091) );
  OR4X2 U439 ( .A(n1081), .B(n1082), .C(n1083), .D(n1084), .Y(N128) );
  OAI221XL U440 ( .A0(n780), .A1(n1231), .B0(n746), .B1(n1229), .C0(n1088), 
        .Y(n1081) );
  OAI221XL U441 ( .A0(n712), .A1(n1239), .B0(n610), .B1(n1237), .C0(n1087), 
        .Y(n1082) );
  OAI221XL U442 ( .A0(n644), .A1(n1247), .B0(n678), .B1(n1245), .C0(n1086), 
        .Y(n1083) );
  OR4X2 U443 ( .A(n1073), .B(n1074), .C(n1075), .D(n1076), .Y(N129) );
  OAI221XL U444 ( .A0(n779), .A1(n1231), .B0(n745), .B1(n1230), .C0(n1080), 
        .Y(n1073) );
  OAI221XL U445 ( .A0(n711), .A1(n1239), .B0(n609), .B1(n889), .C0(n1079), .Y(
        n1074) );
  OAI221XL U446 ( .A0(n643), .A1(n1247), .B0(n677), .B1(n884), .C0(n1078), .Y(
        n1075) );
  OR4X2 U447 ( .A(n1065), .B(n1066), .C(n1067), .D(n1068), .Y(N130) );
  OAI221XL U448 ( .A0(n778), .A1(n1231), .B0(n744), .B1(n1230), .C0(n1072), 
        .Y(n1065) );
  OAI221XL U449 ( .A0(n710), .A1(n1239), .B0(n608), .B1(n889), .C0(n1071), .Y(
        n1066) );
  OAI221XL U450 ( .A0(n642), .A1(n1247), .B0(n676), .B1(n884), .C0(n1070), .Y(
        n1067) );
  OR4X2 U451 ( .A(n1017), .B(n1018), .C(n1019), .D(n1020), .Y(N136) );
  OAI221XL U452 ( .A0(n772), .A1(n1231), .B0(n738), .B1(n1230), .C0(n1024), 
        .Y(n1017) );
  OAI221XL U453 ( .A0(n704), .A1(n1239), .B0(n602), .B1(n889), .C0(n1023), .Y(
        n1018) );
  OAI221XL U454 ( .A0(n636), .A1(n1247), .B0(n670), .B1(n884), .C0(n1022), .Y(
        n1019) );
  OR4X2 U455 ( .A(n1009), .B(n1010), .C(n1011), .D(n1012), .Y(N137) );
  OAI221XL U456 ( .A0(n771), .A1(n1231), .B0(n737), .B1(n1230), .C0(n1016), 
        .Y(n1009) );
  OAI221XL U457 ( .A0(n703), .A1(n1239), .B0(n601), .B1(n1237), .C0(n1015), 
        .Y(n1010) );
  OAI221XL U458 ( .A0(n635), .A1(n1247), .B0(n669), .B1(n884), .C0(n1014), .Y(
        n1011) );
  OR4X2 U459 ( .A(n1001), .B(n1002), .C(n1003), .D(n1004), .Y(N138) );
  OAI221XL U460 ( .A0(n770), .A1(n1231), .B0(n736), .B1(n1230), .C0(n1008), 
        .Y(n1001) );
  OAI221XL U461 ( .A0(n702), .A1(n1239), .B0(n600), .B1(n1237), .C0(n1007), 
        .Y(n1002) );
  OAI221XL U462 ( .A0(n634), .A1(n1247), .B0(n668), .B1(n884), .C0(n1006), .Y(
        n1003) );
  OR4X2 U463 ( .A(n993), .B(n994), .C(n995), .D(n996), .Y(N139) );
  OAI221XL U464 ( .A0(n769), .A1(n1231), .B0(n735), .B1(n1230), .C0(n1000), 
        .Y(n993) );
  OAI221XL U465 ( .A0(n701), .A1(n1239), .B0(n599), .B1(n1237), .C0(n999), .Y(
        n994) );
  OAI221XL U466 ( .A0(n633), .A1(n1247), .B0(n667), .B1(n1245), .C0(n998), .Y(
        n995) );
  OR4X2 U467 ( .A(n985), .B(n986), .C(n987), .D(n988), .Y(N140) );
  OAI221XL U468 ( .A0(n768), .A1(n893), .B0(n734), .B1(n1230), .C0(n992), .Y(
        n985) );
  OAI221XL U469 ( .A0(n700), .A1(n888), .B0(n598), .B1(n1237), .C0(n991), .Y(
        n986) );
  OAI221XL U470 ( .A0(n632), .A1(n883), .B0(n666), .B1(n884), .C0(n990), .Y(
        n987) );
  OR4X2 U471 ( .A(n977), .B(n978), .C(n979), .D(n980), .Y(N141) );
  OAI221XL U472 ( .A0(n767), .A1(n893), .B0(n733), .B1(n1229), .C0(n984), .Y(
        n977) );
  OAI221XL U473 ( .A0(n699), .A1(n888), .B0(n597), .B1(n1237), .C0(n983), .Y(
        n978) );
  OAI221XL U474 ( .A0(n631), .A1(n883), .B0(n665), .B1(n1245), .C0(n982), .Y(
        n979) );
  OR4X2 U475 ( .A(n969), .B(n970), .C(n971), .D(n972), .Y(N142) );
  OAI221XL U476 ( .A0(n766), .A1(n893), .B0(n732), .B1(n1229), .C0(n976), .Y(
        n969) );
  OAI221XL U477 ( .A0(n698), .A1(n888), .B0(n596), .B1(n889), .C0(n975), .Y(
        n970) );
  OAI221XL U478 ( .A0(n630), .A1(n883), .B0(n664), .B1(n1245), .C0(n974), .Y(
        n971) );
  OR4X2 U479 ( .A(n961), .B(n962), .C(n963), .D(n964), .Y(N143) );
  OAI221XL U480 ( .A0(n765), .A1(n893), .B0(n731), .B1(n1229), .C0(n968), .Y(
        n961) );
  OAI221XL U481 ( .A0(n697), .A1(n888), .B0(n595), .B1(n889), .C0(n967), .Y(
        n962) );
  OAI221XL U482 ( .A0(n629), .A1(n883), .B0(n663), .B1(n884), .C0(n966), .Y(
        n963) );
  OR4X2 U483 ( .A(n953), .B(n954), .C(n955), .D(n956), .Y(N144) );
  OAI221XL U484 ( .A0(n764), .A1(n893), .B0(n730), .B1(n1229), .C0(n960), .Y(
        n953) );
  OAI221XL U485 ( .A0(n696), .A1(n888), .B0(n594), .B1(n889), .C0(n959), .Y(
        n954) );
  OAI221XL U486 ( .A0(n628), .A1(n883), .B0(n662), .B1(n884), .C0(n958), .Y(
        n955) );
  OR4X2 U487 ( .A(n945), .B(n946), .C(n947), .D(n948), .Y(N145) );
  OAI221XL U488 ( .A0(n763), .A1(n893), .B0(n729), .B1(n1229), .C0(n952), .Y(
        n945) );
  OAI221XL U489 ( .A0(n695), .A1(n888), .B0(n593), .B1(n889), .C0(n951), .Y(
        n946) );
  OAI221XL U490 ( .A0(n627), .A1(n1247), .B0(n661), .B1(n884), .C0(n950), .Y(
        n947) );
  OR4X2 U491 ( .A(n937), .B(n938), .C(n939), .D(n940), .Y(N146) );
  OAI221XL U492 ( .A0(n762), .A1(n893), .B0(n728), .B1(n1229), .C0(n944), .Y(
        n937) );
  OAI221XL U493 ( .A0(n694), .A1(n888), .B0(n592), .B1(n889), .C0(n943), .Y(
        n938) );
  OAI221XL U494 ( .A0(n626), .A1(n1247), .B0(n660), .B1(n884), .C0(n942), .Y(
        n939) );
  OR4X2 U495 ( .A(n929), .B(n930), .C(n931), .D(n932), .Y(N147) );
  OAI221XL U496 ( .A0(n761), .A1(n1231), .B0(n727), .B1(n1229), .C0(n936), .Y(
        n929) );
  OAI221XL U497 ( .A0(n693), .A1(n1239), .B0(n591), .B1(n889), .C0(n935), .Y(
        n930) );
  OAI221XL U498 ( .A0(n625), .A1(n1247), .B0(n659), .B1(n884), .C0(n934), .Y(
        n931) );
  OR3XL U499 ( .A(counter_1[1]), .B(p_s_flag_in), .C(n585), .Y(n251) );
  INVX1 U500 ( .A(n871), .Y(n1280) );
  AOI221X1 U501 ( .A0(counter_2[0]), .A1(n872), .B0(n862), .B1(counter_2[2]), 
        .C0(n873), .Y(n871) );
  NAND2X1 U502 ( .A(n868), .B(n869), .Y(N52) );
  OAI2BB1X1 U503 ( .A0N(n870), .A1N(counter_2[0]), .B0(counter_2[3]), .Y(n869)
         );
  XNOR2X1 U504 ( .A(counter_1[1]), .B(n585), .Y(N26) );
  XNOR2X1 U505 ( .A(n1281), .B(counter_2[0]), .Y(N50) );
endmodule


module fft ( clk, rst_n, data_in, data_out );
  input [33:0] data_in;
  output [33:0] data_out;
  input clk, rst_n;
  wire   s_p_flag, mux_flag, demux_flag, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48;
  wire   [2:0] rotation;
  wire   [135:0] data_1;
  wire   [135:0] data_2;
  wire   [135:0] data_4;
  wire   [135:0] data_3;

  ctrl ctrl0 ( .clk(clk), .rst_n(rst_n), .s_p_flag_in(s_p_flag), .mux_flag(
        mux_flag), .rotation(rotation), .demux_flag(demux_flag) );
  s_p s_p0 ( .clk(clk), .rst_n(rst_n), .data_in_1(data_in), .data_out_1(data_1), .s_p_flag_out(s_p_flag) );
  mux mux0 ( .mux_flag(mux_flag), .clk(clk), .rst_n(rst_n), .data_in_1(data_2), 
        .data_in_2(data_1), .data_out(data_3), .data_in_3_33_(n45), 
        .data_in_3_32_(n42), .data_in_3_31_(n41), .data_in_3_30_(n27), 
        .data_in_3_29_(n2), .data_in_3_28_(data_4[28]), .data_in_3_27_(n14), 
        .data_in_3_26_(n44), .data_in_3_25_(data_4[25]), .data_in_3_24_(n12), 
        .data_in_3_23_(data_4[23]), .data_in_3_22_(data_4[22]), 
        .data_in_3_21_(data_4[21]), .data_in_3_20_(data_4[20]), 
        .data_in_3_19_(data_4[19]), .data_in_3_18_(data_4[18]), 
        .data_in_3_17_(data_4[17]), .data_in_3_16_(n46), .data_in_3_15_(n48), 
        .data_in_3_14_(n36), .data_in_3_13_(data_4[13]), .data_in_3_12_(
        data_4[12]), .data_in_3_11_(n22), .data_in_3_10_(n13), .data_in_3_9_(
        data_4[9]), .data_in_3_8_(n31), .data_in_3_7_(data_4[7]), 
        .data_in_3_6_(n40), .data_in_3_5_(n7), .data_in_3_4_(n9), 
        .data_in_3_3_(data_4[3]), .data_in_3_2_(data_4[2]), .data_in_3_1_(
        data_4[1]), .data_in_3_0_(data_4[0]) );
  butterfly butterfly0 ( .calc_in({data_3[135:88], n34, data_3[86:0]}), 
        .rotation(rotation), .calc_out(data_4) );
  reg1 reg10 ( .clk(clk), .rst_n(rst_n), .data_in_2({n33, data_4[134:131], n11, 
        data_4[129:128], n19, data_4[126:112], n29, n21, data_4[109:95], n25, 
        n18, data_4[92:82], n5, data_4[80:79], n17, data_4[77], n26, 
        data_4[75:67], n47, data_4[65:62], n23, n35, n20, data_4[58:49], n38, 
        n37, data_4[46:44], n1, n24, data_4[41:32], n41, data_4[30], n32, 
        data_4[28], n16, n44, data_4[25:11], n15, data_4[9], n31, data_4[7], 
        n40, n7, n9, data_4[3:0]}), .reg_datain_flag(demux_flag), .data_out_2(
        data_2) );
  p_s p_s0 ( .clk(clk), .rst_n(rst_n), .data_in_3({n33, data_4[134:128], n19, 
        data_4[126:112], n29, n21, data_4[109:95], n25, n18, data_4[92:82], n3, 
        data_4[80:79], n17, data_4[77], n26, data_4[75:67], n47, data_4[65:62], 
        n23, n35, n20, data_4[58:49], n38, n37, data_4[46:44], n1, n24, 
        data_4[41:32], n41, data_4[30], n32, data_4[28], n14, n44, data_4[25], 
        n12, data_4[23:11], n15, data_4[9], n31, data_4[7], n40, n7, n9, 
        data_4[3:0]}), .p_s_flag_in(demux_flag), .data_out_3(data_out) );
  BUFX12 U1 ( .A(data_4[93]), .Y(n18) );
  BUFX12 U2 ( .A(data_4[10]), .Y(n15) );
  BUFX8 U3 ( .A(data_4[43]), .Y(n1) );
  BUFX16 U4 ( .A(data_4[29]), .Y(n32) );
  DLY1X1 U5 ( .A(n32), .Y(n2) );
  INVX8 U6 ( .A(n4), .Y(n3) );
  CLKINVX8 U7 ( .A(data_4[81]), .Y(n4) );
  INVX8 U8 ( .A(n4), .Y(n5) );
  DLY1X1 U9 ( .A(data_4[46]), .Y(n28) );
  BUFX20 U10 ( .A(data_4[135]), .Y(n33) );
  BUFX12 U11 ( .A(data_4[60]), .Y(n35) );
  BUFX12 U12 ( .A(data_4[127]), .Y(n19) );
  CLKINVX4 U13 ( .A(data_4[5]), .Y(n6) );
  INVX8 U14 ( .A(n6), .Y(n7) );
  CLKINVX4 U15 ( .A(data_4[4]), .Y(n8) );
  INVX8 U16 ( .A(n8), .Y(n9) );
  BUFX12 U17 ( .A(data_4[76]), .Y(n26) );
  CLKINVX8 U18 ( .A(data_4[130]), .Y(n10) );
  INVX8 U19 ( .A(n10), .Y(n11) );
  BUFX8 U20 ( .A(data_4[24]), .Y(n12) );
  CLKINVX8 U21 ( .A(data_4[26]), .Y(n43) );
  BUFX16 U22 ( .A(data_4[61]), .Y(n23) );
  DLY1X1 U23 ( .A(n15), .Y(n13) );
  BUFX8 U24 ( .A(data_4[27]), .Y(n14) );
  BUFX8 U25 ( .A(data_4[27]), .Y(n16) );
  BUFX8 U26 ( .A(data_4[78]), .Y(n17) );
  BUFX8 U27 ( .A(data_4[59]), .Y(n20) );
  BUFX8 U28 ( .A(data_4[110]), .Y(n21) );
  DLY1X1 U29 ( .A(data_4[11]), .Y(n22) );
  BUFX8 U30 ( .A(data_4[42]), .Y(n24) );
  BUFX8 U31 ( .A(data_4[94]), .Y(n25) );
  DLY1X1 U32 ( .A(data_4[30]), .Y(n27) );
  BUFX20 U33 ( .A(data_4[31]), .Y(n41) );
  BUFX8 U34 ( .A(data_4[111]), .Y(n29) );
  CLKINVX4 U35 ( .A(data_4[8]), .Y(n30) );
  INVX8 U36 ( .A(n30), .Y(n31) );
  BUFX12 U37 ( .A(data_3[87]), .Y(n34) );
  BUFX16 U38 ( .A(data_4[47]), .Y(n37) );
  DLY1X1 U39 ( .A(data_4[14]), .Y(n36) );
  BUFX20 U40 ( .A(data_4[48]), .Y(n38) );
  CLKINVX4 U41 ( .A(data_4[6]), .Y(n39) );
  INVX8 U42 ( .A(n39), .Y(n40) );
  BUFX16 U43 ( .A(data_4[66]), .Y(n47) );
  DLY1X1 U44 ( .A(data_4[32]), .Y(n42) );
  INVX8 U45 ( .A(n43), .Y(n44) );
  DLY1X1 U46 ( .A(data_4[33]), .Y(n45) );
  DLY1X1 U47 ( .A(data_4[16]), .Y(n46) );
  DLY1X1 U48 ( .A(data_4[15]), .Y(n48) );
endmodule


module fft_chip ( clk, rst_n, data_in, data_out );
  input [33:0] data_in;
  output [33:0] data_out;
  input clk, rst_n;
  wire   net_clk, net_rst_n;
  wire   [33:0] net_data_in;
  wire   [33:0] net_data_out;

  PIW PIW_clk ( .PAD(clk), .C(net_clk) );
  PIW PIW_rst_n ( .PAD(rst_n), .C(net_rst_n) );
  PIW PIW_data_in0 ( .PAD(data_in[0]), .C(net_data_in[0]) );
  PIW PIW_data_in1 ( .PAD(data_in[1]), .C(net_data_in[1]) );
  PIW PIW_data_in2 ( .PAD(data_in[2]), .C(net_data_in[2]) );
  PIW PIW_data_in3 ( .PAD(data_in[3]), .C(net_data_in[3]) );
  PIW PIW_data_in4 ( .PAD(data_in[4]), .C(net_data_in[4]) );
  PIW PIW_data_in5 ( .PAD(data_in[5]), .C(net_data_in[5]) );
  PIW PIW_data_in6 ( .PAD(data_in[6]), .C(net_data_in[6]) );
  PIW PIW_data_in7 ( .PAD(data_in[7]), .C(net_data_in[7]) );
  PIW PIW_data_in8 ( .PAD(data_in[8]), .C(net_data_in[8]) );
  PIW PIW_data_in9 ( .PAD(data_in[9]), .C(net_data_in[9]) );
  PIW PIW_data_in10 ( .PAD(data_in[10]), .C(net_data_in[10]) );
  PIW PIW_data_in11 ( .PAD(data_in[11]), .C(net_data_in[11]) );
  PIW PIW_data_in12 ( .PAD(data_in[12]), .C(net_data_in[12]) );
  PIW PIW_data_in13 ( .PAD(data_in[13]), .C(net_data_in[13]) );
  PIW PIW_data_in14 ( .PAD(data_in[14]), .C(net_data_in[14]) );
  PIW PIW_data_in15 ( .PAD(data_in[15]), .C(net_data_in[15]) );
  PIW PIW_data_in16 ( .PAD(data_in[16]), .C(net_data_in[16]) );
  PIW PIW_data_in17 ( .PAD(data_in[17]), .C(net_data_in[17]) );
  PIW PIW_data_in18 ( .PAD(data_in[18]), .C(net_data_in[18]) );
  PIW PIW_data_in19 ( .PAD(data_in[19]), .C(net_data_in[19]) );
  PIW PIW_data_in20 ( .PAD(data_in[20]), .C(net_data_in[20]) );
  PIW PIW_data_in21 ( .PAD(data_in[21]), .C(net_data_in[21]) );
  PIW PIW_data_in22 ( .PAD(data_in[22]), .C(net_data_in[22]) );
  PIW PIW_data_in23 ( .PAD(data_in[23]), .C(net_data_in[23]) );
  PIW PIW_data_in24 ( .PAD(data_in[24]), .C(net_data_in[24]) );
  PIW PIW_data_in25 ( .PAD(data_in[25]), .C(net_data_in[25]) );
  PIW PIW_data_in26 ( .PAD(data_in[26]), .C(net_data_in[26]) );
  PIW PIW_data_in27 ( .PAD(data_in[27]), .C(net_data_in[27]) );
  PIW PIW_data_in28 ( .PAD(data_in[28]), .C(net_data_in[28]) );
  PIW PIW_data_in29 ( .PAD(data_in[29]), .C(net_data_in[29]) );
  PIW PIW_data_in30 ( .PAD(data_in[30]), .C(net_data_in[30]) );
  PIW PIW_data_in31 ( .PAD(data_in[31]), .C(net_data_in[31]) );
  PIW PIW_data_in32 ( .PAD(data_in[32]), .C(net_data_in[32]) );
  PIW PIW_data_in33 ( .PAD(data_in[33]), .C(net_data_in[33]) );
  PO8W PO8W_data_out0 ( .I(net_data_out[0]), .PAD(data_out[0]) );
  PO8W PO8W_data_out1 ( .I(net_data_out[1]), .PAD(data_out[1]) );
  PO8W PO8W_data_out2 ( .I(net_data_out[2]), .PAD(data_out[2]) );
  PO8W PO8W_data_out3 ( .I(net_data_out[3]), .PAD(data_out[3]) );
  PO8W PO8W_data_out4 ( .I(net_data_out[4]), .PAD(data_out[4]) );
  PO8W PO8W_data_out5 ( .I(net_data_out[5]), .PAD(data_out[5]) );
  PO8W PO8W_data_out6 ( .I(net_data_out[6]), .PAD(data_out[6]) );
  PO8W PO8W_data_out7 ( .I(net_data_out[7]), .PAD(data_out[7]) );
  PO8W PO8W_data_out8 ( .I(net_data_out[8]), .PAD(data_out[8]) );
  PO8W PO8W_data_out9 ( .I(net_data_out[9]), .PAD(data_out[9]) );
  PO8W PO8W_data_out10 ( .I(net_data_out[10]), .PAD(data_out[10]) );
  PO8W PO8W_data_out11 ( .I(net_data_out[11]), .PAD(data_out[11]) );
  PO8W PO8W_data_out12 ( .I(net_data_out[12]), .PAD(data_out[12]) );
  PO8W PO8W_data_out13 ( .I(net_data_out[13]), .PAD(data_out[13]) );
  PO8W PO8W_data_out14 ( .I(net_data_out[14]), .PAD(data_out[14]) );
  PO8W PO8W_data_out15 ( .I(net_data_out[15]), .PAD(data_out[15]) );
  PO8W PO8W_data_out16 ( .I(net_data_out[16]), .PAD(data_out[16]) );
  PO8W PO8W_data_out17 ( .I(net_data_out[17]), .PAD(data_out[17]) );
  PO8W PO8W_data_out18 ( .I(net_data_out[18]), .PAD(data_out[18]) );
  PO8W PO8W_data_out19 ( .I(net_data_out[19]), .PAD(data_out[19]) );
  PO8W PO8W_data_out20 ( .I(net_data_out[20]), .PAD(data_out[20]) );
  PO8W PO8W_data_out21 ( .I(net_data_out[21]), .PAD(data_out[21]) );
  PO8W PO8W_data_out22 ( .I(net_data_out[22]), .PAD(data_out[22]) );
  PO8W PO8W_data_out23 ( .I(net_data_out[23]), .PAD(data_out[23]) );
  PO8W PO8W_data_out24 ( .I(net_data_out[24]), .PAD(data_out[24]) );
  PO8W PO8W_data_out25 ( .I(net_data_out[25]), .PAD(data_out[25]) );
  PO8W PO8W_data_out26 ( .I(net_data_out[26]), .PAD(data_out[26]) );
  PO8W PO8W_data_out27 ( .I(net_data_out[27]), .PAD(data_out[27]) );
  PO8W PO8W_data_out28 ( .I(net_data_out[28]), .PAD(data_out[28]) );
  PO8W PO8W_data_out29 ( .I(net_data_out[29]), .PAD(data_out[29]) );
  PO8W PO8W_data_out30 ( .I(net_data_out[30]), .PAD(data_out[30]) );
  PO8W PO8W_data_out31 ( .I(net_data_out[31]), .PAD(data_out[31]) );
  PO8W PO8W_data_out32 ( .I(net_data_out[32]), .PAD(data_out[32]) );
  PO8W PO8W_data_out33 ( .I(net_data_out[33]), .PAD(data_out[33]) );
  fft inst_fft ( .clk(net_clk), .rst_n(net_rst_n), .data_in(net_data_in), 
        .data_out(net_data_out) );
endmodule

