
module ctrl ( clk, rst_n, s_p_flag_in, mux_flag, rotation, demux_flag );
  output [2:0] rotation;
  input clk, rst_n, s_p_flag_in;
  output mux_flag, demux_flag;
  wire   N17, N18, N19, n3, n4, n1, n2;
  wire   [2:0] core_tick;

  DFFRHQX4 mux_flag_reg ( .D(core_tick[2]), .CK(clk), .RN(rst_n), .Q(mux_flag)
         );
  DFFRHQX4 rotation_reg_2_ ( .D(core_tick[2]), .CK(clk), .RN(rst_n), .Q(
        rotation[2]) );
  DFFRHQX4 rotation_reg_1_ ( .D(core_tick[1]), .CK(clk), .RN(rst_n), .Q(
        rotation[1]) );
  DFFRHQX4 rotation_reg_0_ ( .D(core_tick[0]), .CK(clk), .RN(rst_n), .Q(
        rotation[0]) );
  DFFRHQX1 core_tick_reg_2_ ( .D(N19), .CK(clk), .RN(rst_n), .Q(core_tick[2])
         );
  DFFRHQX1 core_tick_reg_1_ ( .D(N18), .CK(clk), .RN(rst_n), .Q(core_tick[1])
         );
  DFFRHQX1 core_tick_reg_0_ ( .D(N17), .CK(clk), .RN(rst_n), .Q(core_tick[0])
         );
  DFFRHQX1 demux_flag_reg ( .D(n2), .CK(clk), .RN(rst_n), .Q(demux_flag) );
  AOI21X1 U3 ( .A0(n4), .A1(n1), .B0(core_tick[0]), .Y(N17) );
  NOR2X1 U4 ( .A(s_p_flag_in), .B(core_tick[2]), .Y(n4) );
  INVX1 U5 ( .A(core_tick[1]), .Y(n1) );
  INVX1 U6 ( .A(core_tick[2]), .Y(n2) );
  XOR2X1 U7 ( .A(core_tick[1]), .B(core_tick[0]), .Y(N18) );
  XOR2X1 U8 ( .A(n2), .B(n3), .Y(N19) );
  NAND2X1 U9 ( .A(core_tick[1]), .B(core_tick[0]), .Y(n3) );
endmodule


module s_p ( clk, rst_n, data_in_1, data_out_1, s_p_flag_out );
  input [33:0] data_in_1;
  output [135:0] data_out_1;
  input clk, rst_n;
  output s_p_flag_out;
  wire   N13, N14, N15, N171, n550, n551, n552, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006;
  wire   [3:0] counter;
  wire   [33:0] R15;
  wire   [33:0] R11;
  wire   [33:0] R7;
  wire   [33:0] R3;
  wire   [33:0] R12;
  wire   [33:0] R8;
  wire   [33:0] R4;
  wire   [33:0] R0;
  wire   [33:0] R13;
  wire   [33:0] R9;
  wire   [33:0] R5;
  wire   [33:0] R1;
  wire   [33:0] R14;
  wire   [33:0] R10;
  wire   [33:0] R6;
  wire   [33:0] R2;

  EDFFX1 R13_reg_33_ ( .D(data_in_1[33]), .E(n980), .CK(clk), .Q(R13[33]) );
  EDFFX1 R13_reg_32_ ( .D(data_in_1[32]), .E(n980), .CK(clk), .Q(R13[32]) );
  EDFFX1 R13_reg_31_ ( .D(data_in_1[31]), .E(n980), .CK(clk), .Q(R13[31]) );
  EDFFX1 R13_reg_30_ ( .D(data_in_1[30]), .E(n980), .CK(clk), .Q(R13[30]) );
  EDFFX1 R13_reg_29_ ( .D(data_in_1[29]), .E(n980), .CK(clk), .Q(R13[29]) );
  EDFFX1 R13_reg_28_ ( .D(data_in_1[28]), .E(n980), .CK(clk), .Q(R13[28]) );
  EDFFX1 R13_reg_27_ ( .D(data_in_1[27]), .E(n980), .CK(clk), .Q(R13[27]) );
  EDFFX1 R13_reg_26_ ( .D(data_in_1[26]), .E(n980), .CK(clk), .Q(R13[26]) );
  EDFFX1 R13_reg_25_ ( .D(data_in_1[25]), .E(n980), .CK(clk), .Q(R13[25]) );
  EDFFX1 R13_reg_24_ ( .D(data_in_1[24]), .E(n980), .CK(clk), .Q(R13[24]) );
  EDFFX1 R13_reg_23_ ( .D(data_in_1[23]), .E(n980), .CK(clk), .Q(R13[23]) );
  EDFFX1 R13_reg_22_ ( .D(data_in_1[22]), .E(n980), .CK(clk), .Q(R13[22]) );
  EDFFX1 R13_reg_21_ ( .D(data_in_1[21]), .E(n980), .CK(clk), .Q(R13[21]) );
  EDFFX1 R13_reg_20_ ( .D(data_in_1[20]), .E(n980), .CK(clk), .Q(R13[20]) );
  EDFFX1 R13_reg_19_ ( .D(data_in_1[19]), .E(n980), .CK(clk), .Q(R13[19]) );
  EDFFX1 R13_reg_18_ ( .D(data_in_1[18]), .E(n980), .CK(clk), .Q(R13[18]) );
  EDFFX1 R13_reg_17_ ( .D(data_in_1[17]), .E(n980), .CK(clk), .Q(R13[17]) );
  EDFFX1 R13_reg_16_ ( .D(data_in_1[16]), .E(n980), .CK(clk), .Q(R13[16]) );
  EDFFX1 R13_reg_15_ ( .D(data_in_1[15]), .E(n980), .CK(clk), .Q(R13[15]) );
  EDFFX1 R13_reg_14_ ( .D(data_in_1[14]), .E(n980), .CK(clk), .Q(R13[14]) );
  EDFFX1 R13_reg_13_ ( .D(data_in_1[13]), .E(n980), .CK(clk), .Q(R13[13]) );
  EDFFX1 R13_reg_12_ ( .D(data_in_1[12]), .E(n980), .CK(clk), .Q(R13[12]) );
  EDFFX1 R13_reg_11_ ( .D(data_in_1[11]), .E(n980), .CK(clk), .Q(R13[11]) );
  EDFFX1 R13_reg_10_ ( .D(data_in_1[10]), .E(n980), .CK(clk), .Q(R13[10]) );
  EDFFX1 R13_reg_9_ ( .D(data_in_1[9]), .E(n980), .CK(clk), .Q(R13[9]) );
  EDFFX1 R13_reg_8_ ( .D(data_in_1[8]), .E(n980), .CK(clk), .Q(R13[8]) );
  EDFFX1 R13_reg_7_ ( .D(data_in_1[7]), .E(n980), .CK(clk), .Q(R13[7]) );
  EDFFX1 R13_reg_6_ ( .D(data_in_1[6]), .E(n980), .CK(clk), .Q(R13[6]) );
  EDFFX1 R13_reg_5_ ( .D(data_in_1[5]), .E(n980), .CK(clk), .Q(R13[5]) );
  EDFFX1 R13_reg_4_ ( .D(data_in_1[4]), .E(n980), .CK(clk), .Q(R13[4]) );
  EDFFX1 R13_reg_3_ ( .D(data_in_1[3]), .E(n980), .CK(clk), .Q(R13[3]) );
  EDFFX1 R13_reg_2_ ( .D(data_in_1[2]), .E(n980), .CK(clk), .Q(R13[2]) );
  EDFFX1 R13_reg_1_ ( .D(data_in_1[1]), .E(n980), .CK(clk), .Q(R13[1]) );
  EDFFX1 R13_reg_0_ ( .D(data_in_1[0]), .E(n980), .CK(clk), .Q(R13[0]) );
  EDFFX1 R1_reg_33_ ( .D(data_in_1[33]), .E(n13), .CK(clk), .Q(R1[33]) );
  EDFFX1 R1_reg_32_ ( .D(data_in_1[32]), .E(n13), .CK(clk), .Q(R1[32]) );
  EDFFX1 R1_reg_31_ ( .D(data_in_1[31]), .E(n13), .CK(clk), .Q(R1[31]) );
  EDFFX1 R1_reg_30_ ( .D(data_in_1[30]), .E(n13), .CK(clk), .Q(R1[30]) );
  EDFFX1 R1_reg_29_ ( .D(data_in_1[29]), .E(n13), .CK(clk), .Q(R1[29]) );
  EDFFX1 R1_reg_28_ ( .D(data_in_1[28]), .E(n13), .CK(clk), .Q(R1[28]) );
  EDFFX1 R1_reg_27_ ( .D(data_in_1[27]), .E(n13), .CK(clk), .Q(R1[27]) );
  EDFFX1 R1_reg_26_ ( .D(data_in_1[26]), .E(n13), .CK(clk), .Q(R1[26]) );
  EDFFX1 R1_reg_25_ ( .D(data_in_1[25]), .E(n13), .CK(clk), .Q(R1[25]) );
  EDFFX1 R1_reg_24_ ( .D(data_in_1[24]), .E(n13), .CK(clk), .Q(R1[24]) );
  EDFFX1 R1_reg_23_ ( .D(data_in_1[23]), .E(n13), .CK(clk), .Q(R1[23]) );
  EDFFX1 R1_reg_22_ ( .D(data_in_1[22]), .E(n13), .CK(clk), .Q(R1[22]) );
  EDFFX1 R1_reg_21_ ( .D(data_in_1[21]), .E(n13), .CK(clk), .Q(R1[21]) );
  EDFFX1 R1_reg_20_ ( .D(data_in_1[20]), .E(n13), .CK(clk), .Q(R1[20]) );
  EDFFX1 R1_reg_19_ ( .D(data_in_1[19]), .E(n13), .CK(clk), .Q(R1[19]) );
  EDFFX1 R1_reg_18_ ( .D(data_in_1[18]), .E(n13), .CK(clk), .Q(R1[18]) );
  EDFFX1 R1_reg_17_ ( .D(data_in_1[17]), .E(n13), .CK(clk), .Q(R1[17]) );
  EDFFX1 R1_reg_16_ ( .D(data_in_1[16]), .E(n13), .CK(clk), .Q(R1[16]) );
  EDFFX1 R1_reg_15_ ( .D(data_in_1[15]), .E(n13), .CK(clk), .Q(R1[15]) );
  EDFFX1 R1_reg_14_ ( .D(data_in_1[14]), .E(n13), .CK(clk), .Q(R1[14]) );
  EDFFX1 R1_reg_13_ ( .D(data_in_1[13]), .E(n13), .CK(clk), .Q(R1[13]) );
  EDFFX1 R1_reg_12_ ( .D(data_in_1[12]), .E(n13), .CK(clk), .Q(R1[12]) );
  EDFFX1 R1_reg_11_ ( .D(data_in_1[11]), .E(n13), .CK(clk), .Q(R1[11]) );
  EDFFX1 R1_reg_10_ ( .D(data_in_1[10]), .E(n13), .CK(clk), .Q(R1[10]) );
  EDFFX1 R1_reg_9_ ( .D(data_in_1[9]), .E(n13), .CK(clk), .Q(R1[9]) );
  EDFFX1 R1_reg_8_ ( .D(data_in_1[8]), .E(n13), .CK(clk), .Q(R1[8]) );
  EDFFX1 R1_reg_7_ ( .D(data_in_1[7]), .E(n13), .CK(clk), .Q(R1[7]) );
  EDFFX1 R1_reg_6_ ( .D(data_in_1[6]), .E(n13), .CK(clk), .Q(R1[6]) );
  EDFFX1 R1_reg_5_ ( .D(data_in_1[5]), .E(n13), .CK(clk), .Q(R1[5]) );
  EDFFX1 R1_reg_4_ ( .D(data_in_1[4]), .E(n13), .CK(clk), .Q(R1[4]) );
  EDFFX1 R1_reg_3_ ( .D(data_in_1[3]), .E(n13), .CK(clk), .Q(R1[3]) );
  EDFFX1 R1_reg_2_ ( .D(data_in_1[2]), .E(n13), .CK(clk), .Q(R1[2]) );
  EDFFX1 R1_reg_1_ ( .D(data_in_1[1]), .E(n13), .CK(clk), .Q(R1[1]) );
  EDFFX1 R1_reg_0_ ( .D(data_in_1[0]), .E(n13), .CK(clk), .Q(R1[0]) );
  EDFFX1 R5_reg_33_ ( .D(data_in_1[33]), .E(n12), .CK(clk), .Q(R5[33]) );
  EDFFX1 R5_reg_32_ ( .D(data_in_1[32]), .E(n12), .CK(clk), .Q(R5[32]) );
  EDFFX1 R5_reg_31_ ( .D(data_in_1[31]), .E(n12), .CK(clk), .Q(R5[31]) );
  EDFFX1 R5_reg_30_ ( .D(data_in_1[30]), .E(n12), .CK(clk), .Q(R5[30]) );
  EDFFX1 R5_reg_29_ ( .D(data_in_1[29]), .E(n12), .CK(clk), .Q(R5[29]) );
  EDFFX1 R5_reg_28_ ( .D(data_in_1[28]), .E(n12), .CK(clk), .Q(R5[28]) );
  EDFFX1 R5_reg_27_ ( .D(data_in_1[27]), .E(n12), .CK(clk), .Q(R5[27]) );
  EDFFX1 R5_reg_26_ ( .D(data_in_1[26]), .E(n12), .CK(clk), .Q(R5[26]) );
  EDFFX1 R5_reg_25_ ( .D(data_in_1[25]), .E(n12), .CK(clk), .Q(R5[25]) );
  EDFFX1 R5_reg_24_ ( .D(data_in_1[24]), .E(n12), .CK(clk), .Q(R5[24]) );
  EDFFX1 R5_reg_23_ ( .D(data_in_1[23]), .E(n12), .CK(clk), .Q(R5[23]) );
  EDFFX1 R5_reg_22_ ( .D(data_in_1[22]), .E(n12), .CK(clk), .Q(R5[22]) );
  EDFFX1 R5_reg_21_ ( .D(data_in_1[21]), .E(n12), .CK(clk), .Q(R5[21]) );
  EDFFX1 R5_reg_20_ ( .D(data_in_1[20]), .E(n12), .CK(clk), .Q(R5[20]) );
  EDFFX1 R5_reg_19_ ( .D(data_in_1[19]), .E(n12), .CK(clk), .Q(R5[19]) );
  EDFFX1 R5_reg_18_ ( .D(data_in_1[18]), .E(n12), .CK(clk), .Q(R5[18]) );
  EDFFX1 R5_reg_17_ ( .D(data_in_1[17]), .E(n12), .CK(clk), .Q(R5[17]) );
  EDFFX1 R5_reg_16_ ( .D(data_in_1[16]), .E(n12), .CK(clk), .Q(R5[16]) );
  EDFFX1 R5_reg_15_ ( .D(data_in_1[15]), .E(n12), .CK(clk), .Q(R5[15]) );
  EDFFX1 R5_reg_14_ ( .D(data_in_1[14]), .E(n12), .CK(clk), .Q(R5[14]) );
  EDFFX1 R5_reg_13_ ( .D(data_in_1[13]), .E(n12), .CK(clk), .Q(R5[13]) );
  EDFFX1 R5_reg_12_ ( .D(data_in_1[12]), .E(n12), .CK(clk), .Q(R5[12]) );
  EDFFX1 R5_reg_11_ ( .D(data_in_1[11]), .E(n12), .CK(clk), .Q(R5[11]) );
  EDFFX1 R5_reg_10_ ( .D(data_in_1[10]), .E(n12), .CK(clk), .Q(R5[10]) );
  EDFFX1 R5_reg_9_ ( .D(data_in_1[9]), .E(n12), .CK(clk), .Q(R5[9]) );
  EDFFX1 R5_reg_8_ ( .D(data_in_1[8]), .E(n12), .CK(clk), .Q(R5[8]) );
  EDFFX1 R5_reg_7_ ( .D(data_in_1[7]), .E(n12), .CK(clk), .Q(R5[7]) );
  EDFFX1 R5_reg_6_ ( .D(data_in_1[6]), .E(n12), .CK(clk), .Q(R5[6]) );
  EDFFX1 R5_reg_5_ ( .D(data_in_1[5]), .E(n12), .CK(clk), .Q(R5[5]) );
  EDFFX1 R5_reg_4_ ( .D(data_in_1[4]), .E(n12), .CK(clk), .Q(R5[4]) );
  EDFFX1 R5_reg_3_ ( .D(data_in_1[3]), .E(n12), .CK(clk), .Q(R5[3]) );
  EDFFX1 R5_reg_2_ ( .D(data_in_1[2]), .E(n12), .CK(clk), .Q(R5[2]) );
  EDFFX1 R5_reg_1_ ( .D(data_in_1[1]), .E(n12), .CK(clk), .Q(R5[1]) );
  EDFFX1 R5_reg_0_ ( .D(data_in_1[0]), .E(n12), .CK(clk), .Q(R5[0]) );
  EDFFX1 R9_reg_33_ ( .D(data_in_1[33]), .E(n11), .CK(clk), .Q(R9[33]) );
  EDFFX1 R9_reg_32_ ( .D(data_in_1[32]), .E(n11), .CK(clk), .Q(R9[32]) );
  EDFFX1 R9_reg_31_ ( .D(data_in_1[31]), .E(n11), .CK(clk), .Q(R9[31]) );
  EDFFX1 R9_reg_30_ ( .D(data_in_1[30]), .E(n11), .CK(clk), .Q(R9[30]) );
  EDFFX1 R9_reg_29_ ( .D(data_in_1[29]), .E(n11), .CK(clk), .Q(R9[29]) );
  EDFFX1 R9_reg_28_ ( .D(data_in_1[28]), .E(n11), .CK(clk), .Q(R9[28]) );
  EDFFX1 R9_reg_27_ ( .D(data_in_1[27]), .E(n11), .CK(clk), .Q(R9[27]) );
  EDFFX1 R9_reg_26_ ( .D(data_in_1[26]), .E(n11), .CK(clk), .Q(R9[26]) );
  EDFFX1 R9_reg_25_ ( .D(data_in_1[25]), .E(n11), .CK(clk), .Q(R9[25]) );
  EDFFX1 R9_reg_24_ ( .D(data_in_1[24]), .E(n11), .CK(clk), .Q(R9[24]) );
  EDFFX1 R9_reg_23_ ( .D(data_in_1[23]), .E(n11), .CK(clk), .Q(R9[23]) );
  EDFFX1 R9_reg_22_ ( .D(data_in_1[22]), .E(n11), .CK(clk), .Q(R9[22]) );
  EDFFX1 R9_reg_21_ ( .D(data_in_1[21]), .E(n11), .CK(clk), .Q(R9[21]) );
  EDFFX1 R9_reg_20_ ( .D(data_in_1[20]), .E(n11), .CK(clk), .Q(R9[20]) );
  EDFFX1 R9_reg_19_ ( .D(data_in_1[19]), .E(n11), .CK(clk), .Q(R9[19]) );
  EDFFX1 R9_reg_18_ ( .D(data_in_1[18]), .E(n11), .CK(clk), .Q(R9[18]) );
  EDFFX1 R9_reg_17_ ( .D(data_in_1[17]), .E(n11), .CK(clk), .Q(R9[17]) );
  EDFFX1 R9_reg_16_ ( .D(data_in_1[16]), .E(n11), .CK(clk), .Q(R9[16]) );
  EDFFX1 R9_reg_15_ ( .D(data_in_1[15]), .E(n11), .CK(clk), .Q(R9[15]) );
  EDFFX1 R9_reg_14_ ( .D(data_in_1[14]), .E(n11), .CK(clk), .Q(R9[14]) );
  EDFFX1 R9_reg_13_ ( .D(data_in_1[13]), .E(n11), .CK(clk), .Q(R9[13]) );
  EDFFX1 R9_reg_12_ ( .D(data_in_1[12]), .E(n11), .CK(clk), .Q(R9[12]) );
  EDFFX1 R9_reg_11_ ( .D(data_in_1[11]), .E(n11), .CK(clk), .Q(R9[11]) );
  EDFFX1 R9_reg_10_ ( .D(data_in_1[10]), .E(n11), .CK(clk), .Q(R9[10]) );
  EDFFX1 R9_reg_9_ ( .D(data_in_1[9]), .E(n11), .CK(clk), .Q(R9[9]) );
  EDFFX1 R9_reg_8_ ( .D(data_in_1[8]), .E(n11), .CK(clk), .Q(R9[8]) );
  EDFFX1 R9_reg_7_ ( .D(data_in_1[7]), .E(n11), .CK(clk), .Q(R9[7]) );
  EDFFX1 R9_reg_6_ ( .D(data_in_1[6]), .E(n11), .CK(clk), .Q(R9[6]) );
  EDFFX1 R9_reg_5_ ( .D(data_in_1[5]), .E(n11), .CK(clk), .Q(R9[5]) );
  EDFFX1 R9_reg_4_ ( .D(data_in_1[4]), .E(n11), .CK(clk), .Q(R9[4]) );
  EDFFX1 R9_reg_3_ ( .D(data_in_1[3]), .E(n11), .CK(clk), .Q(R9[3]) );
  EDFFX1 R9_reg_2_ ( .D(data_in_1[2]), .E(n11), .CK(clk), .Q(R9[2]) );
  EDFFX1 R9_reg_1_ ( .D(data_in_1[1]), .E(n11), .CK(clk), .Q(R9[1]) );
  EDFFX1 R9_reg_0_ ( .D(data_in_1[0]), .E(n11), .CK(clk), .Q(R9[0]) );
  EDFFX1 R14_reg_33_ ( .D(data_in_1[33]), .E(n982), .CK(clk), .Q(R14[33]) );
  EDFFX1 R14_reg_32_ ( .D(data_in_1[32]), .E(n982), .CK(clk), .Q(R14[32]) );
  EDFFX1 R14_reg_31_ ( .D(data_in_1[31]), .E(n982), .CK(clk), .Q(R14[31]) );
  EDFFX1 R14_reg_30_ ( .D(data_in_1[30]), .E(n982), .CK(clk), .Q(R14[30]) );
  EDFFX1 R14_reg_29_ ( .D(data_in_1[29]), .E(n982), .CK(clk), .Q(R14[29]) );
  EDFFX1 R14_reg_28_ ( .D(data_in_1[28]), .E(n982), .CK(clk), .Q(R14[28]) );
  EDFFX1 R14_reg_27_ ( .D(data_in_1[27]), .E(n982), .CK(clk), .Q(R14[27]) );
  EDFFX1 R14_reg_26_ ( .D(data_in_1[26]), .E(n982), .CK(clk), .Q(R14[26]) );
  EDFFX1 R14_reg_25_ ( .D(data_in_1[25]), .E(n982), .CK(clk), .Q(R14[25]) );
  EDFFX1 R14_reg_24_ ( .D(data_in_1[24]), .E(n982), .CK(clk), .Q(R14[24]) );
  EDFFX1 R14_reg_23_ ( .D(data_in_1[23]), .E(n982), .CK(clk), .Q(R14[23]) );
  EDFFX1 R14_reg_22_ ( .D(data_in_1[22]), .E(n982), .CK(clk), .Q(R14[22]) );
  EDFFX1 R14_reg_21_ ( .D(data_in_1[21]), .E(n982), .CK(clk), .Q(R14[21]) );
  EDFFX1 R14_reg_20_ ( .D(data_in_1[20]), .E(n982), .CK(clk), .Q(R14[20]) );
  EDFFX1 R14_reg_19_ ( .D(data_in_1[19]), .E(n982), .CK(clk), .Q(R14[19]) );
  EDFFX1 R14_reg_18_ ( .D(data_in_1[18]), .E(n982), .CK(clk), .Q(R14[18]) );
  EDFFX1 R14_reg_17_ ( .D(data_in_1[17]), .E(n982), .CK(clk), .Q(R14[17]) );
  EDFFX1 R14_reg_16_ ( .D(data_in_1[16]), .E(n982), .CK(clk), .Q(R14[16]) );
  EDFFX1 R14_reg_15_ ( .D(data_in_1[15]), .E(n982), .CK(clk), .Q(R14[15]) );
  EDFFX1 R14_reg_14_ ( .D(data_in_1[14]), .E(n982), .CK(clk), .Q(R14[14]) );
  EDFFX1 R14_reg_13_ ( .D(data_in_1[13]), .E(n982), .CK(clk), .Q(R14[13]) );
  EDFFX1 R14_reg_12_ ( .D(data_in_1[12]), .E(n982), .CK(clk), .Q(R14[12]) );
  EDFFX1 R14_reg_11_ ( .D(data_in_1[11]), .E(n982), .CK(clk), .Q(R14[11]) );
  EDFFX1 R14_reg_10_ ( .D(data_in_1[10]), .E(n982), .CK(clk), .Q(R14[10]) );
  EDFFX1 R14_reg_9_ ( .D(data_in_1[9]), .E(n982), .CK(clk), .Q(R14[9]) );
  EDFFX1 R14_reg_8_ ( .D(data_in_1[8]), .E(n982), .CK(clk), .Q(R14[8]) );
  EDFFX1 R14_reg_7_ ( .D(data_in_1[7]), .E(n982), .CK(clk), .Q(R14[7]) );
  EDFFX1 R14_reg_6_ ( .D(data_in_1[6]), .E(n982), .CK(clk), .Q(R14[6]) );
  EDFFX1 R14_reg_5_ ( .D(data_in_1[5]), .E(n982), .CK(clk), .Q(R14[5]) );
  EDFFX1 R14_reg_4_ ( .D(data_in_1[4]), .E(n982), .CK(clk), .Q(R14[4]) );
  EDFFX1 R14_reg_3_ ( .D(data_in_1[3]), .E(n982), .CK(clk), .Q(R14[3]) );
  EDFFX1 R14_reg_2_ ( .D(data_in_1[2]), .E(n982), .CK(clk), .Q(R14[2]) );
  EDFFX1 R14_reg_1_ ( .D(data_in_1[1]), .E(n982), .CK(clk), .Q(R14[1]) );
  EDFFX1 R14_reg_0_ ( .D(data_in_1[0]), .E(n982), .CK(clk), .Q(R14[0]) );
  EDFFX1 R2_reg_33_ ( .D(data_in_1[33]), .E(n10), .CK(clk), .Q(R2[33]) );
  EDFFX1 R2_reg_32_ ( .D(data_in_1[32]), .E(n10), .CK(clk), .Q(R2[32]) );
  EDFFX1 R2_reg_31_ ( .D(data_in_1[31]), .E(n10), .CK(clk), .Q(R2[31]) );
  EDFFX1 R2_reg_30_ ( .D(data_in_1[30]), .E(n10), .CK(clk), .Q(R2[30]) );
  EDFFX1 R2_reg_29_ ( .D(data_in_1[29]), .E(n10), .CK(clk), .Q(R2[29]) );
  EDFFX1 R2_reg_28_ ( .D(data_in_1[28]), .E(n10), .CK(clk), .Q(R2[28]) );
  EDFFX1 R2_reg_27_ ( .D(data_in_1[27]), .E(n10), .CK(clk), .Q(R2[27]) );
  EDFFX1 R2_reg_26_ ( .D(data_in_1[26]), .E(n10), .CK(clk), .Q(R2[26]) );
  EDFFX1 R2_reg_25_ ( .D(data_in_1[25]), .E(n10), .CK(clk), .Q(R2[25]) );
  EDFFX1 R2_reg_24_ ( .D(data_in_1[24]), .E(n10), .CK(clk), .Q(R2[24]) );
  EDFFX1 R2_reg_23_ ( .D(data_in_1[23]), .E(n10), .CK(clk), .Q(R2[23]) );
  EDFFX1 R2_reg_22_ ( .D(data_in_1[22]), .E(n10), .CK(clk), .Q(R2[22]) );
  EDFFX1 R2_reg_21_ ( .D(data_in_1[21]), .E(n10), .CK(clk), .Q(R2[21]) );
  EDFFX1 R2_reg_20_ ( .D(data_in_1[20]), .E(n10), .CK(clk), .Q(R2[20]) );
  EDFFX1 R2_reg_19_ ( .D(data_in_1[19]), .E(n10), .CK(clk), .Q(R2[19]) );
  EDFFX1 R2_reg_18_ ( .D(data_in_1[18]), .E(n10), .CK(clk), .Q(R2[18]) );
  EDFFX1 R2_reg_17_ ( .D(data_in_1[17]), .E(n10), .CK(clk), .Q(R2[17]) );
  EDFFX1 R2_reg_16_ ( .D(data_in_1[16]), .E(n10), .CK(clk), .Q(R2[16]) );
  EDFFX1 R2_reg_15_ ( .D(data_in_1[15]), .E(n10), .CK(clk), .Q(R2[15]) );
  EDFFX1 R2_reg_14_ ( .D(data_in_1[14]), .E(n10), .CK(clk), .Q(R2[14]) );
  EDFFX1 R2_reg_13_ ( .D(data_in_1[13]), .E(n10), .CK(clk), .Q(R2[13]) );
  EDFFX1 R2_reg_12_ ( .D(data_in_1[12]), .E(n10), .CK(clk), .Q(R2[12]) );
  EDFFX1 R2_reg_11_ ( .D(data_in_1[11]), .E(n10), .CK(clk), .Q(R2[11]) );
  EDFFX1 R2_reg_10_ ( .D(data_in_1[10]), .E(n10), .CK(clk), .Q(R2[10]) );
  EDFFX1 R2_reg_9_ ( .D(data_in_1[9]), .E(n10), .CK(clk), .Q(R2[9]) );
  EDFFX1 R2_reg_8_ ( .D(data_in_1[8]), .E(n10), .CK(clk), .Q(R2[8]) );
  EDFFX1 R2_reg_7_ ( .D(data_in_1[7]), .E(n10), .CK(clk), .Q(R2[7]) );
  EDFFX1 R2_reg_6_ ( .D(data_in_1[6]), .E(n10), .CK(clk), .Q(R2[6]) );
  EDFFX1 R2_reg_5_ ( .D(data_in_1[5]), .E(n10), .CK(clk), .Q(R2[5]) );
  EDFFX1 R2_reg_4_ ( .D(data_in_1[4]), .E(n10), .CK(clk), .Q(R2[4]) );
  EDFFX1 R2_reg_3_ ( .D(data_in_1[3]), .E(n10), .CK(clk), .Q(R2[3]) );
  EDFFX1 R2_reg_2_ ( .D(data_in_1[2]), .E(n10), .CK(clk), .Q(R2[2]) );
  EDFFX1 R2_reg_1_ ( .D(data_in_1[1]), .E(n10), .CK(clk), .Q(R2[1]) );
  EDFFX1 R2_reg_0_ ( .D(data_in_1[0]), .E(n10), .CK(clk), .Q(R2[0]) );
  EDFFX1 R6_reg_33_ ( .D(data_in_1[33]), .E(n9), .CK(clk), .Q(R6[33]) );
  EDFFX1 R6_reg_32_ ( .D(data_in_1[32]), .E(n9), .CK(clk), .Q(R6[32]) );
  EDFFX1 R6_reg_31_ ( .D(data_in_1[31]), .E(n9), .CK(clk), .Q(R6[31]) );
  EDFFX1 R6_reg_30_ ( .D(data_in_1[30]), .E(n9), .CK(clk), .Q(R6[30]) );
  EDFFX1 R6_reg_29_ ( .D(data_in_1[29]), .E(n9), .CK(clk), .Q(R6[29]) );
  EDFFX1 R6_reg_28_ ( .D(data_in_1[28]), .E(n9), .CK(clk), .Q(R6[28]) );
  EDFFX1 R6_reg_27_ ( .D(data_in_1[27]), .E(n9), .CK(clk), .Q(R6[27]) );
  EDFFX1 R6_reg_26_ ( .D(data_in_1[26]), .E(n9), .CK(clk), .Q(R6[26]) );
  EDFFX1 R6_reg_25_ ( .D(data_in_1[25]), .E(n9), .CK(clk), .Q(R6[25]) );
  EDFFX1 R6_reg_24_ ( .D(data_in_1[24]), .E(n9), .CK(clk), .Q(R6[24]) );
  EDFFX1 R6_reg_23_ ( .D(data_in_1[23]), .E(n9), .CK(clk), .Q(R6[23]) );
  EDFFX1 R6_reg_22_ ( .D(data_in_1[22]), .E(n9), .CK(clk), .Q(R6[22]) );
  EDFFX1 R6_reg_21_ ( .D(data_in_1[21]), .E(n9), .CK(clk), .Q(R6[21]) );
  EDFFX1 R6_reg_20_ ( .D(data_in_1[20]), .E(n9), .CK(clk), .Q(R6[20]) );
  EDFFX1 R6_reg_19_ ( .D(data_in_1[19]), .E(n9), .CK(clk), .Q(R6[19]) );
  EDFFX1 R6_reg_18_ ( .D(data_in_1[18]), .E(n9), .CK(clk), .Q(R6[18]) );
  EDFFX1 R6_reg_17_ ( .D(data_in_1[17]), .E(n9), .CK(clk), .Q(R6[17]) );
  EDFFX1 R6_reg_16_ ( .D(data_in_1[16]), .E(n9), .CK(clk), .Q(R6[16]) );
  EDFFX1 R6_reg_15_ ( .D(data_in_1[15]), .E(n9), .CK(clk), .Q(R6[15]) );
  EDFFX1 R6_reg_14_ ( .D(data_in_1[14]), .E(n9), .CK(clk), .Q(R6[14]) );
  EDFFX1 R6_reg_13_ ( .D(data_in_1[13]), .E(n9), .CK(clk), .Q(R6[13]) );
  EDFFX1 R6_reg_12_ ( .D(data_in_1[12]), .E(n9), .CK(clk), .Q(R6[12]) );
  EDFFX1 R6_reg_11_ ( .D(data_in_1[11]), .E(n9), .CK(clk), .Q(R6[11]) );
  EDFFX1 R6_reg_10_ ( .D(data_in_1[10]), .E(n9), .CK(clk), .Q(R6[10]) );
  EDFFX1 R6_reg_9_ ( .D(data_in_1[9]), .E(n9), .CK(clk), .Q(R6[9]) );
  EDFFX1 R6_reg_8_ ( .D(data_in_1[8]), .E(n9), .CK(clk), .Q(R6[8]) );
  EDFFX1 R6_reg_7_ ( .D(data_in_1[7]), .E(n9), .CK(clk), .Q(R6[7]) );
  EDFFX1 R6_reg_6_ ( .D(data_in_1[6]), .E(n9), .CK(clk), .Q(R6[6]) );
  EDFFX1 R6_reg_5_ ( .D(data_in_1[5]), .E(n9), .CK(clk), .Q(R6[5]) );
  EDFFX1 R6_reg_4_ ( .D(data_in_1[4]), .E(n9), .CK(clk), .Q(R6[4]) );
  EDFFX1 R6_reg_3_ ( .D(data_in_1[3]), .E(n9), .CK(clk), .Q(R6[3]) );
  EDFFX1 R6_reg_2_ ( .D(data_in_1[2]), .E(n9), .CK(clk), .Q(R6[2]) );
  EDFFX1 R6_reg_1_ ( .D(data_in_1[1]), .E(n9), .CK(clk), .Q(R6[1]) );
  EDFFX1 R6_reg_0_ ( .D(data_in_1[0]), .E(n9), .CK(clk), .Q(R6[0]) );
  EDFFX1 R10_reg_33_ ( .D(data_in_1[33]), .E(n8), .CK(clk), .Q(R10[33]) );
  EDFFX1 R10_reg_32_ ( .D(data_in_1[32]), .E(n8), .CK(clk), .Q(R10[32]) );
  EDFFX1 R10_reg_31_ ( .D(data_in_1[31]), .E(n8), .CK(clk), .Q(R10[31]) );
  EDFFX1 R10_reg_30_ ( .D(data_in_1[30]), .E(n8), .CK(clk), .Q(R10[30]) );
  EDFFX1 R10_reg_29_ ( .D(data_in_1[29]), .E(n8), .CK(clk), .Q(R10[29]) );
  EDFFX1 R10_reg_28_ ( .D(data_in_1[28]), .E(n8), .CK(clk), .Q(R10[28]) );
  EDFFX1 R10_reg_27_ ( .D(data_in_1[27]), .E(n8), .CK(clk), .Q(R10[27]) );
  EDFFX1 R10_reg_26_ ( .D(data_in_1[26]), .E(n8), .CK(clk), .Q(R10[26]) );
  EDFFX1 R10_reg_25_ ( .D(data_in_1[25]), .E(n8), .CK(clk), .Q(R10[25]) );
  EDFFX1 R10_reg_24_ ( .D(data_in_1[24]), .E(n8), .CK(clk), .Q(R10[24]) );
  EDFFX1 R10_reg_23_ ( .D(data_in_1[23]), .E(n8), .CK(clk), .Q(R10[23]) );
  EDFFX1 R10_reg_22_ ( .D(data_in_1[22]), .E(n8), .CK(clk), .Q(R10[22]) );
  EDFFX1 R10_reg_21_ ( .D(data_in_1[21]), .E(n8), .CK(clk), .Q(R10[21]) );
  EDFFX1 R10_reg_20_ ( .D(data_in_1[20]), .E(n8), .CK(clk), .Q(R10[20]) );
  EDFFX1 R10_reg_19_ ( .D(data_in_1[19]), .E(n8), .CK(clk), .Q(R10[19]) );
  EDFFX1 R10_reg_18_ ( .D(data_in_1[18]), .E(n8), .CK(clk), .Q(R10[18]) );
  EDFFX1 R10_reg_17_ ( .D(data_in_1[17]), .E(n8), .CK(clk), .Q(R10[17]) );
  EDFFX1 R10_reg_16_ ( .D(data_in_1[16]), .E(n8), .CK(clk), .Q(R10[16]) );
  EDFFX1 R10_reg_15_ ( .D(data_in_1[15]), .E(n8), .CK(clk), .Q(R10[15]) );
  EDFFX1 R10_reg_14_ ( .D(data_in_1[14]), .E(n8), .CK(clk), .Q(R10[14]) );
  EDFFX1 R10_reg_13_ ( .D(data_in_1[13]), .E(n8), .CK(clk), .Q(R10[13]) );
  EDFFX1 R10_reg_12_ ( .D(data_in_1[12]), .E(n8), .CK(clk), .Q(R10[12]) );
  EDFFX1 R10_reg_11_ ( .D(data_in_1[11]), .E(n8), .CK(clk), .Q(R10[11]) );
  EDFFX1 R10_reg_10_ ( .D(data_in_1[10]), .E(n8), .CK(clk), .Q(R10[10]) );
  EDFFX1 R10_reg_9_ ( .D(data_in_1[9]), .E(n8), .CK(clk), .Q(R10[9]) );
  EDFFX1 R10_reg_8_ ( .D(data_in_1[8]), .E(n8), .CK(clk), .Q(R10[8]) );
  EDFFX1 R10_reg_7_ ( .D(data_in_1[7]), .E(n8), .CK(clk), .Q(R10[7]) );
  EDFFX1 R10_reg_6_ ( .D(data_in_1[6]), .E(n8), .CK(clk), .Q(R10[6]) );
  EDFFX1 R10_reg_5_ ( .D(data_in_1[5]), .E(n8), .CK(clk), .Q(R10[5]) );
  EDFFX1 R10_reg_4_ ( .D(data_in_1[4]), .E(n8), .CK(clk), .Q(R10[4]) );
  EDFFX1 R10_reg_3_ ( .D(data_in_1[3]), .E(n8), .CK(clk), .Q(R10[3]) );
  EDFFX1 R10_reg_2_ ( .D(data_in_1[2]), .E(n8), .CK(clk), .Q(R10[2]) );
  EDFFX1 R10_reg_1_ ( .D(data_in_1[1]), .E(n8), .CK(clk), .Q(R10[1]) );
  EDFFX1 R10_reg_0_ ( .D(data_in_1[0]), .E(n8), .CK(clk), .Q(R10[0]) );
  EDFFX1 R0_reg_33_ ( .D(data_in_1[33]), .E(n1002), .CK(clk), .Q(R0[33]) );
  EDFFX1 R0_reg_32_ ( .D(data_in_1[32]), .E(n1002), .CK(clk), .Q(R0[32]) );
  EDFFX1 R0_reg_31_ ( .D(data_in_1[31]), .E(n1002), .CK(clk), .Q(R0[31]) );
  EDFFX1 R0_reg_30_ ( .D(data_in_1[30]), .E(n1002), .CK(clk), .Q(R0[30]) );
  EDFFX1 R0_reg_29_ ( .D(data_in_1[29]), .E(n1002), .CK(clk), .Q(R0[29]) );
  EDFFX1 R0_reg_28_ ( .D(data_in_1[28]), .E(n1002), .CK(clk), .Q(R0[28]) );
  EDFFX1 R0_reg_27_ ( .D(data_in_1[27]), .E(n1002), .CK(clk), .Q(R0[27]) );
  EDFFX1 R0_reg_26_ ( .D(data_in_1[26]), .E(n1002), .CK(clk), .Q(R0[26]) );
  EDFFX1 R0_reg_25_ ( .D(data_in_1[25]), .E(n1002), .CK(clk), .Q(R0[25]) );
  EDFFX1 R0_reg_24_ ( .D(data_in_1[24]), .E(n1002), .CK(clk), .Q(R0[24]) );
  EDFFX1 R0_reg_23_ ( .D(data_in_1[23]), .E(n1002), .CK(clk), .Q(R0[23]) );
  EDFFX1 R0_reg_22_ ( .D(data_in_1[22]), .E(n1002), .CK(clk), .Q(R0[22]) );
  EDFFX1 R0_reg_21_ ( .D(data_in_1[21]), .E(n1002), .CK(clk), .Q(R0[21]) );
  EDFFX1 R0_reg_20_ ( .D(data_in_1[20]), .E(n1002), .CK(clk), .Q(R0[20]) );
  EDFFX1 R0_reg_19_ ( .D(data_in_1[19]), .E(n1002), .CK(clk), .Q(R0[19]) );
  EDFFX1 R0_reg_18_ ( .D(data_in_1[18]), .E(n1002), .CK(clk), .Q(R0[18]) );
  EDFFX1 R0_reg_17_ ( .D(data_in_1[17]), .E(n1002), .CK(clk), .Q(R0[17]) );
  EDFFX1 R0_reg_16_ ( .D(data_in_1[16]), .E(n1002), .CK(clk), .Q(R0[16]) );
  EDFFX1 R0_reg_15_ ( .D(data_in_1[15]), .E(n1001), .CK(clk), .Q(R0[15]) );
  EDFFX1 R0_reg_14_ ( .D(data_in_1[14]), .E(n996), .CK(clk), .Q(R0[14]) );
  EDFFX1 R0_reg_13_ ( .D(data_in_1[13]), .E(n998), .CK(clk), .Q(R0[13]) );
  EDFFX1 R0_reg_12_ ( .D(data_in_1[12]), .E(n999), .CK(clk), .Q(R0[12]) );
  EDFFX1 R0_reg_11_ ( .D(data_in_1[11]), .E(n1000), .CK(clk), .Q(R0[11]) );
  EDFFX1 R0_reg_10_ ( .D(data_in_1[10]), .E(n1001), .CK(clk), .Q(R0[10]) );
  EDFFX1 R0_reg_9_ ( .D(data_in_1[9]), .E(n998), .CK(clk), .Q(R0[9]) );
  EDFFX1 R0_reg_8_ ( .D(data_in_1[8]), .E(n999), .CK(clk), .Q(R0[8]) );
  EDFFX1 R0_reg_7_ ( .D(data_in_1[7]), .E(n1000), .CK(clk), .Q(R0[7]) );
  EDFFX1 R0_reg_6_ ( .D(data_in_1[6]), .E(n1001), .CK(clk), .Q(R0[6]) );
  EDFFX1 R0_reg_5_ ( .D(data_in_1[5]), .E(n998), .CK(clk), .Q(R0[5]) );
  EDFFX1 R0_reg_4_ ( .D(data_in_1[4]), .E(n999), .CK(clk), .Q(R0[4]) );
  EDFFX1 R0_reg_3_ ( .D(data_in_1[3]), .E(n1000), .CK(clk), .Q(R0[3]) );
  EDFFX1 R0_reg_2_ ( .D(data_in_1[2]), .E(n1001), .CK(clk), .Q(R0[2]) );
  EDFFX1 R0_reg_1_ ( .D(data_in_1[1]), .E(n998), .CK(clk), .Q(R0[1]) );
  EDFFX1 R0_reg_0_ ( .D(data_in_1[0]), .E(n999), .CK(clk), .Q(R0[0]) );
  EDFFX1 R4_reg_33_ ( .D(data_in_1[33]), .E(n7), .CK(clk), .Q(R4[33]) );
  EDFFX1 R4_reg_32_ ( .D(data_in_1[32]), .E(n7), .CK(clk), .Q(R4[32]) );
  EDFFX1 R4_reg_31_ ( .D(data_in_1[31]), .E(n7), .CK(clk), .Q(R4[31]) );
  EDFFX1 R4_reg_30_ ( .D(data_in_1[30]), .E(n7), .CK(clk), .Q(R4[30]) );
  EDFFX1 R4_reg_29_ ( .D(data_in_1[29]), .E(n7), .CK(clk), .Q(R4[29]) );
  EDFFX1 R4_reg_28_ ( .D(data_in_1[28]), .E(n7), .CK(clk), .Q(R4[28]) );
  EDFFX1 R4_reg_27_ ( .D(data_in_1[27]), .E(n7), .CK(clk), .Q(R4[27]) );
  EDFFX1 R4_reg_26_ ( .D(data_in_1[26]), .E(n7), .CK(clk), .Q(R4[26]) );
  EDFFX1 R4_reg_25_ ( .D(data_in_1[25]), .E(n7), .CK(clk), .Q(R4[25]) );
  EDFFX1 R4_reg_24_ ( .D(data_in_1[24]), .E(n7), .CK(clk), .Q(R4[24]) );
  EDFFX1 R4_reg_23_ ( .D(data_in_1[23]), .E(n7), .CK(clk), .Q(R4[23]) );
  EDFFX1 R4_reg_22_ ( .D(data_in_1[22]), .E(n7), .CK(clk), .Q(R4[22]) );
  EDFFX1 R4_reg_21_ ( .D(data_in_1[21]), .E(n7), .CK(clk), .Q(R4[21]) );
  EDFFX1 R4_reg_20_ ( .D(data_in_1[20]), .E(n7), .CK(clk), .Q(R4[20]) );
  EDFFX1 R4_reg_19_ ( .D(data_in_1[19]), .E(n7), .CK(clk), .Q(R4[19]) );
  EDFFX1 R4_reg_18_ ( .D(data_in_1[18]), .E(n7), .CK(clk), .Q(R4[18]) );
  EDFFX1 R4_reg_17_ ( .D(data_in_1[17]), .E(n7), .CK(clk), .Q(R4[17]) );
  EDFFX1 R4_reg_16_ ( .D(data_in_1[16]), .E(n7), .CK(clk), .Q(R4[16]) );
  EDFFX1 R4_reg_15_ ( .D(data_in_1[15]), .E(n7), .CK(clk), .Q(R4[15]) );
  EDFFX1 R4_reg_14_ ( .D(data_in_1[14]), .E(n7), .CK(clk), .Q(R4[14]) );
  EDFFX1 R4_reg_13_ ( .D(data_in_1[13]), .E(n7), .CK(clk), .Q(R4[13]) );
  EDFFX1 R4_reg_12_ ( .D(data_in_1[12]), .E(n7), .CK(clk), .Q(R4[12]) );
  EDFFX1 R4_reg_11_ ( .D(data_in_1[11]), .E(n7), .CK(clk), .Q(R4[11]) );
  EDFFX1 R4_reg_10_ ( .D(data_in_1[10]), .E(n7), .CK(clk), .Q(R4[10]) );
  EDFFX1 R4_reg_9_ ( .D(data_in_1[9]), .E(n7), .CK(clk), .Q(R4[9]) );
  EDFFX1 R4_reg_8_ ( .D(data_in_1[8]), .E(n7), .CK(clk), .Q(R4[8]) );
  EDFFX1 R4_reg_7_ ( .D(data_in_1[7]), .E(n7), .CK(clk), .Q(R4[7]) );
  EDFFX1 R4_reg_6_ ( .D(data_in_1[6]), .E(n7), .CK(clk), .Q(R4[6]) );
  EDFFX1 R4_reg_5_ ( .D(data_in_1[5]), .E(n7), .CK(clk), .Q(R4[5]) );
  EDFFX1 R4_reg_4_ ( .D(data_in_1[4]), .E(n7), .CK(clk), .Q(R4[4]) );
  EDFFX1 R4_reg_3_ ( .D(data_in_1[3]), .E(n7), .CK(clk), .Q(R4[3]) );
  EDFFX1 R4_reg_2_ ( .D(data_in_1[2]), .E(n7), .CK(clk), .Q(R4[2]) );
  EDFFX1 R4_reg_1_ ( .D(data_in_1[1]), .E(n7), .CK(clk), .Q(R4[1]) );
  EDFFX1 R4_reg_0_ ( .D(data_in_1[0]), .E(n7), .CK(clk), .Q(R4[0]) );
  EDFFX1 R8_reg_33_ ( .D(data_in_1[33]), .E(n6), .CK(clk), .Q(R8[33]) );
  EDFFX1 R8_reg_32_ ( .D(data_in_1[32]), .E(n6), .CK(clk), .Q(R8[32]) );
  EDFFX1 R8_reg_31_ ( .D(data_in_1[31]), .E(n6), .CK(clk), .Q(R8[31]) );
  EDFFX1 R8_reg_30_ ( .D(data_in_1[30]), .E(n6), .CK(clk), .Q(R8[30]) );
  EDFFX1 R8_reg_29_ ( .D(data_in_1[29]), .E(n6), .CK(clk), .Q(R8[29]) );
  EDFFX1 R8_reg_28_ ( .D(data_in_1[28]), .E(n6), .CK(clk), .Q(R8[28]) );
  EDFFX1 R8_reg_27_ ( .D(data_in_1[27]), .E(n6), .CK(clk), .Q(R8[27]) );
  EDFFX1 R8_reg_26_ ( .D(data_in_1[26]), .E(n6), .CK(clk), .Q(R8[26]) );
  EDFFX1 R8_reg_25_ ( .D(data_in_1[25]), .E(n6), .CK(clk), .Q(R8[25]) );
  EDFFX1 R8_reg_24_ ( .D(data_in_1[24]), .E(n6), .CK(clk), .Q(R8[24]) );
  EDFFX1 R8_reg_23_ ( .D(data_in_1[23]), .E(n6), .CK(clk), .Q(R8[23]) );
  EDFFX1 R8_reg_22_ ( .D(data_in_1[22]), .E(n6), .CK(clk), .Q(R8[22]) );
  EDFFX1 R8_reg_21_ ( .D(data_in_1[21]), .E(n6), .CK(clk), .Q(R8[21]) );
  EDFFX1 R8_reg_20_ ( .D(data_in_1[20]), .E(n6), .CK(clk), .Q(R8[20]) );
  EDFFX1 R8_reg_19_ ( .D(data_in_1[19]), .E(n6), .CK(clk), .Q(R8[19]) );
  EDFFX1 R8_reg_18_ ( .D(data_in_1[18]), .E(n6), .CK(clk), .Q(R8[18]) );
  EDFFX1 R8_reg_17_ ( .D(data_in_1[17]), .E(n6), .CK(clk), .Q(R8[17]) );
  EDFFX1 R8_reg_16_ ( .D(data_in_1[16]), .E(n6), .CK(clk), .Q(R8[16]) );
  EDFFX1 R8_reg_15_ ( .D(data_in_1[15]), .E(n6), .CK(clk), .Q(R8[15]) );
  EDFFX1 R8_reg_14_ ( .D(data_in_1[14]), .E(n6), .CK(clk), .Q(R8[14]) );
  EDFFX1 R8_reg_13_ ( .D(data_in_1[13]), .E(n6), .CK(clk), .Q(R8[13]) );
  EDFFX1 R8_reg_12_ ( .D(data_in_1[12]), .E(n6), .CK(clk), .Q(R8[12]) );
  EDFFX1 R8_reg_11_ ( .D(data_in_1[11]), .E(n6), .CK(clk), .Q(R8[11]) );
  EDFFX1 R8_reg_10_ ( .D(data_in_1[10]), .E(n6), .CK(clk), .Q(R8[10]) );
  EDFFX1 R8_reg_9_ ( .D(data_in_1[9]), .E(n6), .CK(clk), .Q(R8[9]) );
  EDFFX1 R8_reg_8_ ( .D(data_in_1[8]), .E(n6), .CK(clk), .Q(R8[8]) );
  EDFFX1 R8_reg_7_ ( .D(data_in_1[7]), .E(n6), .CK(clk), .Q(R8[7]) );
  EDFFX1 R8_reg_6_ ( .D(data_in_1[6]), .E(n6), .CK(clk), .Q(R8[6]) );
  EDFFX1 R8_reg_5_ ( .D(data_in_1[5]), .E(n6), .CK(clk), .Q(R8[5]) );
  EDFFX1 R8_reg_4_ ( .D(data_in_1[4]), .E(n6), .CK(clk), .Q(R8[4]) );
  EDFFX1 R8_reg_3_ ( .D(data_in_1[3]), .E(n6), .CK(clk), .Q(R8[3]) );
  EDFFX1 R8_reg_2_ ( .D(data_in_1[2]), .E(n6), .CK(clk), .Q(R8[2]) );
  EDFFX1 R8_reg_1_ ( .D(data_in_1[1]), .E(n6), .CK(clk), .Q(R8[1]) );
  EDFFX1 R8_reg_0_ ( .D(data_in_1[0]), .E(n6), .CK(clk), .Q(R8[0]) );
  EDFFX1 R12_reg_33_ ( .D(data_in_1[33]), .E(n3), .CK(clk), .Q(R12[33]) );
  EDFFX1 R12_reg_32_ ( .D(data_in_1[32]), .E(n3), .CK(clk), .Q(R12[32]) );
  EDFFX1 R12_reg_31_ ( .D(data_in_1[31]), .E(n3), .CK(clk), .Q(R12[31]) );
  EDFFX1 R12_reg_30_ ( .D(data_in_1[30]), .E(n3), .CK(clk), .Q(R12[30]) );
  EDFFX1 R12_reg_29_ ( .D(data_in_1[29]), .E(n3), .CK(clk), .Q(R12[29]) );
  EDFFX1 R12_reg_28_ ( .D(data_in_1[28]), .E(n3), .CK(clk), .Q(R12[28]) );
  EDFFX1 R12_reg_27_ ( .D(data_in_1[27]), .E(n3), .CK(clk), .Q(R12[27]) );
  EDFFX1 R12_reg_26_ ( .D(data_in_1[26]), .E(n3), .CK(clk), .Q(R12[26]) );
  EDFFX1 R12_reg_25_ ( .D(data_in_1[25]), .E(n3), .CK(clk), .Q(R12[25]) );
  EDFFX1 R12_reg_24_ ( .D(data_in_1[24]), .E(n3), .CK(clk), .Q(R12[24]) );
  EDFFX1 R12_reg_23_ ( .D(data_in_1[23]), .E(n3), .CK(clk), .Q(R12[23]) );
  EDFFX1 R12_reg_22_ ( .D(data_in_1[22]), .E(n3), .CK(clk), .Q(R12[22]) );
  EDFFX1 R12_reg_21_ ( .D(data_in_1[21]), .E(n3), .CK(clk), .Q(R12[21]) );
  EDFFX1 R12_reg_20_ ( .D(data_in_1[20]), .E(n3), .CK(clk), .Q(R12[20]) );
  EDFFX1 R12_reg_19_ ( .D(data_in_1[19]), .E(n3), .CK(clk), .Q(R12[19]) );
  EDFFX1 R12_reg_18_ ( .D(data_in_1[18]), .E(n3), .CK(clk), .Q(R12[18]) );
  EDFFX1 R12_reg_17_ ( .D(data_in_1[17]), .E(n3), .CK(clk), .Q(R12[17]) );
  EDFFX1 R12_reg_16_ ( .D(data_in_1[16]), .E(n3), .CK(clk), .Q(R12[16]) );
  EDFFX1 R12_reg_15_ ( .D(data_in_1[15]), .E(n3), .CK(clk), .Q(R12[15]) );
  EDFFX1 R12_reg_14_ ( .D(data_in_1[14]), .E(n3), .CK(clk), .Q(R12[14]) );
  EDFFX1 R12_reg_13_ ( .D(data_in_1[13]), .E(n3), .CK(clk), .Q(R12[13]) );
  EDFFX1 R12_reg_12_ ( .D(data_in_1[12]), .E(n3), .CK(clk), .Q(R12[12]) );
  EDFFX1 R12_reg_11_ ( .D(data_in_1[11]), .E(n3), .CK(clk), .Q(R12[11]) );
  EDFFX1 R12_reg_10_ ( .D(data_in_1[10]), .E(n3), .CK(clk), .Q(R12[10]) );
  EDFFX1 R12_reg_9_ ( .D(data_in_1[9]), .E(n3), .CK(clk), .Q(R12[9]) );
  EDFFX1 R12_reg_8_ ( .D(data_in_1[8]), .E(n3), .CK(clk), .Q(R12[8]) );
  EDFFX1 R12_reg_7_ ( .D(data_in_1[7]), .E(n3), .CK(clk), .Q(R12[7]) );
  EDFFX1 R12_reg_6_ ( .D(data_in_1[6]), .E(n3), .CK(clk), .Q(R12[6]) );
  EDFFX1 R12_reg_5_ ( .D(data_in_1[5]), .E(n3), .CK(clk), .Q(R12[5]) );
  EDFFX1 R12_reg_4_ ( .D(data_in_1[4]), .E(n3), .CK(clk), .Q(R12[4]) );
  EDFFX1 R12_reg_3_ ( .D(data_in_1[3]), .E(n3), .CK(clk), .Q(R12[3]) );
  EDFFX1 R12_reg_2_ ( .D(data_in_1[2]), .E(n3), .CK(clk), .Q(R12[2]) );
  EDFFX1 R12_reg_1_ ( .D(data_in_1[1]), .E(n3), .CK(clk), .Q(R12[1]) );
  EDFFX1 R12_reg_0_ ( .D(data_in_1[0]), .E(n3), .CK(clk), .Q(R12[0]) );
  EDFFX1 R15_reg_33_ ( .D(data_in_1[33]), .E(n993), .CK(clk), .Q(R15[33]) );
  EDFFX1 R15_reg_32_ ( .D(data_in_1[32]), .E(n993), .CK(clk), .Q(R15[32]) );
  EDFFX1 R15_reg_31_ ( .D(data_in_1[31]), .E(n993), .CK(clk), .Q(R15[31]) );
  EDFFX1 R15_reg_30_ ( .D(data_in_1[30]), .E(n993), .CK(clk), .Q(R15[30]) );
  EDFFX1 R15_reg_29_ ( .D(data_in_1[29]), .E(n993), .CK(clk), .Q(R15[29]) );
  EDFFX1 R15_reg_28_ ( .D(data_in_1[28]), .E(n993), .CK(clk), .Q(R15[28]) );
  EDFFX1 R15_reg_27_ ( .D(data_in_1[27]), .E(n993), .CK(clk), .Q(R15[27]) );
  EDFFX1 R15_reg_26_ ( .D(data_in_1[26]), .E(n993), .CK(clk), .Q(R15[26]) );
  EDFFX1 R15_reg_25_ ( .D(data_in_1[25]), .E(n993), .CK(clk), .Q(R15[25]) );
  EDFFX1 R15_reg_24_ ( .D(data_in_1[24]), .E(n993), .CK(clk), .Q(R15[24]) );
  EDFFX1 R15_reg_23_ ( .D(data_in_1[23]), .E(n993), .CK(clk), .Q(R15[23]) );
  EDFFX1 R15_reg_22_ ( .D(data_in_1[22]), .E(n993), .CK(clk), .Q(R15[22]) );
  EDFFX1 R15_reg_21_ ( .D(data_in_1[21]), .E(n993), .CK(clk), .Q(R15[21]) );
  EDFFX1 R15_reg_20_ ( .D(data_in_1[20]), .E(n993), .CK(clk), .Q(R15[20]) );
  EDFFX1 R15_reg_19_ ( .D(data_in_1[19]), .E(n993), .CK(clk), .Q(R15[19]) );
  EDFFX1 R15_reg_18_ ( .D(data_in_1[18]), .E(n993), .CK(clk), .Q(R15[18]) );
  EDFFX1 R15_reg_17_ ( .D(data_in_1[17]), .E(n993), .CK(clk), .Q(R15[17]) );
  EDFFX1 R15_reg_16_ ( .D(data_in_1[16]), .E(n993), .CK(clk), .Q(R15[16]) );
  EDFFX1 R15_reg_15_ ( .D(data_in_1[15]), .E(n993), .CK(clk), .Q(R15[15]) );
  EDFFX1 R15_reg_14_ ( .D(data_in_1[14]), .E(n993), .CK(clk), .Q(R15[14]) );
  EDFFX1 R15_reg_13_ ( .D(data_in_1[13]), .E(n993), .CK(clk), .Q(R15[13]) );
  EDFFX1 R15_reg_12_ ( .D(data_in_1[12]), .E(n993), .CK(clk), .Q(R15[12]) );
  EDFFX1 R15_reg_11_ ( .D(data_in_1[11]), .E(n993), .CK(clk), .Q(R15[11]) );
  EDFFX1 R15_reg_10_ ( .D(data_in_1[10]), .E(n993), .CK(clk), .Q(R15[10]) );
  EDFFX1 R15_reg_9_ ( .D(data_in_1[9]), .E(n993), .CK(clk), .Q(R15[9]) );
  EDFFX1 R15_reg_8_ ( .D(data_in_1[8]), .E(n993), .CK(clk), .Q(R15[8]) );
  EDFFX1 R15_reg_7_ ( .D(data_in_1[7]), .E(n993), .CK(clk), .Q(R15[7]) );
  EDFFX1 R15_reg_6_ ( .D(data_in_1[6]), .E(n993), .CK(clk), .Q(R15[6]) );
  EDFFX1 R15_reg_5_ ( .D(data_in_1[5]), .E(n993), .CK(clk), .Q(R15[5]) );
  EDFFX1 R15_reg_4_ ( .D(data_in_1[4]), .E(n993), .CK(clk), .Q(R15[4]) );
  EDFFX1 R15_reg_3_ ( .D(data_in_1[3]), .E(n993), .CK(clk), .Q(R15[3]) );
  EDFFX1 R15_reg_2_ ( .D(data_in_1[2]), .E(n993), .CK(clk), .Q(R15[2]) );
  EDFFX1 R15_reg_1_ ( .D(data_in_1[1]), .E(n993), .CK(clk), .Q(R15[1]) );
  EDFFX1 R15_reg_0_ ( .D(data_in_1[0]), .E(n993), .CK(clk), .Q(R15[0]) );
  EDFFX1 R3_reg_33_ ( .D(data_in_1[33]), .E(n5), .CK(clk), .Q(R3[33]) );
  EDFFX1 R3_reg_32_ ( .D(data_in_1[32]), .E(n5), .CK(clk), .Q(R3[32]) );
  EDFFX1 R3_reg_31_ ( .D(data_in_1[31]), .E(n5), .CK(clk), .Q(R3[31]) );
  EDFFX1 R3_reg_30_ ( .D(data_in_1[30]), .E(n5), .CK(clk), .Q(R3[30]) );
  EDFFX1 R3_reg_29_ ( .D(data_in_1[29]), .E(n5), .CK(clk), .Q(R3[29]) );
  EDFFX1 R3_reg_28_ ( .D(data_in_1[28]), .E(n5), .CK(clk), .Q(R3[28]) );
  EDFFX1 R3_reg_27_ ( .D(data_in_1[27]), .E(n5), .CK(clk), .Q(R3[27]) );
  EDFFX1 R3_reg_26_ ( .D(data_in_1[26]), .E(n5), .CK(clk), .Q(R3[26]) );
  EDFFX1 R3_reg_25_ ( .D(data_in_1[25]), .E(n5), .CK(clk), .Q(R3[25]) );
  EDFFX1 R3_reg_24_ ( .D(data_in_1[24]), .E(n5), .CK(clk), .Q(R3[24]) );
  EDFFX1 R3_reg_23_ ( .D(data_in_1[23]), .E(n5), .CK(clk), .Q(R3[23]) );
  EDFFX1 R3_reg_22_ ( .D(data_in_1[22]), .E(n5), .CK(clk), .Q(R3[22]) );
  EDFFX1 R3_reg_21_ ( .D(data_in_1[21]), .E(n5), .CK(clk), .Q(R3[21]) );
  EDFFX1 R3_reg_20_ ( .D(data_in_1[20]), .E(n5), .CK(clk), .Q(R3[20]) );
  EDFFX1 R3_reg_19_ ( .D(data_in_1[19]), .E(n5), .CK(clk), .Q(R3[19]) );
  EDFFX1 R3_reg_18_ ( .D(data_in_1[18]), .E(n5), .CK(clk), .Q(R3[18]) );
  EDFFX1 R3_reg_17_ ( .D(data_in_1[17]), .E(n5), .CK(clk), .Q(R3[17]) );
  EDFFX1 R3_reg_16_ ( .D(data_in_1[16]), .E(n5), .CK(clk), .Q(R3[16]) );
  EDFFX1 R3_reg_15_ ( .D(data_in_1[15]), .E(n5), .CK(clk), .Q(R3[15]) );
  EDFFX1 R3_reg_14_ ( .D(data_in_1[14]), .E(n5), .CK(clk), .Q(R3[14]) );
  EDFFX1 R3_reg_13_ ( .D(data_in_1[13]), .E(n5), .CK(clk), .Q(R3[13]) );
  EDFFX1 R3_reg_12_ ( .D(data_in_1[12]), .E(n5), .CK(clk), .Q(R3[12]) );
  EDFFX1 R3_reg_11_ ( .D(data_in_1[11]), .E(n5), .CK(clk), .Q(R3[11]) );
  EDFFX1 R3_reg_10_ ( .D(data_in_1[10]), .E(n5), .CK(clk), .Q(R3[10]) );
  EDFFX1 R3_reg_9_ ( .D(data_in_1[9]), .E(n5), .CK(clk), .Q(R3[9]) );
  EDFFX1 R3_reg_8_ ( .D(data_in_1[8]), .E(n5), .CK(clk), .Q(R3[8]) );
  EDFFX1 R3_reg_7_ ( .D(data_in_1[7]), .E(n5), .CK(clk), .Q(R3[7]) );
  EDFFX1 R3_reg_6_ ( .D(data_in_1[6]), .E(n5), .CK(clk), .Q(R3[6]) );
  EDFFX1 R3_reg_5_ ( .D(data_in_1[5]), .E(n5), .CK(clk), .Q(R3[5]) );
  EDFFX1 R3_reg_4_ ( .D(data_in_1[4]), .E(n5), .CK(clk), .Q(R3[4]) );
  EDFFX1 R3_reg_3_ ( .D(data_in_1[3]), .E(n5), .CK(clk), .Q(R3[3]) );
  EDFFX1 R3_reg_2_ ( .D(data_in_1[2]), .E(n5), .CK(clk), .Q(R3[2]) );
  EDFFX1 R3_reg_1_ ( .D(data_in_1[1]), .E(n5), .CK(clk), .Q(R3[1]) );
  EDFFX1 R3_reg_0_ ( .D(data_in_1[0]), .E(n5), .CK(clk), .Q(R3[0]) );
  EDFFX1 R7_reg_33_ ( .D(data_in_1[33]), .E(n979), .CK(clk), .Q(R7[33]) );
  EDFFX1 R7_reg_32_ ( .D(data_in_1[32]), .E(n979), .CK(clk), .Q(R7[32]) );
  EDFFX1 R7_reg_31_ ( .D(data_in_1[31]), .E(n979), .CK(clk), .Q(R7[31]) );
  EDFFX1 R7_reg_30_ ( .D(data_in_1[30]), .E(n979), .CK(clk), .Q(R7[30]) );
  EDFFX1 R7_reg_29_ ( .D(data_in_1[29]), .E(n979), .CK(clk), .Q(R7[29]) );
  EDFFX1 R7_reg_28_ ( .D(data_in_1[28]), .E(n979), .CK(clk), .Q(R7[28]) );
  EDFFX1 R7_reg_27_ ( .D(data_in_1[27]), .E(n979), .CK(clk), .Q(R7[27]) );
  EDFFX1 R7_reg_26_ ( .D(data_in_1[26]), .E(n979), .CK(clk), .Q(R7[26]) );
  EDFFX1 R7_reg_25_ ( .D(data_in_1[25]), .E(n979), .CK(clk), .Q(R7[25]) );
  EDFFX1 R7_reg_24_ ( .D(data_in_1[24]), .E(n979), .CK(clk), .Q(R7[24]) );
  EDFFX1 R7_reg_23_ ( .D(data_in_1[23]), .E(n979), .CK(clk), .Q(R7[23]) );
  EDFFX1 R7_reg_22_ ( .D(data_in_1[22]), .E(n979), .CK(clk), .Q(R7[22]) );
  EDFFX1 R7_reg_21_ ( .D(data_in_1[21]), .E(n979), .CK(clk), .Q(R7[21]) );
  EDFFX1 R7_reg_20_ ( .D(data_in_1[20]), .E(n979), .CK(clk), .Q(R7[20]) );
  EDFFX1 R7_reg_19_ ( .D(data_in_1[19]), .E(n979), .CK(clk), .Q(R7[19]) );
  EDFFX1 R7_reg_18_ ( .D(data_in_1[18]), .E(n979), .CK(clk), .Q(R7[18]) );
  EDFFX1 R7_reg_17_ ( .D(data_in_1[17]), .E(n979), .CK(clk), .Q(R7[17]) );
  EDFFX1 R7_reg_16_ ( .D(data_in_1[16]), .E(n979), .CK(clk), .Q(R7[16]) );
  EDFFX1 R7_reg_15_ ( .D(data_in_1[15]), .E(n979), .CK(clk), .Q(R7[15]) );
  EDFFX1 R7_reg_14_ ( .D(data_in_1[14]), .E(n979), .CK(clk), .Q(R7[14]) );
  EDFFX1 R7_reg_13_ ( .D(data_in_1[13]), .E(n979), .CK(clk), .Q(R7[13]) );
  EDFFX1 R7_reg_12_ ( .D(data_in_1[12]), .E(n979), .CK(clk), .Q(R7[12]) );
  EDFFX1 R7_reg_11_ ( .D(data_in_1[11]), .E(n979), .CK(clk), .Q(R7[11]) );
  EDFFX1 R7_reg_10_ ( .D(data_in_1[10]), .E(n979), .CK(clk), .Q(R7[10]) );
  EDFFX1 R7_reg_9_ ( .D(data_in_1[9]), .E(n979), .CK(clk), .Q(R7[9]) );
  EDFFX1 R7_reg_8_ ( .D(data_in_1[8]), .E(n979), .CK(clk), .Q(R7[8]) );
  EDFFX1 R7_reg_7_ ( .D(data_in_1[7]), .E(n979), .CK(clk), .Q(R7[7]) );
  EDFFX1 R7_reg_6_ ( .D(data_in_1[6]), .E(n979), .CK(clk), .Q(R7[6]) );
  EDFFX1 R7_reg_5_ ( .D(data_in_1[5]), .E(n979), .CK(clk), .Q(R7[5]) );
  EDFFX1 R7_reg_4_ ( .D(data_in_1[4]), .E(n979), .CK(clk), .Q(R7[4]) );
  EDFFX1 R7_reg_3_ ( .D(data_in_1[3]), .E(n979), .CK(clk), .Q(R7[3]) );
  EDFFX1 R7_reg_2_ ( .D(data_in_1[2]), .E(n979), .CK(clk), .Q(R7[2]) );
  EDFFX1 R7_reg_1_ ( .D(data_in_1[1]), .E(n979), .CK(clk), .Q(R7[1]) );
  EDFFX1 R7_reg_0_ ( .D(data_in_1[0]), .E(n979), .CK(clk), .Q(R7[0]) );
  EDFFX1 R11_reg_33_ ( .D(data_in_1[33]), .E(n4), .CK(clk), .Q(R11[33]) );
  EDFFX1 R11_reg_32_ ( .D(data_in_1[32]), .E(n4), .CK(clk), .Q(R11[32]) );
  EDFFX1 R11_reg_31_ ( .D(data_in_1[31]), .E(n4), .CK(clk), .Q(R11[31]) );
  EDFFX1 R11_reg_30_ ( .D(data_in_1[30]), .E(n4), .CK(clk), .Q(R11[30]) );
  EDFFX1 R11_reg_29_ ( .D(data_in_1[29]), .E(n4), .CK(clk), .Q(R11[29]) );
  EDFFX1 R11_reg_28_ ( .D(data_in_1[28]), .E(n4), .CK(clk), .Q(R11[28]) );
  EDFFX1 R11_reg_27_ ( .D(data_in_1[27]), .E(n4), .CK(clk), .Q(R11[27]) );
  EDFFX1 R11_reg_26_ ( .D(data_in_1[26]), .E(n4), .CK(clk), .Q(R11[26]) );
  EDFFX1 R11_reg_25_ ( .D(data_in_1[25]), .E(n4), .CK(clk), .Q(R11[25]) );
  EDFFX1 R11_reg_24_ ( .D(data_in_1[24]), .E(n4), .CK(clk), .Q(R11[24]) );
  EDFFX1 R11_reg_23_ ( .D(data_in_1[23]), .E(n4), .CK(clk), .Q(R11[23]) );
  EDFFX1 R11_reg_22_ ( .D(data_in_1[22]), .E(n4), .CK(clk), .Q(R11[22]) );
  EDFFX1 R11_reg_21_ ( .D(data_in_1[21]), .E(n4), .CK(clk), .Q(R11[21]) );
  EDFFX1 R11_reg_20_ ( .D(data_in_1[20]), .E(n4), .CK(clk), .Q(R11[20]) );
  EDFFX1 R11_reg_19_ ( .D(data_in_1[19]), .E(n4), .CK(clk), .Q(R11[19]) );
  EDFFX1 R11_reg_18_ ( .D(data_in_1[18]), .E(n4), .CK(clk), .Q(R11[18]) );
  EDFFX1 R11_reg_17_ ( .D(data_in_1[17]), .E(n4), .CK(clk), .Q(R11[17]) );
  EDFFX1 R11_reg_16_ ( .D(data_in_1[16]), .E(n4), .CK(clk), .Q(R11[16]) );
  EDFFX1 R11_reg_15_ ( .D(data_in_1[15]), .E(n4), .CK(clk), .Q(R11[15]) );
  EDFFX1 R11_reg_14_ ( .D(data_in_1[14]), .E(n4), .CK(clk), .Q(R11[14]) );
  EDFFX1 R11_reg_13_ ( .D(data_in_1[13]), .E(n4), .CK(clk), .Q(R11[13]) );
  EDFFX1 R11_reg_12_ ( .D(data_in_1[12]), .E(n4), .CK(clk), .Q(R11[12]) );
  EDFFX1 R11_reg_11_ ( .D(data_in_1[11]), .E(n4), .CK(clk), .Q(R11[11]) );
  EDFFX1 R11_reg_10_ ( .D(data_in_1[10]), .E(n4), .CK(clk), .Q(R11[10]) );
  EDFFX1 R11_reg_9_ ( .D(data_in_1[9]), .E(n4), .CK(clk), .Q(R11[9]) );
  EDFFX1 R11_reg_8_ ( .D(data_in_1[8]), .E(n4), .CK(clk), .Q(R11[8]) );
  EDFFX1 R11_reg_7_ ( .D(data_in_1[7]), .E(n4), .CK(clk), .Q(R11[7]) );
  EDFFX1 R11_reg_6_ ( .D(data_in_1[6]), .E(n4), .CK(clk), .Q(R11[6]) );
  EDFFX1 R11_reg_5_ ( .D(data_in_1[5]), .E(n4), .CK(clk), .Q(R11[5]) );
  EDFFX1 R11_reg_4_ ( .D(data_in_1[4]), .E(n4), .CK(clk), .Q(R11[4]) );
  EDFFX1 R11_reg_3_ ( .D(data_in_1[3]), .E(n4), .CK(clk), .Q(R11[3]) );
  EDFFX1 R11_reg_2_ ( .D(data_in_1[2]), .E(n4), .CK(clk), .Q(R11[2]) );
  EDFFX1 R11_reg_1_ ( .D(data_in_1[1]), .E(n4), .CK(clk), .Q(R11[1]) );
  EDFFX1 R11_reg_0_ ( .D(data_in_1[0]), .E(n4), .CK(clk), .Q(R11[0]) );
  DFFRHQX1 s_p_flag_out_reg ( .D(n3), .CK(clk), .RN(rst_n), .Q(s_p_flag_out)
         );
  DFFHQX1 data_out_1_reg_33_ ( .D(n934), .CK(clk), .Q(data_out_1[33]) );
  DFFHQX1 data_out_1_reg_32_ ( .D(n935), .CK(clk), .Q(data_out_1[32]) );
  DFFHQX1 data_out_1_reg_16_ ( .D(n951), .CK(clk), .Q(data_out_1[16]) );
  DFFHQX1 data_out_1_reg_15_ ( .D(n952), .CK(clk), .Q(data_out_1[15]) );
  DFFHQX1 data_out_1_reg_30_ ( .D(n937), .CK(clk), .Q(data_out_1[30]) );
  DFFHQX1 data_out_1_reg_13_ ( .D(n954), .CK(clk), .Q(data_out_1[13]) );
  JKFFRXL counter_reg_0_ ( .J(1'b1), .K(1'b1), .CK(clk), .RN(rst_n), .Q(
        counter[0]), .QN(n550) );
  DFFHQX1 data_out_1_reg_31_ ( .D(n936), .CK(clk), .Q(data_out_1[31]) );
  DFFHQX1 data_out_1_reg_29_ ( .D(n938), .CK(clk), .Q(data_out_1[29]) );
  DFFHQX1 data_out_1_reg_28_ ( .D(n939), .CK(clk), .Q(data_out_1[28]) );
  DFFHQX1 data_out_1_reg_27_ ( .D(n940), .CK(clk), .Q(data_out_1[27]) );
  DFFHQX1 data_out_1_reg_14_ ( .D(n953), .CK(clk), .Q(data_out_1[14]) );
  DFFHQX1 data_out_1_reg_12_ ( .D(n955), .CK(clk), .Q(data_out_1[12]) );
  DFFHQX1 data_out_1_reg_11_ ( .D(n956), .CK(clk), .Q(data_out_1[11]) );
  DFFHQX1 data_out_1_reg_10_ ( .D(n957), .CK(clk), .Q(data_out_1[10]) );
  DFFRHQX1 counter_reg_3_ ( .D(N15), .CK(clk), .RN(rst_n), .Q(counter[3]) );
  DFFRHQX1 counter_reg_1_ ( .D(N13), .CK(clk), .RN(rst_n), .Q(counter[1]) );
  DFFRHQX1 counter_reg_2_ ( .D(N14), .CK(clk), .RN(rst_n), .Q(counter[2]) );
  DFFHQX1 data_out_1_reg_26_ ( .D(n941), .CK(clk), .Q(data_out_1[26]) );
  DFFHQX1 data_out_1_reg_25_ ( .D(n942), .CK(clk), .Q(data_out_1[25]) );
  DFFHQX1 data_out_1_reg_24_ ( .D(n943), .CK(clk), .Q(data_out_1[24]) );
  DFFHQX1 data_out_1_reg_23_ ( .D(n944), .CK(clk), .Q(data_out_1[23]) );
  DFFHQX1 data_out_1_reg_22_ ( .D(n945), .CK(clk), .Q(data_out_1[22]) );
  DFFHQX1 data_out_1_reg_21_ ( .D(n946), .CK(clk), .Q(data_out_1[21]) );
  DFFHQX1 data_out_1_reg_9_ ( .D(n958), .CK(clk), .Q(data_out_1[9]) );
  DFFHQX1 data_out_1_reg_8_ ( .D(n959), .CK(clk), .Q(data_out_1[8]) );
  DFFHQX1 data_out_1_reg_7_ ( .D(n960), .CK(clk), .Q(data_out_1[7]) );
  DFFHQX1 data_out_1_reg_6_ ( .D(n961), .CK(clk), .Q(data_out_1[6]) );
  DFFHQX1 data_out_1_reg_5_ ( .D(n962), .CK(clk), .Q(data_out_1[5]) );
  DFFHQX1 data_out_1_reg_4_ ( .D(n963), .CK(clk), .Q(data_out_1[4]) );
  DFFHQX1 data_out_1_reg_20_ ( .D(n947), .CK(clk), .Q(data_out_1[20]) );
  DFFHQX1 data_out_1_reg_19_ ( .D(n948), .CK(clk), .Q(data_out_1[19]) );
  DFFHQX1 data_out_1_reg_18_ ( .D(n949), .CK(clk), .Q(data_out_1[18]) );
  DFFHQX1 data_out_1_reg_17_ ( .D(n950), .CK(clk), .Q(data_out_1[17]) );
  DFFHQX1 data_out_1_reg_3_ ( .D(n964), .CK(clk), .Q(data_out_1[3]) );
  DFFHQX1 data_out_1_reg_2_ ( .D(n965), .CK(clk), .Q(data_out_1[2]) );
  DFFHQX1 data_out_1_reg_1_ ( .D(n966), .CK(clk), .Q(data_out_1[1]) );
  DFFHQX1 data_out_1_reg_0_ ( .D(n967), .CK(clk), .Q(data_out_1[0]) );
  DFFHQX1 data_out_1_reg_66_ ( .D(n901), .CK(clk), .Q(data_out_1[66]) );
  DFFHQX1 data_out_1_reg_65_ ( .D(n902), .CK(clk), .Q(data_out_1[65]) );
  DFFHQX1 data_out_1_reg_64_ ( .D(n903), .CK(clk), .Q(data_out_1[64]) );
  DFFHQX1 data_out_1_reg_49_ ( .D(n918), .CK(clk), .Q(data_out_1[49]) );
  DFFHQX1 data_out_1_reg_48_ ( .D(n919), .CK(clk), .Q(data_out_1[48]) );
  DFFHQX1 data_out_1_reg_47_ ( .D(n920), .CK(clk), .Q(data_out_1[47]) );
  DFFHQX1 data_out_1_reg_100_ ( .D(n867), .CK(clk), .Q(data_out_1[100]) );
  DFFHQX1 data_out_1_reg_99_ ( .D(n868), .CK(clk), .Q(data_out_1[99]) );
  DFFHQX1 data_out_1_reg_98_ ( .D(n869), .CK(clk), .Q(data_out_1[98]) );
  DFFHQX1 data_out_1_reg_83_ ( .D(n884), .CK(clk), .Q(data_out_1[83]) );
  DFFHQX1 data_out_1_reg_82_ ( .D(n885), .CK(clk), .Q(data_out_1[82]) );
  DFFHQX1 data_out_1_reg_134_ ( .D(n833), .CK(clk), .Q(data_out_1[134]) );
  DFFHQX1 data_out_1_reg_133_ ( .D(n834), .CK(clk), .Q(data_out_1[133]) );
  DFFHQX1 data_out_1_reg_132_ ( .D(n835), .CK(clk), .Q(data_out_1[132]) );
  DFFHQX1 data_out_1_reg_117_ ( .D(n850), .CK(clk), .Q(data_out_1[117]) );
  DFFHQX1 data_out_1_reg_116_ ( .D(n851), .CK(clk), .Q(data_out_1[116]) );
  DFFHQX1 data_out_1_reg_63_ ( .D(n904), .CK(clk), .Q(data_out_1[63]) );
  DFFHQX1 data_out_1_reg_62_ ( .D(n905), .CK(clk), .Q(data_out_1[62]) );
  DFFHQX1 data_out_1_reg_61_ ( .D(n906), .CK(clk), .Q(data_out_1[61]) );
  DFFHQX1 data_out_1_reg_60_ ( .D(n907), .CK(clk), .Q(data_out_1[60]) );
  DFFHQX1 data_out_1_reg_46_ ( .D(n921), .CK(clk), .Q(data_out_1[46]) );
  DFFHQX1 data_out_1_reg_45_ ( .D(n922), .CK(clk), .Q(data_out_1[45]) );
  DFFHQX1 data_out_1_reg_44_ ( .D(n923), .CK(clk), .Q(data_out_1[44]) );
  DFFHQX1 data_out_1_reg_43_ ( .D(n924), .CK(clk), .Q(data_out_1[43]) );
  DFFHQX1 data_out_1_reg_97_ ( .D(n870), .CK(clk), .Q(data_out_1[97]) );
  DFFHQX1 data_out_1_reg_96_ ( .D(n871), .CK(clk), .Q(data_out_1[96]) );
  DFFHQX1 data_out_1_reg_95_ ( .D(n872), .CK(clk), .Q(data_out_1[95]) );
  DFFHQX1 data_out_1_reg_94_ ( .D(n873), .CK(clk), .Q(data_out_1[94]) );
  DFFHQX1 data_out_1_reg_81_ ( .D(n886), .CK(clk), .Q(data_out_1[81]) );
  DFFHQX1 data_out_1_reg_80_ ( .D(n887), .CK(clk), .Q(data_out_1[80]) );
  DFFHQX1 data_out_1_reg_79_ ( .D(n888), .CK(clk), .Q(data_out_1[79]) );
  DFFHQX1 data_out_1_reg_78_ ( .D(n889), .CK(clk), .Q(data_out_1[78]) );
  DFFHQX1 data_out_1_reg_77_ ( .D(n890), .CK(clk), .Q(data_out_1[77]) );
  DFFHQX1 data_out_1_reg_131_ ( .D(n836), .CK(clk), .Q(data_out_1[131]) );
  DFFHQX1 data_out_1_reg_130_ ( .D(n837), .CK(clk), .Q(data_out_1[130]) );
  DFFHQX1 data_out_1_reg_129_ ( .D(n838), .CK(clk), .Q(data_out_1[129]) );
  DFFHQX1 data_out_1_reg_128_ ( .D(n839), .CK(clk), .Q(data_out_1[128]) );
  DFFHQX1 data_out_1_reg_115_ ( .D(n852), .CK(clk), .Q(data_out_1[115]) );
  DFFHQX1 data_out_1_reg_114_ ( .D(n853), .CK(clk), .Q(data_out_1[114]) );
  DFFHQX1 data_out_1_reg_113_ ( .D(n854), .CK(clk), .Q(data_out_1[113]) );
  DFFHQX1 data_out_1_reg_112_ ( .D(n855), .CK(clk), .Q(data_out_1[112]) );
  DFFHQX1 data_out_1_reg_111_ ( .D(n856), .CK(clk), .Q(data_out_1[111]) );
  DFFHQX1 data_out_1_reg_59_ ( .D(n908), .CK(clk), .Q(data_out_1[59]) );
  DFFHQX1 data_out_1_reg_58_ ( .D(n909), .CK(clk), .Q(data_out_1[58]) );
  DFFHQX1 data_out_1_reg_57_ ( .D(n910), .CK(clk), .Q(data_out_1[57]) );
  DFFHQX1 data_out_1_reg_42_ ( .D(n925), .CK(clk), .Q(data_out_1[42]) );
  DFFHQX1 data_out_1_reg_41_ ( .D(n926), .CK(clk), .Q(data_out_1[41]) );
  DFFHQX1 data_out_1_reg_40_ ( .D(n927), .CK(clk), .Q(data_out_1[40]) );
  DFFHQX1 data_out_1_reg_93_ ( .D(n874), .CK(clk), .Q(data_out_1[93]) );
  DFFHQX1 data_out_1_reg_92_ ( .D(n875), .CK(clk), .Q(data_out_1[92]) );
  DFFHQX1 data_out_1_reg_91_ ( .D(n876), .CK(clk), .Q(data_out_1[91]) );
  DFFHQX1 data_out_1_reg_76_ ( .D(n891), .CK(clk), .Q(data_out_1[76]) );
  DFFHQX1 data_out_1_reg_75_ ( .D(n892), .CK(clk), .Q(data_out_1[75]) );
  DFFHQX1 data_out_1_reg_74_ ( .D(n893), .CK(clk), .Q(data_out_1[74]) );
  DFFHQX1 data_out_1_reg_127_ ( .D(n840), .CK(clk), .Q(data_out_1[127]) );
  DFFHQX1 data_out_1_reg_126_ ( .D(n841), .CK(clk), .Q(data_out_1[126]) );
  DFFHQX1 data_out_1_reg_125_ ( .D(n842), .CK(clk), .Q(data_out_1[125]) );
  DFFHQX1 data_out_1_reg_110_ ( .D(n857), .CK(clk), .Q(data_out_1[110]) );
  DFFHQX1 data_out_1_reg_109_ ( .D(n858), .CK(clk), .Q(data_out_1[109]) );
  DFFHQX1 data_out_1_reg_108_ ( .D(n859), .CK(clk), .Q(data_out_1[108]) );
  DFFHQX1 data_out_1_reg_56_ ( .D(n911), .CK(clk), .Q(data_out_1[56]) );
  DFFHQX1 data_out_1_reg_55_ ( .D(n912), .CK(clk), .Q(data_out_1[55]) );
  DFFHQX1 data_out_1_reg_54_ ( .D(n913), .CK(clk), .Q(data_out_1[54]) );
  DFFHQX1 data_out_1_reg_39_ ( .D(n928), .CK(clk), .Q(data_out_1[39]) );
  DFFHQX1 data_out_1_reg_38_ ( .D(n929), .CK(clk), .Q(data_out_1[38]) );
  DFFHQX1 data_out_1_reg_37_ ( .D(n930), .CK(clk), .Q(data_out_1[37]) );
  DFFHQX1 data_out_1_reg_90_ ( .D(n877), .CK(clk), .Q(data_out_1[90]) );
  DFFHQX1 data_out_1_reg_89_ ( .D(n878), .CK(clk), .Q(data_out_1[89]) );
  DFFHQX1 data_out_1_reg_88_ ( .D(n879), .CK(clk), .Q(data_out_1[88]) );
  DFFHQX1 data_out_1_reg_73_ ( .D(n894), .CK(clk), .Q(data_out_1[73]) );
  DFFHQX1 data_out_1_reg_72_ ( .D(n895), .CK(clk), .Q(data_out_1[72]) );
  DFFHQX1 data_out_1_reg_71_ ( .D(n896), .CK(clk), .Q(data_out_1[71]) );
  DFFHQX1 data_out_1_reg_124_ ( .D(n843), .CK(clk), .Q(data_out_1[124]) );
  DFFHQX1 data_out_1_reg_123_ ( .D(n844), .CK(clk), .Q(data_out_1[123]) );
  DFFHQX1 data_out_1_reg_122_ ( .D(n845), .CK(clk), .Q(data_out_1[122]) );
  DFFHQX1 data_out_1_reg_107_ ( .D(n860), .CK(clk), .Q(data_out_1[107]) );
  DFFHQX1 data_out_1_reg_106_ ( .D(n861), .CK(clk), .Q(data_out_1[106]) );
  DFFHQX1 data_out_1_reg_105_ ( .D(n862), .CK(clk), .Q(data_out_1[105]) );
  DFFHQX1 data_out_1_reg_87_ ( .D(n880), .CK(clk), .Q(data_out_1[87]) );
  DFFHQX1 data_out_1_reg_121_ ( .D(n846), .CK(clk), .Q(data_out_1[121]) );
  DFFHQX1 data_out_1_reg_119_ ( .D(n848), .CK(clk), .Q(data_out_1[119]) );
  DFFHQX1 data_out_1_reg_86_ ( .D(n881), .CK(clk), .Q(data_out_1[86]) );
  DFFHQX1 data_out_1_reg_135_ ( .D(n832), .CK(clk), .Q(data_out_1[135]) );
  DFFHQX1 data_out_1_reg_101_ ( .D(n866), .CK(clk), .Q(data_out_1[101]) );
  DFFHQX1 data_out_1_reg_84_ ( .D(n883), .CK(clk), .Q(data_out_1[84]) );
  DFFHQX1 data_out_1_reg_52_ ( .D(n915), .CK(clk), .Q(data_out_1[52]) );
  DFFHQX1 data_out_1_reg_120_ ( .D(n847), .CK(clk), .Q(data_out_1[120]) );
  DFFHQX1 data_out_1_reg_103_ ( .D(n864), .CK(clk), .Q(data_out_1[103]) );
  DFFHQX1 data_out_1_reg_35_ ( .D(n932), .CK(clk), .Q(data_out_1[35]) );
  DFFHQX1 data_out_1_reg_70_ ( .D(n897), .CK(clk), .Q(data_out_1[70]) );
  DFFHQX1 data_out_1_reg_69_ ( .D(n898), .CK(clk), .Q(data_out_1[69]) );
  DFFHQX1 data_out_1_reg_102_ ( .D(n865), .CK(clk), .Q(data_out_1[102]) );
  DFFHQX1 data_out_1_reg_36_ ( .D(n931), .CK(clk), .Q(data_out_1[36]) );
  DFFHQX1 data_out_1_reg_104_ ( .D(n863), .CK(clk), .Q(data_out_1[104]) );
  DFFHQX1 data_out_1_reg_53_ ( .D(n914), .CK(clk), .Q(data_out_1[53]) );
  DFFHQX1 data_out_1_reg_51_ ( .D(n916), .CK(clk), .Q(data_out_1[51]) );
  DFFHQX1 data_out_1_reg_50_ ( .D(n917), .CK(clk), .Q(data_out_1[50]) );
  DFFHQXL data_out_1_reg_85_ ( .D(n882), .CK(clk), .Q(data_out_1[85]) );
  DFFHQXL data_out_1_reg_68_ ( .D(n899), .CK(clk), .Q(data_out_1[68]) );
  DFFHQXL data_out_1_reg_67_ ( .D(n900), .CK(clk), .Q(data_out_1[67]) );
  DFFHQXL data_out_1_reg_118_ ( .D(n849), .CK(clk), .Q(data_out_1[118]) );
  DFFHQXL data_out_1_reg_34_ ( .D(n933), .CK(clk), .Q(data_out_1[34]) );
  OR4X2 U4 ( .A(n982), .B(n980), .C(n993), .D(n995), .Y(n1) );
  OR3XL U5 ( .A(n1006), .B(n1005), .C(n825), .Y(n2) );
  NOR3X2 U6 ( .A(n1006), .B(n1005), .C(n828), .Y(n3) );
  NOR2X1 U7 ( .A(n826), .B(n827), .Y(n4) );
  NOR2X1 U8 ( .A(n826), .B(n830), .Y(n5) );
  NOR2X1 U9 ( .A(n828), .B(n827), .Y(n6) );
  NOR2X1 U10 ( .A(n828), .B(n829), .Y(n7) );
  NOR2X1 U11 ( .A(n824), .B(n827), .Y(n8) );
  NOR2X1 U12 ( .A(n824), .B(n829), .Y(n9) );
  NOR2X1 U13 ( .A(n824), .B(n830), .Y(n10) );
  NOR2X1 U14 ( .A(n825), .B(n827), .Y(n11) );
  NOR2X1 U15 ( .A(n825), .B(n829), .Y(n12) );
  NOR2X1 U16 ( .A(n825), .B(n830), .Y(n13) );
  OR2X2 U17 ( .A(n829), .B(n826), .Y(n14) );
  AOI22XL U18 ( .A0(R11[1]), .A1(n998), .B0(data_out_1[69]), .B1(n988), .Y(
        n684) );
  AOI22XL U19 ( .A0(R11[2]), .A1(n998), .B0(data_out_1[70]), .B1(n988), .Y(
        n682) );
  AOI22XL U20 ( .A0(R15[16]), .A1(n996), .B0(data_out_1[118]), .B1(n991), .Y(
        n586) );
  AOI22XL U21 ( .A0(R11[0]), .A1(n998), .B0(data_out_1[68]), .B1(n988), .Y(
        n686) );
  AOI22XL U22 ( .A0(R11[17]), .A1(n1001), .B0(data_out_1[85]), .B1(n989), .Y(
        n652) );
  AOI22XL U23 ( .A0(R7[33]), .A1(n998), .B0(data_out_1[67]), .B1(n988), .Y(
        n688) );
  AOI22XL U24 ( .A0(R15[0]), .A1(n997), .B0(data_out_1[102]), .B1(n990), .Y(
        n618) );
  AOI22XL U25 ( .A0(R15[1]), .A1(n997), .B0(data_out_1[103]), .B1(n990), .Y(
        n616) );
  AOI22XL U26 ( .A0(R15[2]), .A1(n997), .B0(data_out_1[104]), .B1(n990), .Y(
        n614) );
  AOI22XL U27 ( .A0(R15[3]), .A1(n997), .B0(data_out_1[105]), .B1(n990), .Y(
        n612) );
  AOI22XL U28 ( .A0(R15[4]), .A1(n997), .B0(data_out_1[106]), .B1(n990), .Y(
        n610) );
  AOI22XL U29 ( .A0(R15[5]), .A1(n997), .B0(data_out_1[107]), .B1(n990), .Y(
        n608) );
  AOI22XL U30 ( .A0(R15[6]), .A1(n997), .B0(data_out_1[108]), .B1(n991), .Y(
        n606) );
  AOI22XL U31 ( .A0(R15[17]), .A1(n996), .B0(data_out_1[119]), .B1(n991), .Y(
        n584) );
  AOI22XL U32 ( .A0(R15[18]), .A1(n996), .B0(data_out_1[120]), .B1(n992), .Y(
        n582) );
  AOI22XL U33 ( .A0(R15[19]), .A1(n996), .B0(data_out_1[121]), .B1(n992), .Y(
        n580) );
  AOI22XL U34 ( .A0(R15[20]), .A1(n996), .B0(data_out_1[122]), .B1(n992), .Y(
        n578) );
  AOI22XL U35 ( .A0(R15[21]), .A1(n995), .B0(data_out_1[123]), .B1(n992), .Y(
        n576) );
  AOI22XL U36 ( .A0(R15[22]), .A1(n995), .B0(data_out_1[124]), .B1(n992), .Y(
        n574) );
  AOI22XL U37 ( .A0(R15[23]), .A1(n995), .B0(data_out_1[125]), .B1(n992), .Y(
        n572) );
  AOI22XL U38 ( .A0(R15[33]), .A1(n997), .B0(data_out_1[135]), .B1(n992), .Y(
        n551) );
  AOI22XL U39 ( .A0(R11[3]), .A1(n998), .B0(data_out_1[71]), .B1(n988), .Y(
        n680) );
  AOI22XL U40 ( .A0(R11[4]), .A1(n1000), .B0(data_out_1[72]), .B1(n990), .Y(
        n678) );
  AOI22XL U41 ( .A0(R11[5]), .A1(n1001), .B0(data_out_1[73]), .B1(n989), .Y(
        n676) );
  AOI22XL U42 ( .A0(R11[6]), .A1(n999), .B0(data_out_1[74]), .B1(n990), .Y(
        n674) );
  AOI22XL U43 ( .A0(R11[18]), .A1(n999), .B0(data_out_1[86]), .B1(n989), .Y(
        n650) );
  AOI22XL U44 ( .A0(R11[19]), .A1(n997), .B0(data_out_1[87]), .B1(n989), .Y(
        n648) );
  AOI22XL U45 ( .A0(R11[20]), .A1(n996), .B0(data_out_1[88]), .B1(n989), .Y(
        n646) );
  AOI22XL U46 ( .A0(R11[21]), .A1(n999), .B0(data_out_1[89]), .B1(n989), .Y(
        n644) );
  AOI22XL U47 ( .A0(R11[22]), .A1(n998), .B0(data_out_1[90]), .B1(n989), .Y(
        n642) );
  AOI22XL U48 ( .A0(R11[23]), .A1(n999), .B0(data_out_1[91]), .B1(n989), .Y(
        n640) );
  AOI22XL U49 ( .A0(R11[33]), .A1(n997), .B0(data_out_1[101]), .B1(n990), .Y(
        n620) );
  AOI22XL U50 ( .A0(R7[0]), .A1(n999), .B0(data_out_1[34]), .B1(n986), .Y(n754) );
  AOI22XL U51 ( .A0(R7[1]), .A1(n999), .B0(data_out_1[35]), .B1(n986), .Y(n752) );
  AOI22XL U52 ( .A0(R7[2]), .A1(n999), .B0(data_out_1[36]), .B1(n987), .Y(n750) );
  AOI22XL U53 ( .A0(R7[3]), .A1(n999), .B0(data_out_1[37]), .B1(n987), .Y(n748) );
  AOI22XL U54 ( .A0(R7[4]), .A1(n999), .B0(data_out_1[38]), .B1(n987), .Y(n746) );
  AOI22XL U55 ( .A0(R7[5]), .A1(n999), .B0(data_out_1[39]), .B1(n987), .Y(n744) );
  AOI22XL U56 ( .A0(R7[6]), .A1(n999), .B0(data_out_1[40]), .B1(n987), .Y(n742) );
  AOI22XL U57 ( .A0(R7[16]), .A1(n997), .B0(data_out_1[50]), .B1(n989), .Y(
        n722) );
  AOI22XL U58 ( .A0(R7[17]), .A1(n996), .B0(data_out_1[51]), .B1(n987), .Y(
        n720) );
  AOI22XL U59 ( .A0(R7[18]), .A1(n997), .B0(data_out_1[52]), .B1(n990), .Y(
        n718) );
  AOI22XL U60 ( .A0(R7[19]), .A1(n996), .B0(data_out_1[53]), .B1(n990), .Y(
        n716) );
  AOI22XL U61 ( .A0(R7[20]), .A1(n997), .B0(data_out_1[54]), .B1(n989), .Y(
        n714) );
  AOI22XL U62 ( .A0(R7[21]), .A1(n996), .B0(data_out_1[55]), .B1(n989), .Y(
        n712) );
  AOI22XL U63 ( .A0(R7[22]), .A1(n997), .B0(data_out_1[56]), .B1(n988), .Y(
        n710) );
  AOI22XL U64 ( .A0(R7[23]), .A1(n996), .B0(data_out_1[57]), .B1(n988), .Y(
        n708) );
  INVX1 U65 ( .A(n1), .Y(n991) );
  INVX1 U66 ( .A(n1), .Y(n992) );
  INVX1 U67 ( .A(n1), .Y(n989) );
  INVX1 U68 ( .A(n1), .Y(n990) );
  INVX1 U69 ( .A(n1), .Y(n987) );
  INVX1 U70 ( .A(n1), .Y(n988) );
  INVX1 U71 ( .A(n1), .Y(n984) );
  INVX1 U72 ( .A(n1), .Y(n985) );
  INVX1 U73 ( .A(n1), .Y(n986) );
  INVX1 U74 ( .A(n1003), .Y(n995) );
  INVX1 U75 ( .A(n1003), .Y(n996) );
  INVX1 U76 ( .A(n1003), .Y(n997) );
  INVX1 U77 ( .A(n1003), .Y(n998) );
  INVX1 U78 ( .A(n1003), .Y(n1001) );
  INVX1 U79 ( .A(n1003), .Y(n1000) );
  INVX1 U80 ( .A(n1003), .Y(n999) );
  INVX1 U81 ( .A(n1003), .Y(n1002) );
  CLKINVX3 U82 ( .A(n2), .Y(n981) );
  INVX1 U83 ( .A(n14), .Y(n979) );
  INVX1 U84 ( .A(n2), .Y(n980) );
  INVX1 U85 ( .A(n15), .Y(n993) );
  INVX1 U86 ( .A(N171), .Y(n1003) );
  CLKINVX3 U87 ( .A(n15), .Y(n994) );
  CLKINVX3 U88 ( .A(n16), .Y(n983) );
  INVX1 U89 ( .A(n16), .Y(n982) );
  NOR2X1 U90 ( .A(n830), .B(n828), .Y(N171) );
  NAND2X1 U91 ( .A(n1005), .B(n1006), .Y(n830) );
  OR3XL U92 ( .A(n1005), .B(n826), .C(n1006), .Y(n15) );
  OR3XL U93 ( .A(n1006), .B(n1005), .C(n824), .Y(n16) );
  OAI211X1 U94 ( .A0(n831), .A1(n1006), .B0(n827), .C0(n14), .Y(N15) );
  NAND2X1 U95 ( .A(n824), .B(n825), .Y(N13) );
  NAND2X1 U96 ( .A(counter[1]), .B(counter[0]), .Y(n826) );
  NAND2X1 U97 ( .A(counter[0]), .B(n1004), .Y(n825) );
  NAND2X1 U98 ( .A(n550), .B(n1004), .Y(n828) );
  INVX1 U99 ( .A(counter[2]), .Y(n1005) );
  INVX1 U100 ( .A(counter[3]), .Y(n1006) );
  INVX1 U101 ( .A(counter[1]), .Y(n1004) );
  NAND2X1 U102 ( .A(n618), .B(n619), .Y(n865) );
  AOI222X1 U103 ( .A0(R12[0]), .A1(n981), .B0(R14[0]), .B1(n994), .C0(R13[0]), 
        .C1(n983), .Y(n619) );
  NAND2X1 U104 ( .A(n616), .B(n617), .Y(n864) );
  AOI222X1 U105 ( .A0(R12[1]), .A1(n981), .B0(R14[1]), .B1(n994), .C0(R13[1]), 
        .C1(n983), .Y(n617) );
  NAND2X1 U106 ( .A(n614), .B(n615), .Y(n863) );
  AOI222X1 U107 ( .A0(R12[2]), .A1(n981), .B0(R14[2]), .B1(n994), .C0(R13[2]), 
        .C1(n983), .Y(n615) );
  NAND2X1 U108 ( .A(n612), .B(n613), .Y(n862) );
  AOI222X1 U109 ( .A0(R12[3]), .A1(n981), .B0(R14[3]), .B1(n994), .C0(R13[3]), 
        .C1(n983), .Y(n613) );
  NAND2X1 U110 ( .A(n610), .B(n611), .Y(n861) );
  AOI222X1 U111 ( .A0(R12[4]), .A1(n981), .B0(R14[4]), .B1(n994), .C0(R13[4]), 
        .C1(n983), .Y(n611) );
  NAND2X1 U112 ( .A(n608), .B(n609), .Y(n860) );
  AOI222X1 U113 ( .A0(R12[5]), .A1(n981), .B0(R14[5]), .B1(n994), .C0(R13[5]), 
        .C1(n983), .Y(n609) );
  NAND2X1 U114 ( .A(n606), .B(n607), .Y(n859) );
  AOI222X1 U115 ( .A0(R12[6]), .A1(n981), .B0(R14[6]), .B1(n994), .C0(R13[6]), 
        .C1(n983), .Y(n607) );
  NAND2X1 U116 ( .A(n604), .B(n605), .Y(n858) );
  AOI222X1 U117 ( .A0(R12[7]), .A1(n981), .B0(R14[7]), .B1(n994), .C0(R13[7]), 
        .C1(n983), .Y(n605) );
  AOI22X1 U118 ( .A0(R15[7]), .A1(n997), .B0(data_out_1[109]), .B1(n991), .Y(
        n604) );
  NAND2X1 U119 ( .A(n602), .B(n603), .Y(n857) );
  AOI222X1 U120 ( .A0(R12[8]), .A1(n981), .B0(R14[8]), .B1(n994), .C0(R13[8]), 
        .C1(n983), .Y(n603) );
  AOI22X1 U121 ( .A0(R15[8]), .A1(n996), .B0(data_out_1[110]), .B1(n991), .Y(
        n602) );
  NAND2X1 U122 ( .A(n600), .B(n601), .Y(n856) );
  AOI222X1 U123 ( .A0(R12[9]), .A1(n981), .B0(R14[9]), .B1(n994), .C0(R13[9]), 
        .C1(n983), .Y(n601) );
  AOI22X1 U124 ( .A0(R15[9]), .A1(n996), .B0(data_out_1[111]), .B1(n991), .Y(
        n600) );
  NAND2X1 U125 ( .A(n598), .B(n599), .Y(n855) );
  AOI222X1 U126 ( .A0(R12[10]), .A1(n981), .B0(R14[10]), .B1(n994), .C0(
        R13[10]), .C1(n983), .Y(n599) );
  AOI22X1 U127 ( .A0(R15[10]), .A1(n996), .B0(data_out_1[112]), .B1(n991), .Y(
        n598) );
  NAND2X1 U128 ( .A(n596), .B(n597), .Y(n854) );
  AOI222X1 U129 ( .A0(R12[11]), .A1(n981), .B0(R14[11]), .B1(n994), .C0(
        R13[11]), .C1(n983), .Y(n597) );
  AOI22X1 U130 ( .A0(R15[11]), .A1(n996), .B0(data_out_1[113]), .B1(n991), .Y(
        n596) );
  NAND2X1 U131 ( .A(n594), .B(n595), .Y(n853) );
  AOI222X1 U132 ( .A0(R12[12]), .A1(n981), .B0(R14[12]), .B1(n994), .C0(
        R13[12]), .C1(n983), .Y(n595) );
  AOI22X1 U133 ( .A0(R15[12]), .A1(n996), .B0(data_out_1[114]), .B1(n991), .Y(
        n594) );
  NAND2X1 U134 ( .A(n592), .B(n593), .Y(n852) );
  AOI222X1 U135 ( .A0(R12[13]), .A1(n981), .B0(R14[13]), .B1(n994), .C0(
        R13[13]), .C1(n983), .Y(n593) );
  AOI22X1 U136 ( .A0(R15[13]), .A1(n996), .B0(data_out_1[115]), .B1(n991), .Y(
        n592) );
  NAND2X1 U137 ( .A(n590), .B(n591), .Y(n851) );
  AOI222X1 U138 ( .A0(R12[14]), .A1(n981), .B0(R14[14]), .B1(n994), .C0(
        R13[14]), .C1(n983), .Y(n591) );
  AOI22X1 U139 ( .A0(R15[14]), .A1(n996), .B0(data_out_1[116]), .B1(n991), .Y(
        n590) );
  NAND2X1 U140 ( .A(n588), .B(n589), .Y(n850) );
  AOI222X1 U141 ( .A0(R12[15]), .A1(n981), .B0(R14[15]), .B1(n994), .C0(
        R13[15]), .C1(n983), .Y(n589) );
  AOI22X1 U142 ( .A0(R15[15]), .A1(n996), .B0(data_out_1[117]), .B1(n991), .Y(
        n588) );
  NAND2X1 U143 ( .A(n586), .B(n587), .Y(n849) );
  AOI222X1 U144 ( .A0(R12[16]), .A1(n981), .B0(R14[16]), .B1(n994), .C0(
        R13[16]), .C1(n983), .Y(n587) );
  NAND2X1 U145 ( .A(n584), .B(n585), .Y(n848) );
  AOI222X1 U146 ( .A0(R12[17]), .A1(n981), .B0(R14[17]), .B1(n994), .C0(
        R13[17]), .C1(n983), .Y(n585) );
  NAND2X1 U147 ( .A(n582), .B(n583), .Y(n847) );
  AOI222X1 U148 ( .A0(R12[18]), .A1(n981), .B0(R14[18]), .B1(n994), .C0(
        R13[18]), .C1(n983), .Y(n583) );
  NAND2X1 U149 ( .A(n580), .B(n581), .Y(n846) );
  AOI222X1 U150 ( .A0(R12[19]), .A1(n981), .B0(R14[19]), .B1(n994), .C0(
        R13[19]), .C1(n983), .Y(n581) );
  NAND2X1 U151 ( .A(n578), .B(n579), .Y(n845) );
  AOI222X1 U152 ( .A0(R12[20]), .A1(n981), .B0(R14[20]), .B1(n994), .C0(
        R13[20]), .C1(n983), .Y(n579) );
  NAND2X1 U153 ( .A(n576), .B(n577), .Y(n844) );
  AOI222X1 U154 ( .A0(R12[21]), .A1(n981), .B0(R14[21]), .B1(n994), .C0(
        R13[21]), .C1(n983), .Y(n577) );
  NAND2X1 U155 ( .A(n574), .B(n575), .Y(n843) );
  AOI222X1 U156 ( .A0(R12[22]), .A1(n981), .B0(R14[22]), .B1(n994), .C0(
        R13[22]), .C1(n983), .Y(n575) );
  NAND2X1 U157 ( .A(n572), .B(n573), .Y(n842) );
  AOI222X1 U158 ( .A0(R12[23]), .A1(n981), .B0(R14[23]), .B1(n994), .C0(
        R13[23]), .C1(n983), .Y(n573) );
  NAND2X1 U159 ( .A(n570), .B(n571), .Y(n841) );
  AOI222X1 U160 ( .A0(R12[24]), .A1(n981), .B0(R14[24]), .B1(n994), .C0(
        R13[24]), .C1(n983), .Y(n571) );
  AOI22X1 U161 ( .A0(R15[24]), .A1(n995), .B0(data_out_1[126]), .B1(n992), .Y(
        n570) );
  NAND2X1 U162 ( .A(n568), .B(n569), .Y(n840) );
  AOI222X1 U163 ( .A0(R12[25]), .A1(n981), .B0(R14[25]), .B1(n994), .C0(
        R13[25]), .C1(n983), .Y(n569) );
  AOI22X1 U164 ( .A0(R15[25]), .A1(n995), .B0(data_out_1[127]), .B1(n992), .Y(
        n568) );
  NAND2X1 U165 ( .A(n566), .B(n567), .Y(n839) );
  AOI222X1 U166 ( .A0(R12[26]), .A1(n981), .B0(R14[26]), .B1(n994), .C0(
        R13[26]), .C1(n983), .Y(n567) );
  AOI22X1 U167 ( .A0(R15[26]), .A1(n995), .B0(data_out_1[128]), .B1(n992), .Y(
        n566) );
  NAND2X1 U168 ( .A(n564), .B(n565), .Y(n838) );
  AOI222X1 U169 ( .A0(R12[27]), .A1(n981), .B0(R14[27]), .B1(n994), .C0(
        R13[27]), .C1(n983), .Y(n565) );
  AOI22X1 U170 ( .A0(R15[27]), .A1(n995), .B0(data_out_1[129]), .B1(n992), .Y(
        n564) );
  NAND2X1 U171 ( .A(n562), .B(n563), .Y(n837) );
  AOI222X1 U172 ( .A0(R12[28]), .A1(n981), .B0(R14[28]), .B1(n994), .C0(
        R13[28]), .C1(n983), .Y(n563) );
  AOI22X1 U173 ( .A0(R15[28]), .A1(n995), .B0(data_out_1[130]), .B1(n992), .Y(
        n562) );
  NAND2X1 U174 ( .A(n560), .B(n561), .Y(n836) );
  AOI222X1 U175 ( .A0(R12[29]), .A1(n981), .B0(R14[29]), .B1(n994), .C0(
        R13[29]), .C1(n983), .Y(n561) );
  AOI22X1 U176 ( .A0(R15[29]), .A1(n995), .B0(data_out_1[131]), .B1(n992), .Y(
        n560) );
  NAND2X1 U177 ( .A(n558), .B(n559), .Y(n835) );
  AOI222X1 U178 ( .A0(R12[30]), .A1(n981), .B0(R14[30]), .B1(n994), .C0(
        R13[30]), .C1(n983), .Y(n559) );
  AOI22X1 U179 ( .A0(R15[30]), .A1(n995), .B0(data_out_1[132]), .B1(n992), .Y(
        n558) );
  NAND2X1 U180 ( .A(n556), .B(n557), .Y(n834) );
  AOI222X1 U181 ( .A0(R12[31]), .A1(n981), .B0(R14[31]), .B1(n994), .C0(
        R13[31]), .C1(n983), .Y(n557) );
  AOI22X1 U182 ( .A0(R15[31]), .A1(n995), .B0(data_out_1[133]), .B1(n991), .Y(
        n556) );
  NAND2X1 U183 ( .A(n554), .B(n555), .Y(n833) );
  AOI222X1 U184 ( .A0(R12[32]), .A1(n981), .B0(R14[32]), .B1(n994), .C0(
        R13[32]), .C1(n983), .Y(n555) );
  AOI22X1 U185 ( .A0(R15[32]), .A1(n995), .B0(data_out_1[134]), .B1(n986), .Y(
        n554) );
  NAND2X1 U186 ( .A(n551), .B(n552), .Y(n832) );
  AOI222X1 U187 ( .A0(R12[33]), .A1(n981), .B0(R14[33]), .B1(n994), .C0(
        R13[33]), .C1(n983), .Y(n552) );
  NAND2X1 U188 ( .A(n686), .B(n687), .Y(n899) );
  AOI222X1 U189 ( .A0(R8[0]), .A1(n981), .B0(R10[0]), .B1(n994), .C0(R9[0]), 
        .C1(n983), .Y(n687) );
  NAND2X1 U190 ( .A(n684), .B(n685), .Y(n898) );
  AOI222X1 U191 ( .A0(R8[1]), .A1(n980), .B0(R10[1]), .B1(n993), .C0(R9[1]), 
        .C1(n983), .Y(n685) );
  NAND2X1 U192 ( .A(n682), .B(n683), .Y(n897) );
  AOI222X1 U193 ( .A0(R8[2]), .A1(n980), .B0(R10[2]), .B1(n993), .C0(R9[2]), 
        .C1(n983), .Y(n683) );
  NAND2X1 U194 ( .A(n680), .B(n681), .Y(n896) );
  AOI222X1 U195 ( .A0(R8[3]), .A1(n981), .B0(R10[3]), .B1(n994), .C0(R9[3]), 
        .C1(n983), .Y(n681) );
  NAND2X1 U196 ( .A(n678), .B(n679), .Y(n895) );
  AOI222X1 U197 ( .A0(R8[4]), .A1(n981), .B0(R10[4]), .B1(n994), .C0(R9[4]), 
        .C1(n983), .Y(n679) );
  NAND2X1 U198 ( .A(n676), .B(n677), .Y(n894) );
  AOI222X1 U199 ( .A0(R8[5]), .A1(n981), .B0(R10[5]), .B1(n994), .C0(R9[5]), 
        .C1(n983), .Y(n677) );
  NAND2X1 U200 ( .A(n674), .B(n675), .Y(n893) );
  AOI222X1 U201 ( .A0(R8[6]), .A1(n981), .B0(R10[6]), .B1(n994), .C0(R9[6]), 
        .C1(n983), .Y(n675) );
  NAND2X1 U202 ( .A(n672), .B(n673), .Y(n892) );
  AOI222X1 U203 ( .A0(R8[7]), .A1(n981), .B0(R10[7]), .B1(n994), .C0(R9[7]), 
        .C1(n983), .Y(n673) );
  AOI22X1 U204 ( .A0(R11[7]), .A1(n998), .B0(data_out_1[75]), .B1(n987), .Y(
        n672) );
  NAND2X1 U205 ( .A(n670), .B(n671), .Y(n891) );
  AOI222X1 U206 ( .A0(R8[8]), .A1(n981), .B0(R10[8]), .B1(n994), .C0(R9[8]), 
        .C1(n983), .Y(n671) );
  AOI22X1 U207 ( .A0(R11[8]), .A1(n997), .B0(data_out_1[76]), .B1(n984), .Y(
        n670) );
  NAND2X1 U208 ( .A(n668), .B(n669), .Y(n890) );
  AOI222X1 U209 ( .A0(R8[9]), .A1(n981), .B0(R10[9]), .B1(n994), .C0(R9[9]), 
        .C1(n983), .Y(n669) );
  AOI22X1 U210 ( .A0(R11[9]), .A1(n1000), .B0(data_out_1[77]), .B1(n984), .Y(
        n668) );
  NAND2X1 U211 ( .A(n666), .B(n667), .Y(n889) );
  AOI222X1 U212 ( .A0(R8[10]), .A1(n981), .B0(R10[10]), .B1(n994), .C0(R9[10]), 
        .C1(n983), .Y(n667) );
  AOI22X1 U213 ( .A0(R11[10]), .A1(n1001), .B0(data_out_1[78]), .B1(n985), .Y(
        n666) );
  NAND2X1 U214 ( .A(n664), .B(n665), .Y(n888) );
  AOI222X1 U215 ( .A0(R8[11]), .A1(n981), .B0(R10[11]), .B1(n994), .C0(R9[11]), 
        .C1(n983), .Y(n665) );
  AOI22X1 U216 ( .A0(R11[11]), .A1(n996), .B0(data_out_1[79]), .B1(n992), .Y(
        n664) );
  NAND2X1 U217 ( .A(n662), .B(n663), .Y(n887) );
  AOI222X1 U218 ( .A0(R8[12]), .A1(n981), .B0(R10[12]), .B1(n994), .C0(R9[12]), 
        .C1(n983), .Y(n663) );
  AOI22X1 U219 ( .A0(R11[12]), .A1(n999), .B0(data_out_1[80]), .B1(n989), .Y(
        n662) );
  NAND2X1 U220 ( .A(n660), .B(n661), .Y(n886) );
  AOI222X1 U221 ( .A0(R8[13]), .A1(n981), .B0(R10[13]), .B1(n994), .C0(R9[13]), 
        .C1(n983), .Y(n661) );
  AOI22X1 U222 ( .A0(R11[13]), .A1(n998), .B0(data_out_1[81]), .B1(n986), .Y(
        n660) );
  NAND2X1 U223 ( .A(n658), .B(n659), .Y(n885) );
  AOI222X1 U224 ( .A0(R8[14]), .A1(n981), .B0(R10[14]), .B1(n994), .C0(R9[14]), 
        .C1(n983), .Y(n659) );
  AOI22X1 U225 ( .A0(R11[14]), .A1(n997), .B0(data_out_1[82]), .B1(n988), .Y(
        n658) );
  NAND2X1 U226 ( .A(n656), .B(n657), .Y(n884) );
  AOI222X1 U227 ( .A0(R8[15]), .A1(n981), .B0(R10[15]), .B1(n994), .C0(R9[15]), 
        .C1(n983), .Y(n657) );
  AOI22X1 U228 ( .A0(R11[15]), .A1(n1000), .B0(data_out_1[83]), .B1(n991), .Y(
        n656) );
  NAND2X1 U229 ( .A(n654), .B(n655), .Y(n883) );
  AOI222X1 U230 ( .A0(R8[16]), .A1(n981), .B0(R10[16]), .B1(n994), .C0(R9[16]), 
        .C1(n983), .Y(n655) );
  AOI22XL U231 ( .A0(R11[16]), .A1(n997), .B0(data_out_1[84]), .B1(n989), .Y(
        n654) );
  NAND2X1 U232 ( .A(n652), .B(n653), .Y(n882) );
  AOI222X1 U233 ( .A0(R8[17]), .A1(n981), .B0(R10[17]), .B1(n994), .C0(R9[17]), 
        .C1(n983), .Y(n653) );
  NAND2X1 U234 ( .A(n650), .B(n651), .Y(n881) );
  AOI222X1 U235 ( .A0(R8[18]), .A1(n981), .B0(R10[18]), .B1(n994), .C0(R9[18]), 
        .C1(n983), .Y(n651) );
  NAND2X1 U236 ( .A(n648), .B(n649), .Y(n880) );
  AOI222X1 U237 ( .A0(R8[19]), .A1(n981), .B0(R10[19]), .B1(n994), .C0(R9[19]), 
        .C1(n983), .Y(n649) );
  NAND2X1 U238 ( .A(n646), .B(n647), .Y(n879) );
  AOI222X1 U239 ( .A0(R8[20]), .A1(n981), .B0(R10[20]), .B1(n994), .C0(R9[20]), 
        .C1(n983), .Y(n647) );
  NAND2X1 U240 ( .A(n644), .B(n645), .Y(n878) );
  AOI222X1 U241 ( .A0(R8[21]), .A1(n981), .B0(R10[21]), .B1(n994), .C0(R9[21]), 
        .C1(n983), .Y(n645) );
  NAND2X1 U242 ( .A(n642), .B(n643), .Y(n877) );
  AOI222X1 U243 ( .A0(R8[22]), .A1(n981), .B0(R10[22]), .B1(n994), .C0(R9[22]), 
        .C1(n983), .Y(n643) );
  NAND2X1 U244 ( .A(n640), .B(n641), .Y(n876) );
  AOI222X1 U245 ( .A0(R8[23]), .A1(n981), .B0(R10[23]), .B1(n994), .C0(R9[23]), 
        .C1(n983), .Y(n641) );
  NAND2X1 U246 ( .A(n638), .B(n639), .Y(n875) );
  AOI222X1 U247 ( .A0(R8[24]), .A1(n981), .B0(R10[24]), .B1(n994), .C0(R9[24]), 
        .C1(n983), .Y(n639) );
  AOI22X1 U248 ( .A0(R11[24]), .A1(n1000), .B0(data_out_1[92]), .B1(n989), .Y(
        n638) );
  NAND2X1 U249 ( .A(n636), .B(n637), .Y(n874) );
  AOI222X1 U250 ( .A0(R8[25]), .A1(n981), .B0(R10[25]), .B1(n994), .C0(R9[25]), 
        .C1(n983), .Y(n637) );
  AOI22X1 U251 ( .A0(R11[25]), .A1(n1001), .B0(data_out_1[93]), .B1(n989), .Y(
        n636) );
  NAND2X1 U252 ( .A(n634), .B(n635), .Y(n873) );
  AOI222X1 U253 ( .A0(R8[26]), .A1(n981), .B0(R10[26]), .B1(n994), .C0(R9[26]), 
        .C1(n983), .Y(n635) );
  AOI22X1 U254 ( .A0(R11[26]), .A1(n996), .B0(data_out_1[94]), .B1(n989), .Y(
        n634) );
  NAND2X1 U255 ( .A(n632), .B(n633), .Y(n872) );
  AOI222X1 U256 ( .A0(R8[27]), .A1(n981), .B0(R10[27]), .B1(n994), .C0(R9[27]), 
        .C1(n983), .Y(n633) );
  AOI22X1 U257 ( .A0(R11[27]), .A1(n999), .B0(data_out_1[95]), .B1(n989), .Y(
        n632) );
  NAND2X1 U258 ( .A(n630), .B(n631), .Y(n871) );
  AOI222X1 U259 ( .A0(R8[28]), .A1(n981), .B0(R10[28]), .B1(n994), .C0(R9[28]), 
        .C1(n983), .Y(n631) );
  AOI22X1 U260 ( .A0(R11[28]), .A1(n998), .B0(data_out_1[96]), .B1(n990), .Y(
        n630) );
  NAND2X1 U261 ( .A(n628), .B(n629), .Y(n870) );
  AOI222X1 U262 ( .A0(R8[29]), .A1(n981), .B0(R10[29]), .B1(n994), .C0(R9[29]), 
        .C1(n983), .Y(n629) );
  AOI22X1 U263 ( .A0(R11[29]), .A1(n997), .B0(data_out_1[97]), .B1(n990), .Y(
        n628) );
  NAND2X1 U264 ( .A(n626), .B(n627), .Y(n869) );
  AOI222X1 U265 ( .A0(R8[30]), .A1(n981), .B0(R10[30]), .B1(n994), .C0(R9[30]), 
        .C1(n983), .Y(n627) );
  AOI22X1 U266 ( .A0(R11[30]), .A1(n997), .B0(data_out_1[98]), .B1(n990), .Y(
        n626) );
  NAND2X1 U267 ( .A(n624), .B(n625), .Y(n868) );
  AOI222X1 U268 ( .A0(R8[31]), .A1(n981), .B0(R10[31]), .B1(n994), .C0(R9[31]), 
        .C1(n983), .Y(n625) );
  AOI22X1 U269 ( .A0(R11[31]), .A1(n997), .B0(data_out_1[99]), .B1(n990), .Y(
        n624) );
  NAND2X1 U270 ( .A(n622), .B(n623), .Y(n867) );
  AOI222X1 U271 ( .A0(R8[32]), .A1(n981), .B0(R10[32]), .B1(n994), .C0(R9[32]), 
        .C1(n983), .Y(n623) );
  AOI22X1 U272 ( .A0(R11[32]), .A1(n997), .B0(data_out_1[100]), .B1(n990), .Y(
        n622) );
  NAND2X1 U273 ( .A(n620), .B(n621), .Y(n866) );
  AOI222X1 U274 ( .A0(R8[33]), .A1(n981), .B0(R10[33]), .B1(n994), .C0(R9[33]), 
        .C1(n983), .Y(n621) );
  NAND2X1 U275 ( .A(n688), .B(n689), .Y(n900) );
  AOI222X1 U276 ( .A0(R4[33]), .A1(n981), .B0(R6[33]), .B1(n994), .C0(R5[33]), 
        .C1(n983), .Y(n689) );
  NAND2X1 U277 ( .A(n822), .B(n823), .Y(n967) );
  AOI222X1 U278 ( .A0(R0[0]), .A1(n980), .B0(R2[0]), .B1(n993), .C0(R1[0]), 
        .C1(n983), .Y(n823) );
  AOI22X1 U279 ( .A0(R3[0]), .A1(n1002), .B0(data_out_1[0]), .B1(n984), .Y(
        n822) );
  NAND2X1 U280 ( .A(n754), .B(n755), .Y(n933) );
  AOI222X1 U281 ( .A0(R4[0]), .A1(n981), .B0(R6[0]), .B1(n994), .C0(R5[0]), 
        .C1(n983), .Y(n755) );
  NAND2X1 U282 ( .A(n752), .B(n753), .Y(n932) );
  AOI222X1 U283 ( .A0(R4[1]), .A1(n981), .B0(R6[1]), .B1(n994), .C0(R5[1]), 
        .C1(n983), .Y(n753) );
  NAND2X1 U284 ( .A(n750), .B(n751), .Y(n931) );
  AOI222X1 U285 ( .A0(R4[2]), .A1(n981), .B0(R6[2]), .B1(n994), .C0(R5[2]), 
        .C1(n983), .Y(n751) );
  NAND2X1 U286 ( .A(n748), .B(n749), .Y(n930) );
  AOI222X1 U287 ( .A0(R4[3]), .A1(n981), .B0(R6[3]), .B1(n994), .C0(R5[3]), 
        .C1(n983), .Y(n749) );
  NAND2X1 U288 ( .A(n746), .B(n747), .Y(n929) );
  AOI222X1 U289 ( .A0(R4[4]), .A1(n981), .B0(R6[4]), .B1(n994), .C0(R5[4]), 
        .C1(n983), .Y(n747) );
  NAND2X1 U290 ( .A(n744), .B(n745), .Y(n928) );
  AOI222X1 U291 ( .A0(R4[5]), .A1(n981), .B0(R6[5]), .B1(n994), .C0(R5[5]), 
        .C1(n983), .Y(n745) );
  NAND2X1 U292 ( .A(n742), .B(n743), .Y(n927) );
  AOI222X1 U293 ( .A0(R4[6]), .A1(n981), .B0(R6[6]), .B1(n994), .C0(R5[6]), 
        .C1(n983), .Y(n743) );
  NAND2X1 U294 ( .A(n740), .B(n741), .Y(n926) );
  AOI222X1 U295 ( .A0(R4[7]), .A1(n981), .B0(R6[7]), .B1(n994), .C0(R5[7]), 
        .C1(n983), .Y(n741) );
  AOI22X1 U296 ( .A0(R7[7]), .A1(n999), .B0(data_out_1[41]), .B1(n987), .Y(
        n740) );
  NAND2X1 U297 ( .A(n738), .B(n739), .Y(n925) );
  AOI222X1 U298 ( .A0(R4[8]), .A1(n981), .B0(R6[8]), .B1(n994), .C0(R5[8]), 
        .C1(n983), .Y(n739) );
  AOI22X1 U299 ( .A0(R7[8]), .A1(n999), .B0(data_out_1[42]), .B1(n987), .Y(
        n738) );
  NAND2X1 U300 ( .A(n736), .B(n737), .Y(n924) );
  AOI222X1 U301 ( .A0(R4[9]), .A1(n981), .B0(R6[9]), .B1(n994), .C0(R5[9]), 
        .C1(n983), .Y(n737) );
  AOI22X1 U302 ( .A0(R7[9]), .A1(n999), .B0(data_out_1[43]), .B1(n987), .Y(
        n736) );
  NAND2X1 U303 ( .A(n734), .B(n735), .Y(n923) );
  AOI222X1 U304 ( .A0(R4[10]), .A1(n981), .B0(R6[10]), .B1(n994), .C0(R5[10]), 
        .C1(n983), .Y(n735) );
  AOI22X1 U305 ( .A0(R7[10]), .A1(n999), .B0(data_out_1[44]), .B1(n987), .Y(
        n734) );
  NAND2X1 U306 ( .A(n732), .B(n733), .Y(n922) );
  AOI222X1 U307 ( .A0(R4[11]), .A1(n981), .B0(R6[11]), .B1(n994), .C0(R5[11]), 
        .C1(n983), .Y(n733) );
  AOI22X1 U308 ( .A0(R7[11]), .A1(n999), .B0(data_out_1[45]), .B1(n987), .Y(
        n732) );
  NAND2X1 U309 ( .A(n730), .B(n731), .Y(n921) );
  AOI222X1 U310 ( .A0(R4[12]), .A1(n981), .B0(R6[12]), .B1(n994), .C0(R5[12]), 
        .C1(n983), .Y(n731) );
  AOI22X1 U311 ( .A0(R7[12]), .A1(n997), .B0(data_out_1[46]), .B1(n987), .Y(
        n730) );
  NAND2X1 U312 ( .A(n728), .B(n729), .Y(n920) );
  AOI222X1 U313 ( .A0(R4[13]), .A1(n981), .B0(R6[13]), .B1(n994), .C0(R5[13]), 
        .C1(n983), .Y(n729) );
  AOI22X1 U314 ( .A0(R7[13]), .A1(n996), .B0(data_out_1[47]), .B1(n987), .Y(
        n728) );
  NAND2X1 U315 ( .A(n726), .B(n727), .Y(n919) );
  AOI222X1 U316 ( .A0(R4[14]), .A1(n981), .B0(R6[14]), .B1(n994), .C0(R5[14]), 
        .C1(n983), .Y(n727) );
  AOI22X1 U317 ( .A0(R7[14]), .A1(n997), .B0(data_out_1[48]), .B1(n985), .Y(
        n726) );
  NAND2X1 U318 ( .A(n724), .B(n725), .Y(n918) );
  AOI222X1 U319 ( .A0(R4[15]), .A1(n981), .B0(R6[15]), .B1(n994), .C0(R5[15]), 
        .C1(n983), .Y(n725) );
  AOI22X1 U320 ( .A0(R7[15]), .A1(n996), .B0(data_out_1[49]), .B1(n984), .Y(
        n724) );
  NAND2X1 U321 ( .A(n722), .B(n723), .Y(n917) );
  AOI222X1 U322 ( .A0(R4[16]), .A1(n981), .B0(R6[16]), .B1(n994), .C0(R5[16]), 
        .C1(n983), .Y(n723) );
  NAND2X1 U323 ( .A(n720), .B(n721), .Y(n916) );
  AOI222X1 U324 ( .A0(R4[17]), .A1(n981), .B0(R6[17]), .B1(n994), .C0(R5[17]), 
        .C1(n983), .Y(n721) );
  NAND2X1 U325 ( .A(n718), .B(n719), .Y(n915) );
  AOI222X1 U326 ( .A0(R4[18]), .A1(n981), .B0(R6[18]), .B1(n994), .C0(R5[18]), 
        .C1(n983), .Y(n719) );
  NAND2X1 U327 ( .A(n716), .B(n717), .Y(n914) );
  AOI222X1 U328 ( .A0(R4[19]), .A1(n981), .B0(R6[19]), .B1(n994), .C0(R5[19]), 
        .C1(n983), .Y(n717) );
  NAND2X1 U329 ( .A(n714), .B(n715), .Y(n913) );
  AOI222X1 U330 ( .A0(R4[20]), .A1(n981), .B0(R6[20]), .B1(n994), .C0(R5[20]), 
        .C1(n983), .Y(n715) );
  NAND2X1 U331 ( .A(n712), .B(n713), .Y(n912) );
  AOI222X1 U332 ( .A0(R4[21]), .A1(n981), .B0(R6[21]), .B1(n994), .C0(R5[21]), 
        .C1(n983), .Y(n713) );
  NAND2X1 U333 ( .A(n710), .B(n711), .Y(n911) );
  AOI222X1 U334 ( .A0(R4[22]), .A1(n981), .B0(R6[22]), .B1(n994), .C0(R5[22]), 
        .C1(n983), .Y(n711) );
  NAND2X1 U335 ( .A(n708), .B(n709), .Y(n910) );
  AOI222X1 U336 ( .A0(R4[23]), .A1(n981), .B0(R6[23]), .B1(n994), .C0(R5[23]), 
        .C1(n983), .Y(n709) );
  NAND2X1 U337 ( .A(n706), .B(n707), .Y(n909) );
  AOI222X1 U338 ( .A0(R4[24]), .A1(n981), .B0(R6[24]), .B1(n994), .C0(R5[24]), 
        .C1(n983), .Y(n707) );
  AOI22X1 U339 ( .A0(R7[24]), .A1(n998), .B0(data_out_1[58]), .B1(n985), .Y(
        n706) );
  NAND2X1 U340 ( .A(n704), .B(n705), .Y(n908) );
  AOI222X1 U341 ( .A0(R4[25]), .A1(n981), .B0(R6[25]), .B1(n994), .C0(R5[25]), 
        .C1(n983), .Y(n705) );
  AOI22X1 U342 ( .A0(R7[25]), .A1(n998), .B0(data_out_1[59]), .B1(n987), .Y(
        n704) );
  NAND2X1 U343 ( .A(n702), .B(n703), .Y(n907) );
  AOI222X1 U344 ( .A0(R4[26]), .A1(n981), .B0(R6[26]), .B1(n994), .C0(R5[26]), 
        .C1(n983), .Y(n703) );
  AOI22X1 U345 ( .A0(R7[26]), .A1(n998), .B0(data_out_1[60]), .B1(n988), .Y(
        n702) );
  NAND2X1 U346 ( .A(n700), .B(n701), .Y(n906) );
  AOI222X1 U347 ( .A0(R4[27]), .A1(n981), .B0(R6[27]), .B1(n994), .C0(R5[27]), 
        .C1(n983), .Y(n701) );
  AOI22X1 U348 ( .A0(R7[27]), .A1(n998), .B0(data_out_1[61]), .B1(n988), .Y(
        n700) );
  NAND2X1 U349 ( .A(n698), .B(n699), .Y(n905) );
  AOI222X1 U350 ( .A0(R4[28]), .A1(n981), .B0(R6[28]), .B1(n994), .C0(R5[28]), 
        .C1(n983), .Y(n699) );
  AOI22X1 U351 ( .A0(R7[28]), .A1(n998), .B0(data_out_1[62]), .B1(n988), .Y(
        n698) );
  NAND2X1 U352 ( .A(n696), .B(n697), .Y(n904) );
  AOI222X1 U353 ( .A0(R4[29]), .A1(n981), .B0(R6[29]), .B1(n994), .C0(R5[29]), 
        .C1(n983), .Y(n697) );
  AOI22X1 U354 ( .A0(R7[29]), .A1(n998), .B0(data_out_1[63]), .B1(n988), .Y(
        n696) );
  NAND2X1 U355 ( .A(n694), .B(n695), .Y(n903) );
  AOI222X1 U356 ( .A0(R4[30]), .A1(n981), .B0(R6[30]), .B1(n994), .C0(R5[30]), 
        .C1(n983), .Y(n695) );
  AOI22X1 U357 ( .A0(R7[30]), .A1(n998), .B0(data_out_1[64]), .B1(n988), .Y(
        n694) );
  NAND2X1 U358 ( .A(n692), .B(n693), .Y(n902) );
  AOI222X1 U359 ( .A0(R4[31]), .A1(n981), .B0(R6[31]), .B1(n994), .C0(R5[31]), 
        .C1(n983), .Y(n693) );
  AOI22X1 U360 ( .A0(R7[31]), .A1(n998), .B0(data_out_1[65]), .B1(n988), .Y(
        n692) );
  NAND2X1 U361 ( .A(n690), .B(n691), .Y(n901) );
  AOI222X1 U362 ( .A0(R4[32]), .A1(n981), .B0(R6[32]), .B1(n994), .C0(R5[32]), 
        .C1(n983), .Y(n691) );
  AOI22X1 U363 ( .A0(R7[32]), .A1(n998), .B0(data_out_1[66]), .B1(n988), .Y(
        n690) );
  NAND2X1 U364 ( .A(n820), .B(n821), .Y(n966) );
  AOI222X1 U365 ( .A0(R0[1]), .A1(n981), .B0(R2[1]), .B1(n994), .C0(R1[1]), 
        .C1(n983), .Y(n821) );
  AOI22X1 U366 ( .A0(R3[1]), .A1(n1002), .B0(data_out_1[1]), .B1(n984), .Y(
        n820) );
  NAND2X1 U367 ( .A(n818), .B(n819), .Y(n965) );
  AOI222X1 U368 ( .A0(R0[2]), .A1(n981), .B0(R2[2]), .B1(n994), .C0(R1[2]), 
        .C1(n982), .Y(n819) );
  AOI22X1 U369 ( .A0(R3[2]), .A1(n1002), .B0(data_out_1[2]), .B1(n984), .Y(
        n818) );
  NAND2X1 U370 ( .A(n816), .B(n817), .Y(n964) );
  AOI222X1 U371 ( .A0(R0[3]), .A1(n981), .B0(R2[3]), .B1(n994), .C0(R1[3]), 
        .C1(n983), .Y(n817) );
  AOI22X1 U372 ( .A0(R3[3]), .A1(n1002), .B0(data_out_1[3]), .B1(n984), .Y(
        n816) );
  NAND2X1 U373 ( .A(n814), .B(n815), .Y(n963) );
  AOI222X1 U374 ( .A0(R0[4]), .A1(n981), .B0(R2[4]), .B1(n994), .C0(R1[4]), 
        .C1(n983), .Y(n815) );
  AOI22X1 U375 ( .A0(R3[4]), .A1(n1002), .B0(data_out_1[4]), .B1(n984), .Y(
        n814) );
  NAND2X1 U376 ( .A(n812), .B(n813), .Y(n962) );
  AOI222X1 U377 ( .A0(R0[5]), .A1(n981), .B0(R2[5]), .B1(n994), .C0(R1[5]), 
        .C1(n983), .Y(n813) );
  AOI22X1 U378 ( .A0(R3[5]), .A1(n1002), .B0(data_out_1[5]), .B1(n984), .Y(
        n812) );
  NAND2X1 U379 ( .A(n810), .B(n811), .Y(n961) );
  AOI222X1 U380 ( .A0(R0[6]), .A1(n981), .B0(R2[6]), .B1(n994), .C0(R1[6]), 
        .C1(n983), .Y(n811) );
  AOI22X1 U381 ( .A0(R3[6]), .A1(n1002), .B0(data_out_1[6]), .B1(n984), .Y(
        n810) );
  NAND2X1 U382 ( .A(n808), .B(n809), .Y(n960) );
  AOI222X1 U383 ( .A0(R0[7]), .A1(n981), .B0(R2[7]), .B1(n994), .C0(R1[7]), 
        .C1(n983), .Y(n809) );
  AOI22X1 U384 ( .A0(R3[7]), .A1(n1001), .B0(data_out_1[7]), .B1(n984), .Y(
        n808) );
  NAND2X1 U385 ( .A(n806), .B(n807), .Y(n959) );
  AOI222X1 U386 ( .A0(R0[8]), .A1(n981), .B0(R2[8]), .B1(n994), .C0(R1[8]), 
        .C1(n983), .Y(n807) );
  AOI22X1 U387 ( .A0(R3[8]), .A1(n1001), .B0(data_out_1[8]), .B1(n984), .Y(
        n806) );
  NAND2X1 U388 ( .A(n804), .B(n805), .Y(n958) );
  AOI222X1 U389 ( .A0(R0[9]), .A1(n981), .B0(R2[9]), .B1(n994), .C0(R1[9]), 
        .C1(n983), .Y(n805) );
  AOI22X1 U390 ( .A0(R3[9]), .A1(n1001), .B0(data_out_1[9]), .B1(n984), .Y(
        n804) );
  NAND2X1 U391 ( .A(n802), .B(n803), .Y(n957) );
  AOI222X1 U392 ( .A0(R0[10]), .A1(n981), .B0(R2[10]), .B1(n994), .C0(R1[10]), 
        .C1(n983), .Y(n803) );
  AOI22X1 U393 ( .A0(R3[10]), .A1(n1001), .B0(data_out_1[10]), .B1(n984), .Y(
        n802) );
  NAND2X1 U394 ( .A(n800), .B(n801), .Y(n956) );
  AOI222X1 U395 ( .A0(R0[11]), .A1(n981), .B0(R2[11]), .B1(n994), .C0(R1[11]), 
        .C1(n983), .Y(n801) );
  AOI22X1 U396 ( .A0(R3[11]), .A1(n1001), .B0(data_out_1[11]), .B1(n984), .Y(
        n800) );
  NAND2X1 U397 ( .A(n798), .B(n799), .Y(n955) );
  AOI222X1 U398 ( .A0(R0[12]), .A1(n981), .B0(R2[12]), .B1(n994), .C0(R1[12]), 
        .C1(n983), .Y(n799) );
  AOI22X1 U399 ( .A0(R3[12]), .A1(n1001), .B0(data_out_1[12]), .B1(n985), .Y(
        n798) );
  NAND2X1 U400 ( .A(n796), .B(n797), .Y(n954) );
  AOI222X1 U401 ( .A0(R0[13]), .A1(n981), .B0(R2[13]), .B1(n994), .C0(R1[13]), 
        .C1(n983), .Y(n797) );
  AOI22X1 U402 ( .A0(R3[13]), .A1(n1001), .B0(data_out_1[13]), .B1(n985), .Y(
        n796) );
  NAND2X1 U403 ( .A(n794), .B(n795), .Y(n953) );
  AOI222X1 U404 ( .A0(R0[14]), .A1(n981), .B0(R2[14]), .B1(n994), .C0(R1[14]), 
        .C1(n983), .Y(n795) );
  AOI22X1 U405 ( .A0(R3[14]), .A1(n1001), .B0(data_out_1[14]), .B1(n985), .Y(
        n794) );
  NAND2X1 U406 ( .A(n792), .B(n793), .Y(n952) );
  AOI222X1 U407 ( .A0(R0[15]), .A1(n981), .B0(R2[15]), .B1(n994), .C0(R1[15]), 
        .C1(n983), .Y(n793) );
  AOI22X1 U408 ( .A0(R3[15]), .A1(n1001), .B0(data_out_1[15]), .B1(n985), .Y(
        n792) );
  NAND2X1 U409 ( .A(n790), .B(n791), .Y(n951) );
  AOI222X1 U410 ( .A0(R0[16]), .A1(n981), .B0(R2[16]), .B1(n994), .C0(R1[16]), 
        .C1(n983), .Y(n791) );
  AOI22X1 U411 ( .A0(R3[16]), .A1(n1001), .B0(data_out_1[16]), .B1(n985), .Y(
        n790) );
  NAND2X1 U412 ( .A(n788), .B(n789), .Y(n950) );
  AOI222X1 U413 ( .A0(R0[17]), .A1(n981), .B0(R2[17]), .B1(n994), .C0(R1[17]), 
        .C1(n983), .Y(n789) );
  AOI22X1 U414 ( .A0(R3[17]), .A1(n1001), .B0(data_out_1[17]), .B1(n985), .Y(
        n788) );
  NAND2X1 U415 ( .A(n786), .B(n787), .Y(n949) );
  AOI222X1 U416 ( .A0(R0[18]), .A1(n981), .B0(R2[18]), .B1(n994), .C0(R1[18]), 
        .C1(n983), .Y(n787) );
  AOI22X1 U417 ( .A0(R3[18]), .A1(n1001), .B0(data_out_1[18]), .B1(n985), .Y(
        n786) );
  NAND2X1 U418 ( .A(n784), .B(n785), .Y(n948) );
  AOI222X1 U419 ( .A0(R0[19]), .A1(n981), .B0(R2[19]), .B1(n994), .C0(R1[19]), 
        .C1(n983), .Y(n785) );
  AOI22X1 U420 ( .A0(R3[19]), .A1(n1001), .B0(data_out_1[19]), .B1(n985), .Y(
        n784) );
  NAND2X1 U421 ( .A(n782), .B(n783), .Y(n947) );
  AOI222X1 U422 ( .A0(R0[20]), .A1(n981), .B0(R2[20]), .B1(n994), .C0(R1[20]), 
        .C1(n983), .Y(n783) );
  AOI22X1 U423 ( .A0(R3[20]), .A1(n1000), .B0(data_out_1[20]), .B1(n985), .Y(
        n782) );
  NAND2X1 U424 ( .A(n780), .B(n781), .Y(n946) );
  AOI222X1 U425 ( .A0(R0[21]), .A1(n981), .B0(R2[21]), .B1(n994), .C0(R1[21]), 
        .C1(n983), .Y(n781) );
  AOI22X1 U426 ( .A0(R3[21]), .A1(n1000), .B0(data_out_1[21]), .B1(n985), .Y(
        n780) );
  NAND2X1 U427 ( .A(n778), .B(n779), .Y(n945) );
  AOI222X1 U428 ( .A0(R0[22]), .A1(n981), .B0(R2[22]), .B1(n994), .C0(R1[22]), 
        .C1(n983), .Y(n779) );
  AOI22X1 U429 ( .A0(R3[22]), .A1(n1000), .B0(data_out_1[22]), .B1(n985), .Y(
        n778) );
  NAND2X1 U430 ( .A(n776), .B(n777), .Y(n944) );
  AOI222X1 U431 ( .A0(R0[23]), .A1(n981), .B0(R2[23]), .B1(n994), .C0(R1[23]), 
        .C1(n983), .Y(n777) );
  AOI22X1 U432 ( .A0(R3[23]), .A1(n1000), .B0(data_out_1[23]), .B1(n985), .Y(
        n776) );
  NAND2X1 U433 ( .A(n774), .B(n775), .Y(n943) );
  AOI222X1 U434 ( .A0(R0[24]), .A1(n981), .B0(R2[24]), .B1(n994), .C0(R1[24]), 
        .C1(n983), .Y(n775) );
  AOI22X1 U435 ( .A0(R3[24]), .A1(n1000), .B0(data_out_1[24]), .B1(n986), .Y(
        n774) );
  NAND2X1 U436 ( .A(n772), .B(n773), .Y(n942) );
  AOI222X1 U437 ( .A0(R0[25]), .A1(n981), .B0(R2[25]), .B1(n994), .C0(R1[25]), 
        .C1(n983), .Y(n773) );
  AOI22X1 U438 ( .A0(R3[25]), .A1(n1000), .B0(data_out_1[25]), .B1(n986), .Y(
        n772) );
  NAND2X1 U439 ( .A(n770), .B(n771), .Y(n941) );
  AOI222X1 U440 ( .A0(R0[26]), .A1(n981), .B0(R2[26]), .B1(n994), .C0(R1[26]), 
        .C1(n983), .Y(n771) );
  AOI22X1 U441 ( .A0(R3[26]), .A1(n1000), .B0(data_out_1[26]), .B1(n986), .Y(
        n770) );
  NAND2X1 U442 ( .A(n768), .B(n769), .Y(n940) );
  AOI222X1 U443 ( .A0(R0[27]), .A1(n981), .B0(R2[27]), .B1(n994), .C0(R1[27]), 
        .C1(n983), .Y(n769) );
  AOI22X1 U444 ( .A0(R3[27]), .A1(n1000), .B0(data_out_1[27]), .B1(n986), .Y(
        n768) );
  NAND2X1 U445 ( .A(n766), .B(n767), .Y(n939) );
  AOI222X1 U446 ( .A0(R0[28]), .A1(n981), .B0(R2[28]), .B1(n994), .C0(R1[28]), 
        .C1(n983), .Y(n767) );
  AOI22X1 U447 ( .A0(R3[28]), .A1(n1000), .B0(data_out_1[28]), .B1(n986), .Y(
        n766) );
  NAND2X1 U448 ( .A(n764), .B(n765), .Y(n938) );
  AOI222X1 U449 ( .A0(R0[29]), .A1(n981), .B0(R2[29]), .B1(n994), .C0(R1[29]), 
        .C1(n983), .Y(n765) );
  AOI22X1 U450 ( .A0(R3[29]), .A1(n1000), .B0(data_out_1[29]), .B1(n986), .Y(
        n764) );
  NAND2X1 U451 ( .A(n762), .B(n763), .Y(n937) );
  AOI222X1 U452 ( .A0(R0[30]), .A1(n981), .B0(R2[30]), .B1(n994), .C0(R1[30]), 
        .C1(n983), .Y(n763) );
  AOI22X1 U453 ( .A0(R3[30]), .A1(n1000), .B0(data_out_1[30]), .B1(n986), .Y(
        n762) );
  NAND2X1 U454 ( .A(n760), .B(n761), .Y(n936) );
  AOI222X1 U455 ( .A0(R0[31]), .A1(n981), .B0(R2[31]), .B1(n994), .C0(R1[31]), 
        .C1(n982), .Y(n761) );
  AOI22X1 U456 ( .A0(R3[31]), .A1(n1000), .B0(data_out_1[31]), .B1(n986), .Y(
        n760) );
  NAND2X1 U457 ( .A(n758), .B(n759), .Y(n935) );
  AOI222X1 U458 ( .A0(R0[32]), .A1(n981), .B0(R2[32]), .B1(n994), .C0(R1[32]), 
        .C1(n983), .Y(n759) );
  AOI22X1 U459 ( .A0(R3[32]), .A1(n1000), .B0(data_out_1[32]), .B1(n986), .Y(
        n758) );
  NAND2X1 U460 ( .A(n756), .B(n757), .Y(n934) );
  AOI222X1 U461 ( .A0(R0[33]), .A1(n981), .B0(R2[33]), .B1(n994), .C0(R1[33]), 
        .C1(n983), .Y(n757) );
  AOI22X1 U462 ( .A0(R3[33]), .A1(n999), .B0(data_out_1[33]), .B1(n986), .Y(
        n756) );
  NAND2X1 U463 ( .A(counter[1]), .B(n550), .Y(n824) );
  NAND2X1 U464 ( .A(counter[3]), .B(n1005), .Y(n827) );
  NAND2X1 U465 ( .A(counter[2]), .B(n1006), .Y(n829) );
  OAI22X1 U466 ( .A0(n831), .A1(n1005), .B0(counter[2]), .B1(n826), .Y(N14) );
  NOR2X1 U467 ( .A(n550), .B(n1004), .Y(n831) );
endmodule


module mux ( mux_flag, clk, rst_n, data_in_1, data_in_2, data_out, 
        data_in_3_33_, data_in_3_32_, data_in_3_31_, data_in_3_30_, 
        data_in_3_29_, data_in_3_28_, data_in_3_27_, data_in_3_26_, 
        data_in_3_25_, data_in_3_24_, data_in_3_23_, data_in_3_22_, 
        data_in_3_21_, data_in_3_20_, data_in_3_19_, data_in_3_18_, 
        data_in_3_17_, data_in_3_16_, data_in_3_15_, data_in_3_14_, 
        data_in_3_13_, data_in_3_12_, data_in_3_11_, data_in_3_10_, 
        data_in_3_9_, data_in_3_8_, data_in_3_7_, data_in_3_6_, data_in_3_5_, 
        data_in_3_4_, data_in_3_3_, data_in_3_2_, data_in_3_1_, data_in_3_0_
 );
  input [135:0] data_in_1;
  input [135:0] data_in_2;
  output [135:0] data_out;
  input mux_flag, clk, rst_n, data_in_3_33_, data_in_3_32_, data_in_3_31_,
         data_in_3_30_, data_in_3_29_, data_in_3_28_, data_in_3_27_,
         data_in_3_26_, data_in_3_25_, data_in_3_24_, data_in_3_23_,
         data_in_3_22_, data_in_3_21_, data_in_3_20_, data_in_3_19_,
         data_in_3_18_, data_in_3_17_, data_in_3_16_, data_in_3_15_,
         data_in_3_14_, data_in_3_13_, data_in_3_12_, data_in_3_11_,
         data_in_3_10_, data_in_3_9_, data_in_3_8_, data_in_3_7_, data_in_3_6_,
         data_in_3_5_, data_in_3_4_, data_in_3_3_, data_in_3_2_, data_in_3_1_,
         data_in_3_0_;
  wire   N6, N7, N8, n140, n141, n281, n282, n285, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n242, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n283, n284, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n720;
  wire   [3:1] counter;
  wire   [33:0] R4;
  wire   [33:0] R3;
  wire   [33:0] R2;
  wire   [33:0] R1;

  JKFFRX4 counter_reg_0_ ( .J(1'b1), .K(1'b1), .CK(clk), .RN(rst_n), .QN(n140)
         );
  DFFRHQX4 counter_reg_1_ ( .D(N6), .CK(clk), .RN(rst_n), .Q(counter[1]) );
  DFFRHQX4 counter_reg_3_ ( .D(N8), .CK(clk), .RN(rst_n), .Q(counter[3]) );
  TLATXL R4_reg_33_ ( .G(n276), .D(data_in_3_33_), .Q(R4[33]) );
  TLATXL R3_reg_33_ ( .G(n82), .D(data_in_3_33_), .Q(R3[33]) );
  TLATXL R2_reg_33_ ( .G(n81), .D(data_in_3_33_), .Q(R2[33]) );
  TLATXL R1_reg_33_ ( .G(n285), .D(data_in_3_33_), .Q(R1[33]) );
  TLATXL R4_reg_14_ ( .G(n276), .D(data_in_3_14_), .Q(R4[14]) );
  TLATXL R3_reg_14_ ( .G(n82), .D(data_in_3_14_), .Q(R3[14]) );
  TLATXL R2_reg_14_ ( .G(n81), .D(data_in_3_14_), .Q(R2[14]) );
  TLATXL R1_reg_14_ ( .G(n274), .D(data_in_3_14_), .Q(R1[14]) );
  TLATXL R3_reg_16_ ( .G(n82), .D(data_in_3_16_), .Q(R3[16]) );
  TLATX1 R2_reg_1_ ( .G(n81), .D(data_in_3_1_), .Q(R2[1]) );
  TLATX1 R2_reg_0_ ( .G(n81), .D(data_in_3_0_), .Q(R2[0]) );
  TLATX1 R3_reg_2_ ( .G(n82), .D(data_in_3_2_), .Q(R3[2]) );
  TLATX1 R3_reg_0_ ( .G(n82), .D(data_in_3_0_), .Q(R3[0]) );
  TLATX1 R4_reg_0_ ( .G(n276), .D(data_in_3_0_), .Q(R4[0]) );
  TLATX1 R2_reg_17_ ( .G(n81), .D(data_in_3_17_), .Q(R2[17]) );
  TLATX1 R2_reg_19_ ( .G(n81), .D(data_in_3_19_), .Q(R2[19]) );
  TLATX1 R1_reg_5_ ( .G(n285), .D(data_in_3_5_), .Q(R1[5]) );
  TLATX1 R1_reg_4_ ( .G(n285), .D(data_in_3_4_), .Q(R1[4]) );
  TLATX1 R1_reg_3_ ( .G(n285), .D(data_in_3_3_), .Q(R1[3]) );
  TLATX1 R1_reg_2_ ( .G(n285), .D(data_in_3_2_), .Q(R1[2]) );
  TLATX1 R1_reg_1_ ( .G(n285), .D(data_in_3_1_), .Q(R1[1]) );
  TLATX1 R1_reg_0_ ( .G(n285), .D(data_in_3_0_), .Q(R1[0]) );
  TLATX1 R2_reg_5_ ( .G(n81), .D(data_in_3_5_), .Q(R2[5]) );
  TLATX1 R2_reg_4_ ( .G(n81), .D(data_in_3_4_), .Q(R2[4]) );
  TLATX1 R2_reg_3_ ( .G(n81), .D(data_in_3_3_), .Q(R2[3]) );
  TLATX1 R2_reg_2_ ( .G(n81), .D(data_in_3_2_), .Q(R2[2]) );
  TLATX1 R3_reg_5_ ( .G(n82), .D(data_in_3_5_), .Q(R3[5]) );
  TLATX1 R3_reg_4_ ( .G(n82), .D(data_in_3_4_), .Q(R3[4]) );
  TLATX1 R3_reg_3_ ( .G(n82), .D(data_in_3_3_), .Q(R3[3]) );
  TLATX1 R4_reg_5_ ( .G(n276), .D(data_in_3_5_), .Q(R4[5]) );
  TLATX1 R4_reg_4_ ( .G(n276), .D(data_in_3_4_), .Q(R4[4]) );
  TLATX1 R4_reg_3_ ( .G(n276), .D(data_in_3_3_), .Q(R4[3]) );
  TLATX1 R4_reg_1_ ( .G(n276), .D(data_in_3_1_), .Q(R4[1]) );
  TLATXL R1_reg_32_ ( .G(n274), .D(data_in_3_32_), .Q(R1[32]) );
  TLATXL R1_reg_31_ ( .G(n285), .D(data_in_3_31_), .Q(R1[31]) );
  TLATXL R1_reg_30_ ( .G(n274), .D(data_in_3_30_), .Q(R1[30]) );
  TLATXL R1_reg_29_ ( .G(n285), .D(data_in_3_29_), .Q(R1[29]) );
  TLATX1 R1_reg_22_ ( .G(n285), .D(data_in_3_22_), .Q(R1[22]) );
  TLATX1 R1_reg_21_ ( .G(n274), .D(data_in_3_21_), .Q(R1[21]) );
  TLATX1 R1_reg_20_ ( .G(n274), .D(data_in_3_20_), .Q(R1[20]) );
  TLATX1 R1_reg_19_ ( .G(n274), .D(data_in_3_19_), .Q(R1[19]) );
  TLATX1 R1_reg_18_ ( .G(n274), .D(data_in_3_18_), .Q(R1[18]) );
  TLATX1 R1_reg_17_ ( .G(n274), .D(data_in_3_17_), .Q(R1[17]) );
  TLATXL R1_reg_16_ ( .G(n274), .D(data_in_3_16_), .Q(R1[16]) );
  TLATXL R1_reg_15_ ( .G(n274), .D(data_in_3_15_), .Q(R1[15]) );
  TLATXL R1_reg_13_ ( .G(n274), .D(data_in_3_13_), .Q(n156) );
  TLATXL R1_reg_12_ ( .G(n274), .D(data_in_3_12_), .Q(R1[12]) );
  TLATXL R2_reg_32_ ( .G(n81), .D(data_in_3_32_), .Q(R2[32]) );
  TLATXL R2_reg_31_ ( .G(n81), .D(data_in_3_31_), .Q(R2[31]) );
  TLATXL R2_reg_30_ ( .G(n81), .D(data_in_3_30_), .Q(R2[30]) );
  TLATXL R2_reg_29_ ( .G(n81), .D(data_in_3_29_), .Q(R2[29]) );
  TLATX1 R2_reg_22_ ( .G(n81), .D(data_in_3_22_), .Q(R2[22]) );
  TLATX1 R2_reg_21_ ( .G(n81), .D(data_in_3_21_), .Q(R2[21]) );
  TLATX1 R2_reg_20_ ( .G(n81), .D(data_in_3_20_), .Q(R2[20]) );
  TLATX1 R2_reg_18_ ( .G(n81), .D(data_in_3_18_), .Q(R2[18]) );
  TLATXL R2_reg_16_ ( .G(n81), .D(data_in_3_16_), .Q(R2[16]) );
  TLATXL R2_reg_15_ ( .G(n81), .D(data_in_3_15_), .Q(R2[15]) );
  TLATXL R2_reg_13_ ( .G(n81), .D(data_in_3_13_), .Q(R2[13]) );
  TLATXL R2_reg_12_ ( .G(n81), .D(data_in_3_12_), .Q(R2[12]) );
  TLATXL R3_reg_32_ ( .G(n82), .D(data_in_3_32_), .Q(R3[32]) );
  TLATXL R3_reg_31_ ( .G(n82), .D(data_in_3_31_), .Q(R3[31]) );
  TLATXL R3_reg_30_ ( .G(n82), .D(data_in_3_30_), .Q(R3[30]) );
  TLATXL R3_reg_29_ ( .G(n82), .D(data_in_3_29_), .Q(R3[29]) );
  TLATX1 R3_reg_22_ ( .G(n82), .D(data_in_3_22_), .Q(R3[22]) );
  TLATX1 R3_reg_21_ ( .G(n82), .D(data_in_3_21_), .Q(R3[21]) );
  TLATX1 R3_reg_20_ ( .G(n82), .D(data_in_3_20_), .Q(R3[20]) );
  TLATX1 R3_reg_19_ ( .G(n82), .D(data_in_3_19_), .Q(R3[19]) );
  TLATX1 R3_reg_18_ ( .G(n82), .D(data_in_3_18_), .Q(R3[18]) );
  TLATX1 R3_reg_17_ ( .G(n82), .D(data_in_3_17_), .Q(R3[17]) );
  TLATXL R3_reg_15_ ( .G(n82), .D(data_in_3_15_), .Q(R3[15]) );
  TLATXL R3_reg_13_ ( .G(n82), .D(data_in_3_13_), .Q(R3[13]) );
  TLATXL R3_reg_12_ ( .G(n82), .D(data_in_3_12_), .Q(R3[12]) );
  TLATXL R4_reg_32_ ( .G(n276), .D(data_in_3_32_), .Q(R4[32]) );
  TLATXL R4_reg_31_ ( .G(n276), .D(data_in_3_31_), .Q(R4[31]) );
  TLATXL R4_reg_30_ ( .G(n276), .D(data_in_3_30_), .Q(R4[30]) );
  TLATXL R4_reg_29_ ( .G(n276), .D(data_in_3_29_), .Q(R4[29]) );
  TLATX1 R4_reg_22_ ( .G(n276), .D(data_in_3_22_), .Q(R4[22]) );
  TLATX1 R4_reg_21_ ( .G(n276), .D(data_in_3_21_), .Q(R4[21]) );
  TLATX1 R4_reg_20_ ( .G(n276), .D(data_in_3_20_), .Q(R4[20]) );
  TLATX1 R4_reg_19_ ( .G(n276), .D(data_in_3_19_), .Q(R4[19]) );
  TLATX1 R4_reg_18_ ( .G(n276), .D(data_in_3_18_), .Q(R4[18]) );
  TLATX1 R4_reg_17_ ( .G(n276), .D(data_in_3_17_), .Q(R4[17]) );
  TLATXL R4_reg_16_ ( .G(n276), .D(data_in_3_16_), .Q(R4[16]) );
  TLATXL R4_reg_15_ ( .G(n276), .D(data_in_3_15_), .Q(R4[15]) );
  TLATXL R4_reg_13_ ( .G(n276), .D(data_in_3_13_), .Q(R4[13]) );
  TLATXL R4_reg_12_ ( .G(n276), .D(data_in_3_12_), .Q(R4[12]) );
  TLATX1 R3_reg_1_ ( .G(n82), .D(data_in_3_1_), .Q(R3[1]) );
  TLATX1 R4_reg_2_ ( .G(n276), .D(data_in_3_2_), .Q(R4[2]) );
  TLATXL R2_reg_28_ ( .G(n81), .D(data_in_3_28_), .Q(R2[28]) );
  TLATXL R2_reg_26_ ( .G(n81), .D(data_in_3_26_), .Q(R2[26]) );
  TLATXL R2_reg_24_ ( .G(n81), .D(data_in_3_24_), .Q(R2[24]) );
  TLATXL R2_reg_10_ ( .G(n81), .D(data_in_3_10_), .Q(R2[10]) );
  TLATXL R1_reg_23_ ( .G(n274), .D(data_in_3_23_), .Q(R1[23]) );
  TLATXL R3_reg_27_ ( .G(n82), .D(data_in_3_27_), .Q(R3[27]) );
  TLATXL R3_reg_10_ ( .G(n82), .D(data_in_3_10_), .Q(R3[10]) );
  TLATXL R4_reg_27_ ( .G(n276), .D(data_in_3_27_), .Q(R4[27]) );
  TLATXL R4_reg_25_ ( .G(n276), .D(data_in_3_25_), .Q(R4[25]) );
  TLATXL R4_reg_24_ ( .G(n276), .D(data_in_3_24_), .Q(R4[24]) );
  TLATXL R4_reg_23_ ( .G(n276), .D(data_in_3_23_), .Q(R4[23]) );
  TLATXL R4_reg_10_ ( .G(n276), .D(data_in_3_10_), .Q(R4[10]) );
  TLATXL R3_reg_23_ ( .G(n82), .D(data_in_3_23_), .Q(R3[23]) );
  TLATXL R3_reg_25_ ( .G(n82), .D(data_in_3_25_), .Q(R3[25]) );
  TLATXL R2_reg_23_ ( .G(n81), .D(data_in_3_23_), .Q(R2[23]) );
  TLATXL R2_reg_11_ ( .G(n81), .D(data_in_3_11_), .Q(R2[11]) );
  TLATXL R3_reg_11_ ( .G(n82), .D(data_in_3_11_), .Q(R3[11]) );
  TLATXL R3_reg_24_ ( .G(n82), .D(data_in_3_24_), .Q(R3[24]) );
  TLATXL R2_reg_25_ ( .G(n81), .D(data_in_3_25_), .Q(R2[25]) );
  TLATXL R1_reg_27_ ( .G(n285), .D(data_in_3_27_), .Q(R1[27]) );
  TLATXL R4_reg_28_ ( .G(n276), .D(data_in_3_28_), .Q(R4[28]) );
  TLATXL R3_reg_28_ ( .G(n82), .D(data_in_3_28_), .Q(R3[28]) );
  TLATXL R4_reg_11_ ( .G(n276), .D(data_in_3_11_), .Q(R4[11]) );
  TLATXL R2_reg_27_ ( .G(n81), .D(data_in_3_27_), .Q(R2[27]) );
  TLATXL R3_reg_26_ ( .G(n82), .D(data_in_3_26_), .Q(R3[26]) );
  TLATXL R4_reg_26_ ( .G(n276), .D(data_in_3_26_), .Q(R4[26]) );
  TLATXL R2_reg_6_ ( .G(n81), .D(data_in_3_6_), .Q(R2[6]) );
  TLATXL R2_reg_7_ ( .G(n81), .D(data_in_3_7_), .Q(R2[7]) );
  TLATXL R2_reg_9_ ( .G(n81), .D(data_in_3_9_), .Q(R2[9]) );
  TLATXL R2_reg_8_ ( .G(n81), .D(data_in_3_8_), .Q(R2[8]) );
  TLATXL R3_reg_8_ ( .G(n82), .D(data_in_3_8_), .Q(R3[8]) );
  TLATXL R3_reg_7_ ( .G(n82), .D(data_in_3_7_), .Q(R3[7]) );
  TLATXL R4_reg_9_ ( .G(n276), .D(data_in_3_9_), .Q(R4[9]) );
  TLATXL R4_reg_6_ ( .G(n276), .D(data_in_3_6_), .Q(R4[6]) );
  TLATXL R4_reg_7_ ( .G(n276), .D(data_in_3_7_), .Q(R4[7]) );
  TLATXL R3_reg_6_ ( .G(n82), .D(data_in_3_6_), .Q(R3[6]) );
  TLATXL R3_reg_9_ ( .G(n82), .D(data_in_3_9_), .Q(R3[9]) );
  TLATXL R4_reg_8_ ( .G(n276), .D(data_in_3_8_), .Q(R4[8]) );
  TLATXL R1_reg_24_ ( .G(n274), .D(data_in_3_24_), .Q(R1[24]) );
  TLATXL R1_reg_10_ ( .G(n274), .D(data_in_3_10_), .Q(R1[10]) );
  TLATXL R1_reg_26_ ( .G(n285), .D(data_in_3_26_), .Q(R1[26]) );
  TLATXL R1_reg_25_ ( .G(n274), .D(data_in_3_25_), .Q(R1[25]) );
  TLATXL R1_reg_28_ ( .G(n274), .D(data_in_3_28_), .Q(R1[28]) );
  TLATXL R1_reg_11_ ( .G(n274), .D(data_in_3_11_), .Q(R1[11]) );
  TLATXL R1_reg_8_ ( .G(n285), .D(data_in_3_8_), .Q(R1[8]) );
  TLATXL R1_reg_6_ ( .G(n285), .D(data_in_3_6_), .Q(R1[6]) );
  TLATXL R1_reg_7_ ( .G(n285), .D(data_in_3_7_), .Q(R1[7]) );
  TLATXL R1_reg_9_ ( .G(n285), .D(data_in_3_9_), .Q(R1[9]) );
  DFFRHQX2 counter_reg_2_ ( .D(N7), .CK(clk), .RN(rst_n), .Q(counter[2]) );
  INVX2 U4 ( .A(counter[3]), .Y(n286) );
  AOI22X2 U5 ( .A0(R4[2]), .A1(n614), .B0(data_in_2[104]), .B1(n86), .Y(n615)
         );
  NOR2X1 U6 ( .A(n656), .B(n446), .Y(n447) );
  BUFX8 U7 ( .A(n253), .Y(n88) );
  CLKINVX1 U8 ( .A(n261), .Y(n253) );
  OAI2BB1X1 U9 ( .A0N(n605), .A1N(n659), .B0(n604), .Y(data_out[101]) );
  AND2X2 U10 ( .A(n277), .B(n659), .Y(n157) );
  NAND2X4 U11 ( .A(R3[18]), .B(n559), .Y(n561) );
  NAND3X4 U12 ( .A(data_in_1[120]), .B(n278), .C(n251), .Y(n663) );
  INVX2 U13 ( .A(n260), .Y(n261) );
  NAND3BX4 U14 ( .AN(n149), .B(n617), .C(n616), .Y(data_out[105]) );
  NAND3X4 U15 ( .A(n452), .B(n451), .C(n450), .Y(data_out[52]) );
  NAND3X1 U16 ( .A(n283), .B(data_in_2[52]), .C(n251), .Y(n452) );
  NAND2X2 U17 ( .A(R4[17]), .B(n614), .Y(n660) );
  INVX1 U18 ( .A(n262), .Y(n1) );
  INVX1 U19 ( .A(n262), .Y(n2) );
  INVX1 U20 ( .A(n262), .Y(n3) );
  BUFX3 U21 ( .A(n3), .Y(n4) );
  BUFX3 U22 ( .A(n3), .Y(n5) );
  INVX1 U23 ( .A(n263), .Y(n6) );
  BUFX3 U24 ( .A(n6), .Y(n7) );
  BUFX3 U25 ( .A(n6), .Y(n8) );
  INVX4 U26 ( .A(n157), .Y(n9) );
  INVXL U27 ( .A(n157), .Y(n10) );
  INVXL U28 ( .A(n157), .Y(n11) );
  INVXL U29 ( .A(n157), .Y(n12) );
  INVXL U30 ( .A(n9), .Y(n13) );
  CLKINVX1 U31 ( .A(n9), .Y(n14) );
  CLKINVXL U32 ( .A(n9), .Y(n15) );
  INVXL U33 ( .A(n9), .Y(n16) );
  INVXL U34 ( .A(n9), .Y(n17) );
  INVX1 U35 ( .A(n10), .Y(n18) );
  INVX1 U36 ( .A(n10), .Y(n19) );
  INVXL U37 ( .A(n10), .Y(n20) );
  INVXL U38 ( .A(n10), .Y(n21) );
  INVXL U39 ( .A(n10), .Y(n22) );
  INVX1 U40 ( .A(n11), .Y(n23) );
  INVX1 U41 ( .A(n11), .Y(n24) );
  INVX1 U42 ( .A(n11), .Y(n25) );
  INVX1 U43 ( .A(n11), .Y(n26) );
  INVX1 U44 ( .A(n11), .Y(n27) );
  INVX1 U45 ( .A(n12), .Y(n28) );
  INVX1 U46 ( .A(n12), .Y(n29) );
  INVX1 U47 ( .A(n12), .Y(n30) );
  INVX1 U48 ( .A(n12), .Y(n31) );
  INVX1 U49 ( .A(n12), .Y(n32) );
  INVX1 U50 ( .A(n1), .Y(n33) );
  INVX1 U51 ( .A(n1), .Y(n34) );
  INVX1 U52 ( .A(n1), .Y(n35) );
  INVX1 U53 ( .A(n1), .Y(n36) );
  INVX1 U54 ( .A(n33), .Y(n37) );
  INVX1 U55 ( .A(n33), .Y(n38) );
  INVX1 U56 ( .A(n33), .Y(n39) );
  INVX1 U57 ( .A(n33), .Y(n40) );
  INVX1 U58 ( .A(n33), .Y(n41) );
  INVX1 U59 ( .A(n34), .Y(n42) );
  INVX1 U60 ( .A(n34), .Y(n43) );
  INVX1 U61 ( .A(n34), .Y(n44) );
  INVX1 U62 ( .A(n34), .Y(n45) );
  INVX1 U63 ( .A(n34), .Y(n46) );
  INVX1 U64 ( .A(n35), .Y(n47) );
  INVX1 U65 ( .A(n35), .Y(n48) );
  INVX1 U66 ( .A(n35), .Y(n49) );
  INVX1 U67 ( .A(n35), .Y(n50) );
  INVX1 U68 ( .A(n35), .Y(n51) );
  INVX1 U69 ( .A(n36), .Y(n52) );
  INVX1 U70 ( .A(n36), .Y(n53) );
  INVX1 U71 ( .A(n36), .Y(n54) );
  INVX1 U72 ( .A(n36), .Y(n55) );
  INVX1 U73 ( .A(n36), .Y(n56) );
  INVX1 U74 ( .A(n2), .Y(n57) );
  INVX1 U75 ( .A(n2), .Y(n58) );
  INVX1 U76 ( .A(n2), .Y(n59) );
  INVX1 U77 ( .A(n2), .Y(n60) );
  INVX1 U78 ( .A(n57), .Y(n61) );
  INVX1 U79 ( .A(n57), .Y(n62) );
  INVX1 U80 ( .A(n57), .Y(n63) );
  INVX1 U81 ( .A(n57), .Y(n64) );
  INVX1 U82 ( .A(n57), .Y(n65) );
  INVX1 U83 ( .A(n58), .Y(n66) );
  INVX1 U84 ( .A(n58), .Y(n67) );
  INVX1 U85 ( .A(n58), .Y(n68) );
  INVX1 U86 ( .A(n58), .Y(n69) );
  INVX1 U87 ( .A(n58), .Y(n70) );
  INVX1 U88 ( .A(n59), .Y(n71) );
  INVX1 U89 ( .A(n59), .Y(n72) );
  INVX1 U90 ( .A(n59), .Y(n73) );
  INVX1 U91 ( .A(n59), .Y(n74) );
  INVX1 U92 ( .A(n59), .Y(n75) );
  INVX1 U93 ( .A(n60), .Y(n76) );
  INVX1 U94 ( .A(n60), .Y(n77) );
  INVX1 U95 ( .A(n60), .Y(n78) );
  INVX1 U96 ( .A(n60), .Y(n79) );
  INVX1 U97 ( .A(n60), .Y(n80) );
  INVXL U98 ( .A(n157), .Y(n263) );
  NAND2X2 U99 ( .A(data_in_1[54]), .B(n17), .Y(n456) );
  NAND2XL U100 ( .A(data_in_1[88]), .B(n18), .Y(n150) );
  NAND2XL U101 ( .A(data_in_1[122]), .B(n16), .Y(n153) );
  NAND3XL U102 ( .A(n280), .B(data_in_2[103]), .C(n251), .Y(n613) );
  NAND2X2 U103 ( .A(R4[19]), .B(n265), .Y(n666) );
  OR2X2 U104 ( .A(n95), .B(n391), .Y(n147) );
  NAND3X2 U105 ( .A(n404), .B(n403), .C(n402), .Y(data_out[37]) );
  NAND3X2 U106 ( .A(n514), .B(n513), .C(n512), .Y(data_out[71]) );
  INVXL U107 ( .A(data_in_2[67]), .Y(n495) );
  INVX1 U108 ( .A(data_in_2[50]), .Y(n442) );
  NAND2BX1 U109 ( .AN(n278), .B(data_in_2[34]), .Y(n392) );
  NAND2BX1 U110 ( .AN(n278), .B(data_in_2[51]), .Y(n446) );
  BUFX3 U111 ( .A(n252), .Y(n90) );
  NAND2X1 U112 ( .A(data_in_1[13]), .B(n50), .Y(n329) );
  NAND2X1 U113 ( .A(R3[33]), .B(n708), .Y(n604) );
  BUFX3 U114 ( .A(n258), .Y(n93) );
  BUFX3 U115 ( .A(n256), .Y(n92) );
  BUFX3 U116 ( .A(n257), .Y(n91) );
  OAI2BB1X1 U117 ( .A0N(n711), .A1N(n710), .B0(n709), .Y(data_out[135]) );
  BUFX3 U118 ( .A(n259), .Y(n94) );
  BUFX3 U119 ( .A(n255), .Y(n89) );
  BUFX3 U120 ( .A(n254), .Y(n87) );
  OAI2BB1X2 U121 ( .A0N(n554), .A1N(n659), .B0(n553), .Y(data_out[84]) );
  NAND2X1 U122 ( .A(R3[16]), .B(n708), .Y(n553) );
  OAI2BB1X1 U123 ( .A0N(n658), .A1N(n710), .B0(n657), .Y(data_out[118]) );
  OR3XL U124 ( .A(counter[1]), .B(counter[2]), .C(counter[3]), .Y(n141) );
  INVXL U125 ( .A(n702), .Y(n271) );
  NOR3X1 U126 ( .A(n282), .B(n720), .C(n286), .Y(n81) );
  BUFX3 U127 ( .A(n260), .Y(n86) );
  CLKINVX4 U128 ( .A(n702), .Y(n273) );
  NOR2X1 U129 ( .A(n83), .B(n141), .Y(n82) );
  NAND2X1 U130 ( .A(n659), .B(n279), .Y(n379) );
  INVX4 U131 ( .A(mux_flag), .Y(n284) );
  INVX8 U132 ( .A(n284), .Y(n278) );
  INVX2 U133 ( .A(n272), .Y(n267) );
  CLKINVX3 U134 ( .A(n272), .Y(n265) );
  AND2X4 U135 ( .A(n147), .B(n148), .Y(n393) );
  XOR2X1 U136 ( .A(counter[1]), .B(n83), .Y(N6) );
  NAND2X1 U137 ( .A(R2[20]), .B(n268), .Y(n455) );
  INVX1 U138 ( .A(n271), .Y(n268) );
  DLY1X1 U139 ( .A(n242), .Y(n83) );
  CLKINVX4 U140 ( .A(n140), .Y(n242) );
  NAND2X1 U141 ( .A(R3[17]), .B(n614), .Y(n557) );
  INVX2 U142 ( .A(n702), .Y(n272) );
  NAND3X2 U143 ( .A(n668), .B(n667), .C(n666), .Y(data_out[121]) );
  NAND3X1 U144 ( .A(data_in_1[86]), .B(n710), .C(n278), .Y(n560) );
  INVX4 U145 ( .A(n659), .Y(n708) );
  INVX3 U146 ( .A(n273), .Y(n264) );
  OAI2BB1X4 U147 ( .A0N(data_in_1[104]), .A1N(n14), .B0(n615), .Y(
        data_out[104]) );
  NAND2X1 U148 ( .A(R4[1]), .B(n614), .Y(n611) );
  NOR2X1 U149 ( .A(n95), .B(n606), .Y(n609) );
  INVX4 U150 ( .A(n273), .Y(n95) );
  NAND3X4 U151 ( .A(n280), .B(data_in_2[120]), .C(n251), .Y(n664) );
  BUFX12 U152 ( .A(n710), .Y(n251) );
  NAND2X2 U153 ( .A(data_in_1[36]), .B(n13), .Y(n400) );
  NAND3X1 U154 ( .A(data_in_1[103]), .B(n278), .C(n251), .Y(n612) );
  NOR2X1 U155 ( .A(n95), .B(n607), .Y(n608) );
  NAND3X1 U156 ( .A(data_in_1[52]), .B(n278), .C(n251), .Y(n451) );
  NOR2X1 U157 ( .A(n448), .B(n447), .Y(n449) );
  INVX4 U158 ( .A(n251), .Y(n559) );
  AND3X2 U159 ( .A(n283), .B(data_in_2[119]), .C(n659), .Y(n158) );
  NAND2X2 U160 ( .A(R4[18]), .B(n614), .Y(n662) );
  NAND3X4 U161 ( .A(n664), .B(n663), .C(n662), .Y(data_out[120]) );
  NAND2X1 U162 ( .A(data_in_1[101]), .B(n278), .Y(n602) );
  INVX4 U163 ( .A(n665), .Y(n702) );
  NAND2X1 U164 ( .A(R4[16]), .B(n656), .Y(n657) );
  OAI21X1 U165 ( .A0(n277), .A1(n552), .B0(n551), .Y(n554) );
  NAND2X1 U166 ( .A(data_in_1[84]), .B(n278), .Y(n551) );
  OAI21X1 U167 ( .A0(n277), .A1(n603), .B0(n602), .Y(n605) );
  NAND2X1 U168 ( .A(R2[18]), .B(n614), .Y(n450) );
  AOI21X2 U169 ( .A0(R3[1]), .A1(n614), .B0(n504), .Y(n505) );
  NOR2X2 U170 ( .A(n614), .B(n503), .Y(n504) );
  NAND2BX1 U171 ( .AN(n665), .B(R2[19]), .Y(n160) );
  INVX4 U172 ( .A(n665), .Y(n614) );
  CLKBUFXL U173 ( .A(n379), .Y(n84) );
  BUFX3 U174 ( .A(n86), .Y(n85) );
  INVXL U175 ( .A(n261), .Y(n255) );
  INVXL U176 ( .A(n261), .Y(n257) );
  INVXL U177 ( .A(n261), .Y(n256) );
  INVXL U178 ( .A(n84), .Y(n258) );
  INVXL U179 ( .A(n84), .Y(n259) );
  INVX2 U180 ( .A(n710), .Y(n656) );
  OAI2BB1X1 U181 ( .A0N(n444), .A1N(n710), .B0(n443), .Y(data_out[50]) );
  OAI2BB1X1 U182 ( .A0N(n497), .A1N(n710), .B0(n496), .Y(data_out[67]) );
  NAND2BX4 U183 ( .AN(n242), .B(n390), .Y(n710) );
  CLKINVX8 U184 ( .A(n284), .Y(n277) );
  INVX2 U185 ( .A(n271), .Y(n269) );
  NAND2X1 U186 ( .A(data_in_1[135]), .B(n277), .Y(n706) );
  NAND3BX2 U187 ( .AN(n159), .B(n150), .C(n151), .Y(data_out[88]) );
  NAND2X1 U188 ( .A(R2[33]), .B(n656), .Y(n496) );
  NOR2X1 U189 ( .A(n510), .B(n509), .Y(n511) );
  NAND2BXL U190 ( .AN(n278), .B(data_in_2[69]), .Y(n503) );
  NAND2XL U191 ( .A(R2[16]), .B(n559), .Y(n443) );
  INVXL U192 ( .A(n157), .Y(n262) );
  OR2XL U193 ( .A(n656), .B(n392), .Y(n148) );
  NOR2X1 U194 ( .A(n397), .B(n396), .Y(n398) );
  NOR2XL U195 ( .A(n614), .B(n395), .Y(n396) );
  NOR2X1 U196 ( .A(n609), .B(n608), .Y(n610) );
  NOR2XL U197 ( .A(n656), .B(n445), .Y(n448) );
  NAND2X1 U198 ( .A(R4[33]), .B(n708), .Y(n709) );
  INVX1 U199 ( .A(n160), .Y(n453) );
  AND2X2 U200 ( .A(data_in_2[105]), .B(n90), .Y(n149) );
  NAND2XL U201 ( .A(R3[20]), .B(n267), .Y(n151) );
  NAND3X2 U202 ( .A(n152), .B(n153), .C(n154), .Y(data_out[122]) );
  NAND2XL U203 ( .A(data_in_2[122]), .B(n85), .Y(n152) );
  NAND2XL U204 ( .A(R4[20]), .B(n265), .Y(n154) );
  NAND2BXL U205 ( .AN(n278), .B(data_in_2[35]), .Y(n395) );
  OAI21XL U206 ( .A0(n277), .A1(n655), .B0(n654), .Y(n658) );
  NAND2BXL U207 ( .AN(n278), .B(data_in_2[102]), .Y(n607) );
  NAND2XL U208 ( .A(R3[4]), .B(n268), .Y(n515) );
  NAND2XL U209 ( .A(R4[4]), .B(n266), .Y(n618) );
  NAND2XL U210 ( .A(R3[5]), .B(n269), .Y(n518) );
  NAND2XL U211 ( .A(R4[5]), .B(n266), .Y(n621) );
  NAND2XL U212 ( .A(R3[22]), .B(n266), .Y(n569) );
  NAND2XL U213 ( .A(data_in_1[56]), .B(n31), .Y(n462) );
  NAND2XL U214 ( .A(data_in_1[57]), .B(n27), .Y(n465) );
  NAND2XL U215 ( .A(R3[6]), .B(n269), .Y(n521) );
  NAND2XL U216 ( .A(R2[24]), .B(n266), .Y(n467) );
  NAND2XL U217 ( .A(data_in_1[58]), .B(n40), .Y(n468) );
  NAND2XL U218 ( .A(R3[24]), .B(n266), .Y(n575) );
  NAND2XL U219 ( .A(data_in_1[59]), .B(n48), .Y(n471) );
  NAND2XL U220 ( .A(R3[25]), .B(n266), .Y(n578) );
  NAND2XL U221 ( .A(R2[26]), .B(n268), .Y(n473) );
  NAND2XL U222 ( .A(data_in_1[60]), .B(n52), .Y(n474) );
  NAND2XL U223 ( .A(R2[27]), .B(n269), .Y(n476) );
  NAND2XL U224 ( .A(data_in_1[61]), .B(n63), .Y(n477) );
  NAND2XL U225 ( .A(R3[26]), .B(n266), .Y(n581) );
  NAND2XL U226 ( .A(R3[27]), .B(n266), .Y(n584) );
  NAND2XL U227 ( .A(R3[28]), .B(n266), .Y(n587) );
  NAND2XL U228 ( .A(R3[29]), .B(n266), .Y(n590) );
  NAND2XL U229 ( .A(R3[30]), .B(n266), .Y(n593) );
  NAND2XL U230 ( .A(R2[29]), .B(n269), .Y(n482) );
  NAND2XL U231 ( .A(data_in_1[63]), .B(n72), .Y(n483) );
  NAND2XL U232 ( .A(R2[30]), .B(n268), .Y(n485) );
  NAND2XL U233 ( .A(data_in_1[64]), .B(n13), .Y(n486) );
  NAND2XL U234 ( .A(R2[28]), .B(n266), .Y(n479) );
  NAND2XL U235 ( .A(data_in_1[62]), .B(n70), .Y(n480) );
  NAND2XL U236 ( .A(R3[31]), .B(n266), .Y(n596) );
  NAND2XL U237 ( .A(R4[32]), .B(n269), .Y(n703) );
  NAND2XL U238 ( .A(data_in_1[134]), .B(n27), .Y(n704) );
  NAND2XL U239 ( .A(R3[32]), .B(n266), .Y(n599) );
  NAND2XL U240 ( .A(R2[31]), .B(n269), .Y(n488) );
  NAND2XL U241 ( .A(data_in_1[65]), .B(n21), .Y(n489) );
  NAND2XL U242 ( .A(R2[32]), .B(n266), .Y(n491) );
  NAND2XL U243 ( .A(data_in_1[66]), .B(n25), .Y(n492) );
  OR2X2 U244 ( .A(n380), .B(n155), .Y(data_out[30]) );
  AND2X1 U245 ( .A(R1[30]), .B(n269), .Y(n155) );
  NAND2X1 U246 ( .A(n156), .B(n266), .Y(n328) );
  INVX1 U247 ( .A(n84), .Y(n252) );
  INVX1 U248 ( .A(n261), .Y(n254) );
  INVX1 U249 ( .A(n272), .Y(n266) );
  INVX1 U250 ( .A(n273), .Y(n270) );
  INVX1 U251 ( .A(n379), .Y(n260) );
  INVXL U252 ( .A(mux_flag), .Y(n279) );
  INVXL U253 ( .A(mux_flag), .Y(n280) );
  INVXL U254 ( .A(mux_flag), .Y(n283) );
  XOR2X1 U255 ( .A(n720), .B(n282), .Y(N7) );
  INVX1 U256 ( .A(n162), .Y(n276) );
  INVX1 U257 ( .A(n275), .Y(n274) );
  NAND3BX4 U258 ( .AN(n158), .B(n661), .C(n660), .Y(data_out[119]) );
  OAI21XL U259 ( .A0(n277), .A1(n556), .B0(n555), .Y(n558) );
  INVX1 U260 ( .A(data_in_2[85]), .Y(n556) );
  NOR2BXL U261 ( .AN(data_in_1[69]), .B(n279), .Y(n506) );
  NAND2X1 U262 ( .A(R3[3]), .B(n269), .Y(n512) );
  NAND2X2 U263 ( .A(data_in_1[71]), .B(n21), .Y(n513) );
  NAND2X2 U264 ( .A(data_in_2[71]), .B(n91), .Y(n514) );
  AND2X2 U265 ( .A(data_in_2[88]), .B(n87), .Y(n159) );
  NOR2X1 U266 ( .A(n559), .B(n394), .Y(n397) );
  NAND2XL U267 ( .A(R2[3]), .B(n269), .Y(n402) );
  NAND2XL U268 ( .A(data_in_1[37]), .B(n20), .Y(n403) );
  NAND2XL U269 ( .A(data_in_2[37]), .B(n92), .Y(n404) );
  NAND2X1 U270 ( .A(R4[3]), .B(n266), .Y(n616) );
  NAND2X2 U271 ( .A(data_in_1[105]), .B(n19), .Y(n617) );
  OAI2BB1X2 U272 ( .A0N(R3[2]), .A1N(n270), .B0(n511), .Y(data_out[70]) );
  NOR2X2 U273 ( .A(n264), .B(n507), .Y(n510) );
  NOR2X2 U274 ( .A(n264), .B(n508), .Y(n509) );
  NAND3X1 U275 ( .A(n568), .B(n567), .C(n566), .Y(data_out[89]) );
  NAND2XL U276 ( .A(R3[21]), .B(n267), .Y(n566) );
  NAND2XL U277 ( .A(data_in_1[89]), .B(n22), .Y(n567) );
  NAND2XL U278 ( .A(data_in_2[89]), .B(n85), .Y(n568) );
  NAND3X1 U279 ( .A(n517), .B(n516), .C(n515), .Y(data_out[72]) );
  NAND2XL U280 ( .A(data_in_1[72]), .B(n24), .Y(n516) );
  NAND2XL U281 ( .A(data_in_2[72]), .B(n93), .Y(n517) );
  NAND3X1 U282 ( .A(n671), .B(n670), .C(n669), .Y(data_out[123]) );
  NAND2XL U283 ( .A(R4[21]), .B(n264), .Y(n669) );
  NAND2XL U284 ( .A(data_in_1[123]), .B(n23), .Y(n670) );
  NAND2XL U285 ( .A(data_in_2[123]), .B(n89), .Y(n671) );
  NAND3X1 U286 ( .A(n407), .B(n406), .C(n405), .Y(data_out[38]) );
  NAND2XL U287 ( .A(R2[4]), .B(n269), .Y(n405) );
  NAND2XL U288 ( .A(data_in_1[38]), .B(n28), .Y(n406) );
  NAND2XL U289 ( .A(data_in_2[38]), .B(n87), .Y(n407) );
  NAND3X1 U290 ( .A(n460), .B(n459), .C(n458), .Y(data_out[55]) );
  NAND2XL U291 ( .A(R2[21]), .B(n268), .Y(n458) );
  NAND2X1 U292 ( .A(data_in_1[55]), .B(n25), .Y(n459) );
  NAND2XL U293 ( .A(data_in_2[55]), .B(n88), .Y(n460) );
  NAND3X1 U294 ( .A(n410), .B(n409), .C(n408), .Y(data_out[39]) );
  NAND2XL U295 ( .A(R2[5]), .B(n269), .Y(n408) );
  NAND2XL U296 ( .A(data_in_1[39]), .B(n29), .Y(n409) );
  NAND2XL U297 ( .A(data_in_2[39]), .B(n94), .Y(n410) );
  NAND3X1 U298 ( .A(n520), .B(n519), .C(n518), .Y(data_out[73]) );
  NAND2XL U299 ( .A(data_in_1[73]), .B(n38), .Y(n519) );
  NAND2XL U300 ( .A(data_in_2[73]), .B(n91), .Y(n520) );
  NAND3X1 U301 ( .A(n463), .B(n462), .C(n461), .Y(data_out[56]) );
  NAND2XL U302 ( .A(R2[22]), .B(n268), .Y(n461) );
  NAND2XL U303 ( .A(data_in_2[56]), .B(n89), .Y(n463) );
  NAND3X1 U304 ( .A(n413), .B(n412), .C(n411), .Y(data_out[40]) );
  NAND2XL U305 ( .A(R2[6]), .B(n269), .Y(n411) );
  NAND2XL U306 ( .A(data_in_1[40]), .B(n4), .Y(n412) );
  NAND2XL U307 ( .A(data_in_2[40]), .B(n91), .Y(n413) );
  NAND3X1 U308 ( .A(n620), .B(n619), .C(n618), .Y(data_out[106]) );
  NAND2XL U309 ( .A(data_in_1[106]), .B(n26), .Y(n619) );
  NAND2XL U310 ( .A(data_in_2[106]), .B(n86), .Y(n620) );
  NAND3X1 U311 ( .A(n523), .B(n522), .C(n521), .Y(data_out[74]) );
  NAND2XL U312 ( .A(data_in_1[74]), .B(n7), .Y(n522) );
  NAND2XL U313 ( .A(data_in_2[74]), .B(n87), .Y(n523) );
  NAND3X1 U314 ( .A(n466), .B(n465), .C(n464), .Y(data_out[57]) );
  NAND2XL U315 ( .A(R2[23]), .B(n268), .Y(n464) );
  NAND2XL U316 ( .A(data_in_2[57]), .B(n88), .Y(n466) );
  NAND3X1 U317 ( .A(n571), .B(n570), .C(n569), .Y(data_out[90]) );
  NAND2XL U318 ( .A(data_in_1[90]), .B(n5), .Y(n570) );
  NAND2XL U319 ( .A(data_in_2[90]), .B(n90), .Y(n571) );
  NAND3X1 U320 ( .A(n623), .B(n622), .C(n621), .Y(data_out[107]) );
  NAND2XL U321 ( .A(data_in_1[107]), .B(n37), .Y(n622) );
  NAND2XL U322 ( .A(data_in_2[107]), .B(n93), .Y(n623) );
  NAND3X1 U323 ( .A(n674), .B(n673), .C(n672), .Y(data_out[124]) );
  NAND2XL U324 ( .A(R4[22]), .B(n265), .Y(n672) );
  NAND2XL U325 ( .A(data_in_1[124]), .B(n32), .Y(n673) );
  NAND2XL U326 ( .A(data_in_2[124]), .B(n92), .Y(n674) );
  NAND3X1 U327 ( .A(n574), .B(n573), .C(n572), .Y(data_out[91]) );
  NAND2XL U328 ( .A(R3[23]), .B(n267), .Y(n572) );
  NAND2XL U329 ( .A(data_in_1[91]), .B(n8), .Y(n573) );
  NAND2XL U330 ( .A(data_in_2[91]), .B(n85), .Y(n574) );
  NAND3X1 U331 ( .A(n677), .B(n676), .C(n675), .Y(data_out[125]) );
  NAND2XL U332 ( .A(R4[23]), .B(n264), .Y(n675) );
  NAND2XL U333 ( .A(data_in_1[125]), .B(n39), .Y(n676) );
  NAND2XL U334 ( .A(data_in_2[125]), .B(n86), .Y(n677) );
  NAND2X4 U335 ( .A(n140), .B(n390), .Y(n659) );
  NAND2XL U336 ( .A(data_in_1[51]), .B(n277), .Y(n445) );
  NAND2XL U337 ( .A(data_in_1[34]), .B(n277), .Y(n391) );
  NAND2XL U338 ( .A(data_in_1[35]), .B(n278), .Y(n394) );
  NAND2XL U339 ( .A(data_in_1[50]), .B(n277), .Y(n441) );
  NAND2BXL U340 ( .AN(n278), .B(data_in_2[70]), .Y(n508) );
  NAND2XL U341 ( .A(data_in_1[118]), .B(n278), .Y(n654) );
  OAI21XL U342 ( .A0(n277), .A1(n495), .B0(n494), .Y(n497) );
  OAI21XL U343 ( .A0(n277), .A1(n707), .B0(n706), .Y(n711) );
  INVX1 U344 ( .A(data_in_2[118]), .Y(n655) );
  INVX1 U345 ( .A(data_in_2[84]), .Y(n552) );
  INVX1 U346 ( .A(data_in_2[101]), .Y(n603) );
  OAI21XL U347 ( .A0(n277), .A1(n442), .B0(n441), .Y(n444) );
  NAND2BXL U348 ( .AN(n278), .B(data_in_2[68]), .Y(n498) );
  INVX1 U349 ( .A(data_in_2[135]), .Y(n707) );
  NAND3X1 U350 ( .A(n641), .B(n640), .C(n639), .Y(data_out[113]) );
  NAND2XL U351 ( .A(R4[11]), .B(n265), .Y(n639) );
  NAND2XL U352 ( .A(data_in_1[113]), .B(n68), .Y(n640) );
  NAND2XL U353 ( .A(data_in_2[113]), .B(n88), .Y(n641) );
  NAND3X1 U354 ( .A(n538), .B(n537), .C(n536), .Y(data_out[79]) );
  NAND2XL U355 ( .A(R3[11]), .B(n267), .Y(n536) );
  NAND2XL U356 ( .A(data_in_1[79]), .B(n69), .Y(n537) );
  NAND2XL U357 ( .A(data_in_2[79]), .B(n94), .Y(n538) );
  NAND3X1 U358 ( .A(n416), .B(n415), .C(n414), .Y(data_out[41]) );
  NAND2XL U359 ( .A(R2[7]), .B(n269), .Y(n414) );
  NAND2XL U360 ( .A(data_in_1[41]), .B(n45), .Y(n415) );
  NAND2XL U361 ( .A(data_in_2[41]), .B(n85), .Y(n416) );
  NAND3X1 U362 ( .A(n526), .B(n525), .C(n524), .Y(data_out[75]) );
  NAND2XL U363 ( .A(R3[7]), .B(n267), .Y(n524) );
  NAND2XL U364 ( .A(data_in_1[75]), .B(n42), .Y(n525) );
  NAND2XL U365 ( .A(data_in_2[75]), .B(n93), .Y(n526) );
  NAND3X1 U366 ( .A(n469), .B(n468), .C(n467), .Y(data_out[58]) );
  NAND2XL U367 ( .A(data_in_2[58]), .B(n88), .Y(n469) );
  NAND3X1 U368 ( .A(n419), .B(n418), .C(n417), .Y(data_out[42]) );
  NAND2XL U369 ( .A(R2[8]), .B(n268), .Y(n417) );
  NAND2XL U370 ( .A(data_in_1[42]), .B(n51), .Y(n418) );
  NAND2XL U371 ( .A(data_in_2[42]), .B(n90), .Y(n419) );
  NAND3X1 U372 ( .A(n626), .B(n625), .C(n624), .Y(data_out[108]) );
  NAND2XL U373 ( .A(R4[6]), .B(n265), .Y(n624) );
  NAND2XL U374 ( .A(data_in_1[108]), .B(n30), .Y(n625) );
  NAND2XL U375 ( .A(data_in_2[108]), .B(n90), .Y(n626) );
  NAND3X1 U376 ( .A(n529), .B(n528), .C(n527), .Y(data_out[76]) );
  NAND2XL U377 ( .A(R3[8]), .B(n267), .Y(n527) );
  NAND2XL U378 ( .A(data_in_1[76]), .B(n49), .Y(n528) );
  NAND2XL U379 ( .A(data_in_2[76]), .B(n87), .Y(n529) );
  NAND3X1 U380 ( .A(n472), .B(n471), .C(n470), .Y(data_out[59]) );
  NAND2XL U381 ( .A(R2[25]), .B(n268), .Y(n470) );
  NAND2XL U382 ( .A(data_in_2[59]), .B(n91), .Y(n472) );
  NAND3X1 U383 ( .A(n422), .B(n421), .C(n420), .Y(data_out[43]) );
  NAND2XL U384 ( .A(R2[9]), .B(n268), .Y(n420) );
  NAND2XL U385 ( .A(data_in_1[43]), .B(n61), .Y(n421) );
  NAND2XL U386 ( .A(data_in_2[43]), .B(n86), .Y(n422) );
  NAND3X1 U387 ( .A(n577), .B(n576), .C(n575), .Y(data_out[92]) );
  NAND2XL U388 ( .A(data_in_1[92]), .B(n43), .Y(n576) );
  NAND2XL U389 ( .A(data_in_2[92]), .B(n92), .Y(n577) );
  NAND3X1 U390 ( .A(n629), .B(n628), .C(n627), .Y(data_out[109]) );
  NAND2XL U391 ( .A(R4[7]), .B(n265), .Y(n627) );
  NAND2XL U392 ( .A(data_in_1[109]), .B(n44), .Y(n628) );
  NAND2XL U393 ( .A(data_in_2[109]), .B(n94), .Y(n629) );
  NAND3X1 U394 ( .A(n680), .B(n679), .C(n678), .Y(data_out[126]) );
  NAND2XL U395 ( .A(R4[24]), .B(n264), .Y(n678) );
  NAND2XL U396 ( .A(data_in_1[126]), .B(n41), .Y(n679) );
  NAND2XL U397 ( .A(data_in_2[126]), .B(n86), .Y(n680) );
  NAND3X1 U398 ( .A(n532), .B(n531), .C(n530), .Y(data_out[77]) );
  NAND2XL U399 ( .A(R3[9]), .B(n267), .Y(n530) );
  NAND2XL U400 ( .A(data_in_1[77]), .B(n55), .Y(n531) );
  NAND2XL U401 ( .A(data_in_2[77]), .B(n85), .Y(n532) );
  NAND3X1 U402 ( .A(n475), .B(n474), .C(n473), .Y(data_out[60]) );
  NAND2XL U403 ( .A(data_in_2[60]), .B(n88), .Y(n475) );
  NAND3X1 U404 ( .A(n580), .B(n579), .C(n578), .Y(data_out[93]) );
  NAND2XL U405 ( .A(data_in_1[93]), .B(n47), .Y(n579) );
  NAND2XL U406 ( .A(data_in_2[93]), .B(n89), .Y(n580) );
  NAND3X1 U407 ( .A(n632), .B(n631), .C(n630), .Y(data_out[110]) );
  NAND2XL U408 ( .A(R4[8]), .B(n265), .Y(n630) );
  NAND2XL U409 ( .A(data_in_1[110]), .B(n50), .Y(n631) );
  NAND2XL U410 ( .A(data_in_2[110]), .B(n92), .Y(n632) );
  NAND3X1 U411 ( .A(n683), .B(n682), .C(n681), .Y(data_out[127]) );
  NAND2XL U412 ( .A(R4[25]), .B(n264), .Y(n681) );
  NAND2XL U413 ( .A(data_in_1[127]), .B(n46), .Y(n682) );
  NAND2XL U414 ( .A(data_in_2[127]), .B(n93), .Y(n683) );
  NAND3X1 U415 ( .A(n535), .B(n534), .C(n533), .Y(data_out[78]) );
  NAND2XL U416 ( .A(R3[10]), .B(n267), .Y(n533) );
  NAND2XL U417 ( .A(data_in_1[78]), .B(n66), .Y(n534) );
  NAND2XL U418 ( .A(data_in_2[78]), .B(n90), .Y(n535) );
  NAND3X1 U419 ( .A(n583), .B(n582), .C(n581), .Y(data_out[94]) );
  NAND2XL U420 ( .A(data_in_1[94]), .B(n56), .Y(n582) );
  NAND2XL U421 ( .A(data_in_2[94]), .B(n94), .Y(n583) );
  NAND3X1 U422 ( .A(n635), .B(n634), .C(n633), .Y(data_out[111]) );
  NAND2XL U423 ( .A(R4[9]), .B(n265), .Y(n633) );
  NAND2XL U424 ( .A(data_in_1[111]), .B(n54), .Y(n634) );
  NAND2XL U425 ( .A(data_in_2[111]), .B(n89), .Y(n635) );
  NAND3X1 U426 ( .A(n686), .B(n685), .C(n684), .Y(data_out[128]) );
  NAND2XL U427 ( .A(R4[26]), .B(n264), .Y(n684) );
  NAND2XL U428 ( .A(data_in_1[128]), .B(n53), .Y(n685) );
  NAND2XL U429 ( .A(data_in_2[128]), .B(n87), .Y(n686) );
  NAND3X1 U430 ( .A(n638), .B(n637), .C(n636), .Y(data_out[112]) );
  NAND2XL U431 ( .A(R4[10]), .B(n265), .Y(n636) );
  NAND2XL U432 ( .A(data_in_1[112]), .B(n67), .Y(n637) );
  NAND2XL U433 ( .A(data_in_2[112]), .B(n89), .Y(n638) );
  NAND3X1 U434 ( .A(n428), .B(n427), .C(n426), .Y(data_out[45]) );
  NAND2XL U435 ( .A(R2[11]), .B(n268), .Y(n426) );
  NAND2XL U436 ( .A(data_in_1[45]), .B(n74), .Y(n427) );
  NAND2XL U437 ( .A(data_in_2[45]), .B(n85), .Y(n428) );
  NAND3X1 U438 ( .A(n541), .B(n540), .C(n539), .Y(data_out[80]) );
  NAND2XL U439 ( .A(R3[12]), .B(n267), .Y(n539) );
  NAND2XL U440 ( .A(data_in_1[80]), .B(n78), .Y(n540) );
  NAND2XL U441 ( .A(data_in_2[80]), .B(n94), .Y(n541) );
  NAND3X1 U442 ( .A(n487), .B(n486), .C(n485), .Y(data_out[64]) );
  NAND2XL U443 ( .A(data_in_2[64]), .B(n88), .Y(n487) );
  NAND3X1 U444 ( .A(n695), .B(n694), .C(n693), .Y(data_out[131]) );
  NAND2XL U445 ( .A(R4[29]), .B(n264), .Y(n693) );
  NAND2XL U446 ( .A(data_in_1[131]), .B(n77), .Y(n694) );
  NAND2XL U447 ( .A(data_in_2[131]), .B(n86), .Y(n695) );
  NAND3X1 U448 ( .A(n692), .B(n691), .C(n690), .Y(data_out[130]) );
  NAND2XL U449 ( .A(R4[28]), .B(n264), .Y(n690) );
  NAND2XL U450 ( .A(data_in_1[130]), .B(n65), .Y(n691) );
  NAND2XL U451 ( .A(data_in_2[130]), .B(n90), .Y(n692) );
  NAND3X1 U452 ( .A(n589), .B(n588), .C(n587), .Y(data_out[96]) );
  NAND2XL U453 ( .A(data_in_1[96]), .B(n73), .Y(n588) );
  NAND2XL U454 ( .A(data_in_2[96]), .B(n87), .Y(n589) );
  NAND3X1 U455 ( .A(n425), .B(n424), .C(n423), .Y(data_out[44]) );
  NAND2XL U456 ( .A(R2[10]), .B(n268), .Y(n423) );
  NAND2XL U457 ( .A(data_in_1[44]), .B(n71), .Y(n424) );
  NAND2XL U458 ( .A(data_in_2[44]), .B(n93), .Y(n425) );
  NAND3X1 U459 ( .A(n478), .B(n477), .C(n476), .Y(data_out[61]) );
  NAND2XL U460 ( .A(data_in_2[61]), .B(n92), .Y(n478) );
  NAND3X1 U461 ( .A(n481), .B(n480), .C(n479), .Y(data_out[62]) );
  NAND2XL U462 ( .A(data_in_2[62]), .B(n86), .Y(n481) );
  NAND3X1 U463 ( .A(n586), .B(n585), .C(n584), .Y(data_out[95]) );
  NAND2XL U464 ( .A(data_in_1[95]), .B(n64), .Y(n585) );
  NAND2XL U465 ( .A(data_in_2[95]), .B(n91), .Y(n586) );
  NAND3X1 U466 ( .A(n689), .B(n688), .C(n687), .Y(data_out[129]) );
  NAND2XL U467 ( .A(R4[27]), .B(n264), .Y(n687) );
  NAND2XL U468 ( .A(data_in_1[129]), .B(n62), .Y(n688) );
  NAND2XL U469 ( .A(data_in_2[129]), .B(n92), .Y(n689) );
  NAND3X1 U470 ( .A(n698), .B(n697), .C(n696), .Y(data_out[132]) );
  NAND2XL U471 ( .A(R4[30]), .B(n264), .Y(n696) );
  NAND2XL U472 ( .A(data_in_1[132]), .B(n15), .Y(n697) );
  NAND2XL U473 ( .A(data_in_2[132]), .B(n92), .Y(n698) );
  NAND3X1 U474 ( .A(n592), .B(n591), .C(n590), .Y(data_out[97]) );
  NAND2XL U475 ( .A(data_in_1[97]), .B(n76), .Y(n591) );
  NAND2XL U476 ( .A(data_in_2[97]), .B(n91), .Y(n592) );
  NAND3X1 U477 ( .A(n431), .B(n430), .C(n429), .Y(data_out[46]) );
  NAND2XL U478 ( .A(R2[12]), .B(n268), .Y(n429) );
  NAND2XL U479 ( .A(data_in_1[46]), .B(n79), .Y(n430) );
  NAND2XL U480 ( .A(data_in_2[46]), .B(n87), .Y(n431) );
  NAND3X1 U481 ( .A(n434), .B(n433), .C(n432), .Y(data_out[47]) );
  NAND2XL U482 ( .A(R2[13]), .B(n268), .Y(n432) );
  NAND2XL U483 ( .A(data_in_1[47]), .B(n17), .Y(n433) );
  NAND2XL U484 ( .A(data_in_2[47]), .B(n91), .Y(n434) );
  NAND3X1 U485 ( .A(n644), .B(n643), .C(n642), .Y(data_out[114]) );
  NAND2XL U486 ( .A(R4[12]), .B(n265), .Y(n642) );
  NAND2XL U487 ( .A(data_in_1[114]), .B(n75), .Y(n643) );
  NAND2XL U488 ( .A(data_in_2[114]), .B(n85), .Y(n644) );
  NAND3X1 U489 ( .A(n595), .B(n594), .C(n593), .Y(data_out[98]) );
  NAND2XL U490 ( .A(data_in_1[98]), .B(n14), .Y(n594) );
  NAND2XL U491 ( .A(data_in_2[98]), .B(n89), .Y(n595) );
  NAND3X1 U492 ( .A(n484), .B(n483), .C(n482), .Y(data_out[63]) );
  NAND2XL U493 ( .A(data_in_2[63]), .B(n93), .Y(n484) );
  NAND3X1 U494 ( .A(n647), .B(n646), .C(n645), .Y(data_out[115]) );
  NAND2XL U495 ( .A(R4[13]), .B(n265), .Y(n645) );
  NAND2XL U496 ( .A(data_in_1[115]), .B(n80), .Y(n646) );
  NAND2XL U497 ( .A(data_in_2[115]), .B(n90), .Y(n647) );
  NAND3X1 U498 ( .A(n544), .B(n543), .C(n542), .Y(data_out[81]) );
  NAND2XL U499 ( .A(R3[13]), .B(n267), .Y(n542) );
  NAND2XL U500 ( .A(data_in_1[81]), .B(n16), .Y(n543) );
  NAND2XL U501 ( .A(data_in_2[81]), .B(n93), .Y(n544) );
  NAND3X1 U502 ( .A(n547), .B(n546), .C(n545), .Y(data_out[82]) );
  NAND2XL U503 ( .A(R3[14]), .B(n267), .Y(n545) );
  NAND2XL U504 ( .A(data_in_1[82]), .B(n23), .Y(n546) );
  NAND2XL U505 ( .A(data_in_2[82]), .B(n87), .Y(n547) );
  NAND3X1 U506 ( .A(n650), .B(n649), .C(n648), .Y(data_out[116]) );
  NAND2XL U507 ( .A(R4[14]), .B(n265), .Y(n648) );
  NAND2XL U508 ( .A(data_in_1[116]), .B(n18), .Y(n649) );
  NAND2XL U509 ( .A(data_in_2[116]), .B(n90), .Y(n650) );
  NAND3X1 U510 ( .A(n701), .B(n700), .C(n699), .Y(data_out[133]) );
  NAND2XL U511 ( .A(R4[31]), .B(n264), .Y(n699) );
  NAND2XL U512 ( .A(data_in_1[133]), .B(n20), .Y(n700) );
  NAND2XL U513 ( .A(data_in_2[133]), .B(n86), .Y(n701) );
  NAND3X1 U514 ( .A(n653), .B(n652), .C(n651), .Y(data_out[117]) );
  NAND2XL U515 ( .A(R4[15]), .B(n265), .Y(n651) );
  NAND2XL U516 ( .A(data_in_1[117]), .B(n28), .Y(n652) );
  NAND2XL U517 ( .A(data_in_2[117]), .B(n94), .Y(n653) );
  NAND3X1 U518 ( .A(n598), .B(n597), .C(n596), .Y(data_out[99]) );
  NAND2XL U519 ( .A(data_in_1[99]), .B(n22), .Y(n597) );
  NAND2XL U520 ( .A(data_in_2[99]), .B(n85), .Y(n598) );
  NAND3X1 U521 ( .A(n705), .B(n704), .C(n703), .Y(data_out[134]) );
  NAND2XL U522 ( .A(data_in_2[134]), .B(n85), .Y(n705) );
  NAND3X1 U523 ( .A(n550), .B(n549), .C(n548), .Y(data_out[83]) );
  NAND2XL U524 ( .A(R3[15]), .B(n267), .Y(n548) );
  NAND2XL U525 ( .A(data_in_1[83]), .B(n26), .Y(n549) );
  NAND2XL U526 ( .A(data_in_2[83]), .B(n92), .Y(n550) );
  NAND3X1 U527 ( .A(n601), .B(n600), .C(n599), .Y(data_out[100]) );
  NAND2XL U528 ( .A(data_in_1[100]), .B(n24), .Y(n600) );
  NAND2XL U529 ( .A(data_in_2[100]), .B(n93), .Y(n601) );
  NAND3X1 U530 ( .A(n490), .B(n489), .C(n488), .Y(data_out[65]) );
  NAND2XL U531 ( .A(data_in_2[65]), .B(n94), .Y(n490) );
  NAND3X1 U532 ( .A(n437), .B(n436), .C(n435), .Y(data_out[48]) );
  NAND2XL U533 ( .A(R2[14]), .B(n268), .Y(n435) );
  NAND2XL U534 ( .A(data_in_1[48]), .B(n19), .Y(n436) );
  NAND2XL U535 ( .A(data_in_2[48]), .B(n88), .Y(n437) );
  NAND3X1 U536 ( .A(n493), .B(n492), .C(n491), .Y(data_out[66]) );
  NAND2XL U537 ( .A(data_in_2[66]), .B(n89), .Y(n493) );
  NAND3X1 U538 ( .A(n440), .B(n439), .C(n438), .Y(data_out[49]) );
  NAND2XL U539 ( .A(R2[15]), .B(n268), .Y(n438) );
  NAND2XL U540 ( .A(data_in_1[49]), .B(n29), .Y(n439) );
  NAND2XL U541 ( .A(data_in_2[49]), .B(n91), .Y(n440) );
  NAND3X1 U542 ( .A(n296), .B(n295), .C(n294), .Y(data_out[2]) );
  NAND2X1 U543 ( .A(R1[2]), .B(n269), .Y(n294) );
  NAND2XL U544 ( .A(data_in_1[2]), .B(n31), .Y(n295) );
  NAND2X1 U545 ( .A(data_in_2[2]), .B(n92), .Y(n296) );
  NAND3X1 U546 ( .A(n293), .B(n292), .C(n291), .Y(data_out[1]) );
  NAND2X1 U547 ( .A(R1[1]), .B(n269), .Y(n291) );
  NAND2X1 U548 ( .A(data_in_2[1]), .B(n86), .Y(n293) );
  NAND2XL U549 ( .A(data_in_1[1]), .B(n8), .Y(n292) );
  NAND3X1 U550 ( .A(n299), .B(n298), .C(n297), .Y(data_out[3]) );
  NAND2X1 U551 ( .A(R1[3]), .B(n269), .Y(n297) );
  NAND2XL U552 ( .A(data_in_1[3]), .B(n7), .Y(n298) );
  NAND2X1 U553 ( .A(data_in_2[3]), .B(n91), .Y(n299) );
  NAND3X1 U554 ( .A(n290), .B(n289), .C(n288), .Y(data_out[0]) );
  NAND2XL U555 ( .A(R1[0]), .B(n264), .Y(n288) );
  NAND2XL U556 ( .A(data_in_1[0]), .B(n38), .Y(n289) );
  NAND2XL U557 ( .A(data_in_2[0]), .B(n89), .Y(n290) );
  NAND3X1 U558 ( .A(n356), .B(n355), .C(n354), .Y(data_out[22]) );
  NAND2X1 U559 ( .A(R1[22]), .B(n269), .Y(n354) );
  NAND2X1 U560 ( .A(data_in_1[22]), .B(n37), .Y(n355) );
  NAND2X1 U561 ( .A(data_in_2[22]), .B(n94), .Y(n356) );
  NAND3X1 U562 ( .A(n344), .B(n343), .C(n342), .Y(data_out[18]) );
  NAND2X1 U563 ( .A(R1[18]), .B(n269), .Y(n342) );
  NAND2X1 U564 ( .A(data_in_1[18]), .B(n5), .Y(n343) );
  NAND2X1 U565 ( .A(data_in_2[18]), .B(n88), .Y(n344) );
  NAND3X1 U566 ( .A(n347), .B(n346), .C(n345), .Y(data_out[19]) );
  NAND2X1 U567 ( .A(R1[19]), .B(n266), .Y(n345) );
  NAND2X1 U568 ( .A(data_in_1[19]), .B(n4), .Y(n346) );
  NAND2X1 U569 ( .A(data_in_2[19]), .B(n90), .Y(n347) );
  NAND3X1 U570 ( .A(n341), .B(n340), .C(n339), .Y(data_out[17]) );
  NAND2X1 U571 ( .A(R1[17]), .B(n266), .Y(n339) );
  NAND2X1 U572 ( .A(data_in_1[17]), .B(n32), .Y(n340) );
  NAND2X1 U573 ( .A(data_in_2[17]), .B(n87), .Y(n341) );
  NAND3X1 U574 ( .A(n350), .B(n349), .C(n348), .Y(data_out[20]) );
  NAND2X1 U575 ( .A(R1[20]), .B(n266), .Y(n348) );
  NAND2X1 U576 ( .A(data_in_1[20]), .B(n30), .Y(n349) );
  NAND2X1 U577 ( .A(data_in_2[20]), .B(n93), .Y(n350) );
  NAND3X1 U578 ( .A(n302), .B(n301), .C(n300), .Y(data_out[4]) );
  NAND2X1 U579 ( .A(R1[4]), .B(n266), .Y(n300) );
  NAND2XL U580 ( .A(data_in_1[4]), .B(n40), .Y(n301) );
  NAND2X1 U581 ( .A(data_in_2[4]), .B(n87), .Y(n302) );
  NAND3X1 U582 ( .A(n305), .B(n304), .C(n303), .Y(data_out[5]) );
  NAND2X1 U583 ( .A(R1[5]), .B(n270), .Y(n303) );
  NAND2XL U584 ( .A(data_in_1[5]), .B(n39), .Y(n304) );
  NAND2X1 U585 ( .A(data_in_2[5]), .B(n91), .Y(n305) );
  NAND3X1 U586 ( .A(n314), .B(n313), .C(n312), .Y(data_out[8]) );
  NAND2X1 U587 ( .A(R1[8]), .B(n265), .Y(n312) );
  NAND2XL U588 ( .A(data_in_1[8]), .B(n46), .Y(n313) );
  NAND2X1 U589 ( .A(data_in_2[8]), .B(n93), .Y(n314) );
  NAND3X1 U590 ( .A(n311), .B(n310), .C(n309), .Y(data_out[7]) );
  NAND2X1 U591 ( .A(R1[7]), .B(n270), .Y(n309) );
  NAND2XL U592 ( .A(data_in_1[7]), .B(n44), .Y(n310) );
  NAND2X1 U593 ( .A(data_in_2[7]), .B(n90), .Y(n311) );
  NAND3X1 U594 ( .A(n308), .B(n307), .C(n306), .Y(data_out[6]) );
  NAND2X1 U595 ( .A(R1[6]), .B(n269), .Y(n306) );
  NAND2X1 U596 ( .A(data_in_1[6]), .B(n42), .Y(n307) );
  NAND2X1 U597 ( .A(data_in_2[6]), .B(n88), .Y(n308) );
  NAND3X1 U598 ( .A(n317), .B(n316), .C(n315), .Y(data_out[9]) );
  NAND2X1 U599 ( .A(R1[9]), .B(n268), .Y(n315) );
  NAND2X1 U600 ( .A(data_in_1[9]), .B(n48), .Y(n316) );
  NAND2X1 U601 ( .A(data_in_2[9]), .B(n92), .Y(n317) );
  NAND3X1 U602 ( .A(n362), .B(n361), .C(n360), .Y(data_out[24]) );
  NAND2X1 U603 ( .A(R1[24]), .B(n266), .Y(n360) );
  NAND2X1 U604 ( .A(data_in_1[24]), .B(n45), .Y(n361) );
  NAND2X1 U605 ( .A(data_in_2[24]), .B(n89), .Y(n362) );
  NAND3X1 U606 ( .A(n365), .B(n364), .C(n363), .Y(data_out[25]) );
  NAND2X1 U607 ( .A(R1[25]), .B(n269), .Y(n363) );
  NAND2XL U608 ( .A(data_in_1[25]), .B(n47), .Y(n364) );
  NAND2X1 U609 ( .A(data_in_2[25]), .B(n94), .Y(n365) );
  NAND3X1 U610 ( .A(n353), .B(n352), .C(n351), .Y(data_out[21]) );
  NAND2X1 U611 ( .A(R1[21]), .B(n269), .Y(n351) );
  NAND2XL U612 ( .A(data_in_1[21]), .B(n41), .Y(n352) );
  NAND2X1 U613 ( .A(data_in_2[21]), .B(n85), .Y(n353) );
  NAND3X1 U614 ( .A(n359), .B(n358), .C(n357), .Y(data_out[23]) );
  NAND2XL U615 ( .A(R1[23]), .B(n269), .Y(n357) );
  NAND2XL U616 ( .A(data_in_1[23]), .B(n43), .Y(n358) );
  NAND2X1 U617 ( .A(data_in_2[23]), .B(n86), .Y(n359) );
  NAND3X1 U618 ( .A(n368), .B(n367), .C(n366), .Y(data_out[26]) );
  NAND2X1 U619 ( .A(R1[26]), .B(n265), .Y(n366) );
  NAND2XL U620 ( .A(data_in_1[26]), .B(n49), .Y(n367) );
  NAND2X1 U621 ( .A(data_in_2[26]), .B(n85), .Y(n368) );
  NAND3X1 U622 ( .A(n320), .B(n319), .C(n318), .Y(data_out[10]) );
  NAND2X1 U623 ( .A(R1[10]), .B(n265), .Y(n318) );
  NAND2XL U624 ( .A(data_in_1[10]), .B(n53), .Y(n319) );
  NAND2X1 U625 ( .A(data_in_2[10]), .B(n88), .Y(n320) );
  NAND3X1 U626 ( .A(n371), .B(n370), .C(n369), .Y(data_out[27]) );
  NAND2XL U627 ( .A(R1[27]), .B(n269), .Y(n369) );
  NAND2XL U628 ( .A(data_in_1[27]), .B(n52), .Y(n370) );
  NAND2X1 U629 ( .A(data_in_2[27]), .B(n86), .Y(n371) );
  NAND3X1 U630 ( .A(n383), .B(n382), .C(n381), .Y(data_out[31]) );
  NAND2XL U631 ( .A(R1[31]), .B(n269), .Y(n381) );
  NAND2X1 U632 ( .A(data_in_2[31]), .B(n93), .Y(n383) );
  NAND2XL U633 ( .A(data_in_1[31]), .B(n64), .Y(n382) );
  NAND3X1 U634 ( .A(n374), .B(n373), .C(n372), .Y(data_out[28]) );
  NAND2X1 U635 ( .A(R1[28]), .B(n270), .Y(n372) );
  NAND2X1 U636 ( .A(data_in_2[28]), .B(n90), .Y(n374) );
  NAND2XL U637 ( .A(data_in_1[28]), .B(n54), .Y(n373) );
  INVX1 U638 ( .A(data_in_2[30]), .Y(n378) );
  NAND3X1 U639 ( .A(n326), .B(n325), .C(n324), .Y(data_out[12]) );
  NAND2X1 U640 ( .A(R1[12]), .B(n265), .Y(n324) );
  NAND2X1 U641 ( .A(data_in_2[12]), .B(n89), .Y(n326) );
  NAND2X1 U642 ( .A(data_in_1[12]), .B(n55), .Y(n325) );
  NAND3X1 U643 ( .A(n377), .B(n376), .C(n375), .Y(data_out[29]) );
  NAND2XL U644 ( .A(R1[29]), .B(n269), .Y(n375) );
  NAND2XL U645 ( .A(data_in_1[29]), .B(n56), .Y(n376) );
  NAND2X1 U646 ( .A(data_in_2[29]), .B(n91), .Y(n377) );
  NAND3X1 U647 ( .A(n335), .B(n334), .C(n333), .Y(data_out[15]) );
  NAND2X1 U648 ( .A(R1[15]), .B(n267), .Y(n333) );
  NAND2X1 U649 ( .A(data_in_1[15]), .B(n63), .Y(n334) );
  NAND2X1 U650 ( .A(data_in_2[15]), .B(n94), .Y(n335) );
  NAND3X1 U651 ( .A(n386), .B(n385), .C(n384), .Y(data_out[32]) );
  NAND2XL U652 ( .A(R1[32]), .B(n269), .Y(n384) );
  NAND2XL U653 ( .A(data_in_1[32]), .B(n65), .Y(n385) );
  NAND2XL U654 ( .A(data_in_2[32]), .B(n86), .Y(n386) );
  NAND3X1 U655 ( .A(n323), .B(n322), .C(n321), .Y(data_out[11]) );
  NAND2X1 U656 ( .A(R1[11]), .B(n269), .Y(n321) );
  NAND2X1 U657 ( .A(data_in_1[11]), .B(n51), .Y(n322) );
  NAND2X1 U658 ( .A(data_in_2[11]), .B(n87), .Y(n323) );
  NAND3X1 U659 ( .A(n332), .B(n331), .C(n330), .Y(data_out[14]) );
  NAND2X1 U660 ( .A(R1[14]), .B(n268), .Y(n330) );
  NAND2X1 U661 ( .A(data_in_1[14]), .B(n61), .Y(n331) );
  NAND2X1 U662 ( .A(data_in_2[14]), .B(n92), .Y(n332) );
  NAND3X1 U663 ( .A(n161), .B(n329), .C(n328), .Y(data_out[13]) );
  OR2XL U664 ( .A(n84), .B(n327), .Y(n161) );
  NAND3X1 U665 ( .A(n389), .B(n388), .C(n387), .Y(data_out[33]) );
  NAND2XL U666 ( .A(R1[33]), .B(n269), .Y(n387) );
  NAND2XL U667 ( .A(data_in_1[33]), .B(n67), .Y(n388) );
  NAND2XL U668 ( .A(data_in_2[33]), .B(n87), .Y(n389) );
  NAND3X1 U669 ( .A(n338), .B(n337), .C(n336), .Y(data_out[16]) );
  NAND2X1 U670 ( .A(R1[16]), .B(n266), .Y(n336) );
  NAND2XL U671 ( .A(data_in_1[16]), .B(n66), .Y(n337) );
  NAND2X1 U672 ( .A(data_in_2[16]), .B(n85), .Y(n338) );
  INVX1 U673 ( .A(data_in_2[13]), .Y(n327) );
  NOR2X1 U674 ( .A(n720), .B(n282), .Y(n281) );
  INVXL U675 ( .A(counter[2]), .Y(n720) );
  INVX1 U676 ( .A(n285), .Y(n275) );
  OR2XL U677 ( .A(n140), .B(n141), .Y(n162) );
  NAND3XL U678 ( .A(data_in_2[86]), .B(n710), .C(n283), .Y(n562) );
  INVX8 U679 ( .A(n287), .Y(n390) );
  NOR2X1 U680 ( .A(n501), .B(n500), .Y(n502) );
  NAND2BX4 U681 ( .AN(n242), .B(n390), .Y(n665) );
  OAI2BB2XL U682 ( .B0(n84), .B1(n378), .A0N(data_in_1[30]), .A1N(n62), .Y(
        n380) );
  NAND3XL U683 ( .A(n283), .B(data_in_2[121]), .C(n665), .Y(n667) );
  NAND3XL U684 ( .A(n280), .B(data_in_2[87]), .C(n665), .Y(n565) );
  NOR2XL U685 ( .A(n708), .B(n498), .Y(n501) );
  NOR2X1 U686 ( .A(n708), .B(n499), .Y(n500) );
  XOR2X1 U687 ( .A(counter[3]), .B(n281), .Y(N8) );
  NOR4BXL U688 ( .AN(counter[1]), .B(n720), .C(n286), .D(n83), .Y(n285) );
  NAND2XL U689 ( .A(counter[1]), .B(n83), .Y(n282) );
  NAND3XL U690 ( .A(data_in_1[87]), .B(n278), .C(n665), .Y(n564) );
  NAND3XL U691 ( .A(data_in_1[121]), .B(n278), .C(n665), .Y(n668) );
  NAND2XL U692 ( .A(data_in_1[70]), .B(n278), .Y(n507) );
  NAND3XL U693 ( .A(data_in_1[119]), .B(n278), .C(n659), .Y(n661) );
  NAND2XL U694 ( .A(data_in_1[102]), .B(n278), .Y(n606) );
  NAND2XL U695 ( .A(data_in_1[68]), .B(n278), .Y(n499) );
  NAND2XL U696 ( .A(data_in_1[85]), .B(n278), .Y(n555) );
  NAND2X1 U697 ( .A(data_in_1[67]), .B(n278), .Y(n494) );
  NAND3BX4 U698 ( .AN(counter[2]), .B(n286), .C(counter[1]), .Y(n287) );
  OAI2BB1X4 U699 ( .A0N(R2[0]), .A1N(n614), .B0(n393), .Y(data_out[34]) );
  OAI2BB1X4 U700 ( .A0N(R2[1]), .A1N(n270), .B0(n398), .Y(data_out[35]) );
  NAND2X4 U701 ( .A(data_in_2[36]), .B(n89), .Y(n401) );
  NAND2X4 U702 ( .A(R2[2]), .B(n269), .Y(n399) );
  NAND3X4 U703 ( .A(n401), .B(n400), .C(n399), .Y(data_out[36]) );
  OAI2BB1X4 U704 ( .A0N(R2[17]), .A1N(n559), .B0(n449), .Y(data_out[51]) );
  AOI21X4 U705 ( .A0(data_in_2[53]), .A1(n88), .B0(n453), .Y(n454) );
  OAI2BB1X4 U706 ( .A0N(data_in_1[53]), .A1N(n15), .B0(n454), .Y(data_out[53])
         );
  NAND2X4 U707 ( .A(data_in_2[54]), .B(n94), .Y(n457) );
  NAND3X4 U708 ( .A(n457), .B(n456), .C(n455), .Y(data_out[54]) );
  OAI2BB1X4 U709 ( .A0N(R3[0]), .A1N(n614), .B0(n502), .Y(data_out[68]) );
  OAI2BB1X4 U710 ( .A0N(n506), .A1N(n251), .B0(n505), .Y(data_out[69]) );
  OAI2BB1X4 U711 ( .A0N(n558), .A1N(n251), .B0(n557), .Y(data_out[85]) );
  NAND3X4 U712 ( .A(n562), .B(n561), .C(n560), .Y(data_out[86]) );
  NAND2X4 U713 ( .A(R3[19]), .B(n267), .Y(n563) );
  NAND3X4 U714 ( .A(n565), .B(n564), .C(n563), .Y(data_out[87]) );
  OAI2BB1X4 U715 ( .A0N(R4[0]), .A1N(n614), .B0(n610), .Y(data_out[102]) );
  NAND3X4 U716 ( .A(n613), .B(n612), .C(n611), .Y(data_out[103]) );
endmodule


module multi16_11_DW01_add_0 ( A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, 
        A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, 
        B_20_, B_19_, B_18_, B_17_, B_16_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, 
        SUM_17_, SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, 
        SUM_9_, SUM_8_, SUM_7_, SUM_6_, SUM_5_ );
  input A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_,
         A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, B_20_, B_19_,
         B_18_, B_17_, B_16_;
  output SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, SUM_15_,
         SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, SUM_7_,
         SUM_6_, SUM_5_;
  wire   n1, n2, n3, n4, n5, n7, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44;

  INVX4 U2 ( .A(n24), .Y(SUM_15_) );
  AOI21X2 U3 ( .A0(n23), .A1(n22), .B0(n21), .Y(n42) );
  INVX4 U4 ( .A(n38), .Y(n23) );
  OAI21X1 U5 ( .A0(n42), .A1(n35), .B0(n37), .Y(n40) );
  BUFX3 U6 ( .A(A_14_), .Y(SUM_14_) );
  CLKINVX3 U7 ( .A(n39), .Y(n21) );
  NOR2X1 U8 ( .A(B_18_), .B(A_18_), .Y(n35) );
  XOR2X1 U9 ( .A(n40), .B(n41), .Y(SUM_19_) );
  NOR2BX1 U10 ( .AN(n33), .B(n32), .Y(n41) );
  NAND2X2 U11 ( .A(B_17_), .B(A_17_), .Y(n39) );
  NAND2X2 U12 ( .A(B_16_), .B(A_16_), .Y(n38) );
  INVX1 U13 ( .A(n35), .Y(n19) );
  NOR2X2 U14 ( .A(B_17_), .B(A_17_), .Y(n34) );
  NOR2X1 U15 ( .A(B_17_), .B(A_17_), .Y(n5) );
  NAND2X1 U16 ( .A(n3), .B(n4), .Y(SUM_18_) );
  OAI21X1 U17 ( .A0(n31), .A1(n32), .B0(n33), .Y(n27) );
  AOI21XL U18 ( .A0(n19), .A1(n36), .B0(n20), .Y(n31) );
  INVXL U19 ( .A(n43), .Y(n1) );
  NOR2X2 U20 ( .A(B_16_), .B(A_16_), .Y(n7) );
  NOR2BX4 U21 ( .AN(n38), .B(n7), .Y(SUM_16_) );
  INVX1 U22 ( .A(n42), .Y(n2) );
  NAND2XL U23 ( .A(n1), .B(n42), .Y(n4) );
  INVX1 U24 ( .A(n5), .Y(n22) );
  NAND2X1 U25 ( .A(B_19_), .B(A_19_), .Y(n33) );
  NOR2X1 U26 ( .A(B_19_), .B(A_19_), .Y(n32) );
  NAND2X1 U27 ( .A(n43), .B(n2), .Y(n3) );
  XOR2X4 U28 ( .A(n23), .B(n44), .Y(SUM_17_) );
  INVX2 U29 ( .A(A_15_), .Y(n24) );
  INVXL U30 ( .A(n29), .Y(n18) );
  BUFX3 U31 ( .A(A_13_), .Y(SUM_13_) );
  BUFX3 U32 ( .A(A_12_), .Y(SUM_12_) );
  BUFX3 U33 ( .A(A_11_), .Y(SUM_11_) );
  BUFX3 U34 ( .A(A_10_), .Y(SUM_10_) );
  BUFX3 U35 ( .A(A_9_), .Y(SUM_9_) );
  BUFX3 U36 ( .A(A_8_), .Y(SUM_8_) );
  BUFX3 U37 ( .A(A_7_), .Y(SUM_7_) );
  BUFX3 U38 ( .A(A_6_), .Y(SUM_6_) );
  BUFX3 U39 ( .A(A_5_), .Y(SUM_5_) );
  INVXL U40 ( .A(n37), .Y(n20) );
  NOR2X4 U41 ( .A(n34), .B(n21), .Y(n44) );
  XOR2X1 U42 ( .A(n25), .B(n26), .Y(SUM_21_) );
  AOI21X1 U43 ( .A0(n27), .A1(n28), .B0(n18), .Y(n26) );
  XNOR2X1 U44 ( .A(B_21_), .B(A_21_), .Y(n25) );
  XNOR2X1 U45 ( .A(n30), .B(n27), .Y(SUM_20_) );
  OAI21XL U46 ( .A0(n34), .A1(n38), .B0(n39), .Y(n36) );
  NAND2X1 U47 ( .A(n29), .B(n28), .Y(n30) );
  OR2X1 U48 ( .A(B_20_), .B(A_20_), .Y(n28) );
  NAND2X1 U49 ( .A(B_20_), .B(A_20_), .Y(n29) );
  NAND2X1 U50 ( .A(n37), .B(n19), .Y(n43) );
  NAND2X1 U51 ( .A(B_18_), .B(A_18_), .Y(n37) );
endmodule


module multi16_11_DW02_mult_0 ( A, B, PRODUCT_23_, PRODUCT_22_, PRODUCT_21_, 
        PRODUCT_20_, PRODUCT_19_, PRODUCT_18_, PRODUCT_17_, PRODUCT_16_, 
        PRODUCT_15_, PRODUCT_14_, PRODUCT_13_, PRODUCT_12_, PRODUCT_11_, 
        PRODUCT_10_, PRODUCT_9_, PRODUCT_8_, PRODUCT_7_ );
  input [16:0] A;
  input [7:0] B;
  output PRODUCT_23_, PRODUCT_22_, PRODUCT_21_, PRODUCT_20_, PRODUCT_19_,
         PRODUCT_18_, PRODUCT_17_, PRODUCT_16_, PRODUCT_15_, PRODUCT_14_,
         PRODUCT_13_, PRODUCT_12_, PRODUCT_11_, PRODUCT_10_, PRODUCT_9_,
         PRODUCT_8_, PRODUCT_7_;
  wire   ab_16__7_, ab_16__6_, ab_16__5_, ab_16__4_, ab_16__3_, ab_16__2_,
         ab_16__1_, ab_16__0_, ab_15__7_, ab_15__6_, ab_15__5_, ab_15__4_,
         ab_15__3_, ab_15__2_, ab_15__1_, ab_15__0_, ab_14__7_, ab_14__6_,
         ab_14__5_, ab_14__4_, ab_14__3_, ab_14__2_, ab_14__1_, ab_14__0_,
         ab_13__7_, ab_13__6_, ab_13__5_, ab_13__4_, ab_13__3_, ab_13__2_,
         ab_13__1_, ab_13__0_, ab_12__7_, ab_12__6_, ab_12__5_, ab_12__4_,
         ab_12__3_, ab_12__2_, ab_12__1_, ab_12__0_, ab_11__7_, ab_11__6_,
         ab_11__5_, ab_11__4_, ab_11__3_, ab_11__2_, ab_11__1_, ab_11__0_,
         ab_10__7_, ab_10__6_, ab_10__5_, ab_10__4_, ab_10__3_, ab_10__2_,
         ab_10__1_, ab_10__0_, ab_9__7_, ab_9__6_, ab_9__5_, ab_9__4_,
         ab_9__3_, ab_9__2_, ab_9__1_, ab_9__0_, ab_8__7_, ab_8__6_, ab_8__5_,
         ab_8__4_, ab_8__3_, ab_8__2_, ab_8__1_, ab_8__0_, ab_7__7_, ab_7__6_,
         ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_, ab_7__0_, ab_6__7_,
         ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_, ab_6__1_, ab_6__0_,
         ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_, ab_5__2_, ab_5__1_,
         ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_, ab_4__3_, ab_4__2_,
         ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_, ab_3__4_, ab_3__3_,
         ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_, ab_2__5_, ab_2__4_,
         ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_, ab_1__6_, ab_1__5_,
         ab_1__4_, ab_1__3_, ab_1__2_, ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_,
         ab_0__3_, ab_0__2_, CARRYB_16__6_, CARRYB_16__5_, CARRYB_16__4_,
         CARRYB_16__3_, CARRYB_16__2_, CARRYB_16__1_, CARRYB_16__0_,
         CARRYB_15__6_, CARRYB_15__5_, CARRYB_15__4_, CARRYB_15__3_,
         CARRYB_15__2_, CARRYB_15__1_, CARRYB_15__0_, CARRYB_14__6_,
         CARRYB_14__5_, CARRYB_14__4_, CARRYB_14__3_, CARRYB_14__2_,
         CARRYB_14__1_, CARRYB_14__0_, CARRYB_13__6_, CARRYB_13__5_,
         CARRYB_13__4_, CARRYB_13__3_, CARRYB_13__2_, CARRYB_13__1_,
         CARRYB_13__0_, CARRYB_12__6_, CARRYB_12__5_, CARRYB_12__4_,
         CARRYB_12__3_, CARRYB_12__2_, CARRYB_12__1_, CARRYB_12__0_,
         CARRYB_11__6_, CARRYB_11__5_, CARRYB_11__4_, CARRYB_11__3_,
         CARRYB_11__2_, CARRYB_11__1_, CARRYB_11__0_, CARRYB_10__6_,
         CARRYB_10__5_, CARRYB_10__4_, CARRYB_10__3_, CARRYB_10__2_,
         CARRYB_10__1_, CARRYB_10__0_, CARRYB_9__6_, CARRYB_9__5_,
         CARRYB_9__4_, CARRYB_9__3_, CARRYB_9__2_, CARRYB_9__1_, CARRYB_9__0_,
         CARRYB_8__6_, CARRYB_8__5_, CARRYB_8__4_, CARRYB_8__3_, CARRYB_8__2_,
         CARRYB_8__1_, CARRYB_8__0_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_,
         CARRYB_7__3_, CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_,
         CARRYB_6__5_, CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_,
         CARRYB_6__0_, CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_,
         CARRYB_5__2_, CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_,
         CARRYB_4__4_, CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_,
         CARRYB_3__6_, CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_,
         CARRYB_3__1_, CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_,
         CARRYB_2__3_, CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__6_,
         CARRYB_1__5_, CARRYB_1__0_, SUMB_16__6_, SUMB_16__5_, SUMB_16__4_,
         SUMB_16__3_, SUMB_16__2_, SUMB_16__1_, SUMB_16__0_, SUMB_15__6_,
         SUMB_15__5_, SUMB_15__4_, SUMB_15__3_, SUMB_15__2_, SUMB_15__1_,
         SUMB_14__6_, SUMB_14__5_, SUMB_14__4_, SUMB_14__3_, SUMB_14__2_,
         SUMB_14__1_, SUMB_13__6_, SUMB_13__5_, SUMB_13__4_, SUMB_13__3_,
         SUMB_13__2_, SUMB_13__1_, SUMB_12__6_, SUMB_12__5_, SUMB_12__4_,
         SUMB_12__3_, SUMB_12__2_, SUMB_12__1_, SUMB_11__6_, SUMB_11__5_,
         SUMB_11__4_, SUMB_11__3_, SUMB_11__2_, SUMB_11__1_, SUMB_10__6_,
         SUMB_10__5_, SUMB_10__4_, SUMB_10__3_, SUMB_10__2_, SUMB_10__1_,
         SUMB_9__6_, SUMB_9__5_, SUMB_9__4_, SUMB_9__3_, SUMB_9__2_,
         SUMB_9__1_, SUMB_8__6_, SUMB_8__5_, SUMB_8__4_, SUMB_8__3_,
         SUMB_8__2_, SUMB_8__1_, SUMB_7__6_, SUMB_7__5_, SUMB_7__4_,
         SUMB_7__3_, SUMB_7__2_, SUMB_7__1_, SUMB_6__6_, SUMB_6__5_,
         SUMB_6__4_, SUMB_6__3_, SUMB_6__2_, SUMB_6__1_, SUMB_5__6_,
         SUMB_5__5_, SUMB_5__4_, SUMB_5__3_, SUMB_5__2_, SUMB_5__1_,
         SUMB_4__6_, SUMB_4__5_, SUMB_4__4_, SUMB_4__3_, SUMB_4__2_,
         SUMB_4__1_, SUMB_3__6_, SUMB_3__5_, SUMB_3__4_, SUMB_3__3_,
         SUMB_3__2_, SUMB_3__1_, SUMB_2__6_, SUMB_2__5_, SUMB_2__4_,
         SUMB_2__3_, SUMB_2__2_, SUMB_2__1_, SUMB_1__6_, SUMB_1__5_,
         SUMB_1__4_, SUMB_1__3_, SUMB_1__2_, SUMB_1__1_, PROD1_7_, A1_21_,
         A1_20_, A1_19_, A1_18_, A1_17_, A1_16_, A1_15_, A1_13_, A1_12_,
         A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, A1_4_, A1_3_, A1_2_,
         A1_1_, A1_0_, n3, n4, n5, n6, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80;

  ADDFHX4 S2_14_1 ( .A(ab_14__1_), .B(CARRYB_13__1_), .CI(SUMB_13__2_), .CO(
        CARRYB_14__1_), .S(SUMB_14__1_) );
  ADDFHX4 S1_13_0 ( .A(ab_13__0_), .B(CARRYB_12__0_), .CI(SUMB_12__1_), .CO(
        CARRYB_13__0_), .S(A1_11_) );
  ADDFHX4 S2_13_1 ( .A(ab_13__1_), .B(CARRYB_12__1_), .CI(SUMB_12__2_), .CO(
        CARRYB_13__1_), .S(SUMB_13__1_) );
  ADDFHX4 S1_12_0 ( .A(ab_12__0_), .B(CARRYB_11__0_), .CI(SUMB_11__1_), .CO(
        CARRYB_12__0_), .S(A1_10_) );
  ADDFHX4 S2_11_1 ( .A(ab_11__1_), .B(CARRYB_10__1_), .CI(SUMB_10__2_), .CO(
        CARRYB_11__1_), .S(SUMB_11__1_) );
  ADDFHX4 S2_10_2 ( .A(ab_10__2_), .B(CARRYB_9__2_), .CI(SUMB_9__3_), .CO(
        CARRYB_10__2_), .S(SUMB_10__2_) );
  multi16_11_DW01_add_0 FS_1 ( .A_21_(A1_21_), .A_20_(A1_20_), .A_19_(A1_19_), 
        .A_18_(A1_18_), .A_17_(A1_17_), .A_16_(A1_16_), .A_15_(A1_15_), 
        .A_14_(SUMB_16__0_), .A_13_(A1_13_), .A_12_(A1_12_), .A_11_(A1_11_), 
        .A_10_(A1_10_), .A_9_(A1_9_), .A_8_(A1_8_), .A_7_(A1_7_), .A_6_(A1_6_), 
        .A_5_(PROD1_7_), .B_21_(n60), .B_20_(n59), .B_19_(n56), .B_18_(n58), 
        .B_17_(n55), .B_16_(n57), .SUM_21_(PRODUCT_23_), .SUM_20_(PRODUCT_22_), 
        .SUM_19_(PRODUCT_21_), .SUM_18_(PRODUCT_20_), .SUM_17_(PRODUCT_19_), 
        .SUM_16_(PRODUCT_18_), .SUM_15_(PRODUCT_17_), .SUM_14_(PRODUCT_16_), 
        .SUM_13_(PRODUCT_15_), .SUM_12_(PRODUCT_14_), .SUM_11_(PRODUCT_13_), 
        .SUM_10_(PRODUCT_12_), .SUM_9_(PRODUCT_11_), .SUM_8_(PRODUCT_10_), 
        .SUM_7_(PRODUCT_9_), .SUM_6_(PRODUCT_8_), .SUM_5_(PRODUCT_7_) );
  ADDFHX1 S3_15_6 ( .A(ab_15__6_), .B(CARRYB_14__6_), .CI(ab_14__7_), .CO(
        CARRYB_15__6_), .S(SUMB_15__6_) );
  ADDFHX2 S4_0 ( .A(ab_16__0_), .B(CARRYB_15__0_), .CI(SUMB_15__1_), .CO(
        CARRYB_16__0_), .S(SUMB_16__0_) );
  ADDFX2 S5_6 ( .A(ab_16__6_), .B(CARRYB_15__6_), .CI(ab_15__7_), .CO(
        CARRYB_16__6_), .S(SUMB_16__6_) );
  ADDFHX1 S4_5 ( .A(ab_16__5_), .B(CARRYB_15__5_), .CI(SUMB_15__6_), .CO(
        CARRYB_16__5_), .S(SUMB_16__5_) );
  ADDFHX4 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  ADDFHX4 S3_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(ab_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  ADDFHX2 S2_15_4 ( .A(ab_15__4_), .B(CARRYB_14__4_), .CI(SUMB_14__5_), .CO(
        CARRYB_15__4_), .S(SUMB_15__4_) );
  ADDFHX2 S4_4 ( .A(ab_16__4_), .B(CARRYB_15__4_), .CI(SUMB_15__5_), .CO(
        CARRYB_16__4_), .S(SUMB_16__4_) );
  ADDFHX2 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  ADDFHX2 S4_1 ( .A(ab_16__1_), .B(CARRYB_15__1_), .CI(SUMB_15__2_), .CO(
        CARRYB_16__1_), .S(SUMB_16__1_) );
  ADDFHX4 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  ADDFHX2 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  ADDFHX2 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  ADDFHX4 S2_8_3 ( .A(ab_8__3_), .B(CARRYB_7__3_), .CI(SUMB_7__4_), .CO(
        CARRYB_8__3_), .S(SUMB_8__3_) );
  ADDFHX4 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  ADDFHX2 S2_11_5 ( .A(ab_11__5_), .B(CARRYB_10__5_), .CI(SUMB_10__6_), .CO(
        CARRYB_11__5_), .S(SUMB_11__5_) );
  ADDFHX4 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  ADDFHX4 S2_9_1 ( .A(ab_9__1_), .B(CARRYB_8__1_), .CI(SUMB_8__2_), .CO(
        CARRYB_9__1_), .S(SUMB_9__1_) );
  ADDFHX4 S2_10_1 ( .A(ab_10__1_), .B(CARRYB_9__1_), .CI(SUMB_9__2_), .CO(
        CARRYB_10__1_), .S(SUMB_10__1_) );
  ADDFHX4 S1_8_0 ( .A(ab_8__0_), .B(CARRYB_7__0_), .CI(SUMB_7__1_), .CO(
        CARRYB_8__0_), .S(A1_6_) );
  ADDFHX4 S2_7_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  ADDFHX2 S2_14_5 ( .A(ab_14__5_), .B(CARRYB_13__5_), .CI(SUMB_13__6_), .CO(
        CARRYB_14__5_), .S(SUMB_14__5_) );
  ADDFHX2 S2_15_5 ( .A(ab_15__5_), .B(CARRYB_14__5_), .CI(SUMB_14__6_), .CO(
        CARRYB_15__5_), .S(SUMB_15__5_) );
  ADDFHX4 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  ADDFHX4 S2_11_3 ( .A(ab_11__3_), .B(CARRYB_10__3_), .CI(SUMB_10__4_), .CO(
        CARRYB_11__3_), .S(SUMB_11__3_) );
  ADDFHX2 S3_12_6 ( .A(ab_12__6_), .B(CARRYB_11__6_), .CI(ab_11__7_), .CO(
        CARRYB_12__6_), .S(SUMB_12__6_) );
  ADDFHX4 S2_12_3 ( .A(ab_12__3_), .B(CARRYB_11__3_), .CI(SUMB_11__4_), .CO(
        CARRYB_12__3_), .S(SUMB_12__3_) );
  ADDFHX4 S2_13_2 ( .A(ab_13__2_), .B(SUMB_12__3_), .CI(CARRYB_12__2_), .CO(
        CARRYB_13__2_), .S(SUMB_13__2_) );
  ADDFHX4 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  ADDFHX4 S2_12_5 ( .A(ab_12__5_), .B(CARRYB_11__5_), .CI(SUMB_11__6_), .CO(
        CARRYB_12__5_), .S(SUMB_12__5_) );
  ADDFHX4 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  ADDFHX2 S2_2_2 ( .A(ab_2__2_), .B(n10), .CI(SUMB_1__3_), .CO(CARRYB_2__2_), 
        .S(SUMB_2__2_) );
  ADDFHX4 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  ADDFHX4 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  ADDFHX4 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  ADDFHX4 S2_14_3 ( .A(ab_14__3_), .B(CARRYB_13__3_), .CI(SUMB_13__4_), .CO(
        CARRYB_14__3_), .S(SUMB_14__3_) );
  ADDFHX4 S2_14_2 ( .A(ab_14__2_), .B(CARRYB_13__2_), .CI(SUMB_13__3_), .CO(
        CARRYB_14__2_), .S(SUMB_14__2_) );
  ADDFHX4 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  ADDFHX4 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  ADDFHX4 S2_9_5 ( .A(ab_9__5_), .B(CARRYB_8__5_), .CI(SUMB_8__6_), .CO(
        CARRYB_9__5_), .S(SUMB_9__5_) );
  ADDFHX4 S2_10_4 ( .A(ab_10__4_), .B(CARRYB_9__4_), .CI(SUMB_9__5_), .CO(
        CARRYB_10__4_), .S(SUMB_10__4_) );
  ADDFHX4 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  ADDFHX4 S2_8_4 ( .A(ab_8__4_), .B(CARRYB_7__4_), .CI(SUMB_7__5_), .CO(
        CARRYB_8__4_), .S(SUMB_8__4_) );
  ADDFHX4 S2_2_1 ( .A(ab_2__1_), .B(n8), .CI(SUMB_1__2_), .CO(CARRYB_2__1_), 
        .S(SUMB_2__1_) );
  ADDFHX4 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  ADDFHX4 S4_3 ( .A(ab_16__3_), .B(CARRYB_15__3_), .CI(SUMB_15__4_), .CO(
        CARRYB_16__3_), .S(SUMB_16__3_) );
  ADDFHX4 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  ADDFHX2 S2_2_3 ( .A(ab_2__3_), .B(n11), .CI(SUMB_1__4_), .CO(CARRYB_2__3_), 
        .S(SUMB_2__3_) );
  ADDFHX2 S3_11_6 ( .A(ab_11__6_), .B(CARRYB_10__6_), .CI(ab_10__7_), .CO(
        CARRYB_11__6_), .S(SUMB_11__6_) );
  ADDFHX2 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  ADDFHX2 S2_13_5 ( .A(ab_13__5_), .B(CARRYB_12__5_), .CI(SUMB_12__6_), .CO(
        CARRYB_13__5_), .S(SUMB_13__5_) );
  ADDFHX2 S2_15_3 ( .A(ab_15__3_), .B(CARRYB_14__3_), .CI(SUMB_14__4_), .CO(
        CARRYB_15__3_), .S(SUMB_15__3_) );
  ADDFHX2 S2_15_1 ( .A(ab_15__1_), .B(CARRYB_14__1_), .CI(SUMB_14__2_), .CO(
        CARRYB_15__1_), .S(SUMB_15__1_) );
  ADDFHX2 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  ADDFHX2 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  ADDFHX2 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  ADDFHX2 S1_11_0 ( .A(ab_11__0_), .B(CARRYB_10__0_), .CI(SUMB_10__1_), .CO(
        CARRYB_11__0_), .S(A1_9_) );
  ADDFHX2 S3_8_6 ( .A(ab_8__6_), .B(CARRYB_7__6_), .CI(ab_7__7_), .CO(
        CARRYB_8__6_), .S(SUMB_8__6_) );
  ADDFHX2 S2_11_4 ( .A(ab_11__4_), .B(CARRYB_10__4_), .CI(SUMB_10__5_), .CO(
        CARRYB_11__4_), .S(SUMB_11__4_) );
  ADDFHX2 S2_2_4 ( .A(ab_2__4_), .B(n9), .CI(SUMB_1__5_), .CO(CARRYB_2__4_), 
        .S(SUMB_2__4_) );
  ADDFHX1 S2_12_2 ( .A(ab_12__2_), .B(CARRYB_11__2_), .CI(SUMB_11__3_), .CO(
        CARRYB_12__2_), .S(SUMB_12__2_) );
  ADDFHX2 S3_10_6 ( .A(ab_10__6_), .B(CARRYB_9__6_), .CI(ab_9__7_), .CO(
        CARRYB_10__6_), .S(SUMB_10__6_) );
  ADDFHX2 S4_2 ( .A(ab_16__2_), .B(CARRYB_15__2_), .CI(SUMB_15__3_), .CO(
        CARRYB_16__2_), .S(SUMB_16__2_) );
  ADDFHX2 S2_14_4 ( .A(ab_14__4_), .B(CARRYB_13__4_), .CI(SUMB_13__5_), .CO(
        CARRYB_14__4_), .S(SUMB_14__4_) );
  ADDFHX2 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  ADDFHX2 S3_7_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(
        CARRYB_7__6_), .S(SUMB_7__6_) );
  ADDFHX2 S2_10_5 ( .A(ab_10__5_), .B(CARRYB_9__5_), .CI(SUMB_9__6_), .CO(
        CARRYB_10__5_), .S(SUMB_10__5_) );
  ADDFHX2 S2_11_2 ( .A(ab_11__2_), .B(CARRYB_10__2_), .CI(SUMB_10__3_), .CO(
        CARRYB_11__2_), .S(SUMB_11__2_) );
  ADDFHX2 S3_13_6 ( .A(ab_13__6_), .B(CARRYB_12__6_), .CI(ab_12__7_), .CO(
        CARRYB_13__6_), .S(SUMB_13__6_) );
  ADDFHX2 S3_9_6 ( .A(ab_9__6_), .B(CARRYB_8__6_), .CI(ab_8__7_), .CO(
        CARRYB_9__6_), .S(SUMB_9__6_) );
  ADDFHX2 S2_9_4 ( .A(ab_9__4_), .B(CARRYB_8__4_), .CI(SUMB_8__5_), .CO(
        CARRYB_9__4_), .S(SUMB_9__4_) );
  ADDFHX2 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  ADDFHX2 S2_8_5 ( .A(ab_8__5_), .B(CARRYB_7__5_), .CI(SUMB_7__6_), .CO(
        CARRYB_8__5_), .S(SUMB_8__5_) );
  ADDFHX4 S2_13_4 ( .A(ab_13__4_), .B(CARRYB_12__4_), .CI(SUMB_12__5_), .CO(
        CARRYB_13__4_), .S(SUMB_13__4_) );
  ADDFHX4 S1_7_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(PROD1_7_) );
  ADDFHX4 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  ADDFHX4 S2_12_1 ( .A(ab_12__1_), .B(CARRYB_11__1_), .CI(SUMB_11__2_), .CO(
        CARRYB_12__1_), .S(SUMB_12__1_) );
  ADDFHX2 S2_7_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  ADDFHX4 S2_7_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  ADDFHX4 S2_8_1 ( .A(ab_8__1_), .B(CARRYB_7__1_), .CI(SUMB_7__2_), .CO(
        CARRYB_8__1_), .S(SUMB_8__1_) );
  ADDFHX4 S2_8_2 ( .A(ab_8__2_), .B(CARRYB_7__2_), .CI(SUMB_7__3_), .CO(
        CARRYB_8__2_), .S(SUMB_8__2_) );
  ADDFHX4 S2_9_2 ( .A(ab_9__2_), .B(CARRYB_8__2_), .CI(SUMB_8__3_), .CO(
        CARRYB_9__2_), .S(SUMB_9__2_) );
  ADDFHX4 S2_15_2 ( .A(ab_15__2_), .B(CARRYB_14__2_), .CI(SUMB_14__3_), .CO(
        CARRYB_15__2_), .S(SUMB_15__2_) );
  ADDFHX4 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  ADDFHX4 S1_14_0 ( .A(ab_14__0_), .B(CARRYB_13__0_), .CI(SUMB_13__1_), .CO(
        CARRYB_14__0_), .S(A1_12_) );
  ADDFHX4 S1_15_0 ( .A(ab_15__0_), .B(CARRYB_14__0_), .CI(SUMB_14__1_), .CO(
        CARRYB_15__0_), .S(A1_13_) );
  AND2X2 U2 ( .A(A[2]), .B(B[6]), .Y(ab_2__6_) );
  NAND3X2 U3 ( .A(n19), .B(n20), .C(n21), .Y(CARRYB_9__0_) );
  AND2X1 U4 ( .A(A[2]), .B(B[2]), .Y(ab_2__2_) );
  NAND2X2 U5 ( .A(ab_6__1_), .B(CARRYB_5__1_), .Y(n35) );
  AND2X2 U6 ( .A(A[1]), .B(B[6]), .Y(ab_1__6_) );
  XOR2X1 U7 ( .A(ab_14__6_), .B(ab_13__7_), .Y(n3) );
  XOR2X1 U8 ( .A(CARRYB_13__6_), .B(n3), .Y(SUMB_14__6_) );
  NAND2X1 U9 ( .A(ab_14__6_), .B(CARRYB_13__6_), .Y(n4) );
  NAND2X1 U10 ( .A(ab_13__7_), .B(CARRYB_13__6_), .Y(n5) );
  NAND2X1 U11 ( .A(ab_13__7_), .B(ab_14__6_), .Y(n6) );
  NAND3X1 U12 ( .A(n6), .B(n4), .C(n5), .Y(CARRYB_14__6_) );
  XOR2X2 U13 ( .A(CARRYB_16__1_), .B(SUMB_16__2_), .Y(A1_16_) );
  NAND3X4 U14 ( .A(n48), .B(n46), .C(n47), .Y(CARRYB_4__6_) );
  INVX3 U15 ( .A(n67), .Y(n41) );
  INVX4 U16 ( .A(B[4]), .Y(n69) );
  XOR3X2 U17 ( .A(CARRYB_5__1_), .B(ab_6__1_), .C(n26), .Y(SUMB_6__1_) );
  NAND3X4 U18 ( .A(n13), .B(n14), .C(n15), .Y(CARRYB_12__4_) );
  NAND2XL U19 ( .A(A[1]), .B(B[1]), .Y(n66) );
  XOR2X2 U20 ( .A(ab_1__3_), .B(ab_0__4_), .Y(SUMB_1__3_) );
  NOR2X2 U21 ( .A(n69), .B(n64), .Y(ab_0__4_) );
  XOR2X1 U22 ( .A(ab_1__2_), .B(ab_0__3_), .Y(SUMB_1__2_) );
  CLKINVX3 U23 ( .A(B[2]), .Y(n71) );
  NAND2XL U24 ( .A(ab_3__7_), .B(ab_4__6_), .Y(n48) );
  XOR3X2 U25 ( .A(CARRYB_6__4_), .B(ab_7__4_), .C(SUMB_6__5_), .Y(SUMB_7__4_)
         );
  INVX2 U26 ( .A(A[0]), .Y(n64) );
  XOR2X1 U27 ( .A(n30), .B(CARRYB_9__3_), .Y(SUMB_10__3_) );
  XOR2X1 U28 ( .A(ab_10__3_), .B(SUMB_9__4_), .Y(n30) );
  XOR2X1 U29 ( .A(CARRYB_16__0_), .B(SUMB_16__1_), .Y(A1_15_) );
  NOR2X2 U30 ( .A(n70), .B(n64), .Y(ab_0__3_) );
  NAND2X1 U31 ( .A(CARRYB_11__4_), .B(SUMB_11__5_), .Y(n15) );
  NAND2X1 U32 ( .A(ab_12__4_), .B(SUMB_11__5_), .Y(n14) );
  XOR3X2 U33 ( .A(SUMB_4__5_), .B(ab_5__4_), .C(CARRYB_4__4_), .Y(SUMB_5__4_)
         );
  AND2X2 U34 ( .A(CARRYB_16__1_), .B(SUMB_16__2_), .Y(n55) );
  XOR2X1 U35 ( .A(CARRYB_16__3_), .B(SUMB_16__4_), .Y(A1_18_) );
  AND2X2 U37 ( .A(ab_0__2_), .B(n74), .Y(n8) );
  AND2X2 U38 ( .A(ab_0__5_), .B(ab_1__4_), .Y(n9) );
  AND2X2 U39 ( .A(ab_0__3_), .B(ab_1__2_), .Y(n10) );
  AND2X2 U40 ( .A(ab_0__4_), .B(ab_1__3_), .Y(n11) );
  NAND2X1 U41 ( .A(ab_10__3_), .B(CARRYB_9__3_), .Y(n32) );
  XOR3X4 U42 ( .A(ab_12__4_), .B(CARRYB_11__4_), .C(SUMB_11__5_), .Y(
        SUMB_12__4_) );
  XOR2X4 U43 ( .A(ab_13__3_), .B(CARRYB_12__3_), .Y(n12) );
  XOR2X2 U44 ( .A(n12), .B(SUMB_12__4_), .Y(SUMB_13__3_) );
  NAND2X1 U45 ( .A(ab_12__4_), .B(CARRYB_11__4_), .Y(n13) );
  NAND2X1 U46 ( .A(ab_13__3_), .B(CARRYB_12__3_), .Y(n16) );
  NAND2X1 U47 ( .A(ab_13__3_), .B(SUMB_12__4_), .Y(n17) );
  NAND2X1 U48 ( .A(CARRYB_12__3_), .B(SUMB_12__4_), .Y(n18) );
  NAND3X2 U49 ( .A(n16), .B(n17), .C(n18), .Y(CARRYB_13__3_) );
  XOR3X2 U50 ( .A(ab_9__0_), .B(CARRYB_8__0_), .C(SUMB_8__1_), .Y(A1_7_) );
  NAND2X1 U51 ( .A(ab_9__0_), .B(CARRYB_8__0_), .Y(n19) );
  NAND2X1 U52 ( .A(ab_9__0_), .B(SUMB_8__1_), .Y(n20) );
  NAND2X1 U53 ( .A(CARRYB_8__0_), .B(SUMB_8__1_), .Y(n21) );
  XOR2X1 U54 ( .A(ab_10__0_), .B(SUMB_9__1_), .Y(n22) );
  XOR2X1 U55 ( .A(n22), .B(CARRYB_9__0_), .Y(A1_8_) );
  NAND2X1 U56 ( .A(ab_10__0_), .B(SUMB_9__1_), .Y(n23) );
  NAND2X1 U57 ( .A(ab_10__0_), .B(CARRYB_9__0_), .Y(n24) );
  NAND2X1 U58 ( .A(SUMB_9__1_), .B(CARRYB_9__0_), .Y(n25) );
  NAND3X2 U59 ( .A(n23), .B(n24), .C(n25), .Y(CARRYB_10__0_) );
  AND2X2 U60 ( .A(B[5]), .B(A[0]), .Y(ab_0__5_) );
  BUFX3 U61 ( .A(SUMB_5__2_), .Y(n26) );
  AND2X2 U62 ( .A(A[4]), .B(n41), .Y(ab_4__6_) );
  NAND3X2 U63 ( .A(n54), .B(n52), .C(n53), .Y(CARRYB_7__3_) );
  XOR3X2 U64 ( .A(ab_9__3_), .B(SUMB_8__4_), .C(CARRYB_8__3_), .Y(SUMB_9__3_)
         );
  NAND2X2 U65 ( .A(ab_9__3_), .B(SUMB_8__4_), .Y(n27) );
  NAND2X2 U66 ( .A(ab_9__3_), .B(CARRYB_8__3_), .Y(n28) );
  NAND2X4 U67 ( .A(SUMB_8__4_), .B(CARRYB_8__3_), .Y(n29) );
  NAND3X4 U68 ( .A(n27), .B(n28), .C(n29), .Y(CARRYB_9__3_) );
  NAND2X1 U69 ( .A(ab_10__3_), .B(SUMB_9__4_), .Y(n31) );
  NAND2X1 U70 ( .A(SUMB_9__4_), .B(CARRYB_9__3_), .Y(n33) );
  NAND3X2 U71 ( .A(n31), .B(n32), .C(n33), .Y(CARRYB_10__3_) );
  NAND2X2 U72 ( .A(SUMB_5__2_), .B(CARRYB_5__1_), .Y(n34) );
  NAND2X2 U73 ( .A(ab_6__1_), .B(SUMB_5__2_), .Y(n36) );
  NAND3X4 U74 ( .A(n36), .B(n34), .C(n35), .Y(CARRYB_6__1_) );
  INVX4 U75 ( .A(B[3]), .Y(n70) );
  XOR2X4 U76 ( .A(SUMB_6__4_), .B(ab_7__3_), .Y(n37) );
  XOR2X2 U77 ( .A(CARRYB_6__3_), .B(n37), .Y(SUMB_7__3_) );
  NAND2X2 U78 ( .A(SUMB_6__5_), .B(CARRYB_6__4_), .Y(n38) );
  NAND2X1 U79 ( .A(ab_7__4_), .B(CARRYB_6__4_), .Y(n39) );
  NAND2X2 U80 ( .A(ab_7__4_), .B(SUMB_6__5_), .Y(n40) );
  NAND3X4 U81 ( .A(n40), .B(n38), .C(n39), .Y(CARRYB_7__4_) );
  AND2X2 U82 ( .A(A[1]), .B(B[5]), .Y(ab_1__5_) );
  INVX4 U83 ( .A(B[6]), .Y(n67) );
  XOR2X2 U84 ( .A(ab_1__6_), .B(ab_0__7_), .Y(SUMB_1__6_) );
  XOR2X4 U85 ( .A(CARRYB_16__2_), .B(SUMB_16__3_), .Y(A1_17_) );
  NOR2X4 U86 ( .A(n73), .B(n64), .Y(ab_0__7_) );
  XOR3X4 U87 ( .A(CARRYB_2__5_), .B(ab_3__5_), .C(SUMB_2__6_), .Y(SUMB_3__5_)
         );
  XOR2X2 U88 ( .A(ab_1__5_), .B(ab_0__6_), .Y(SUMB_1__5_) );
  INVX4 U89 ( .A(n62), .Y(CARRYB_1__5_) );
  INVX4 U90 ( .A(n61), .Y(CARRYB_1__6_) );
  NAND2X2 U91 ( .A(ab_0__6_), .B(ab_1__5_), .Y(n62) );
  NAND2X1 U92 ( .A(ab_3__7_), .B(CARRYB_3__6_), .Y(n47) );
  NAND2X2 U93 ( .A(ab_1__6_), .B(ab_0__7_), .Y(n61) );
  NOR2X2 U94 ( .A(n71), .B(n64), .Y(ab_0__2_) );
  INVX2 U95 ( .A(n63), .Y(n73) );
  AND2X2 U96 ( .A(A[3]), .B(B[2]), .Y(ab_3__2_) );
  AND2X1 U97 ( .A(A[6]), .B(B[2]), .Y(ab_6__2_) );
  AND2X1 U98 ( .A(A[9]), .B(B[2]), .Y(ab_9__2_) );
  NAND2X2 U99 ( .A(SUMB_2__6_), .B(CARRYB_2__5_), .Y(n42) );
  NAND2X2 U100 ( .A(ab_3__5_), .B(CARRYB_2__5_), .Y(n43) );
  NAND2X2 U101 ( .A(SUMB_2__6_), .B(ab_3__5_), .Y(n44) );
  NAND3X4 U102 ( .A(n44), .B(n42), .C(n43), .Y(CARRYB_3__5_) );
  AND2X2 U103 ( .A(A[3]), .B(B[5]), .Y(ab_3__5_) );
  XOR2X1 U104 ( .A(ab_4__6_), .B(ab_3__7_), .Y(n45) );
  XOR2X1 U105 ( .A(CARRYB_3__6_), .B(n45), .Y(SUMB_4__6_) );
  NAND2X1 U106 ( .A(ab_4__6_), .B(CARRYB_3__6_), .Y(n46) );
  NAND2X2 U107 ( .A(CARRYB_4__4_), .B(SUMB_4__5_), .Y(n49) );
  NAND2X2 U108 ( .A(CARRYB_4__4_), .B(ab_5__4_), .Y(n50) );
  NAND2X2 U109 ( .A(ab_5__4_), .B(SUMB_4__5_), .Y(n51) );
  NAND3X4 U110 ( .A(n51), .B(n50), .C(n49), .Y(CARRYB_5__4_) );
  NAND2X1 U111 ( .A(SUMB_6__4_), .B(CARRYB_6__3_), .Y(n52) );
  NAND2X1 U112 ( .A(ab_7__3_), .B(CARRYB_6__3_), .Y(n53) );
  NAND2X1 U113 ( .A(ab_7__3_), .B(SUMB_6__4_), .Y(n54) );
  AND2X1 U114 ( .A(A[7]), .B(B[3]), .Y(ab_7__3_) );
  AND2X2 U115 ( .A(A[1]), .B(B[2]), .Y(ab_1__2_) );
  NOR2X4 U116 ( .A(n67), .B(n64), .Y(ab_0__6_) );
  AND2X2 U117 ( .A(CARRYB_16__0_), .B(SUMB_16__1_), .Y(n57) );
  AND2X1 U118 ( .A(CARRYB_16__2_), .B(SUMB_16__3_), .Y(n58) );
  BUFX3 U119 ( .A(B[7]), .Y(n63) );
  XOR2X1 U120 ( .A(CARRYB_16__4_), .B(SUMB_16__5_), .Y(A1_19_) );
  NOR2XL U121 ( .A(n79), .B(n68), .Y(ab_12__5_) );
  AND2X1 U122 ( .A(A[11]), .B(n63), .Y(ab_11__7_) );
  NOR2XL U123 ( .A(n79), .B(n71), .Y(ab_12__2_) );
  NOR2XL U124 ( .A(n79), .B(n72), .Y(ab_12__1_) );
  AND2X1 U125 ( .A(A[10]), .B(B[0]), .Y(ab_10__0_) );
  AND2X1 U126 ( .A(A[7]), .B(B[2]), .Y(ab_7__2_) );
  AND2X1 U127 ( .A(A[7]), .B(B[0]), .Y(ab_7__0_) );
  AND2X1 U128 ( .A(A[6]), .B(B[0]), .Y(ab_6__0_) );
  AND2X1 U129 ( .A(A[7]), .B(B[1]), .Y(ab_7__1_) );
  AND2X1 U130 ( .A(A[8]), .B(B[0]), .Y(ab_8__0_) );
  AND2X1 U131 ( .A(A[6]), .B(B[1]), .Y(ab_6__1_) );
  AND2X1 U132 ( .A(A[8]), .B(B[1]), .Y(ab_8__1_) );
  AND2X1 U133 ( .A(A[5]), .B(B[2]), .Y(ab_5__2_) );
  AND2X1 U134 ( .A(A[5]), .B(B[1]), .Y(ab_5__1_) );
  AND2X1 U135 ( .A(A[2]), .B(B[1]), .Y(ab_2__1_) );
  AND2X1 U136 ( .A(A[11]), .B(B[0]), .Y(ab_11__0_) );
  AND2X1 U137 ( .A(A[8]), .B(B[2]), .Y(ab_8__2_) );
  AND2X1 U138 ( .A(A[10]), .B(B[2]), .Y(ab_10__2_) );
  AND2X1 U139 ( .A(A[11]), .B(B[1]), .Y(ab_11__1_) );
  AND2X1 U140 ( .A(A[11]), .B(B[2]), .Y(ab_11__2_) );
  AND2X1 U141 ( .A(A[4]), .B(B[2]), .Y(ab_4__2_) );
  AND2X1 U142 ( .A(A[2]), .B(B[0]), .Y(ab_2__0_) );
  AND2X1 U143 ( .A(A[10]), .B(B[1]), .Y(ab_10__1_) );
  AND2X1 U144 ( .A(A[9]), .B(B[1]), .Y(ab_9__1_) );
  INVXL U145 ( .A(B[0]), .Y(n80) );
  INVXL U146 ( .A(B[1]), .Y(n72) );
  NOR2X1 U147 ( .A(n75), .B(n68), .Y(ab_16__5_) );
  AND2X2 U148 ( .A(CARRYB_16__3_), .B(SUMB_16__4_), .Y(n56) );
  XOR2X1 U149 ( .A(n74), .B(ab_0__2_), .Y(SUMB_1__1_) );
  XOR2X1 U150 ( .A(CARRYB_16__5_), .B(SUMB_16__6_), .Y(A1_20_) );
  XOR2X1 U151 ( .A(CARRYB_16__6_), .B(ab_16__7_), .Y(A1_21_) );
  AND2X1 U152 ( .A(CARRYB_16__4_), .B(SUMB_16__5_), .Y(n59) );
  AND2X2 U153 ( .A(CARRYB_16__5_), .B(SUMB_16__6_), .Y(n60) );
  NOR2X1 U154 ( .A(n75), .B(n73), .Y(ab_16__7_) );
  NOR2X1 U155 ( .A(n75), .B(n72), .Y(ab_16__1_) );
  NOR2X1 U156 ( .A(n75), .B(n71), .Y(ab_16__2_) );
  NOR2XL U157 ( .A(n75), .B(n69), .Y(ab_16__4_) );
  NOR2X1 U158 ( .A(n76), .B(n73), .Y(ab_15__7_) );
  AND2X2 U159 ( .A(A[1]), .B(B[3]), .Y(ab_1__3_) );
  INVX1 U160 ( .A(n66), .Y(n74) );
  NOR2X1 U161 ( .A(n77), .B(n72), .Y(ab_14__1_) );
  NOR2X1 U162 ( .A(n76), .B(n72), .Y(ab_15__1_) );
  NOR2X1 U163 ( .A(n78), .B(n72), .Y(ab_13__1_) );
  NOR2X1 U164 ( .A(n78), .B(n71), .Y(ab_13__2_) );
  NOR2X1 U165 ( .A(n77), .B(n71), .Y(ab_14__2_) );
  AND2X2 U166 ( .A(A[11]), .B(B[3]), .Y(ab_11__3_) );
  AND2X2 U167 ( .A(A[10]), .B(B[3]), .Y(ab_10__3_) );
  AND2X2 U168 ( .A(A[9]), .B(B[3]), .Y(ab_9__3_) );
  AND2X2 U169 ( .A(A[8]), .B(B[3]), .Y(ab_8__3_) );
  NOR2XL U170 ( .A(n78), .B(n69), .Y(ab_13__4_) );
  NOR2XL U171 ( .A(n77), .B(n69), .Y(ab_14__4_) );
  NOR2XL U172 ( .A(n79), .B(n69), .Y(ab_12__4_) );
  NOR2X1 U173 ( .A(n77), .B(n68), .Y(ab_14__5_) );
  AND2X1 U174 ( .A(A[11]), .B(B[5]), .Y(ab_11__5_) );
  NOR2X1 U175 ( .A(n78), .B(n68), .Y(ab_13__5_) );
  AND2X1 U176 ( .A(A[10]), .B(B[5]), .Y(ab_10__5_) );
  AND2X1 U177 ( .A(A[9]), .B(B[5]), .Y(ab_9__5_) );
  AND2X1 U178 ( .A(A[8]), .B(B[5]), .Y(ab_8__5_) );
  NOR2XL U179 ( .A(n79), .B(n73), .Y(ab_12__7_) );
  AND2X2 U180 ( .A(A[6]), .B(B[3]), .Y(ab_6__3_) );
  AND2X1 U181 ( .A(A[7]), .B(B[5]), .Y(ab_7__5_) );
  AND2X1 U182 ( .A(A[6]), .B(B[5]), .Y(ab_6__5_) );
  AND2X1 U183 ( .A(A[4]), .B(B[3]), .Y(ab_4__3_) );
  AND2X1 U184 ( .A(A[4]), .B(B[5]), .Y(ab_4__5_) );
  AND2X1 U185 ( .A(A[5]), .B(B[5]), .Y(ab_5__5_) );
  AND2X2 U186 ( .A(A[5]), .B(B[3]), .Y(ab_5__3_) );
  AND2X2 U187 ( .A(A[3]), .B(B[3]), .Y(ab_3__3_) );
  AND2X2 U188 ( .A(A[2]), .B(B[3]), .Y(ab_2__3_) );
  XOR2X1 U189 ( .A(ab_1__4_), .B(ab_0__5_), .Y(SUMB_1__4_) );
  NOR2XL U190 ( .A(n78), .B(n73), .Y(ab_13__7_) );
  AND2X1 U191 ( .A(A[2]), .B(B[5]), .Y(ab_2__5_) );
  NOR2XL U192 ( .A(n77), .B(n73), .Y(ab_14__7_) );
  NOR2X1 U193 ( .A(n76), .B(n71), .Y(ab_15__2_) );
  NOR2XL U194 ( .A(n76), .B(n69), .Y(ab_15__4_) );
  NOR2X1 U195 ( .A(n76), .B(n68), .Y(ab_15__5_) );
  INVX1 U196 ( .A(A[16]), .Y(n75) );
  INVXL U197 ( .A(B[5]), .Y(n68) );
  AND2X1 U198 ( .A(A[2]), .B(B[4]), .Y(ab_2__4_) );
  AND2X2 U199 ( .A(A[1]), .B(B[4]), .Y(ab_1__4_) );
  NAND2XL U200 ( .A(A[0]), .B(B[0]), .Y(n65) );
  AND2X1 U201 ( .A(A[3]), .B(B[4]), .Y(ab_3__4_) );
  AND2X1 U202 ( .A(A[11]), .B(B[4]), .Y(ab_11__4_) );
  AND2X1 U203 ( .A(A[10]), .B(B[4]), .Y(ab_10__4_) );
  AND2X1 U204 ( .A(A[9]), .B(B[4]), .Y(ab_9__4_) );
  AND2X1 U205 ( .A(A[8]), .B(B[4]), .Y(ab_8__4_) );
  AND2X1 U206 ( .A(A[7]), .B(B[4]), .Y(ab_7__4_) );
  AND2X1 U207 ( .A(A[10]), .B(n63), .Y(ab_10__7_) );
  AND2X1 U208 ( .A(A[6]), .B(B[4]), .Y(ab_6__4_) );
  AND2X2 U209 ( .A(A[9]), .B(B[0]), .Y(ab_9__0_) );
  AND2X1 U210 ( .A(A[4]), .B(B[4]), .Y(ab_4__4_) );
  AND2X1 U211 ( .A(A[5]), .B(B[4]), .Y(ab_5__4_) );
  AND2X1 U212 ( .A(A[9]), .B(n63), .Y(ab_9__7_) );
  AND2X1 U213 ( .A(A[8]), .B(n63), .Y(ab_8__7_) );
  AND2X1 U214 ( .A(A[7]), .B(n63), .Y(ab_7__7_) );
  AND2X1 U215 ( .A(A[2]), .B(n63), .Y(ab_2__7_) );
  AND2X1 U216 ( .A(A[3]), .B(B[1]), .Y(ab_3__1_) );
  AND2X1 U217 ( .A(A[4]), .B(B[1]), .Y(ab_4__1_) );
  AND2X1 U218 ( .A(A[3]), .B(n63), .Y(ab_3__7_) );
  AND2X1 U219 ( .A(A[6]), .B(n63), .Y(ab_6__7_) );
  AND2X1 U220 ( .A(A[4]), .B(n63), .Y(ab_4__7_) );
  AND2X1 U221 ( .A(A[5]), .B(n63), .Y(ab_5__7_) );
  AND2X1 U222 ( .A(A[3]), .B(B[0]), .Y(ab_3__0_) );
  NOR2XL U223 ( .A(n66), .B(n65), .Y(CARRYB_1__0_) );
  AND2X2 U224 ( .A(A[5]), .B(B[0]), .Y(ab_5__0_) );
  AND2X1 U225 ( .A(A[4]), .B(B[0]), .Y(ab_4__0_) );
  AND2X1 U226 ( .A(A[1]), .B(n63), .Y(ab_1__7_) );
  INVX1 U227 ( .A(A[14]), .Y(n77) );
  INVX1 U228 ( .A(A[15]), .Y(n76) );
  INVX1 U229 ( .A(A[12]), .Y(n79) );
  INVX1 U230 ( .A(A[13]), .Y(n78) );
  NOR2XL U231 ( .A(n75), .B(n67), .Y(ab_16__6_) );
  NOR2XL U232 ( .A(n76), .B(n67), .Y(ab_15__6_) );
  NOR2XL U233 ( .A(n77), .B(n67), .Y(ab_14__6_) );
  NOR2XL U234 ( .A(n78), .B(n67), .Y(ab_13__6_) );
  NOR2XL U235 ( .A(n79), .B(n67), .Y(ab_12__6_) );
  AND2X1 U236 ( .A(A[11]), .B(n41), .Y(ab_11__6_) );
  AND2X1 U237 ( .A(A[10]), .B(n41), .Y(ab_10__6_) );
  AND2X1 U238 ( .A(A[9]), .B(n41), .Y(ab_9__6_) );
  AND2X1 U239 ( .A(A[8]), .B(n41), .Y(ab_8__6_) );
  AND2X1 U240 ( .A(A[7]), .B(n41), .Y(ab_7__6_) );
  AND2X1 U241 ( .A(A[6]), .B(n41), .Y(ab_6__6_) );
  AND2X1 U242 ( .A(A[5]), .B(n41), .Y(ab_5__6_) );
  AND2X1 U243 ( .A(A[3]), .B(n41), .Y(ab_3__6_) );
  NOR2XL U244 ( .A(n75), .B(n70), .Y(ab_16__3_) );
  NOR2XL U245 ( .A(n76), .B(n70), .Y(ab_15__3_) );
  NOR2XL U246 ( .A(n77), .B(n70), .Y(ab_14__3_) );
  NOR2XL U247 ( .A(n78), .B(n70), .Y(ab_13__3_) );
  NOR2XL U248 ( .A(n79), .B(n70), .Y(ab_12__3_) );
  NOR2X1 U250 ( .A(n80), .B(n75), .Y(ab_16__0_) );
  NOR2X1 U251 ( .A(n80), .B(n76), .Y(ab_15__0_) );
  NOR2X1 U252 ( .A(n80), .B(n77), .Y(ab_14__0_) );
  NOR2X1 U253 ( .A(n80), .B(n78), .Y(ab_13__0_) );
  NOR2X1 U254 ( .A(n80), .B(n79), .Y(ab_12__0_) );
endmodule


module multi16_11 ( in_17bit, in_8bit, out );
  input [16:0] in_17bit;
  input [7:0] in_8bit;
  output [16:0] out;
  wire   N19, N20, N21, N32, N33, n54, n62, n70, n77, n1, n2, n3, n4, n5, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n55, n56, n57, n58, n59, n60, n61, n63, n64,
         n65, n66, n67, n68, n69, n71, n72, n73, n74, n75, n76, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120;
  wire   [16:1] in_17bit_b;
  wire   [7:0] in_8bit_b;
  wire   [23:8] mul;
  wire   [16:13] sub_add_52_b0_carry;

  multi16_11_DW02_mult_0 mult_55 ( .A({in_17bit_b, in_17bit[0]}), .B(in_8bit_b), .PRODUCT_23_(mul[23]), .PRODUCT_22_(mul[22]), .PRODUCT_21_(mul[21]), 
        .PRODUCT_20_(mul[20]), .PRODUCT_19_(mul[19]), .PRODUCT_18_(mul[18]), 
        .PRODUCT_17_(mul[17]), .PRODUCT_16_(mul[16]), .PRODUCT_15_(mul[15]), 
        .PRODUCT_14_(mul[14]), .PRODUCT_13_(mul[13]), .PRODUCT_12_(mul[12]), 
        .PRODUCT_11_(mul[11]), .PRODUCT_10_(mul[10]), .PRODUCT_9_(mul[9]), 
        .PRODUCT_8_(mul[8]), .PRODUCT_7_(N32) );
  INVX12 U2 ( .A(in_17bit[16]), .Y(n26) );
  NAND2BX2 U3 ( .AN(mul[21]), .B(n109), .Y(n110) );
  NOR3BX2 U4 ( .AN(n41), .B(n40), .C(n39), .Y(in_17bit_b[1]) );
  NAND3X1 U5 ( .A(in_17bit[0]), .B(n25), .C(in_17bit[1]), .Y(n41) );
  NOR2X1 U6 ( .A(n104), .B(mul[18]), .Y(n5) );
  INVX4 U7 ( .A(n27), .Y(n25) );
  NAND2X4 U8 ( .A(in_8bit[6]), .B(n2), .Y(n3) );
  NAND2X2 U9 ( .A(n1), .B(n22), .Y(n4) );
  NAND2X4 U10 ( .A(n3), .B(n4), .Y(in_8bit_b[6]) );
  CLKINVXL U11 ( .A(in_8bit[6]), .Y(n1) );
  CLKINVX4 U12 ( .A(n22), .Y(n2) );
  NOR2X4 U13 ( .A(n6), .B(mul[19]), .Y(n106) );
  CLKINVX3 U14 ( .A(n5), .Y(n6) );
  NOR2X2 U15 ( .A(n120), .B(n31), .Y(n16) );
  XOR2X4 U16 ( .A(n32), .B(in_8bit[4]), .Y(in_8bit_b[4]) );
  AND2X2 U17 ( .A(n45), .B(n25), .Y(n13) );
  NAND2XL U18 ( .A(n52), .B(n25), .Y(n51) );
  XOR2X4 U19 ( .A(n7), .B(n105), .Y(out[13]) );
  AOI21X2 U20 ( .A0(n31), .A1(n30), .B0(n120), .Y(n32) );
  NOR3X2 U21 ( .A(in_8bit[0]), .B(in_8bit[2]), .C(in_8bit[1]), .Y(n31) );
  XOR2X1 U22 ( .A(n108), .B(mul[21]), .Y(out[14]) );
  NOR2X2 U23 ( .A(n19), .B(n99), .Y(n98) );
  NAND2X2 U24 ( .A(n10), .B(n11), .Y(in_8bit_b[2]) );
  NAND2XL U25 ( .A(n9), .B(in_8bit[2]), .Y(n11) );
  NOR2X2 U26 ( .A(n26), .B(n21), .Y(n42) );
  NOR2XL U27 ( .A(n26), .B(n50), .Y(n48) );
  XNOR2X1 U28 ( .A(in_8bit[1]), .B(n28), .Y(in_8bit_b[1]) );
  INVX1 U29 ( .A(n77), .Y(in_8bit_b[0]) );
  INVX1 U30 ( .A(n23), .Y(n9) );
  INVX1 U31 ( .A(n89), .Y(n91) );
  NAND2BX1 U32 ( .AN(mul[12]), .B(n88), .Y(n89) );
  INVX1 U33 ( .A(n95), .Y(n96) );
  NAND2BX1 U34 ( .AN(mul[14]), .B(n94), .Y(n95) );
  NAND2BX2 U35 ( .AN(mul[15]), .B(n96), .Y(n97) );
  XOR2X1 U36 ( .A(mul[14]), .B(n93), .Y(out[7]) );
  NOR2X2 U37 ( .A(mul[16]), .B(n97), .Y(n12) );
  XNOR2X2 U38 ( .A(n35), .B(n36), .Y(in_8bit_b[5]) );
  INVX1 U39 ( .A(mul[8]), .Y(n114) );
  NOR2X2 U40 ( .A(n19), .B(n106), .Y(n105) );
  CLKINVX3 U41 ( .A(mul[22]), .Y(n112) );
  CLKINVX3 U42 ( .A(in_17bit[16]), .Y(n27) );
  INVX1 U43 ( .A(in_8bit[2]), .Y(n24) );
  CLKINVX3 U44 ( .A(n97), .Y(n99) );
  NOR2XL U45 ( .A(in_17bit[1]), .B(in_17bit[0]), .Y(n40) );
  NAND2X1 U46 ( .A(n23), .B(n24), .Y(n10) );
  INVX1 U47 ( .A(n29), .Y(n23) );
  CLKINVX4 U48 ( .A(n107), .Y(n109) );
  BUFX1 U49 ( .A(mul[20]), .Y(n7) );
  AND2X4 U50 ( .A(n110), .B(n54), .Y(n111) );
  AOI21X1 U51 ( .A0(n8), .A1(n112), .B0(n19), .Y(n113) );
  NOR2BX4 U52 ( .AN(n54), .B(n109), .Y(n108) );
  OAI21XL U53 ( .A0(in_8bit[1]), .A1(in_8bit[0]), .B0(in_8bit[7]), .Y(n29) );
  INVXL U54 ( .A(n110), .Y(n8) );
  NOR2X2 U55 ( .A(n19), .B(n12), .Y(n100) );
  XOR2X4 U56 ( .A(n102), .B(mul[18]), .Y(out[11]) );
  INVX8 U57 ( .A(n34), .Y(n37) );
  NOR3X2 U58 ( .A(in_8bit[6]), .B(n38), .C(n120), .Y(in_8bit_b[7]) );
  NAND2X4 U59 ( .A(n37), .B(n36), .Y(n38) );
  OAI21X2 U60 ( .A0(mul[18]), .A1(n104), .B0(n54), .Y(n103) );
  OR2X4 U61 ( .A(n19), .B(n96), .Y(n20) );
  NOR2X4 U62 ( .A(n101), .B(n19), .Y(n102) );
  INVX4 U63 ( .A(n104), .Y(n101) );
  NOR2X4 U64 ( .A(n120), .B(n37), .Y(n35) );
  XOR2X2 U65 ( .A(mul[17]), .B(n100), .Y(out[10]) );
  XNOR2X4 U66 ( .A(n16), .B(n30), .Y(in_8bit_b[3]) );
  NAND2BX4 U67 ( .AN(mul[17]), .B(n12), .Y(n104) );
  NAND2BX4 U68 ( .AN(in_8bit[0]), .B(n33), .Y(n34) );
  NOR2X2 U69 ( .A(in_17bit[1]), .B(in_17bit[0]), .Y(n21) );
  XOR2X2 U70 ( .A(n15), .B(in_17bit[3]), .Y(in_17bit_b[3]) );
  NOR2X2 U71 ( .A(n26), .B(n44), .Y(n15) );
  XOR2X1 U72 ( .A(mul[16]), .B(n98), .Y(out[9]) );
  NOR2X1 U73 ( .A(n26), .B(n14), .Y(n72) );
  XNOR2X2 U74 ( .A(n48), .B(n49), .Y(in_17bit_b[5]) );
  XNOR2X1 U75 ( .A(n46), .B(n13), .Y(in_17bit_b[4]) );
  NAND2XL U76 ( .A(n50), .B(n49), .Y(n52) );
  NAND2BXL U77 ( .AN(n45), .B(n46), .Y(n47) );
  NOR2XL U78 ( .A(n26), .B(n66), .Y(n64) );
  NAND2XL U79 ( .A(n60), .B(n25), .Y(n59) );
  NAND2XL U80 ( .A(n58), .B(n57), .Y(n60) );
  NAND2BXL U81 ( .AN(n52), .B(n53), .Y(n55) );
  NAND2BXL U82 ( .AN(n60), .B(n61), .Y(n63) );
  NAND2XL U83 ( .A(n68), .B(n25), .Y(n67) );
  AND2X2 U84 ( .A(n71), .B(n69), .Y(n14) );
  NAND2XL U85 ( .A(n66), .B(n65), .Y(n68) );
  NAND2XL U86 ( .A(n14), .B(n74), .Y(n73) );
  AND2X1 U87 ( .A(N21), .B(n25), .Y(in_17bit_b[16]) );
  INVX1 U88 ( .A(n43), .Y(n44) );
  XOR2X1 U89 ( .A(mul[23]), .B(n113), .Y(out[16]) );
  NOR2XL U90 ( .A(n19), .B(n91), .Y(n90) );
  NOR2XL U91 ( .A(n19), .B(n85), .Y(n84) );
  NOR2XL U92 ( .A(n19), .B(n79), .Y(n78) );
  MX2X1 U93 ( .A(in_17bit[14]), .B(N19), .S0(n25), .Y(in_17bit_b[14]) );
  MX2X1 U94 ( .A(in_17bit[12]), .B(n17), .S0(n25), .Y(in_17bit_b[12]) );
  XNOR2X1 U95 ( .A(n73), .B(n116), .Y(n17) );
  MX2X1 U96 ( .A(in_17bit[13]), .B(n18), .S0(n25), .Y(in_17bit_b[13]) );
  XNOR2X1 U97 ( .A(n75), .B(n117), .Y(n18) );
  MX2X1 U98 ( .A(in_17bit[15]), .B(N20), .S0(n25), .Y(in_17bit_b[15]) );
  AOI22XL U99 ( .A0(mul[8]), .A1(n19), .B0(N33), .B1(n54), .Y(n62) );
  AND2X4 U100 ( .A(n38), .B(in_8bit[7]), .Y(n22) );
  XNOR2X1 U101 ( .A(n25), .B(in_8bit[7]), .Y(n19) );
  INVX1 U102 ( .A(n92), .Y(n94) );
  NAND2BX1 U103 ( .AN(mul[13]), .B(n91), .Y(n92) );
  INVX1 U104 ( .A(n80), .Y(n82) );
  NAND2BX1 U105 ( .AN(mul[9]), .B(n79), .Y(n80) );
  INVX1 U106 ( .A(n83), .Y(n85) );
  NAND2BX1 U107 ( .AN(mul[10]), .B(n82), .Y(n83) );
  INVX1 U108 ( .A(n86), .Y(n88) );
  NAND2BX1 U109 ( .AN(mul[11]), .B(n85), .Y(n86) );
  INVX1 U110 ( .A(n76), .Y(n79) );
  NAND2BX1 U111 ( .AN(mul[8]), .B(n115), .Y(n76) );
  INVX1 U112 ( .A(N32), .Y(n115) );
  INVXL U113 ( .A(in_8bit[3]), .Y(n30) );
  XNOR2X1 U114 ( .A(n56), .B(n57), .Y(in_17bit_b[7]) );
  NOR2X1 U115 ( .A(n26), .B(n58), .Y(n56) );
  XNOR2X1 U116 ( .A(n64), .B(n65), .Y(in_17bit_b[9]) );
  XOR2X1 U117 ( .A(n53), .B(n51), .Y(in_17bit_b[6]) );
  XOR2X1 U118 ( .A(n61), .B(n59), .Y(in_17bit_b[8]) );
  INVX1 U119 ( .A(n47), .Y(n50) );
  INVX1 U120 ( .A(n55), .Y(n58) );
  INVX1 U121 ( .A(n63), .Y(n66) );
  NAND3X1 U122 ( .A(n116), .B(n14), .C(n74), .Y(n75) );
  XOR2X1 U123 ( .A(n69), .B(n67), .Y(in_17bit_b[10]) );
  INVX1 U124 ( .A(n75), .Y(sub_add_52_b0_carry[13]) );
  XNOR2X1 U125 ( .A(n72), .B(n74), .Y(in_17bit_b[11]) );
  INVX1 U126 ( .A(n68), .Y(n71) );
  NOR2X1 U127 ( .A(in_17bit[1]), .B(n25), .Y(n39) );
  INVXL U128 ( .A(in_8bit[5]), .Y(n36) );
  INVX1 U129 ( .A(in_17bit[5]), .Y(n49) );
  XOR2X1 U130 ( .A(mul[13]), .B(n90), .Y(out[6]) );
  XNOR2X1 U131 ( .A(mul[15]), .B(n20), .Y(out[8]) );
  NOR2X1 U132 ( .A(n19), .B(n94), .Y(n93) );
  XOR2X1 U133 ( .A(mul[12]), .B(n87), .Y(out[5]) );
  NOR2X1 U134 ( .A(n19), .B(n88), .Y(n87) );
  XOR2X1 U135 ( .A(mul[11]), .B(n84), .Y(out[4]) );
  XOR2X1 U136 ( .A(mul[9]), .B(n78), .Y(out[2]) );
  XOR2X1 U137 ( .A(mul[10]), .B(n81), .Y(out[3]) );
  NOR2X1 U138 ( .A(n19), .B(n82), .Y(n81) );
  NAND2BXL U139 ( .AN(in_17bit[3]), .B(n44), .Y(n45) );
  INVX1 U140 ( .A(in_17bit[4]), .Y(n46) );
  INVX1 U141 ( .A(n62), .Y(out[1]) );
  INVX1 U142 ( .A(in_17bit[7]), .Y(n57) );
  INVX1 U143 ( .A(in_17bit[6]), .Y(n53) );
  INVX1 U144 ( .A(in_17bit[8]), .Y(n61) );
  INVX1 U145 ( .A(n70), .Y(out[0]) );
  AOI22XL U146 ( .A0(N32), .A1(n19), .B0(N32), .B1(n54), .Y(n70) );
  INVX1 U147 ( .A(in_17bit[11]), .Y(n74) );
  INVX1 U148 ( .A(in_17bit[9]), .Y(n65) );
  INVX1 U149 ( .A(in_17bit[10]), .Y(n69) );
  INVX1 U150 ( .A(in_17bit[12]), .Y(n116) );
  INVXL U151 ( .A(n19), .Y(n54) );
  INVX1 U152 ( .A(in_17bit[13]), .Y(n117) );
  INVX1 U153 ( .A(in_17bit[14]), .Y(n118) );
  INVX1 U154 ( .A(in_17bit[15]), .Y(n119) );
  INVX1 U155 ( .A(in_8bit[7]), .Y(n120) );
  NAND2BX1 U156 ( .AN(in_17bit[2]), .B(n21), .Y(n43) );
  XOR2X2 U157 ( .A(in_17bit[2]), .B(n42), .Y(in_17bit_b[2]) );
  XNOR2X2 U158 ( .A(mul[19]), .B(n103), .Y(out[12]) );
  NOR4X2 U159 ( .A(in_8bit[1]), .B(in_8bit[2]), .C(in_8bit[4]), .D(in_8bit[3]), 
        .Y(n33) );
  NAND2BX2 U160 ( .AN(mul[20]), .B(n106), .Y(n107) );
  AOI22XL U161 ( .A0(in_8bit[0]), .A1(in_8bit[7]), .B0(in_8bit[0]), .B1(n120), 
        .Y(n77) );
  NAND2XL U162 ( .A(in_8bit[0]), .B(in_8bit[7]), .Y(n28) );
  XNOR2X4 U163 ( .A(n111), .B(n112), .Y(out[15]) );
  XOR2X1 U164 ( .A(n114), .B(n115), .Y(N33) );
  XOR2X1 U165 ( .A(n26), .B(sub_add_52_b0_carry[16]), .Y(N21) );
  AND2X1 U166 ( .A(sub_add_52_b0_carry[15]), .B(n119), .Y(
        sub_add_52_b0_carry[16]) );
  XOR2X1 U167 ( .A(n119), .B(sub_add_52_b0_carry[15]), .Y(N20) );
  AND2X1 U168 ( .A(sub_add_52_b0_carry[14]), .B(n118), .Y(
        sub_add_52_b0_carry[15]) );
  XOR2X1 U169 ( .A(n118), .B(sub_add_52_b0_carry[14]), .Y(N19) );
  AND2X1 U170 ( .A(sub_add_52_b0_carry[13]), .B(n117), .Y(
        sub_add_52_b0_carry[14]) );
endmodule


module multi16_10_DW01_add_0 ( A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, 
        A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, 
        B_20_, B_19_, B_18_, B_17_, B_16_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, 
        SUM_17_, SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, 
        SUM_9_, SUM_8_, SUM_7_, SUM_6_, SUM_5_ );
  input A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_,
         A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, B_20_, B_19_,
         B_18_, B_17_, B_16_;
  output SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, SUM_15_,
         SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, SUM_7_,
         SUM_6_, SUM_5_;
  wire   n1, n2, n3, n4, n6, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43;

  CLKINVX4 U2 ( .A(n1), .Y(n2) );
  INVX2 U3 ( .A(n43), .Y(n1) );
  BUFX3 U4 ( .A(A_13_), .Y(SUM_13_) );
  NAND2X4 U5 ( .A(B_16_), .B(A_16_), .Y(n37) );
  OAI21X1 U6 ( .A0(n33), .A1(n37), .B0(n4), .Y(n35) );
  INVX1 U7 ( .A(n33), .Y(n21) );
  CLKINVX4 U8 ( .A(n37), .Y(n22) );
  OAI21XL U9 ( .A0(n30), .A1(n31), .B0(n32), .Y(n26) );
  INVX1 U10 ( .A(n20), .Y(n4) );
  NOR2X1 U11 ( .A(B_16_), .B(A_16_), .Y(n6) );
  NAND2X2 U12 ( .A(n22), .B(n21), .Y(n3) );
  INVX2 U13 ( .A(n38), .Y(n20) );
  NOR2X2 U14 ( .A(B_17_), .B(A_17_), .Y(n33) );
  NAND2X2 U15 ( .A(B_17_), .B(A_17_), .Y(n38) );
  NAND2X2 U16 ( .A(B_18_), .B(A_18_), .Y(n36) );
  NOR2X1 U17 ( .A(n33), .B(n20), .Y(n43) );
  NOR2X4 U18 ( .A(B_18_), .B(A_18_), .Y(n34) );
  OAI21X4 U19 ( .A0(n41), .A1(n34), .B0(n36), .Y(n39) );
  INVX2 U20 ( .A(n34), .Y(n18) );
  NOR2BX2 U21 ( .AN(n32), .B(n31), .Y(n40) );
  NOR2X1 U22 ( .A(B_19_), .B(A_19_), .Y(n31) );
  CLKINVX4 U23 ( .A(n23), .Y(SUM_15_) );
  XOR2X4 U24 ( .A(n42), .B(n41), .Y(SUM_18_) );
  XOR2X4 U25 ( .A(n39), .B(n40), .Y(SUM_19_) );
  NOR2BX2 U26 ( .AN(n37), .B(n6), .Y(SUM_16_) );
  AND2X4 U27 ( .A(n3), .B(n4), .Y(n41) );
  INVXL U28 ( .A(n28), .Y(n17) );
  BUFX4 U29 ( .A(A_14_), .Y(SUM_14_) );
  AOI21XL U30 ( .A0(n26), .A1(n27), .B0(n17), .Y(n25) );
  BUFX3 U31 ( .A(A_12_), .Y(SUM_12_) );
  INVX1 U32 ( .A(n36), .Y(n19) );
  NAND2X1 U33 ( .A(n36), .B(n18), .Y(n42) );
  BUFX3 U34 ( .A(A_5_), .Y(SUM_5_) );
  BUFX3 U35 ( .A(A_6_), .Y(SUM_6_) );
  BUFX3 U36 ( .A(A_7_), .Y(SUM_7_) );
  BUFX3 U37 ( .A(A_8_), .Y(SUM_8_) );
  BUFX3 U38 ( .A(A_10_), .Y(SUM_10_) );
  BUFX3 U39 ( .A(A_11_), .Y(SUM_11_) );
  BUFX3 U40 ( .A(A_9_), .Y(SUM_9_) );
  INVX4 U41 ( .A(A_15_), .Y(n23) );
  XOR2X4 U42 ( .A(n22), .B(n2), .Y(SUM_17_) );
  XOR2X1 U43 ( .A(n24), .B(n25), .Y(SUM_21_) );
  XNOR2X1 U44 ( .A(B_21_), .B(A_21_), .Y(n24) );
  XNOR2X1 U45 ( .A(n29), .B(n26), .Y(SUM_20_) );
  AOI21X1 U46 ( .A0(n18), .A1(n35), .B0(n19), .Y(n30) );
  NAND2X1 U47 ( .A(n28), .B(n27), .Y(n29) );
  OR2X1 U48 ( .A(B_20_), .B(A_20_), .Y(n27) );
  NAND2X1 U49 ( .A(B_20_), .B(A_20_), .Y(n28) );
  NAND2X1 U50 ( .A(B_19_), .B(A_19_), .Y(n32) );
endmodule


module multi16_10_DW02_mult_0 ( A, B, PRODUCT_23_, PRODUCT_22_, PRODUCT_21_, 
        PRODUCT_20_, PRODUCT_19_, PRODUCT_18_, PRODUCT_17_, PRODUCT_16_, 
        PRODUCT_15_, PRODUCT_14_, PRODUCT_13_, PRODUCT_12_, PRODUCT_11_, 
        PRODUCT_10_, PRODUCT_9_, PRODUCT_8_, PRODUCT_7_ );
  input [16:0] A;
  input [7:0] B;
  output PRODUCT_23_, PRODUCT_22_, PRODUCT_21_, PRODUCT_20_, PRODUCT_19_,
         PRODUCT_18_, PRODUCT_17_, PRODUCT_16_, PRODUCT_15_, PRODUCT_14_,
         PRODUCT_13_, PRODUCT_12_, PRODUCT_11_, PRODUCT_10_, PRODUCT_9_,
         PRODUCT_8_, PRODUCT_7_;
  wire   ab_16__7_, ab_16__6_, ab_16__5_, ab_16__4_, ab_16__3_, ab_16__2_,
         ab_16__1_, ab_16__0_, ab_15__7_, ab_15__6_, ab_15__5_, ab_15__4_,
         ab_15__3_, ab_15__2_, ab_15__1_, ab_15__0_, ab_14__7_, ab_14__6_,
         ab_14__5_, ab_14__4_, ab_14__3_, ab_14__2_, ab_14__1_, ab_14__0_,
         ab_13__7_, ab_13__6_, ab_13__5_, ab_13__4_, ab_13__3_, ab_13__2_,
         ab_13__1_, ab_13__0_, ab_12__7_, ab_12__6_, ab_12__5_, ab_12__4_,
         ab_12__3_, ab_12__2_, ab_12__1_, ab_12__0_, ab_11__7_, ab_11__6_,
         ab_11__5_, ab_11__4_, ab_11__3_, ab_11__2_, ab_11__1_, ab_11__0_,
         ab_10__7_, ab_10__6_, ab_10__5_, ab_10__4_, ab_10__3_, ab_10__2_,
         ab_10__1_, ab_10__0_, ab_9__7_, ab_9__6_, ab_9__5_, ab_9__4_,
         ab_9__3_, ab_9__2_, ab_9__1_, ab_9__0_, ab_8__7_, ab_8__6_, ab_8__5_,
         ab_8__4_, ab_8__3_, ab_8__2_, ab_8__1_, ab_8__0_, ab_7__7_, ab_7__6_,
         ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_, ab_7__0_, ab_6__7_,
         ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_, ab_6__1_, ab_6__0_,
         ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_, ab_5__2_, ab_5__1_,
         ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_, ab_4__3_, ab_4__2_,
         ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_, ab_3__4_, ab_3__3_,
         ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_, ab_2__5_, ab_2__4_,
         ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_, ab_1__6_, ab_1__5_,
         ab_1__4_, ab_1__3_, ab_1__2_, ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_,
         ab_0__3_, ab_0__2_, CARRYB_16__6_, CARRYB_16__5_, CARRYB_16__4_,
         CARRYB_16__3_, CARRYB_16__2_, CARRYB_16__1_, CARRYB_16__0_,
         CARRYB_15__6_, CARRYB_15__5_, CARRYB_15__4_, CARRYB_15__3_,
         CARRYB_15__2_, CARRYB_15__1_, CARRYB_15__0_, CARRYB_14__6_,
         CARRYB_14__5_, CARRYB_14__4_, CARRYB_14__3_, CARRYB_14__2_,
         CARRYB_14__1_, CARRYB_14__0_, CARRYB_13__6_, CARRYB_13__5_,
         CARRYB_13__4_, CARRYB_13__3_, CARRYB_13__2_, CARRYB_13__1_,
         CARRYB_13__0_, CARRYB_12__6_, CARRYB_12__5_, CARRYB_12__4_,
         CARRYB_12__3_, CARRYB_12__2_, CARRYB_12__1_, CARRYB_12__0_,
         CARRYB_11__6_, CARRYB_11__5_, CARRYB_11__4_, CARRYB_11__3_,
         CARRYB_11__2_, CARRYB_11__1_, CARRYB_11__0_, CARRYB_10__6_,
         CARRYB_10__5_, CARRYB_10__4_, CARRYB_10__3_, CARRYB_10__2_,
         CARRYB_10__1_, CARRYB_10__0_, CARRYB_9__6_, CARRYB_9__5_,
         CARRYB_9__4_, CARRYB_9__3_, CARRYB_9__2_, CARRYB_9__1_, CARRYB_9__0_,
         CARRYB_8__6_, CARRYB_8__5_, CARRYB_8__4_, CARRYB_8__3_, CARRYB_8__2_,
         CARRYB_8__1_, CARRYB_8__0_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_,
         CARRYB_7__3_, CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_,
         CARRYB_6__5_, CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_,
         CARRYB_6__0_, CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_,
         CARRYB_5__2_, CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_,
         CARRYB_4__4_, CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_,
         CARRYB_3__6_, CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_,
         CARRYB_3__1_, CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_,
         CARRYB_2__3_, CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__0_,
         SUMB_16__6_, SUMB_16__5_, SUMB_16__4_, SUMB_16__3_, SUMB_16__2_,
         SUMB_16__1_, SUMB_16__0_, SUMB_15__6_, SUMB_15__5_, SUMB_15__4_,
         SUMB_15__3_, SUMB_15__2_, SUMB_15__1_, SUMB_14__6_, SUMB_14__5_,
         SUMB_14__4_, SUMB_14__3_, SUMB_14__2_, SUMB_14__1_, SUMB_13__6_,
         SUMB_13__5_, SUMB_13__4_, SUMB_13__3_, SUMB_13__2_, SUMB_13__1_,
         SUMB_12__6_, SUMB_12__5_, SUMB_12__4_, SUMB_12__3_, SUMB_12__2_,
         SUMB_12__1_, SUMB_11__6_, SUMB_11__5_, SUMB_11__4_, SUMB_11__3_,
         SUMB_11__2_, SUMB_11__1_, SUMB_10__6_, SUMB_10__5_, SUMB_10__4_,
         SUMB_10__3_, SUMB_10__2_, SUMB_10__1_, SUMB_9__6_, SUMB_9__5_,
         SUMB_9__4_, SUMB_9__3_, SUMB_9__2_, SUMB_9__1_, SUMB_8__6_,
         SUMB_8__5_, SUMB_8__4_, SUMB_8__3_, SUMB_8__2_, SUMB_8__1_,
         SUMB_7__6_, SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_,
         SUMB_7__1_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, PROD1_7_, A1_21_, A1_20_, A1_19_, A1_18_,
         A1_17_, A1_16_, A1_15_, A1_13_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_,
         A1_7_, A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79;

  ADDFHX4 S4_1 ( .A(ab_16__1_), .B(CARRYB_15__1_), .CI(SUMB_15__2_), .CO(
        CARRYB_16__1_), .S(SUMB_16__1_) );
  ADDFHX4 S2_15_2 ( .A(ab_15__2_), .B(CARRYB_14__2_), .CI(SUMB_14__3_), .CO(
        CARRYB_15__2_), .S(SUMB_15__2_) );
  ADDFHX4 S1_14_0 ( .A(ab_14__0_), .B(CARRYB_13__0_), .CI(SUMB_13__1_), .CO(
        CARRYB_14__0_), .S(A1_12_) );
  ADDFHX4 S2_14_2 ( .A(ab_14__2_), .B(CARRYB_13__2_), .CI(SUMB_13__3_), .CO(
        CARRYB_14__2_), .S(SUMB_14__2_) );
  ADDFHX4 S1_13_0 ( .A(ab_13__0_), .B(CARRYB_12__0_), .CI(SUMB_12__1_), .CO(
        CARRYB_13__0_), .S(A1_11_) );
  ADDFHX4 S2_13_1 ( .A(ab_13__1_), .B(CARRYB_12__1_), .CI(SUMB_12__2_), .CO(
        CARRYB_13__1_), .S(SUMB_13__1_) );
  ADDFHX4 S2_13_2 ( .A(ab_13__2_), .B(CARRYB_12__2_), .CI(SUMB_12__3_), .CO(
        CARRYB_13__2_), .S(SUMB_13__2_) );
  ADDFHX4 S1_12_0 ( .A(ab_12__0_), .B(CARRYB_11__0_), .CI(SUMB_11__1_), .CO(
        CARRYB_12__0_), .S(A1_10_) );
  ADDFHX4 S2_12_1 ( .A(ab_12__1_), .B(CARRYB_11__1_), .CI(SUMB_11__2_), .CO(
        CARRYB_12__1_), .S(SUMB_12__1_) );
  multi16_10_DW01_add_0 FS_1 ( .A_21_(A1_21_), .A_20_(A1_20_), .A_19_(A1_19_), 
        .A_18_(A1_18_), .A_17_(A1_17_), .A_16_(A1_16_), .A_15_(A1_15_), 
        .A_14_(SUMB_16__0_), .A_13_(A1_13_), .A_12_(A1_12_), .A_11_(A1_11_), 
        .A_10_(A1_10_), .A_9_(A1_9_), .A_8_(A1_8_), .A_7_(A1_7_), .A_6_(A1_6_), 
        .A_5_(PROD1_7_), .B_21_(n61), .B_20_(n60), .B_19_(n59), .B_18_(n56), 
        .B_17_(n57), .B_16_(n58), .SUM_21_(PRODUCT_23_), .SUM_20_(PRODUCT_22_), 
        .SUM_19_(PRODUCT_21_), .SUM_18_(PRODUCT_20_), .SUM_17_(PRODUCT_19_), 
        .SUM_16_(PRODUCT_18_), .SUM_15_(PRODUCT_17_), .SUM_14_(PRODUCT_16_), 
        .SUM_13_(PRODUCT_15_), .SUM_12_(PRODUCT_14_), .SUM_11_(PRODUCT_13_), 
        .SUM_10_(PRODUCT_12_), .SUM_9_(PRODUCT_11_), .SUM_8_(PRODUCT_10_), 
        .SUM_7_(PRODUCT_9_), .SUM_6_(PRODUCT_8_), .SUM_5_(PRODUCT_7_) );
  ADDFHX1 S2_14_5 ( .A(ab_14__5_), .B(CARRYB_13__5_), .CI(SUMB_13__6_), .CO(
        CARRYB_14__5_), .S(SUMB_14__5_) );
  ADDFHX1 S3_15_6 ( .A(ab_15__6_), .B(CARRYB_14__6_), .CI(ab_14__7_), .CO(
        CARRYB_15__6_), .S(SUMB_15__6_) );
  ADDFX2 S5_6 ( .A(ab_16__6_), .B(CARRYB_15__6_), .CI(ab_15__7_), .CO(
        CARRYB_16__6_), .S(SUMB_16__6_) );
  ADDFHX1 S2_15_5 ( .A(ab_15__5_), .B(CARRYB_14__5_), .CI(SUMB_14__6_), .CO(
        CARRYB_15__5_), .S(SUMB_15__5_) );
  ADDFHX1 S4_5 ( .A(ab_16__5_), .B(CARRYB_15__5_), .CI(SUMB_15__6_), .CO(
        CARRYB_16__5_), .S(SUMB_16__5_) );
  ADDFHX4 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  ADDFHX4 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  ADDFHX4 S1_8_0 ( .A(ab_8__0_), .B(CARRYB_7__0_), .CI(SUMB_7__1_), .CO(
        CARRYB_8__0_), .S(A1_6_) );
  ADDFHX4 S2_10_5 ( .A(ab_10__5_), .B(CARRYB_9__5_), .CI(SUMB_9__6_), .CO(
        CARRYB_10__5_), .S(SUMB_10__5_) );
  ADDFHX4 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  ADDFHX4 S2_11_3 ( .A(ab_11__3_), .B(CARRYB_10__3_), .CI(SUMB_10__4_), .CO(
        CARRYB_11__3_), .S(SUMB_11__3_) );
  ADDFHX4 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  ADDFHX4 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  ADDFHX4 S2_15_3 ( .A(ab_15__3_), .B(CARRYB_14__3_), .CI(SUMB_14__4_), .CO(
        CARRYB_15__3_), .S(SUMB_15__3_) );
  ADDFHX2 S3_11_6 ( .A(ab_11__6_), .B(CARRYB_10__6_), .CI(ab_10__7_), .CO(
        CARRYB_11__6_), .S(SUMB_11__6_) );
  ADDFHX4 S3_12_6 ( .A(ab_12__6_), .B(CARRYB_11__6_), .CI(ab_11__7_), .CO(
        CARRYB_12__6_), .S(SUMB_12__6_) );
  ADDFHX2 S3_13_6 ( .A(ab_13__6_), .B(CARRYB_12__6_), .CI(ab_12__7_), .CO(
        CARRYB_13__6_), .S(SUMB_13__6_) );
  ADDFHX4 S2_12_4 ( .A(ab_12__4_), .B(CARRYB_11__4_), .CI(SUMB_11__5_), .CO(
        CARRYB_12__4_), .S(SUMB_12__4_) );
  ADDFHX4 S3_9_6 ( .A(ab_9__6_), .B(CARRYB_8__6_), .CI(ab_8__7_), .CO(
        CARRYB_9__6_), .S(SUMB_9__6_) );
  ADDFHX2 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  ADDFHX4 S2_11_5 ( .A(ab_11__5_), .B(CARRYB_10__5_), .CI(SUMB_10__6_), .CO(
        CARRYB_11__5_), .S(SUMB_11__5_) );
  ADDFHX4 S2_8_2 ( .A(ab_8__2_), .B(CARRYB_7__2_), .CI(SUMB_7__3_), .CO(
        CARRYB_8__2_), .S(SUMB_8__2_) );
  ADDFHX4 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  ADDFHX4 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  ADDFHX4 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  ADDFHX4 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  ADDFHX4 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  ADDFHX4 S2_7_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  ADDFHX2 S2_13_3 ( .A(ab_13__3_), .B(CARRYB_12__3_), .CI(SUMB_12__4_), .CO(
        CARRYB_13__3_), .S(SUMB_13__3_) );
  ADDFHX4 S2_2_4 ( .A(ab_2__4_), .B(n22), .CI(SUMB_1__5_), .CO(CARRYB_2__4_), 
        .S(SUMB_2__4_) );
  ADDFHX4 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  ADDFHX4 S2_7_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  ADDFHX4 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  ADDFHX2 S4_4 ( .A(ab_16__4_), .B(CARRYB_15__4_), .CI(SUMB_15__5_), .CO(
        CARRYB_16__4_), .S(SUMB_16__4_) );
  ADDFHX4 S1_10_0 ( .A(ab_10__0_), .B(CARRYB_9__0_), .CI(SUMB_9__1_), .CO(
        CARRYB_10__0_), .S(A1_8_) );
  ADDFHX4 S2_9_2 ( .A(ab_9__2_), .B(CARRYB_8__2_), .CI(SUMB_8__3_), .CO(
        CARRYB_9__2_), .S(SUMB_9__2_) );
  ADDFHX4 S2_7_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  ADDFHX2 S4_2 ( .A(ab_16__2_), .B(CARRYB_15__2_), .CI(SUMB_15__3_), .CO(
        CARRYB_16__2_), .S(SUMB_16__2_) );
  ADDFHX2 S2_13_5 ( .A(ab_13__5_), .B(CARRYB_12__5_), .CI(SUMB_12__6_), .CO(
        CARRYB_13__5_), .S(SUMB_13__5_) );
  ADDFHX4 S2_7_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  ADDFHX4 S2_10_3 ( .A(ab_10__3_), .B(CARRYB_9__3_), .CI(SUMB_9__4_), .CO(
        CARRYB_10__3_), .S(SUMB_10__3_) );
  ADDFHX2 S3_7_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(
        CARRYB_7__6_), .S(SUMB_7__6_) );
  ADDFHX2 S2_15_4 ( .A(ab_15__4_), .B(CARRYB_14__4_), .CI(SUMB_14__5_), .CO(
        CARRYB_15__4_), .S(SUMB_15__4_) );
  ADDFHX2 S3_8_6 ( .A(ab_8__6_), .B(CARRYB_7__6_), .CI(ab_7__7_), .CO(
        CARRYB_8__6_), .S(SUMB_8__6_) );
  ADDFHX4 S2_14_4 ( .A(ab_14__4_), .B(CARRYB_13__4_), .CI(SUMB_13__5_), .CO(
        CARRYB_14__4_), .S(SUMB_14__4_) );
  ADDFHX4 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  ADDFHX4 S2_7_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  ADDFHX4 S2_11_1 ( .A(ab_11__1_), .B(CARRYB_10__1_), .CI(SUMB_10__2_), .CO(
        CARRYB_11__1_), .S(SUMB_11__1_) );
  ADDFHX4 S2_8_5 ( .A(ab_8__5_), .B(CARRYB_7__5_), .CI(SUMB_7__6_), .CO(
        CARRYB_8__5_), .S(SUMB_8__5_) );
  ADDFHX4 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  ADDFHX4 S2_10_4 ( .A(ab_10__4_), .B(CARRYB_9__4_), .CI(SUMB_9__5_), .CO(
        CARRYB_10__4_), .S(SUMB_10__4_) );
  ADDFHX4 S2_11_4 ( .A(ab_11__4_), .B(CARRYB_10__4_), .CI(SUMB_10__5_), .CO(
        CARRYB_11__4_), .S(SUMB_11__4_) );
  ADDFHX4 S2_9_5 ( .A(ab_9__5_), .B(CARRYB_8__5_), .CI(SUMB_8__6_), .CO(
        CARRYB_9__5_), .S(SUMB_9__5_) );
  ADDFHX2 S2_2_1 ( .A(ab_2__1_), .B(n24), .CI(SUMB_1__2_), .CO(CARRYB_2__1_), 
        .S(SUMB_2__1_) );
  ADDFHX4 S2_14_1 ( .A(ab_14__1_), .B(CARRYB_13__1_), .CI(SUMB_13__2_), .CO(
        CARRYB_14__1_), .S(SUMB_14__1_) );
  ADDFHX4 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  ADDFHX2 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  ADDFHX1 S3_14_6 ( .A(ab_14__6_), .B(CARRYB_13__6_), .CI(ab_13__7_), .CO(
        CARRYB_14__6_), .S(SUMB_14__6_) );
  ADDFHX2 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  ADDFHX2 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  ADDFHX2 S2_12_5 ( .A(ab_12__5_), .B(CARRYB_11__5_), .CI(SUMB_11__6_), .CO(
        CARRYB_12__5_), .S(SUMB_12__5_) );
  ADDFHX2 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  ADDFHX2 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  ADDFHX2 S2_8_1 ( .A(ab_8__1_), .B(CARRYB_7__1_), .CI(SUMB_7__2_), .CO(
        CARRYB_8__1_), .S(SUMB_8__1_) );
  ADDFHX2 S2_13_4 ( .A(ab_13__4_), .B(CARRYB_12__4_), .CI(SUMB_12__5_), .CO(
        CARRYB_13__4_), .S(SUMB_13__4_) );
  ADDFHX2 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  ADDFHX4 S4_3 ( .A(ab_16__3_), .B(CARRYB_15__3_), .CI(SUMB_15__4_), .CO(
        CARRYB_16__3_), .S(SUMB_16__3_) );
  ADDFHX4 S2_12_3 ( .A(ab_12__3_), .B(CARRYB_11__3_), .CI(SUMB_11__4_), .CO(
        CARRYB_12__3_), .S(SUMB_12__3_) );
  ADDFHX4 S2_10_2 ( .A(ab_10__2_), .B(CARRYB_9__2_), .CI(SUMB_9__3_), .CO(
        CARRYB_10__2_), .S(SUMB_10__2_) );
  ADDFHX4 S1_7_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(PROD1_7_) );
  ADDFHX4 S1_9_0 ( .A(ab_9__0_), .B(CARRYB_8__0_), .CI(SUMB_8__1_), .CO(
        CARRYB_9__0_), .S(A1_7_) );
  ADDFHX4 S1_11_0 ( .A(ab_11__0_), .B(CARRYB_10__0_), .CI(SUMB_10__1_), .CO(
        CARRYB_11__0_), .S(A1_9_) );
  ADDFHX4 S3_10_6 ( .A(ab_10__6_), .B(CARRYB_9__6_), .CI(ab_9__7_), .CO(
        CARRYB_10__6_), .S(SUMB_10__6_) );
  ADDFHX4 S3_2_6 ( .A(ab_2__6_), .B(n20), .CI(ab_1__7_), .CO(CARRYB_2__6_), 
        .S(SUMB_2__6_) );
  ADDFHX4 S2_2_5 ( .A(ab_2__5_), .B(n21), .CI(SUMB_1__6_), .CO(CARRYB_2__5_), 
        .S(SUMB_2__5_) );
  ADDFHX4 S1_2_0 ( .A(ab_2__0_), .B(n17), .CI(SUMB_1__1_), .CO(CARRYB_2__0_), 
        .S(A1_0_) );
  ADDFHX4 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  ADDFHX4 S2_2_3 ( .A(ab_2__3_), .B(n23), .CI(SUMB_1__4_), .CO(CARRYB_2__3_), 
        .S(SUMB_2__3_) );
  ADDFHX4 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  ADDFHX4 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  ADDFHX4 S2_8_4 ( .A(ab_8__4_), .B(CARRYB_7__4_), .CI(SUMB_7__5_), .CO(
        CARRYB_8__4_), .S(SUMB_8__4_) );
  ADDFHX4 S1_15_0 ( .A(ab_15__0_), .B(CARRYB_14__0_), .CI(SUMB_14__1_), .CO(
        CARRYB_15__0_), .S(A1_13_) );
  ADDFHX4 S4_0 ( .A(ab_16__0_), .B(CARRYB_15__0_), .CI(SUMB_15__1_), .CO(
        CARRYB_16__0_), .S(SUMB_16__0_) );
  ADDFHX4 S2_9_1 ( .A(ab_9__1_), .B(CARRYB_8__1_), .CI(SUMB_8__2_), .CO(
        CARRYB_9__1_), .S(SUMB_9__1_) );
  AND2X4 U2 ( .A(ab_0__4_), .B(ab_1__3_), .Y(n23) );
  AND2X4 U3 ( .A(ab_0__6_), .B(ab_1__5_), .Y(n21) );
  XOR3X2 U4 ( .A(ab_8__3_), .B(CARRYB_7__3_), .C(SUMB_7__4_), .Y(SUMB_8__3_)
         );
  NAND3X4 U5 ( .A(n6), .B(n4), .C(n5), .Y(CARRYB_15__1_) );
  NAND3X2 U6 ( .A(n37), .B(n35), .C(n36), .Y(CARRYB_2__2_) );
  NAND2X2 U7 ( .A(SUMB_1__3_), .B(n19), .Y(n37) );
  NAND2X2 U8 ( .A(SUMB_1__3_), .B(ab_2__2_), .Y(n36) );
  AND2X4 U9 ( .A(CARRYB_16__0_), .B(SUMB_16__1_), .Y(n58) );
  AND2X2 U10 ( .A(A[2]), .B(B[6]), .Y(ab_2__6_) );
  XOR2X4 U11 ( .A(CARRYB_9__1_), .B(n52), .Y(SUMB_10__1_) );
  NAND2X1 U12 ( .A(SUMB_8__4_), .B(CARRYB_8__3_), .Y(n13) );
  NAND2XL U13 ( .A(SUMB_5__4_), .B(CARRYB_5__3_), .Y(n25) );
  NAND2XL U14 ( .A(ab_6__3_), .B(CARRYB_5__3_), .Y(n26) );
  NAND2XL U15 ( .A(A[1]), .B(B[1]), .Y(n64) );
  XOR2X4 U16 ( .A(SUMB_14__2_), .B(ab_15__1_), .Y(n3) );
  XOR2X2 U17 ( .A(CARRYB_14__1_), .B(n3), .Y(SUMB_15__1_) );
  NAND2X2 U18 ( .A(SUMB_14__2_), .B(CARRYB_14__1_), .Y(n4) );
  NAND2X2 U19 ( .A(ab_15__1_), .B(CARRYB_14__1_), .Y(n5) );
  NAND2XL U20 ( .A(ab_15__1_), .B(SUMB_14__2_), .Y(n6) );
  NOR2X4 U21 ( .A(n74), .B(n70), .Y(ab_15__1_) );
  NAND2X2 U22 ( .A(ab_8__3_), .B(CARRYB_7__3_), .Y(n7) );
  NAND2X2 U23 ( .A(ab_8__3_), .B(SUMB_7__4_), .Y(n8) );
  NAND2X2 U24 ( .A(CARRYB_7__3_), .B(SUMB_7__4_), .Y(n9) );
  NAND3X4 U25 ( .A(n7), .B(n8), .C(n9), .Y(CARRYB_8__3_) );
  XOR2X2 U26 ( .A(ab_9__3_), .B(SUMB_8__4_), .Y(n10) );
  XOR2X2 U27 ( .A(n10), .B(CARRYB_8__3_), .Y(SUMB_9__3_) );
  NAND2XL U28 ( .A(ab_9__3_), .B(SUMB_8__4_), .Y(n11) );
  NAND2X2 U29 ( .A(ab_9__3_), .B(CARRYB_8__3_), .Y(n12) );
  NAND3X2 U30 ( .A(n11), .B(n12), .C(n13), .Y(CARRYB_9__3_) );
  XOR3X4 U31 ( .A(CARRYB_11__2_), .B(ab_12__2_), .C(SUMB_11__3_), .Y(
        SUMB_12__2_) );
  NAND2X2 U32 ( .A(SUMB_11__3_), .B(CARRYB_11__2_), .Y(n14) );
  NAND2X2 U33 ( .A(ab_12__2_), .B(CARRYB_11__2_), .Y(n15) );
  NAND2X2 U34 ( .A(ab_12__2_), .B(SUMB_11__3_), .Y(n16) );
  NAND3X4 U35 ( .A(n16), .B(n14), .C(n15), .Y(CARRYB_12__2_) );
  AND2X1 U36 ( .A(A[2]), .B(B[2]), .Y(ab_2__2_) );
  NAND3X2 U37 ( .A(n44), .B(n42), .C(n43), .Y(CARRYB_14__3_) );
  AND2X2 U38 ( .A(A[1]), .B(B[4]), .Y(ab_1__4_) );
  AND2X1 U39 ( .A(A[1]), .B(B[2]), .Y(ab_1__2_) );
  BUFX3 U40 ( .A(CARRYB_1__0_), .Y(n17) );
  NAND3X4 U41 ( .A(n48), .B(n46), .C(n47), .Y(CARRYB_4__6_) );
  NAND2X2 U42 ( .A(ab_4__6_), .B(CARRYB_3__6_), .Y(n46) );
  INVX4 U43 ( .A(B[4]), .Y(n67) );
  AND2X2 U44 ( .A(A[2]), .B(B[4]), .Y(ab_2__4_) );
  AND2X1 U45 ( .A(A[3]), .B(B[4]), .Y(ab_3__4_) );
  NOR2X4 U46 ( .A(n71), .B(n62), .Y(ab_0__7_) );
  INVX4 U47 ( .A(B[7]), .Y(n71) );
  NOR2X4 U48 ( .A(n65), .B(n62), .Y(ab_0__6_) );
  INVX4 U49 ( .A(B[6]), .Y(n65) );
  INVX1 U50 ( .A(A[0]), .Y(n62) );
  NOR2X1 U51 ( .A(n68), .B(n62), .Y(ab_0__3_) );
  NOR2X1 U52 ( .A(n78), .B(n69), .Y(ab_11__2_) );
  INVX1 U53 ( .A(B[2]), .Y(n69) );
  INVX1 U54 ( .A(B[5]), .Y(n66) );
  AND2X2 U56 ( .A(ab_0__3_), .B(ab_1__2_), .Y(n19) );
  AND2X2 U57 ( .A(ab_0__7_), .B(ab_1__6_), .Y(n20) );
  AND2X2 U58 ( .A(ab_0__5_), .B(ab_1__4_), .Y(n22) );
  AND2X2 U59 ( .A(ab_0__2_), .B(n72), .Y(n24) );
  AND2X1 U60 ( .A(CARRYB_16__4_), .B(SUMB_16__5_), .Y(n60) );
  AND2X1 U61 ( .A(A[9]), .B(B[6]), .Y(ab_9__6_) );
  AND2X1 U62 ( .A(A[8]), .B(B[6]), .Y(ab_8__6_) );
  NAND3X2 U63 ( .A(n51), .B(n49), .C(n50), .Y(CARRYB_6__5_) );
  NAND2X1 U64 ( .A(SUMB_16__2_), .B(n29), .Y(n30) );
  CLKINVX2 U65 ( .A(SUMB_16__2_), .Y(n28) );
  XOR2X2 U66 ( .A(ab_1__5_), .B(ab_0__6_), .Y(SUMB_1__5_) );
  XOR3X4 U67 ( .A(CARRYB_5__3_), .B(ab_6__3_), .C(SUMB_5__4_), .Y(SUMB_6__3_)
         );
  NAND2X1 U68 ( .A(ab_6__3_), .B(SUMB_5__4_), .Y(n27) );
  NAND3X2 U69 ( .A(n27), .B(n25), .C(n26), .Y(CARRYB_6__3_) );
  AND2X2 U70 ( .A(A[6]), .B(B[3]), .Y(ab_6__3_) );
  NAND2X1 U71 ( .A(n28), .B(CARRYB_16__1_), .Y(n31) );
  NAND2X2 U72 ( .A(n30), .B(n31), .Y(A1_16_) );
  CLKINVX2 U73 ( .A(CARRYB_16__1_), .Y(n29) );
  AND2X2 U74 ( .A(A[2]), .B(B[1]), .Y(ab_2__1_) );
  XOR2X4 U75 ( .A(CARRYB_16__2_), .B(SUMB_16__3_), .Y(A1_17_) );
  XOR3X4 U76 ( .A(CARRYB_10__2_), .B(ab_11__2_), .C(SUMB_10__3_), .Y(
        SUMB_11__2_) );
  NAND2X2 U77 ( .A(SUMB_10__3_), .B(CARRYB_10__2_), .Y(n32) );
  NAND2X1 U78 ( .A(ab_11__2_), .B(CARRYB_10__2_), .Y(n33) );
  NAND2X2 U79 ( .A(ab_11__2_), .B(SUMB_10__3_), .Y(n34) );
  NAND3X4 U80 ( .A(n34), .B(n32), .C(n33), .Y(CARRYB_11__2_) );
  XOR3X2 U81 ( .A(ab_2__2_), .B(SUMB_1__3_), .C(n19), .Y(SUMB_2__2_) );
  NAND2XL U82 ( .A(n19), .B(ab_2__2_), .Y(n35) );
  XOR2X4 U83 ( .A(ab_1__3_), .B(ab_0__4_), .Y(SUMB_1__3_) );
  XOR3X4 U84 ( .A(CARRYB_8__4_), .B(ab_9__4_), .C(SUMB_8__5_), .Y(SUMB_9__4_)
         );
  NAND2X1 U85 ( .A(SUMB_8__5_), .B(CARRYB_8__4_), .Y(n38) );
  NAND2X1 U86 ( .A(ab_9__4_), .B(CARRYB_8__4_), .Y(n39) );
  NAND2X2 U87 ( .A(ab_9__4_), .B(SUMB_8__5_), .Y(n40) );
  NAND3X4 U88 ( .A(n40), .B(n38), .C(n39), .Y(CARRYB_9__4_) );
  XOR2X2 U89 ( .A(CARRYB_13__3_), .B(n41), .Y(SUMB_14__3_) );
  AND2X2 U90 ( .A(CARRYB_16__1_), .B(SUMB_16__2_), .Y(n57) );
  NAND2X1 U91 ( .A(ab_10__1_), .B(SUMB_9__2_), .Y(n55) );
  XOR2X4 U92 ( .A(SUMB_13__4_), .B(ab_14__3_), .Y(n41) );
  NAND2XL U93 ( .A(ab_3__7_), .B(ab_4__6_), .Y(n48) );
  AND2X1 U94 ( .A(A[4]), .B(B[0]), .Y(ab_4__0_) );
  AND2X1 U95 ( .A(A[4]), .B(B[1]), .Y(ab_4__1_) );
  XOR2X1 U96 ( .A(ab_4__6_), .B(ab_3__7_), .Y(n45) );
  XOR2X4 U97 ( .A(SUMB_9__2_), .B(ab_10__1_), .Y(n52) );
  NAND2X2 U98 ( .A(SUMB_9__2_), .B(CARRYB_9__1_), .Y(n53) );
  NAND2X2 U99 ( .A(ab_10__1_), .B(CARRYB_9__1_), .Y(n54) );
  AND2X2 U100 ( .A(A[2]), .B(B[3]), .Y(ab_2__3_) );
  XOR2X1 U101 ( .A(n72), .B(ab_0__2_), .Y(SUMB_1__1_) );
  AND2X2 U102 ( .A(A[2]), .B(B[5]), .Y(ab_2__5_) );
  NAND2X1 U103 ( .A(ab_6__5_), .B(CARRYB_5__5_), .Y(n50) );
  NAND2X1 U104 ( .A(SUMB_5__6_), .B(CARRYB_5__5_), .Y(n49) );
  XOR2X2 U105 ( .A(CARRYB_16__3_), .B(SUMB_16__4_), .Y(A1_18_) );
  NAND2X1 U106 ( .A(SUMB_13__4_), .B(CARRYB_13__3_), .Y(n42) );
  NAND2X1 U107 ( .A(ab_14__3_), .B(CARRYB_13__3_), .Y(n43) );
  NAND2X1 U108 ( .A(ab_14__3_), .B(SUMB_13__4_), .Y(n44) );
  XOR2X1 U109 ( .A(CARRYB_3__6_), .B(n45), .Y(SUMB_4__6_) );
  NAND2X2 U110 ( .A(ab_3__7_), .B(CARRYB_3__6_), .Y(n47) );
  XOR3X4 U111 ( .A(CARRYB_5__5_), .B(ab_6__5_), .C(SUMB_5__6_), .Y(SUMB_6__5_)
         );
  NAND2XL U112 ( .A(ab_6__5_), .B(SUMB_5__6_), .Y(n51) );
  NAND3X4 U113 ( .A(n55), .B(n53), .C(n54), .Y(CARRYB_10__1_) );
  AND2X1 U114 ( .A(A[3]), .B(B[6]), .Y(ab_3__6_) );
  AND2X1 U115 ( .A(A[5]), .B(B[6]), .Y(ab_5__6_) );
  AND2X1 U116 ( .A(CARRYB_16__2_), .B(SUMB_16__3_), .Y(n56) );
  AND2X1 U117 ( .A(A[10]), .B(B[1]), .Y(ab_10__1_) );
  AND2X1 U118 ( .A(A[9]), .B(B[1]), .Y(ab_9__1_) );
  AND2X1 U119 ( .A(A[7]), .B(B[1]), .Y(ab_7__1_) );
  AND2X1 U120 ( .A(A[8]), .B(B[0]), .Y(ab_8__0_) );
  AND2X1 U121 ( .A(A[10]), .B(B[0]), .Y(ab_10__0_) );
  INVXL U122 ( .A(B[3]), .Y(n68) );
  AND2X1 U123 ( .A(CARRYB_16__5_), .B(SUMB_16__6_), .Y(n61) );
  INVXL U124 ( .A(B[0]), .Y(n79) );
  INVXL U125 ( .A(B[1]), .Y(n70) );
  AND2X2 U126 ( .A(A[1]), .B(B[3]), .Y(ab_1__3_) );
  AND2X1 U127 ( .A(A[7]), .B(B[6]), .Y(ab_7__6_) );
  AND2X1 U128 ( .A(A[10]), .B(B[6]), .Y(ab_10__6_) );
  AND2X1 U129 ( .A(A[6]), .B(B[6]), .Y(ab_6__6_) );
  NOR2XL U130 ( .A(n78), .B(n70), .Y(ab_11__1_) );
  NOR2XL U131 ( .A(n76), .B(n70), .Y(ab_13__1_) );
  NOR2XL U132 ( .A(n77), .B(n70), .Y(ab_12__1_) );
  AND2X1 U133 ( .A(A[3]), .B(B[0]), .Y(ab_3__0_) );
  XOR2X1 U134 ( .A(CARRYB_16__6_), .B(ab_16__7_), .Y(A1_21_) );
  NOR2X1 U135 ( .A(n73), .B(n70), .Y(ab_16__1_) );
  NOR2X1 U136 ( .A(n73), .B(n68), .Y(ab_16__3_) );
  INVX1 U137 ( .A(n64), .Y(n72) );
  AND2X2 U138 ( .A(A[8]), .B(B[1]), .Y(ab_8__1_) );
  AND2X2 U139 ( .A(A[6]), .B(B[1]), .Y(ab_6__1_) );
  AND2X2 U140 ( .A(A[9]), .B(B[0]), .Y(ab_9__0_) );
  AND2X2 U141 ( .A(A[5]), .B(B[1]), .Y(ab_5__1_) );
  AND2X2 U142 ( .A(A[5]), .B(B[0]), .Y(ab_5__0_) );
  AND2X2 U143 ( .A(A[7]), .B(B[0]), .Y(ab_7__0_) );
  AND2X2 U144 ( .A(A[6]), .B(B[0]), .Y(ab_6__0_) );
  XOR2X1 U145 ( .A(CARRYB_16__4_), .B(SUMB_16__5_), .Y(A1_19_) );
  XOR2X1 U146 ( .A(CARRYB_16__5_), .B(SUMB_16__6_), .Y(A1_20_) );
  AND2X2 U147 ( .A(CARRYB_16__3_), .B(SUMB_16__4_), .Y(n59) );
  NOR2X1 U148 ( .A(n73), .B(n71), .Y(ab_16__7_) );
  NOR2X2 U149 ( .A(n67), .B(n62), .Y(ab_0__4_) );
  NOR2X1 U150 ( .A(n66), .B(n62), .Y(ab_0__5_) );
  NOR2XL U151 ( .A(n73), .B(n67), .Y(ab_16__4_) );
  NOR2X1 U152 ( .A(n74), .B(n71), .Y(ab_15__7_) );
  NOR2X1 U153 ( .A(n73), .B(n65), .Y(ab_16__6_) );
  NOR2X1 U154 ( .A(n75), .B(n70), .Y(ab_14__1_) );
  NOR2XL U155 ( .A(n76), .B(n68), .Y(ab_13__3_) );
  NOR2XL U156 ( .A(n77), .B(n68), .Y(ab_12__3_) );
  NOR2XL U157 ( .A(n74), .B(n68), .Y(ab_15__3_) );
  NOR2XL U158 ( .A(n78), .B(n68), .Y(ab_11__3_) );
  NOR2XL U159 ( .A(n75), .B(n68), .Y(ab_14__3_) );
  AND2X1 U160 ( .A(A[10]), .B(B[3]), .Y(ab_10__3_) );
  AND2X1 U161 ( .A(A[9]), .B(B[3]), .Y(ab_9__3_) );
  AND2X1 U162 ( .A(A[8]), .B(B[3]), .Y(ab_8__3_) );
  NOR2XL U163 ( .A(n75), .B(n67), .Y(ab_14__4_) );
  NOR2XL U164 ( .A(n77), .B(n67), .Y(ab_12__4_) );
  AND2X1 U165 ( .A(A[7]), .B(B[3]), .Y(ab_7__3_) );
  NOR2XL U166 ( .A(n78), .B(n67), .Y(ab_11__4_) );
  NOR2XL U167 ( .A(n76), .B(n67), .Y(ab_13__4_) );
  AND2X1 U168 ( .A(A[3]), .B(B[3]), .Y(ab_3__3_) );
  AND2X1 U169 ( .A(A[3]), .B(B[1]), .Y(ab_3__1_) );
  AND2X1 U170 ( .A(A[4]), .B(B[3]), .Y(ab_4__3_) );
  AND2X1 U171 ( .A(A[5]), .B(B[3]), .Y(ab_5__3_) );
  NOR2XL U172 ( .A(n78), .B(n71), .Y(ab_11__7_) );
  AND2X1 U173 ( .A(A[9]), .B(B[7]), .Y(ab_9__7_) );
  NOR2XL U174 ( .A(n76), .B(n71), .Y(ab_13__7_) );
  AND2X1 U175 ( .A(A[10]), .B(B[7]), .Y(ab_10__7_) );
  AND2X1 U176 ( .A(A[8]), .B(B[7]), .Y(ab_8__7_) );
  AND2X1 U177 ( .A(A[7]), .B(B[7]), .Y(ab_7__7_) );
  AND2X1 U178 ( .A(A[6]), .B(B[7]), .Y(ab_6__7_) );
  AND2X1 U179 ( .A(A[3]), .B(B[7]), .Y(ab_3__7_) );
  AND2X1 U180 ( .A(A[4]), .B(B[6]), .Y(ab_4__6_) );
  AND2X1 U181 ( .A(A[4]), .B(B[7]), .Y(ab_4__7_) );
  AND2X1 U182 ( .A(A[5]), .B(B[7]), .Y(ab_5__7_) );
  NOR2XL U183 ( .A(n64), .B(n63), .Y(CARRYB_1__0_) );
  XOR2X1 U184 ( .A(ab_1__2_), .B(ab_0__3_), .Y(SUMB_1__2_) );
  XOR2X1 U185 ( .A(ab_1__4_), .B(ab_0__5_), .Y(SUMB_1__4_) );
  NOR2XL U186 ( .A(n75), .B(n71), .Y(ab_14__7_) );
  NOR2XL U187 ( .A(n77), .B(n71), .Y(ab_12__7_) );
  AND2X1 U188 ( .A(A[2]), .B(B[7]), .Y(ab_2__7_) );
  NOR2XL U189 ( .A(n74), .B(n67), .Y(ab_15__4_) );
  AND2X2 U190 ( .A(A[2]), .B(B[0]), .Y(ab_2__0_) );
  INVX1 U191 ( .A(A[16]), .Y(n73) );
  AND2X1 U192 ( .A(A[10]), .B(B[4]), .Y(ab_10__4_) );
  AND2X1 U193 ( .A(A[9]), .B(B[4]), .Y(ab_9__4_) );
  AND2X1 U194 ( .A(A[8]), .B(B[4]), .Y(ab_8__4_) );
  AND2X1 U195 ( .A(A[7]), .B(B[4]), .Y(ab_7__4_) );
  AND2X1 U196 ( .A(A[6]), .B(B[4]), .Y(ab_6__4_) );
  AND2X1 U197 ( .A(A[4]), .B(B[4]), .Y(ab_4__4_) );
  AND2X1 U198 ( .A(A[5]), .B(B[4]), .Y(ab_5__4_) );
  NAND2XL U199 ( .A(A[0]), .B(B[0]), .Y(n63) );
  XOR2X1 U200 ( .A(ab_1__6_), .B(ab_0__7_), .Y(SUMB_1__6_) );
  INVX1 U201 ( .A(A[11]), .Y(n78) );
  INVX1 U202 ( .A(A[12]), .Y(n77) );
  INVX1 U203 ( .A(A[13]), .Y(n76) );
  INVX1 U204 ( .A(A[14]), .Y(n75) );
  INVX1 U205 ( .A(A[15]), .Y(n74) );
  XOR2X4 U206 ( .A(CARRYB_16__0_), .B(SUMB_16__1_), .Y(A1_15_) );
  NOR2XL U207 ( .A(n78), .B(n65), .Y(ab_11__6_) );
  NOR2XL U208 ( .A(n77), .B(n65), .Y(ab_12__6_) );
  NOR2XL U209 ( .A(n76), .B(n65), .Y(ab_13__6_) );
  NOR2XL U210 ( .A(n75), .B(n65), .Y(ab_14__6_) );
  NOR2XL U211 ( .A(n74), .B(n65), .Y(ab_15__6_) );
  NOR2XL U212 ( .A(n73), .B(n66), .Y(ab_16__5_) );
  NOR2XL U213 ( .A(n74), .B(n66), .Y(ab_15__5_) );
  NOR2XL U214 ( .A(n75), .B(n66), .Y(ab_14__5_) );
  NOR2XL U215 ( .A(n76), .B(n66), .Y(ab_13__5_) );
  NOR2XL U216 ( .A(n77), .B(n66), .Y(ab_12__5_) );
  NOR2XL U217 ( .A(n78), .B(n66), .Y(ab_11__5_) );
  AND2X1 U218 ( .A(A[10]), .B(B[5]), .Y(ab_10__5_) );
  AND2X1 U219 ( .A(A[9]), .B(B[5]), .Y(ab_9__5_) );
  AND2X1 U220 ( .A(A[8]), .B(B[5]), .Y(ab_8__5_) );
  AND2X1 U221 ( .A(A[7]), .B(B[5]), .Y(ab_7__5_) );
  AND2X1 U222 ( .A(A[6]), .B(B[5]), .Y(ab_6__5_) );
  AND2X1 U223 ( .A(A[5]), .B(B[5]), .Y(ab_5__5_) );
  AND2X1 U224 ( .A(A[4]), .B(B[5]), .Y(ab_4__5_) );
  AND2X1 U225 ( .A(A[3]), .B(B[5]), .Y(ab_3__5_) );
  AND2X2 U226 ( .A(A[1]), .B(B[5]), .Y(ab_1__5_) );
  NOR2X2 U227 ( .A(n69), .B(n62), .Y(ab_0__2_) );
  NOR2XL U228 ( .A(n73), .B(n69), .Y(ab_16__2_) );
  NOR2XL U229 ( .A(n74), .B(n69), .Y(ab_15__2_) );
  NOR2XL U230 ( .A(n75), .B(n69), .Y(ab_14__2_) );
  NOR2XL U231 ( .A(n76), .B(n69), .Y(ab_13__2_) );
  NOR2XL U232 ( .A(n77), .B(n69), .Y(ab_12__2_) );
  AND2X1 U233 ( .A(A[1]), .B(B[7]), .Y(ab_1__7_) );
  AND2X2 U234 ( .A(A[1]), .B(B[6]), .Y(ab_1__6_) );
  AND2X1 U235 ( .A(A[10]), .B(B[2]), .Y(ab_10__2_) );
  AND2X1 U236 ( .A(A[9]), .B(B[2]), .Y(ab_9__2_) );
  AND2X1 U237 ( .A(A[8]), .B(B[2]), .Y(ab_8__2_) );
  AND2X1 U238 ( .A(A[7]), .B(B[2]), .Y(ab_7__2_) );
  AND2X1 U239 ( .A(A[6]), .B(B[2]), .Y(ab_6__2_) );
  AND2X1 U240 ( .A(A[5]), .B(B[2]), .Y(ab_5__2_) );
  AND2X1 U241 ( .A(A[4]), .B(B[2]), .Y(ab_4__2_) );
  AND2X1 U242 ( .A(A[3]), .B(B[2]), .Y(ab_3__2_) );
  NOR2X1 U244 ( .A(n79), .B(n73), .Y(ab_16__0_) );
  NOR2X1 U245 ( .A(n79), .B(n74), .Y(ab_15__0_) );
  NOR2X1 U246 ( .A(n79), .B(n75), .Y(ab_14__0_) );
  NOR2X1 U247 ( .A(n79), .B(n76), .Y(ab_13__0_) );
  NOR2X1 U248 ( .A(n79), .B(n77), .Y(ab_12__0_) );
  NOR2X1 U249 ( .A(n79), .B(n78), .Y(ab_11__0_) );
endmodule


module multi16_10 ( in_17bit, in_8bit, out );
  input [16:0] in_17bit;
  input [7:0] in_8bit;
  output [16:0] out;
  wire   N18, N19, N20, N21, N32, N33, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n55, n56, n57, n58, n59, n60, n61, n63, n64, n65, n66, n67, n68,
         n69, n71, n72, n73, n74, n75, n76, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n133,
         n134, n135, n136;
  wire   [16:1] in_17bit_b;
  wire   [6:0] in_8bit_b;
  wire   [23:8] mul;
  wire   [16:12] sub_add_52_b0_carry;

  multi16_10_DW02_mult_0 mult_55 ( .A({in_17bit_b, in_17bit[0]}), .B({n22, n23, 
        n8, in_8bit_b[4:0]}), .PRODUCT_23_(mul[23]), .PRODUCT_22_(mul[22]), 
        .PRODUCT_21_(mul[21]), .PRODUCT_20_(mul[20]), .PRODUCT_19_(mul[19]), 
        .PRODUCT_18_(mul[18]), .PRODUCT_17_(mul[17]), .PRODUCT_16_(mul[16]), 
        .PRODUCT_15_(mul[15]), .PRODUCT_14_(mul[14]), .PRODUCT_13_(mul[13]), 
        .PRODUCT_12_(mul[12]), .PRODUCT_11_(mul[11]), .PRODUCT_10_(mul[10]), 
        .PRODUCT_9_(mul[9]), .PRODUCT_8_(mul[8]), .PRODUCT_7_(N32) );
  NAND2X2 U2 ( .A(n3), .B(n28), .Y(n6) );
  INVX1 U3 ( .A(n120), .Y(n123) );
  INVX2 U4 ( .A(n116), .Y(n11) );
  NAND2X2 U5 ( .A(n21), .B(n136), .Y(n116) );
  NAND2X2 U6 ( .A(n19), .B(n20), .Y(n21) );
  NOR2X2 U7 ( .A(n123), .B(n25), .Y(n121) );
  NOR2XL U8 ( .A(in_8bit[4]), .B(in_8bit[1]), .Y(n1) );
  NOR2X2 U9 ( .A(n2), .B(n48), .Y(n49) );
  CLKINVX3 U10 ( .A(n1), .Y(n2) );
  NAND2BX2 U11 ( .AN(in_8bit[0]), .B(n47), .Y(n48) );
  NAND3BX1 U12 ( .AN(in_8bit[2]), .B(n50), .C(n49), .Y(n51) );
  NAND2X2 U13 ( .A(in_17bit[2]), .B(n4), .Y(n5) );
  NAND2X4 U14 ( .A(n5), .B(n6), .Y(in_17bit_b[2]) );
  INVXL U15 ( .A(in_17bit[2]), .Y(n3) );
  INVX2 U16 ( .A(n28), .Y(n4) );
  NAND2BXL U17 ( .AN(in_17bit[2]), .B(n32), .Y(n55) );
  NAND2BXL U18 ( .AN(mul[21]), .B(n119), .Y(n120) );
  NOR3BX2 U19 ( .AN(n53), .B(n52), .C(n32), .Y(in_17bit_b[1]) );
  INVX2 U20 ( .A(in_8bit_b[5]), .Y(n7) );
  CLKINVX4 U21 ( .A(n7), .Y(n8) );
  XOR2X2 U22 ( .A(n43), .B(in_8bit[4]), .Y(in_8bit_b[4]) );
  OR3X1 U23 ( .A(in_8bit[6]), .B(n34), .C(n51), .Y(n9) );
  INVXL U24 ( .A(in_8bit[0]), .Y(n38) );
  NOR2X1 U25 ( .A(in_17bit[1]), .B(in_17bit[16]), .Y(n52) );
  NAND3XL U26 ( .A(in_17bit[0]), .B(in_17bit[16]), .C(in_17bit[1]), .Y(n53) );
  XNOR2X1 U27 ( .A(n61), .B(n63), .Y(in_17bit_b[5]) );
  NOR2XL U28 ( .A(n36), .B(n64), .Y(n61) );
  NAND2BX1 U29 ( .AN(in_8bit[1]), .B(n38), .Y(n39) );
  XOR2X2 U30 ( .A(n40), .B(n47), .Y(in_8bit_b[3]) );
  OAI21XL U31 ( .A0(in_8bit[2]), .A1(n39), .B0(n33), .Y(n40) );
  XOR2X2 U32 ( .A(in_8bit[2]), .B(n26), .Y(in_8bit_b[2]) );
  NOR2XL U33 ( .A(n34), .B(n41), .Y(n26) );
  INVX1 U34 ( .A(N32), .Y(n126) );
  BUFX3 U35 ( .A(mul[18]), .Y(n18) );
  BUFX3 U36 ( .A(in_8bit_b[6]), .Y(n23) );
  CLKINVX2 U37 ( .A(n9), .Y(n22) );
  AOI21X1 U38 ( .A0(n42), .A1(n41), .B0(n34), .Y(n43) );
  NAND2BX1 U39 ( .AN(mul[12]), .B(n98), .Y(n99) );
  NOR2X1 U40 ( .A(mul[15]), .B(n105), .Y(n24) );
  XNOR2X1 U41 ( .A(n46), .B(n50), .Y(in_8bit_b[5]) );
  INVX1 U42 ( .A(mul[8]), .Y(n125) );
  INVX4 U43 ( .A(n112), .Y(n114) );
  INVX1 U44 ( .A(n117), .Y(n20) );
  INVX1 U45 ( .A(mul[19]), .Y(n19) );
  NAND2X2 U46 ( .A(n12), .B(n13), .Y(out[13]) );
  NAND2X1 U47 ( .A(mul[20]), .B(n116), .Y(n12) );
  NAND2X2 U48 ( .A(n10), .B(n11), .Y(n13) );
  INVX1 U49 ( .A(mul[20]), .Y(n10) );
  CLKINVX3 U50 ( .A(n34), .Y(n33) );
  INVX1 U51 ( .A(in_8bit[1]), .Y(n35) );
  INVX1 U52 ( .A(n25), .Y(n136) );
  INVX2 U53 ( .A(in_17bit[16]), .Y(n36) );
  NAND2X1 U54 ( .A(mul[21]), .B(n15), .Y(n16) );
  NAND2X1 U55 ( .A(n14), .B(n118), .Y(n17) );
  NAND2X2 U56 ( .A(n16), .B(n17), .Y(out[14]) );
  INVXL U57 ( .A(mul[21]), .Y(n14) );
  CLKINVX2 U58 ( .A(n118), .Y(n15) );
  AND2X2 U59 ( .A(n136), .B(n117), .Y(n115) );
  NAND2BX4 U60 ( .AN(mul[17]), .B(n111), .Y(n112) );
  XOR2X2 U61 ( .A(n115), .B(mul[19]), .Y(out[12]) );
  NOR2X4 U62 ( .A(in_17bit[1]), .B(in_17bit[0]), .Y(n32) );
  NOR2X4 U63 ( .A(n36), .B(n32), .Y(n28) );
  CLKINVX8 U64 ( .A(n109), .Y(n111) );
  NAND2BX4 U65 ( .AN(mul[16]), .B(n24), .Y(n109) );
  NAND2BX4 U66 ( .AN(mul[18]), .B(n114), .Y(n117) );
  XNOR2X4 U67 ( .A(n121), .B(n122), .Y(out[15]) );
  NOR2X2 U68 ( .A(n25), .B(n119), .Y(n118) );
  NOR3X2 U69 ( .A(mul[20]), .B(mul[19]), .C(n117), .Y(n119) );
  INVX2 U70 ( .A(in_8bit[3]), .Y(n47) );
  CLKINVX1 U71 ( .A(n105), .Y(n107) );
  XOR2X2 U72 ( .A(mul[17]), .B(n110), .Y(out[10]) );
  NAND2BXL U73 ( .AN(mul[14]), .B(n104), .Y(n105) );
  NOR2XL U74 ( .A(n25), .B(n92), .Y(n91) );
  INVX2 U75 ( .A(n39), .Y(n41) );
  XNOR2X1 U76 ( .A(in_17bit[16]), .B(n33), .Y(n25) );
  XNOR2XL U77 ( .A(n27), .B(in_8bit[6]), .Y(in_8bit_b[6]) );
  NAND2X1 U78 ( .A(n51), .B(n33), .Y(n27) );
  NAND2BXL U79 ( .AN(in_17bit[3]), .B(n56), .Y(n58) );
  INVX2 U80 ( .A(mul[22]), .Y(n122) );
  AOI21XL U81 ( .A0(n123), .A1(n122), .B0(n25), .Y(n124) );
  NOR2XL U82 ( .A(n25), .B(n95), .Y(n94) );
  NOR2XL U83 ( .A(n25), .B(n89), .Y(n88) );
  AOI22XL U84 ( .A0(mul[8]), .A1(n25), .B0(N33), .B1(n136), .Y(n135) );
  XOR2X1 U85 ( .A(mul[23]), .B(n124), .Y(out[16]) );
  NAND2XL U86 ( .A(n66), .B(in_17bit[16]), .Y(n65) );
  INVXL U87 ( .A(in_8bit[5]), .Y(n50) );
  NAND2XL U88 ( .A(n64), .B(n63), .Y(n66) );
  NAND2BXL U89 ( .AN(n58), .B(n59), .Y(n60) );
  NAND2BXL U90 ( .AN(n66), .B(n67), .Y(n68) );
  NAND2XL U91 ( .A(n74), .B(in_17bit[16]), .Y(n73) );
  NAND2XL U92 ( .A(n72), .B(n71), .Y(n74) );
  NAND2BXL U93 ( .AN(n74), .B(n75), .Y(n76) );
  NAND2XL U94 ( .A(n82), .B(in_17bit[16]), .Y(n81) );
  INVXL U95 ( .A(n86), .Y(sub_add_52_b0_carry[12]) );
  NAND2XL U96 ( .A(n80), .B(n79), .Y(n82) );
  AND2X1 U97 ( .A(N21), .B(in_17bit[16]), .Y(in_17bit_b[16]) );
  XOR2X2 U98 ( .A(n29), .B(in_17bit[3]), .Y(in_17bit_b[3]) );
  NOR2X2 U99 ( .A(n36), .B(n56), .Y(n29) );
  INVX1 U100 ( .A(n55), .Y(n56) );
  MX2X1 U101 ( .A(in_17bit[13]), .B(N18), .S0(in_17bit[16]), .Y(in_17bit_b[13]) );
  MX2X1 U102 ( .A(in_17bit[14]), .B(N19), .S0(in_17bit[16]), .Y(in_17bit_b[14]) );
  MX2X1 U103 ( .A(in_17bit[15]), .B(N20), .S0(in_17bit[16]), .Y(in_17bit_b[15]) );
  MX2X1 U104 ( .A(in_17bit[11]), .B(n30), .S0(in_17bit[16]), .Y(in_17bit_b[11]) );
  XNOR2X1 U105 ( .A(n84), .B(n127), .Y(n30) );
  MX2X1 U106 ( .A(in_17bit[12]), .B(n31), .S0(in_17bit[16]), .Y(in_17bit_b[12]) );
  XNOR2X1 U107 ( .A(n86), .B(n128), .Y(n31) );
  INVX1 U108 ( .A(n93), .Y(n95) );
  NAND2BX1 U109 ( .AN(mul[10]), .B(n92), .Y(n93) );
  INVX1 U110 ( .A(n87), .Y(n89) );
  NAND2BX1 U111 ( .AN(mul[8]), .B(n126), .Y(n87) );
  INVX1 U112 ( .A(n90), .Y(n92) );
  NAND2BX1 U113 ( .AN(mul[9]), .B(n89), .Y(n90) );
  XOR2X1 U114 ( .A(mul[16]), .B(n108), .Y(out[9]) );
  NOR2X1 U115 ( .A(n25), .B(n24), .Y(n108) );
  XOR2X1 U116 ( .A(mul[13]), .B(n100), .Y(out[6]) );
  NOR2X1 U117 ( .A(n25), .B(n101), .Y(n100) );
  XOR2X1 U118 ( .A(mul[15]), .B(n106), .Y(out[8]) );
  NOR2X1 U119 ( .A(n25), .B(n107), .Y(n106) );
  XOR2X1 U120 ( .A(mul[14]), .B(n103), .Y(out[7]) );
  NOR2X1 U121 ( .A(n25), .B(n104), .Y(n103) );
  XOR2X1 U122 ( .A(mul[12]), .B(n97), .Y(out[5]) );
  NOR2X1 U123 ( .A(n25), .B(n98), .Y(n97) );
  XOR2X1 U124 ( .A(mul[11]), .B(n94), .Y(out[4]) );
  XOR2X1 U125 ( .A(mul[9]), .B(n88), .Y(out[2]) );
  XOR2X1 U126 ( .A(mul[10]), .B(n91), .Y(out[3]) );
  INVX1 U127 ( .A(n99), .Y(n101) );
  INVX1 U128 ( .A(n102), .Y(n104) );
  NAND2BX1 U129 ( .AN(mul[13]), .B(n101), .Y(n102) );
  INVX1 U130 ( .A(n96), .Y(n98) );
  NAND2BX1 U131 ( .AN(mul[11]), .B(n95), .Y(n96) );
  INVX1 U132 ( .A(n135), .Y(out[1]) );
  INVX1 U133 ( .A(n134), .Y(out[0]) );
  AOI22XL U134 ( .A0(N32), .A1(n25), .B0(N32), .B1(n136), .Y(n134) );
  XOR2X1 U135 ( .A(n35), .B(n37), .Y(in_8bit_b[1]) );
  NAND2XL U136 ( .A(in_8bit[0]), .B(n33), .Y(n37) );
  INVX1 U137 ( .A(n133), .Y(in_8bit_b[0]) );
  AOI22XL U138 ( .A0(in_8bit[0]), .A1(n33), .B0(in_8bit[0]), .B1(n34), .Y(n133) );
  XNOR2X1 U139 ( .A(n69), .B(n71), .Y(in_17bit_b[7]) );
  NOR2X1 U140 ( .A(n36), .B(n72), .Y(n69) );
  XNOR2X1 U141 ( .A(n78), .B(n79), .Y(in_17bit_b[9]) );
  NOR2X1 U142 ( .A(n36), .B(n80), .Y(n78) );
  XOR2X1 U143 ( .A(n59), .B(n57), .Y(in_17bit_b[4]) );
  NAND2X1 U144 ( .A(n58), .B(in_17bit[16]), .Y(n57) );
  XOR2X1 U145 ( .A(n67), .B(n65), .Y(in_17bit_b[6]) );
  XOR2X1 U146 ( .A(n75), .B(n73), .Y(in_17bit_b[8]) );
  INVX1 U147 ( .A(n60), .Y(n64) );
  INVX1 U148 ( .A(n68), .Y(n72) );
  INVX1 U149 ( .A(n76), .Y(n80) );
  INVX1 U150 ( .A(in_8bit[7]), .Y(n34) );
  XOR2X1 U151 ( .A(n83), .B(n81), .Y(in_17bit_b[10]) );
  NAND2BX1 U152 ( .AN(n82), .B(n83), .Y(n84) );
  NAND2X1 U153 ( .A(n127), .B(n85), .Y(n86) );
  INVX1 U154 ( .A(n84), .Y(n85) );
  INVX1 U155 ( .A(in_17bit[5]), .Y(n63) );
  INVX1 U156 ( .A(in_17bit[4]), .Y(n59) );
  INVX1 U157 ( .A(in_17bit[7]), .Y(n71) );
  INVX1 U158 ( .A(in_17bit[6]), .Y(n67) );
  INVX1 U159 ( .A(in_17bit[8]), .Y(n75) );
  INVX1 U160 ( .A(in_17bit[9]), .Y(n79) );
  INVX1 U161 ( .A(in_17bit[10]), .Y(n83) );
  INVX1 U162 ( .A(in_17bit[11]), .Y(n127) );
  INVX1 U163 ( .A(in_17bit[12]), .Y(n128) );
  INVX1 U164 ( .A(in_17bit[13]), .Y(n129) );
  INVX1 U165 ( .A(in_17bit[14]), .Y(n130) );
  INVX1 U166 ( .A(in_17bit[15]), .Y(n131) );
  AOI21X1 U167 ( .A0(n45), .A1(n44), .B0(n34), .Y(n46) );
  NOR3XL U168 ( .A(in_8bit[0]), .B(in_8bit[3]), .C(in_8bit[1]), .Y(n44) );
  NOR2X1 U169 ( .A(in_8bit[4]), .B(in_8bit[2]), .Y(n45) );
  NOR2XL U170 ( .A(in_8bit[3]), .B(in_8bit[2]), .Y(n42) );
  NOR2X4 U171 ( .A(n25), .B(n111), .Y(n110) );
  NOR2X4 U172 ( .A(n25), .B(n114), .Y(n113) );
  XOR2X4 U173 ( .A(n18), .B(n113), .Y(out[11]) );
  XOR2X1 U174 ( .A(n125), .B(n126), .Y(N33) );
  XOR2X1 U175 ( .A(n36), .B(sub_add_52_b0_carry[16]), .Y(N21) );
  AND2X1 U176 ( .A(sub_add_52_b0_carry[15]), .B(n131), .Y(
        sub_add_52_b0_carry[16]) );
  XOR2X1 U177 ( .A(n131), .B(sub_add_52_b0_carry[15]), .Y(N20) );
  AND2X1 U178 ( .A(sub_add_52_b0_carry[14]), .B(n130), .Y(
        sub_add_52_b0_carry[15]) );
  XOR2X1 U179 ( .A(n130), .B(sub_add_52_b0_carry[14]), .Y(N19) );
  AND2X1 U180 ( .A(sub_add_52_b0_carry[13]), .B(n129), .Y(
        sub_add_52_b0_carry[14]) );
  XOR2X1 U181 ( .A(n129), .B(sub_add_52_b0_carry[13]), .Y(N18) );
  AND2X1 U182 ( .A(sub_add_52_b0_carry[12]), .B(n128), .Y(
        sub_add_52_b0_carry[13]) );
endmodule


module multi16_9_DW01_add_0 ( A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, 
        A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, 
        B_20_, B_19_, B_18_, B_17_, B_16_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, 
        SUM_17_, SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, 
        SUM_9_, SUM_8_, SUM_7_, SUM_6_, SUM_5_ );
  input A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_,
         A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, B_20_, B_19_,
         B_18_, B_17_, B_16_;
  output SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, SUM_15_,
         SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, SUM_7_,
         SUM_6_, SUM_5_;
  wire   n1, n2, n3, n4, n5, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41;

  INVX4 U2 ( .A(n35), .Y(n19) );
  NAND2X2 U3 ( .A(n1), .B(n2), .Y(n3) );
  NAND2X2 U4 ( .A(n3), .B(n33), .Y(n36) );
  INVX2 U5 ( .A(n38), .Y(n1) );
  INVXL U6 ( .A(n31), .Y(n2) );
  INVX2 U7 ( .A(n41), .Y(SUM_16_) );
  NAND2X2 U8 ( .A(n34), .B(n40), .Y(n41) );
  XOR2X2 U9 ( .A(n4), .B(n38), .Y(SUM_18_) );
  AOI2BB1X4 U10 ( .A0N(n34), .A1N(n30), .B0(n19), .Y(n38) );
  XOR2X2 U11 ( .A(n36), .B(n37), .Y(SUM_19_) );
  OR2X2 U12 ( .A(B_16_), .B(A_16_), .Y(n40) );
  BUFX3 U13 ( .A(A_13_), .Y(SUM_13_) );
  BUFX3 U14 ( .A(A_14_), .Y(SUM_14_) );
  NAND2X1 U15 ( .A(n33), .B(n17), .Y(n4) );
  NOR2X1 U16 ( .A(B_18_), .B(A_18_), .Y(n31) );
  NOR2BX1 U17 ( .AN(n29), .B(n28), .Y(n37) );
  INVX1 U18 ( .A(n31), .Y(n17) );
  INVX1 U19 ( .A(n34), .Y(n20) );
  NAND2X2 U20 ( .A(B_16_), .B(A_16_), .Y(n34) );
  INVX4 U21 ( .A(n21), .Y(SUM_15_) );
  OAI21X1 U22 ( .A0(n27), .A1(n28), .B0(n29), .Y(n24) );
  AOI21XL U23 ( .A0(n17), .A1(n32), .B0(n18), .Y(n27) );
  NOR2X4 U24 ( .A(B_17_), .B(A_17_), .Y(n30) );
  NAND2X2 U25 ( .A(B_17_), .B(A_17_), .Y(n35) );
  NAND2X2 U26 ( .A(B_19_), .B(A_19_), .Y(n29) );
  NOR2X1 U27 ( .A(B_19_), .B(A_19_), .Y(n28) );
  INVXL U28 ( .A(n26), .Y(n16) );
  NAND2X1 U29 ( .A(n26), .B(n25), .Y(n5) );
  NOR2X4 U30 ( .A(n30), .B(n19), .Y(n39) );
  XNOR2X1 U31 ( .A(n5), .B(n24), .Y(SUM_20_) );
  BUFX4 U32 ( .A(A_12_), .Y(SUM_12_) );
  BUFX3 U33 ( .A(A_11_), .Y(SUM_11_) );
  INVXL U34 ( .A(n33), .Y(n18) );
  INVX2 U35 ( .A(A_15_), .Y(n21) );
  BUFX3 U36 ( .A(A_6_), .Y(SUM_6_) );
  BUFX3 U37 ( .A(A_7_), .Y(SUM_7_) );
  BUFX3 U38 ( .A(A_8_), .Y(SUM_8_) );
  BUFX3 U39 ( .A(A_9_), .Y(SUM_9_) );
  BUFX3 U40 ( .A(A_10_), .Y(SUM_10_) );
  BUFX3 U41 ( .A(A_5_), .Y(SUM_5_) );
  XOR2X2 U42 ( .A(n20), .B(n39), .Y(SUM_17_) );
  XOR2X1 U43 ( .A(n22), .B(n23), .Y(SUM_21_) );
  AOI21X1 U44 ( .A0(n24), .A1(n25), .B0(n16), .Y(n23) );
  XNOR2X1 U45 ( .A(B_21_), .B(A_21_), .Y(n22) );
  OAI21XL U46 ( .A0(n30), .A1(n34), .B0(n35), .Y(n32) );
  OR2X1 U47 ( .A(B_20_), .B(A_20_), .Y(n25) );
  NAND2X1 U48 ( .A(B_20_), .B(A_20_), .Y(n26) );
  NAND2X1 U49 ( .A(B_18_), .B(A_18_), .Y(n33) );
endmodule


module multi16_9_DW02_mult_0 ( A, B, PRODUCT_23_, PRODUCT_22_, PRODUCT_21_, 
        PRODUCT_20_, PRODUCT_19_, PRODUCT_18_, PRODUCT_17_, PRODUCT_16_, 
        PRODUCT_15_, PRODUCT_14_, PRODUCT_13_, PRODUCT_12_, PRODUCT_11_, 
        PRODUCT_10_, PRODUCT_9_, PRODUCT_8_, PRODUCT_7_ );
  input [16:0] A;
  input [7:0] B;
  output PRODUCT_23_, PRODUCT_22_, PRODUCT_21_, PRODUCT_20_, PRODUCT_19_,
         PRODUCT_18_, PRODUCT_17_, PRODUCT_16_, PRODUCT_15_, PRODUCT_14_,
         PRODUCT_13_, PRODUCT_12_, PRODUCT_11_, PRODUCT_10_, PRODUCT_9_,
         PRODUCT_8_, PRODUCT_7_;
  wire   ab_16__7_, ab_16__6_, ab_16__5_, ab_16__4_, ab_16__3_, ab_16__2_,
         ab_16__1_, ab_16__0_, ab_15__7_, ab_15__6_, ab_15__5_, ab_15__4_,
         ab_15__3_, ab_15__2_, ab_15__1_, ab_15__0_, ab_14__7_, ab_14__6_,
         ab_14__5_, ab_14__4_, ab_14__3_, ab_14__2_, ab_14__1_, ab_14__0_,
         ab_13__7_, ab_13__6_, ab_13__5_, ab_13__4_, ab_13__3_, ab_13__2_,
         ab_13__1_, ab_13__0_, ab_12__7_, ab_12__6_, ab_12__5_, ab_12__4_,
         ab_12__3_, ab_12__2_, ab_12__1_, ab_12__0_, ab_11__7_, ab_11__6_,
         ab_11__5_, ab_11__4_, ab_11__3_, ab_11__2_, ab_11__1_, ab_11__0_,
         ab_10__7_, ab_10__6_, ab_10__5_, ab_10__4_, ab_10__3_, ab_10__2_,
         ab_10__1_, ab_10__0_, ab_9__7_, ab_9__6_, ab_9__5_, ab_9__4_,
         ab_9__3_, ab_9__2_, ab_9__1_, ab_9__0_, ab_8__7_, ab_8__6_, ab_8__5_,
         ab_8__4_, ab_8__3_, ab_8__2_, ab_8__1_, ab_8__0_, ab_7__7_, ab_7__6_,
         ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_, ab_7__0_, ab_6__7_,
         ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_, ab_6__1_, ab_6__0_,
         ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_, ab_5__2_, ab_5__1_,
         ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_, ab_4__3_, ab_4__2_,
         ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_, ab_3__4_, ab_3__3_,
         ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_, ab_2__5_, ab_2__4_,
         ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_, ab_1__6_, ab_1__5_,
         ab_1__4_, ab_1__3_, ab_1__2_, ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_,
         ab_0__3_, ab_0__2_, CARRYB_16__6_, CARRYB_16__5_, CARRYB_16__4_,
         CARRYB_16__3_, CARRYB_16__2_, CARRYB_16__1_, CARRYB_16__0_,
         CARRYB_15__6_, CARRYB_15__5_, CARRYB_15__4_, CARRYB_15__3_,
         CARRYB_15__2_, CARRYB_15__1_, CARRYB_15__0_, CARRYB_14__6_,
         CARRYB_14__5_, CARRYB_14__4_, CARRYB_14__3_, CARRYB_14__2_,
         CARRYB_14__1_, CARRYB_14__0_, CARRYB_13__6_, CARRYB_13__5_,
         CARRYB_13__4_, CARRYB_13__3_, CARRYB_13__2_, CARRYB_13__1_,
         CARRYB_13__0_, CARRYB_12__6_, CARRYB_12__5_, CARRYB_12__4_,
         CARRYB_12__3_, CARRYB_12__2_, CARRYB_12__1_, CARRYB_12__0_,
         CARRYB_11__6_, CARRYB_11__5_, CARRYB_11__4_, CARRYB_11__3_,
         CARRYB_11__2_, CARRYB_11__1_, CARRYB_11__0_, CARRYB_10__6_,
         CARRYB_10__5_, CARRYB_10__4_, CARRYB_10__3_, CARRYB_10__2_,
         CARRYB_10__1_, CARRYB_10__0_, CARRYB_9__6_, CARRYB_9__5_,
         CARRYB_9__4_, CARRYB_9__3_, CARRYB_9__2_, CARRYB_9__1_, CARRYB_9__0_,
         CARRYB_8__6_, CARRYB_8__5_, CARRYB_8__4_, CARRYB_8__3_, CARRYB_8__2_,
         CARRYB_8__1_, CARRYB_8__0_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_,
         CARRYB_7__3_, CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_,
         CARRYB_6__5_, CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_,
         CARRYB_6__0_, CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_,
         CARRYB_5__2_, CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_,
         CARRYB_4__4_, CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_,
         CARRYB_3__6_, CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_,
         CARRYB_3__1_, CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_,
         CARRYB_2__3_, CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__0_,
         SUMB_16__6_, SUMB_16__5_, SUMB_16__4_, SUMB_16__3_, SUMB_16__2_,
         SUMB_16__1_, SUMB_16__0_, SUMB_15__6_, SUMB_15__5_, SUMB_15__4_,
         SUMB_15__3_, SUMB_15__2_, SUMB_15__1_, SUMB_14__6_, SUMB_14__5_,
         SUMB_14__4_, SUMB_14__3_, SUMB_14__2_, SUMB_14__1_, SUMB_13__6_,
         SUMB_13__5_, SUMB_13__4_, SUMB_13__3_, SUMB_13__2_, SUMB_13__1_,
         SUMB_12__6_, SUMB_12__5_, SUMB_12__4_, SUMB_12__3_, SUMB_12__2_,
         SUMB_12__1_, SUMB_11__6_, SUMB_11__5_, SUMB_11__4_, SUMB_11__3_,
         SUMB_11__2_, SUMB_11__1_, SUMB_10__6_, SUMB_10__5_, SUMB_10__4_,
         SUMB_10__3_, SUMB_10__2_, SUMB_10__1_, SUMB_9__6_, SUMB_9__5_,
         SUMB_9__4_, SUMB_9__3_, SUMB_9__2_, SUMB_9__1_, SUMB_8__6_,
         SUMB_8__5_, SUMB_8__4_, SUMB_8__3_, SUMB_8__2_, SUMB_8__1_,
         SUMB_7__6_, SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_,
         SUMB_7__1_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, PROD1_7_, A1_21_, A1_20_, A1_19_, A1_18_,
         A1_17_, A1_16_, A1_15_, A1_13_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_,
         A1_7_, A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, n3, n4, n5, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37;

  ADDFHX4 S1_14_0 ( .A(ab_14__0_), .B(CARRYB_13__0_), .CI(SUMB_13__1_), .CO(
        CARRYB_14__0_), .S(A1_12_) );
  ADDFHX4 S2_14_3 ( .A(ab_14__3_), .B(CARRYB_13__3_), .CI(SUMB_13__4_), .CO(
        CARRYB_14__3_), .S(SUMB_14__3_) );
  ADDFHX4 S1_13_0 ( .A(ab_13__0_), .B(CARRYB_12__0_), .CI(SUMB_12__1_), .CO(
        CARRYB_13__0_), .S(A1_11_) );
  ADDFHX4 S2_13_1 ( .A(ab_13__1_), .B(CARRYB_12__1_), .CI(SUMB_12__2_), .CO(
        CARRYB_13__1_), .S(SUMB_13__1_) );
  ADDFHX4 S2_12_3 ( .A(ab_12__3_), .B(CARRYB_11__3_), .CI(SUMB_11__4_), .CO(
        CARRYB_12__3_), .S(SUMB_12__3_) );
  ADDFHX4 S1_11_0 ( .A(ab_11__0_), .B(CARRYB_10__0_), .CI(SUMB_10__1_), .CO(
        CARRYB_11__0_), .S(A1_9_) );
  ADDFHX4 S2_11_3 ( .A(ab_11__3_), .B(CARRYB_10__3_), .CI(SUMB_10__4_), .CO(
        CARRYB_11__3_), .S(SUMB_11__3_) );
  ADDFHX4 S1_10_0 ( .A(ab_10__0_), .B(CARRYB_9__0_), .CI(SUMB_9__1_), .CO(
        CARRYB_10__0_), .S(A1_8_) );
  ADDFHX4 S2_10_1 ( .A(ab_10__1_), .B(CARRYB_9__1_), .CI(SUMB_9__2_), .CO(
        CARRYB_10__1_), .S(SUMB_10__1_) );
  ADDFHX4 S2_10_2 ( .A(ab_10__2_), .B(CARRYB_9__2_), .CI(SUMB_9__3_), .CO(
        CARRYB_10__2_), .S(SUMB_10__2_) );
  ADDFHX4 S2_10_3 ( .A(ab_10__3_), .B(CARRYB_9__3_), .CI(SUMB_9__4_), .CO(
        CARRYB_10__3_), .S(SUMB_10__3_) );
  ADDFHX4 S2_10_5 ( .A(ab_10__5_), .B(CARRYB_9__5_), .CI(SUMB_9__6_), .CO(
        CARRYB_10__5_), .S(SUMB_10__5_) );
  ADDFHX4 S2_9_1 ( .A(ab_9__1_), .B(CARRYB_8__1_), .CI(SUMB_8__2_), .CO(
        CARRYB_9__1_), .S(SUMB_9__1_) );
  ADDFHX4 S2_9_5 ( .A(ab_9__5_), .B(CARRYB_8__5_), .CI(SUMB_8__6_), .CO(
        CARRYB_9__5_), .S(SUMB_9__5_) );
  ADDFHX4 S1_8_0 ( .A(ab_8__0_), .B(CARRYB_7__0_), .CI(SUMB_7__1_), .CO(
        CARRYB_8__0_), .S(A1_6_) );
  ADDFHX4 S2_8_1 ( .A(ab_8__1_), .B(CARRYB_7__1_), .CI(SUMB_7__2_), .CO(
        CARRYB_8__1_), .S(SUMB_8__1_) );
  ADDFHX4 S2_8_2 ( .A(ab_8__2_), .B(CARRYB_7__2_), .CI(SUMB_7__3_), .CO(
        CARRYB_8__2_), .S(SUMB_8__2_) );
  ADDFHX4 S2_8_3 ( .A(ab_8__3_), .B(CARRYB_7__3_), .CI(SUMB_7__4_), .CO(
        CARRYB_8__3_), .S(SUMB_8__3_) );
  ADDFHX4 S2_7_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  ADDFHX4 S2_7_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  ADDFHX4 S2_7_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  ADDFHX4 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  ADDFHX4 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  ADDFHX4 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  ADDFHX4 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  ADDFHX4 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  ADDFHX4 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  ADDFHX4 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  ADDFHX4 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  ADDFHX4 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  ADDFHX4 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  ADDFHX4 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  multi16_9_DW01_add_0 FS_1 ( .A_21_(A1_21_), .A_20_(A1_20_), .A_19_(A1_19_), 
        .A_18_(A1_18_), .A_17_(A1_17_), .A_16_(A1_16_), .A_15_(A1_15_), 
        .A_14_(SUMB_16__0_), .A_13_(A1_13_), .A_12_(A1_12_), .A_11_(A1_11_), 
        .A_10_(A1_10_), .A_9_(A1_9_), .A_8_(A1_8_), .A_7_(A1_7_), .A_6_(A1_6_), 
        .A_5_(PROD1_7_), .B_21_(n18), .B_20_(n17), .B_19_(n16), .B_18_(n15), 
        .B_17_(n14), .B_16_(n13), .SUM_21_(PRODUCT_23_), .SUM_20_(PRODUCT_22_), 
        .SUM_19_(PRODUCT_21_), .SUM_18_(PRODUCT_20_), .SUM_17_(PRODUCT_19_), 
        .SUM_16_(PRODUCT_18_), .SUM_15_(PRODUCT_17_), .SUM_14_(PRODUCT_16_), 
        .SUM_13_(PRODUCT_15_), .SUM_12_(PRODUCT_14_), .SUM_11_(PRODUCT_13_), 
        .SUM_10_(PRODUCT_12_), .SUM_9_(PRODUCT_11_), .SUM_8_(PRODUCT_10_), 
        .SUM_7_(PRODUCT_9_), .SUM_6_(PRODUCT_8_), .SUM_5_(PRODUCT_7_) );
  ADDFHX2 S2_8_5 ( .A(ab_8__5_), .B(CARRYB_7__5_), .CI(SUMB_7__6_), .CO(
        CARRYB_8__5_), .S(SUMB_8__5_) );
  ADDFHX1 S3_15_6 ( .A(ab_15__6_), .B(CARRYB_14__6_), .CI(ab_14__7_), .CO(
        CARRYB_15__6_), .S(SUMB_15__6_) );
  ADDFHX2 S2_15_4 ( .A(ab_15__4_), .B(CARRYB_14__4_), .CI(SUMB_14__5_), .CO(
        CARRYB_15__4_), .S(SUMB_15__4_) );
  ADDFHX2 S2_15_5 ( .A(ab_15__5_), .B(CARRYB_14__5_), .CI(SUMB_14__6_), .CO(
        CARRYB_15__5_), .S(SUMB_15__5_) );
  ADDFX2 S5_6 ( .A(ab_16__6_), .B(CARRYB_15__6_), .CI(ab_15__7_), .CO(
        CARRYB_16__6_), .S(SUMB_16__6_) );
  ADDFHX4 S2_11_2 ( .A(ab_11__2_), .B(CARRYB_10__2_), .CI(SUMB_10__3_), .CO(
        CARRYB_11__2_), .S(SUMB_11__2_) );
  ADDFHX2 S3_2_6 ( .A(ab_2__6_), .B(n11), .CI(ab_1__7_), .CO(CARRYB_2__6_), 
        .S(SUMB_2__6_) );
  ADDFHX4 S3_9_6 ( .A(ab_9__6_), .B(CARRYB_8__6_), .CI(ab_8__7_), .CO(
        CARRYB_9__6_), .S(SUMB_9__6_) );
  ADDFHX4 S2_12_2 ( .A(ab_12__2_), .B(CARRYB_11__2_), .CI(SUMB_11__3_), .CO(
        CARRYB_12__2_), .S(SUMB_12__2_) );
  ADDFHX4 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  ADDFHX4 S2_7_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  ADDFHX2 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  ADDFHX4 S2_14_2 ( .A(ab_14__2_), .B(CARRYB_13__2_), .CI(SUMB_13__3_), .CO(
        CARRYB_14__2_), .S(SUMB_14__2_) );
  ADDFHX4 S3_7_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(
        CARRYB_7__6_), .S(SUMB_7__6_) );
  ADDFHX2 S3_12_6 ( .A(ab_12__6_), .B(CARRYB_11__6_), .CI(ab_11__7_), .CO(
        CARRYB_12__6_), .S(SUMB_12__6_) );
  ADDFHX4 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  ADDFHX2 S2_14_5 ( .A(ab_14__5_), .B(CARRYB_13__5_), .CI(SUMB_13__6_), .CO(
        CARRYB_14__5_), .S(SUMB_14__5_) );
  ADDFHX4 S2_10_4 ( .A(ab_10__4_), .B(CARRYB_9__4_), .CI(SUMB_9__5_), .CO(
        CARRYB_10__4_), .S(SUMB_10__4_) );
  ADDFHX4 S2_11_4 ( .A(ab_11__4_), .B(CARRYB_10__4_), .CI(SUMB_10__5_), .CO(
        CARRYB_11__4_), .S(SUMB_11__4_) );
  ADDFHX2 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  ADDFHX4 S2_14_1 ( .A(ab_14__1_), .B(CARRYB_13__1_), .CI(SUMB_13__2_), .CO(
        CARRYB_14__1_), .S(SUMB_14__1_) );
  ADDFHX4 S3_10_6 ( .A(ab_10__6_), .B(CARRYB_9__6_), .CI(ab_9__7_), .CO(
        CARRYB_10__6_), .S(SUMB_10__6_) );
  ADDFHX2 S2_2_5 ( .A(ab_2__5_), .B(n9), .CI(SUMB_1__6_), .CO(CARRYB_2__5_), 
        .S(SUMB_2__5_) );
  ADDFHX4 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  ADDFHX4 S2_11_1 ( .A(ab_11__1_), .B(CARRYB_10__1_), .CI(SUMB_10__2_), .CO(
        CARRYB_11__1_), .S(SUMB_11__1_) );
  ADDFHX4 S2_15_1 ( .A(ab_15__1_), .B(CARRYB_14__1_), .CI(SUMB_14__2_), .CO(
        CARRYB_15__1_), .S(SUMB_15__1_) );
  ADDFHX4 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  ADDFHX4 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  ADDFHX4 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  ADDFHX1 S3_14_6 ( .A(ab_14__6_), .B(CARRYB_13__6_), .CI(ab_13__7_), .CO(
        CARRYB_14__6_), .S(SUMB_14__6_) );
  ADDFHX1 S4_5 ( .A(ab_16__5_), .B(CARRYB_15__5_), .CI(SUMB_15__6_), .CO(
        CARRYB_16__5_), .S(SUMB_16__5_) );
  ADDFHX2 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  ADDFHX2 S1_7_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(PROD1_7_) );
  ADDFHX2 S3_11_6 ( .A(ab_11__6_), .B(CARRYB_10__6_), .CI(ab_10__7_), .CO(
        CARRYB_11__6_), .S(SUMB_11__6_) );
  ADDFHX2 S4_4 ( .A(ab_16__4_), .B(CARRYB_15__4_), .CI(SUMB_15__5_), .CO(
        CARRYB_16__4_), .S(SUMB_16__4_) );
  ADDFHX2 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  ADDFHX2 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  ADDFHX2 S4_1 ( .A(ab_16__1_), .B(CARRYB_15__1_), .CI(SUMB_15__2_), .CO(
        CARRYB_16__1_), .S(SUMB_16__1_) );
  ADDFHX1 S4_0 ( .A(ab_16__0_), .B(CARRYB_15__0_), .CI(SUMB_15__1_), .CO(
        CARRYB_16__0_), .S(SUMB_16__0_) );
  ADDFHX2 S2_2_2 ( .A(ab_2__2_), .B(n10), .CI(SUMB_1__3_), .CO(CARRYB_2__2_), 
        .S(SUMB_2__2_) );
  ADDFHX2 S1_9_0 ( .A(ab_9__0_), .B(CARRYB_8__0_), .CI(SUMB_8__1_), .CO(
        CARRYB_9__0_), .S(A1_7_) );
  ADDFHX2 S1_12_0 ( .A(ab_12__0_), .B(CARRYB_11__0_), .CI(SUMB_11__1_), .CO(
        CARRYB_12__0_), .S(A1_10_) );
  ADDFHX2 S3_8_6 ( .A(ab_8__6_), .B(CARRYB_7__6_), .CI(ab_7__7_), .CO(
        CARRYB_8__6_), .S(SUMB_8__6_) );
  ADDFHX2 S2_12_1 ( .A(ab_12__1_), .B(CARRYB_11__1_), .CI(SUMB_11__2_), .CO(
        CARRYB_12__1_), .S(SUMB_12__1_) );
  ADDFHX2 S2_9_2 ( .A(ab_9__2_), .B(CARRYB_8__2_), .CI(SUMB_8__3_), .CO(
        CARRYB_9__2_), .S(SUMB_9__2_) );
  ADDFHX2 S2_13_2 ( .A(ab_13__2_), .B(CARRYB_12__2_), .CI(SUMB_12__3_), .CO(
        CARRYB_13__2_), .S(SUMB_13__2_) );
  ADDFHX2 S2_13_3 ( .A(ab_13__3_), .B(CARRYB_12__3_), .CI(SUMB_12__4_), .CO(
        CARRYB_13__3_), .S(SUMB_13__3_) );
  ADDFHX2 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  ADDFHX2 S2_2_1 ( .A(ab_2__1_), .B(n12), .CI(SUMB_1__2_), .CO(CARRYB_2__1_), 
        .S(SUMB_2__1_) );
  ADDFHX2 S1_15_0 ( .A(ab_15__0_), .B(CARRYB_14__0_), .CI(SUMB_14__1_), .CO(
        CARRYB_15__0_), .S(A1_13_) );
  ADDFHX2 S3_13_6 ( .A(ab_13__6_), .B(CARRYB_12__6_), .CI(ab_12__7_), .CO(
        CARRYB_13__6_), .S(SUMB_13__6_) );
  ADDFHX4 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  ADDFHX2 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  ADDFHX4 S2_15_2 ( .A(ab_15__2_), .B(CARRYB_14__2_), .CI(SUMB_14__3_), .CO(
        CARRYB_15__2_), .S(SUMB_15__2_) );
  ADDFHX2 S4_2 ( .A(ab_16__2_), .B(CARRYB_15__2_), .CI(SUMB_15__3_), .CO(
        CARRYB_16__2_), .S(SUMB_16__2_) );
  ADDFHX4 S4_3 ( .A(ab_16__3_), .B(CARRYB_15__3_), .CI(SUMB_15__4_), .CO(
        CARRYB_16__3_), .S(SUMB_16__3_) );
  ADDFHX4 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  ADDFHX4 S2_9_4 ( .A(ab_9__4_), .B(CARRYB_8__4_), .CI(SUMB_8__5_), .CO(
        CARRYB_9__4_), .S(SUMB_9__4_) );
  ADDFHX4 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  ADDFHX4 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  ADDFHX4 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  ADDFHX4 S2_11_5 ( .A(ab_11__5_), .B(CARRYB_10__5_), .CI(SUMB_10__6_), .CO(
        CARRYB_11__5_), .S(SUMB_11__5_) );
  ADDFHX4 S2_13_5 ( .A(ab_13__5_), .B(CARRYB_12__5_), .CI(SUMB_12__6_), .CO(
        CARRYB_13__5_), .S(SUMB_13__5_) );
  ADDFHX4 S2_2_3 ( .A(ab_2__3_), .B(n7), .CI(SUMB_1__4_), .CO(CARRYB_2__3_), 
        .S(SUMB_2__3_) );
  ADDFHX2 S2_8_4 ( .A(ab_8__4_), .B(CARRYB_7__4_), .CI(SUMB_7__5_), .CO(
        CARRYB_8__4_), .S(SUMB_8__4_) );
  ADDFHX4 S2_9_3 ( .A(ab_9__3_), .B(CARRYB_8__3_), .CI(SUMB_8__4_), .CO(
        CARRYB_9__3_), .S(SUMB_9__3_) );
  ADDFHX4 S2_14_4 ( .A(ab_14__4_), .B(CARRYB_13__4_), .CI(SUMB_13__5_), .CO(
        CARRYB_14__4_), .S(SUMB_14__4_) );
  ADDFHX4 S2_2_4 ( .A(ab_2__4_), .B(n8), .CI(SUMB_1__5_), .CO(CARRYB_2__4_), 
        .S(SUMB_2__4_) );
  ADDFHX2 S2_12_4 ( .A(ab_12__4_), .B(CARRYB_11__4_), .CI(SUMB_11__5_), .CO(
        CARRYB_12__4_), .S(SUMB_12__4_) );
  ADDFHX2 S2_12_5 ( .A(ab_12__5_), .B(CARRYB_11__5_), .CI(SUMB_11__6_), .CO(
        CARRYB_12__5_), .S(SUMB_12__5_) );
  ADDFHX4 S2_13_4 ( .A(ab_13__4_), .B(CARRYB_12__4_), .CI(SUMB_12__5_), .CO(
        CARRYB_13__4_), .S(SUMB_13__4_) );
  ADDFHX2 S2_15_3 ( .A(ab_15__3_), .B(CARRYB_14__3_), .CI(SUMB_14__4_), .CO(
        CARRYB_15__3_), .S(SUMB_15__3_) );
  AND2X2 U2 ( .A(A[2]), .B(B[3]), .Y(ab_2__3_) );
  AND2X2 U3 ( .A(A[3]), .B(B[0]), .Y(ab_3__0_) );
  XOR3X4 U4 ( .A(CARRYB_6__2_), .B(ab_7__2_), .C(SUMB_6__3_), .Y(SUMB_7__2_)
         );
  NAND2X1 U5 ( .A(SUMB_6__3_), .B(CARRYB_6__2_), .Y(n3) );
  NAND2X1 U6 ( .A(ab_7__2_), .B(CARRYB_6__2_), .Y(n4) );
  NAND2X1 U7 ( .A(ab_7__2_), .B(SUMB_6__3_), .Y(n5) );
  NAND3X2 U8 ( .A(n5), .B(n3), .C(n4), .Y(CARRYB_7__2_) );
  AND2X2 U9 ( .A(A[7]), .B(B[2]), .Y(ab_7__2_) );
  AND2X2 U10 ( .A(A[1]), .B(B[5]), .Y(ab_1__5_) );
  NOR2X2 U11 ( .A(n27), .B(n21), .Y(ab_0__3_) );
  INVX2 U12 ( .A(A[0]), .Y(n21) );
  NOR2X1 U13 ( .A(n28), .B(n21), .Y(ab_0__2_) );
  AND2X2 U14 ( .A(A[1]), .B(B[2]), .Y(ab_1__2_) );
  CLKINVX3 U15 ( .A(B[3]), .Y(n27) );
  INVX2 U16 ( .A(B[2]), .Y(n28) );
  XOR2X1 U17 ( .A(ab_1__2_), .B(ab_0__3_), .Y(SUMB_1__2_) );
  XOR2X1 U18 ( .A(CARRYB_16__3_), .B(SUMB_16__4_), .Y(A1_18_) );
  BUFX3 U19 ( .A(B[7]), .Y(n19) );
  XOR2X2 U20 ( .A(CARRYB_16__1_), .B(SUMB_16__2_), .Y(A1_16_) );
  CLKINVX3 U21 ( .A(B[6]), .Y(n24) );
  AND2X2 U23 ( .A(ab_0__4_), .B(ab_1__3_), .Y(n7) );
  AND2X2 U24 ( .A(ab_0__5_), .B(ab_1__4_), .Y(n8) );
  AND2X2 U25 ( .A(ab_0__6_), .B(ab_1__5_), .Y(n9) );
  AND2X2 U26 ( .A(ab_0__3_), .B(ab_1__2_), .Y(n10) );
  AND2X2 U27 ( .A(ab_0__7_), .B(ab_1__6_), .Y(n11) );
  AND2X2 U28 ( .A(ab_0__2_), .B(n31), .Y(n12) );
  NOR2X2 U29 ( .A(n26), .B(n21), .Y(ab_0__4_) );
  NOR2X2 U30 ( .A(n24), .B(n21), .Y(ab_0__6_) );
  AND2X2 U31 ( .A(A[2]), .B(B[1]), .Y(ab_2__1_) );
  NOR2X1 U32 ( .A(n30), .B(n21), .Y(ab_0__7_) );
  INVX2 U33 ( .A(n19), .Y(n30) );
  XOR2X1 U34 ( .A(ab_1__6_), .B(ab_0__7_), .Y(SUMB_1__6_) );
  AND2X2 U35 ( .A(CARRYB_16__0_), .B(SUMB_16__1_), .Y(n13) );
  AND2X1 U36 ( .A(A[6]), .B(n19), .Y(ab_6__7_) );
  AND2X1 U37 ( .A(A[8]), .B(n19), .Y(ab_8__7_) );
  AND2X1 U38 ( .A(A[10]), .B(n19), .Y(ab_10__7_) );
  AND2X1 U39 ( .A(A[11]), .B(B[0]), .Y(ab_11__0_) );
  AND2X1 U40 ( .A(A[10]), .B(B[0]), .Y(ab_10__0_) );
  AND2X1 U41 ( .A(A[9]), .B(B[0]), .Y(ab_9__0_) );
  AND2X1 U42 ( .A(A[8]), .B(B[0]), .Y(ab_8__0_) );
  AND2X1 U43 ( .A(A[6]), .B(B[0]), .Y(ab_6__0_) );
  AND2X1 U44 ( .A(A[7]), .B(B[0]), .Y(ab_7__0_) );
  AND2X1 U45 ( .A(A[9]), .B(n19), .Y(ab_9__7_) );
  INVXL U46 ( .A(B[0]), .Y(n37) );
  INVX4 U47 ( .A(B[4]), .Y(n26) );
  NOR2XL U48 ( .A(n36), .B(n29), .Y(ab_12__1_) );
  XOR2X2 U49 ( .A(CARRYB_16__0_), .B(SUMB_16__1_), .Y(A1_15_) );
  AND2X2 U50 ( .A(CARRYB_16__1_), .B(SUMB_16__2_), .Y(n14) );
  AND2X1 U51 ( .A(CARRYB_16__2_), .B(SUMB_16__3_), .Y(n15) );
  AND2X1 U52 ( .A(CARRYB_16__3_), .B(SUMB_16__4_), .Y(n16) );
  NOR2X1 U53 ( .A(n32), .B(n28), .Y(ab_16__2_) );
  NOR2XL U54 ( .A(n32), .B(n27), .Y(ab_16__3_) );
  NOR2X1 U55 ( .A(n32), .B(n29), .Y(ab_16__1_) );
  AND2X1 U56 ( .A(A[11]), .B(B[1]), .Y(ab_11__1_) );
  AND2X1 U57 ( .A(A[11]), .B(B[3]), .Y(ab_11__3_) );
  AND2X1 U58 ( .A(A[10]), .B(B[3]), .Y(ab_10__3_) );
  AND2X1 U59 ( .A(A[10]), .B(B[1]), .Y(ab_10__1_) );
  AND2X1 U60 ( .A(A[9]), .B(B[3]), .Y(ab_9__3_) );
  AND2X1 U61 ( .A(A[8]), .B(B[3]), .Y(ab_8__3_) );
  AND2X1 U62 ( .A(A[9]), .B(B[1]), .Y(ab_9__1_) );
  AND2X1 U63 ( .A(A[7]), .B(B[3]), .Y(ab_7__3_) );
  AND2X1 U64 ( .A(A[8]), .B(B[1]), .Y(ab_8__1_) );
  AND2X1 U65 ( .A(A[6]), .B(B[3]), .Y(ab_6__3_) );
  AND2X1 U66 ( .A(A[7]), .B(B[1]), .Y(ab_7__1_) );
  AND2X2 U67 ( .A(A[7]), .B(n19), .Y(ab_7__7_) );
  AND2X1 U68 ( .A(A[5]), .B(n19), .Y(ab_5__7_) );
  AND2X1 U69 ( .A(A[5]), .B(B[3]), .Y(ab_5__3_) );
  AND2X2 U70 ( .A(A[4]), .B(n19), .Y(ab_4__7_) );
  AND2X1 U71 ( .A(A[6]), .B(B[1]), .Y(ab_6__1_) );
  AND2X1 U72 ( .A(A[4]), .B(B[3]), .Y(ab_4__3_) );
  AND2X1 U73 ( .A(A[5]), .B(B[1]), .Y(ab_5__1_) );
  AND2X1 U74 ( .A(A[4]), .B(B[1]), .Y(ab_4__1_) );
  AND2X1 U75 ( .A(A[5]), .B(B[0]), .Y(ab_5__0_) );
  AND2X2 U76 ( .A(A[4]), .B(B[0]), .Y(ab_4__0_) );
  XOR2X1 U77 ( .A(n31), .B(ab_0__2_), .Y(SUMB_1__1_) );
  XOR2X2 U78 ( .A(CARRYB_16__4_), .B(SUMB_16__5_), .Y(A1_19_) );
  XOR2X1 U79 ( .A(CARRYB_16__5_), .B(SUMB_16__6_), .Y(A1_20_) );
  XOR2X1 U80 ( .A(CARRYB_16__6_), .B(ab_16__7_), .Y(A1_21_) );
  AND2X1 U81 ( .A(CARRYB_16__4_), .B(SUMB_16__5_), .Y(n17) );
  AND2X2 U82 ( .A(CARRYB_16__5_), .B(SUMB_16__6_), .Y(n18) );
  INVXL U83 ( .A(B[1]), .Y(n29) );
  NOR2XL U84 ( .A(n32), .B(n30), .Y(ab_16__7_) );
  NOR2X1 U85 ( .A(n24), .B(n20), .Y(ab_1__6_) );
  NOR2XL U86 ( .A(n33), .B(n30), .Y(ab_15__7_) );
  NOR2X1 U87 ( .A(n34), .B(n29), .Y(ab_14__1_) );
  NOR2X1 U88 ( .A(n35), .B(n29), .Y(ab_13__1_) );
  NOR2XL U89 ( .A(n36), .B(n28), .Y(ab_12__2_) );
  NOR2XL U90 ( .A(n35), .B(n28), .Y(ab_13__2_) );
  NOR2XL U91 ( .A(n33), .B(n28), .Y(ab_15__2_) );
  NOR2XL U92 ( .A(n36), .B(n27), .Y(ab_12__3_) );
  NOR2XL U93 ( .A(n35), .B(n27), .Y(ab_13__3_) );
  NOR2XL U94 ( .A(n34), .B(n27), .Y(ab_14__3_) );
  NOR2XL U95 ( .A(n33), .B(n27), .Y(ab_15__3_) );
  AND2X1 U96 ( .A(A[11]), .B(n19), .Y(ab_11__7_) );
  AND2X1 U97 ( .A(A[2]), .B(n19), .Y(ab_2__7_) );
  NOR2X1 U98 ( .A(n23), .B(n22), .Y(CARRYB_1__0_) );
  XOR2X1 U99 ( .A(ab_1__5_), .B(ab_0__6_), .Y(SUMB_1__5_) );
  AND2X1 U100 ( .A(A[2]), .B(B[4]), .Y(ab_2__4_) );
  XOR2X1 U101 ( .A(ab_1__4_), .B(ab_0__5_), .Y(SUMB_1__4_) );
  XOR2X1 U102 ( .A(ab_1__3_), .B(ab_0__4_), .Y(SUMB_1__3_) );
  NOR2X1 U103 ( .A(n33), .B(n29), .Y(ab_15__1_) );
  NOR2XL U104 ( .A(n34), .B(n28), .Y(ab_14__2_) );
  NOR2XL U105 ( .A(n35), .B(n30), .Y(ab_13__7_) );
  NOR2XL U106 ( .A(n34), .B(n30), .Y(ab_14__7_) );
  NOR2XL U107 ( .A(n36), .B(n30), .Y(ab_12__7_) );
  AND2X2 U108 ( .A(A[2]), .B(B[0]), .Y(ab_2__0_) );
  INVX1 U109 ( .A(A[16]), .Y(n32) );
  AND2X1 U110 ( .A(A[2]), .B(B[5]), .Y(ab_2__5_) );
  AND2X1 U111 ( .A(A[8]), .B(B[5]), .Y(ab_8__5_) );
  AND2X1 U112 ( .A(A[7]), .B(B[5]), .Y(ab_7__5_) );
  AND2X1 U113 ( .A(A[9]), .B(B[5]), .Y(ab_9__5_) );
  AND2X1 U114 ( .A(A[10]), .B(B[5]), .Y(ab_10__5_) );
  AND2X1 U115 ( .A(A[6]), .B(B[5]), .Y(ab_6__5_) );
  AND2X1 U116 ( .A(A[11]), .B(B[5]), .Y(ab_11__5_) );
  NAND2XL U117 ( .A(A[0]), .B(B[0]), .Y(n22) );
  AND2X1 U118 ( .A(A[5]), .B(B[5]), .Y(ab_5__5_) );
  AND2X1 U119 ( .A(A[4]), .B(B[5]), .Y(ab_4__5_) );
  INVX1 U120 ( .A(A[12]), .Y(n36) );
  INVX1 U121 ( .A(A[13]), .Y(n35) );
  INVX1 U122 ( .A(A[14]), .Y(n34) );
  INVX1 U123 ( .A(A[15]), .Y(n33) );
  XOR2X4 U124 ( .A(CARRYB_16__2_), .B(SUMB_16__3_), .Y(A1_17_) );
  AND2X2 U125 ( .A(A[1]), .B(B[1]), .Y(n31) );
  AND2X2 U126 ( .A(A[1]), .B(B[4]), .Y(ab_1__4_) );
  INVXL U127 ( .A(A[1]), .Y(n20) );
  INVX4 U128 ( .A(B[5]), .Y(n25) );
  AND2X1 U129 ( .A(A[3]), .B(n19), .Y(ab_3__7_) );
  AND2X1 U130 ( .A(A[3]), .B(B[5]), .Y(ab_3__5_) );
  AND2X1 U131 ( .A(A[3]), .B(B[4]), .Y(ab_3__4_) );
  AND2X1 U132 ( .A(A[3]), .B(B[3]), .Y(ab_3__3_) );
  AND2X1 U133 ( .A(A[3]), .B(B[1]), .Y(ab_3__1_) );
  NOR2X2 U134 ( .A(n25), .B(n21), .Y(ab_0__5_) );
  AND2X1 U135 ( .A(A[11]), .B(B[6]), .Y(ab_11__6_) );
  AND2X1 U136 ( .A(A[10]), .B(B[6]), .Y(ab_10__6_) );
  AND2X1 U137 ( .A(A[9]), .B(B[6]), .Y(ab_9__6_) );
  AND2X1 U138 ( .A(A[8]), .B(B[6]), .Y(ab_8__6_) );
  AND2X1 U139 ( .A(A[7]), .B(B[6]), .Y(ab_7__6_) );
  AND2X1 U140 ( .A(A[6]), .B(B[6]), .Y(ab_6__6_) );
  AND2X1 U141 ( .A(A[5]), .B(B[6]), .Y(ab_5__6_) );
  AND2X1 U142 ( .A(A[4]), .B(B[6]), .Y(ab_4__6_) );
  AND2X1 U143 ( .A(A[3]), .B(B[6]), .Y(ab_3__6_) );
  AND2X1 U144 ( .A(A[2]), .B(B[6]), .Y(ab_2__6_) );
  NOR2XL U145 ( .A(n32), .B(n26), .Y(ab_16__4_) );
  NOR2XL U146 ( .A(n33), .B(n26), .Y(ab_15__4_) );
  NOR2XL U147 ( .A(n34), .B(n26), .Y(ab_14__4_) );
  NOR2XL U148 ( .A(n35), .B(n26), .Y(ab_13__4_) );
  NOR2XL U149 ( .A(n36), .B(n26), .Y(ab_12__4_) );
  AND2X1 U150 ( .A(A[11]), .B(B[2]), .Y(ab_11__2_) );
  AND2X1 U151 ( .A(A[10]), .B(B[2]), .Y(ab_10__2_) );
  AND2X1 U152 ( .A(A[9]), .B(B[2]), .Y(ab_9__2_) );
  AND2X1 U153 ( .A(A[8]), .B(B[2]), .Y(ab_8__2_) );
  AND2X1 U154 ( .A(A[6]), .B(B[2]), .Y(ab_6__2_) );
  AND2X1 U155 ( .A(A[5]), .B(B[2]), .Y(ab_5__2_) );
  AND2X1 U156 ( .A(A[4]), .B(B[2]), .Y(ab_4__2_) );
  AND2X1 U157 ( .A(A[3]), .B(B[2]), .Y(ab_3__2_) );
  AND2X2 U158 ( .A(A[2]), .B(B[2]), .Y(ab_2__2_) );
  NOR2XL U159 ( .A(n32), .B(n24), .Y(ab_16__6_) );
  NOR2XL U160 ( .A(n33), .B(n24), .Y(ab_15__6_) );
  NOR2XL U161 ( .A(n34), .B(n24), .Y(ab_14__6_) );
  NOR2XL U162 ( .A(n35), .B(n24), .Y(ab_13__6_) );
  NOR2XL U163 ( .A(n36), .B(n24), .Y(ab_12__6_) );
  NOR2XL U164 ( .A(n32), .B(n25), .Y(ab_16__5_) );
  NOR2XL U165 ( .A(n33), .B(n25), .Y(ab_15__5_) );
  NOR2XL U166 ( .A(n34), .B(n25), .Y(ab_14__5_) );
  NOR2XL U167 ( .A(n35), .B(n25), .Y(ab_13__5_) );
  NOR2XL U168 ( .A(n36), .B(n25), .Y(ab_12__5_) );
  AND2X1 U169 ( .A(A[11]), .B(B[4]), .Y(ab_11__4_) );
  AND2X1 U170 ( .A(A[10]), .B(B[4]), .Y(ab_10__4_) );
  AND2X1 U171 ( .A(A[9]), .B(B[4]), .Y(ab_9__4_) );
  AND2X1 U172 ( .A(A[8]), .B(B[4]), .Y(ab_8__4_) );
  AND2X1 U173 ( .A(A[7]), .B(B[4]), .Y(ab_7__4_) );
  AND2X1 U174 ( .A(A[6]), .B(B[4]), .Y(ab_6__4_) );
  AND2X1 U175 ( .A(A[5]), .B(B[4]), .Y(ab_5__4_) );
  AND2X1 U176 ( .A(A[4]), .B(B[4]), .Y(ab_4__4_) );
  AND2X2 U177 ( .A(A[1]), .B(B[3]), .Y(ab_1__3_) );
  AND2X1 U178 ( .A(A[1]), .B(n19), .Y(ab_1__7_) );
  NAND2XL U179 ( .A(A[1]), .B(B[1]), .Y(n23) );
  NOR2X1 U181 ( .A(n37), .B(n32), .Y(ab_16__0_) );
  NOR2X1 U182 ( .A(n37), .B(n33), .Y(ab_15__0_) );
  NOR2X1 U183 ( .A(n37), .B(n34), .Y(ab_14__0_) );
  NOR2X1 U184 ( .A(n37), .B(n35), .Y(ab_13__0_) );
  NOR2X1 U185 ( .A(n37), .B(n36), .Y(ab_12__0_) );
endmodule


module multi16_9 ( in_17bit, in_8bit, out );
  input [16:0] in_17bit;
  input [7:0] in_8bit;
  output [16:0] out;
  wire   N19, N20, N21, N32, N33, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n55, n56, n57, n58, n59, n60, n61, n63, n64, n65, n66, n67, n68, n69,
         n71, n72, n73, n74, n75, n76, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n126, n127, n128, n129;
  wire   [16:1] in_17bit_b;
  wire   [7:0] in_8bit_b;
  wire   [23:8] mul;
  wire   [16:13] sub_add_52_b0_carry;

  multi16_9_DW02_mult_0 mult_55 ( .A({in_17bit_b, in_17bit[0]}), .B(in_8bit_b), 
        .PRODUCT_23_(mul[23]), .PRODUCT_22_(mul[22]), .PRODUCT_21_(mul[21]), 
        .PRODUCT_20_(mul[20]), .PRODUCT_19_(mul[19]), .PRODUCT_18_(mul[18]), 
        .PRODUCT_17_(mul[17]), .PRODUCT_16_(mul[16]), .PRODUCT_15_(mul[15]), 
        .PRODUCT_14_(mul[14]), .PRODUCT_13_(mul[13]), .PRODUCT_12_(mul[12]), 
        .PRODUCT_11_(mul[11]), .PRODUCT_10_(mul[10]), .PRODUCT_9_(mul[9]), 
        .PRODUCT_8_(mul[8]), .PRODUCT_7_(N32) );
  INVX4 U2 ( .A(n110), .Y(n4) );
  NAND2BX2 U3 ( .AN(mul[20]), .B(n3), .Y(n112) );
  NAND4BX2 U4 ( .AN(in_8bit[2]), .B(n37), .C(n36), .D(n35), .Y(n40) );
  INVX2 U5 ( .A(n32), .Y(n36) );
  NOR2X2 U6 ( .A(n15), .B(n44), .Y(n1) );
  NOR2X4 U7 ( .A(n2), .B(n43), .Y(in_17bit_b[1]) );
  INVX4 U8 ( .A(n1), .Y(n2) );
  NOR2X4 U9 ( .A(n42), .B(n41), .Y(n43) );
  NOR2X4 U10 ( .A(n9), .B(n107), .Y(n106) );
  INVX2 U11 ( .A(n115), .Y(n117) );
  XOR2X4 U12 ( .A(mul[19]), .B(n109), .Y(out[12]) );
  NOR2X4 U13 ( .A(n9), .B(n110), .Y(n109) );
  CLKINVX4 U14 ( .A(n108), .Y(n110) );
  NOR2X4 U15 ( .A(mul[19]), .B(n4), .Y(n3) );
  AOI21X1 U16 ( .A0(n33), .A1(n36), .B0(n17), .Y(n34) );
  NOR2XL U17 ( .A(in_8bit[4]), .B(in_8bit[2]), .Y(n33) );
  NOR3XL U18 ( .A(in_8bit[6]), .B(n18), .C(n40), .Y(in_8bit_b[7]) );
  NAND2XL U19 ( .A(in_8bit[0]), .B(n16), .Y(n23) );
  CLKINVX2 U20 ( .A(in_8bit[0]), .Y(n30) );
  INVX1 U21 ( .A(n10), .Y(n14) );
  OAI21XL U22 ( .A0(in_8bit[2]), .A1(n25), .B0(n16), .Y(n26) );
  INVX2 U23 ( .A(in_17bit[3]), .Y(n45) );
  NOR2X2 U24 ( .A(n21), .B(n14), .Y(n46) );
  XOR2X2 U25 ( .A(in_8bit[2]), .B(n24), .Y(in_8bit_b[2]) );
  NOR2X2 U26 ( .A(n17), .B(n27), .Y(n24) );
  XNOR2X1 U27 ( .A(n50), .B(n51), .Y(in_17bit_b[5]) );
  NOR2XL U28 ( .A(n21), .B(n52), .Y(n50) );
  XNOR2X2 U29 ( .A(n34), .B(n37), .Y(in_8bit_b[5]) );
  XNOR2X1 U30 ( .A(n57), .B(n58), .Y(in_17bit_b[7]) );
  INVX1 U31 ( .A(n96), .Y(n98) );
  NAND2BX1 U32 ( .AN(mul[12]), .B(n89), .Y(n90) );
  XNOR2X1 U33 ( .A(n48), .B(n7), .Y(in_17bit_b[4]) );
  XOR2X1 U34 ( .A(n19), .B(n23), .Y(in_8bit_b[1]) );
  NAND2BX2 U35 ( .AN(mul[18]), .B(n107), .Y(n108) );
  INVX1 U36 ( .A(n112), .Y(n114) );
  INVX1 U37 ( .A(in_8bit[5]), .Y(n37) );
  NAND2BX1 U38 ( .AN(mul[21]), .B(n114), .Y(n115) );
  INVX1 U39 ( .A(mul[22]), .Y(n116) );
  INVX1 U40 ( .A(n18), .Y(n16) );
  INVX2 U41 ( .A(in_17bit[16]), .Y(n21) );
  NOR2X4 U42 ( .A(n9), .B(n117), .Y(n5) );
  NAND2X2 U43 ( .A(in_17bit[0]), .B(n20), .Y(n41) );
  XOR2X2 U44 ( .A(mul[18]), .B(n106), .Y(out[11]) );
  INVX1 U45 ( .A(in_17bit[1]), .Y(n42) );
  NOR2X4 U46 ( .A(n21), .B(n15), .Y(n11) );
  NOR2X4 U47 ( .A(in_17bit[1]), .B(in_17bit[0]), .Y(n15) );
  NAND2BX1 U48 ( .AN(in_8bit[1]), .B(n30), .Y(n25) );
  XOR2X2 U49 ( .A(in_17bit[2]), .B(n11), .Y(in_17bit_b[2]) );
  CLKINVX8 U50 ( .A(in_8bit[3]), .Y(n31) );
  XOR2X2 U51 ( .A(mul[17]), .B(n103), .Y(out[10]) );
  NOR2X2 U52 ( .A(n9), .B(n104), .Y(n103) );
  CLKINVX3 U53 ( .A(n102), .Y(n104) );
  NOR2X1 U54 ( .A(in_17bit[1]), .B(n20), .Y(n44) );
  INVX8 U55 ( .A(n22), .Y(n20) );
  CLKINVX8 U56 ( .A(in_17bit[16]), .Y(n22) );
  AOI21X2 U57 ( .A0(n28), .A1(n27), .B0(n17), .Y(n29) );
  NOR2X2 U58 ( .A(n9), .B(n114), .Y(n113) );
  NAND2X2 U59 ( .A(n40), .B(n16), .Y(n38) );
  NAND2BX1 U60 ( .AN(mul[14]), .B(n95), .Y(n96) );
  INVXL U61 ( .A(in_8bit[6]), .Y(n39) );
  NAND2BXL U62 ( .AN(mul[8]), .B(n120), .Y(n78) );
  INVX2 U63 ( .A(n25), .Y(n27) );
  XNOR2X4 U64 ( .A(n5), .B(n116), .Y(out[15]) );
  NOR2XL U65 ( .A(n9), .B(n92), .Y(n91) );
  XNOR2X2 U66 ( .A(n55), .B(n6), .Y(in_17bit_b[6]) );
  AND2X1 U67 ( .A(n53), .B(n20), .Y(n6) );
  AND2X1 U68 ( .A(n47), .B(n20), .Y(n7) );
  NAND2X1 U69 ( .A(n52), .B(n51), .Y(n53) );
  NAND2BXL U70 ( .AN(n47), .B(n48), .Y(n49) );
  NAND2BXL U71 ( .AN(n53), .B(n55), .Y(n56) );
  NAND2XL U72 ( .A(n69), .B(n20), .Y(n68) );
  AND2X2 U73 ( .A(n72), .B(n71), .Y(n8) );
  NAND2XL U74 ( .A(n67), .B(n66), .Y(n69) );
  NAND2XL U75 ( .A(n59), .B(n58), .Y(n61) );
  NAND2XL U76 ( .A(n8), .B(n75), .Y(n74) );
  NAND2BXL U77 ( .AN(n61), .B(n63), .Y(n64) );
  AND2X1 U78 ( .A(N21), .B(n20), .Y(in_17bit_b[16]) );
  XNOR2X1 U79 ( .A(n20), .B(n16), .Y(n9) );
  NAND2BXL U80 ( .AN(in_17bit[2]), .B(n15), .Y(n10) );
  INVXL U81 ( .A(in_17bit[5]), .Y(n51) );
  INVXL U82 ( .A(in_17bit[4]), .Y(n48) );
  MX2X1 U83 ( .A(in_17bit[13]), .B(n12), .S0(n20), .Y(in_17bit_b[13]) );
  XNOR2X1 U84 ( .A(n76), .B(n122), .Y(n12) );
  MX2X1 U85 ( .A(in_17bit[14]), .B(N19), .S0(n20), .Y(in_17bit_b[14]) );
  MX2X1 U86 ( .A(in_17bit[15]), .B(N20), .S0(n20), .Y(in_17bit_b[15]) );
  INVXL U87 ( .A(in_17bit[7]), .Y(n58) );
  INVXL U88 ( .A(in_17bit[6]), .Y(n55) );
  INVXL U89 ( .A(in_17bit[8]), .Y(n63) );
  MX2X1 U90 ( .A(in_17bit[12]), .B(n13), .S0(n20), .Y(in_17bit_b[12]) );
  XNOR2X1 U91 ( .A(n74), .B(n121), .Y(n13) );
  NAND2BX1 U92 ( .AN(mul[16]), .B(n101), .Y(n102) );
  INVX1 U93 ( .A(n81), .Y(n83) );
  NAND2BX1 U94 ( .AN(mul[9]), .B(n80), .Y(n81) );
  INVX1 U95 ( .A(n84), .Y(n86) );
  NAND2BX1 U96 ( .AN(mul[10]), .B(n83), .Y(n84) );
  INVX1 U97 ( .A(n87), .Y(n89) );
  NAND2BX1 U98 ( .AN(mul[11]), .B(n86), .Y(n87) );
  INVX1 U99 ( .A(n78), .Y(n80) );
  INVX1 U100 ( .A(N32), .Y(n120) );
  INVX1 U101 ( .A(n99), .Y(n101) );
  NAND2BX1 U102 ( .AN(mul[15]), .B(n98), .Y(n99) );
  INVX1 U103 ( .A(n93), .Y(n95) );
  NAND2BX1 U104 ( .AN(mul[13]), .B(n92), .Y(n93) );
  INVX1 U105 ( .A(n90), .Y(n92) );
  XOR2X1 U106 ( .A(mul[16]), .B(n100), .Y(out[9]) );
  NOR2XL U107 ( .A(n9), .B(n101), .Y(n100) );
  XOR2X1 U108 ( .A(mul[14]), .B(n94), .Y(out[7]) );
  NOR2XL U109 ( .A(n9), .B(n95), .Y(n94) );
  XOR2X1 U110 ( .A(mul[15]), .B(n97), .Y(out[8]) );
  NOR2XL U111 ( .A(n9), .B(n98), .Y(n97) );
  XOR2X1 U112 ( .A(mul[11]), .B(n85), .Y(out[4]) );
  NOR2X1 U113 ( .A(n9), .B(n86), .Y(n85) );
  XOR2X1 U114 ( .A(mul[9]), .B(n79), .Y(out[2]) );
  NOR2X1 U115 ( .A(n9), .B(n80), .Y(n79) );
  XOR2X1 U116 ( .A(mul[12]), .B(n88), .Y(out[5]) );
  NOR2X1 U117 ( .A(n9), .B(n89), .Y(n88) );
  XOR2X1 U118 ( .A(mul[10]), .B(n82), .Y(out[3]) );
  NOR2X1 U119 ( .A(n9), .B(n83), .Y(n82) );
  XOR2X1 U120 ( .A(mul[13]), .B(n91), .Y(out[6]) );
  XOR2X1 U121 ( .A(mul[23]), .B(n118), .Y(out[16]) );
  INVX1 U122 ( .A(n128), .Y(out[1]) );
  AOI22X1 U123 ( .A0(mul[8]), .A1(n9), .B0(N33), .B1(n129), .Y(n128) );
  INVX1 U124 ( .A(mul[8]), .Y(n119) );
  INVX1 U125 ( .A(n127), .Y(out[0]) );
  AOI22XL U126 ( .A0(N32), .A1(n9), .B0(N32), .B1(n129), .Y(n127) );
  INVXL U127 ( .A(n9), .Y(n129) );
  INVXL U128 ( .A(in_8bit[1]), .Y(n19) );
  INVX1 U129 ( .A(n126), .Y(in_8bit_b[0]) );
  AOI22XL U130 ( .A0(in_8bit[0]), .A1(n16), .B0(in_8bit[0]), .B1(n17), .Y(n126) );
  XNOR2X1 U131 ( .A(n65), .B(n66), .Y(in_17bit_b[9]) );
  NOR2X1 U132 ( .A(n21), .B(n67), .Y(n65) );
  NOR2X1 U133 ( .A(n21), .B(n59), .Y(n57) );
  XNOR2X1 U134 ( .A(n73), .B(n75), .Y(in_17bit_b[11]) );
  NOR2X1 U135 ( .A(n21), .B(n8), .Y(n73) );
  XOR2X1 U136 ( .A(n63), .B(n60), .Y(in_17bit_b[8]) );
  XOR2X1 U137 ( .A(n71), .B(n68), .Y(in_17bit_b[10]) );
  INVX1 U138 ( .A(n49), .Y(n52) );
  INVX1 U139 ( .A(n56), .Y(n59) );
  INVX1 U140 ( .A(n64), .Y(n67) );
  NAND3BXL U141 ( .AN(in_8bit[1]), .B(n31), .C(n30), .Y(n32) );
  INVX1 U142 ( .A(n69), .Y(n72) );
  INVX1 U143 ( .A(in_8bit[7]), .Y(n17) );
  INVX1 U144 ( .A(in_8bit[7]), .Y(n18) );
  NAND3X1 U145 ( .A(n121), .B(n8), .C(n75), .Y(n76) );
  INVX1 U146 ( .A(n76), .Y(sub_add_52_b0_carry[13]) );
  NOR2XL U147 ( .A(in_8bit[3]), .B(in_8bit[2]), .Y(n28) );
  NAND2BXL U148 ( .AN(in_17bit[3]), .B(n14), .Y(n47) );
  INVX1 U149 ( .A(in_17bit[9]), .Y(n66) );
  INVX1 U150 ( .A(in_17bit[11]), .Y(n75) );
  INVX1 U151 ( .A(in_17bit[10]), .Y(n71) );
  INVX1 U152 ( .A(in_17bit[12]), .Y(n121) );
  INVX1 U153 ( .A(in_17bit[13]), .Y(n122) );
  INVX1 U154 ( .A(in_17bit[14]), .Y(n123) );
  INVX1 U155 ( .A(in_17bit[15]), .Y(n124) );
  INVX1 U156 ( .A(in_8bit[4]), .Y(n35) );
  NAND2XL U157 ( .A(n61), .B(n20), .Y(n60) );
  AOI21XL U158 ( .A0(n117), .A1(n116), .B0(n9), .Y(n118) );
  INVX4 U159 ( .A(n105), .Y(n107) );
  XOR2X4 U160 ( .A(n26), .B(n31), .Y(in_8bit_b[3]) );
  XNOR2X4 U161 ( .A(n29), .B(n35), .Y(in_8bit_b[4]) );
  XOR2X4 U162 ( .A(n39), .B(n38), .Y(in_8bit_b[6]) );
  XNOR2X4 U163 ( .A(n46), .B(n45), .Y(in_17bit_b[3]) );
  NAND2BX4 U164 ( .AN(mul[17]), .B(n104), .Y(n105) );
  NOR2X4 U165 ( .A(n9), .B(n3), .Y(n111) );
  XOR2X4 U166 ( .A(mul[20]), .B(n111), .Y(out[13]) );
  XOR2X4 U167 ( .A(n113), .B(mul[21]), .Y(out[14]) );
  XOR2X1 U168 ( .A(n119), .B(n120), .Y(N33) );
  XOR2X1 U169 ( .A(n21), .B(sub_add_52_b0_carry[16]), .Y(N21) );
  AND2X1 U170 ( .A(sub_add_52_b0_carry[15]), .B(n124), .Y(
        sub_add_52_b0_carry[16]) );
  XOR2X1 U171 ( .A(n124), .B(sub_add_52_b0_carry[15]), .Y(N20) );
  AND2X1 U172 ( .A(sub_add_52_b0_carry[14]), .B(n123), .Y(
        sub_add_52_b0_carry[15]) );
  XOR2X1 U173 ( .A(n123), .B(sub_add_52_b0_carry[14]), .Y(N19) );
  AND2X1 U174 ( .A(sub_add_52_b0_carry[13]), .B(n122), .Y(
        sub_add_52_b0_carry[14]) );
endmodule


module multi16_8_DW01_add_0 ( A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, 
        A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, 
        B_20_, B_19_, B_18_, B_17_, B_16_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, 
        SUM_17_, SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, 
        SUM_9_, SUM_8_, SUM_7_, SUM_6_, SUM_5_ );
  input A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_,
         A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, B_20_, B_19_,
         B_18_, B_17_, B_16_;
  output SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, SUM_15_,
         SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, SUM_7_,
         SUM_6_, SUM_5_;
  wire   n1, n2, n3, n4, n5, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43;

  NAND2X4 U2 ( .A(B_16_), .B(A_16_), .Y(n37) );
  AOI21X4 U3 ( .A0(n22), .A1(n23), .B0(n21), .Y(n41) );
  NOR2X4 U4 ( .A(n21), .B(n33), .Y(n43) );
  NAND2X1 U5 ( .A(n42), .B(n2), .Y(n3) );
  NAND2X2 U6 ( .A(n1), .B(n41), .Y(n4) );
  NAND2X4 U7 ( .A(n3), .B(n4), .Y(SUM_18_) );
  INVX1 U8 ( .A(n42), .Y(n1) );
  INVXL U9 ( .A(n41), .Y(n2) );
  NAND2X1 U10 ( .A(n36), .B(n19), .Y(n42) );
  XOR2X2 U11 ( .A(n23), .B(n43), .Y(SUM_17_) );
  BUFX3 U12 ( .A(A_13_), .Y(SUM_13_) );
  BUFX3 U13 ( .A(A_14_), .Y(SUM_14_) );
  NOR2X1 U14 ( .A(B_18_), .B(A_18_), .Y(n34) );
  INVX1 U15 ( .A(n34), .Y(n19) );
  XOR2X1 U16 ( .A(n39), .B(n40), .Y(SUM_19_) );
  NOR2BX1 U17 ( .AN(n32), .B(n31), .Y(n40) );
  OAI21XL U18 ( .A0(n41), .A1(n34), .B0(n36), .Y(n39) );
  NOR2X2 U19 ( .A(B_16_), .B(A_16_), .Y(n17) );
  NOR2X4 U20 ( .A(n23), .B(n17), .Y(SUM_16_) );
  INVX4 U21 ( .A(n37), .Y(n23) );
  OAI21X1 U22 ( .A0(n30), .A1(n31), .B0(n32), .Y(n27) );
  AOI21XL U23 ( .A0(n19), .A1(n35), .B0(n20), .Y(n30) );
  INVX4 U24 ( .A(n24), .Y(SUM_15_) );
  CLKINVX4 U25 ( .A(A_15_), .Y(n24) );
  NAND2X4 U26 ( .A(B_17_), .B(A_17_), .Y(n38) );
  INVX4 U27 ( .A(n33), .Y(n22) );
  INVXL U28 ( .A(n29), .Y(n18) );
  XOR2X1 U29 ( .A(n5), .B(n27), .Y(SUM_20_) );
  NAND2XL U30 ( .A(B_18_), .B(A_18_), .Y(n36) );
  BUFX4 U31 ( .A(A_12_), .Y(SUM_12_) );
  INVX1 U32 ( .A(n36), .Y(n20) );
  AND2X2 U33 ( .A(n29), .B(n28), .Y(n5) );
  BUFX3 U34 ( .A(A_10_), .Y(SUM_10_) );
  BUFX3 U35 ( .A(A_11_), .Y(SUM_11_) );
  BUFX3 U36 ( .A(A_9_), .Y(SUM_9_) );
  BUFX3 U37 ( .A(A_5_), .Y(SUM_5_) );
  BUFX3 U38 ( .A(A_6_), .Y(SUM_6_) );
  BUFX3 U39 ( .A(A_7_), .Y(SUM_7_) );
  BUFX3 U40 ( .A(A_8_), .Y(SUM_8_) );
  INVX4 U41 ( .A(n38), .Y(n21) );
  NOR2X4 U42 ( .A(B_17_), .B(A_17_), .Y(n33) );
  XOR2X1 U43 ( .A(n25), .B(n26), .Y(SUM_21_) );
  AOI21X1 U44 ( .A0(n27), .A1(n28), .B0(n18), .Y(n26) );
  XNOR2X1 U45 ( .A(B_21_), .B(A_21_), .Y(n25) );
  OAI21XL U46 ( .A0(n33), .A1(n37), .B0(n38), .Y(n35) );
  OR2X1 U47 ( .A(B_20_), .B(A_20_), .Y(n28) );
  NAND2X1 U48 ( .A(B_20_), .B(A_20_), .Y(n29) );
  NOR2X1 U49 ( .A(B_19_), .B(A_19_), .Y(n31) );
  NAND2X1 U50 ( .A(B_19_), .B(A_19_), .Y(n32) );
endmodule


module multi16_8_DW02_mult_0 ( A, B, PRODUCT_23_, PRODUCT_22_, PRODUCT_21_, 
        PRODUCT_20_, PRODUCT_19_, PRODUCT_18_, PRODUCT_17_, PRODUCT_16_, 
        PRODUCT_15_, PRODUCT_14_, PRODUCT_13_, PRODUCT_12_, PRODUCT_11_, 
        PRODUCT_10_, PRODUCT_9_, PRODUCT_8_, PRODUCT_7_ );
  input [16:0] A;
  input [7:0] B;
  output PRODUCT_23_, PRODUCT_22_, PRODUCT_21_, PRODUCT_20_, PRODUCT_19_,
         PRODUCT_18_, PRODUCT_17_, PRODUCT_16_, PRODUCT_15_, PRODUCT_14_,
         PRODUCT_13_, PRODUCT_12_, PRODUCT_11_, PRODUCT_10_, PRODUCT_9_,
         PRODUCT_8_, PRODUCT_7_;
  wire   ab_16__7_, ab_16__6_, ab_16__5_, ab_16__4_, ab_16__3_, ab_16__2_,
         ab_16__1_, ab_16__0_, ab_15__7_, ab_15__6_, ab_15__5_, ab_15__4_,
         ab_15__3_, ab_15__2_, ab_15__1_, ab_15__0_, ab_14__7_, ab_14__6_,
         ab_14__5_, ab_14__4_, ab_14__3_, ab_14__2_, ab_14__1_, ab_14__0_,
         ab_13__7_, ab_13__6_, ab_13__5_, ab_13__4_, ab_13__3_, ab_13__2_,
         ab_13__1_, ab_13__0_, ab_12__7_, ab_12__6_, ab_12__5_, ab_12__4_,
         ab_12__3_, ab_12__2_, ab_12__1_, ab_12__0_, ab_11__7_, ab_11__6_,
         ab_11__5_, ab_11__4_, ab_11__3_, ab_11__2_, ab_11__1_, ab_11__0_,
         ab_10__7_, ab_10__6_, ab_10__5_, ab_10__4_, ab_10__3_, ab_10__2_,
         ab_10__1_, ab_10__0_, ab_9__7_, ab_9__6_, ab_9__5_, ab_9__4_,
         ab_9__3_, ab_9__2_, ab_9__1_, ab_9__0_, ab_8__7_, ab_8__6_, ab_8__5_,
         ab_8__4_, ab_8__3_, ab_8__2_, ab_8__1_, ab_8__0_, ab_7__7_, ab_7__6_,
         ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_, ab_7__0_, ab_6__7_,
         ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_, ab_6__1_, ab_6__0_,
         ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_, ab_5__2_, ab_5__1_,
         ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_, ab_4__3_, ab_4__2_,
         ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_, ab_3__4_, ab_3__3_,
         ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_, ab_2__5_, ab_2__4_,
         ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_, ab_1__6_, ab_1__5_,
         ab_1__4_, ab_1__3_, ab_1__2_, ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_,
         ab_0__3_, ab_0__2_, CARRYB_16__6_, CARRYB_16__5_, CARRYB_16__4_,
         CARRYB_16__3_, CARRYB_16__2_, CARRYB_16__1_, CARRYB_16__0_,
         CARRYB_15__6_, CARRYB_15__5_, CARRYB_15__4_, CARRYB_15__3_,
         CARRYB_15__2_, CARRYB_15__1_, CARRYB_15__0_, CARRYB_14__6_,
         CARRYB_14__5_, CARRYB_14__4_, CARRYB_14__3_, CARRYB_14__2_,
         CARRYB_14__1_, CARRYB_14__0_, CARRYB_13__6_, CARRYB_13__5_,
         CARRYB_13__4_, CARRYB_13__3_, CARRYB_13__2_, CARRYB_13__1_,
         CARRYB_13__0_, CARRYB_12__6_, CARRYB_12__5_, CARRYB_12__4_,
         CARRYB_12__3_, CARRYB_12__2_, CARRYB_12__1_, CARRYB_12__0_,
         CARRYB_11__6_, CARRYB_11__5_, CARRYB_11__4_, CARRYB_11__3_,
         CARRYB_11__2_, CARRYB_11__1_, CARRYB_11__0_, CARRYB_10__6_,
         CARRYB_10__5_, CARRYB_10__4_, CARRYB_10__3_, CARRYB_10__2_,
         CARRYB_10__1_, CARRYB_10__0_, CARRYB_9__6_, CARRYB_9__5_,
         CARRYB_9__4_, CARRYB_9__3_, CARRYB_9__2_, CARRYB_9__1_, CARRYB_9__0_,
         CARRYB_8__6_, CARRYB_8__5_, CARRYB_8__4_, CARRYB_8__3_, CARRYB_8__2_,
         CARRYB_8__1_, CARRYB_8__0_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_,
         CARRYB_7__3_, CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_,
         CARRYB_6__5_, CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_,
         CARRYB_6__0_, CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_,
         CARRYB_5__2_, CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_,
         CARRYB_4__4_, CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_,
         CARRYB_3__6_, CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_,
         CARRYB_3__1_, CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_,
         CARRYB_2__3_, CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__1_,
         CARRYB_1__0_, SUMB_16__6_, SUMB_16__5_, SUMB_16__4_, SUMB_16__3_,
         SUMB_16__2_, SUMB_16__1_, SUMB_16__0_, SUMB_15__6_, SUMB_15__5_,
         SUMB_15__4_, SUMB_15__3_, SUMB_15__2_, SUMB_15__1_, SUMB_14__6_,
         SUMB_14__5_, SUMB_14__4_, SUMB_14__3_, SUMB_14__2_, SUMB_14__1_,
         SUMB_13__6_, SUMB_13__5_, SUMB_13__4_, SUMB_13__3_, SUMB_13__2_,
         SUMB_13__1_, SUMB_12__6_, SUMB_12__5_, SUMB_12__4_, SUMB_12__3_,
         SUMB_12__2_, SUMB_12__1_, SUMB_11__6_, SUMB_11__5_, SUMB_11__4_,
         SUMB_11__3_, SUMB_11__2_, SUMB_11__1_, SUMB_10__6_, SUMB_10__5_,
         SUMB_10__4_, SUMB_10__3_, SUMB_10__2_, SUMB_10__1_, SUMB_9__6_,
         SUMB_9__5_, SUMB_9__4_, SUMB_9__3_, SUMB_9__2_, SUMB_9__1_,
         SUMB_8__6_, SUMB_8__5_, SUMB_8__4_, SUMB_8__3_, SUMB_8__2_,
         SUMB_8__1_, SUMB_7__6_, SUMB_7__5_, SUMB_7__4_, SUMB_7__3_,
         SUMB_7__2_, SUMB_7__1_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_,
         SUMB_6__3_, SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_,
         SUMB_5__4_, SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_,
         SUMB_4__5_, SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_,
         SUMB_3__6_, SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_,
         SUMB_3__1_, SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_,
         SUMB_2__2_, SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_,
         SUMB_1__3_, SUMB_1__2_, SUMB_1__1_, PROD1_7_, A1_21_, A1_20_, A1_19_,
         A1_18_, A1_17_, A1_16_, A1_15_, A1_13_, A1_12_, A1_11_, A1_10_, A1_9_,
         A1_8_, A1_7_, A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, n4, n5, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34;

  ADDFHX4 S1_15_0 ( .A(ab_15__0_), .B(CARRYB_14__0_), .CI(SUMB_14__1_), .CO(
        CARRYB_15__0_), .S(A1_13_) );
  ADDFHX4 S1_14_0 ( .A(ab_14__0_), .B(CARRYB_13__0_), .CI(SUMB_13__1_), .CO(
        CARRYB_14__0_), .S(A1_12_) );
  ADDFHX4 S1_13_0 ( .A(ab_13__0_), .B(CARRYB_12__0_), .CI(SUMB_12__1_), .CO(
        CARRYB_13__0_), .S(A1_11_) );
  ADDFHX4 S2_13_1 ( .A(ab_13__1_), .B(CARRYB_12__1_), .CI(SUMB_12__2_), .CO(
        CARRYB_13__1_), .S(SUMB_13__1_) );
  ADDFHX4 S1_12_0 ( .A(ab_12__0_), .B(CARRYB_11__0_), .CI(SUMB_11__1_), .CO(
        CARRYB_12__0_), .S(A1_10_) );
  ADDFHX4 S2_12_1 ( .A(ab_12__1_), .B(CARRYB_11__1_), .CI(SUMB_11__2_), .CO(
        CARRYB_12__1_), .S(SUMB_12__1_) );
  ADDFHX4 S2_12_2 ( .A(ab_12__2_), .B(CARRYB_11__2_), .CI(SUMB_11__3_), .CO(
        CARRYB_12__2_), .S(SUMB_12__2_) );
  ADDFHX4 S1_11_0 ( .A(ab_11__0_), .B(CARRYB_10__0_), .CI(SUMB_10__1_), .CO(
        CARRYB_11__0_), .S(A1_9_) );
  ADDFHX4 S2_11_1 ( .A(ab_11__1_), .B(CARRYB_10__1_), .CI(SUMB_10__2_), .CO(
        CARRYB_11__1_), .S(SUMB_11__1_) );
  ADDFHX4 S2_11_2 ( .A(ab_11__2_), .B(CARRYB_10__2_), .CI(SUMB_10__3_), .CO(
        CARRYB_11__2_), .S(SUMB_11__2_) );
  ADDFHX4 S1_10_0 ( .A(ab_10__0_), .B(CARRYB_9__0_), .CI(SUMB_9__1_), .CO(
        CARRYB_10__0_), .S(A1_8_) );
  ADDFHX4 S2_10_1 ( .A(ab_10__1_), .B(CARRYB_9__1_), .CI(SUMB_9__2_), .CO(
        CARRYB_10__1_), .S(SUMB_10__1_) );
  ADDFHX4 S1_9_0 ( .A(ab_9__0_), .B(CARRYB_8__0_), .CI(SUMB_8__1_), .CO(
        CARRYB_9__0_), .S(A1_7_) );
  ADDFHX4 S2_9_1 ( .A(ab_9__1_), .B(CARRYB_8__1_), .CI(SUMB_8__2_), .CO(
        CARRYB_9__1_), .S(SUMB_9__1_) );
  ADDFHX4 S2_9_2 ( .A(ab_9__2_), .B(CARRYB_8__2_), .CI(SUMB_8__3_), .CO(
        CARRYB_9__2_), .S(SUMB_9__2_) );
  ADDFHX4 S2_9_3 ( .A(ab_9__3_), .B(CARRYB_8__3_), .CI(SUMB_8__4_), .CO(
        CARRYB_9__3_), .S(SUMB_9__3_) );
  ADDFHX4 S2_9_4 ( .A(ab_9__4_), .B(CARRYB_8__4_), .CI(SUMB_8__5_), .CO(
        CARRYB_9__4_), .S(SUMB_9__4_) );
  ADDFHX4 S1_8_0 ( .A(ab_8__0_), .B(CARRYB_7__0_), .CI(SUMB_7__1_), .CO(
        CARRYB_8__0_), .S(A1_6_) );
  ADDFHX4 S2_8_1 ( .A(ab_8__1_), .B(CARRYB_7__1_), .CI(SUMB_7__2_), .CO(
        CARRYB_8__1_), .S(SUMB_8__1_) );
  ADDFHX4 S2_8_2 ( .A(ab_8__2_), .B(CARRYB_7__2_), .CI(SUMB_7__3_), .CO(
        CARRYB_8__2_), .S(SUMB_8__2_) );
  ADDFHX4 S2_8_4 ( .A(ab_8__4_), .B(CARRYB_7__4_), .CI(SUMB_7__5_), .CO(
        CARRYB_8__4_), .S(SUMB_8__4_) );
  ADDFHX4 S2_7_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  ADDFHX4 S3_7_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(
        CARRYB_7__6_), .S(SUMB_7__6_) );
  ADDFHX4 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  ADDFHX4 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  ADDFHX4 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  ADDFHX4 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  ADDFHX4 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  ADDFHX4 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  ADDFHX4 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  ADDFHX4 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  ADDFHX4 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  ADDFHX4 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  ADDFHX4 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  ADDFHX4 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  ADDFHX4 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  ADDFHX4 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  ADDFHX4 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  ADDFHX4 S2_2_4 ( .A(ab_2__4_), .B(n4), .CI(SUMB_1__5_), .CO(CARRYB_2__4_), 
        .S(SUMB_2__4_) );
  multi16_8_DW01_add_0 FS_1 ( .A_21_(A1_21_), .A_20_(A1_20_), .A_19_(A1_19_), 
        .A_18_(A1_18_), .A_17_(A1_17_), .A_16_(A1_16_), .A_15_(A1_15_), 
        .A_14_(SUMB_16__0_), .A_13_(A1_13_), .A_12_(A1_12_), .A_11_(A1_11_), 
        .A_10_(A1_10_), .A_9_(A1_9_), .A_8_(A1_8_), .A_7_(A1_7_), .A_6_(A1_6_), 
        .A_5_(PROD1_7_), .B_21_(n14), .B_20_(n13), .B_19_(n12), .B_18_(n10), 
        .B_17_(n11), .B_16_(n9), .SUM_21_(PRODUCT_23_), .SUM_20_(PRODUCT_22_), 
        .SUM_19_(PRODUCT_21_), .SUM_18_(PRODUCT_20_), .SUM_17_(PRODUCT_19_), 
        .SUM_16_(PRODUCT_18_), .SUM_15_(PRODUCT_17_), .SUM_14_(PRODUCT_16_), 
        .SUM_13_(PRODUCT_15_), .SUM_12_(PRODUCT_14_), .SUM_11_(PRODUCT_13_), 
        .SUM_10_(PRODUCT_12_), .SUM_9_(PRODUCT_11_), .SUM_8_(PRODUCT_10_), 
        .SUM_7_(PRODUCT_9_), .SUM_6_(PRODUCT_8_), .SUM_5_(PRODUCT_7_) );
  ADDFHX2 S2_15_4 ( .A(ab_15__4_), .B(CARRYB_14__4_), .CI(SUMB_14__5_), .CO(
        CARRYB_15__4_), .S(SUMB_15__4_) );
  ADDFHX4 S2_11_4 ( .A(ab_11__4_), .B(CARRYB_10__4_), .CI(SUMB_10__5_), .CO(
        CARRYB_11__4_), .S(SUMB_11__4_) );
  ADDFHX4 S2_11_3 ( .A(ab_11__3_), .B(CARRYB_10__3_), .CI(SUMB_10__4_), .CO(
        CARRYB_11__3_), .S(SUMB_11__3_) );
  ADDFHX4 S2_12_3 ( .A(ab_12__3_), .B(CARRYB_11__3_), .CI(SUMB_11__4_), .CO(
        CARRYB_12__3_), .S(SUMB_12__3_) );
  ADDFHX4 S4_1 ( .A(ab_16__1_), .B(CARRYB_15__1_), .CI(SUMB_15__2_), .CO(
        CARRYB_16__1_), .S(SUMB_16__1_) );
  ADDFHX2 S2_8_5 ( .A(ab_8__5_), .B(CARRYB_7__5_), .CI(SUMB_7__6_), .CO(
        CARRYB_8__5_), .S(SUMB_8__5_) );
  ADDFHX4 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  ADDFHX4 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  ADDFHX4 S1_7_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(PROD1_7_) );
  ADDFHX4 S4_3 ( .A(ab_16__3_), .B(CARRYB_15__3_), .CI(SUMB_15__4_), .CO(
        CARRYB_16__3_), .S(SUMB_16__3_) );
  ADDFHX4 S2_14_2 ( .A(ab_14__2_), .B(CARRYB_13__2_), .CI(SUMB_13__3_), .CO(
        CARRYB_14__2_), .S(SUMB_14__2_) );
  ADDFHX4 S2_14_1 ( .A(ab_14__1_), .B(CARRYB_13__1_), .CI(SUMB_13__2_), .CO(
        CARRYB_14__1_), .S(SUMB_14__1_) );
  ADDFHX4 S2_15_1 ( .A(ab_15__1_), .B(CARRYB_14__1_), .CI(SUMB_14__2_), .CO(
        CARRYB_15__1_), .S(SUMB_15__1_) );
  ADDFHX4 S3_8_6 ( .A(ab_8__6_), .B(CARRYB_7__6_), .CI(ab_7__7_), .CO(
        CARRYB_8__6_), .S(SUMB_8__6_) );
  ADDFHX2 S2_15_5 ( .A(ab_15__5_), .B(CARRYB_14__5_), .CI(SUMB_14__6_), .CO(
        CARRYB_15__5_), .S(SUMB_15__5_) );
  ADDFHX4 S3_11_6 ( .A(ab_11__6_), .B(CARRYB_10__6_), .CI(ab_10__7_), .CO(
        CARRYB_11__6_), .S(SUMB_11__6_) );
  ADDFHX4 S3_2_6 ( .A(ab_2__6_), .B(n7), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  ADDFHX4 S2_9_5 ( .A(ab_9__5_), .B(CARRYB_8__5_), .CI(SUMB_8__6_), .CO(
        CARRYB_9__5_), .S(SUMB_9__5_) );
  ADDFHX2 S4_0 ( .A(ab_16__0_), .B(CARRYB_15__0_), .CI(SUMB_15__1_), .CO(
        CARRYB_16__0_), .S(SUMB_16__0_) );
  ADDFHX4 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  ADDFHX4 S2_14_4 ( .A(ab_14__4_), .B(CARRYB_13__4_), .CI(SUMB_13__5_), .CO(
        CARRYB_14__4_), .S(SUMB_14__4_) );
  ADDFHX4 S2_14_3 ( .A(ab_14__3_), .B(CARRYB_13__3_), .CI(SUMB_13__4_), .CO(
        CARRYB_14__3_), .S(SUMB_14__3_) );
  ADDFHX4 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  ADDFHX4 S2_15_2 ( .A(ab_15__2_), .B(CARRYB_14__2_), .CI(SUMB_14__3_), .CO(
        CARRYB_15__2_), .S(SUMB_15__2_) );
  ADDFHX4 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  ADDFHX4 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  ADDFHX4 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  ADDFHX4 S2_11_5 ( .A(ab_11__5_), .B(CARRYB_10__5_), .CI(SUMB_10__6_), .CO(
        CARRYB_11__5_), .S(SUMB_11__5_) );
  ADDFHX4 S2_12_4 ( .A(ab_12__4_), .B(CARRYB_11__4_), .CI(SUMB_11__5_), .CO(
        CARRYB_12__4_), .S(SUMB_12__4_) );
  ADDFHX4 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  ADDFHX4 S3_9_6 ( .A(ab_9__6_), .B(CARRYB_8__6_), .CI(ab_8__7_), .CO(
        CARRYB_9__6_), .S(SUMB_9__6_) );
  ADDFHX4 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  ADDFHX4 S2_12_5 ( .A(ab_12__5_), .B(CARRYB_11__5_), .CI(SUMB_11__6_), .CO(
        CARRYB_12__5_), .S(SUMB_12__5_) );
  ADDFHX4 S2_8_3 ( .A(ab_8__3_), .B(CARRYB_7__3_), .CI(SUMB_7__4_), .CO(
        CARRYB_8__3_), .S(SUMB_8__3_) );
  ADDFHX4 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  ADDFX2 S5_6 ( .A(ab_16__6_), .B(CARRYB_15__6_), .CI(ab_15__7_), .CO(
        CARRYB_16__6_), .S(SUMB_16__6_) );
  ADDFHX1 S4_5 ( .A(ab_16__5_), .B(CARRYB_15__5_), .CI(SUMB_15__6_), .CO(
        CARRYB_16__5_), .S(SUMB_16__5_) );
  ADDFHX2 S3_10_6 ( .A(ab_10__6_), .B(CARRYB_9__6_), .CI(ab_9__7_), .CO(
        CARRYB_10__6_), .S(SUMB_10__6_) );
  ADDFHX2 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  ADDFX1 S4_4 ( .A(ab_16__4_), .B(CARRYB_15__4_), .CI(SUMB_15__5_), .CO(
        CARRYB_16__4_), .S(SUMB_16__4_) );
  ADDFHX2 S2_2_2 ( .A(ab_2__2_), .B(n8), .CI(SUMB_1__3_), .CO(CARRYB_2__2_), 
        .S(SUMB_2__2_) );
  ADDFHX2 S4_2 ( .A(ab_16__2_), .B(CARRYB_15__2_), .CI(SUMB_15__3_), .CO(
        CARRYB_16__2_), .S(SUMB_16__2_) );
  ADDFHX2 S2_13_5 ( .A(ab_13__5_), .B(CARRYB_12__5_), .CI(SUMB_12__6_), .CO(
        CARRYB_13__5_), .S(SUMB_13__5_) );
  ADDFHX2 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  ADDFHX2 S2_2_3 ( .A(ab_2__3_), .B(n5), .CI(SUMB_1__4_), .CO(CARRYB_2__3_), 
        .S(SUMB_2__3_) );
  ADDFHX2 S2_13_2 ( .A(ab_13__2_), .B(CARRYB_12__2_), .CI(SUMB_12__3_), .CO(
        CARRYB_13__2_), .S(SUMB_13__2_) );
  ADDFHX2 S2_7_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  ADDFHX2 S2_10_5 ( .A(ab_10__5_), .B(CARRYB_9__5_), .CI(SUMB_9__6_), .CO(
        CARRYB_10__5_), .S(SUMB_10__5_) );
  ADDFHX2 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  ADDFHX2 S2_10_4 ( .A(ab_10__4_), .B(CARRYB_9__4_), .CI(SUMB_9__5_), .CO(
        CARRYB_10__4_), .S(SUMB_10__4_) );
  ADDFHX1 S3_15_6 ( .A(ab_15__6_), .B(CARRYB_14__6_), .CI(ab_14__7_), .CO(
        CARRYB_15__6_), .S(SUMB_15__6_) );
  ADDFHX2 S3_12_6 ( .A(ab_12__6_), .B(CARRYB_11__6_), .CI(ab_11__7_), .CO(
        CARRYB_12__6_), .S(SUMB_12__6_) );
  ADDFHX2 S2_2_5 ( .A(ab_2__5_), .B(n6), .CI(SUMB_1__6_), .CO(CARRYB_2__5_), 
        .S(SUMB_2__5_) );
  ADDFHX2 S2_14_5 ( .A(ab_14__5_), .B(CARRYB_13__5_), .CI(SUMB_13__6_), .CO(
        CARRYB_14__5_), .S(SUMB_14__5_) );
  ADDFHX2 S2_15_3 ( .A(ab_15__3_), .B(CARRYB_14__3_), .CI(SUMB_14__4_), .CO(
        CARRYB_15__3_), .S(SUMB_15__3_) );
  ADDFHX2 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  ADDFHX4 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  ADDFHX4 S2_7_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  ADDFHX2 S3_13_6 ( .A(ab_13__6_), .B(CARRYB_12__6_), .CI(ab_12__7_), .CO(
        CARRYB_13__6_), .S(SUMB_13__6_) );
  ADDFHX2 S3_14_6 ( .A(ab_14__6_), .B(CARRYB_13__6_), .CI(ab_13__7_), .CO(
        CARRYB_14__6_), .S(SUMB_14__6_) );
  ADDFHX4 S2_13_3 ( .A(ab_13__3_), .B(CARRYB_12__3_), .CI(SUMB_12__4_), .CO(
        CARRYB_13__3_), .S(SUMB_13__3_) );
  ADDFHX4 S2_10_3 ( .A(ab_10__3_), .B(CARRYB_9__3_), .CI(SUMB_9__4_), .CO(
        CARRYB_10__3_), .S(SUMB_10__3_) );
  ADDFHX4 S2_10_2 ( .A(ab_10__2_), .B(CARRYB_9__2_), .CI(SUMB_9__3_), .CO(
        CARRYB_10__2_), .S(SUMB_10__2_) );
  ADDFHX4 S2_7_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  ADDFHX4 S2_7_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  ADDFHX4 S2_13_4 ( .A(ab_13__4_), .B(CARRYB_12__4_), .CI(SUMB_12__5_), .CO(
        CARRYB_13__4_), .S(SUMB_13__4_) );
  NOR2X1 U2 ( .A(n24), .B(n18), .Y(ab_0__3_) );
  XOR2X2 U3 ( .A(ab_1__5_), .B(ab_0__6_), .Y(SUMB_1__5_) );
  NOR2X4 U4 ( .A(n21), .B(n18), .Y(ab_0__6_) );
  AND2X2 U5 ( .A(A[2]), .B(B[5]), .Y(ab_2__5_) );
  AND2X4 U6 ( .A(ab_0__4_), .B(ab_1__3_), .Y(n5) );
  AND2X1 U7 ( .A(A[1]), .B(B[6]), .Y(ab_1__6_) );
  NAND2XL U8 ( .A(A[1]), .B(B[1]), .Y(n20) );
  INVX4 U9 ( .A(B[3]), .Y(n24) );
  XOR2X1 U10 ( .A(CARRYB_16__4_), .B(SUMB_16__5_), .Y(A1_19_) );
  NOR2X1 U11 ( .A(n16), .B(n18), .Y(ab_0__7_) );
  INVX1 U12 ( .A(n20), .Y(n26) );
  XOR2X1 U13 ( .A(CARRYB_16__3_), .B(SUMB_16__4_), .Y(A1_18_) );
  AND2X2 U15 ( .A(ab_0__5_), .B(ab_1__4_), .Y(n4) );
  AND2X2 U16 ( .A(ab_0__6_), .B(ab_1__5_), .Y(n6) );
  AND2X2 U17 ( .A(ab_0__7_), .B(ab_1__6_), .Y(n7) );
  AND2X2 U18 ( .A(ab_0__3_), .B(ab_1__2_), .Y(n8) );
  INVX1 U19 ( .A(n16), .Y(n17) );
  INVX1 U20 ( .A(B[7]), .Y(n16) );
  AND2X2 U21 ( .A(CARRYB_16__0_), .B(SUMB_16__1_), .Y(n9) );
  AND2X2 U22 ( .A(A[2]), .B(B[4]), .Y(ab_2__4_) );
  AND2X2 U23 ( .A(A[2]), .B(B[0]), .Y(ab_2__0_) );
  AND2X4 U24 ( .A(A[2]), .B(B[1]), .Y(ab_2__1_) );
  XOR2X2 U25 ( .A(CARRYB_16__0_), .B(SUMB_16__1_), .Y(A1_15_) );
  NOR2X2 U26 ( .A(n22), .B(n18), .Y(ab_0__5_) );
  INVX4 U27 ( .A(B[5]), .Y(n22) );
  AND2X2 U28 ( .A(A[3]), .B(B[5]), .Y(ab_3__5_) );
  XOR2X4 U29 ( .A(SUMB_16__2_), .B(CARRYB_16__1_), .Y(A1_16_) );
  AND2X2 U30 ( .A(CARRYB_16__1_), .B(SUMB_16__2_), .Y(n11) );
  INVX2 U31 ( .A(B[6]), .Y(n21) );
  AND2X1 U32 ( .A(A[3]), .B(B[1]), .Y(ab_3__1_) );
  INVX2 U33 ( .A(n15), .Y(CARRYB_1__1_) );
  NAND2X1 U34 ( .A(ab_0__2_), .B(n26), .Y(n15) );
  AND2X2 U35 ( .A(A[1]), .B(B[2]), .Y(ab_1__2_) );
  XOR2X1 U36 ( .A(ab_1__6_), .B(ab_0__7_), .Y(SUMB_1__6_) );
  NOR2X1 U37 ( .A(n25), .B(n18), .Y(ab_0__2_) );
  NOR2XL U38 ( .A(n27), .B(n23), .Y(ab_16__4_) );
  AND2X1 U39 ( .A(A[5]), .B(B[0]), .Y(ab_5__0_) );
  AND2X1 U40 ( .A(A[4]), .B(B[0]), .Y(ab_4__0_) );
  INVXL U41 ( .A(A[0]), .Y(n18) );
  AND2X1 U42 ( .A(A[6]), .B(B[0]), .Y(ab_6__0_) );
  AND2X1 U43 ( .A(A[7]), .B(B[0]), .Y(ab_7__0_) );
  AND2X1 U44 ( .A(A[4]), .B(B[1]), .Y(ab_4__1_) );
  AND2X1 U45 ( .A(A[8]), .B(B[0]), .Y(ab_8__0_) );
  AND2X1 U46 ( .A(A[10]), .B(B[1]), .Y(ab_10__1_) );
  AND2X1 U47 ( .A(A[9]), .B(B[1]), .Y(ab_9__1_) );
  AND2X1 U48 ( .A(A[8]), .B(B[1]), .Y(ab_8__1_) );
  AND2X1 U49 ( .A(A[10]), .B(B[0]), .Y(ab_10__0_) );
  AND2X1 U50 ( .A(A[9]), .B(B[0]), .Y(ab_9__0_) );
  AND2X1 U51 ( .A(A[7]), .B(B[1]), .Y(ab_7__1_) );
  AND2X1 U52 ( .A(A[6]), .B(B[1]), .Y(ab_6__1_) );
  INVXL U53 ( .A(B[0]), .Y(n34) );
  AND2X1 U54 ( .A(CARRYB_16__2_), .B(SUMB_16__3_), .Y(n10) );
  NOR2XL U55 ( .A(n27), .B(n24), .Y(ab_16__3_) );
  XOR2X1 U56 ( .A(CARRYB_16__5_), .B(SUMB_16__6_), .Y(A1_20_) );
  XOR2X1 U57 ( .A(CARRYB_16__6_), .B(ab_16__7_), .Y(A1_21_) );
  AND2X1 U58 ( .A(CARRYB_16__3_), .B(SUMB_16__4_), .Y(n12) );
  AND2X1 U59 ( .A(CARRYB_16__4_), .B(SUMB_16__5_), .Y(n13) );
  AND2X2 U60 ( .A(CARRYB_16__5_), .B(SUMB_16__6_), .Y(n14) );
  NOR2X1 U61 ( .A(n27), .B(n16), .Y(ab_16__7_) );
  NOR2X1 U62 ( .A(n23), .B(n18), .Y(ab_0__4_) );
  NOR2XL U63 ( .A(n28), .B(n24), .Y(ab_15__3_) );
  NOR2XL U64 ( .A(n29), .B(n24), .Y(ab_14__3_) );
  NOR2XL U65 ( .A(n28), .B(n16), .Y(ab_15__7_) );
  AND2X1 U66 ( .A(A[10]), .B(B[3]), .Y(ab_10__3_) );
  AND2X1 U67 ( .A(A[9]), .B(B[3]), .Y(ab_9__3_) );
  AND2X1 U68 ( .A(A[8]), .B(B[3]), .Y(ab_8__3_) );
  AND2X1 U69 ( .A(A[7]), .B(B[3]), .Y(ab_7__3_) );
  AND2X1 U70 ( .A(A[6]), .B(B[3]), .Y(ab_6__3_) );
  NOR2XL U71 ( .A(n32), .B(n16), .Y(ab_11__7_) );
  XOR2X1 U72 ( .A(ab_1__4_), .B(ab_0__5_), .Y(SUMB_1__4_) );
  XOR2X1 U73 ( .A(ab_1__3_), .B(ab_0__4_), .Y(SUMB_1__3_) );
  NOR2XL U74 ( .A(n31), .B(n16), .Y(ab_12__7_) );
  NOR2XL U75 ( .A(n29), .B(n16), .Y(ab_14__7_) );
  NOR2XL U76 ( .A(n30), .B(n16), .Y(ab_13__7_) );
  INVX1 U77 ( .A(A[16]), .Y(n27) );
  NAND2XL U78 ( .A(A[0]), .B(B[0]), .Y(n19) );
  AND2X1 U79 ( .A(A[3]), .B(B[4]), .Y(ab_3__4_) );
  INVX1 U80 ( .A(A[13]), .Y(n30) );
  AND2X1 U81 ( .A(A[4]), .B(B[4]), .Y(ab_4__4_) );
  AND2X1 U82 ( .A(A[3]), .B(B[0]), .Y(ab_3__0_) );
  XOR2X1 U83 ( .A(n26), .B(ab_0__2_), .Y(SUMB_1__1_) );
  AND2X1 U84 ( .A(A[9]), .B(B[4]), .Y(ab_9__4_) );
  AND2X1 U85 ( .A(A[10]), .B(B[4]), .Y(ab_10__4_) );
  AND2X1 U86 ( .A(A[8]), .B(B[4]), .Y(ab_8__4_) );
  AND2X1 U87 ( .A(A[7]), .B(B[4]), .Y(ab_7__4_) );
  AND2X1 U88 ( .A(A[6]), .B(B[4]), .Y(ab_6__4_) );
  AND2X1 U89 ( .A(A[5]), .B(B[4]), .Y(ab_5__4_) );
  AND2X1 U90 ( .A(A[8]), .B(B[6]), .Y(ab_8__6_) );
  AND2X1 U91 ( .A(A[7]), .B(B[6]), .Y(ab_7__6_) );
  AND2X1 U92 ( .A(A[9]), .B(B[6]), .Y(ab_9__6_) );
  AND2X1 U93 ( .A(A[6]), .B(B[6]), .Y(ab_6__6_) );
  AND2X1 U94 ( .A(A[5]), .B(B[6]), .Y(ab_5__6_) );
  AND2X1 U95 ( .A(A[3]), .B(n17), .Y(ab_3__7_) );
  AND2X1 U96 ( .A(A[4]), .B(B[6]), .Y(ab_4__6_) );
  AND2X1 U97 ( .A(A[5]), .B(B[1]), .Y(ab_5__1_) );
  AND2X1 U98 ( .A(A[2]), .B(n17), .Y(ab_2__7_) );
  AND2X1 U99 ( .A(A[3]), .B(B[6]), .Y(ab_3__6_) );
  AND2X1 U100 ( .A(A[2]), .B(B[6]), .Y(ab_2__6_) );
  XOR2X1 U101 ( .A(ab_1__2_), .B(ab_0__3_), .Y(SUMB_1__2_) );
  INVX4 U102 ( .A(B[4]), .Y(n23) );
  INVX1 U103 ( .A(A[11]), .Y(n32) );
  AND2X1 U104 ( .A(A[10]), .B(B[6]), .Y(ab_10__6_) );
  INVX1 U105 ( .A(A[14]), .Y(n29) );
  INVX1 U106 ( .A(A[15]), .Y(n28) );
  INVX1 U107 ( .A(A[12]), .Y(n31) );
  INVX1 U108 ( .A(B[1]), .Y(n33) );
  XOR2X4 U109 ( .A(CARRYB_16__2_), .B(SUMB_16__3_), .Y(A1_17_) );
  NOR2XL U110 ( .A(n32), .B(n23), .Y(ab_11__4_) );
  NOR2XL U111 ( .A(n31), .B(n23), .Y(ab_12__4_) );
  NOR2XL U112 ( .A(n30), .B(n23), .Y(ab_13__4_) );
  NOR2XL U113 ( .A(n29), .B(n23), .Y(ab_14__4_) );
  NOR2XL U114 ( .A(n28), .B(n23), .Y(ab_15__4_) );
  NOR2XL U115 ( .A(n27), .B(n21), .Y(ab_16__6_) );
  NOR2XL U116 ( .A(n28), .B(n21), .Y(ab_15__6_) );
  NOR2XL U117 ( .A(n29), .B(n21), .Y(ab_14__6_) );
  NOR2XL U118 ( .A(n30), .B(n21), .Y(ab_13__6_) );
  NOR2XL U119 ( .A(n31), .B(n21), .Y(ab_12__6_) );
  NOR2XL U120 ( .A(n32), .B(n21), .Y(ab_11__6_) );
  AND2X1 U121 ( .A(A[10]), .B(B[5]), .Y(ab_10__5_) );
  AND2X1 U122 ( .A(A[9]), .B(B[5]), .Y(ab_9__5_) );
  AND2X1 U123 ( .A(A[8]), .B(B[5]), .Y(ab_8__5_) );
  AND2X1 U124 ( .A(A[7]), .B(B[5]), .Y(ab_7__5_) );
  AND2X1 U125 ( .A(A[6]), .B(B[5]), .Y(ab_6__5_) );
  AND2X1 U126 ( .A(A[5]), .B(B[5]), .Y(ab_5__5_) );
  AND2X1 U127 ( .A(A[4]), .B(B[5]), .Y(ab_4__5_) );
  NOR2XL U128 ( .A(n27), .B(n25), .Y(ab_16__2_) );
  NOR2XL U129 ( .A(n28), .B(n25), .Y(ab_15__2_) );
  NOR2XL U130 ( .A(n29), .B(n25), .Y(ab_14__2_) );
  NOR2XL U131 ( .A(n30), .B(n25), .Y(ab_13__2_) );
  NOR2XL U132 ( .A(n31), .B(n25), .Y(ab_12__2_) );
  NOR2XL U133 ( .A(n32), .B(n25), .Y(ab_11__2_) );
  AND2X1 U134 ( .A(A[10]), .B(B[2]), .Y(ab_10__2_) );
  AND2X1 U135 ( .A(A[9]), .B(B[2]), .Y(ab_9__2_) );
  AND2X1 U136 ( .A(A[8]), .B(B[2]), .Y(ab_8__2_) );
  AND2X1 U137 ( .A(A[7]), .B(B[2]), .Y(ab_7__2_) );
  AND2X1 U138 ( .A(A[6]), .B(B[2]), .Y(ab_6__2_) );
  AND2X1 U139 ( .A(A[5]), .B(B[2]), .Y(ab_5__2_) );
  AND2X2 U140 ( .A(A[4]), .B(B[2]), .Y(ab_4__2_) );
  AND2X2 U141 ( .A(A[3]), .B(B[2]), .Y(ab_3__2_) );
  AND2X2 U142 ( .A(A[2]), .B(B[2]), .Y(ab_2__2_) );
  INVX4 U143 ( .A(B[2]), .Y(n25) );
  AND2X2 U144 ( .A(A[2]), .B(B[3]), .Y(ab_2__3_) );
  AND2X2 U145 ( .A(A[3]), .B(B[3]), .Y(ab_3__3_) );
  AND2X2 U146 ( .A(A[4]), .B(B[3]), .Y(ab_4__3_) );
  AND2X2 U147 ( .A(A[5]), .B(B[3]), .Y(ab_5__3_) );
  NOR2X1 U148 ( .A(n32), .B(n24), .Y(ab_11__3_) );
  NOR2X1 U149 ( .A(n31), .B(n24), .Y(ab_12__3_) );
  NOR2X1 U150 ( .A(n30), .B(n24), .Y(ab_13__3_) );
  NOR2XL U151 ( .A(n27), .B(n22), .Y(ab_16__5_) );
  NOR2XL U152 ( .A(n28), .B(n22), .Y(ab_15__5_) );
  NOR2XL U153 ( .A(n29), .B(n22), .Y(ab_14__5_) );
  NOR2XL U154 ( .A(n30), .B(n22), .Y(ab_13__5_) );
  NOR2XL U155 ( .A(n31), .B(n22), .Y(ab_12__5_) );
  NOR2XL U156 ( .A(n32), .B(n22), .Y(ab_11__5_) );
  AND2X2 U157 ( .A(A[1]), .B(B[5]), .Y(ab_1__5_) );
  AND2X1 U158 ( .A(A[1]), .B(n17), .Y(ab_1__7_) );
  NOR2XL U159 ( .A(n20), .B(n19), .Y(CARRYB_1__0_) );
  AND2X2 U160 ( .A(A[1]), .B(B[4]), .Y(ab_1__4_) );
  AND2X2 U161 ( .A(A[1]), .B(B[3]), .Y(ab_1__3_) );
  AND2X1 U162 ( .A(A[10]), .B(n17), .Y(ab_10__7_) );
  AND2X1 U163 ( .A(A[9]), .B(n17), .Y(ab_9__7_) );
  AND2X1 U164 ( .A(A[8]), .B(n17), .Y(ab_8__7_) );
  AND2X1 U165 ( .A(A[7]), .B(n17), .Y(ab_7__7_) );
  AND2X1 U166 ( .A(A[6]), .B(n17), .Y(ab_6__7_) );
  AND2X1 U167 ( .A(A[5]), .B(n17), .Y(ab_5__7_) );
  AND2X1 U168 ( .A(A[4]), .B(n17), .Y(ab_4__7_) );
  NOR2X1 U170 ( .A(n33), .B(n27), .Y(ab_16__1_) );
  NOR2X1 U171 ( .A(n34), .B(n27), .Y(ab_16__0_) );
  NOR2X1 U172 ( .A(n33), .B(n28), .Y(ab_15__1_) );
  NOR2X1 U173 ( .A(n34), .B(n28), .Y(ab_15__0_) );
  NOR2X1 U174 ( .A(n33), .B(n29), .Y(ab_14__1_) );
  NOR2X1 U175 ( .A(n34), .B(n29), .Y(ab_14__0_) );
  NOR2X1 U176 ( .A(n33), .B(n30), .Y(ab_13__1_) );
  NOR2X1 U177 ( .A(n34), .B(n30), .Y(ab_13__0_) );
  NOR2X1 U178 ( .A(n33), .B(n31), .Y(ab_12__1_) );
  NOR2X1 U179 ( .A(n34), .B(n31), .Y(ab_12__0_) );
  NOR2X1 U180 ( .A(n33), .B(n32), .Y(ab_11__1_) );
  NOR2X1 U181 ( .A(n34), .B(n32), .Y(ab_11__0_) );
endmodule


module multi16_8 ( in_17bit, in_8bit, out );
  input [16:0] in_17bit;
  input [7:0] in_8bit;
  output [16:0] out;
  wire   N18, N19, N20, N21, N32, N33, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n55, n56, n57, n58, n59, n60, n61, n63, n64, n65, n66, n67, n68,
         n69, n71, n72, n73, n74, n75, n76, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n116, n117, n118, n119;
  wire   [16:1] in_17bit_b;
  wire   [7:0] in_8bit_b;
  wire   [23:8] mul;
  wire   [16:12] sub_add_52_b0_carry;

  multi16_8_DW02_mult_0 mult_55 ( .A({in_17bit_b, in_17bit[0]}), .B(in_8bit_b), 
        .PRODUCT_23_(mul[23]), .PRODUCT_22_(mul[22]), .PRODUCT_21_(mul[21]), 
        .PRODUCT_20_(mul[20]), .PRODUCT_19_(mul[19]), .PRODUCT_18_(mul[18]), 
        .PRODUCT_17_(mul[17]), .PRODUCT_16_(mul[16]), .PRODUCT_15_(mul[15]), 
        .PRODUCT_14_(mul[14]), .PRODUCT_13_(mul[13]), .PRODUCT_12_(mul[12]), 
        .PRODUCT_11_(mul[11]), .PRODUCT_10_(mul[10]), .PRODUCT_9_(mul[9]), 
        .PRODUCT_8_(mul[8]), .PRODUCT_7_(N32) );
  NOR2X2 U2 ( .A(n20), .B(n39), .Y(n38) );
  OAI22X1 U3 ( .A0(in_17bit[1]), .A1(in_17bit[0]), .B0(in_17bit[16]), .B1(
        in_17bit[1]), .Y(n35) );
  CLKINVX2 U4 ( .A(in_17bit[16]), .Y(n19) );
  NAND2XL U5 ( .A(n105), .B(n104), .Y(n1) );
  CLKINVX3 U6 ( .A(n8), .Y(n2) );
  AND2X4 U7 ( .A(n1), .B(n2), .Y(n106) );
  INVX3 U8 ( .A(mul[22]), .Y(n104) );
  XOR2X2 U9 ( .A(mul[23]), .B(n106), .Y(out[16]) );
  NOR2X4 U10 ( .A(mul[20]), .B(n10), .Y(n9) );
  NAND2BX1 U11 ( .AN(in_8bit[2]), .B(n25), .Y(n29) );
  CLKINVX4 U12 ( .A(in_8bit[3]), .Y(n25) );
  XOR2X1 U13 ( .A(mul[19]), .B(n98), .Y(out[12]) );
  XOR2X1 U14 ( .A(n101), .B(mul[21]), .Y(out[14]) );
  OR2X2 U15 ( .A(n114), .B(n31), .Y(n13) );
  INVX2 U16 ( .A(n102), .Y(n105) );
  NAND2BX1 U17 ( .AN(mul[21]), .B(n9), .Y(n102) );
  NOR2BX2 U18 ( .AN(n36), .B(n35), .Y(in_17bit_b[1]) );
  XOR2X1 U19 ( .A(mul[16]), .B(n91), .Y(out[9]) );
  AOI21X2 U20 ( .A0(n14), .A1(n18), .B0(n114), .Y(n24) );
  NOR2X2 U21 ( .A(mul[13]), .B(n83), .Y(n5) );
  NOR2X1 U22 ( .A(n8), .B(n89), .Y(n88) );
  INVX2 U23 ( .A(n93), .Y(n95) );
  NOR2X2 U24 ( .A(n8), .B(n9), .Y(n101) );
  INVX1 U25 ( .A(n37), .Y(n39) );
  AND2X2 U26 ( .A(n15), .B(n22), .Y(n14) );
  INVX1 U27 ( .A(in_8bit[1]), .Y(n22) );
  INVX1 U28 ( .A(n87), .Y(n89) );
  NAND2BX1 U29 ( .AN(mul[14]), .B(n5), .Y(n87) );
  CLKINVX3 U30 ( .A(n90), .Y(n92) );
  NAND2BX2 U31 ( .AN(mul[15]), .B(n89), .Y(n90) );
  NOR2X1 U32 ( .A(n8), .B(n5), .Y(n86) );
  INVX1 U33 ( .A(n116), .Y(in_8bit_b[0]) );
  XNOR2X1 U34 ( .A(n48), .B(n6), .Y(in_17bit_b[6]) );
  INVX1 U35 ( .A(n83), .Y(n85) );
  NAND2BX1 U36 ( .AN(mul[12]), .B(n82), .Y(n83) );
  NAND2X1 U37 ( .A(n31), .B(n30), .Y(n34) );
  XOR2X2 U38 ( .A(mul[17]), .B(n94), .Y(out[10]) );
  INVX4 U39 ( .A(n97), .Y(n99) );
  NAND2BX4 U40 ( .AN(mul[18]), .B(n4), .Y(n97) );
  NOR2X4 U41 ( .A(n8), .B(n4), .Y(n96) );
  NAND2BXL U42 ( .AN(in_17bit[2]), .B(n16), .Y(n37) );
  NOR3XL U43 ( .A(in_8bit[6]), .B(n114), .C(n34), .Y(in_8bit_b[7]) );
  XOR2X4 U44 ( .A(in_17bit[2]), .B(n3), .Y(in_17bit_b[2]) );
  NOR2X4 U45 ( .A(n19), .B(n16), .Y(n3) );
  XOR2X2 U46 ( .A(mul[18]), .B(n96), .Y(out[11]) );
  INVX2 U47 ( .A(n11), .Y(n10) );
  NOR2X4 U48 ( .A(mul[17]), .B(n93), .Y(n4) );
  NOR2X4 U49 ( .A(n8), .B(n99), .Y(n98) );
  NOR2X4 U50 ( .A(in_17bit[1]), .B(in_17bit[0]), .Y(n16) );
  NOR2X4 U51 ( .A(n8), .B(n105), .Y(n103) );
  XOR2X4 U52 ( .A(n38), .B(in_17bit[3]), .Y(in_17bit_b[3]) );
  NAND2X2 U53 ( .A(n34), .B(in_8bit[7]), .Y(n33) );
  NOR2X4 U54 ( .A(mul[19]), .B(n12), .Y(n11) );
  INVX2 U55 ( .A(n99), .Y(n12) );
  NOR2X4 U56 ( .A(n8), .B(n11), .Y(n100) );
  NAND3XL U57 ( .A(in_17bit[0]), .B(in_17bit[16]), .C(in_17bit[1]), .Y(n36) );
  NOR4X1 U58 ( .A(in_8bit[0]), .B(in_8bit[4]), .C(in_8bit[1]), .D(n29), .Y(n31) );
  NOR2X2 U59 ( .A(n8), .B(n92), .Y(n91) );
  INVXL U60 ( .A(in_8bit[2]), .Y(n18) );
  NAND2BX4 U61 ( .AN(mul[16]), .B(n92), .Y(n93) );
  XOR2X4 U62 ( .A(n13), .B(n30), .Y(in_8bit_b[5]) );
  NAND2BXL U63 ( .AN(mul[8]), .B(n108), .Y(n69) );
  XNOR2X2 U64 ( .A(n44), .B(n45), .Y(in_17bit_b[5]) );
  NOR2X2 U65 ( .A(n20), .B(n46), .Y(n44) );
  AND2X1 U66 ( .A(n47), .B(n17), .Y(n6) );
  NAND2XL U67 ( .A(n46), .B(n45), .Y(n47) );
  NAND2XL U68 ( .A(n52), .B(n51), .Y(n55) );
  XOR2X2 U69 ( .A(n42), .B(n40), .Y(in_17bit_b[4]) );
  NAND2BXL U70 ( .AN(n41), .B(n42), .Y(n43) );
  NAND2BXL U71 ( .AN(n47), .B(n48), .Y(n49) );
  NOR2XL U72 ( .A(n19), .B(n60), .Y(n58) );
  INVXL U73 ( .A(n66), .Y(n67) );
  INVXL U74 ( .A(n68), .Y(sub_add_52_b0_carry[12]) );
  AND2X2 U75 ( .A(sub_add_52_b0_carry[13]), .B(n111), .Y(
        sub_add_52_b0_carry[14]) );
  NAND2XL U76 ( .A(n60), .B(n59), .Y(n63) );
  NAND2BXL U77 ( .AN(n55), .B(n56), .Y(n57) );
  XOR2XL U78 ( .A(n111), .B(sub_add_52_b0_carry[13]), .Y(N18) );
  AND2X1 U79 ( .A(N21), .B(n17), .Y(in_17bit_b[16]) );
  INVXL U80 ( .A(in_17bit[16]), .Y(n20) );
  XOR2X1 U81 ( .A(mul[14]), .B(n86), .Y(out[7]) );
  INVXL U82 ( .A(in_17bit[5]), .Y(n45) );
  NOR2X2 U83 ( .A(n114), .B(n14), .Y(n23) );
  INVXL U84 ( .A(in_17bit[4]), .Y(n42) );
  INVXL U85 ( .A(in_8bit[0]), .Y(n15) );
  MX2X1 U86 ( .A(in_17bit[12]), .B(n7), .S0(n17), .Y(in_17bit_b[12]) );
  XNOR2X1 U87 ( .A(n68), .B(n110), .Y(n7) );
  MX2X1 U88 ( .A(in_17bit[13]), .B(N18), .S0(n17), .Y(in_17bit_b[13]) );
  MX2X1 U89 ( .A(in_17bit[14]), .B(N19), .S0(n17), .Y(in_17bit_b[14]) );
  MX2X1 U90 ( .A(in_17bit[15]), .B(N20), .S0(n17), .Y(in_17bit_b[15]) );
  INVXL U91 ( .A(in_17bit[7]), .Y(n51) );
  INVXL U92 ( .A(in_17bit[9]), .Y(n59) );
  INVXL U93 ( .A(in_17bit[6]), .Y(n48) );
  INVXL U94 ( .A(in_17bit[8]), .Y(n56) );
  XOR2X1 U95 ( .A(n22), .B(n21), .Y(in_8bit_b[1]) );
  XNOR2X1 U96 ( .A(n17), .B(in_8bit[7]), .Y(n8) );
  INVX1 U97 ( .A(n80), .Y(n82) );
  NAND2BX1 U98 ( .AN(mul[11]), .B(n79), .Y(n80) );
  INVX1 U99 ( .A(n76), .Y(n79) );
  NAND2BX1 U100 ( .AN(mul[10]), .B(n75), .Y(n76) );
  INVX1 U101 ( .A(n73), .Y(n75) );
  NAND2BX1 U102 ( .AN(mul[9]), .B(n72), .Y(n73) );
  INVX1 U103 ( .A(n69), .Y(n72) );
  INVX1 U104 ( .A(N32), .Y(n108) );
  XNOR2X1 U105 ( .A(n50), .B(n51), .Y(in_17bit_b[7]) );
  NOR2X1 U106 ( .A(n20), .B(n52), .Y(n50) );
  XOR2X1 U107 ( .A(n56), .B(n53), .Y(in_17bit_b[8]) );
  NAND2X1 U108 ( .A(n55), .B(n17), .Y(n53) );
  XOR2X1 U109 ( .A(n64), .B(n61), .Y(in_17bit_b[10]) );
  NAND2X1 U110 ( .A(n63), .B(n17), .Y(n61) );
  NAND2BX1 U111 ( .AN(n63), .B(n64), .Y(n66) );
  XNOR2X1 U112 ( .A(n58), .B(n59), .Y(in_17bit_b[9]) );
  INVX1 U113 ( .A(n43), .Y(n46) );
  INVX1 U114 ( .A(n49), .Y(n52) );
  INVX1 U115 ( .A(n57), .Y(n60) );
  NAND2X1 U116 ( .A(n109), .B(n67), .Y(n68) );
  INVXL U117 ( .A(in_8bit[5]), .Y(n30) );
  XOR2X1 U118 ( .A(mul[15]), .B(n88), .Y(out[8]) );
  XOR2X1 U119 ( .A(mul[11]), .B(n78), .Y(out[4]) );
  NOR2X1 U120 ( .A(n8), .B(n79), .Y(n78) );
  XOR2X1 U121 ( .A(mul[9]), .B(n71), .Y(out[2]) );
  NOR2X1 U122 ( .A(n8), .B(n72), .Y(n71) );
  XOR2X1 U123 ( .A(mul[12]), .B(n81), .Y(out[5]) );
  NOR2X1 U124 ( .A(n8), .B(n82), .Y(n81) );
  XOR2X1 U125 ( .A(mul[10]), .B(n74), .Y(out[3]) );
  NOR2X1 U126 ( .A(n8), .B(n75), .Y(n74) );
  XOR2X1 U127 ( .A(mul[13]), .B(n84), .Y(out[6]) );
  NOR2X1 U128 ( .A(n8), .B(n85), .Y(n84) );
  NAND2BXL U129 ( .AN(in_17bit[3]), .B(n39), .Y(n41) );
  INVX1 U130 ( .A(n118), .Y(out[1]) );
  AOI22XL U131 ( .A0(mul[8]), .A1(n8), .B0(N33), .B1(n119), .Y(n118) );
  INVX1 U132 ( .A(mul[8]), .Y(n107) );
  MXI2X1 U133 ( .A(n109), .B(n65), .S0(n17), .Y(in_17bit_b[11]) );
  XOR2X1 U134 ( .A(n66), .B(n109), .Y(n65) );
  INVX1 U135 ( .A(n117), .Y(out[0]) );
  AOI22XL U136 ( .A0(N32), .A1(n8), .B0(N32), .B1(n119), .Y(n117) );
  INVXL U137 ( .A(n8), .Y(n119) );
  INVX1 U138 ( .A(in_17bit[10]), .Y(n64) );
  INVX1 U139 ( .A(in_17bit[11]), .Y(n109) );
  INVX1 U140 ( .A(in_17bit[12]), .Y(n110) );
  INVX1 U141 ( .A(in_17bit[13]), .Y(n111) );
  INVX1 U142 ( .A(in_17bit[14]), .Y(n112) );
  INVX1 U143 ( .A(in_17bit[15]), .Y(n113) );
  INVXL U144 ( .A(n29), .Y(n26) );
  INVXL U145 ( .A(in_8bit[6]), .Y(n32) );
  INVX1 U146 ( .A(in_8bit[7]), .Y(n114) );
  AOI21X2 U147 ( .A0(n27), .A1(n26), .B0(n114), .Y(n28) );
  INVXL U148 ( .A(n20), .Y(n17) );
  NAND2X1 U149 ( .A(n41), .B(in_17bit[16]), .Y(n40) );
  AOI22XL U150 ( .A0(in_8bit[0]), .A1(in_8bit[7]), .B0(in_8bit[0]), .B1(n114), 
        .Y(n116) );
  NAND2XL U151 ( .A(in_8bit[0]), .B(in_8bit[7]), .Y(n21) );
  NOR2XL U152 ( .A(in_8bit[1]), .B(in_8bit[0]), .Y(n27) );
  XNOR2X4 U153 ( .A(n23), .B(n18), .Y(in_8bit_b[2]) );
  XNOR2X4 U154 ( .A(n24), .B(n25), .Y(in_8bit_b[3]) );
  XOR2X4 U155 ( .A(n28), .B(in_8bit[4]), .Y(in_8bit_b[4]) );
  XOR2X4 U156 ( .A(n33), .B(n32), .Y(in_8bit_b[6]) );
  NOR2X4 U157 ( .A(n8), .B(n95), .Y(n94) );
  XOR2X4 U158 ( .A(mul[20]), .B(n100), .Y(out[13]) );
  XNOR2X4 U159 ( .A(n103), .B(n104), .Y(out[15]) );
  XOR2X1 U160 ( .A(n107), .B(n108), .Y(N33) );
  XOR2X1 U161 ( .A(n19), .B(sub_add_52_b0_carry[16]), .Y(N21) );
  AND2X1 U162 ( .A(sub_add_52_b0_carry[15]), .B(n113), .Y(
        sub_add_52_b0_carry[16]) );
  XOR2X1 U163 ( .A(n113), .B(sub_add_52_b0_carry[15]), .Y(N20) );
  AND2X1 U164 ( .A(sub_add_52_b0_carry[14]), .B(n112), .Y(
        sub_add_52_b0_carry[15]) );
  XOR2X1 U165 ( .A(n112), .B(sub_add_52_b0_carry[14]), .Y(N19) );
  AND2X1 U166 ( .A(sub_add_52_b0_carry[12]), .B(n110), .Y(
        sub_add_52_b0_carry[13]) );
endmodule


module multi16_7_DW01_add_0 ( A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, 
        A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, 
        B_20_, B_19_, B_18_, B_17_, B_16_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, 
        SUM_17_, SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, 
        SUM_9_, SUM_8_, SUM_7_, SUM_6_, SUM_5_ );
  input A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_,
         A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, B_20_, B_19_,
         B_18_, B_17_, B_16_;
  output SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, SUM_15_,
         SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, SUM_7_,
         SUM_6_, SUM_5_;
  wire   n1, n2, n4, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41;

  NOR2X1 U2 ( .A(B_19_), .B(A_19_), .Y(n29) );
  NOR2X1 U3 ( .A(n28), .B(n29), .Y(n1) );
  INVXL U4 ( .A(n30), .Y(n2) );
  OR2X4 U5 ( .A(n1), .B(n2), .Y(n24) );
  AOI21X1 U6 ( .A0(n16), .A1(n33), .B0(n17), .Y(n28) );
  AOI21XL U7 ( .A0(n24), .A1(n25), .B0(n15), .Y(n23) );
  XNOR2X2 U8 ( .A(n27), .B(n24), .Y(SUM_20_) );
  NOR2X4 U9 ( .A(B_17_), .B(A_17_), .Y(n31) );
  BUFX3 U10 ( .A(A_14_), .Y(SUM_14_) );
  BUFX3 U11 ( .A(A_11_), .Y(SUM_11_) );
  NAND2X1 U12 ( .A(n34), .B(n16), .Y(n40) );
  INVX2 U13 ( .A(n31), .Y(n19) );
  INVX4 U14 ( .A(n36), .Y(n18) );
  XOR2X4 U15 ( .A(n40), .B(n39), .Y(SUM_18_) );
  CLKINVX3 U16 ( .A(n35), .Y(n20) );
  NAND2X1 U17 ( .A(B_18_), .B(A_18_), .Y(n34) );
  NOR2BX2 U18 ( .AN(n30), .B(n29), .Y(n38) );
  NOR2X4 U19 ( .A(n31), .B(n18), .Y(n41) );
  XOR2X4 U20 ( .A(n37), .B(n38), .Y(SUM_19_) );
  OAI21X2 U21 ( .A0(n39), .A1(n32), .B0(n34), .Y(n37) );
  AOI21X4 U22 ( .A0(n20), .A1(n19), .B0(n18), .Y(n39) );
  NOR2X2 U23 ( .A(B_18_), .B(A_18_), .Y(n32) );
  INVX2 U24 ( .A(n32), .Y(n16) );
  NAND2X2 U25 ( .A(B_17_), .B(A_17_), .Y(n36) );
  INVX4 U26 ( .A(n21), .Y(SUM_15_) );
  NAND2X2 U27 ( .A(B_16_), .B(A_16_), .Y(n35) );
  NOR2BX2 U28 ( .AN(n35), .B(n4), .Y(SUM_16_) );
  XOR2X2 U29 ( .A(n20), .B(n41), .Y(SUM_17_) );
  INVX2 U30 ( .A(A_15_), .Y(n21) );
  INVXL U31 ( .A(n34), .Y(n17) );
  NOR2XL U32 ( .A(B_16_), .B(A_16_), .Y(n4) );
  INVXL U33 ( .A(n26), .Y(n15) );
  BUFX3 U34 ( .A(A_12_), .Y(SUM_12_) );
  BUFX3 U35 ( .A(A_5_), .Y(SUM_5_) );
  BUFX3 U36 ( .A(A_9_), .Y(SUM_9_) );
  BUFX3 U37 ( .A(A_6_), .Y(SUM_6_) );
  BUFX3 U38 ( .A(A_7_), .Y(SUM_7_) );
  BUFX3 U39 ( .A(A_8_), .Y(SUM_8_) );
  BUFX4 U40 ( .A(A_13_), .Y(SUM_13_) );
  BUFX3 U41 ( .A(A_10_), .Y(SUM_10_) );
  XOR2X1 U42 ( .A(n22), .B(n23), .Y(SUM_21_) );
  XNOR2X1 U43 ( .A(B_21_), .B(A_21_), .Y(n22) );
  OAI21XL U44 ( .A0(n31), .A1(n35), .B0(n36), .Y(n33) );
  NAND2X1 U45 ( .A(n26), .B(n25), .Y(n27) );
  OR2X1 U46 ( .A(B_20_), .B(A_20_), .Y(n25) );
  NAND2X1 U47 ( .A(B_20_), .B(A_20_), .Y(n26) );
  NAND2X1 U48 ( .A(B_19_), .B(A_19_), .Y(n30) );
endmodule


module multi16_7_DW02_mult_0 ( A, B, PRODUCT_23_, PRODUCT_22_, PRODUCT_21_, 
        PRODUCT_20_, PRODUCT_19_, PRODUCT_18_, PRODUCT_17_, PRODUCT_16_, 
        PRODUCT_15_, PRODUCT_14_, PRODUCT_13_, PRODUCT_12_, PRODUCT_11_, 
        PRODUCT_10_, PRODUCT_9_, PRODUCT_8_, PRODUCT_7_ );
  input [16:0] A;
  input [7:0] B;
  output PRODUCT_23_, PRODUCT_22_, PRODUCT_21_, PRODUCT_20_, PRODUCT_19_,
         PRODUCT_18_, PRODUCT_17_, PRODUCT_16_, PRODUCT_15_, PRODUCT_14_,
         PRODUCT_13_, PRODUCT_12_, PRODUCT_11_, PRODUCT_10_, PRODUCT_9_,
         PRODUCT_8_, PRODUCT_7_;
  wire   ab_16__7_, ab_16__6_, ab_16__5_, ab_16__4_, ab_16__3_, ab_16__2_,
         ab_16__1_, ab_16__0_, ab_15__7_, ab_15__6_, ab_15__5_, ab_15__4_,
         ab_15__3_, ab_15__2_, ab_15__1_, ab_15__0_, ab_14__7_, ab_14__6_,
         ab_14__5_, ab_14__4_, ab_14__3_, ab_14__2_, ab_14__1_, ab_14__0_,
         ab_13__7_, ab_13__6_, ab_13__5_, ab_13__4_, ab_13__3_, ab_13__2_,
         ab_13__1_, ab_13__0_, ab_12__7_, ab_12__6_, ab_12__5_, ab_12__4_,
         ab_12__3_, ab_12__2_, ab_12__1_, ab_12__0_, ab_11__7_, ab_11__6_,
         ab_11__5_, ab_11__4_, ab_11__3_, ab_11__2_, ab_11__1_, ab_11__0_,
         ab_10__7_, ab_10__6_, ab_10__5_, ab_10__4_, ab_10__3_, ab_10__2_,
         ab_10__1_, ab_10__0_, ab_9__7_, ab_9__6_, ab_9__5_, ab_9__4_,
         ab_9__3_, ab_9__2_, ab_9__1_, ab_9__0_, ab_8__7_, ab_8__6_, ab_8__5_,
         ab_8__4_, ab_8__3_, ab_8__2_, ab_8__1_, ab_8__0_, ab_7__7_, ab_7__6_,
         ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_, ab_7__0_, ab_6__7_,
         ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_, ab_6__1_, ab_6__0_,
         ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_, ab_5__2_, ab_5__1_,
         ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_, ab_4__3_, ab_4__2_,
         ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_, ab_3__4_, ab_3__3_,
         ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_, ab_2__5_, ab_2__4_,
         ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_, ab_1__6_, ab_1__5_,
         ab_1__4_, ab_1__3_, ab_1__2_, ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_,
         ab_0__3_, ab_0__2_, CARRYB_16__6_, CARRYB_16__5_, CARRYB_16__4_,
         CARRYB_16__3_, CARRYB_16__2_, CARRYB_16__1_, CARRYB_16__0_,
         CARRYB_15__6_, CARRYB_15__5_, CARRYB_15__4_, CARRYB_15__3_,
         CARRYB_15__2_, CARRYB_15__1_, CARRYB_15__0_, CARRYB_14__6_,
         CARRYB_14__5_, CARRYB_14__4_, CARRYB_14__3_, CARRYB_14__2_,
         CARRYB_14__1_, CARRYB_14__0_, CARRYB_13__6_, CARRYB_13__5_,
         CARRYB_13__4_, CARRYB_13__3_, CARRYB_13__2_, CARRYB_13__1_,
         CARRYB_13__0_, CARRYB_12__6_, CARRYB_12__5_, CARRYB_12__4_,
         CARRYB_12__3_, CARRYB_12__2_, CARRYB_12__1_, CARRYB_12__0_,
         CARRYB_11__6_, CARRYB_11__5_, CARRYB_11__4_, CARRYB_11__3_,
         CARRYB_11__2_, CARRYB_11__1_, CARRYB_11__0_, CARRYB_10__6_,
         CARRYB_10__5_, CARRYB_10__4_, CARRYB_10__3_, CARRYB_10__2_,
         CARRYB_10__1_, CARRYB_10__0_, CARRYB_9__6_, CARRYB_9__5_,
         CARRYB_9__4_, CARRYB_9__3_, CARRYB_9__2_, CARRYB_9__1_, CARRYB_9__0_,
         CARRYB_8__6_, CARRYB_8__5_, CARRYB_8__4_, CARRYB_8__3_, CARRYB_8__2_,
         CARRYB_8__1_, CARRYB_8__0_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_,
         CARRYB_7__3_, CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_,
         CARRYB_6__5_, CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_,
         CARRYB_6__0_, CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_,
         CARRYB_5__2_, CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_,
         CARRYB_4__4_, CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_,
         CARRYB_3__6_, CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_,
         CARRYB_3__1_, CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_,
         CARRYB_2__3_, CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__6_,
         CARRYB_1__0_, SUMB_16__6_, SUMB_16__5_, SUMB_16__4_, SUMB_16__3_,
         SUMB_16__2_, SUMB_16__1_, SUMB_16__0_, SUMB_15__6_, SUMB_15__5_,
         SUMB_15__4_, SUMB_15__3_, SUMB_15__2_, SUMB_15__1_, SUMB_14__6_,
         SUMB_14__5_, SUMB_14__4_, SUMB_14__3_, SUMB_14__2_, SUMB_14__1_,
         SUMB_13__6_, SUMB_13__5_, SUMB_13__4_, SUMB_13__3_, SUMB_13__2_,
         SUMB_13__1_, SUMB_12__6_, SUMB_12__5_, SUMB_12__4_, SUMB_12__3_,
         SUMB_12__2_, SUMB_12__1_, SUMB_11__6_, SUMB_11__5_, SUMB_11__4_,
         SUMB_11__3_, SUMB_11__2_, SUMB_11__1_, SUMB_10__6_, SUMB_10__5_,
         SUMB_10__4_, SUMB_10__3_, SUMB_10__2_, SUMB_10__1_, SUMB_9__6_,
         SUMB_9__5_, SUMB_9__4_, SUMB_9__3_, SUMB_9__2_, SUMB_9__1_,
         SUMB_8__6_, SUMB_8__5_, SUMB_8__4_, SUMB_8__3_, SUMB_8__2_,
         SUMB_8__1_, SUMB_7__6_, SUMB_7__5_, SUMB_7__4_, SUMB_7__3_,
         SUMB_7__2_, SUMB_7__1_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_,
         SUMB_6__3_, SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_,
         SUMB_5__4_, SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_,
         SUMB_4__5_, SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_,
         SUMB_3__6_, SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_,
         SUMB_3__1_, SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_,
         SUMB_2__2_, SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_,
         SUMB_1__3_, SUMB_1__2_, SUMB_1__1_, PROD1_7_, A1_21_, A1_20_, A1_19_,
         A1_18_, A1_17_, A1_16_, A1_15_, A1_13_, A1_12_, A1_11_, A1_10_, A1_9_,
         A1_8_, A1_7_, A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, n4, n5, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57;

  ADDFHX4 S1_12_0 ( .A(ab_12__0_), .B(CARRYB_11__0_), .CI(SUMB_11__1_), .CO(
        CARRYB_12__0_), .S(A1_10_) );
  ADDFHX4 S2_12_1 ( .A(ab_12__1_), .B(CARRYB_11__1_), .CI(SUMB_11__2_), .CO(
        CARRYB_12__1_), .S(SUMB_12__1_) );
  multi16_7_DW01_add_0 FS_1 ( .A_21_(A1_21_), .A_20_(A1_20_), .A_19_(A1_19_), 
        .A_18_(A1_18_), .A_17_(A1_17_), .A_16_(A1_16_), .A_15_(A1_15_), 
        .A_14_(SUMB_16__0_), .A_13_(A1_13_), .A_12_(A1_12_), .A_11_(A1_11_), 
        .A_10_(A1_10_), .A_9_(A1_9_), .A_8_(A1_8_), .A_7_(A1_7_), .A_6_(A1_6_), 
        .A_5_(PROD1_7_), .B_21_(n37), .B_20_(n36), .B_19_(n35), .B_18_(n32), 
        .B_17_(n33), .B_16_(n34), .SUM_21_(PRODUCT_23_), .SUM_20_(PRODUCT_22_), 
        .SUM_19_(PRODUCT_21_), .SUM_18_(PRODUCT_20_), .SUM_17_(PRODUCT_19_), 
        .SUM_16_(PRODUCT_18_), .SUM_15_(PRODUCT_17_), .SUM_14_(PRODUCT_16_), 
        .SUM_13_(PRODUCT_15_), .SUM_12_(PRODUCT_14_), .SUM_11_(PRODUCT_13_), 
        .SUM_10_(PRODUCT_12_), .SUM_9_(PRODUCT_11_), .SUM_8_(PRODUCT_10_), 
        .SUM_7_(PRODUCT_9_), .SUM_6_(PRODUCT_8_), .SUM_5_(PRODUCT_7_) );
  ADDFX2 S5_6 ( .A(ab_16__6_), .B(CARRYB_15__6_), .CI(ab_15__7_), .CO(
        CARRYB_16__6_), .S(SUMB_16__6_) );
  ADDFHX4 S2_14_1 ( .A(ab_14__1_), .B(CARRYB_13__1_), .CI(SUMB_13__2_), .CO(
        CARRYB_14__1_), .S(SUMB_14__1_) );
  ADDFHX4 S2_11_1 ( .A(ab_11__1_), .B(CARRYB_10__1_), .CI(SUMB_10__2_), .CO(
        CARRYB_11__1_), .S(SUMB_11__1_) );
  ADDFHX1 S4_4 ( .A(ab_16__4_), .B(CARRYB_15__4_), .CI(SUMB_15__5_), .CO(
        CARRYB_16__4_), .S(SUMB_16__4_) );
  ADDFHX1 S4_5 ( .A(ab_16__5_), .B(CARRYB_15__5_), .CI(SUMB_15__6_), .CO(
        CARRYB_16__5_), .S(SUMB_16__5_) );
  ADDFHX2 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  ADDFHX2 S4_2 ( .A(ab_16__2_), .B(CARRYB_15__2_), .CI(SUMB_15__3_), .CO(
        CARRYB_16__2_), .S(SUMB_16__2_) );
  ADDFHX4 S2_15_2 ( .A(ab_15__2_), .B(CARRYB_14__2_), .CI(SUMB_14__3_), .CO(
        CARRYB_15__2_), .S(SUMB_15__2_) );
  ADDFHX2 S2_13_4 ( .A(ab_13__4_), .B(CARRYB_12__4_), .CI(SUMB_12__5_), .CO(
        CARRYB_13__4_), .S(SUMB_13__4_) );
  ADDFHX2 S2_13_3 ( .A(ab_13__3_), .B(CARRYB_12__3_), .CI(SUMB_12__4_), .CO(
        CARRYB_13__3_), .S(SUMB_13__3_) );
  ADDFHX2 S2_11_5 ( .A(ab_11__5_), .B(CARRYB_10__5_), .CI(SUMB_10__6_), .CO(
        CARRYB_11__5_), .S(SUMB_11__5_) );
  ADDFHX2 S2_11_4 ( .A(ab_11__4_), .B(CARRYB_10__4_), .CI(SUMB_10__5_), .CO(
        CARRYB_11__4_), .S(SUMB_11__4_) );
  ADDFHX4 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  ADDFHX4 S2_15_1 ( .A(ab_15__1_), .B(CARRYB_14__1_), .CI(SUMB_14__2_), .CO(
        CARRYB_15__1_), .S(SUMB_15__1_) );
  ADDFHX4 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  ADDFHX4 S2_15_3 ( .A(ab_15__3_), .B(CARRYB_14__3_), .CI(SUMB_14__4_), .CO(
        CARRYB_15__3_), .S(SUMB_15__3_) );
  ADDFHX4 S3_10_6 ( .A(ab_10__6_), .B(CARRYB_9__6_), .CI(ab_9__7_), .CO(
        CARRYB_10__6_), .S(SUMB_10__6_) );
  ADDFHX4 S3_7_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(
        CARRYB_7__6_), .S(SUMB_7__6_) );
  ADDFHX4 S2_12_5 ( .A(ab_12__5_), .B(CARRYB_11__5_), .CI(SUMB_11__6_), .CO(
        CARRYB_12__5_), .S(SUMB_12__5_) );
  ADDFHX2 S2_13_5 ( .A(ab_13__5_), .B(CARRYB_12__5_), .CI(SUMB_12__6_), .CO(
        CARRYB_13__5_), .S(SUMB_13__5_) );
  ADDFHX4 S2_2_2 ( .A(ab_2__2_), .B(n5), .CI(SUMB_1__3_), .CO(CARRYB_2__2_), 
        .S(SUMB_2__2_) );
  ADDFHX4 S1_8_0 ( .A(ab_8__0_), .B(CARRYB_7__0_), .CI(SUMB_7__1_), .CO(
        CARRYB_8__0_), .S(A1_6_) );
  ADDFHX4 S1_9_0 ( .A(ab_9__0_), .B(CARRYB_8__0_), .CI(SUMB_8__1_), .CO(
        CARRYB_9__0_), .S(A1_7_) );
  ADDFHX4 S1_11_0 ( .A(ab_11__0_), .B(CARRYB_10__0_), .CI(SUMB_10__1_), .CO(
        CARRYB_11__0_), .S(A1_9_) );
  ADDFHX4 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  ADDFHX4 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  ADDFHX4 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  ADDFHX4 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  ADDFHX4 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  ADDFHX4 S3_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(ab_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  ADDFHX4 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  ADDFHX4 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  ADDFHX4 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  ADDFHX4 S2_7_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  ADDFHX4 S2_11_2 ( .A(ab_11__2_), .B(CARRYB_10__2_), .CI(SUMB_10__3_), .CO(
        CARRYB_11__2_), .S(SUMB_11__2_) );
  ADDFHX4 S2_9_2 ( .A(ab_9__2_), .B(CARRYB_8__2_), .CI(SUMB_8__3_), .CO(
        CARRYB_9__2_), .S(SUMB_9__2_) );
  ADDFHX4 S2_10_2 ( .A(ab_10__2_), .B(CARRYB_9__2_), .CI(SUMB_9__3_), .CO(
        CARRYB_10__2_), .S(SUMB_10__2_) );
  ADDFHX4 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  ADDFHX4 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  ADDFHX4 S2_12_2 ( .A(ab_12__2_), .B(CARRYB_11__2_), .CI(SUMB_11__3_), .CO(
        CARRYB_12__2_), .S(SUMB_12__2_) );
  ADDFHX4 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  ADDFHX4 S2_8_3 ( .A(ab_8__3_), .B(CARRYB_7__3_), .CI(SUMB_7__4_), .CO(
        CARRYB_8__3_), .S(SUMB_8__3_) );
  ADDFHX4 S2_9_1 ( .A(ab_9__1_), .B(CARRYB_8__1_), .CI(SUMB_8__2_), .CO(
        CARRYB_9__1_), .S(SUMB_9__1_) );
  ADDFHX4 S2_10_1 ( .A(ab_10__1_), .B(CARRYB_9__1_), .CI(SUMB_9__2_), .CO(
        CARRYB_10__1_), .S(SUMB_10__1_) );
  ADDFHX4 S2_10_4 ( .A(ab_10__4_), .B(CARRYB_9__4_), .CI(SUMB_9__5_), .CO(
        CARRYB_10__4_), .S(SUMB_10__4_) );
  ADDFHX4 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  ADDFHX2 S3_14_6 ( .A(ab_14__6_), .B(CARRYB_13__6_), .CI(ab_13__7_), .CO(
        CARRYB_14__6_), .S(SUMB_14__6_) );
  ADDFHX1 S2_15_5 ( .A(ab_15__5_), .B(CARRYB_14__5_), .CI(SUMB_14__6_), .CO(
        CARRYB_15__5_), .S(SUMB_15__5_) );
  ADDFHX4 S3_13_6 ( .A(ab_13__6_), .B(CARRYB_12__6_), .CI(ab_12__7_), .CO(
        CARRYB_13__6_), .S(SUMB_13__6_) );
  ADDFHX4 S2_2_1 ( .A(ab_2__1_), .B(n4), .CI(SUMB_1__2_), .CO(CARRYB_2__1_), 
        .S(SUMB_2__1_) );
  ADDFHX2 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  ADDFHX4 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  ADDFHX4 S2_11_3 ( .A(ab_11__3_), .B(CARRYB_10__3_), .CI(SUMB_10__4_), .CO(
        CARRYB_11__3_), .S(SUMB_11__3_) );
  ADDFHX4 S2_12_3 ( .A(ab_12__3_), .B(CARRYB_11__3_), .CI(SUMB_11__4_), .CO(
        CARRYB_12__3_), .S(SUMB_12__3_) );
  ADDFHX4 S2_14_4 ( .A(ab_14__4_), .B(CARRYB_13__4_), .CI(SUMB_13__5_), .CO(
        CARRYB_14__4_), .S(SUMB_14__4_) );
  ADDFHX2 S2_15_4 ( .A(ab_15__4_), .B(CARRYB_14__4_), .CI(SUMB_14__5_), .CO(
        CARRYB_15__4_), .S(SUMB_15__4_) );
  ADDFHX4 S2_7_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  ADDFHX4 S2_10_3 ( .A(ab_10__3_), .B(CARRYB_9__3_), .CI(SUMB_9__4_), .CO(
        CARRYB_10__3_), .S(SUMB_10__3_) );
  ADDFHX4 S2_7_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  ADDFHX4 S2_8_2 ( .A(ab_8__2_), .B(CARRYB_7__2_), .CI(SUMB_7__3_), .CO(
        CARRYB_8__2_), .S(SUMB_8__2_) );
  ADDFHX4 S2_7_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  ADDFHX4 S2_8_1 ( .A(ab_8__1_), .B(CARRYB_7__1_), .CI(SUMB_7__2_), .CO(
        CARRYB_8__1_), .S(SUMB_8__1_) );
  ADDFHX2 S1_7_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(PROD1_7_) );
  ADDFHX1 S2_14_5 ( .A(ab_14__5_), .B(CARRYB_13__5_), .CI(SUMB_13__6_), .CO(
        CARRYB_14__5_), .S(SUMB_14__5_) );
  ADDFHX1 S4_0 ( .A(ab_16__0_), .B(CARRYB_15__0_), .CI(SUMB_15__1_), .CO(
        CARRYB_16__0_), .S(SUMB_16__0_) );
  ADDFHX2 S4_3 ( .A(ab_16__3_), .B(CARRYB_15__3_), .CI(SUMB_15__4_), .CO(
        CARRYB_16__3_), .S(SUMB_16__3_) );
  ADDFHX2 S1_13_0 ( .A(ab_13__0_), .B(CARRYB_12__0_), .CI(SUMB_12__1_), .CO(
        CARRYB_13__0_), .S(A1_11_) );
  ADDFHX2 S1_10_0 ( .A(ab_10__0_), .B(CARRYB_9__0_), .CI(SUMB_9__1_), .CO(
        CARRYB_10__0_), .S(A1_8_) );
  ADDFHX2 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  ADDFHX2 S2_2_5 ( .A(ab_2__5_), .B(n8), .CI(SUMB_1__6_), .CO(CARRYB_2__5_), 
        .S(SUMB_2__5_) );
  ADDFHX2 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  ADDFHX2 S2_8_5 ( .A(ab_8__5_), .B(CARRYB_7__5_), .CI(SUMB_7__6_), .CO(
        CARRYB_8__5_), .S(SUMB_8__5_) );
  ADDFHX2 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  ADDFHX2 S1_15_0 ( .A(ab_15__0_), .B(CARRYB_14__0_), .CI(SUMB_14__1_), .CO(
        CARRYB_15__0_), .S(A1_13_) );
  ADDFHX2 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  ADDFHX2 S3_8_6 ( .A(ab_8__6_), .B(CARRYB_7__6_), .CI(ab_7__7_), .CO(
        CARRYB_8__6_), .S(SUMB_8__6_) );
  ADDFHX2 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  ADDFHX2 S2_7_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  ADDFHX2 S2_8_4 ( .A(ab_8__4_), .B(CARRYB_7__4_), .CI(SUMB_7__5_), .CO(
        CARRYB_8__4_), .S(SUMB_8__4_) );
  ADDFHX2 S1_14_0 ( .A(ab_14__0_), .B(CARRYB_13__0_), .CI(SUMB_13__1_), .CO(
        CARRYB_14__0_), .S(A1_12_) );
  ADDFHX2 S2_2_4 ( .A(ab_2__4_), .B(n6), .CI(SUMB_1__5_), .CO(CARRYB_2__4_), 
        .S(SUMB_2__4_) );
  ADDFHX2 S2_10_5 ( .A(ab_10__5_), .B(CARRYB_9__5_), .CI(SUMB_9__6_), .CO(
        CARRYB_10__5_), .S(SUMB_10__5_) );
  ADDFHX4 S3_11_6 ( .A(ab_11__6_), .B(CARRYB_10__6_), .CI(ab_10__7_), .CO(
        CARRYB_11__6_), .S(SUMB_11__6_) );
  ADDFHX4 S3_12_6 ( .A(ab_12__6_), .B(CARRYB_11__6_), .CI(ab_11__7_), .CO(
        CARRYB_12__6_), .S(SUMB_12__6_) );
  ADDFHX4 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  ADDFHX4 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  ADDFHX4 S2_9_3 ( .A(ab_9__3_), .B(CARRYB_8__3_), .CI(SUMB_8__4_), .CO(
        CARRYB_9__3_), .S(SUMB_9__3_) );
  ADDFHX4 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  ADDFHX4 S2_13_1 ( .A(ab_13__1_), .B(CARRYB_12__1_), .CI(SUMB_12__2_), .CO(
        CARRYB_13__1_), .S(SUMB_13__1_) );
  ADDFHX4 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  ADDFHX4 S2_2_3 ( .A(ab_2__3_), .B(n7), .CI(SUMB_1__4_), .CO(CARRYB_2__3_), 
        .S(SUMB_2__3_) );
  ADDFHX4 S3_9_6 ( .A(ab_9__6_), .B(CARRYB_8__6_), .CI(ab_8__7_), .CO(
        CARRYB_9__6_), .S(SUMB_9__6_) );
  ADDFHX1 S3_15_6 ( .A(ab_15__6_), .B(CARRYB_14__6_), .CI(ab_14__7_), .CO(
        CARRYB_15__6_), .S(SUMB_15__6_) );
  ADDFHX4 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  ADDFHX4 S2_13_2 ( .A(ab_13__2_), .B(CARRYB_12__2_), .CI(SUMB_12__3_), .CO(
        CARRYB_13__2_), .S(SUMB_13__2_) );
  ADDFHX4 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  AND2X2 U2 ( .A(A[1]), .B(B[3]), .Y(ab_1__3_) );
  INVX4 U3 ( .A(n38), .Y(CARRYB_1__6_) );
  NAND2X2 U4 ( .A(ab_0__7_), .B(ab_1__6_), .Y(n38) );
  AND2X4 U5 ( .A(CARRYB_16__1_), .B(SUMB_16__2_), .Y(n33) );
  NAND3X2 U6 ( .A(n31), .B(n29), .C(n30), .Y(CARRYB_16__1_) );
  AND2X2 U7 ( .A(A[3]), .B(B[6]), .Y(ab_3__6_) );
  AND2X2 U8 ( .A(A[2]), .B(B[6]), .Y(ab_2__6_) );
  INVX4 U9 ( .A(B[6]), .Y(n45) );
  NOR2X4 U10 ( .A(n47), .B(n42), .Y(ab_0__4_) );
  INVX4 U11 ( .A(B[4]), .Y(n47) );
  XOR2X4 U12 ( .A(CARRYB_16__2_), .B(SUMB_16__3_), .Y(A1_17_) );
  INVX4 U13 ( .A(B[2]), .Y(n49) );
  AND2X1 U14 ( .A(A[1]), .B(B[2]), .Y(ab_1__2_) );
  XOR2X1 U15 ( .A(CARRYB_5__5_), .B(n12), .Y(SUMB_6__5_) );
  NAND3X2 U16 ( .A(n19), .B(n17), .C(n18), .Y(CARRYB_9__5_) );
  INVXL U17 ( .A(A[0]), .Y(n42) );
  NOR2X1 U18 ( .A(n45), .B(n42), .Y(ab_0__6_) );
  NOR2X1 U19 ( .A(n49), .B(n42), .Y(ab_0__2_) );
  CLKINVX3 U20 ( .A(B[3]), .Y(n48) );
  INVX1 U21 ( .A(n41), .Y(n40) );
  NOR2X1 U22 ( .A(n53), .B(n50), .Y(ab_16__1_) );
  AND2X2 U24 ( .A(ab_0__2_), .B(n52), .Y(n4) );
  AND2X2 U25 ( .A(ab_0__3_), .B(ab_1__2_), .Y(n5) );
  AND2X2 U26 ( .A(ab_0__5_), .B(ab_1__4_), .Y(n6) );
  AND2X2 U27 ( .A(ab_0__4_), .B(ab_1__3_), .Y(n7) );
  AND2X2 U28 ( .A(ab_0__6_), .B(ab_1__5_), .Y(n8) );
  XOR3X4 U29 ( .A(CARRYB_11__4_), .B(ab_12__4_), .C(SUMB_11__5_), .Y(
        SUMB_12__4_) );
  NAND3X4 U30 ( .A(n11), .B(n9), .C(n10), .Y(CARRYB_9__4_) );
  NAND3X2 U31 ( .A(n15), .B(n13), .C(n14), .Y(CARRYB_6__5_) );
  NAND2X1 U32 ( .A(CARRYB_8__5_), .B(SUMB_8__6_), .Y(n17) );
  XOR3X4 U33 ( .A(CARRYB_8__4_), .B(ab_9__4_), .C(SUMB_8__5_), .Y(SUMB_9__4_)
         );
  NAND2X1 U34 ( .A(SUMB_8__5_), .B(CARRYB_8__4_), .Y(n9) );
  NAND2X1 U35 ( .A(ab_9__4_), .B(CARRYB_8__4_), .Y(n10) );
  NAND2X1 U36 ( .A(ab_9__4_), .B(SUMB_8__5_), .Y(n11) );
  XOR2X4 U37 ( .A(SUMB_5__6_), .B(ab_6__5_), .Y(n12) );
  NAND2X1 U38 ( .A(SUMB_5__6_), .B(CARRYB_5__5_), .Y(n13) );
  NAND2X1 U39 ( .A(ab_6__5_), .B(CARRYB_5__5_), .Y(n14) );
  NAND2X1 U40 ( .A(ab_6__5_), .B(SUMB_5__6_), .Y(n15) );
  XOR2X4 U41 ( .A(SUMB_8__6_), .B(n16), .Y(SUMB_9__5_) );
  XOR2X2 U42 ( .A(CARRYB_16__0_), .B(SUMB_16__1_), .Y(A1_15_) );
  AND2X1 U43 ( .A(A[10]), .B(n39), .Y(ab_10__7_) );
  AND2X1 U44 ( .A(A[8]), .B(n39), .Y(ab_8__7_) );
  AND2X1 U45 ( .A(A[7]), .B(n39), .Y(ab_7__7_) );
  AND2X1 U46 ( .A(A[6]), .B(n39), .Y(ab_6__7_) );
  AND2X1 U47 ( .A(A[5]), .B(n39), .Y(ab_5__7_) );
  AND2X1 U48 ( .A(A[4]), .B(n39), .Y(ab_4__7_) );
  AND2X2 U49 ( .A(CARRYB_16__0_), .B(SUMB_16__1_), .Y(n34) );
  NAND2XL U50 ( .A(ab_9__5_), .B(CARRYB_8__5_), .Y(n19) );
  XOR2X2 U51 ( .A(CARRYB_16__1_), .B(SUMB_16__2_), .Y(A1_16_) );
  NAND3X4 U52 ( .A(n25), .B(n23), .C(n24), .Y(CARRYB_12__4_) );
  NAND2X1 U53 ( .A(ab_14__3_), .B(CARRYB_13__3_), .Y(n27) );
  NAND3X4 U54 ( .A(n28), .B(n26), .C(n27), .Y(CARRYB_14__3_) );
  XOR2X4 U55 ( .A(CARRYB_8__5_), .B(ab_9__5_), .Y(n16) );
  NAND2X1 U56 ( .A(ab_9__5_), .B(SUMB_8__6_), .Y(n18) );
  AND2X1 U57 ( .A(A[9]), .B(B[5]), .Y(ab_9__5_) );
  XOR3X4 U58 ( .A(CARRYB_13__2_), .B(ab_14__2_), .C(SUMB_13__3_), .Y(
        SUMB_14__2_) );
  NAND2XL U59 ( .A(SUMB_13__3_), .B(CARRYB_13__2_), .Y(n20) );
  NAND2XL U60 ( .A(ab_14__2_), .B(CARRYB_13__2_), .Y(n21) );
  NAND2XL U61 ( .A(ab_14__2_), .B(SUMB_13__3_), .Y(n22) );
  NAND3X2 U62 ( .A(n22), .B(n20), .C(n21), .Y(CARRYB_14__2_) );
  NAND2X1 U63 ( .A(SUMB_11__5_), .B(CARRYB_11__4_), .Y(n23) );
  NAND2X1 U64 ( .A(ab_12__4_), .B(CARRYB_11__4_), .Y(n24) );
  NAND2X1 U65 ( .A(ab_12__4_), .B(SUMB_11__5_), .Y(n25) );
  XOR3X2 U66 ( .A(CARRYB_13__3_), .B(ab_14__3_), .C(SUMB_13__4_), .Y(
        SUMB_14__3_) );
  NAND2X1 U67 ( .A(SUMB_13__4_), .B(CARRYB_13__3_), .Y(n26) );
  NAND2X1 U68 ( .A(ab_14__3_), .B(SUMB_13__4_), .Y(n28) );
  XOR3X4 U69 ( .A(CARRYB_15__1_), .B(ab_16__1_), .C(SUMB_15__2_), .Y(
        SUMB_16__1_) );
  NAND2XL U70 ( .A(SUMB_15__2_), .B(CARRYB_15__1_), .Y(n29) );
  NAND2XL U71 ( .A(ab_16__1_), .B(CARRYB_15__1_), .Y(n30) );
  NAND2XL U72 ( .A(ab_16__1_), .B(SUMB_15__2_), .Y(n31) );
  INVX2 U73 ( .A(B[5]), .Y(n46) );
  AND2X1 U74 ( .A(A[2]), .B(B[3]), .Y(ab_2__3_) );
  INVX4 U75 ( .A(n39), .Y(n51) );
  NOR2X1 U76 ( .A(n46), .B(n42), .Y(ab_0__5_) );
  XOR2X1 U77 ( .A(ab_1__5_), .B(ab_0__6_), .Y(SUMB_1__5_) );
  AND2X1 U78 ( .A(A[9]), .B(n39), .Y(ab_9__7_) );
  AND2X1 U79 ( .A(A[9]), .B(n40), .Y(ab_9__0_) );
  AND2X1 U80 ( .A(A[11]), .B(B[1]), .Y(ab_11__1_) );
  AND2X1 U81 ( .A(A[10]), .B(B[1]), .Y(ab_10__1_) );
  AND2X1 U82 ( .A(A[9]), .B(B[1]), .Y(ab_9__1_) );
  AND2X1 U83 ( .A(A[7]), .B(B[1]), .Y(ab_7__1_) );
  AND2X1 U84 ( .A(A[6]), .B(B[1]), .Y(ab_6__1_) );
  AND2X1 U85 ( .A(A[10]), .B(n40), .Y(ab_10__0_) );
  AND2X1 U86 ( .A(A[7]), .B(n40), .Y(ab_7__0_) );
  AND2X1 U87 ( .A(A[6]), .B(n40), .Y(ab_6__0_) );
  INVXL U88 ( .A(B[1]), .Y(n50) );
  AND2X1 U89 ( .A(A[10]), .B(B[5]), .Y(ab_10__5_) );
  NOR2X1 U90 ( .A(n51), .B(n42), .Y(ab_0__7_) );
  AND2X1 U91 ( .A(A[8]), .B(B[5]), .Y(ab_8__5_) );
  AND2X1 U92 ( .A(A[7]), .B(B[5]), .Y(ab_7__5_) );
  AND2X1 U93 ( .A(A[6]), .B(B[5]), .Y(ab_6__5_) );
  AND2X1 U94 ( .A(A[3]), .B(B[5]), .Y(ab_3__5_) );
  AND2X1 U95 ( .A(A[11]), .B(B[5]), .Y(ab_11__5_) );
  AND2X1 U96 ( .A(A[5]), .B(B[5]), .Y(ab_5__5_) );
  AND2X1 U97 ( .A(A[2]), .B(B[2]), .Y(ab_2__2_) );
  AND2X1 U98 ( .A(A[2]), .B(B[4]), .Y(ab_2__4_) );
  NAND2XL U99 ( .A(A[1]), .B(B[1]), .Y(n44) );
  AND2X1 U100 ( .A(A[2]), .B(B[1]), .Y(ab_2__1_) );
  NOR2XL U101 ( .A(n57), .B(n50), .Y(ab_12__1_) );
  AND2X1 U102 ( .A(A[3]), .B(n40), .Y(ab_3__0_) );
  NOR2XL U103 ( .A(n44), .B(n43), .Y(CARRYB_1__0_) );
  AND2X1 U104 ( .A(A[2]), .B(n40), .Y(ab_2__0_) );
  XOR2X1 U105 ( .A(CARRYB_16__3_), .B(SUMB_16__4_), .Y(A1_18_) );
  AND2X2 U106 ( .A(CARRYB_16__2_), .B(SUMB_16__3_), .Y(n32) );
  XOR2X1 U107 ( .A(CARRYB_16__4_), .B(SUMB_16__5_), .Y(A1_19_) );
  AND2X2 U108 ( .A(CARRYB_16__3_), .B(SUMB_16__4_), .Y(n35) );
  AND2X2 U109 ( .A(CARRYB_16__4_), .B(SUMB_16__5_), .Y(n36) );
  NOR2X1 U110 ( .A(n53), .B(n46), .Y(ab_16__5_) );
  NOR2X1 U111 ( .A(n53), .B(n47), .Y(ab_16__4_) );
  INVX1 U112 ( .A(n44), .Y(n52) );
  AND2X2 U113 ( .A(A[4]), .B(B[1]), .Y(ab_4__1_) );
  AND2X2 U114 ( .A(A[11]), .B(n40), .Y(ab_11__0_) );
  AND2X2 U115 ( .A(A[8]), .B(B[1]), .Y(ab_8__1_) );
  AND2X2 U116 ( .A(A[5]), .B(B[1]), .Y(ab_5__1_) );
  AND2X2 U117 ( .A(A[8]), .B(n40), .Y(ab_8__0_) );
  AND2X2 U118 ( .A(A[5]), .B(n40), .Y(ab_5__0_) );
  AND2X2 U119 ( .A(A[4]), .B(n40), .Y(ab_4__0_) );
  XOR2X1 U120 ( .A(n52), .B(ab_0__2_), .Y(SUMB_1__1_) );
  XOR2X1 U121 ( .A(CARRYB_16__5_), .B(SUMB_16__6_), .Y(A1_20_) );
  XOR2X1 U122 ( .A(CARRYB_16__6_), .B(ab_16__7_), .Y(A1_21_) );
  INVX1 U123 ( .A(B[0]), .Y(n41) );
  AND2X2 U124 ( .A(CARRYB_16__5_), .B(SUMB_16__6_), .Y(n37) );
  NOR2X1 U125 ( .A(n53), .B(n51), .Y(ab_16__7_) );
  NOR2X1 U126 ( .A(n48), .B(n42), .Y(ab_0__3_) );
  AND2X2 U127 ( .A(A[3]), .B(B[1]), .Y(ab_3__1_) );
  AND2X1 U128 ( .A(A[2]), .B(B[5]), .Y(ab_2__5_) );
  XOR2X1 U129 ( .A(ab_1__6_), .B(ab_0__7_), .Y(SUMB_1__6_) );
  NOR2XL U130 ( .A(n54), .B(n51), .Y(ab_15__7_) );
  BUFX3 U131 ( .A(B[7]), .Y(n39) );
  NOR2X1 U132 ( .A(n55), .B(n50), .Y(ab_14__1_) );
  NOR2X1 U133 ( .A(n56), .B(n50), .Y(ab_13__1_) );
  AND2X1 U134 ( .A(A[11]), .B(B[2]), .Y(ab_11__2_) );
  AND2X1 U135 ( .A(A[10]), .B(B[2]), .Y(ab_10__2_) );
  AND2X1 U136 ( .A(A[9]), .B(B[2]), .Y(ab_9__2_) );
  AND2X1 U137 ( .A(A[8]), .B(B[2]), .Y(ab_8__2_) );
  AND2X1 U138 ( .A(A[11]), .B(B[4]), .Y(ab_11__4_) );
  AND2X1 U139 ( .A(A[10]), .B(B[4]), .Y(ab_10__4_) );
  NOR2XL U140 ( .A(n55), .B(n47), .Y(ab_14__4_) );
  AND2X1 U141 ( .A(A[9]), .B(B[4]), .Y(ab_9__4_) );
  NOR2XL U142 ( .A(n56), .B(n47), .Y(ab_13__4_) );
  AND2X1 U143 ( .A(A[7]), .B(B[2]), .Y(ab_7__2_) );
  AND2X1 U144 ( .A(A[8]), .B(B[4]), .Y(ab_8__4_) );
  AND2X1 U145 ( .A(A[7]), .B(B[4]), .Y(ab_7__4_) );
  NOR2XL U146 ( .A(n54), .B(n46), .Y(ab_15__5_) );
  AND2X1 U147 ( .A(A[3]), .B(B[2]), .Y(ab_3__2_) );
  AND2X1 U148 ( .A(A[4]), .B(B[2]), .Y(ab_4__2_) );
  AND2X1 U149 ( .A(A[5]), .B(B[2]), .Y(ab_5__2_) );
  AND2X1 U150 ( .A(A[6]), .B(B[2]), .Y(ab_6__2_) );
  AND2X1 U151 ( .A(A[3]), .B(B[3]), .Y(ab_3__3_) );
  NOR2XL U152 ( .A(n56), .B(n46), .Y(ab_13__5_) );
  AND2X1 U153 ( .A(A[3]), .B(B[4]), .Y(ab_3__4_) );
  AND2X1 U154 ( .A(A[6]), .B(B[4]), .Y(ab_6__4_) );
  AND2X1 U155 ( .A(A[4]), .B(B[4]), .Y(ab_4__4_) );
  AND2X1 U156 ( .A(A[5]), .B(B[4]), .Y(ab_5__4_) );
  NOR2XL U157 ( .A(n57), .B(n46), .Y(ab_12__5_) );
  AND2X1 U158 ( .A(A[4]), .B(B[5]), .Y(ab_4__5_) );
  AND2X1 U159 ( .A(A[2]), .B(n39), .Y(ab_2__7_) );
  AND2X1 U160 ( .A(A[3]), .B(n39), .Y(ab_3__7_) );
  AND2X1 U161 ( .A(A[11]), .B(n39), .Y(ab_11__7_) );
  NOR2XL U162 ( .A(n56), .B(n51), .Y(ab_13__7_) );
  XOR2X1 U163 ( .A(ab_1__2_), .B(ab_0__3_), .Y(SUMB_1__2_) );
  XOR2X1 U164 ( .A(ab_1__4_), .B(ab_0__5_), .Y(SUMB_1__4_) );
  NOR2XL U165 ( .A(n55), .B(n51), .Y(ab_14__7_) );
  NOR2XL U166 ( .A(n57), .B(n51), .Y(ab_12__7_) );
  NOR2X1 U167 ( .A(n54), .B(n50), .Y(ab_15__1_) );
  NOR2XL U168 ( .A(n54), .B(n47), .Y(ab_15__4_) );
  NOR2XL U169 ( .A(n57), .B(n47), .Y(ab_12__4_) );
  NOR2XL U170 ( .A(n55), .B(n46), .Y(ab_14__5_) );
  XOR2X1 U171 ( .A(ab_1__3_), .B(ab_0__4_), .Y(SUMB_1__3_) );
  INVX1 U172 ( .A(A[16]), .Y(n53) );
  NAND2XL U173 ( .A(A[0]), .B(n40), .Y(n43) );
  INVX1 U174 ( .A(A[12]), .Y(n57) );
  INVX1 U175 ( .A(A[13]), .Y(n56) );
  INVX1 U176 ( .A(A[14]), .Y(n55) );
  INVX1 U177 ( .A(A[15]), .Y(n54) );
  NOR2XL U178 ( .A(n53), .B(n49), .Y(ab_16__2_) );
  NOR2XL U179 ( .A(n54), .B(n49), .Y(ab_15__2_) );
  NOR2XL U180 ( .A(n55), .B(n49), .Y(ab_14__2_) );
  NOR2XL U181 ( .A(n56), .B(n49), .Y(ab_13__2_) );
  NOR2XL U182 ( .A(n57), .B(n49), .Y(ab_12__2_) );
  AND2X2 U183 ( .A(A[1]), .B(B[6]), .Y(ab_1__6_) );
  NOR2XL U184 ( .A(n53), .B(n45), .Y(ab_16__6_) );
  NOR2XL U185 ( .A(n54), .B(n45), .Y(ab_15__6_) );
  NOR2XL U186 ( .A(n55), .B(n45), .Y(ab_14__6_) );
  NOR2XL U187 ( .A(n56), .B(n45), .Y(ab_13__6_) );
  NOR2XL U188 ( .A(n57), .B(n45), .Y(ab_12__6_) );
  AND2X1 U189 ( .A(A[11]), .B(B[6]), .Y(ab_11__6_) );
  AND2X1 U190 ( .A(A[10]), .B(B[6]), .Y(ab_10__6_) );
  AND2X1 U191 ( .A(A[9]), .B(B[6]), .Y(ab_9__6_) );
  AND2X1 U192 ( .A(A[8]), .B(B[6]), .Y(ab_8__6_) );
  AND2X1 U193 ( .A(A[7]), .B(B[6]), .Y(ab_7__6_) );
  AND2X1 U194 ( .A(A[6]), .B(B[6]), .Y(ab_6__6_) );
  AND2X1 U195 ( .A(A[5]), .B(B[6]), .Y(ab_5__6_) );
  AND2X1 U196 ( .A(A[4]), .B(B[6]), .Y(ab_4__6_) );
  AND2X1 U197 ( .A(A[1]), .B(n39), .Y(ab_1__7_) );
  AND2X2 U198 ( .A(A[1]), .B(B[5]), .Y(ab_1__5_) );
  AND2X2 U199 ( .A(A[1]), .B(B[4]), .Y(ab_1__4_) );
  NOR2XL U200 ( .A(n53), .B(n48), .Y(ab_16__3_) );
  NOR2XL U201 ( .A(n54), .B(n48), .Y(ab_15__3_) );
  NOR2XL U202 ( .A(n55), .B(n48), .Y(ab_14__3_) );
  NOR2XL U203 ( .A(n56), .B(n48), .Y(ab_13__3_) );
  NOR2XL U204 ( .A(n57), .B(n48), .Y(ab_12__3_) );
  AND2X1 U205 ( .A(A[11]), .B(B[3]), .Y(ab_11__3_) );
  AND2X1 U206 ( .A(A[10]), .B(B[3]), .Y(ab_10__3_) );
  AND2X1 U207 ( .A(A[9]), .B(B[3]), .Y(ab_9__3_) );
  AND2X1 U208 ( .A(A[8]), .B(B[3]), .Y(ab_8__3_) );
  AND2X1 U209 ( .A(A[7]), .B(B[3]), .Y(ab_7__3_) );
  AND2X1 U210 ( .A(A[6]), .B(B[3]), .Y(ab_6__3_) );
  AND2X1 U211 ( .A(A[5]), .B(B[3]), .Y(ab_5__3_) );
  AND2X1 U212 ( .A(A[4]), .B(B[3]), .Y(ab_4__3_) );
  NOR2X1 U214 ( .A(n41), .B(n53), .Y(ab_16__0_) );
  NOR2X1 U215 ( .A(n41), .B(n54), .Y(ab_15__0_) );
  NOR2X1 U216 ( .A(n41), .B(n55), .Y(ab_14__0_) );
  NOR2X1 U217 ( .A(n41), .B(n56), .Y(ab_13__0_) );
  NOR2X1 U218 ( .A(n41), .B(n57), .Y(ab_12__0_) );
endmodule


module multi16_7 ( in_17bit, in_8bit, out );
  input [16:0] in_17bit;
  input [7:0] in_8bit;
  output [16:0] out;
  wire   N19, N20, N21, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114;
  wire   [16:1] in_17bit_b;
  wire   [7:1] in_8bit_b;
  wire   [23:8] mul;
  wire   [16:13] sub_add_52_b0_carry;

  multi16_7_DW02_mult_0 mult_55 ( .A({in_17bit_b, in_17bit[0]}), .B({in_8bit_b, 
        in_8bit[0]}), .PRODUCT_23_(mul[23]), .PRODUCT_22_(mul[22]), 
        .PRODUCT_21_(mul[21]), .PRODUCT_20_(mul[20]), .PRODUCT_19_(mul[19]), 
        .PRODUCT_18_(mul[18]), .PRODUCT_17_(mul[17]), .PRODUCT_16_(mul[16]), 
        .PRODUCT_15_(mul[15]), .PRODUCT_14_(mul[14]), .PRODUCT_13_(mul[13]), 
        .PRODUCT_12_(mul[12]), .PRODUCT_11_(mul[11]), .PRODUCT_10_(mul[10]), 
        .PRODUCT_9_(mul[9]), .PRODUCT_8_(mul[8]), .PRODUCT_7_(out[0]) );
  AND3X4 U2 ( .A(in_17bit[1]), .B(n25), .C(in_17bit[0]), .Y(n18) );
  NOR2X2 U3 ( .A(n37), .B(n36), .Y(n39) );
  NAND2BX2 U4 ( .AN(in_8bit[0]), .B(n29), .Y(n37) );
  NAND2BXL U5 ( .AN(in_8bit[3]), .B(n24), .Y(n36) );
  CLKINVX2 U6 ( .A(in_8bit[4]), .Y(n24) );
  NOR2X4 U7 ( .A(mul[20]), .B(n102), .Y(n5) );
  XNOR2X4 U8 ( .A(n33), .B(n24), .Y(in_8bit_b[4]) );
  OAI21X1 U9 ( .A0(in_8bit[2]), .A1(n37), .B0(n20), .Y(n32) );
  CLKINVX3 U10 ( .A(n22), .Y(n20) );
  NAND2X1 U11 ( .A(n40), .B(in_8bit[6]), .Y(n3) );
  NAND2X2 U12 ( .A(n1), .B(n2), .Y(n4) );
  NAND2X4 U13 ( .A(n3), .B(n4), .Y(in_8bit_b[6]) );
  INVX1 U14 ( .A(n40), .Y(n1) );
  CLKINVXL U15 ( .A(in_8bit[6]), .Y(n2) );
  NAND2X1 U16 ( .A(n41), .B(n20), .Y(n40) );
  NOR2X2 U17 ( .A(in_17bit[1]), .B(n25), .Y(n42) );
  XOR2X2 U18 ( .A(n31), .B(n30), .Y(in_8bit_b[2]) );
  XOR2X2 U19 ( .A(in_17bit[2]), .B(n43), .Y(in_17bit_b[2]) );
  NOR2X2 U20 ( .A(n26), .B(n19), .Y(n43) );
  NOR2X1 U21 ( .A(mul[15]), .B(n93), .Y(n12) );
  NOR2X2 U22 ( .A(n13), .B(n9), .Y(n97) );
  INVX2 U23 ( .A(mul[22]), .Y(n108) );
  NOR2BX2 U24 ( .AN(n14), .B(n21), .Y(n33) );
  XOR2X1 U25 ( .A(n29), .B(n28), .Y(in_8bit_b[1]) );
  NOR2X1 U26 ( .A(mul[13]), .B(n89), .Y(n11) );
  NOR2X2 U27 ( .A(mul[16]), .B(n10), .Y(n9) );
  INVX2 U28 ( .A(n100), .Y(n8) );
  XOR2X1 U29 ( .A(mul[14]), .B(n92), .Y(out[7]) );
  NOR2X1 U30 ( .A(n13), .B(n11), .Y(n92) );
  NOR2X2 U31 ( .A(n13), .B(n5), .Y(n105) );
  INVX1 U32 ( .A(in_17bit[16]), .Y(n27) );
  INVX1 U33 ( .A(n89), .Y(n91) );
  INVXL U34 ( .A(in_8bit[3]), .Y(n23) );
  INVX1 U35 ( .A(n93), .Y(n95) );
  NAND2BX1 U36 ( .AN(mul[14]), .B(n11), .Y(n93) );
  NAND2X1 U37 ( .A(in_8bit[0]), .B(n20), .Y(n28) );
  BUFX1 U38 ( .A(mul[19]), .Y(n6) );
  NOR2BX4 U39 ( .AN(n77), .B(n109), .Y(n107) );
  INVX4 U40 ( .A(n102), .Y(n104) );
  NOR3X1 U41 ( .A(n36), .B(in_8bit[2]), .C(n37), .Y(n34) );
  XOR2X2 U42 ( .A(n23), .B(n32), .Y(in_8bit_b[3]) );
  OR3X2 U43 ( .A(n37), .B(in_8bit[3]), .C(in_8bit[2]), .Y(n14) );
  NOR2X2 U44 ( .A(n13), .B(n7), .Y(n101) );
  NOR2XL U45 ( .A(n27), .B(n46), .Y(n45) );
  NAND2X2 U46 ( .A(n39), .B(n38), .Y(n41) );
  NOR2X4 U47 ( .A(in_8bit[5]), .B(in_8bit[2]), .Y(n38) );
  NOR2X4 U48 ( .A(n13), .B(n104), .Y(n103) );
  XOR2X4 U49 ( .A(n105), .B(mul[21]), .Y(out[14]) );
  XOR2X4 U50 ( .A(mul[18]), .B(n99), .Y(out[11]) );
  NAND2BX4 U51 ( .AN(mul[19]), .B(n7), .Y(n102) );
  INVX4 U52 ( .A(n98), .Y(n100) );
  NAND2BX4 U53 ( .AN(mul[21]), .B(n5), .Y(n106) );
  INVX4 U54 ( .A(n106), .Y(n109) );
  NAND2BX4 U55 ( .AN(mul[17]), .B(n9), .Y(n98) );
  NOR2X4 U56 ( .A(mul[18]), .B(n8), .Y(n7) );
  CLKINVX2 U57 ( .A(in_8bit[1]), .Y(n29) );
  XOR2X2 U58 ( .A(n35), .B(in_8bit[5]), .Y(in_8bit_b[5]) );
  NOR2X1 U59 ( .A(n34), .B(n21), .Y(n35) );
  NAND2X1 U60 ( .A(n66), .B(n25), .Y(n65) );
  INVX4 U61 ( .A(n27), .Y(n25) );
  XNOR2X1 U62 ( .A(n25), .B(n20), .Y(n13) );
  INVX1 U63 ( .A(n12), .Y(n10) );
  NOR2XL U64 ( .A(n13), .B(n12), .Y(n96) );
  XOR2X1 U65 ( .A(in_17bit[3]), .B(n45), .Y(in_17bit_b[3]) );
  NAND2BXL U66 ( .AN(mul[10]), .B(n82), .Y(n83) );
  XOR2X1 U67 ( .A(mul[13]), .B(n90), .Y(out[6]) );
  NOR2XL U68 ( .A(n13), .B(n91), .Y(n90) );
  XOR2X1 U69 ( .A(mul[15]), .B(n94), .Y(out[8]) );
  NOR2XL U70 ( .A(n13), .B(n95), .Y(n94) );
  NOR2XL U71 ( .A(n13), .B(n85), .Y(n84) );
  NOR2XL U72 ( .A(n13), .B(n17), .Y(n79) );
  XNOR2X1 U73 ( .A(mul[8]), .B(n78), .Y(out[1]) );
  INVXL U74 ( .A(in_8bit[7]), .Y(n22) );
  INVXL U75 ( .A(in_8bit[7]), .Y(n21) );
  NAND2XL U76 ( .A(n50), .B(n49), .Y(n52) );
  NAND2BXL U77 ( .AN(n52), .B(n53), .Y(n54) );
  NOR2XL U78 ( .A(n26), .B(n64), .Y(n62) );
  NAND2XL U79 ( .A(n57), .B(n56), .Y(n59) );
  NAND2XL U80 ( .A(n64), .B(n63), .Y(n66) );
  NAND2BXL U81 ( .AN(n59), .B(n60), .Y(n61) );
  NOR2XL U82 ( .A(n26), .B(n71), .Y(n69) );
  NAND2XL U83 ( .A(n75), .B(n25), .Y(n72) );
  NAND2XL U84 ( .A(n71), .B(n70), .Y(n75) );
  NAND2BXL U85 ( .AN(n66), .B(n67), .Y(n68) );
  AND2X1 U86 ( .A(N21), .B(n25), .Y(in_17bit_b[16]) );
  INVX1 U87 ( .A(n44), .Y(n46) );
  NAND2XL U88 ( .A(n20), .B(n37), .Y(n30) );
  NAND2BXL U89 ( .AN(in_17bit[3]), .B(n46), .Y(n47) );
  MX2X1 U90 ( .A(in_17bit[12]), .B(n15), .S0(n25), .Y(in_17bit_b[12]) );
  XNOR2X1 U91 ( .A(in_17bit[12]), .B(n73), .Y(n15) );
  MX2X1 U92 ( .A(in_17bit[13]), .B(n16), .S0(n25), .Y(in_17bit_b[13]) );
  XNOR2X1 U93 ( .A(n76), .B(n112), .Y(n16) );
  MX2X1 U94 ( .A(in_17bit[14]), .B(N19), .S0(n25), .Y(in_17bit_b[14]) );
  MX2X1 U95 ( .A(in_17bit[15]), .B(N20), .S0(n25), .Y(in_17bit_b[15]) );
  NOR2XL U96 ( .A(in_17bit[11]), .B(n75), .Y(n73) );
  INVX1 U97 ( .A(n86), .Y(n88) );
  NAND2BX1 U98 ( .AN(mul[11]), .B(n85), .Y(n86) );
  INVX1 U99 ( .A(n83), .Y(n85) );
  INVX1 U100 ( .A(n80), .Y(n82) );
  NAND2BX1 U101 ( .AN(mul[9]), .B(n17), .Y(n80) );
  NOR2X1 U102 ( .A(mul[8]), .B(out[0]), .Y(n17) );
  NAND2BX1 U103 ( .AN(mul[12]), .B(n88), .Y(n89) );
  XOR2X1 U104 ( .A(mul[16]), .B(n96), .Y(out[9]) );
  XOR2X1 U105 ( .A(mul[10]), .B(n81), .Y(out[3]) );
  NOR2X1 U106 ( .A(n13), .B(n82), .Y(n81) );
  XOR2X1 U107 ( .A(mul[9]), .B(n79), .Y(out[2]) );
  XOR2X1 U108 ( .A(mul[12]), .B(n87), .Y(out[5]) );
  NOR2X1 U109 ( .A(n13), .B(n88), .Y(n87) );
  XOR2X1 U110 ( .A(mul[11]), .B(n84), .Y(out[4]) );
  NAND2X1 U111 ( .A(out[0]), .B(n77), .Y(n78) );
  INVX1 U112 ( .A(n13), .Y(n77) );
  NOR3XL U113 ( .A(n41), .B(in_8bit[6]), .C(n22), .Y(in_8bit_b[7]) );
  XNOR2X1 U114 ( .A(n48), .B(n49), .Y(in_17bit_b[4]) );
  NOR2X1 U115 ( .A(n26), .B(n50), .Y(n48) );
  XNOR2X1 U116 ( .A(n55), .B(n56), .Y(in_17bit_b[6]) );
  NOR2X1 U117 ( .A(n26), .B(n57), .Y(n55) );
  XNOR2X1 U118 ( .A(n62), .B(n63), .Y(in_17bit_b[8]) );
  XOR2X1 U119 ( .A(n53), .B(n51), .Y(in_17bit_b[5]) );
  NAND2X1 U120 ( .A(n52), .B(n25), .Y(n51) );
  XOR2X1 U121 ( .A(n60), .B(n58), .Y(in_17bit_b[7]) );
  NAND2X1 U122 ( .A(n59), .B(n25), .Y(n58) );
  XOR2X1 U123 ( .A(n67), .B(n65), .Y(in_17bit_b[9]) );
  INVX1 U124 ( .A(n54), .Y(n57) );
  INVX1 U125 ( .A(n61), .Y(n64) );
  NAND3BX1 U126 ( .AN(n75), .B(n111), .C(n74), .Y(n76) );
  XNOR2X1 U127 ( .A(n69), .B(n70), .Y(in_17bit_b[10]) );
  XOR2X1 U128 ( .A(n74), .B(n72), .Y(in_17bit_b[11]) );
  INVX1 U129 ( .A(n76), .Y(sub_add_52_b0_carry[13]) );
  INVX1 U130 ( .A(n68), .Y(n71) );
  INVX1 U131 ( .A(in_8bit[2]), .Y(n31) );
  NOR2X4 U132 ( .A(in_17bit[1]), .B(in_17bit[0]), .Y(n19) );
  INVX1 U133 ( .A(in_17bit[4]), .Y(n49) );
  INVX1 U134 ( .A(in_17bit[6]), .Y(n56) );
  INVX1 U135 ( .A(in_17bit[5]), .Y(n53) );
  INVX1 U136 ( .A(n47), .Y(n50) );
  NAND2BXL U137 ( .AN(in_17bit[2]), .B(n19), .Y(n44) );
  INVX1 U138 ( .A(in_17bit[16]), .Y(n26) );
  INVX1 U139 ( .A(in_17bit[8]), .Y(n63) );
  INVX1 U140 ( .A(in_17bit[7]), .Y(n60) );
  INVX1 U141 ( .A(in_17bit[10]), .Y(n70) );
  INVX1 U142 ( .A(in_17bit[11]), .Y(n74) );
  INVX1 U143 ( .A(in_17bit[9]), .Y(n67) );
  INVX1 U144 ( .A(in_17bit[12]), .Y(n111) );
  INVX1 U145 ( .A(in_17bit[13]), .Y(n112) );
  INVX1 U146 ( .A(in_17bit[14]), .Y(n113) );
  INVX1 U147 ( .A(in_17bit[15]), .Y(n114) );
  XOR2X1 U148 ( .A(mul[23]), .B(n110), .Y(out[16]) );
  AOI21XL U149 ( .A0(n109), .A1(n108), .B0(n13), .Y(n110) );
  XOR2X2 U150 ( .A(mul[20]), .B(n103), .Y(out[13]) );
  XOR2X2 U151 ( .A(n6), .B(n101), .Y(out[12]) );
  NOR3X4 U152 ( .A(n18), .B(n19), .C(n42), .Y(in_17bit_b[1]) );
  XOR2X4 U153 ( .A(mul[17]), .B(n97), .Y(out[10]) );
  NOR2X4 U154 ( .A(n13), .B(n100), .Y(n99) );
  XNOR2X4 U155 ( .A(n107), .B(n108), .Y(out[15]) );
  XOR2X1 U156 ( .A(n26), .B(sub_add_52_b0_carry[16]), .Y(N21) );
  AND2X1 U157 ( .A(sub_add_52_b0_carry[15]), .B(n114), .Y(
        sub_add_52_b0_carry[16]) );
  XOR2X1 U158 ( .A(n114), .B(sub_add_52_b0_carry[15]), .Y(N20) );
  AND2X1 U159 ( .A(sub_add_52_b0_carry[14]), .B(n113), .Y(
        sub_add_52_b0_carry[15]) );
  XOR2X1 U160 ( .A(n113), .B(sub_add_52_b0_carry[14]), .Y(N19) );
  AND2X1 U161 ( .A(sub_add_52_b0_carry[13]), .B(n112), .Y(
        sub_add_52_b0_carry[14]) );
endmodule


module multi16_6_DW01_add_0 ( A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, 
        A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, 
        B_20_, B_19_, B_18_, B_17_, B_16_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, 
        SUM_17_, SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, 
        SUM_9_, SUM_8_, SUM_7_, SUM_6_, SUM_5_ );
  input A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_,
         A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, B_20_, B_19_,
         B_18_, B_17_, B_16_;
  output SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, SUM_15_,
         SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, SUM_7_,
         SUM_6_, SUM_5_;
  wire   n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39;

  NAND2X2 U2 ( .A(n31), .B(n13), .Y(n37) );
  NOR2X4 U3 ( .A(B_18_), .B(A_18_), .Y(n29) );
  CLKINVX4 U4 ( .A(n18), .Y(SUM_15_) );
  XOR2X2 U5 ( .A(n17), .B(n38), .Y(SUM_17_) );
  CLKINVX4 U6 ( .A(n32), .Y(n17) );
  NOR2X2 U7 ( .A(n28), .B(n15), .Y(n38) );
  BUFX3 U8 ( .A(A_13_), .Y(SUM_13_) );
  BUFX3 U9 ( .A(A_11_), .Y(SUM_11_) );
  NAND2X1 U10 ( .A(B_19_), .B(A_19_), .Y(n27) );
  NOR2X2 U11 ( .A(B_17_), .B(A_17_), .Y(n28) );
  INVX1 U12 ( .A(A_15_), .Y(n18) );
  XOR2X2 U13 ( .A(n34), .B(n35), .Y(SUM_19_) );
  OAI21XL U14 ( .A0(n25), .A1(n26), .B0(n27), .Y(n21) );
  NAND2X4 U15 ( .A(B_17_), .B(A_17_), .Y(n33) );
  INVX4 U16 ( .A(n33), .Y(n15) );
  OAI21X2 U17 ( .A0(n36), .A1(n29), .B0(n31), .Y(n34) );
  AOI21X4 U18 ( .A0(n17), .A1(n16), .B0(n15), .Y(n36) );
  NOR2BX2 U19 ( .AN(n27), .B(n26), .Y(n35) );
  NOR2X1 U20 ( .A(B_19_), .B(A_19_), .Y(n26) );
  XOR2X2 U21 ( .A(n37), .B(n36), .Y(SUM_18_) );
  INVX2 U22 ( .A(n28), .Y(n16) );
  AND2X4 U23 ( .A(n32), .B(n39), .Y(SUM_16_) );
  NAND2X1 U24 ( .A(B_18_), .B(A_18_), .Y(n31) );
  NAND2X2 U25 ( .A(B_16_), .B(A_16_), .Y(n32) );
  INVXL U26 ( .A(n23), .Y(n12) );
  AOI21XL U27 ( .A0(n21), .A1(n22), .B0(n12), .Y(n20) );
  BUFX3 U28 ( .A(A_12_), .Y(SUM_12_) );
  INVX1 U29 ( .A(n31), .Y(n14) );
  BUFX3 U30 ( .A(A_14_), .Y(SUM_14_) );
  BUFX3 U31 ( .A(A_10_), .Y(SUM_10_) );
  BUFX3 U32 ( .A(A_9_), .Y(SUM_9_) );
  BUFX3 U33 ( .A(A_8_), .Y(SUM_8_) );
  BUFX3 U34 ( .A(A_7_), .Y(SUM_7_) );
  BUFX3 U35 ( .A(A_6_), .Y(SUM_6_) );
  BUFX3 U36 ( .A(A_5_), .Y(SUM_5_) );
  INVX1 U37 ( .A(n29), .Y(n13) );
  OR2X2 U38 ( .A(B_16_), .B(A_16_), .Y(n39) );
  XOR2X1 U39 ( .A(n19), .B(n20), .Y(SUM_21_) );
  XNOR2X1 U40 ( .A(B_21_), .B(A_21_), .Y(n19) );
  XNOR2X1 U41 ( .A(n24), .B(n21), .Y(SUM_20_) );
  AOI21X1 U42 ( .A0(n13), .A1(n30), .B0(n14), .Y(n25) );
  OAI21XL U43 ( .A0(n28), .A1(n32), .B0(n33), .Y(n30) );
  NAND2X1 U44 ( .A(n23), .B(n22), .Y(n24) );
  OR2X1 U45 ( .A(B_20_), .B(A_20_), .Y(n22) );
  NAND2X1 U46 ( .A(B_20_), .B(A_20_), .Y(n23) );
endmodule


module multi16_6_DW02_mult_0 ( A, B, PRODUCT_23_, PRODUCT_22_, PRODUCT_21_, 
        PRODUCT_20_, PRODUCT_19_, PRODUCT_18_, PRODUCT_17_, PRODUCT_16_, 
        PRODUCT_15_, PRODUCT_14_, PRODUCT_13_, PRODUCT_12_, PRODUCT_11_, 
        PRODUCT_10_, PRODUCT_9_, PRODUCT_8_, PRODUCT_7_ );
  input [16:0] A;
  input [7:0] B;
  output PRODUCT_23_, PRODUCT_22_, PRODUCT_21_, PRODUCT_20_, PRODUCT_19_,
         PRODUCT_18_, PRODUCT_17_, PRODUCT_16_, PRODUCT_15_, PRODUCT_14_,
         PRODUCT_13_, PRODUCT_12_, PRODUCT_11_, PRODUCT_10_, PRODUCT_9_,
         PRODUCT_8_, PRODUCT_7_;
  wire   ab_16__7_, ab_16__6_, ab_16__5_, ab_16__4_, ab_16__3_, ab_16__2_,
         ab_16__1_, ab_16__0_, ab_15__7_, ab_15__6_, ab_15__5_, ab_15__4_,
         ab_15__3_, ab_15__2_, ab_15__1_, ab_15__0_, ab_14__7_, ab_14__6_,
         ab_14__5_, ab_14__4_, ab_14__3_, ab_14__2_, ab_14__1_, ab_14__0_,
         ab_13__7_, ab_13__6_, ab_13__5_, ab_13__4_, ab_13__3_, ab_13__2_,
         ab_13__1_, ab_13__0_, ab_12__7_, ab_12__6_, ab_12__5_, ab_12__4_,
         ab_12__3_, ab_12__2_, ab_12__1_, ab_12__0_, ab_11__7_, ab_11__6_,
         ab_11__5_, ab_11__4_, ab_11__3_, ab_11__2_, ab_11__1_, ab_11__0_,
         ab_10__7_, ab_10__6_, ab_10__5_, ab_10__4_, ab_10__3_, ab_10__2_,
         ab_10__1_, ab_10__0_, ab_9__7_, ab_9__6_, ab_9__5_, ab_9__4_,
         ab_9__3_, ab_9__2_, ab_9__1_, ab_9__0_, ab_8__7_, ab_8__6_, ab_8__5_,
         ab_8__4_, ab_8__3_, ab_8__2_, ab_8__1_, ab_8__0_, ab_7__7_, ab_7__6_,
         ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_, ab_7__0_, ab_6__7_,
         ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_, ab_6__1_, ab_6__0_,
         ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_, ab_5__2_, ab_5__1_,
         ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_, ab_4__3_, ab_4__2_,
         ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_, ab_3__4_, ab_3__3_,
         ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_, ab_2__5_, ab_2__4_,
         ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_, ab_1__6_, ab_1__5_,
         ab_1__4_, ab_1__3_, ab_1__2_, ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_,
         ab_0__3_, ab_0__2_, CARRYB_16__6_, CARRYB_16__5_, CARRYB_16__4_,
         CARRYB_16__3_, CARRYB_16__2_, CARRYB_16__1_, CARRYB_16__0_,
         CARRYB_15__6_, CARRYB_15__5_, CARRYB_15__4_, CARRYB_15__3_,
         CARRYB_15__2_, CARRYB_15__1_, CARRYB_15__0_, CARRYB_14__6_,
         CARRYB_14__5_, CARRYB_14__4_, CARRYB_14__3_, CARRYB_14__2_,
         CARRYB_14__1_, CARRYB_14__0_, CARRYB_13__6_, CARRYB_13__5_,
         CARRYB_13__4_, CARRYB_13__3_, CARRYB_13__2_, CARRYB_13__1_,
         CARRYB_13__0_, CARRYB_12__6_, CARRYB_12__5_, CARRYB_12__4_,
         CARRYB_12__3_, CARRYB_12__2_, CARRYB_12__1_, CARRYB_12__0_,
         CARRYB_11__6_, CARRYB_11__5_, CARRYB_11__4_, CARRYB_11__3_,
         CARRYB_11__2_, CARRYB_11__1_, CARRYB_11__0_, CARRYB_10__6_,
         CARRYB_10__5_, CARRYB_10__4_, CARRYB_10__3_, CARRYB_10__2_,
         CARRYB_10__1_, CARRYB_10__0_, CARRYB_9__6_, CARRYB_9__5_,
         CARRYB_9__4_, CARRYB_9__3_, CARRYB_9__2_, CARRYB_9__1_, CARRYB_9__0_,
         CARRYB_8__6_, CARRYB_8__5_, CARRYB_8__4_, CARRYB_8__3_, CARRYB_8__2_,
         CARRYB_8__1_, CARRYB_8__0_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_,
         CARRYB_7__3_, CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_,
         CARRYB_6__5_, CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_,
         CARRYB_6__0_, CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_,
         CARRYB_5__2_, CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_,
         CARRYB_4__4_, CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_,
         CARRYB_3__6_, CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_,
         CARRYB_3__1_, CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_,
         CARRYB_2__3_, CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__1_,
         CARRYB_1__0_, SUMB_16__6_, SUMB_16__5_, SUMB_16__4_, SUMB_16__3_,
         SUMB_16__2_, SUMB_16__1_, SUMB_16__0_, SUMB_15__6_, SUMB_15__5_,
         SUMB_15__4_, SUMB_15__3_, SUMB_15__2_, SUMB_15__1_, SUMB_14__6_,
         SUMB_14__5_, SUMB_14__4_, SUMB_14__3_, SUMB_14__2_, SUMB_14__1_,
         SUMB_13__6_, SUMB_13__5_, SUMB_13__4_, SUMB_13__3_, SUMB_13__2_,
         SUMB_13__1_, SUMB_12__6_, SUMB_12__5_, SUMB_12__4_, SUMB_12__3_,
         SUMB_12__2_, SUMB_12__1_, SUMB_11__6_, SUMB_11__5_, SUMB_11__4_,
         SUMB_11__3_, SUMB_11__2_, SUMB_11__1_, SUMB_10__6_, SUMB_10__5_,
         SUMB_10__4_, SUMB_10__3_, SUMB_10__2_, SUMB_10__1_, SUMB_9__6_,
         SUMB_9__5_, SUMB_9__4_, SUMB_9__3_, SUMB_9__2_, SUMB_9__1_,
         SUMB_8__6_, SUMB_8__5_, SUMB_8__4_, SUMB_8__3_, SUMB_8__2_,
         SUMB_8__1_, SUMB_7__6_, SUMB_7__5_, SUMB_7__4_, SUMB_7__3_,
         SUMB_7__2_, SUMB_7__1_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_,
         SUMB_6__3_, SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_,
         SUMB_5__4_, SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_,
         SUMB_4__5_, SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_,
         SUMB_3__6_, SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_,
         SUMB_3__1_, SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_,
         SUMB_2__2_, SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_,
         SUMB_1__3_, SUMB_1__2_, SUMB_1__1_, PROD1_7_, A1_21_, A1_20_, A1_19_,
         A1_18_, A1_17_, A1_16_, A1_15_, A1_13_, A1_12_, A1_11_, A1_10_, A1_9_,
         A1_8_, A1_7_, A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, n3, n4, n5,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57;

  ADDFHX4 S2_15_2 ( .A(ab_15__2_), .B(CARRYB_14__2_), .CI(SUMB_14__3_), .CO(
        CARRYB_15__2_), .S(SUMB_15__2_) );
  ADDFHX4 S1_14_0 ( .A(ab_14__0_), .B(CARRYB_13__0_), .CI(SUMB_13__1_), .CO(
        CARRYB_14__0_), .S(A1_12_) );
  ADDFHX4 S2_14_2 ( .A(ab_14__2_), .B(CARRYB_13__2_), .CI(SUMB_13__3_), .CO(
        CARRYB_14__2_), .S(SUMB_14__2_) );
  ADDFHX4 S1_12_0 ( .A(ab_12__0_), .B(CARRYB_11__0_), .CI(SUMB_11__1_), .CO(
        CARRYB_12__0_), .S(A1_10_) );
  ADDFHX4 S2_12_1 ( .A(ab_12__1_), .B(CARRYB_11__1_), .CI(SUMB_11__2_), .CO(
        CARRYB_12__1_), .S(SUMB_12__1_) );
  ADDFHX4 S1_11_0 ( .A(ab_11__0_), .B(CARRYB_10__0_), .CI(SUMB_10__1_), .CO(
        CARRYB_11__0_), .S(A1_9_) );
  ADDFHX4 S2_11_1 ( .A(ab_11__1_), .B(CARRYB_10__1_), .CI(SUMB_10__2_), .CO(
        CARRYB_11__1_), .S(SUMB_11__1_) );
  ADDFHX4 S2_11_2 ( .A(ab_11__2_), .B(CARRYB_10__2_), .CI(SUMB_10__3_), .CO(
        CARRYB_11__2_), .S(SUMB_11__2_) );
  multi16_6_DW01_add_0 FS_1 ( .A_21_(A1_21_), .A_20_(A1_20_), .A_19_(A1_19_), 
        .A_18_(A1_18_), .A_17_(A1_17_), .A_16_(A1_16_), .A_15_(A1_15_), 
        .A_14_(SUMB_16__0_), .A_13_(A1_13_), .A_12_(A1_12_), .A_11_(A1_11_), 
        .A_10_(A1_10_), .A_9_(A1_9_), .A_8_(A1_8_), .A_7_(A1_7_), .A_6_(A1_6_), 
        .A_5_(PROD1_7_), .B_21_(n12), .B_20_(n39), .B_19_(n38), .B_18_(n35), 
        .B_17_(n36), .B_16_(n37), .SUM_21_(PRODUCT_23_), .SUM_20_(PRODUCT_22_), 
        .SUM_19_(PRODUCT_21_), .SUM_18_(PRODUCT_20_), .SUM_17_(PRODUCT_19_), 
        .SUM_16_(PRODUCT_18_), .SUM_15_(PRODUCT_17_), .SUM_14_(PRODUCT_16_), 
        .SUM_13_(PRODUCT_15_), .SUM_12_(PRODUCT_14_), .SUM_11_(PRODUCT_13_), 
        .SUM_10_(PRODUCT_12_), .SUM_9_(PRODUCT_11_), .SUM_8_(PRODUCT_10_), 
        .SUM_7_(PRODUCT_9_), .SUM_6_(PRODUCT_8_), .SUM_5_(PRODUCT_7_) );
  ADDFHX1 S3_11_6 ( .A(ab_11__6_), .B(CARRYB_10__6_), .CI(ab_10__7_), .CO(
        CARRYB_11__6_), .S(SUMB_11__6_) );
  ADDFHX1 S3_14_6 ( .A(ab_14__6_), .B(CARRYB_13__6_), .CI(ab_13__7_), .CO(
        CARRYB_14__6_), .S(SUMB_14__6_) );
  ADDFX2 S3_15_6 ( .A(ab_15__6_), .B(CARRYB_14__6_), .CI(ab_14__7_), .CO(
        CARRYB_15__6_), .S(SUMB_15__6_) );
  ADDFHX1 S2_15_5 ( .A(ab_15__5_), .B(CARRYB_14__5_), .CI(SUMB_14__6_), .CO(
        CARRYB_15__5_), .S(SUMB_15__5_) );
  ADDFX2 S5_6 ( .A(ab_16__6_), .B(CARRYB_15__6_), .CI(ab_15__7_), .CO(
        CARRYB_16__6_), .S(SUMB_16__6_) );
  ADDFHX2 S3_2_6 ( .A(ab_2__6_), .B(n10), .CI(ab_1__7_), .CO(CARRYB_2__6_), 
        .S(SUMB_2__6_) );
  ADDFHX2 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  ADDFHX4 S2_15_3 ( .A(ab_15__3_), .B(CARRYB_14__3_), .CI(SUMB_14__4_), .CO(
        CARRYB_15__3_), .S(SUMB_15__3_) );
  ADDFHX2 S2_7_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  ADDFHX2 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  ADDFHX4 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  ADDFHX4 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  ADDFHX2 S2_11_5 ( .A(ab_11__5_), .B(CARRYB_10__5_), .CI(SUMB_10__6_), .CO(
        CARRYB_11__5_), .S(SUMB_11__5_) );
  ADDFHX2 S3_10_6 ( .A(ab_10__6_), .B(CARRYB_9__6_), .CI(ab_9__7_), .CO(
        CARRYB_10__6_), .S(SUMB_10__6_) );
  ADDFHX4 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  ADDFHX2 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  ADDFHX4 S1_9_0 ( .A(ab_9__0_), .B(CARRYB_8__0_), .CI(SUMB_8__1_), .CO(
        CARRYB_9__0_), .S(A1_7_) );
  ADDFHX4 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  ADDFHX4 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  ADDFHX4 S2_10_2 ( .A(ab_10__2_), .B(CARRYB_9__2_), .CI(SUMB_9__3_), .CO(
        CARRYB_10__2_), .S(SUMB_10__2_) );
  ADDFHX4 S2_11_3 ( .A(ab_11__3_), .B(CARRYB_10__3_), .CI(SUMB_10__4_), .CO(
        CARRYB_11__3_), .S(SUMB_11__3_) );
  ADDFHX4 S3_7_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(
        CARRYB_7__6_), .S(SUMB_7__6_) );
  ADDFHX4 S3_8_6 ( .A(ab_8__6_), .B(CARRYB_7__6_), .CI(ab_7__7_), .CO(
        CARRYB_8__6_), .S(SUMB_8__6_) );
  ADDFHX4 S1_8_0 ( .A(ab_8__0_), .B(CARRYB_7__0_), .CI(SUMB_7__1_), .CO(
        CARRYB_8__0_), .S(A1_6_) );
  ADDFHX4 S2_8_2 ( .A(ab_8__2_), .B(CARRYB_7__2_), .CI(SUMB_7__3_), .CO(
        CARRYB_8__2_), .S(SUMB_8__2_) );
  ADDFHX2 S2_10_4 ( .A(ab_10__4_), .B(CARRYB_9__4_), .CI(SUMB_9__5_), .CO(
        CARRYB_10__4_), .S(SUMB_10__4_) );
  ADDFHX2 S2_11_4 ( .A(ab_11__4_), .B(CARRYB_10__4_), .CI(SUMB_10__5_), .CO(
        CARRYB_11__4_), .S(SUMB_11__4_) );
  ADDFHX2 S2_2_3 ( .A(ab_2__3_), .B(n7), .CI(SUMB_1__4_), .CO(CARRYB_2__3_), 
        .S(SUMB_2__3_) );
  ADDFHX4 S2_13_3 ( .A(ab_13__3_), .B(CARRYB_12__3_), .CI(SUMB_12__4_), .CO(
        CARRYB_13__3_), .S(SUMB_13__3_) );
  ADDFHX4 S2_9_2 ( .A(ab_9__2_), .B(CARRYB_8__2_), .CI(SUMB_8__3_), .CO(
        CARRYB_9__2_), .S(SUMB_9__2_) );
  ADDFHX4 S2_7_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  ADDFHX2 S2_15_4 ( .A(ab_15__4_), .B(CARRYB_14__4_), .CI(SUMB_14__5_), .CO(
        CARRYB_15__4_), .S(SUMB_15__4_) );
  ADDFHX4 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  ADDFHX4 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  ADDFHX2 S4_1 ( .A(ab_16__1_), .B(CARRYB_15__1_), .CI(SUMB_15__2_), .CO(
        CARRYB_16__1_), .S(SUMB_16__1_) );
  ADDFHX4 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  ADDFHX4 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  ADDFHX2 S2_2_2 ( .A(ab_2__2_), .B(n8), .CI(SUMB_1__3_), .CO(CARRYB_2__2_), 
        .S(SUMB_2__2_) );
  ADDFHX4 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  ADDFHX2 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  ADDFHX4 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  ADDFHX2 S3_12_6 ( .A(ab_12__6_), .B(CARRYB_11__6_), .CI(ab_11__7_), .CO(
        CARRYB_12__6_), .S(SUMB_12__6_) );
  ADDFHX2 S3_13_6 ( .A(ab_13__6_), .B(CARRYB_12__6_), .CI(ab_12__7_), .CO(
        CARRYB_13__6_), .S(SUMB_13__6_) );
  ADDFHX4 S3_9_6 ( .A(ab_9__6_), .B(CARRYB_8__6_), .CI(ab_8__7_), .CO(
        CARRYB_9__6_), .S(SUMB_9__6_) );
  ADDFHX4 S2_8_3 ( .A(ab_8__3_), .B(CARRYB_7__3_), .CI(SUMB_7__4_), .CO(
        CARRYB_8__3_), .S(SUMB_8__3_) );
  ADDFHX4 S2_14_3 ( .A(ab_14__3_), .B(CARRYB_13__3_), .CI(SUMB_13__4_), .CO(
        CARRYB_14__3_), .S(SUMB_14__3_) );
  ADDFHX2 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  ADDFHX4 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  ADDFHX4 S2_8_1 ( .A(ab_8__1_), .B(CARRYB_7__1_), .CI(SUMB_7__2_), .CO(
        CARRYB_8__1_), .S(SUMB_8__1_) );
  ADDFHX4 S2_14_4 ( .A(ab_14__4_), .B(CARRYB_13__4_), .CI(SUMB_13__5_), .CO(
        CARRYB_14__4_), .S(SUMB_14__4_) );
  ADDFHX2 S2_12_5 ( .A(ab_12__5_), .B(CARRYB_11__5_), .CI(SUMB_11__6_), .CO(
        CARRYB_12__5_), .S(SUMB_12__5_) );
  ADDFHX2 S4_5 ( .A(ab_16__5_), .B(CARRYB_15__5_), .CI(SUMB_15__6_), .CO(
        CARRYB_16__5_), .S(SUMB_16__5_) );
  ADDFHX1 S2_2_4 ( .A(ab_2__4_), .B(n11), .CI(SUMB_1__5_), .CO(CARRYB_2__4_), 
        .S(SUMB_2__4_) );
  ADDFHX2 S2_2_5 ( .A(ab_2__5_), .B(n9), .CI(SUMB_1__6_), .CO(CARRYB_2__5_), 
        .S(SUMB_2__5_) );
  ADDFHX2 S4_2 ( .A(ab_16__2_), .B(CARRYB_15__2_), .CI(SUMB_15__3_), .CO(
        CARRYB_16__2_), .S(SUMB_16__2_) );
  ADDFHX2 S4_3 ( .A(ab_16__3_), .B(CARRYB_15__3_), .CI(SUMB_15__4_), .CO(
        CARRYB_16__3_), .S(SUMB_16__3_) );
  ADDFHX1 S2_13_5 ( .A(ab_13__5_), .B(CARRYB_12__5_), .CI(SUMB_12__6_), .CO(
        CARRYB_13__5_), .S(SUMB_13__5_) );
  ADDFHX2 S1_13_0 ( .A(ab_13__0_), .B(CARRYB_12__0_), .CI(SUMB_12__1_), .CO(
        CARRYB_13__0_), .S(A1_11_) );
  ADDFHX2 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  ADDFHX2 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  ADDFHX2 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  ADDFHX2 S2_13_1 ( .A(ab_13__1_), .B(CARRYB_12__1_), .CI(SUMB_12__2_), .CO(
        CARRYB_13__1_), .S(SUMB_13__1_) );
  ADDFHX2 S2_7_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  ADDFHX2 S2_12_3 ( .A(ab_12__3_), .B(CARRYB_11__3_), .CI(SUMB_11__4_), .CO(
        CARRYB_12__3_), .S(SUMB_12__3_) );
  ADDFHX2 S2_7_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  ADDFHX1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  ADDFHX2 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  ADDFHX1 S2_14_5 ( .A(ab_14__5_), .B(CARRYB_13__5_), .CI(SUMB_13__6_), .CO(
        CARRYB_14__5_), .S(SUMB_14__5_) );
  ADDFHX2 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  ADDFHX4 S2_12_4 ( .A(ab_12__4_), .B(CARRYB_11__4_), .CI(SUMB_11__5_), .CO(
        CARRYB_12__4_), .S(SUMB_12__4_) );
  ADDFHX4 S2_13_4 ( .A(ab_13__4_), .B(CARRYB_12__4_), .CI(SUMB_12__5_), .CO(
        CARRYB_13__4_), .S(SUMB_13__4_) );
  ADDFHX4 S2_8_4 ( .A(ab_8__4_), .B(CARRYB_7__4_), .CI(SUMB_7__5_), .CO(
        CARRYB_8__4_), .S(SUMB_8__4_) );
  ADDFHX4 S2_9_4 ( .A(ab_9__4_), .B(CARRYB_8__4_), .CI(SUMB_8__5_), .CO(
        CARRYB_9__4_), .S(SUMB_9__4_) );
  ADDFHX4 S2_9_5 ( .A(ab_9__5_), .B(CARRYB_8__5_), .CI(SUMB_8__6_), .CO(
        CARRYB_9__5_), .S(SUMB_9__5_) );
  ADDFHX4 S2_10_5 ( .A(ab_10__5_), .B(CARRYB_9__5_), .CI(SUMB_9__6_), .CO(
        CARRYB_10__5_), .S(SUMB_10__5_) );
  ADDFHX2 S2_10_3 ( .A(ab_10__3_), .B(CARRYB_9__3_), .CI(SUMB_9__4_), .CO(
        CARRYB_10__3_), .S(SUMB_10__3_) );
  ADDFHX4 S2_10_1 ( .A(ab_10__1_), .B(CARRYB_9__1_), .CI(SUMB_9__2_), .CO(
        CARRYB_10__1_), .S(SUMB_10__1_) );
  ADDFHX4 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  ADDFHX4 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  ADDFHX4 S2_14_1 ( .A(ab_14__1_), .B(CARRYB_13__1_), .CI(SUMB_13__2_), .CO(
        CARRYB_14__1_), .S(SUMB_14__1_) );
  ADDFHX4 S2_15_1 ( .A(ab_15__1_), .B(CARRYB_14__1_), .CI(SUMB_14__2_), .CO(
        CARRYB_15__1_), .S(SUMB_15__1_) );
  ADDFHX4 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  ADDFHX4 S1_7_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(PROD1_7_) );
  ADDFHX2 S2_9_1 ( .A(ab_9__1_), .B(CARRYB_8__1_), .CI(SUMB_8__2_), .CO(
        CARRYB_9__1_), .S(SUMB_9__1_) );
  ADDFHX4 S1_10_0 ( .A(ab_10__0_), .B(CARRYB_9__0_), .CI(SUMB_9__1_), .CO(
        CARRYB_10__0_), .S(A1_8_) );
  ADDFHX4 S1_15_0 ( .A(ab_15__0_), .B(CARRYB_14__0_), .CI(SUMB_14__1_), .CO(
        CARRYB_15__0_), .S(A1_13_) );
  ADDFHX2 S4_0 ( .A(ab_16__0_), .B(CARRYB_15__0_), .CI(SUMB_15__1_), .CO(
        CARRYB_16__0_), .S(SUMB_16__0_) );
  ADDFHX2 S4_4 ( .A(ab_16__4_), .B(CARRYB_15__4_), .CI(SUMB_15__5_), .CO(
        CARRYB_16__4_), .S(SUMB_16__4_) );
  ADDFHX4 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  ADDFHX4 S2_8_5 ( .A(ab_8__5_), .B(CARRYB_7__5_), .CI(SUMB_7__6_), .CO(
        CARRYB_8__5_), .S(SUMB_8__5_) );
  CLKINVX8 U2 ( .A(n30), .Y(CARRYB_1__1_) );
  XOR3X2 U3 ( .A(n50), .B(1'b0), .C(ab_0__2_), .Y(SUMB_1__1_) );
  NAND2X2 U4 ( .A(A[1]), .B(B[1]), .Y(n42) );
  XOR3X2 U5 ( .A(CARRYB_8__3_), .B(ab_9__3_), .C(SUMB_8__4_), .Y(SUMB_9__3_)
         );
  NAND2X2 U6 ( .A(SUMB_8__4_), .B(CARRYB_8__3_), .Y(n3) );
  NAND2X2 U7 ( .A(ab_9__3_), .B(CARRYB_8__3_), .Y(n4) );
  NAND2X2 U8 ( .A(ab_9__3_), .B(SUMB_8__4_), .Y(n5) );
  NAND3X2 U9 ( .A(n5), .B(n3), .C(n4), .Y(CARRYB_9__3_) );
  AND2X2 U10 ( .A(A[4]), .B(B[5]), .Y(ab_4__5_) );
  INVX4 U11 ( .A(B[3]), .Y(n46) );
  AND2X2 U12 ( .A(A[1]), .B(B[3]), .Y(ab_1__3_) );
  AND2X2 U13 ( .A(A[2]), .B(B[3]), .Y(ab_2__3_) );
  INVX4 U14 ( .A(B[7]), .Y(n49) );
  NOR2X4 U15 ( .A(n43), .B(n40), .Y(ab_0__6_) );
  INVX4 U16 ( .A(B[6]), .Y(n43) );
  NOR2XL U17 ( .A(n56), .B(n46), .Y(ab_11__3_) );
  NAND3X2 U18 ( .A(n25), .B(n23), .C(n24), .Y(CARRYB_6__3_) );
  NOR2X1 U19 ( .A(n47), .B(n40), .Y(ab_0__2_) );
  CLKINVX3 U20 ( .A(n42), .Y(n50) );
  INVX1 U21 ( .A(B[4]), .Y(n45) );
  XOR2X2 U22 ( .A(CARRYB_16__1_), .B(SUMB_16__2_), .Y(A1_16_) );
  XOR2X2 U23 ( .A(CARRYB_16__2_), .B(SUMB_16__3_), .Y(A1_17_) );
  AND2X2 U24 ( .A(A[4]), .B(B[6]), .Y(ab_4__6_) );
  NAND2X1 U25 ( .A(ab_6__3_), .B(CARRYB_5__3_), .Y(n25) );
  NAND2X1 U26 ( .A(CARRYB_5__3_), .B(SUMB_5__4_), .Y(n23) );
  INVX1 U27 ( .A(A[0]), .Y(n40) );
  XOR3X2 U28 ( .A(SUMB_5__4_), .B(ab_6__3_), .C(CARRYB_5__3_), .Y(SUMB_6__3_)
         );
  NAND2X1 U29 ( .A(ab_0__2_), .B(n50), .Y(n30) );
  NOR2X1 U30 ( .A(n46), .B(n40), .Y(ab_0__3_) );
  XOR2X1 U31 ( .A(CARRYB_16__0_), .B(SUMB_16__1_), .Y(A1_15_) );
  AND2X2 U33 ( .A(ab_0__4_), .B(ab_1__3_), .Y(n7) );
  AND2X2 U34 ( .A(ab_0__3_), .B(ab_1__2_), .Y(n8) );
  AND2X2 U35 ( .A(ab_0__6_), .B(ab_1__5_), .Y(n9) );
  AND2X2 U36 ( .A(ab_0__7_), .B(ab_1__6_), .Y(n10) );
  AND2X2 U37 ( .A(ab_0__5_), .B(ab_1__4_), .Y(n11) );
  AND2X2 U38 ( .A(CARRYB_16__5_), .B(SUMB_16__6_), .Y(n12) );
  AND2X2 U39 ( .A(A[2]), .B(B[5]), .Y(ab_2__5_) );
  NAND3X2 U40 ( .A(n17), .B(n18), .C(n19), .Y(CARRYB_13__2_) );
  XOR3X2 U41 ( .A(ab_12__2_), .B(CARRYB_11__2_), .C(SUMB_11__3_), .Y(
        SUMB_12__2_) );
  NAND2X1 U42 ( .A(ab_12__2_), .B(CARRYB_11__2_), .Y(n13) );
  NAND2X1 U43 ( .A(ab_12__2_), .B(SUMB_11__3_), .Y(n14) );
  NAND2X1 U44 ( .A(CARRYB_11__2_), .B(SUMB_11__3_), .Y(n15) );
  NAND3X1 U45 ( .A(n13), .B(n14), .C(n15), .Y(CARRYB_12__2_) );
  XOR2X2 U46 ( .A(ab_13__2_), .B(SUMB_12__3_), .Y(n16) );
  XOR2X1 U47 ( .A(n16), .B(CARRYB_12__2_), .Y(SUMB_13__2_) );
  NAND2X1 U48 ( .A(ab_13__2_), .B(SUMB_12__3_), .Y(n17) );
  NAND2X1 U49 ( .A(ab_13__2_), .B(CARRYB_12__2_), .Y(n18) );
  NAND2X1 U50 ( .A(SUMB_12__3_), .B(CARRYB_12__2_), .Y(n19) );
  XOR3X2 U51 ( .A(ab_3__4_), .B(SUMB_2__5_), .C(CARRYB_2__4_), .Y(SUMB_3__4_)
         );
  NAND2X1 U52 ( .A(CARRYB_2__4_), .B(ab_3__4_), .Y(n20) );
  NAND2XL U53 ( .A(SUMB_2__5_), .B(ab_3__4_), .Y(n21) );
  NAND2X1 U54 ( .A(SUMB_2__5_), .B(CARRYB_2__4_), .Y(n22) );
  NAND3X2 U55 ( .A(n22), .B(n20), .C(n21), .Y(CARRYB_3__4_) );
  AND2X2 U56 ( .A(A[3]), .B(B[2]), .Y(ab_3__2_) );
  AND2X4 U57 ( .A(CARRYB_16__1_), .B(SUMB_16__2_), .Y(n36) );
  NAND3X2 U58 ( .A(n34), .B(n32), .C(n33), .Y(CARRYB_7__4_) );
  NAND2X1 U59 ( .A(ab_7__4_), .B(SUMB_6__5_), .Y(n34) );
  XOR2X2 U60 ( .A(CARRYB_6__4_), .B(n31), .Y(SUMB_7__4_) );
  AND2X2 U61 ( .A(A[3]), .B(B[6]), .Y(ab_3__6_) );
  AND2X2 U62 ( .A(A[3]), .B(B[5]), .Y(ab_3__5_) );
  INVX2 U63 ( .A(B[5]), .Y(n44) );
  XOR2X2 U64 ( .A(CARRYB_16__4_), .B(SUMB_16__5_), .Y(A1_19_) );
  NAND3X4 U65 ( .A(n29), .B(n27), .C(n28), .Y(CARRYB_4__6_) );
  NAND2X2 U66 ( .A(ab_4__6_), .B(CARRYB_3__6_), .Y(n27) );
  NAND2X2 U67 ( .A(ab_3__7_), .B(CARRYB_3__6_), .Y(n28) );
  XOR2X2 U68 ( .A(CARRYB_16__3_), .B(SUMB_16__4_), .Y(A1_18_) );
  NAND2X2 U69 ( .A(ab_6__3_), .B(SUMB_5__4_), .Y(n24) );
  XOR2X1 U70 ( .A(ab_4__6_), .B(ab_3__7_), .Y(n26) );
  XOR2X1 U71 ( .A(CARRYB_3__6_), .B(n26), .Y(SUMB_4__6_) );
  NAND2XL U72 ( .A(ab_3__7_), .B(ab_4__6_), .Y(n29) );
  XOR2X4 U73 ( .A(SUMB_6__5_), .B(ab_7__4_), .Y(n31) );
  NAND2X1 U74 ( .A(SUMB_6__5_), .B(CARRYB_6__4_), .Y(n32) );
  NAND2X1 U75 ( .A(ab_7__4_), .B(CARRYB_6__4_), .Y(n33) );
  NOR2XL U76 ( .A(n55), .B(n43), .Y(ab_12__6_) );
  NOR2XL U77 ( .A(n52), .B(n43), .Y(ab_15__6_) );
  NOR2XL U78 ( .A(n45), .B(n40), .Y(ab_0__4_) );
  INVX2 U79 ( .A(B[2]), .Y(n47) );
  AND2X1 U80 ( .A(A[3]), .B(B[3]), .Y(ab_3__3_) );
  AND2X1 U81 ( .A(A[10]), .B(B[1]), .Y(ab_10__1_) );
  AND2X1 U82 ( .A(A[8]), .B(B[0]), .Y(ab_8__0_) );
  AND2X1 U83 ( .A(A[9]), .B(B[1]), .Y(ab_9__1_) );
  AND2X1 U84 ( .A(A[8]), .B(B[1]), .Y(ab_8__1_) );
  AND2X1 U85 ( .A(A[6]), .B(B[1]), .Y(ab_6__1_) );
  AND2X1 U86 ( .A(A[10]), .B(B[0]), .Y(ab_10__0_) );
  AND2X1 U87 ( .A(A[7]), .B(B[0]), .Y(ab_7__0_) );
  AND2X1 U88 ( .A(A[6]), .B(B[0]), .Y(ab_6__0_) );
  INVXL U89 ( .A(B[0]), .Y(n57) );
  INVXL U90 ( .A(B[1]), .Y(n48) );
  NOR2XL U91 ( .A(n53), .B(n43), .Y(ab_14__6_) );
  NOR2XL U92 ( .A(n56), .B(n48), .Y(ab_11__1_) );
  NOR2XL U93 ( .A(n54), .B(n43), .Y(ab_13__6_) );
  AND2X1 U94 ( .A(A[5]), .B(B[0]), .Y(ab_5__0_) );
  AND2X1 U95 ( .A(A[4]), .B(B[0]), .Y(ab_4__0_) );
  AND2X1 U96 ( .A(A[2]), .B(B[0]), .Y(ab_2__0_) );
  AND2X1 U97 ( .A(A[2]), .B(B[4]), .Y(ab_2__4_) );
  AND2X1 U98 ( .A(A[7]), .B(B[6]), .Y(ab_7__6_) );
  AND2X1 U99 ( .A(A[5]), .B(B[6]), .Y(ab_5__6_) );
  AND2X1 U100 ( .A(A[2]), .B(B[1]), .Y(ab_2__1_) );
  AND2X1 U101 ( .A(CARRYB_16__2_), .B(SUMB_16__3_), .Y(n35) );
  AND2X2 U102 ( .A(CARRYB_16__0_), .B(SUMB_16__1_), .Y(n37) );
  NOR2X1 U103 ( .A(n51), .B(n48), .Y(ab_16__1_) );
  NOR2XL U104 ( .A(n51), .B(n47), .Y(ab_16__2_) );
  NOR2X1 U105 ( .A(n51), .B(n46), .Y(ab_16__3_) );
  NOR2X1 U106 ( .A(n51), .B(n44), .Y(ab_16__5_) );
  AND2X2 U107 ( .A(A[7]), .B(B[1]), .Y(ab_7__1_) );
  AND2X2 U108 ( .A(A[9]), .B(B[0]), .Y(ab_9__0_) );
  AND2X2 U109 ( .A(A[5]), .B(B[1]), .Y(ab_5__1_) );
  AND2X2 U110 ( .A(A[4]), .B(B[1]), .Y(ab_4__1_) );
  XOR2X1 U111 ( .A(CARRYB_16__5_), .B(SUMB_16__6_), .Y(A1_20_) );
  XOR2X1 U112 ( .A(CARRYB_16__6_), .B(ab_16__7_), .Y(A1_21_) );
  AND2X2 U113 ( .A(CARRYB_16__3_), .B(SUMB_16__4_), .Y(n38) );
  AND2X1 U114 ( .A(CARRYB_16__4_), .B(SUMB_16__5_), .Y(n39) );
  NOR2X1 U115 ( .A(n44), .B(n40), .Y(ab_0__5_) );
  NOR2X1 U116 ( .A(n49), .B(n40), .Y(ab_0__7_) );
  NOR2XL U117 ( .A(n51), .B(n45), .Y(ab_16__4_) );
  NOR2XL U118 ( .A(n52), .B(n49), .Y(ab_15__7_) );
  NOR2X1 U119 ( .A(n51), .B(n43), .Y(ab_16__6_) );
  AND2X1 U120 ( .A(A[1]), .B(B[2]), .Y(ab_1__2_) );
  NOR2X1 U121 ( .A(n53), .B(n48), .Y(ab_14__1_) );
  NOR2X1 U122 ( .A(n54), .B(n48), .Y(ab_13__1_) );
  NOR2X1 U123 ( .A(n55), .B(n48), .Y(ab_12__1_) );
  NOR2XL U124 ( .A(n53), .B(n47), .Y(ab_14__2_) );
  NOR2XL U125 ( .A(n54), .B(n47), .Y(ab_13__2_) );
  NOR2XL U126 ( .A(n55), .B(n47), .Y(ab_12__2_) );
  NOR2XL U127 ( .A(n52), .B(n47), .Y(ab_15__2_) );
  NOR2XL U128 ( .A(n56), .B(n47), .Y(ab_11__2_) );
  NOR2XL U129 ( .A(n54), .B(n46), .Y(ab_13__3_) );
  NOR2XL U130 ( .A(n52), .B(n46), .Y(ab_15__3_) );
  NOR2XL U131 ( .A(n55), .B(n46), .Y(ab_12__3_) );
  NOR2XL U132 ( .A(n53), .B(n46), .Y(ab_14__3_) );
  AND2X1 U133 ( .A(A[10]), .B(B[3]), .Y(ab_10__3_) );
  AND2X1 U134 ( .A(A[9]), .B(B[3]), .Y(ab_9__3_) );
  AND2X1 U135 ( .A(A[8]), .B(B[3]), .Y(ab_8__3_) );
  NOR2XL U136 ( .A(n53), .B(n45), .Y(ab_14__4_) );
  NOR2XL U137 ( .A(n55), .B(n45), .Y(ab_12__4_) );
  NOR2XL U138 ( .A(n56), .B(n45), .Y(ab_11__4_) );
  NOR2XL U139 ( .A(n54), .B(n45), .Y(ab_13__4_) );
  AND2X1 U140 ( .A(A[7]), .B(B[3]), .Y(ab_7__3_) );
  AND2X1 U141 ( .A(A[6]), .B(B[3]), .Y(ab_6__3_) );
  AND2X1 U142 ( .A(A[3]), .B(B[1]), .Y(ab_3__1_) );
  NOR2XL U143 ( .A(n54), .B(n44), .Y(ab_13__5_) );
  NOR2XL U144 ( .A(n56), .B(n44), .Y(ab_11__5_) );
  NOR2XL U145 ( .A(n55), .B(n44), .Y(ab_12__5_) );
  AND2X1 U146 ( .A(A[10]), .B(B[5]), .Y(ab_10__5_) );
  AND2X1 U147 ( .A(A[5]), .B(B[3]), .Y(ab_5__3_) );
  AND2X1 U148 ( .A(A[9]), .B(B[5]), .Y(ab_9__5_) );
  AND2X1 U149 ( .A(A[8]), .B(B[5]), .Y(ab_8__5_) );
  AND2X1 U150 ( .A(A[7]), .B(B[5]), .Y(ab_7__5_) );
  AND2X1 U151 ( .A(A[6]), .B(B[5]), .Y(ab_6__5_) );
  AND2X1 U152 ( .A(A[4]), .B(B[3]), .Y(ab_4__3_) );
  AND2X1 U153 ( .A(A[5]), .B(B[5]), .Y(ab_5__5_) );
  NOR2XL U154 ( .A(n56), .B(n49), .Y(ab_11__7_) );
  XOR2X1 U155 ( .A(ab_1__4_), .B(ab_0__5_), .Y(SUMB_1__4_) );
  XOR2X1 U156 ( .A(ab_1__3_), .B(ab_0__4_), .Y(SUMB_1__3_) );
  XOR2X1 U157 ( .A(ab_1__6_), .B(ab_0__7_), .Y(SUMB_1__6_) );
  NOR2X1 U158 ( .A(n52), .B(n48), .Y(ab_15__1_) );
  NOR2XL U159 ( .A(n52), .B(n45), .Y(ab_15__4_) );
  NOR2XL U160 ( .A(n53), .B(n44), .Y(ab_14__5_) );
  NOR2XL U161 ( .A(n52), .B(n44), .Y(ab_15__5_) );
  NOR2XL U162 ( .A(n53), .B(n49), .Y(ab_14__7_) );
  NOR2XL U163 ( .A(n55), .B(n49), .Y(ab_12__7_) );
  NOR2XL U164 ( .A(n54), .B(n49), .Y(ab_13__7_) );
  INVX1 U165 ( .A(A[16]), .Y(n51) );
  NOR2XL U166 ( .A(n51), .B(n49), .Y(ab_16__7_) );
  AND2X1 U167 ( .A(A[10]), .B(B[4]), .Y(ab_10__4_) );
  AND2X1 U168 ( .A(A[9]), .B(B[4]), .Y(ab_9__4_) );
  AND2X1 U169 ( .A(A[8]), .B(B[4]), .Y(ab_8__4_) );
  AND2X1 U170 ( .A(A[7]), .B(B[4]), .Y(ab_7__4_) );
  AND2X1 U171 ( .A(A[6]), .B(B[4]), .Y(ab_6__4_) );
  XOR2X1 U172 ( .A(ab_1__2_), .B(ab_0__3_), .Y(SUMB_1__2_) );
  AND2X1 U173 ( .A(A[5]), .B(B[4]), .Y(ab_5__4_) );
  AND2X1 U174 ( .A(A[3]), .B(B[4]), .Y(ab_3__4_) );
  AND2X1 U175 ( .A(A[4]), .B(B[4]), .Y(ab_4__4_) );
  AND2X2 U176 ( .A(A[3]), .B(B[0]), .Y(ab_3__0_) );
  NOR2X1 U177 ( .A(n42), .B(n41), .Y(CARRYB_1__0_) );
  AND2X2 U178 ( .A(A[10]), .B(B[6]), .Y(ab_10__6_) );
  AND2X1 U179 ( .A(A[2]), .B(B[7]), .Y(ab_2__7_) );
  NOR2XL U180 ( .A(n56), .B(n43), .Y(ab_11__6_) );
  AND2X2 U181 ( .A(A[9]), .B(B[6]), .Y(ab_9__6_) );
  AND2X2 U182 ( .A(A[8]), .B(B[6]), .Y(ab_8__6_) );
  AND2X2 U183 ( .A(A[6]), .B(B[6]), .Y(ab_6__6_) );
  XOR2X1 U184 ( .A(ab_1__5_), .B(ab_0__6_), .Y(SUMB_1__5_) );
  AND2X1 U185 ( .A(A[2]), .B(B[6]), .Y(ab_2__6_) );
  NAND2XL U186 ( .A(A[0]), .B(B[0]), .Y(n41) );
  INVX1 U187 ( .A(A[11]), .Y(n56) );
  INVX1 U188 ( .A(A[12]), .Y(n55) );
  INVX1 U189 ( .A(A[13]), .Y(n54) );
  INVX1 U190 ( .A(A[14]), .Y(n53) );
  INVX1 U191 ( .A(A[15]), .Y(n52) );
  AND2X2 U192 ( .A(A[1]), .B(B[6]), .Y(ab_1__6_) );
  AND2X1 U193 ( .A(A[10]), .B(B[2]), .Y(ab_10__2_) );
  AND2X1 U194 ( .A(A[9]), .B(B[2]), .Y(ab_9__2_) );
  AND2X1 U195 ( .A(A[8]), .B(B[2]), .Y(ab_8__2_) );
  AND2X1 U196 ( .A(A[7]), .B(B[2]), .Y(ab_7__2_) );
  AND2X1 U197 ( .A(A[6]), .B(B[2]), .Y(ab_6__2_) );
  AND2X1 U198 ( .A(A[5]), .B(B[2]), .Y(ab_5__2_) );
  AND2X1 U199 ( .A(A[4]), .B(B[2]), .Y(ab_4__2_) );
  AND2X1 U200 ( .A(A[2]), .B(B[2]), .Y(ab_2__2_) );
  AND2X1 U201 ( .A(A[1]), .B(B[7]), .Y(ab_1__7_) );
  AND2X2 U202 ( .A(A[1]), .B(B[5]), .Y(ab_1__5_) );
  AND2X2 U203 ( .A(A[1]), .B(B[4]), .Y(ab_1__4_) );
  AND2X1 U204 ( .A(A[10]), .B(B[7]), .Y(ab_10__7_) );
  AND2X1 U205 ( .A(A[9]), .B(B[7]), .Y(ab_9__7_) );
  AND2X1 U206 ( .A(A[8]), .B(B[7]), .Y(ab_8__7_) );
  AND2X1 U207 ( .A(A[7]), .B(B[7]), .Y(ab_7__7_) );
  AND2X1 U208 ( .A(A[6]), .B(B[7]), .Y(ab_6__7_) );
  AND2X1 U209 ( .A(A[5]), .B(B[7]), .Y(ab_5__7_) );
  AND2X1 U210 ( .A(A[4]), .B(B[7]), .Y(ab_4__7_) );
  AND2X1 U211 ( .A(A[3]), .B(B[7]), .Y(ab_3__7_) );
  NOR2X1 U213 ( .A(n57), .B(n51), .Y(ab_16__0_) );
  NOR2X1 U214 ( .A(n57), .B(n52), .Y(ab_15__0_) );
  NOR2X1 U215 ( .A(n57), .B(n53), .Y(ab_14__0_) );
  NOR2X1 U216 ( .A(n57), .B(n54), .Y(ab_13__0_) );
  NOR2X1 U217 ( .A(n57), .B(n55), .Y(ab_12__0_) );
  NOR2X1 U218 ( .A(n57), .B(n56), .Y(ab_11__0_) );
endmodule


module multi16_6 ( in_17bit, in_8bit, out );
  input [16:0] in_17bit;
  input [7:0] in_8bit;
  output [16:0] out;
  wire   N18, N19, N20, N21, N32, N33, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n55, n56, n57, n58, n59, n60, n61, n63, n64, n65, n66, n67, n68,
         n69, n71, n72, n73, n74, n75, n76, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n116, n117, n118, n119;
  wire   [16:1] in_17bit_b;
  wire   [7:0] in_8bit_b;
  wire   [23:8] mul;
  wire   [16:12] sub_add_52_b0_carry;

  multi16_6_DW02_mult_0 mult_55 ( .A({in_17bit_b, in_17bit[0]}), .B(in_8bit_b), 
        .PRODUCT_23_(mul[23]), .PRODUCT_22_(mul[22]), .PRODUCT_21_(mul[21]), 
        .PRODUCT_20_(mul[20]), .PRODUCT_19_(mul[19]), .PRODUCT_18_(mul[18]), 
        .PRODUCT_17_(mul[17]), .PRODUCT_16_(mul[16]), .PRODUCT_15_(mul[15]), 
        .PRODUCT_14_(mul[14]), .PRODUCT_13_(mul[13]), .PRODUCT_12_(mul[12]), 
        .PRODUCT_11_(mul[11]), .PRODUCT_10_(mul[10]), .PRODUCT_9_(mul[9]), 
        .PRODUCT_8_(mul[8]), .PRODUCT_7_(N32) );
  NOR2X4 U2 ( .A(n13), .B(n33), .Y(in_17bit_b[1]) );
  NAND2X1 U3 ( .A(n31), .B(n2), .Y(n3) );
  NAND2X1 U4 ( .A(n1), .B(n29), .Y(n4) );
  NAND2X2 U5 ( .A(n3), .B(n4), .Y(in_8bit_b[5]) );
  INVXL U6 ( .A(n31), .Y(n1) );
  INVX1 U7 ( .A(n29), .Y(n2) );
  INVXL U8 ( .A(in_8bit[5]), .Y(n31) );
  XOR2X2 U9 ( .A(in_17bit[2]), .B(n34), .Y(in_17bit_b[2]) );
  NAND2BXL U10 ( .AN(in_17bit[2]), .B(n15), .Y(n35) );
  XOR2X2 U11 ( .A(n27), .B(n23), .Y(in_8bit_b[3]) );
  INVX8 U12 ( .A(n92), .Y(n94) );
  INVX2 U13 ( .A(in_17bit[16]), .Y(n19) );
  OAI22X2 U14 ( .A0(in_17bit[16]), .A1(in_17bit[1]), .B0(in_17bit[0]), .B1(
        in_17bit[1]), .Y(n33) );
  INVX3 U15 ( .A(n89), .Y(n91) );
  NAND2XL U16 ( .A(n24), .B(n21), .Y(n25) );
  NAND2BXL U17 ( .AN(in_8bit[0]), .B(n21), .Y(n22) );
  NOR2X2 U18 ( .A(in_8bit[2]), .B(in_8bit[1]), .Y(n21) );
  NOR3X4 U19 ( .A(in_8bit[6]), .B(n17), .C(n32), .Y(in_8bit_b[7]) );
  NAND2BX4 U20 ( .AN(n30), .B(n31), .Y(n32) );
  AND3X2 U21 ( .A(in_17bit[1]), .B(in_17bit[0]), .C(in_17bit[16]), .Y(n13) );
  NAND2XL U22 ( .A(n22), .B(n16), .Y(n23) );
  NAND2X1 U23 ( .A(n25), .B(n16), .Y(n26) );
  INVX1 U24 ( .A(n85), .Y(n87) );
  XOR2X1 U25 ( .A(mul[13]), .B(n80), .Y(out[6]) );
  NOR2XL U26 ( .A(n7), .B(n81), .Y(n80) );
  NOR2XL U27 ( .A(n7), .B(n5), .Y(n88) );
  NOR2X2 U28 ( .A(n7), .B(n91), .Y(n90) );
  INVX1 U29 ( .A(n79), .Y(n81) );
  INVX1 U30 ( .A(n82), .Y(n84) );
  NAND2BX1 U31 ( .AN(mul[13]), .B(n81), .Y(n82) );
  NOR2X1 U32 ( .A(mul[15]), .B(n6), .Y(n5) );
  NAND2BX1 U33 ( .AN(mul[16]), .B(n5), .Y(n89) );
  CLKINVX3 U34 ( .A(n95), .Y(n97) );
  XOR2X1 U35 ( .A(mul[14]), .B(n83), .Y(out[7]) );
  NOR2X1 U36 ( .A(n7), .B(n84), .Y(n83) );
  INVX4 U37 ( .A(n98), .Y(n100) );
  NAND2BX2 U38 ( .AN(mul[19]), .B(n97), .Y(n98) );
  NAND4BX2 U39 ( .AN(in_8bit[0]), .B(n28), .C(n21), .D(n27), .Y(n30) );
  CLKINVX3 U40 ( .A(n18), .Y(n16) );
  OR2X2 U41 ( .A(n19), .B(n36), .Y(n14) );
  INVX1 U42 ( .A(n35), .Y(n36) );
  NAND2X4 U43 ( .A(n32), .B(n16), .Y(n10) );
  NOR2X4 U44 ( .A(n19), .B(n15), .Y(n34) );
  XNOR2X4 U45 ( .A(n38), .B(n39), .Y(in_17bit_b[4]) );
  NOR2X2 U46 ( .A(n19), .B(n40), .Y(n38) );
  XOR2X4 U47 ( .A(in_8bit[1]), .B(n12), .Y(in_8bit_b[1]) );
  NAND2BX4 U48 ( .AN(mul[20]), .B(n100), .Y(n101) );
  XNOR2X2 U49 ( .A(in_8bit[2]), .B(n20), .Y(in_8bit_b[2]) );
  INVX2 U50 ( .A(n104), .Y(n106) );
  NAND2BX4 U51 ( .AN(mul[18]), .B(n94), .Y(n95) );
  NAND2BX2 U52 ( .AN(mul[21]), .B(n103), .Y(n104) );
  OR2X4 U53 ( .A(n7), .B(n106), .Y(n11) );
  XOR2X4 U54 ( .A(n11), .B(n105), .Y(out[15]) );
  NAND2BX1 U55 ( .AN(mul[10]), .B(n71), .Y(n72) );
  INVXL U56 ( .A(n87), .Y(n6) );
  NAND2XL U57 ( .A(n30), .B(n16), .Y(n29) );
  XNOR2X1 U58 ( .A(in_17bit[16]), .B(n16), .Y(n7) );
  NAND2BX4 U59 ( .AN(mul[17]), .B(n91), .Y(n92) );
  INVX2 U60 ( .A(mul[22]), .Y(n105) );
  NAND2BXL U61 ( .AN(mul[8]), .B(n109), .Y(n65) );
  XOR2X1 U62 ( .A(mul[15]), .B(n86), .Y(out[8]) );
  NOR2XL U63 ( .A(n7), .B(n87), .Y(n86) );
  NOR2XL U64 ( .A(n7), .B(n74), .Y(n73) );
  NOR2XL U65 ( .A(n7), .B(n67), .Y(n66) );
  NAND2XL U66 ( .A(n40), .B(n39), .Y(n42) );
  NAND2BXL U67 ( .AN(n42), .B(n43), .Y(n44) );
  NOR2XL U68 ( .A(n19), .B(n55), .Y(n52) );
  NAND2XL U69 ( .A(n55), .B(n53), .Y(n57) );
  NAND2XL U70 ( .A(n47), .B(n46), .Y(n49) );
  NAND2BXL U71 ( .AN(n49), .B(n50), .Y(n51) );
  NOR2XL U72 ( .A(n19), .B(n63), .Y(n60) );
  NAND2XL U73 ( .A(n63), .B(n61), .Y(n64) );
  NAND2BXL U74 ( .AN(n57), .B(n58), .Y(n59) );
  NOR2X2 U75 ( .A(in_17bit[1]), .B(in_17bit[0]), .Y(n15) );
  NAND2BX1 U76 ( .AN(in_17bit[3]), .B(n36), .Y(n37) );
  MX2X1 U77 ( .A(in_17bit[11]), .B(n8), .S0(in_17bit[16]), .Y(in_17bit_b[11])
         );
  XNOR2X1 U78 ( .A(n64), .B(n110), .Y(n8) );
  MX2X1 U79 ( .A(in_17bit[12]), .B(n9), .S0(in_17bit[16]), .Y(in_17bit_b[12])
         );
  XOR2X1 U80 ( .A(n111), .B(sub_add_52_b0_carry[12]), .Y(n9) );
  MX2X1 U81 ( .A(in_17bit[13]), .B(N18), .S0(in_17bit[16]), .Y(in_17bit_b[13])
         );
  MX2X1 U82 ( .A(in_17bit[14]), .B(N19), .S0(in_17bit[16]), .Y(in_17bit_b[14])
         );
  MX2X1 U83 ( .A(in_17bit[15]), .B(N20), .S0(in_17bit[16]), .Y(in_17bit_b[15])
         );
  XNOR2X4 U84 ( .A(n10), .B(in_8bit[6]), .Y(in_8bit_b[6]) );
  INVX1 U85 ( .A(n68), .Y(n71) );
  NAND2BX1 U86 ( .AN(mul[9]), .B(n67), .Y(n68) );
  INVX1 U87 ( .A(n72), .Y(n74) );
  INVX1 U88 ( .A(n65), .Y(n67) );
  INVX1 U89 ( .A(N32), .Y(n109) );
  XOR2X1 U90 ( .A(mul[23]), .B(n107), .Y(out[16]) );
  NAND2BXL U91 ( .AN(mul[14]), .B(n84), .Y(n85) );
  INVX1 U92 ( .A(n75), .Y(n78) );
  NAND2BX1 U93 ( .AN(mul[11]), .B(n74), .Y(n75) );
  NAND2BX1 U94 ( .AN(mul[12]), .B(n78), .Y(n79) );
  AOI21X1 U95 ( .A0(n106), .A1(n105), .B0(n7), .Y(n107) );
  XOR2X1 U96 ( .A(mul[16]), .B(n88), .Y(out[9]) );
  XOR2X1 U97 ( .A(mul[9]), .B(n66), .Y(out[2]) );
  XOR2X1 U98 ( .A(mul[12]), .B(n76), .Y(out[5]) );
  NOR2X1 U99 ( .A(n7), .B(n78), .Y(n76) );
  XOR2X1 U100 ( .A(mul[10]), .B(n69), .Y(out[3]) );
  NOR2X1 U101 ( .A(n7), .B(n71), .Y(n69) );
  XOR2X1 U102 ( .A(mul[11]), .B(n73), .Y(out[4]) );
  XOR2X4 U103 ( .A(n102), .B(mul[21]), .Y(out[14]) );
  INVX1 U104 ( .A(n118), .Y(out[1]) );
  AOI22XL U105 ( .A0(mul[8]), .A1(n7), .B0(N33), .B1(n119), .Y(n118) );
  INVX1 U106 ( .A(mul[8]), .Y(n108) );
  INVX1 U107 ( .A(n117), .Y(out[0]) );
  AOI22XL U108 ( .A0(N32), .A1(n7), .B0(N32), .B1(n119), .Y(n117) );
  INVXL U109 ( .A(n7), .Y(n119) );
  AND2X2 U110 ( .A(in_8bit[0]), .B(n16), .Y(n12) );
  INVX1 U111 ( .A(n116), .Y(in_8bit_b[0]) );
  AOI22X1 U112 ( .A0(in_8bit[0]), .A1(n16), .B0(in_8bit[0]), .B1(n17), .Y(n116) );
  XNOR2X1 U113 ( .A(n45), .B(n46), .Y(in_17bit_b[6]) );
  NOR2X1 U114 ( .A(n19), .B(n47), .Y(n45) );
  XNOR2X1 U115 ( .A(n52), .B(n53), .Y(in_17bit_b[8]) );
  XOR2X1 U116 ( .A(n43), .B(n41), .Y(in_17bit_b[5]) );
  NAND2X1 U117 ( .A(n42), .B(in_17bit[16]), .Y(n41) );
  XOR2X1 U118 ( .A(n50), .B(n48), .Y(in_17bit_b[7]) );
  NAND2X1 U119 ( .A(n49), .B(in_17bit[16]), .Y(n48) );
  XOR2X1 U120 ( .A(n58), .B(n56), .Y(in_17bit_b[9]) );
  NAND2X1 U121 ( .A(n57), .B(in_17bit[16]), .Y(n56) );
  INVX1 U122 ( .A(n44), .Y(n47) );
  INVX1 U123 ( .A(n51), .Y(n55) );
  INVXL U124 ( .A(in_8bit[7]), .Y(n17) );
  AND2X2 U125 ( .A(N21), .B(in_17bit[16]), .Y(in_17bit_b[16]) );
  NOR2X1 U126 ( .A(n64), .B(in_17bit[11]), .Y(sub_add_52_b0_carry[12]) );
  XNOR2X1 U127 ( .A(n60), .B(n61), .Y(in_17bit_b[10]) );
  INVX1 U128 ( .A(n59), .Y(n63) );
  INVX1 U129 ( .A(in_17bit[4]), .Y(n39) );
  INVX1 U130 ( .A(in_17bit[6]), .Y(n46) );
  XNOR2X2 U131 ( .A(in_17bit[3]), .B(n14), .Y(in_17bit_b[3]) );
  INVX1 U132 ( .A(in_17bit[5]), .Y(n43) );
  INVX1 U133 ( .A(n37), .Y(n40) );
  INVX1 U134 ( .A(in_17bit[8]), .Y(n53) );
  INVX1 U135 ( .A(in_17bit[7]), .Y(n50) );
  INVX1 U136 ( .A(in_17bit[10]), .Y(n61) );
  INVX1 U137 ( .A(in_17bit[9]), .Y(n58) );
  INVX1 U138 ( .A(in_17bit[11]), .Y(n110) );
  INVX1 U139 ( .A(in_17bit[12]), .Y(n111) );
  INVX1 U140 ( .A(in_17bit[13]), .Y(n112) );
  INVX1 U141 ( .A(in_17bit[14]), .Y(n113) );
  INVX1 U142 ( .A(in_17bit[15]), .Y(n114) );
  NOR2X1 U143 ( .A(in_8bit[3]), .B(in_8bit[0]), .Y(n24) );
  INVX1 U144 ( .A(in_8bit[3]), .Y(n27) );
  INVX1 U145 ( .A(in_8bit[4]), .Y(n28) );
  INVX1 U146 ( .A(in_8bit[7]), .Y(n18) );
  INVX4 U147 ( .A(n101), .Y(n103) );
  XOR2X2 U148 ( .A(mul[20]), .B(n99), .Y(out[13]) );
  XOR2X2 U149 ( .A(mul[19]), .B(n96), .Y(out[12]) );
  OAI21XL U150 ( .A0(in_8bit[1]), .A1(in_8bit[0]), .B0(n16), .Y(n20) );
  XOR2X4 U151 ( .A(n28), .B(n26), .Y(in_8bit_b[4]) );
  XOR2X4 U152 ( .A(mul[17]), .B(n90), .Y(out[10]) );
  NOR2X4 U153 ( .A(n7), .B(n94), .Y(n93) );
  XOR2X4 U154 ( .A(mul[18]), .B(n93), .Y(out[11]) );
  NOR2X4 U155 ( .A(n7), .B(n97), .Y(n96) );
  NOR2X4 U156 ( .A(n7), .B(n100), .Y(n99) );
  NOR2X4 U157 ( .A(n7), .B(n103), .Y(n102) );
  XOR2X1 U158 ( .A(n108), .B(n109), .Y(N33) );
  XOR2X1 U159 ( .A(n19), .B(sub_add_52_b0_carry[16]), .Y(N21) );
  AND2X1 U160 ( .A(sub_add_52_b0_carry[15]), .B(n114), .Y(
        sub_add_52_b0_carry[16]) );
  XOR2X1 U161 ( .A(n114), .B(sub_add_52_b0_carry[15]), .Y(N20) );
  AND2X1 U162 ( .A(sub_add_52_b0_carry[14]), .B(n113), .Y(
        sub_add_52_b0_carry[15]) );
  XOR2X1 U163 ( .A(n113), .B(sub_add_52_b0_carry[14]), .Y(N19) );
  AND2X1 U164 ( .A(sub_add_52_b0_carry[13]), .B(n112), .Y(
        sub_add_52_b0_carry[14]) );
  XOR2X1 U165 ( .A(n112), .B(sub_add_52_b0_carry[13]), .Y(N18) );
  AND2X1 U166 ( .A(sub_add_52_b0_carry[12]), .B(n111), .Y(
        sub_add_52_b0_carry[13]) );
endmodule


module multi16_5_DW01_add_0 ( A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, 
        A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, 
        B_20_, B_19_, B_18_, B_17_, B_16_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, 
        SUM_17_, SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, 
        SUM_9_, SUM_8_, SUM_7_, SUM_6_, SUM_5_ );
  input A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_,
         A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, B_20_, B_19_,
         B_18_, B_17_, B_16_;
  output SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, SUM_15_,
         SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, SUM_7_,
         SUM_6_, SUM_5_;
  wire   n1, n3, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39;

  AOI21X4 U2 ( .A0(n19), .A1(n18), .B0(n17), .Y(n38) );
  CLKINVX3 U3 ( .A(n30), .Y(n18) );
  XOR2X1 U4 ( .A(n36), .B(n37), .Y(SUM_19_) );
  OAI21X1 U5 ( .A0(n38), .A1(n31), .B0(n33), .Y(n36) );
  NOR2XL U6 ( .A(B_19_), .B(A_19_), .Y(n28) );
  XOR2X4 U7 ( .A(n19), .B(n39), .Y(SUM_17_) );
  NOR2X1 U8 ( .A(B_18_), .B(A_18_), .Y(n31) );
  AOI21X1 U9 ( .A0(n15), .A1(n32), .B0(n16), .Y(n27) );
  NAND2X2 U10 ( .A(B_18_), .B(A_18_), .Y(n33) );
  INVX2 U11 ( .A(n31), .Y(n15) );
  NOR2BX2 U12 ( .AN(n34), .B(n3), .Y(SUM_16_) );
  BUFX4 U13 ( .A(A_12_), .Y(SUM_12_) );
  CLKINVX3 U14 ( .A(n20), .Y(SUM_15_) );
  NOR2X4 U15 ( .A(n30), .B(n17), .Y(n39) );
  INVX4 U16 ( .A(n35), .Y(n17) );
  CLKINVX4 U17 ( .A(n34), .Y(n19) );
  NAND2X4 U18 ( .A(B_16_), .B(A_16_), .Y(n34) );
  NOR2XL U19 ( .A(B_16_), .B(A_16_), .Y(n3) );
  XOR2X2 U20 ( .A(n1), .B(n38), .Y(SUM_18_) );
  NAND2X2 U21 ( .A(n33), .B(n15), .Y(n1) );
  CLKINVX2 U22 ( .A(A_15_), .Y(n20) );
  INVXL U23 ( .A(n25), .Y(n14) );
  BUFX3 U24 ( .A(A_11_), .Y(SUM_11_) );
  OAI21XL U25 ( .A0(n27), .A1(n28), .B0(n29), .Y(n23) );
  BUFX3 U26 ( .A(A_5_), .Y(SUM_5_) );
  BUFX3 U27 ( .A(A_6_), .Y(SUM_6_) );
  BUFX8 U28 ( .A(A_14_), .Y(SUM_14_) );
  BUFX3 U29 ( .A(A_7_), .Y(SUM_7_) );
  BUFX3 U30 ( .A(A_8_), .Y(SUM_8_) );
  BUFX3 U31 ( .A(A_9_), .Y(SUM_9_) );
  BUFX8 U32 ( .A(A_13_), .Y(SUM_13_) );
  BUFX3 U33 ( .A(A_10_), .Y(SUM_10_) );
  INVXL U34 ( .A(n33), .Y(n16) );
  NAND2X2 U35 ( .A(B_17_), .B(A_17_), .Y(n35) );
  NOR2X4 U36 ( .A(B_17_), .B(A_17_), .Y(n30) );
  XOR2X1 U37 ( .A(n21), .B(n22), .Y(SUM_21_) );
  AOI21X1 U38 ( .A0(n23), .A1(n24), .B0(n14), .Y(n22) );
  XNOR2X1 U39 ( .A(B_21_), .B(A_21_), .Y(n21) );
  XNOR2X1 U40 ( .A(n26), .B(n23), .Y(SUM_20_) );
  OAI21XL U41 ( .A0(n30), .A1(n34), .B0(n35), .Y(n32) );
  NAND2X1 U42 ( .A(n25), .B(n24), .Y(n26) );
  OR2X1 U43 ( .A(B_20_), .B(A_20_), .Y(n24) );
  NAND2X1 U44 ( .A(B_20_), .B(A_20_), .Y(n25) );
  NOR2BX1 U45 ( .AN(n29), .B(n28), .Y(n37) );
  NAND2X1 U46 ( .A(B_19_), .B(A_19_), .Y(n29) );
endmodule


module multi16_5_DW02_mult_0 ( A, B, PRODUCT_23_, PRODUCT_22_, PRODUCT_21_, 
        PRODUCT_20_, PRODUCT_19_, PRODUCT_18_, PRODUCT_17_, PRODUCT_16_, 
        PRODUCT_15_, PRODUCT_14_, PRODUCT_13_, PRODUCT_12_, PRODUCT_11_, 
        PRODUCT_10_, PRODUCT_9_, PRODUCT_8_, PRODUCT_7_ );
  input [16:0] A;
  input [7:0] B;
  output PRODUCT_23_, PRODUCT_22_, PRODUCT_21_, PRODUCT_20_, PRODUCT_19_,
         PRODUCT_18_, PRODUCT_17_, PRODUCT_16_, PRODUCT_15_, PRODUCT_14_,
         PRODUCT_13_, PRODUCT_12_, PRODUCT_11_, PRODUCT_10_, PRODUCT_9_,
         PRODUCT_8_, PRODUCT_7_;
  wire   ab_16__7_, ab_16__6_, ab_16__5_, ab_16__4_, ab_16__3_, ab_16__2_,
         ab_16__1_, ab_16__0_, ab_15__7_, ab_15__6_, ab_15__5_, ab_15__4_,
         ab_15__3_, ab_15__2_, ab_15__1_, ab_15__0_, ab_14__7_, ab_14__6_,
         ab_14__5_, ab_14__4_, ab_14__3_, ab_14__2_, ab_14__1_, ab_14__0_,
         ab_13__7_, ab_13__6_, ab_13__5_, ab_13__4_, ab_13__3_, ab_13__2_,
         ab_13__1_, ab_13__0_, ab_12__7_, ab_12__6_, ab_12__5_, ab_12__4_,
         ab_12__3_, ab_12__2_, ab_12__1_, ab_12__0_, ab_11__7_, ab_11__6_,
         ab_11__5_, ab_11__4_, ab_11__3_, ab_11__2_, ab_11__1_, ab_11__0_,
         ab_10__7_, ab_10__6_, ab_10__5_, ab_10__4_, ab_10__3_, ab_10__2_,
         ab_10__1_, ab_10__0_, ab_9__7_, ab_9__6_, ab_9__5_, ab_9__4_,
         ab_9__3_, ab_9__2_, ab_9__1_, ab_9__0_, ab_8__7_, ab_8__6_, ab_8__5_,
         ab_8__4_, ab_8__3_, ab_8__2_, ab_8__1_, ab_8__0_, ab_7__7_, ab_7__6_,
         ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_, ab_7__0_, ab_6__7_,
         ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_, ab_6__1_, ab_6__0_,
         ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_, ab_5__2_, ab_5__1_,
         ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_, ab_4__3_, ab_4__2_,
         ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_, ab_3__4_, ab_3__3_,
         ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_, ab_2__5_, ab_2__4_,
         ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_, ab_1__6_, ab_1__5_,
         ab_1__4_, ab_1__3_, ab_1__2_, ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_,
         ab_0__3_, ab_0__2_, CARRYB_16__6_, CARRYB_16__5_, CARRYB_16__4_,
         CARRYB_16__3_, CARRYB_16__2_, CARRYB_16__1_, CARRYB_16__0_,
         CARRYB_15__6_, CARRYB_15__5_, CARRYB_15__4_, CARRYB_15__3_,
         CARRYB_15__2_, CARRYB_15__1_, CARRYB_15__0_, CARRYB_14__6_,
         CARRYB_14__5_, CARRYB_14__4_, CARRYB_14__3_, CARRYB_14__2_,
         CARRYB_14__1_, CARRYB_14__0_, CARRYB_13__6_, CARRYB_13__5_,
         CARRYB_13__4_, CARRYB_13__3_, CARRYB_13__2_, CARRYB_13__1_,
         CARRYB_13__0_, CARRYB_12__6_, CARRYB_12__5_, CARRYB_12__4_,
         CARRYB_12__3_, CARRYB_12__2_, CARRYB_12__1_, CARRYB_12__0_,
         CARRYB_11__6_, CARRYB_11__5_, CARRYB_11__4_, CARRYB_11__3_,
         CARRYB_11__2_, CARRYB_11__1_, CARRYB_11__0_, CARRYB_10__6_,
         CARRYB_10__5_, CARRYB_10__4_, CARRYB_10__3_, CARRYB_10__2_,
         CARRYB_10__1_, CARRYB_10__0_, CARRYB_9__6_, CARRYB_9__5_,
         CARRYB_9__4_, CARRYB_9__3_, CARRYB_9__2_, CARRYB_9__1_, CARRYB_9__0_,
         CARRYB_8__6_, CARRYB_8__5_, CARRYB_8__4_, CARRYB_8__3_, CARRYB_8__2_,
         CARRYB_8__1_, CARRYB_8__0_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_,
         CARRYB_7__3_, CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_,
         CARRYB_6__5_, CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_,
         CARRYB_6__0_, CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_,
         CARRYB_5__2_, CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_,
         CARRYB_4__4_, CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_,
         CARRYB_3__6_, CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_,
         CARRYB_3__1_, CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_,
         CARRYB_2__3_, CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__0_,
         SUMB_16__6_, SUMB_16__5_, SUMB_16__4_, SUMB_16__3_, SUMB_16__2_,
         SUMB_16__1_, SUMB_16__0_, SUMB_15__6_, SUMB_15__5_, SUMB_15__4_,
         SUMB_15__3_, SUMB_15__2_, SUMB_15__1_, SUMB_14__6_, SUMB_14__5_,
         SUMB_14__4_, SUMB_14__3_, SUMB_14__2_, SUMB_14__1_, SUMB_13__6_,
         SUMB_13__5_, SUMB_13__4_, SUMB_13__3_, SUMB_13__2_, SUMB_13__1_,
         SUMB_12__6_, SUMB_12__5_, SUMB_12__4_, SUMB_12__3_, SUMB_12__2_,
         SUMB_12__1_, SUMB_11__6_, SUMB_11__5_, SUMB_11__4_, SUMB_11__3_,
         SUMB_11__2_, SUMB_11__1_, SUMB_10__6_, SUMB_10__5_, SUMB_10__4_,
         SUMB_10__3_, SUMB_10__2_, SUMB_10__1_, SUMB_9__6_, SUMB_9__5_,
         SUMB_9__4_, SUMB_9__3_, SUMB_9__2_, SUMB_9__1_, SUMB_8__6_,
         SUMB_8__5_, SUMB_8__4_, SUMB_8__3_, SUMB_8__2_, SUMB_8__1_,
         SUMB_7__6_, SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_,
         SUMB_7__1_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, PROD1_7_, A1_21_, A1_20_, A1_19_, A1_18_,
         A1_17_, A1_16_, A1_15_, A1_13_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_,
         A1_7_, A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_18_, n4, n5, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34;

  ADDFHX4 S2_15_2 ( .A(ab_15__2_), .B(CARRYB_14__2_), .CI(SUMB_14__3_), .CO(
        CARRYB_15__2_), .S(SUMB_15__2_) );
  ADDFHX4 S1_14_0 ( .A(ab_14__0_), .B(CARRYB_13__0_), .CI(SUMB_13__1_), .CO(
        CARRYB_14__0_), .S(A1_12_) );
  ADDFHX4 S2_14_1 ( .A(ab_14__1_), .B(CARRYB_13__1_), .CI(SUMB_13__2_), .CO(
        CARRYB_14__1_), .S(SUMB_14__1_) );
  ADDFHX4 S2_14_2 ( .A(ab_14__2_), .B(CARRYB_13__2_), .CI(SUMB_13__3_), .CO(
        CARRYB_14__2_), .S(SUMB_14__2_) );
  ADDFHX4 S2_14_3 ( .A(ab_14__3_), .B(CARRYB_13__3_), .CI(SUMB_13__4_), .CO(
        CARRYB_14__3_), .S(SUMB_14__3_) );
  ADDFHX4 S1_13_0 ( .A(ab_13__0_), .B(CARRYB_12__0_), .CI(SUMB_12__1_), .CO(
        CARRYB_13__0_), .S(A1_11_) );
  ADDFHX4 S2_13_1 ( .A(ab_13__1_), .B(CARRYB_12__1_), .CI(SUMB_12__2_), .CO(
        CARRYB_13__1_), .S(SUMB_13__1_) );
  ADDFHX4 S2_13_2 ( .A(ab_13__2_), .B(CARRYB_12__2_), .CI(SUMB_12__3_), .CO(
        CARRYB_13__2_), .S(SUMB_13__2_) );
  ADDFHX4 S2_12_1 ( .A(ab_12__1_), .B(CARRYB_11__1_), .CI(SUMB_11__2_), .CO(
        CARRYB_12__1_), .S(SUMB_12__1_) );
  ADDFHX4 S2_12_2 ( .A(ab_12__2_), .B(CARRYB_11__2_), .CI(SUMB_11__3_), .CO(
        CARRYB_12__2_), .S(SUMB_12__2_) );
  ADDFHX4 S2_12_3 ( .A(ab_12__3_), .B(CARRYB_11__3_), .CI(SUMB_11__4_), .CO(
        CARRYB_12__3_), .S(SUMB_12__3_) );
  ADDFHX4 S2_11_3 ( .A(ab_11__3_), .B(CARRYB_10__3_), .CI(SUMB_10__4_), .CO(
        CARRYB_11__3_), .S(SUMB_11__3_) );
  ADDFHX4 S2_11_5 ( .A(ab_11__5_), .B(CARRYB_10__5_), .CI(SUMB_10__6_), .CO(
        CARRYB_11__5_), .S(SUMB_11__5_) );
  ADDFHX4 S2_10_1 ( .A(ab_10__1_), .B(CARRYB_9__1_), .CI(SUMB_9__2_), .CO(
        CARRYB_10__1_), .S(SUMB_10__1_) );
  ADDFHX4 S2_10_2 ( .A(ab_10__2_), .B(CARRYB_9__2_), .CI(SUMB_9__3_), .CO(
        CARRYB_10__2_), .S(SUMB_10__2_) );
  ADDFHX4 S1_9_0 ( .A(ab_9__0_), .B(CARRYB_8__0_), .CI(SUMB_8__1_), .CO(
        CARRYB_9__0_), .S(A1_7_) );
  ADDFHX4 S2_9_3 ( .A(ab_9__3_), .B(CARRYB_8__3_), .CI(SUMB_8__4_), .CO(
        CARRYB_9__3_), .S(SUMB_9__3_) );
  ADDFHX4 S2_9_5 ( .A(ab_9__5_), .B(CARRYB_8__5_), .CI(SUMB_8__6_), .CO(
        CARRYB_9__5_), .S(SUMB_9__5_) );
  ADDFHX4 S2_8_5 ( .A(ab_8__5_), .B(CARRYB_7__5_), .CI(SUMB_7__6_), .CO(
        CARRYB_8__5_), .S(SUMB_8__5_) );
  ADDFHX4 S2_7_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  ADDFHX4 S2_7_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  ADDFHX4 S2_7_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  ADDFHX4 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  ADDFHX4 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  ADDFHX4 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  ADDFHX4 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  ADDFHX4 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  ADDFHX4 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  ADDFHX4 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  ADDFHX4 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  multi16_5_DW01_add_0 FS_1 ( .A_21_(A1_21_), .A_20_(A1_20_), .A_19_(A1_19_), 
        .A_18_(A1_18_), .A_17_(A1_17_), .A_16_(A1_16_), .A_15_(A1_15_), 
        .A_14_(SUMB_16__0_), .A_13_(A1_13_), .A_12_(A1_12_), .A_11_(A1_11_), 
        .A_10_(A1_10_), .A_9_(A1_9_), .A_8_(A1_8_), .A_7_(A1_7_), .A_6_(A1_6_), 
        .A_5_(PROD1_7_), .B_21_(n17), .B_20_(n16), .B_19_(n15), .B_18_(A2_18_), 
        .B_17_(n14), .B_16_(n10), .SUM_21_(PRODUCT_23_), .SUM_20_(PRODUCT_22_), 
        .SUM_19_(PRODUCT_21_), .SUM_18_(PRODUCT_20_), .SUM_17_(PRODUCT_19_), 
        .SUM_16_(PRODUCT_18_), .SUM_15_(PRODUCT_17_), .SUM_14_(PRODUCT_16_), 
        .SUM_13_(PRODUCT_15_), .SUM_12_(PRODUCT_14_), .SUM_11_(PRODUCT_13_), 
        .SUM_10_(PRODUCT_12_), .SUM_9_(PRODUCT_11_), .SUM_8_(PRODUCT_10_), 
        .SUM_7_(PRODUCT_9_), .SUM_6_(PRODUCT_8_), .SUM_5_(PRODUCT_7_) );
  ADDFHX2 S4_3 ( .A(ab_16__3_), .B(CARRYB_15__3_), .CI(SUMB_15__4_), .CO(
        CARRYB_16__3_), .S(SUMB_16__3_) );
  ADDFHX2 S2_15_4 ( .A(ab_15__4_), .B(CARRYB_14__4_), .CI(SUMB_14__5_), .CO(
        CARRYB_15__4_), .S(SUMB_15__4_) );
  ADDFHX2 S2_15_5 ( .A(ab_15__5_), .B(CARRYB_14__5_), .CI(SUMB_14__6_), .CO(
        CARRYB_15__5_), .S(SUMB_15__5_) );
  ADDFHX4 S2_7_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  ADDFHX4 S2_9_4 ( .A(ab_9__4_), .B(CARRYB_8__4_), .CI(SUMB_8__5_), .CO(
        CARRYB_9__4_), .S(SUMB_9__4_) );
  ADDFHX4 S2_11_4 ( .A(ab_11__4_), .B(CARRYB_10__4_), .CI(SUMB_10__5_), .CO(
        CARRYB_11__4_), .S(SUMB_11__4_) );
  ADDFHX2 S3_11_6 ( .A(ab_11__6_), .B(CARRYB_10__6_), .CI(ab_10__7_), .CO(
        CARRYB_11__6_), .S(SUMB_11__6_) );
  ADDFHX4 S3_9_6 ( .A(ab_9__6_), .B(CARRYB_8__6_), .CI(ab_8__7_), .CO(
        CARRYB_9__6_), .S(SUMB_9__6_) );
  ADDFHX4 S3_2_6 ( .A(ab_2__6_), .B(n9), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  ADDFHX4 S1_7_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(PROD1_7_) );
  ADDFHX4 S1_8_0 ( .A(ab_8__0_), .B(CARRYB_7__0_), .CI(SUMB_7__1_), .CO(
        CARRYB_8__0_), .S(A1_6_) );
  ADDFHX4 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  ADDFHX4 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  ADDFHX4 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  ADDFHX4 S1_10_0 ( .A(ab_10__0_), .B(CARRYB_9__0_), .CI(SUMB_9__1_), .CO(
        CARRYB_10__0_), .S(A1_8_) );
  ADDFHX4 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  ADDFHX4 S3_8_6 ( .A(ab_8__6_), .B(CARRYB_7__6_), .CI(ab_7__7_), .CO(
        CARRYB_8__6_), .S(SUMB_8__6_) );
  ADDFHX4 S1_11_0 ( .A(ab_11__0_), .B(CARRYB_10__0_), .CI(SUMB_10__1_), .CO(
        CARRYB_11__0_), .S(A1_9_) );
  ADDFHX4 S1_12_0 ( .A(ab_12__0_), .B(CARRYB_11__0_), .CI(SUMB_11__1_), .CO(
        CARRYB_12__0_), .S(A1_10_) );
  ADDFHX4 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  ADDFHX4 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  ADDFHX2 S3_7_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(
        CARRYB_7__6_), .S(SUMB_7__6_) );
  ADDFHX4 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  ADDFHX4 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  ADDFHX4 S2_14_4 ( .A(ab_14__4_), .B(CARRYB_13__4_), .CI(SUMB_13__5_), .CO(
        CARRYB_14__4_), .S(SUMB_14__4_) );
  ADDFHX4 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  ADDFHX4 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  ADDFHX2 S3_15_6 ( .A(ab_15__6_), .B(CARRYB_14__6_), .CI(ab_14__7_), .CO(
        CARRYB_15__6_), .S(SUMB_15__6_) );
  ADDFHX4 S2_2_3 ( .A(ab_2__3_), .B(n4), .CI(SUMB_1__4_), .CO(CARRYB_2__3_), 
        .S(SUMB_2__3_) );
  ADDFHX4 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  ADDFHX2 S4_0 ( .A(ab_16__0_), .B(CARRYB_15__0_), .CI(SUMB_15__1_), .CO(
        CARRYB_16__0_), .S(SUMB_16__0_) );
  ADDFHX4 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  ADDFHX2 S4_1 ( .A(ab_16__1_), .B(CARRYB_15__1_), .CI(SUMB_15__2_), .CO(
        CARRYB_16__1_), .S(SUMB_16__1_) );
  ADDFHX4 S2_9_1 ( .A(ab_9__1_), .B(CARRYB_8__1_), .CI(SUMB_8__2_), .CO(
        CARRYB_9__1_), .S(SUMB_9__1_) );
  ADDFHX2 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  ADDFX2 S5_6 ( .A(ab_16__6_), .B(CARRYB_15__6_), .CI(ab_15__7_), .CO(
        CARRYB_16__6_), .S(SUMB_16__6_) );
  ADDFHX1 S4_5 ( .A(ab_16__5_), .B(CARRYB_15__5_), .CI(SUMB_15__6_), .CO(
        CARRYB_16__5_), .S(SUMB_16__5_) );
  ADDFHX2 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  ADDFHX2 S3_10_6 ( .A(ab_10__6_), .B(CARRYB_9__6_), .CI(ab_9__7_), .CO(
        CARRYB_10__6_), .S(SUMB_10__6_) );
  ADDFHX2 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  ADDFHX2 S2_2_1 ( .A(ab_2__1_), .B(n5), .CI(SUMB_1__2_), .CO(CARRYB_2__1_), 
        .S(SUMB_2__1_) );
  ADDFHX2 S1_15_0 ( .A(ab_15__0_), .B(CARRYB_14__0_), .CI(SUMB_14__1_), .CO(
        CARRYB_15__0_), .S(A1_13_) );
  ADDFHX2 S2_13_5 ( .A(ab_13__5_), .B(CARRYB_12__5_), .CI(SUMB_12__6_), .CO(
        CARRYB_13__5_), .S(SUMB_13__5_) );
  ADDFHX2 S2_15_1 ( .A(ab_15__1_), .B(CARRYB_14__1_), .CI(SUMB_14__2_), .CO(
        CARRYB_15__1_), .S(SUMB_15__1_) );
  ADDFHX2 S2_10_5 ( .A(ab_10__5_), .B(CARRYB_9__5_), .CI(SUMB_9__6_), .CO(
        CARRYB_10__5_), .S(SUMB_10__5_) );
  ADDFHX2 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  ADDFHX2 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  ADDFHX1 S3_14_6 ( .A(ab_14__6_), .B(CARRYB_13__6_), .CI(ab_13__7_), .CO(
        CARRYB_14__6_), .S(SUMB_14__6_) );
  ADDFHX2 S2_14_5 ( .A(ab_14__5_), .B(CARRYB_13__5_), .CI(SUMB_13__6_), .CO(
        CARRYB_14__5_), .S(SUMB_14__5_) );
  ADDFHX2 S2_2_2 ( .A(ab_2__2_), .B(n8), .CI(SUMB_1__3_), .CO(CARRYB_2__2_), 
        .S(SUMB_2__2_) );
  ADDFHX2 S2_7_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  ADDFHX2 S3_12_6 ( .A(ab_12__6_), .B(CARRYB_11__6_), .CI(ab_11__7_), .CO(
        CARRYB_12__6_), .S(SUMB_12__6_) );
  ADDFHX4 S2_2_4 ( .A(ab_2__4_), .B(n7), .CI(SUMB_1__5_), .CO(CARRYB_2__4_), 
        .S(SUMB_2__4_) );
  ADDFHX4 S2_10_4 ( .A(ab_10__4_), .B(CARRYB_9__4_), .CI(SUMB_9__5_), .CO(
        CARRYB_10__4_), .S(SUMB_10__4_) );
  ADDFHX4 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  ADDFHX4 S2_13_4 ( .A(ab_13__4_), .B(CARRYB_12__4_), .CI(SUMB_12__5_), .CO(
        CARRYB_13__4_), .S(SUMB_13__4_) );
  ADDFHX4 S2_8_4 ( .A(ab_8__4_), .B(CARRYB_7__4_), .CI(SUMB_7__5_), .CO(
        CARRYB_8__4_), .S(SUMB_8__4_) );
  ADDFHX4 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  ADDFHX4 S2_2_5 ( .A(ab_2__5_), .B(n6), .CI(SUMB_1__6_), .CO(CARRYB_2__5_), 
        .S(SUMB_2__5_) );
  ADDFHX4 S2_8_2 ( .A(ab_8__2_), .B(CARRYB_7__2_), .CI(SUMB_7__3_), .CO(
        CARRYB_8__2_), .S(SUMB_8__2_) );
  ADDFHX4 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  ADDFHX4 S2_15_3 ( .A(ab_15__3_), .B(CARRYB_14__3_), .CI(SUMB_14__4_), .CO(
        CARRYB_15__3_), .S(SUMB_15__3_) );
  ADDFHX4 S2_12_5 ( .A(ab_12__5_), .B(CARRYB_11__5_), .CI(SUMB_11__6_), .CO(
        CARRYB_12__5_), .S(SUMB_12__5_) );
  ADDFHX4 S2_11_1 ( .A(ab_11__1_), .B(CARRYB_10__1_), .CI(SUMB_10__2_), .CO(
        CARRYB_11__1_), .S(SUMB_11__1_) );
  ADDFHX4 S2_8_1 ( .A(ab_8__1_), .B(CARRYB_7__1_), .CI(SUMB_7__2_), .CO(
        CARRYB_8__1_), .S(SUMB_8__1_) );
  ADDFHX2 S4_4 ( .A(ab_16__4_), .B(CARRYB_15__4_), .CI(SUMB_15__5_), .CO(
        CARRYB_16__4_), .S(SUMB_16__4_) );
  ADDFHX2 S2_12_4 ( .A(ab_12__4_), .B(CARRYB_11__4_), .CI(SUMB_11__5_), .CO(
        CARRYB_12__4_), .S(SUMB_12__4_) );
  ADDFHX4 S2_13_3 ( .A(ab_13__3_), .B(CARRYB_12__3_), .CI(SUMB_12__4_), .CO(
        CARRYB_13__3_), .S(SUMB_13__3_) );
  ADDFHX4 S4_2 ( .A(ab_16__2_), .B(CARRYB_15__2_), .CI(SUMB_15__3_), .CO(
        CARRYB_16__2_), .S(SUMB_16__2_) );
  ADDFHX4 S2_8_3 ( .A(ab_8__3_), .B(CARRYB_7__3_), .CI(SUMB_7__4_), .CO(
        CARRYB_8__3_), .S(SUMB_8__3_) );
  ADDFHX2 S3_13_6 ( .A(ab_13__6_), .B(CARRYB_12__6_), .CI(ab_12__7_), .CO(
        CARRYB_13__6_), .S(SUMB_13__6_) );
  ADDFHX2 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  ADDFHX2 S2_10_3 ( .A(ab_10__3_), .B(CARRYB_9__3_), .CI(SUMB_9__4_), .CO(
        CARRYB_10__3_), .S(SUMB_10__3_) );
  ADDFHX4 S2_11_2 ( .A(ab_11__2_), .B(CARRYB_10__2_), .CI(SUMB_10__3_), .CO(
        CARRYB_11__2_), .S(SUMB_11__2_) );
  ADDFHX2 S14_19 ( .A(1'b0), .B(CARRYB_16__2_), .CI(SUMB_16__3_), .CO(A2_18_), 
        .S(A1_17_) );
  AND2X4 U2 ( .A(ab_0__3_), .B(ab_1__2_), .Y(n8) );
  AND2X2 U3 ( .A(A[1]), .B(B[5]), .Y(ab_1__5_) );
  AND2X2 U4 ( .A(A[1]), .B(B[6]), .Y(ab_1__6_) );
  INVX3 U5 ( .A(B[6]), .Y(n21) );
  XOR2X1 U6 ( .A(CARRYB_16__3_), .B(SUMB_16__4_), .Y(A1_18_) );
  NOR2X4 U7 ( .A(n21), .B(n18), .Y(ab_0__6_) );
  NAND2X2 U8 ( .A(ab_9__2_), .B(CARRYB_8__2_), .Y(n12) );
  NAND2XL U9 ( .A(A[1]), .B(B[1]), .Y(n20) );
  INVXL U10 ( .A(A[0]), .Y(n18) );
  INVX2 U11 ( .A(B[4]), .Y(n23) );
  XOR2X1 U12 ( .A(CARRYB_16__4_), .B(SUMB_16__5_), .Y(A1_19_) );
  CLKINVX3 U13 ( .A(B[5]), .Y(n22) );
  NOR2X1 U14 ( .A(n22), .B(n18), .Y(ab_0__5_) );
  AND2X2 U16 ( .A(ab_0__4_), .B(ab_1__3_), .Y(n4) );
  AND2X2 U17 ( .A(ab_0__2_), .B(n28), .Y(n5) );
  AND2X2 U18 ( .A(ab_0__6_), .B(ab_1__5_), .Y(n6) );
  AND2X2 U19 ( .A(ab_0__5_), .B(ab_1__4_), .Y(n7) );
  AND2X2 U20 ( .A(ab_0__7_), .B(ab_1__6_), .Y(n9) );
  AND2X2 U21 ( .A(CARRYB_16__0_), .B(SUMB_16__1_), .Y(n10) );
  AND2X2 U22 ( .A(A[2]), .B(B[4]), .Y(ab_2__4_) );
  XOR3X2 U23 ( .A(CARRYB_8__2_), .B(ab_9__2_), .C(SUMB_8__3_), .Y(SUMB_9__2_)
         );
  NOR2X1 U24 ( .A(n27), .B(n18), .Y(ab_0__7_) );
  INVX1 U25 ( .A(B[7]), .Y(n27) );
  AND2X2 U26 ( .A(A[2]), .B(B[2]), .Y(ab_2__2_) );
  NAND3X4 U27 ( .A(n13), .B(n11), .C(n12), .Y(CARRYB_9__2_) );
  AND2X2 U28 ( .A(A[2]), .B(B[3]), .Y(ab_2__3_) );
  NAND2X2 U29 ( .A(SUMB_8__3_), .B(CARRYB_8__2_), .Y(n11) );
  NAND2X2 U30 ( .A(ab_9__2_), .B(SUMB_8__3_), .Y(n13) );
  AND2X2 U31 ( .A(A[1]), .B(B[2]), .Y(ab_1__2_) );
  NOR2X1 U32 ( .A(n25), .B(n18), .Y(ab_0__2_) );
  AND2X2 U33 ( .A(CARRYB_16__3_), .B(SUMB_16__4_), .Y(n15) );
  AND2X1 U34 ( .A(A[8]), .B(B[0]), .Y(ab_8__0_) );
  AND2X1 U35 ( .A(A[5]), .B(B[1]), .Y(ab_5__1_) );
  INVXL U36 ( .A(B[2]), .Y(n25) );
  AND2X1 U37 ( .A(A[7]), .B(B[0]), .Y(ab_7__0_) );
  AND2X1 U38 ( .A(A[6]), .B(B[0]), .Y(ab_6__0_) );
  AND2X1 U39 ( .A(A[5]), .B(B[0]), .Y(ab_5__0_) );
  AND2X1 U40 ( .A(A[4]), .B(B[0]), .Y(ab_4__0_) );
  AND2X1 U41 ( .A(A[4]), .B(B[1]), .Y(ab_4__1_) );
  AND2X1 U42 ( .A(A[9]), .B(B[0]), .Y(ab_9__0_) );
  AND2X1 U43 ( .A(A[11]), .B(B[1]), .Y(ab_11__1_) );
  AND2X1 U44 ( .A(A[10]), .B(B[1]), .Y(ab_10__1_) );
  AND2X1 U45 ( .A(A[9]), .B(B[1]), .Y(ab_9__1_) );
  AND2X1 U46 ( .A(A[11]), .B(B[0]), .Y(ab_11__0_) );
  AND2X1 U47 ( .A(A[8]), .B(B[1]), .Y(ab_8__1_) );
  AND2X1 U48 ( .A(A[10]), .B(B[0]), .Y(ab_10__0_) );
  AND2X1 U49 ( .A(A[7]), .B(B[1]), .Y(ab_7__1_) );
  AND2X1 U50 ( .A(A[6]), .B(B[1]), .Y(ab_6__1_) );
  INVXL U51 ( .A(B[0]), .Y(n34) );
  INVXL U52 ( .A(B[1]), .Y(n26) );
  AND2X1 U53 ( .A(A[10]), .B(B[7]), .Y(ab_10__7_) );
  AND2X1 U54 ( .A(A[8]), .B(B[7]), .Y(ab_8__7_) );
  AND2X1 U55 ( .A(A[6]), .B(B[7]), .Y(ab_6__7_) );
  AND2X1 U56 ( .A(A[5]), .B(B[7]), .Y(ab_5__7_) );
  AND2X1 U57 ( .A(A[3]), .B(B[0]), .Y(ab_3__0_) );
  AND2X1 U58 ( .A(A[2]), .B(B[1]), .Y(ab_2__1_) );
  XOR2X1 U59 ( .A(ab_1__6_), .B(ab_0__7_), .Y(SUMB_1__6_) );
  AND2X1 U60 ( .A(A[3]), .B(B[5]), .Y(ab_3__5_) );
  XOR2X1 U61 ( .A(ab_1__5_), .B(ab_0__6_), .Y(SUMB_1__5_) );
  INVX4 U62 ( .A(B[3]), .Y(n24) );
  XOR2X1 U63 ( .A(ab_1__4_), .B(ab_0__5_), .Y(SUMB_1__4_) );
  AND2X2 U64 ( .A(CARRYB_16__1_), .B(SUMB_16__2_), .Y(n14) );
  XOR2X2 U65 ( .A(CARRYB_16__0_), .B(SUMB_16__1_), .Y(A1_15_) );
  NOR2X1 U66 ( .A(n29), .B(n26), .Y(ab_16__1_) );
  NOR2X1 U67 ( .A(n29), .B(n22), .Y(ab_16__5_) );
  INVX1 U68 ( .A(n20), .Y(n28) );
  NOR2X1 U69 ( .A(n29), .B(n25), .Y(ab_16__2_) );
  XOR2X1 U70 ( .A(CARRYB_16__6_), .B(ab_16__7_), .Y(A1_21_) );
  XOR2X1 U71 ( .A(n28), .B(ab_0__2_), .Y(SUMB_1__1_) );
  XOR2X1 U72 ( .A(CARRYB_16__5_), .B(SUMB_16__6_), .Y(A1_20_) );
  AND2X1 U73 ( .A(CARRYB_16__4_), .B(SUMB_16__5_), .Y(n16) );
  AND2X2 U74 ( .A(CARRYB_16__5_), .B(SUMB_16__6_), .Y(n17) );
  NOR2XL U75 ( .A(n23), .B(n18), .Y(ab_0__4_) );
  NOR2XL U76 ( .A(n24), .B(n18), .Y(ab_0__3_) );
  NOR2XL U77 ( .A(n29), .B(n23), .Y(ab_16__4_) );
  NOR2XL U78 ( .A(n30), .B(n25), .Y(ab_15__2_) );
  NOR2XL U79 ( .A(n31), .B(n25), .Y(ab_14__2_) );
  NOR2X1 U80 ( .A(n30), .B(n26), .Y(ab_15__1_) );
  NOR2XL U81 ( .A(n32), .B(n25), .Y(ab_13__2_) );
  NOR2X1 U82 ( .A(n31), .B(n26), .Y(ab_14__1_) );
  NOR2XL U83 ( .A(n33), .B(n25), .Y(ab_12__2_) );
  NOR2XL U84 ( .A(n31), .B(n23), .Y(ab_14__4_) );
  NOR2X1 U85 ( .A(n32), .B(n26), .Y(ab_13__1_) );
  NOR2XL U86 ( .A(n32), .B(n23), .Y(ab_13__4_) );
  NOR2XL U87 ( .A(n33), .B(n23), .Y(ab_12__4_) );
  AND2X1 U88 ( .A(A[11]), .B(B[2]), .Y(ab_11__2_) );
  NOR2X1 U89 ( .A(n33), .B(n26), .Y(ab_12__1_) );
  AND2X1 U90 ( .A(A[10]), .B(B[2]), .Y(ab_10__2_) );
  NOR2X1 U91 ( .A(n33), .B(n22), .Y(ab_12__5_) );
  NOR2X1 U92 ( .A(n32), .B(n22), .Y(ab_13__5_) );
  AND2X1 U93 ( .A(A[11]), .B(B[5]), .Y(ab_11__5_) );
  AND2X1 U94 ( .A(A[9]), .B(B[2]), .Y(ab_9__2_) );
  AND2X1 U95 ( .A(A[10]), .B(B[5]), .Y(ab_10__5_) );
  AND2X1 U96 ( .A(A[8]), .B(B[2]), .Y(ab_8__2_) );
  AND2X1 U97 ( .A(A[9]), .B(B[5]), .Y(ab_9__5_) );
  AND2X1 U98 ( .A(A[11]), .B(B[6]), .Y(ab_11__6_) );
  AND2X1 U99 ( .A(A[8]), .B(B[5]), .Y(ab_8__5_) );
  AND2X1 U100 ( .A(A[7]), .B(B[2]), .Y(ab_7__2_) );
  AND2X1 U101 ( .A(A[7]), .B(B[5]), .Y(ab_7__5_) );
  AND2X1 U102 ( .A(A[6]), .B(B[5]), .Y(ab_6__5_) );
  AND2X1 U103 ( .A(A[6]), .B(B[2]), .Y(ab_6__2_) );
  AND2X2 U104 ( .A(A[9]), .B(B[7]), .Y(ab_9__7_) );
  AND2X1 U105 ( .A(A[10]), .B(B[6]), .Y(ab_10__6_) );
  AND2X1 U106 ( .A(A[5]), .B(B[5]), .Y(ab_5__5_) );
  AND2X1 U107 ( .A(A[5]), .B(B[2]), .Y(ab_5__2_) );
  AND2X1 U108 ( .A(A[4]), .B(B[5]), .Y(ab_4__5_) );
  AND2X1 U109 ( .A(A[9]), .B(B[6]), .Y(ab_9__6_) );
  AND2X1 U110 ( .A(A[4]), .B(B[2]), .Y(ab_4__2_) );
  AND2X2 U111 ( .A(A[7]), .B(B[7]), .Y(ab_7__7_) );
  AND2X1 U112 ( .A(A[8]), .B(B[6]), .Y(ab_8__6_) );
  AND2X2 U113 ( .A(A[3]), .B(B[2]), .Y(ab_3__2_) );
  AND2X1 U114 ( .A(A[7]), .B(B[6]), .Y(ab_7__6_) );
  AND2X2 U115 ( .A(A[3]), .B(B[1]), .Y(ab_3__1_) );
  AND2X2 U116 ( .A(A[2]), .B(B[7]), .Y(ab_2__7_) );
  AND2X1 U117 ( .A(A[3]), .B(B[6]), .Y(ab_3__6_) );
  AND2X1 U118 ( .A(A[3]), .B(B[7]), .Y(ab_3__7_) );
  AND2X1 U119 ( .A(A[4]), .B(B[6]), .Y(ab_4__6_) );
  AND2X1 U120 ( .A(A[4]), .B(B[7]), .Y(ab_4__7_) );
  AND2X1 U121 ( .A(A[5]), .B(B[6]), .Y(ab_5__6_) );
  AND2X1 U122 ( .A(A[6]), .B(B[6]), .Y(ab_6__6_) );
  NOR2XL U123 ( .A(n20), .B(n19), .Y(CARRYB_1__0_) );
  AND2X2 U124 ( .A(A[11]), .B(B[7]), .Y(ab_11__7_) );
  XOR2X1 U125 ( .A(ab_1__3_), .B(ab_0__4_), .Y(SUMB_1__3_) );
  XOR2X1 U126 ( .A(ab_1__2_), .B(ab_0__3_), .Y(SUMB_1__2_) );
  AND2X1 U127 ( .A(A[2]), .B(B[6]), .Y(ab_2__6_) );
  AND2X1 U128 ( .A(A[2]), .B(B[5]), .Y(ab_2__5_) );
  NOR2XL U129 ( .A(n30), .B(n22), .Y(ab_15__5_) );
  NOR2XL U130 ( .A(n31), .B(n22), .Y(ab_14__5_) );
  NOR2XL U131 ( .A(n30), .B(n23), .Y(ab_15__4_) );
  AND2X2 U132 ( .A(A[2]), .B(B[0]), .Y(ab_2__0_) );
  INVX1 U133 ( .A(A[16]), .Y(n29) );
  AND2X1 U134 ( .A(A[11]), .B(B[3]), .Y(ab_11__3_) );
  AND2X1 U135 ( .A(A[10]), .B(B[3]), .Y(ab_10__3_) );
  AND2X1 U136 ( .A(A[11]), .B(B[4]), .Y(ab_11__4_) );
  AND2X1 U137 ( .A(A[10]), .B(B[4]), .Y(ab_10__4_) );
  AND2X1 U138 ( .A(A[9]), .B(B[3]), .Y(ab_9__3_) );
  AND2X1 U139 ( .A(A[9]), .B(B[4]), .Y(ab_9__4_) );
  AND2X1 U140 ( .A(A[8]), .B(B[3]), .Y(ab_8__3_) );
  AND2X1 U141 ( .A(A[8]), .B(B[4]), .Y(ab_8__4_) );
  AND2X1 U142 ( .A(A[7]), .B(B[3]), .Y(ab_7__3_) );
  AND2X1 U143 ( .A(A[7]), .B(B[4]), .Y(ab_7__4_) );
  AND2X1 U144 ( .A(A[6]), .B(B[4]), .Y(ab_6__4_) );
  AND2X1 U145 ( .A(A[6]), .B(B[3]), .Y(ab_6__3_) );
  AND2X1 U146 ( .A(A[5]), .B(B[4]), .Y(ab_5__4_) );
  AND2X1 U147 ( .A(A[5]), .B(B[3]), .Y(ab_5__3_) );
  AND2X1 U148 ( .A(A[4]), .B(B[4]), .Y(ab_4__4_) );
  AND2X1 U149 ( .A(A[4]), .B(B[3]), .Y(ab_4__3_) );
  AND2X1 U150 ( .A(A[3]), .B(B[3]), .Y(ab_3__3_) );
  NAND2XL U151 ( .A(A[0]), .B(B[0]), .Y(n19) );
  AND2X1 U152 ( .A(A[3]), .B(B[4]), .Y(ab_3__4_) );
  INVX1 U153 ( .A(A[12]), .Y(n33) );
  INVX1 U154 ( .A(A[13]), .Y(n32) );
  INVX1 U155 ( .A(A[14]), .Y(n31) );
  INVX1 U156 ( .A(A[15]), .Y(n30) );
  XOR2X4 U157 ( .A(CARRYB_16__1_), .B(SUMB_16__2_), .Y(A1_16_) );
  NOR2XL U158 ( .A(n29), .B(n24), .Y(ab_16__3_) );
  NOR2XL U159 ( .A(n30), .B(n24), .Y(ab_15__3_) );
  NOR2XL U160 ( .A(n31), .B(n24), .Y(ab_14__3_) );
  NOR2XL U161 ( .A(n32), .B(n24), .Y(ab_13__3_) );
  NOR2XL U162 ( .A(n33), .B(n24), .Y(ab_12__3_) );
  NOR2XL U163 ( .A(n29), .B(n27), .Y(ab_16__7_) );
  NOR2XL U164 ( .A(n30), .B(n27), .Y(ab_15__7_) );
  NOR2XL U165 ( .A(n31), .B(n27), .Y(ab_14__7_) );
  NOR2XL U166 ( .A(n32), .B(n27), .Y(ab_13__7_) );
  NOR2XL U167 ( .A(n33), .B(n27), .Y(ab_12__7_) );
  NOR2XL U168 ( .A(n29), .B(n21), .Y(ab_16__6_) );
  NOR2XL U169 ( .A(n30), .B(n21), .Y(ab_15__6_) );
  NOR2XL U170 ( .A(n31), .B(n21), .Y(ab_14__6_) );
  NOR2XL U171 ( .A(n32), .B(n21), .Y(ab_13__6_) );
  NOR2XL U172 ( .A(n33), .B(n21), .Y(ab_12__6_) );
  AND2X1 U173 ( .A(A[1]), .B(B[7]), .Y(ab_1__7_) );
  AND2X2 U174 ( .A(A[1]), .B(B[4]), .Y(ab_1__4_) );
  AND2X2 U175 ( .A(A[1]), .B(B[3]), .Y(ab_1__3_) );
  NOR2X1 U177 ( .A(n34), .B(n29), .Y(ab_16__0_) );
  NOR2X1 U178 ( .A(n34), .B(n30), .Y(ab_15__0_) );
  NOR2X1 U179 ( .A(n34), .B(n31), .Y(ab_14__0_) );
  NOR2X1 U180 ( .A(n34), .B(n32), .Y(ab_13__0_) );
  NOR2X1 U181 ( .A(n34), .B(n33), .Y(ab_12__0_) );
endmodule


module multi16_5 ( in_17bit, in_8bit, out );
  input [16:0] in_17bit;
  input [7:0] in_8bit;
  output [16:0] out;
  wire   N19, N20, N21, N32, N33, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n55, n56, n57, n58, n59, n60, n61, n63, n64, n65, n66, n67, n68, n69,
         n71, n72, n73, n74, n75, n76, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n124, n125, n126, n127;
  wire   [16:1] in_17bit_b;
  wire   [7:0] in_8bit_b;
  wire   [23:8] mul;
  wire   [16:13] sub_add_52_b0_carry;

  multi16_5_DW02_mult_0 mult_55 ( .A({in_17bit_b, in_17bit[0]}), .B(in_8bit_b), 
        .PRODUCT_23_(mul[23]), .PRODUCT_22_(mul[22]), .PRODUCT_21_(mul[21]), 
        .PRODUCT_20_(mul[20]), .PRODUCT_19_(mul[19]), .PRODUCT_18_(mul[18]), 
        .PRODUCT_17_(mul[17]), .PRODUCT_16_(mul[16]), .PRODUCT_15_(mul[15]), 
        .PRODUCT_14_(mul[14]), .PRODUCT_13_(mul[13]), .PRODUCT_12_(mul[12]), 
        .PRODUCT_11_(mul[11]), .PRODUCT_10_(mul[10]), .PRODUCT_9_(mul[9]), 
        .PRODUCT_8_(mul[8]), .PRODUCT_7_(N32) );
  NAND3X1 U2 ( .A(n19), .B(in_17bit[0]), .C(in_17bit[1]), .Y(n41) );
  CLKINVX3 U3 ( .A(in_17bit[16]), .Y(n22) );
  XOR2X2 U4 ( .A(mul[17]), .B(n101), .Y(out[10]) );
  NAND2X1 U5 ( .A(mul[18]), .B(n2), .Y(n3) );
  NAND2X1 U6 ( .A(n1), .B(n103), .Y(n4) );
  NAND2X2 U7 ( .A(n3), .B(n4), .Y(out[11]) );
  INVXL U8 ( .A(mul[18]), .Y(n1) );
  INVX2 U9 ( .A(n103), .Y(n2) );
  OAI22X1 U10 ( .A0(in_17bit[0]), .A1(in_17bit[1]), .B0(in_17bit[1]), .B1(n19), 
        .Y(n40) );
  NOR2X4 U11 ( .A(in_17bit[1]), .B(in_17bit[0]), .Y(n16) );
  CLKINVX3 U12 ( .A(n37), .Y(n5) );
  NOR2X2 U13 ( .A(n18), .B(n39), .Y(n37) );
  NOR2X2 U14 ( .A(n10), .B(n104), .Y(n103) );
  XOR2X2 U15 ( .A(n35), .B(n33), .Y(in_8bit_b[5]) );
  INVX2 U16 ( .A(n106), .Y(n108) );
  INVX4 U17 ( .A(n112), .Y(n115) );
  INVX2 U18 ( .A(n36), .Y(n39) );
  NOR2X4 U19 ( .A(n10), .B(n111), .Y(n110) );
  NOR3X4 U20 ( .A(in_8bit[1]), .B(in_8bit[3]), .C(in_8bit[2]), .Y(n31) );
  INVX3 U21 ( .A(n18), .Y(n17) );
  NAND2X2 U22 ( .A(n32), .B(n31), .Y(n34) );
  INVX4 U23 ( .A(n5), .Y(n6) );
  NOR2BX2 U24 ( .AN(n41), .B(n40), .Y(in_17bit_b[1]) );
  XOR2X2 U25 ( .A(n27), .B(n26), .Y(in_8bit_b[3]) );
  NAND2XL U26 ( .A(n34), .B(n17), .Y(n33) );
  XOR2X2 U27 ( .A(n30), .B(in_8bit[4]), .Y(in_8bit_b[4]) );
  NOR2X2 U28 ( .A(n21), .B(n44), .Y(n43) );
  NOR2X1 U29 ( .A(n10), .B(n7), .Y(n101) );
  NOR2X2 U30 ( .A(in_8bit[4]), .B(in_8bit[0]), .Y(n32) );
  INVX1 U31 ( .A(n42), .Y(n44) );
  XNOR2X2 U32 ( .A(in_8bit[2]), .B(n23), .Y(in_8bit_b[2]) );
  OAI21X2 U33 ( .A0(in_8bit[1]), .A1(in_8bit[0]), .B0(n17), .Y(n23) );
  INVX1 U34 ( .A(n91), .Y(n93) );
  NAND2BX1 U35 ( .AN(mul[12]), .B(n90), .Y(n91) );
  XOR2X1 U36 ( .A(n51), .B(n49), .Y(in_17bit_b[5]) );
  INVX1 U37 ( .A(n9), .Y(n8) );
  NAND2BX2 U38 ( .AN(mul[18]), .B(n104), .Y(n106) );
  XOR2X2 U39 ( .A(mul[21]), .B(n110), .Y(out[14]) );
  INVX1 U40 ( .A(in_8bit[7]), .Y(n18) );
  NAND2BX2 U41 ( .AN(n34), .B(n35), .Y(n36) );
  INVX1 U42 ( .A(n97), .Y(n99) );
  NAND2BX1 U43 ( .AN(mul[14]), .B(n96), .Y(n97) );
  INVXL U44 ( .A(in_17bit[16]), .Y(n20) );
  AND3X2 U45 ( .A(n39), .B(n17), .C(n38), .Y(in_8bit_b[7]) );
  AOI21X1 U46 ( .A0(n115), .A1(n114), .B0(n10), .Y(n116) );
  NAND2BXL U47 ( .AN(in_17bit[2]), .B(n16), .Y(n42) );
  OAI21X2 U48 ( .A0(mul[19]), .A1(n106), .B0(n127), .Y(n107) );
  CLKINVX4 U49 ( .A(mul[19]), .Y(n105) );
  INVX4 U50 ( .A(n22), .Y(n19) );
  XNOR2X2 U51 ( .A(mul[20]), .B(n107), .Y(out[13]) );
  XNOR2X4 U52 ( .A(in_17bit[2]), .B(n15), .Y(in_17bit_b[2]) );
  OR2X4 U53 ( .A(n21), .B(n16), .Y(n15) );
  INVX4 U54 ( .A(n109), .Y(n111) );
  XOR2X2 U55 ( .A(in_8bit[1]), .B(n14), .Y(in_8bit_b[1]) );
  INVX4 U56 ( .A(n102), .Y(n104) );
  NAND2BX4 U57 ( .AN(mul[17]), .B(n7), .Y(n102) );
  NAND2BX2 U58 ( .AN(mul[21]), .B(n111), .Y(n112) );
  XNOR2X1 U59 ( .A(n46), .B(n47), .Y(in_17bit_b[4]) );
  NAND2XL U60 ( .A(n50), .B(n19), .Y(n49) );
  XNOR2X1 U61 ( .A(n19), .B(n17), .Y(n10) );
  NOR2X4 U62 ( .A(mul[16]), .B(n8), .Y(n7) );
  NAND2BXL U63 ( .AN(mul[10]), .B(n84), .Y(n85) );
  NAND2BXL U64 ( .AN(mul[8]), .B(n118), .Y(n79) );
  NOR2X4 U65 ( .A(mul[15]), .B(n97), .Y(n9) );
  INVX2 U66 ( .A(mul[22]), .Y(n114) );
  XOR2X1 U67 ( .A(mul[23]), .B(n116), .Y(out[16]) );
  NOR2XL U68 ( .A(n10), .B(n93), .Y(n92) );
  XOR2X1 U69 ( .A(mul[15]), .B(n98), .Y(out[8]) );
  XOR2X1 U70 ( .A(mul[14]), .B(n95), .Y(out[7]) );
  NOR2XL U71 ( .A(n10), .B(n96), .Y(n95) );
  NOR2XL U72 ( .A(n10), .B(n81), .Y(n80) );
  NOR2XL U73 ( .A(n20), .B(n64), .Y(n61) );
  NAND2XL U74 ( .A(n58), .B(n19), .Y(n57) );
  NAND2XL U75 ( .A(n56), .B(n55), .Y(n58) );
  NAND2BXL U76 ( .AN(n50), .B(n51), .Y(n52) );
  NAND2BXL U77 ( .AN(n58), .B(n59), .Y(n60) );
  NOR2XL U78 ( .A(n20), .B(n72), .Y(n69) );
  NAND2XL U79 ( .A(n66), .B(n19), .Y(n65) );
  NAND2XL U80 ( .A(n72), .B(n71), .Y(n76) );
  NAND2XL U81 ( .A(n76), .B(n19), .Y(n73) );
  NAND2XL U82 ( .A(n64), .B(n63), .Y(n66) );
  NAND2BXL U83 ( .AN(n66), .B(n67), .Y(n68) );
  AND2X1 U84 ( .A(N21), .B(n19), .Y(in_17bit_b[16]) );
  INVX1 U85 ( .A(n45), .Y(n48) );
  INVXL U86 ( .A(in_17bit[4]), .Y(n47) );
  INVXL U87 ( .A(in_17bit[6]), .Y(n55) );
  INVXL U88 ( .A(in_17bit[5]), .Y(n51) );
  MX2X1 U89 ( .A(in_17bit[13]), .B(n11), .S0(n19), .Y(in_17bit_b[13]) );
  XNOR2X1 U90 ( .A(n78), .B(n120), .Y(n11) );
  MX2X1 U91 ( .A(in_17bit[14]), .B(N19), .S0(n19), .Y(in_17bit_b[14]) );
  MX2X1 U92 ( .A(in_17bit[15]), .B(N20), .S0(n19), .Y(in_17bit_b[15]) );
  INVXL U93 ( .A(in_17bit[8]), .Y(n63) );
  INVXL U94 ( .A(in_17bit[7]), .Y(n59) );
  MX2X1 U95 ( .A(in_17bit[12]), .B(n12), .S0(n19), .Y(in_17bit_b[12]) );
  XNOR2X1 U96 ( .A(in_17bit[12]), .B(n74), .Y(n12) );
  INVX1 U97 ( .A(n85), .Y(n87) );
  INVX1 U98 ( .A(n88), .Y(n90) );
  NAND2BX1 U99 ( .AN(mul[11]), .B(n87), .Y(n88) );
  INVX1 U100 ( .A(n79), .Y(n81) );
  INVX1 U101 ( .A(n82), .Y(n84) );
  NAND2BX1 U102 ( .AN(mul[9]), .B(n81), .Y(n82) );
  INVX1 U103 ( .A(N32), .Y(n118) );
  INVX1 U104 ( .A(n94), .Y(n96) );
  NAND2BX1 U105 ( .AN(mul[13]), .B(n93), .Y(n94) );
  NOR2XL U106 ( .A(n10), .B(n99), .Y(n98) );
  XOR2X1 U107 ( .A(mul[9]), .B(n80), .Y(out[2]) );
  XOR2X1 U108 ( .A(mul[11]), .B(n86), .Y(out[4]) );
  NOR2X1 U109 ( .A(n10), .B(n87), .Y(n86) );
  XOR2X1 U110 ( .A(mul[12]), .B(n89), .Y(out[5]) );
  NOR2X1 U111 ( .A(n10), .B(n90), .Y(n89) );
  XOR2X1 U112 ( .A(mul[13]), .B(n92), .Y(out[6]) );
  XOR2X1 U113 ( .A(mul[10]), .B(n83), .Y(out[3]) );
  NOR2X1 U114 ( .A(n10), .B(n84), .Y(n83) );
  XOR2X4 U115 ( .A(n13), .B(n105), .Y(out[12]) );
  OR2X4 U116 ( .A(n10), .B(n108), .Y(n13) );
  INVX1 U117 ( .A(n126), .Y(out[1]) );
  AOI22X1 U118 ( .A0(mul[8]), .A1(n10), .B0(N33), .B1(n127), .Y(n126) );
  INVX1 U119 ( .A(mul[8]), .Y(n117) );
  INVX1 U120 ( .A(n125), .Y(out[0]) );
  AOI22XL U121 ( .A0(N32), .A1(n10), .B0(N32), .B1(n127), .Y(n125) );
  INVXL U122 ( .A(n10), .Y(n127) );
  AND2X1 U123 ( .A(in_8bit[0]), .B(n17), .Y(n14) );
  INVX1 U124 ( .A(n124), .Y(in_8bit_b[0]) );
  AOI22XL U125 ( .A0(in_8bit[0]), .A1(n17), .B0(in_8bit[0]), .B1(n18), .Y(n124) );
  NOR2X1 U126 ( .A(n20), .B(n48), .Y(n46) );
  XNOR2X1 U127 ( .A(n53), .B(n55), .Y(in_17bit_b[6]) );
  NOR2X1 U128 ( .A(n20), .B(n56), .Y(n53) );
  XNOR2X1 U129 ( .A(n61), .B(n63), .Y(in_17bit_b[8]) );
  XNOR2X1 U130 ( .A(n69), .B(n71), .Y(in_17bit_b[10]) );
  XOR2X1 U131 ( .A(n59), .B(n57), .Y(in_17bit_b[7]) );
  XOR2X1 U132 ( .A(n67), .B(n65), .Y(in_17bit_b[9]) );
  INVX1 U133 ( .A(in_8bit[5]), .Y(n35) );
  NAND2X1 U134 ( .A(n48), .B(n47), .Y(n50) );
  INVX1 U135 ( .A(n52), .Y(n56) );
  INVX1 U136 ( .A(n60), .Y(n64) );
  INVX1 U137 ( .A(n68), .Y(n72) );
  NAND3BX1 U138 ( .AN(n76), .B(n119), .C(n75), .Y(n78) );
  XOR2X1 U139 ( .A(n75), .B(n73), .Y(in_17bit_b[11]) );
  INVX1 U140 ( .A(n78), .Y(sub_add_52_b0_carry[13]) );
  NAND2BXL U141 ( .AN(in_17bit[3]), .B(n44), .Y(n45) );
  INVX1 U142 ( .A(in_17bit[16]), .Y(n21) );
  NOR2X1 U143 ( .A(in_17bit[11]), .B(n76), .Y(n74) );
  INVX1 U144 ( .A(in_17bit[9]), .Y(n67) );
  INVX1 U145 ( .A(in_17bit[10]), .Y(n71) );
  INVX1 U146 ( .A(in_17bit[11]), .Y(n75) );
  INVX1 U147 ( .A(in_17bit[12]), .Y(n119) );
  INVX1 U148 ( .A(in_17bit[13]), .Y(n120) );
  INVX1 U149 ( .A(in_17bit[14]), .Y(n121) );
  INVX1 U150 ( .A(in_17bit[15]), .Y(n122) );
  INVX1 U151 ( .A(in_8bit[3]), .Y(n27) );
  NAND2X1 U152 ( .A(n25), .B(n17), .Y(n26) );
  NAND2BXL U153 ( .AN(in_8bit[0]), .B(n24), .Y(n25) );
  AOI21X1 U154 ( .A0(n29), .A1(n28), .B0(n18), .Y(n30) );
  NOR2XL U155 ( .A(in_8bit[3]), .B(in_8bit[0]), .Y(n29) );
  INVX1 U156 ( .A(in_8bit[6]), .Y(n38) );
  NAND3BX2 U157 ( .AN(mul[20]), .B(n108), .C(n105), .Y(n109) );
  NOR2XL U158 ( .A(in_8bit[2]), .B(in_8bit[1]), .Y(n28) );
  NOR2XL U159 ( .A(in_8bit[2]), .B(in_8bit[1]), .Y(n24) );
  XNOR2X4 U160 ( .A(n6), .B(n38), .Y(in_8bit_b[6]) );
  XOR2X4 U161 ( .A(in_17bit[3]), .B(n43), .Y(in_17bit_b[3]) );
  NOR2X4 U162 ( .A(n10), .B(n9), .Y(n100) );
  XOR2X4 U163 ( .A(mul[16]), .B(n100), .Y(out[9]) );
  NOR2X4 U164 ( .A(n10), .B(n115), .Y(n113) );
  XNOR2X4 U165 ( .A(n113), .B(n114), .Y(out[15]) );
  XOR2X1 U166 ( .A(n117), .B(n118), .Y(N33) );
  XOR2X1 U167 ( .A(n20), .B(sub_add_52_b0_carry[16]), .Y(N21) );
  AND2X1 U168 ( .A(sub_add_52_b0_carry[15]), .B(n122), .Y(
        sub_add_52_b0_carry[16]) );
  XOR2X1 U169 ( .A(n122), .B(sub_add_52_b0_carry[15]), .Y(N20) );
  AND2X1 U170 ( .A(sub_add_52_b0_carry[14]), .B(n121), .Y(
        sub_add_52_b0_carry[15]) );
  XOR2X1 U171 ( .A(n121), .B(sub_add_52_b0_carry[14]), .Y(N19) );
  AND2X1 U172 ( .A(sub_add_52_b0_carry[13]), .B(n120), .Y(
        sub_add_52_b0_carry[14]) );
endmodule


module multi16_4_DW01_add_0 ( A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, 
        A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, 
        B_20_, B_19_, B_18_, B_17_, B_16_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, 
        SUM_17_, SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, 
        SUM_9_, SUM_8_, SUM_7_, SUM_6_, SUM_5_ );
  input A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_,
         A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, B_20_, B_19_,
         B_18_, B_17_, B_16_;
  output SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, SUM_15_,
         SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, SUM_7_,
         SUM_6_, SUM_5_;
  wire   n1, n2, n3, n4, n5, n6, n7, n9, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41;

  CLKINVX4 U2 ( .A(n25), .Y(SUM_15_) );
  NAND2X2 U3 ( .A(B_19_), .B(A_19_), .Y(n33) );
  INVX2 U4 ( .A(n37), .Y(n24) );
  NOR2BX2 U5 ( .AN(n33), .B(n32), .Y(n40) );
  NAND2X2 U6 ( .A(n3), .B(n1), .Y(n2) );
  NAND2X1 U7 ( .A(B_18_), .B(A_18_), .Y(n36) );
  BUFX3 U8 ( .A(A_12_), .Y(SUM_12_) );
  BUFX3 U9 ( .A(A_13_), .Y(SUM_13_) );
  BUFX3 U10 ( .A(A_14_), .Y(SUM_14_) );
  INVX1 U11 ( .A(n34), .Y(n23) );
  AND2X2 U12 ( .A(n37), .B(n7), .Y(SUM_16_) );
  OAI21XL U13 ( .A0(n31), .A1(n32), .B0(n33), .Y(n28) );
  OR2X2 U14 ( .A(B_18_), .B(A_18_), .Y(n1) );
  NOR2X4 U15 ( .A(A_17_), .B(B_17_), .Y(n34) );
  NAND2X1 U16 ( .A(B_16_), .B(A_16_), .Y(n37) );
  CLKINVX4 U17 ( .A(n3), .Y(n4) );
  INVX1 U18 ( .A(n38), .Y(n22) );
  NAND2BX2 U19 ( .AN(n34), .B(n38), .Y(n5) );
  OR2X2 U20 ( .A(A_16_), .B(B_16_), .Y(n7) );
  XOR2X4 U21 ( .A(n6), .B(n4), .Y(SUM_18_) );
  NOR2X2 U22 ( .A(B_19_), .B(A_19_), .Y(n32) );
  INVX3 U23 ( .A(n41), .Y(n3) );
  AOI21X2 U24 ( .A0(n24), .A1(n23), .B0(n22), .Y(n41) );
  NAND2X4 U25 ( .A(n2), .B(n36), .Y(n39) );
  XOR2X4 U26 ( .A(n39), .B(n40), .Y(SUM_19_) );
  NAND2X2 U27 ( .A(B_17_), .B(A_17_), .Y(n38) );
  NAND2X2 U28 ( .A(n36), .B(n1), .Y(n6) );
  AND2X2 U29 ( .A(n30), .B(n29), .Y(n9) );
  XNOR2X4 U30 ( .A(n24), .B(n5), .Y(SUM_17_) );
  XOR2X1 U31 ( .A(n9), .B(n28), .Y(SUM_20_) );
  INVXL U32 ( .A(n30), .Y(n20) );
  OR2X2 U33 ( .A(B_20_), .B(A_20_), .Y(n29) );
  AOI21XL U34 ( .A0(n28), .A1(n29), .B0(n20), .Y(n27) );
  CLKINVX2 U35 ( .A(A_15_), .Y(n25) );
  INVXL U36 ( .A(n36), .Y(n21) );
  BUFX3 U37 ( .A(A_5_), .Y(SUM_5_) );
  BUFX3 U38 ( .A(A_7_), .Y(SUM_7_) );
  BUFX3 U39 ( .A(A_8_), .Y(SUM_8_) );
  BUFX3 U40 ( .A(A_6_), .Y(SUM_6_) );
  BUFX3 U41 ( .A(A_10_), .Y(SUM_10_) );
  BUFX3 U42 ( .A(A_11_), .Y(SUM_11_) );
  BUFX3 U43 ( .A(A_9_), .Y(SUM_9_) );
  XOR2X1 U44 ( .A(n26), .B(n27), .Y(SUM_21_) );
  XNOR2X1 U45 ( .A(B_21_), .B(A_21_), .Y(n26) );
  AOI21X1 U46 ( .A0(n1), .A1(n35), .B0(n21), .Y(n31) );
  OAI21XL U47 ( .A0(n34), .A1(n37), .B0(n38), .Y(n35) );
  NAND2X1 U48 ( .A(B_20_), .B(A_20_), .Y(n30) );
endmodule


module multi16_4_DW02_mult_0 ( A, B, PRODUCT_23_, PRODUCT_22_, PRODUCT_21_, 
        PRODUCT_20_, PRODUCT_19_, PRODUCT_18_, PRODUCT_17_, PRODUCT_16_, 
        PRODUCT_15_, PRODUCT_14_, PRODUCT_13_, PRODUCT_12_, PRODUCT_11_, 
        PRODUCT_10_, PRODUCT_9_, PRODUCT_8_, PRODUCT_7_ );
  input [16:0] A;
  input [7:0] B;
  output PRODUCT_23_, PRODUCT_22_, PRODUCT_21_, PRODUCT_20_, PRODUCT_19_,
         PRODUCT_18_, PRODUCT_17_, PRODUCT_16_, PRODUCT_15_, PRODUCT_14_,
         PRODUCT_13_, PRODUCT_12_, PRODUCT_11_, PRODUCT_10_, PRODUCT_9_,
         PRODUCT_8_, PRODUCT_7_;
  wire   ab_16__7_, ab_16__6_, ab_16__5_, ab_16__4_, ab_16__3_, ab_16__2_,
         ab_16__1_, ab_16__0_, ab_15__7_, ab_15__6_, ab_15__5_, ab_15__4_,
         ab_15__3_, ab_15__2_, ab_15__1_, ab_15__0_, ab_14__7_, ab_14__6_,
         ab_14__5_, ab_14__4_, ab_14__3_, ab_14__2_, ab_14__1_, ab_14__0_,
         ab_13__7_, ab_13__6_, ab_13__5_, ab_13__4_, ab_13__3_, ab_13__2_,
         ab_13__1_, ab_13__0_, ab_12__7_, ab_12__6_, ab_12__5_, ab_12__4_,
         ab_12__3_, ab_12__2_, ab_12__1_, ab_12__0_, ab_11__7_, ab_11__6_,
         ab_11__5_, ab_11__4_, ab_11__3_, ab_11__2_, ab_11__1_, ab_11__0_,
         ab_10__7_, ab_10__6_, ab_10__5_, ab_10__4_, ab_10__3_, ab_10__2_,
         ab_10__1_, ab_10__0_, ab_9__7_, ab_9__6_, ab_9__5_, ab_9__4_,
         ab_9__3_, ab_9__2_, ab_9__1_, ab_9__0_, ab_8__7_, ab_8__6_, ab_8__5_,
         ab_8__4_, ab_8__3_, ab_8__2_, ab_8__1_, ab_8__0_, ab_7__7_, ab_7__6_,
         ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_, ab_7__0_, ab_6__7_,
         ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_, ab_6__1_, ab_6__0_,
         ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_, ab_5__2_, ab_5__1_,
         ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_, ab_4__3_, ab_4__2_,
         ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_, ab_3__4_, ab_3__3_,
         ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_, ab_2__5_, ab_2__4_,
         ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_, ab_1__6_, ab_1__5_,
         ab_1__4_, ab_1__3_, ab_1__2_, ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_,
         ab_0__3_, ab_0__2_, CARRYB_16__6_, CARRYB_16__5_, CARRYB_16__4_,
         CARRYB_16__3_, CARRYB_16__2_, CARRYB_16__1_, CARRYB_16__0_,
         CARRYB_15__6_, CARRYB_15__5_, CARRYB_15__4_, CARRYB_15__3_,
         CARRYB_15__2_, CARRYB_15__1_, CARRYB_15__0_, CARRYB_14__6_,
         CARRYB_14__5_, CARRYB_14__4_, CARRYB_14__3_, CARRYB_14__2_,
         CARRYB_14__1_, CARRYB_14__0_, CARRYB_13__6_, CARRYB_13__5_,
         CARRYB_13__4_, CARRYB_13__3_, CARRYB_13__2_, CARRYB_13__1_,
         CARRYB_13__0_, CARRYB_12__6_, CARRYB_12__5_, CARRYB_12__4_,
         CARRYB_12__3_, CARRYB_12__2_, CARRYB_12__1_, CARRYB_12__0_,
         CARRYB_11__6_, CARRYB_11__5_, CARRYB_11__4_, CARRYB_11__3_,
         CARRYB_11__2_, CARRYB_11__1_, CARRYB_11__0_, CARRYB_10__6_,
         CARRYB_10__5_, CARRYB_10__4_, CARRYB_10__3_, CARRYB_10__2_,
         CARRYB_10__1_, CARRYB_10__0_, CARRYB_9__6_, CARRYB_9__5_,
         CARRYB_9__4_, CARRYB_9__3_, CARRYB_9__2_, CARRYB_9__1_, CARRYB_9__0_,
         CARRYB_8__6_, CARRYB_8__5_, CARRYB_8__4_, CARRYB_8__3_, CARRYB_8__2_,
         CARRYB_8__1_, CARRYB_8__0_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_,
         CARRYB_7__3_, CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_,
         CARRYB_6__5_, CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_,
         CARRYB_6__0_, CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_,
         CARRYB_5__2_, CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_,
         CARRYB_4__4_, CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_,
         CARRYB_3__6_, CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_,
         CARRYB_3__1_, CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_,
         CARRYB_2__3_, CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__1_,
         CARRYB_1__0_, SUMB_16__6_, SUMB_16__5_, SUMB_16__4_, SUMB_16__3_,
         SUMB_16__2_, SUMB_16__1_, SUMB_16__0_, SUMB_15__6_, SUMB_15__5_,
         SUMB_15__4_, SUMB_15__3_, SUMB_15__2_, SUMB_15__1_, SUMB_14__6_,
         SUMB_14__5_, SUMB_14__4_, SUMB_14__3_, SUMB_14__2_, SUMB_14__1_,
         SUMB_13__6_, SUMB_13__5_, SUMB_13__4_, SUMB_13__3_, SUMB_13__2_,
         SUMB_13__1_, SUMB_12__6_, SUMB_12__5_, SUMB_12__4_, SUMB_12__3_,
         SUMB_12__2_, SUMB_12__1_, SUMB_11__6_, SUMB_11__5_, SUMB_11__4_,
         SUMB_11__3_, SUMB_11__2_, SUMB_11__1_, SUMB_10__6_, SUMB_10__5_,
         SUMB_10__4_, SUMB_10__3_, SUMB_10__2_, SUMB_10__1_, SUMB_9__6_,
         SUMB_9__5_, SUMB_9__4_, SUMB_9__3_, SUMB_9__2_, SUMB_9__1_,
         SUMB_8__6_, SUMB_8__5_, SUMB_8__4_, SUMB_8__3_, SUMB_8__2_,
         SUMB_8__1_, SUMB_7__6_, SUMB_7__5_, SUMB_7__4_, SUMB_7__3_,
         SUMB_7__2_, SUMB_7__1_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_,
         SUMB_6__3_, SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_,
         SUMB_5__4_, SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_,
         SUMB_4__5_, SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_,
         SUMB_3__6_, SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_,
         SUMB_3__1_, SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_,
         SUMB_2__2_, SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_,
         SUMB_1__3_, SUMB_1__2_, SUMB_1__1_, PROD1_7_, A1_21_, A1_20_, A1_19_,
         A1_18_, A1_17_, A1_16_, A1_15_, A1_13_, A1_12_, A1_11_, A1_10_, A1_9_,
         A1_8_, A1_7_, A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, n4, n5, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41;

  ADDFHX4 S2_15_1 ( .A(ab_15__1_), .B(CARRYB_14__1_), .CI(SUMB_14__2_), .CO(
        CARRYB_15__1_), .S(SUMB_15__1_) );
  ADDFHX4 S1_14_0 ( .A(ab_14__0_), .B(CARRYB_13__0_), .CI(SUMB_13__1_), .CO(
        CARRYB_14__0_), .S(A1_12_) );
  ADDFHX4 S2_14_1 ( .A(ab_14__1_), .B(CARRYB_13__1_), .CI(SUMB_13__2_), .CO(
        CARRYB_14__1_), .S(SUMB_14__1_) );
  ADDFHX4 S1_13_0 ( .A(ab_13__0_), .B(CARRYB_12__0_), .CI(SUMB_12__1_), .CO(
        CARRYB_13__0_), .S(A1_11_) );
  ADDFHX4 S2_13_1 ( .A(ab_13__1_), .B(CARRYB_12__1_), .CI(SUMB_12__2_), .CO(
        CARRYB_13__1_), .S(SUMB_13__1_) );
  ADDFHX4 S2_12_1 ( .A(ab_12__1_), .B(CARRYB_11__1_), .CI(SUMB_11__2_), .CO(
        CARRYB_12__1_), .S(SUMB_12__1_) );
  ADDFHX4 S2_12_2 ( .A(ab_12__2_), .B(CARRYB_11__2_), .CI(SUMB_11__3_), .CO(
        CARRYB_12__2_), .S(SUMB_12__2_) );
  ADDFHX4 S2_12_3 ( .A(ab_12__3_), .B(CARRYB_11__3_), .CI(SUMB_11__4_), .CO(
        CARRYB_12__3_), .S(SUMB_12__3_) );
  ADDFHX4 S2_12_4 ( .A(ab_12__4_), .B(CARRYB_11__4_), .CI(SUMB_11__5_), .CO(
        CARRYB_12__4_), .S(SUMB_12__4_) );
  ADDFHX4 S1_11_0 ( .A(ab_11__0_), .B(CARRYB_10__0_), .CI(SUMB_10__1_), .CO(
        CARRYB_11__0_), .S(A1_9_) );
  ADDFHX4 S2_11_1 ( .A(ab_11__1_), .B(CARRYB_10__1_), .CI(SUMB_10__2_), .CO(
        CARRYB_11__1_), .S(SUMB_11__1_) );
  ADDFHX4 S2_11_2 ( .A(ab_11__2_), .B(CARRYB_10__2_), .CI(SUMB_10__3_), .CO(
        CARRYB_11__2_), .S(SUMB_11__2_) );
  ADDFHX4 S2_11_3 ( .A(ab_11__3_), .B(CARRYB_10__3_), .CI(SUMB_10__4_), .CO(
        CARRYB_11__3_), .S(SUMB_11__3_) );
  ADDFHX4 S1_10_0 ( .A(ab_10__0_), .B(CARRYB_9__0_), .CI(SUMB_9__1_), .CO(
        CARRYB_10__0_), .S(A1_8_) );
  ADDFHX4 S2_10_1 ( .A(ab_10__1_), .B(CARRYB_9__1_), .CI(SUMB_9__2_), .CO(
        CARRYB_10__1_), .S(SUMB_10__1_) );
  ADDFHX4 S2_9_1 ( .A(ab_9__1_), .B(CARRYB_8__1_), .CI(SUMB_8__2_), .CO(
        CARRYB_9__1_), .S(SUMB_9__1_) );
  ADDFHX4 S2_9_2 ( .A(ab_9__2_), .B(CARRYB_8__2_), .CI(SUMB_8__3_), .CO(
        CARRYB_9__2_), .S(SUMB_9__2_) );
  ADDFHX4 S2_9_3 ( .A(ab_9__3_), .B(CARRYB_8__3_), .CI(SUMB_8__4_), .CO(
        CARRYB_9__3_), .S(SUMB_9__3_) );
  ADDFHX4 S2_9_4 ( .A(ab_9__4_), .B(CARRYB_8__4_), .CI(SUMB_8__5_), .CO(
        CARRYB_9__4_), .S(SUMB_9__4_) );
  ADDFHX4 S2_8_1 ( .A(ab_8__1_), .B(CARRYB_7__1_), .CI(SUMB_7__2_), .CO(
        CARRYB_8__1_), .S(SUMB_8__1_) );
  ADDFHX4 S2_8_2 ( .A(ab_8__2_), .B(CARRYB_7__2_), .CI(SUMB_7__3_), .CO(
        CARRYB_8__2_), .S(SUMB_8__2_) );
  ADDFHX4 S2_8_3 ( .A(ab_8__3_), .B(CARRYB_7__3_), .CI(SUMB_7__4_), .CO(
        CARRYB_8__3_), .S(SUMB_8__3_) );
  ADDFHX4 S2_8_4 ( .A(ab_8__4_), .B(CARRYB_7__4_), .CI(SUMB_7__5_), .CO(
        CARRYB_8__4_), .S(SUMB_8__4_) );
  ADDFHX4 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  ADDFHX4 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  ADDFHX4 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  ADDFHX4 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  multi16_4_DW01_add_0 FS_1 ( .A_21_(A1_21_), .A_20_(A1_20_), .A_19_(A1_19_), 
        .A_18_(A1_18_), .A_17_(A1_17_), .A_16_(A1_16_), .A_15_(A1_15_), 
        .A_14_(SUMB_16__0_), .A_13_(A1_13_), .A_12_(A1_12_), .A_11_(A1_11_), 
        .A_10_(A1_10_), .A_9_(A1_9_), .A_8_(A1_8_), .A_7_(A1_7_), .A_6_(A1_6_), 
        .A_5_(PROD1_7_), .B_21_(n10), .B_20_(n22), .B_19_(n21), .B_18_(n20), 
        .B_17_(n4), .B_16_(n19), .SUM_21_(PRODUCT_23_), .SUM_20_(PRODUCT_22_), 
        .SUM_19_(PRODUCT_21_), .SUM_18_(PRODUCT_20_), .SUM_17_(PRODUCT_19_), 
        .SUM_16_(PRODUCT_18_), .SUM_15_(PRODUCT_17_), .SUM_14_(PRODUCT_16_), 
        .SUM_13_(PRODUCT_15_), .SUM_12_(PRODUCT_14_), .SUM_11_(PRODUCT_13_), 
        .SUM_10_(PRODUCT_12_), .SUM_9_(PRODUCT_11_), .SUM_8_(PRODUCT_10_), 
        .SUM_7_(PRODUCT_9_), .SUM_6_(PRODUCT_8_), .SUM_5_(PRODUCT_7_) );
  ADDFHX1 S3_15_6 ( .A(ab_15__6_), .B(CARRYB_14__6_), .CI(ab_14__7_), .CO(
        CARRYB_15__6_), .S(SUMB_15__6_) );
  ADDFHX1 S3_14_6 ( .A(ab_14__6_), .B(CARRYB_13__6_), .CI(ab_13__7_), .CO(
        CARRYB_14__6_), .S(SUMB_14__6_) );
  ADDFX2 S5_6 ( .A(ab_16__6_), .B(CARRYB_15__6_), .CI(ab_15__7_), .CO(
        CARRYB_16__6_), .S(SUMB_16__6_) );
  ADDFX2 S4_5 ( .A(ab_16__5_), .B(CARRYB_15__5_), .CI(SUMB_15__6_), .CO(
        CARRYB_16__5_), .S(SUMB_16__5_) );
  ADDFHX1 S3_13_6 ( .A(ab_13__6_), .B(CARRYB_12__6_), .CI(ab_12__7_), .CO(
        CARRYB_13__6_), .S(SUMB_13__6_) );
  ADDFHX2 S2_14_5 ( .A(ab_14__5_), .B(CARRYB_13__5_), .CI(SUMB_13__6_), .CO(
        CARRYB_14__5_), .S(SUMB_14__5_) );
  ADDFHX4 S2_14_2 ( .A(ab_14__2_), .B(CARRYB_13__2_), .CI(SUMB_13__3_), .CO(
        CARRYB_14__2_), .S(SUMB_14__2_) );
  ADDFHX4 S3_7_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(
        CARRYB_7__6_), .S(SUMB_7__6_) );
  ADDFHX4 S3_8_6 ( .A(ab_8__6_), .B(CARRYB_7__6_), .CI(ab_7__7_), .CO(
        CARRYB_8__6_), .S(SUMB_8__6_) );
  ADDFHX2 S3_2_6 ( .A(ab_2__6_), .B(n5), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  ADDFHX2 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  ADDFHX4 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  ADDFHX2 S4_4 ( .A(ab_16__4_), .B(CARRYB_15__4_), .CI(SUMB_15__5_), .CO(
        CARRYB_16__4_), .S(SUMB_16__4_) );
  ADDFHX2 S2_2_4 ( .A(ab_2__4_), .B(n7), .CI(SUMB_1__5_), .CO(CARRYB_2__4_), 
        .S(SUMB_2__4_) );
  ADDFHX4 S1_8_0 ( .A(ab_8__0_), .B(CARRYB_7__0_), .CI(SUMB_7__1_), .CO(
        CARRYB_8__0_), .S(A1_6_) );
  ADDFHX4 S2_7_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  ADDFHX4 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  ADDFHX2 S2_15_4 ( .A(ab_15__4_), .B(CARRYB_14__4_), .CI(SUMB_14__5_), .CO(
        CARRYB_15__4_), .S(SUMB_15__4_) );
  ADDFHX4 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  ADDFHX2 S4_0 ( .A(ab_16__0_), .B(CARRYB_15__0_), .CI(SUMB_15__1_), .CO(
        CARRYB_16__0_), .S(SUMB_16__0_) );
  ADDFHX4 S4_3 ( .A(ab_16__3_), .B(CARRYB_15__3_), .CI(SUMB_15__4_), .CO(
        CARRYB_16__3_), .S(SUMB_16__3_) );
  ADDFHX4 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  ADDFHX2 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  ADDFHX4 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  ADDFHX2 S2_2_5 ( .A(ab_2__5_), .B(n8), .CI(SUMB_1__6_), .CO(CARRYB_2__5_), 
        .S(SUMB_2__5_) );
  ADDFHX4 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  ADDFHX4 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  ADDFHX2 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  ADDFHX4 S2_8_5 ( .A(ab_8__5_), .B(CARRYB_7__5_), .CI(SUMB_7__6_), .CO(
        CARRYB_8__5_), .S(SUMB_8__5_) );
  ADDFHX4 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  ADDFHX4 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  ADDFHX4 S2_11_4 ( .A(ab_11__4_), .B(CARRYB_10__4_), .CI(SUMB_10__5_), .CO(
        CARRYB_11__4_), .S(SUMB_11__4_) );
  ADDFHX4 S2_10_5 ( .A(ab_10__5_), .B(CARRYB_9__5_), .CI(SUMB_9__6_), .CO(
        CARRYB_10__5_), .S(SUMB_10__5_) );
  ADDFHX4 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  ADDFHX4 S2_15_3 ( .A(ab_15__3_), .B(CARRYB_14__3_), .CI(SUMB_14__4_), .CO(
        CARRYB_15__3_), .S(SUMB_15__3_) );
  ADDFHX4 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  ADDFHX4 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  ADDFHX4 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  ADDFHX2 S4_1 ( .A(ab_16__1_), .B(CARRYB_15__1_), .CI(SUMB_15__2_), .CO(
        CARRYB_16__1_), .S(SUMB_16__1_) );
  ADDFHX4 S2_9_5 ( .A(ab_9__5_), .B(CARRYB_8__5_), .CI(SUMB_8__6_), .CO(
        CARRYB_9__5_), .S(SUMB_9__5_) );
  ADDFHX4 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  ADDFHX4 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  ADDFHX4 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  ADDFHX2 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  ADDFHX2 S1_7_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(PROD1_7_) );
  ADDFHX2 S3_12_6 ( .A(ab_12__6_), .B(CARRYB_11__6_), .CI(ab_11__7_), .CO(
        CARRYB_12__6_), .S(SUMB_12__6_) );
  ADDFHX1 S2_15_5 ( .A(ab_15__5_), .B(CARRYB_14__5_), .CI(SUMB_14__6_), .CO(
        CARRYB_15__5_), .S(SUMB_15__5_) );
  ADDFHX2 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  ADDFHX2 S2_2_2 ( .A(ab_2__2_), .B(n6), .CI(SUMB_1__3_), .CO(CARRYB_2__2_), 
        .S(SUMB_2__2_) );
  ADDFHX2 S4_2 ( .A(ab_16__2_), .B(CARRYB_15__2_), .CI(SUMB_15__3_), .CO(
        CARRYB_16__2_), .S(SUMB_16__2_) );
  ADDFHX2 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  ADDFHX2 S1_9_0 ( .A(ab_9__0_), .B(CARRYB_8__0_), .CI(SUMB_8__1_), .CO(
        CARRYB_9__0_), .S(A1_7_) );
  ADDFHX2 S1_12_0 ( .A(ab_12__0_), .B(CARRYB_11__0_), .CI(SUMB_11__1_), .CO(
        CARRYB_12__0_), .S(A1_10_) );
  ADDFHX2 S1_15_0 ( .A(ab_15__0_), .B(CARRYB_14__0_), .CI(SUMB_14__1_), .CO(
        CARRYB_15__0_), .S(A1_13_) );
  ADDFHX2 S2_14_4 ( .A(ab_14__4_), .B(CARRYB_13__4_), .CI(SUMB_13__5_), .CO(
        CARRYB_14__4_), .S(SUMB_14__4_) );
  ADDFHX2 S2_11_5 ( .A(ab_11__5_), .B(CARRYB_10__5_), .CI(SUMB_10__6_), .CO(
        CARRYB_11__5_), .S(SUMB_11__5_) );
  ADDFHX2 S2_10_2 ( .A(ab_10__2_), .B(CARRYB_9__2_), .CI(SUMB_9__3_), .CO(
        CARRYB_10__2_), .S(SUMB_10__2_) );
  ADDFHX2 S2_7_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  ADDFHX2 S2_10_4 ( .A(ab_10__4_), .B(CARRYB_9__4_), .CI(SUMB_9__5_), .CO(
        CARRYB_10__4_), .S(SUMB_10__4_) );
  ADDFHX2 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  ADDFHX2 S2_7_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  ADDFHX2 S2_13_5 ( .A(ab_13__5_), .B(SUMB_12__6_), .CI(CARRYB_12__5_), .CO(
        CARRYB_13__5_), .S(SUMB_13__5_) );
  ADDFHX2 S3_9_6 ( .A(ab_9__6_), .B(CARRYB_8__6_), .CI(ab_8__7_), .CO(
        CARRYB_9__6_), .S(SUMB_9__6_) );
  ADDFHX2 S2_15_2 ( .A(ab_15__2_), .B(CARRYB_14__2_), .CI(SUMB_14__3_), .CO(
        CARRYB_15__2_), .S(SUMB_15__2_) );
  ADDFHX1 S2_12_5 ( .A(ab_12__5_), .B(CARRYB_11__5_), .CI(SUMB_11__6_), .CO(
        CARRYB_12__5_), .S(SUMB_12__5_) );
  ADDFHX2 S2_14_3 ( .A(ab_14__3_), .B(CARRYB_13__3_), .CI(SUMB_13__4_), .CO(
        CARRYB_14__3_), .S(SUMB_14__3_) );
  ADDFHX4 S3_11_6 ( .A(ab_11__6_), .B(CARRYB_10__6_), .CI(ab_10__7_), .CO(
        CARRYB_11__6_), .S(SUMB_11__6_) );
  ADDFHX4 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  ADDFHX4 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  ADDFHX4 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  ADDFHX4 S2_7_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  ADDFHX4 S2_13_2 ( .A(ab_13__2_), .B(CARRYB_12__2_), .CI(SUMB_12__3_), .CO(
        CARRYB_13__2_), .S(SUMB_13__2_) );
  ADDFHX4 S2_13_3 ( .A(ab_13__3_), .B(CARRYB_12__3_), .CI(SUMB_12__4_), .CO(
        CARRYB_13__3_), .S(SUMB_13__3_) );
  ADDFHX4 S2_13_4 ( .A(ab_13__4_), .B(CARRYB_12__4_), .CI(SUMB_12__5_), .CO(
        CARRYB_13__4_), .S(SUMB_13__4_) );
  ADDFHX4 S2_7_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  ADDFHX4 S2_10_3 ( .A(ab_10__3_), .B(CARRYB_9__3_), .CI(SUMB_9__4_), .CO(
        CARRYB_10__3_), .S(SUMB_10__3_) );
  ADDFHX2 S2_2_3 ( .A(ab_2__3_), .B(n9), .CI(SUMB_1__4_), .CO(CARRYB_2__3_), 
        .S(SUMB_2__3_) );
  CLKINVX3 U2 ( .A(SUMB_16__2_), .Y(n12) );
  NAND3X4 U3 ( .A(n18), .B(n16), .C(n17), .Y(CARRYB_10__6_) );
  AND2X1 U4 ( .A(A[2]), .B(B[2]), .Y(ab_2__2_) );
  AND2X2 U5 ( .A(A[2]), .B(B[6]), .Y(ab_2__6_) );
  NOR2X4 U6 ( .A(n32), .B(n25), .Y(ab_0__2_) );
  INVX3 U7 ( .A(B[2]), .Y(n32) );
  XOR2X1 U8 ( .A(ab_1__5_), .B(ab_0__6_), .Y(SUMB_1__5_) );
  AND2X2 U9 ( .A(CARRYB_16__2_), .B(SUMB_16__3_), .Y(n20) );
  NAND2X1 U10 ( .A(n13), .B(n14), .Y(A1_16_) );
  NAND2X2 U11 ( .A(CARRYB_16__1_), .B(n12), .Y(n13) );
  NAND2X1 U12 ( .A(ab_9__7_), .B(CARRYB_9__6_), .Y(n17) );
  NAND2X1 U13 ( .A(ab_10__6_), .B(CARRYB_9__6_), .Y(n16) );
  XOR2X1 U14 ( .A(CARRYB_16__5_), .B(SUMB_16__6_), .Y(A1_20_) );
  AND2X2 U16 ( .A(CARRYB_16__1_), .B(SUMB_16__2_), .Y(n4) );
  AND2X2 U17 ( .A(ab_0__7_), .B(ab_1__6_), .Y(n5) );
  AND2X2 U18 ( .A(ab_0__3_), .B(ab_1__2_), .Y(n6) );
  AND2X2 U19 ( .A(ab_0__5_), .B(ab_1__4_), .Y(n7) );
  AND2X2 U20 ( .A(ab_0__6_), .B(ab_1__5_), .Y(n8) );
  AND2X2 U21 ( .A(ab_0__4_), .B(ab_1__3_), .Y(n9) );
  AND2X2 U22 ( .A(CARRYB_16__5_), .B(SUMB_16__6_), .Y(n10) );
  NOR2X2 U23 ( .A(n34), .B(n25), .Y(ab_0__7_) );
  NOR2X2 U24 ( .A(n30), .B(n25), .Y(ab_0__4_) );
  INVX1 U25 ( .A(A[0]), .Y(n25) );
  INVX2 U26 ( .A(n23), .Y(CARRYB_1__1_) );
  NAND2X2 U27 ( .A(n11), .B(SUMB_16__2_), .Y(n14) );
  CLKINVX3 U28 ( .A(CARRYB_16__1_), .Y(n11) );
  AND2X1 U29 ( .A(A[3]), .B(B[5]), .Y(ab_3__5_) );
  AND2X1 U30 ( .A(A[1]), .B(B[5]), .Y(ab_1__5_) );
  NOR2XL U31 ( .A(n36), .B(n34), .Y(ab_16__7_) );
  INVX4 U32 ( .A(B[5]), .Y(n29) );
  XOR2X2 U33 ( .A(CARRYB_16__4_), .B(SUMB_16__5_), .Y(A1_19_) );
  NOR2X4 U34 ( .A(n28), .B(n25), .Y(ab_0__6_) );
  INVX3 U35 ( .A(B[6]), .Y(n28) );
  AND2X1 U36 ( .A(A[1]), .B(B[4]), .Y(ab_1__4_) );
  INVX4 U37 ( .A(B[4]), .Y(n30) );
  AND2X2 U38 ( .A(A[1]), .B(B[2]), .Y(ab_1__2_) );
  XOR2X1 U39 ( .A(CARRYB_16__0_), .B(SUMB_16__1_), .Y(A1_15_) );
  XOR2X1 U40 ( .A(ab_1__6_), .B(ab_0__7_), .Y(SUMB_1__6_) );
  XOR2X4 U41 ( .A(CARRYB_16__2_), .B(SUMB_16__3_), .Y(A1_17_) );
  NAND2X1 U42 ( .A(ab_0__2_), .B(n35), .Y(n23) );
  NOR2X2 U43 ( .A(n31), .B(n25), .Y(ab_0__3_) );
  NOR2X2 U44 ( .A(n29), .B(n25), .Y(ab_0__5_) );
  INVX2 U45 ( .A(B[3]), .Y(n31) );
  XOR2XL U46 ( .A(ab_10__6_), .B(ab_9__7_), .Y(n15) );
  XOR2X1 U47 ( .A(CARRYB_9__6_), .B(n15), .Y(SUMB_10__6_) );
  NAND2XL U48 ( .A(ab_9__7_), .B(ab_10__6_), .Y(n18) );
  NOR2XL U49 ( .A(n40), .B(n29), .Y(ab_12__5_) );
  INVX4 U50 ( .A(B[7]), .Y(n34) );
  NAND2XL U51 ( .A(A[1]), .B(B[1]), .Y(n27) );
  AND2X2 U52 ( .A(A[2]), .B(B[0]), .Y(ab_2__0_) );
  AND2X2 U53 ( .A(CARRYB_16__0_), .B(SUMB_16__1_), .Y(n19) );
  INVXL U54 ( .A(B[0]), .Y(n24) );
  AND2X1 U55 ( .A(A[9]), .B(B[0]), .Y(ab_9__0_) );
  AND2X1 U56 ( .A(A[8]), .B(B[0]), .Y(ab_8__0_) );
  AND2X1 U57 ( .A(A[5]), .B(B[1]), .Y(ab_5__1_) );
  AND2X1 U58 ( .A(A[6]), .B(B[1]), .Y(ab_6__1_) );
  AND2X1 U59 ( .A(A[7]), .B(B[0]), .Y(ab_7__0_) );
  AND2X1 U60 ( .A(A[6]), .B(B[0]), .Y(ab_6__0_) );
  AND2X1 U61 ( .A(A[10]), .B(B[0]), .Y(ab_10__0_) );
  AND2X1 U62 ( .A(A[10]), .B(B[1]), .Y(ab_10__1_) );
  AND2X1 U63 ( .A(A[9]), .B(B[1]), .Y(ab_9__1_) );
  AND2X1 U64 ( .A(A[7]), .B(B[1]), .Y(ab_7__1_) );
  AND2X1 U65 ( .A(A[8]), .B(B[1]), .Y(ab_8__1_) );
  INVXL U66 ( .A(B[1]), .Y(n33) );
  AND2X1 U67 ( .A(A[10]), .B(B[5]), .Y(ab_10__5_) );
  NOR2X1 U68 ( .A(n41), .B(n29), .Y(ab_11__5_) );
  AND2X1 U69 ( .A(A[3]), .B(B[0]), .Y(ab_3__0_) );
  AND2X1 U70 ( .A(A[2]), .B(B[5]), .Y(ab_2__5_) );
  NOR2XL U71 ( .A(n39), .B(n33), .Y(ab_13__1_) );
  NOR2XL U72 ( .A(n40), .B(n33), .Y(ab_12__1_) );
  NOR2XL U73 ( .A(n41), .B(n33), .Y(ab_11__1_) );
  AND2X1 U74 ( .A(A[9]), .B(B[5]), .Y(ab_9__5_) );
  AND2X1 U75 ( .A(A[8]), .B(B[5]), .Y(ab_8__5_) );
  AND2X1 U76 ( .A(A[7]), .B(B[5]), .Y(ab_7__5_) );
  AND2X1 U77 ( .A(A[6]), .B(B[5]), .Y(ab_6__5_) );
  AND2X1 U78 ( .A(A[2]), .B(B[1]), .Y(ab_2__1_) );
  AND2X1 U79 ( .A(CARRYB_16__3_), .B(SUMB_16__4_), .Y(n21) );
  AND2X2 U80 ( .A(CARRYB_16__4_), .B(SUMB_16__5_), .Y(n22) );
  NOR2X1 U81 ( .A(n36), .B(n33), .Y(ab_16__1_) );
  NOR2X1 U82 ( .A(n36), .B(n29), .Y(ab_16__5_) );
  INVX1 U83 ( .A(n27), .Y(n35) );
  AND2X1 U84 ( .A(A[10]), .B(B[6]), .Y(ab_10__6_) );
  AND2X1 U85 ( .A(A[9]), .B(B[6]), .Y(ab_9__6_) );
  AND2X1 U86 ( .A(A[8]), .B(B[6]), .Y(ab_8__6_) );
  AND2X1 U87 ( .A(A[7]), .B(B[6]), .Y(ab_7__6_) );
  AND2X1 U88 ( .A(A[6]), .B(B[6]), .Y(ab_6__6_) );
  AND2X1 U89 ( .A(A[5]), .B(B[6]), .Y(ab_5__6_) );
  AND2X2 U90 ( .A(A[4]), .B(B[1]), .Y(ab_4__1_) );
  AND2X2 U91 ( .A(A[5]), .B(B[0]), .Y(ab_5__0_) );
  AND2X1 U92 ( .A(A[4]), .B(B[0]), .Y(ab_4__0_) );
  NOR2BX1 U93 ( .AN(B[0]), .B(n36), .Y(ab_16__0_) );
  XOR2X1 U94 ( .A(CARRYB_16__6_), .B(ab_16__7_), .Y(A1_21_) );
  XOR2X1 U95 ( .A(ab_1__4_), .B(ab_0__5_), .Y(SUMB_1__4_) );
  NOR2XL U96 ( .A(n37), .B(n34), .Y(ab_15__7_) );
  AND2X2 U97 ( .A(A[1]), .B(B[3]), .Y(ab_1__3_) );
  AND2X1 U98 ( .A(A[4]), .B(B[5]), .Y(ab_4__5_) );
  XOR2X1 U99 ( .A(n35), .B(ab_0__2_), .Y(SUMB_1__1_) );
  NOR2X1 U100 ( .A(n37), .B(n33), .Y(ab_15__1_) );
  NOR2X1 U101 ( .A(n38), .B(n33), .Y(ab_14__1_) );
  AND2X1 U102 ( .A(A[10]), .B(B[4]), .Y(ab_10__4_) );
  AND2X1 U103 ( .A(A[9]), .B(B[4]), .Y(ab_9__4_) );
  NOR2XL U104 ( .A(n39), .B(n29), .Y(ab_13__5_) );
  AND2X1 U105 ( .A(A[8]), .B(B[4]), .Y(ab_8__4_) );
  AND2X1 U106 ( .A(A[7]), .B(B[4]), .Y(ab_7__4_) );
  AND2X1 U107 ( .A(A[6]), .B(B[4]), .Y(ab_6__4_) );
  NOR2XL U108 ( .A(n41), .B(n34), .Y(ab_11__7_) );
  AND2X1 U109 ( .A(A[5]), .B(B[5]), .Y(ab_5__5_) );
  AND2X1 U110 ( .A(A[5]), .B(B[4]), .Y(ab_5__4_) );
  AND2X1 U111 ( .A(A[4]), .B(B[4]), .Y(ab_4__4_) );
  AND2X1 U112 ( .A(A[4]), .B(B[6]), .Y(ab_4__6_) );
  AND2X1 U113 ( .A(A[3]), .B(B[4]), .Y(ab_3__4_) );
  AND2X1 U114 ( .A(A[3]), .B(B[6]), .Y(ab_3__6_) );
  AND2X2 U115 ( .A(A[3]), .B(B[1]), .Y(ab_3__1_) );
  AND2X1 U116 ( .A(A[2]), .B(B[4]), .Y(ab_2__4_) );
  XOR2X1 U117 ( .A(ab_1__2_), .B(ab_0__3_), .Y(SUMB_1__2_) );
  XOR2X1 U118 ( .A(ab_1__3_), .B(ab_0__4_), .Y(SUMB_1__3_) );
  NOR2XL U119 ( .A(n38), .B(n29), .Y(ab_14__5_) );
  NOR2XL U120 ( .A(n37), .B(n29), .Y(ab_15__5_) );
  NOR2XL U121 ( .A(n40), .B(n34), .Y(ab_12__7_) );
  NOR2XL U122 ( .A(n39), .B(n34), .Y(ab_13__7_) );
  NOR2XL U123 ( .A(n38), .B(n34), .Y(ab_14__7_) );
  INVX1 U124 ( .A(A[16]), .Y(n36) );
  NAND2XL U125 ( .A(A[0]), .B(B[0]), .Y(n26) );
  INVX1 U126 ( .A(A[11]), .Y(n41) );
  INVX1 U127 ( .A(A[12]), .Y(n40) );
  INVX1 U128 ( .A(A[13]), .Y(n39) );
  INVX1 U129 ( .A(A[14]), .Y(n38) );
  INVX1 U130 ( .A(A[15]), .Y(n37) );
  XOR2X4 U131 ( .A(CARRYB_16__3_), .B(SUMB_16__4_), .Y(A1_18_) );
  NOR2XL U132 ( .A(n36), .B(n30), .Y(ab_16__4_) );
  NOR2XL U133 ( .A(n37), .B(n30), .Y(ab_15__4_) );
  NOR2XL U134 ( .A(n38), .B(n30), .Y(ab_14__4_) );
  NOR2XL U135 ( .A(n39), .B(n30), .Y(ab_13__4_) );
  NOR2XL U136 ( .A(n40), .B(n30), .Y(ab_12__4_) );
  NOR2XL U137 ( .A(n41), .B(n30), .Y(ab_11__4_) );
  NOR2XL U138 ( .A(n27), .B(n26), .Y(CARRYB_1__0_) );
  NOR2XL U139 ( .A(n36), .B(n32), .Y(ab_16__2_) );
  NOR2XL U140 ( .A(n37), .B(n32), .Y(ab_15__2_) );
  NOR2XL U141 ( .A(n38), .B(n32), .Y(ab_14__2_) );
  NOR2XL U142 ( .A(n39), .B(n32), .Y(ab_13__2_) );
  NOR2XL U143 ( .A(n40), .B(n32), .Y(ab_12__2_) );
  NOR2XL U144 ( .A(n41), .B(n32), .Y(ab_11__2_) );
  AND2X1 U145 ( .A(A[10]), .B(B[2]), .Y(ab_10__2_) );
  AND2X1 U146 ( .A(A[9]), .B(B[2]), .Y(ab_9__2_) );
  AND2X1 U147 ( .A(A[8]), .B(B[2]), .Y(ab_8__2_) );
  AND2X1 U148 ( .A(A[7]), .B(B[2]), .Y(ab_7__2_) );
  AND2X1 U149 ( .A(A[6]), .B(B[2]), .Y(ab_6__2_) );
  AND2X1 U150 ( .A(A[5]), .B(B[2]), .Y(ab_5__2_) );
  AND2X1 U151 ( .A(A[4]), .B(B[2]), .Y(ab_4__2_) );
  AND2X1 U152 ( .A(A[3]), .B(B[2]), .Y(ab_3__2_) );
  NOR2XL U153 ( .A(n36), .B(n31), .Y(ab_16__3_) );
  NOR2XL U154 ( .A(n37), .B(n31), .Y(ab_15__3_) );
  NOR2XL U155 ( .A(n38), .B(n31), .Y(ab_14__3_) );
  NOR2XL U156 ( .A(n39), .B(n31), .Y(ab_13__3_) );
  NOR2XL U157 ( .A(n40), .B(n31), .Y(ab_12__3_) );
  NOR2XL U158 ( .A(n41), .B(n31), .Y(ab_11__3_) );
  AND2X1 U159 ( .A(A[10]), .B(B[3]), .Y(ab_10__3_) );
  AND2X1 U160 ( .A(A[9]), .B(B[3]), .Y(ab_9__3_) );
  AND2X1 U161 ( .A(A[8]), .B(B[3]), .Y(ab_8__3_) );
  AND2X1 U162 ( .A(A[7]), .B(B[3]), .Y(ab_7__3_) );
  AND2X1 U163 ( .A(A[6]), .B(B[3]), .Y(ab_6__3_) );
  AND2X1 U164 ( .A(A[5]), .B(B[3]), .Y(ab_5__3_) );
  AND2X1 U165 ( .A(A[4]), .B(B[3]), .Y(ab_4__3_) );
  AND2X1 U166 ( .A(A[3]), .B(B[3]), .Y(ab_3__3_) );
  AND2X1 U167 ( .A(A[2]), .B(B[3]), .Y(ab_2__3_) );
  NOR2XL U168 ( .A(n36), .B(n28), .Y(ab_16__6_) );
  NOR2XL U169 ( .A(n37), .B(n28), .Y(ab_15__6_) );
  NOR2XL U170 ( .A(n38), .B(n28), .Y(ab_14__6_) );
  NOR2XL U171 ( .A(n39), .B(n28), .Y(ab_13__6_) );
  NOR2XL U172 ( .A(n40), .B(n28), .Y(ab_12__6_) );
  NOR2XL U173 ( .A(n41), .B(n28), .Y(ab_11__6_) );
  AND2X1 U174 ( .A(A[10]), .B(B[7]), .Y(ab_10__7_) );
  AND2X1 U175 ( .A(A[9]), .B(B[7]), .Y(ab_9__7_) );
  AND2X1 U176 ( .A(A[8]), .B(B[7]), .Y(ab_8__7_) );
  AND2X1 U177 ( .A(A[7]), .B(B[7]), .Y(ab_7__7_) );
  AND2X1 U178 ( .A(A[6]), .B(B[7]), .Y(ab_6__7_) );
  AND2X1 U179 ( .A(A[5]), .B(B[7]), .Y(ab_5__7_) );
  AND2X1 U180 ( .A(A[4]), .B(B[7]), .Y(ab_4__7_) );
  AND2X1 U181 ( .A(A[3]), .B(B[7]), .Y(ab_3__7_) );
  AND2X1 U182 ( .A(A[2]), .B(B[7]), .Y(ab_2__7_) );
  AND2X2 U183 ( .A(A[1]), .B(B[6]), .Y(ab_1__6_) );
  AND2X1 U184 ( .A(A[1]), .B(B[7]), .Y(ab_1__7_) );
  NOR2X1 U186 ( .A(n24), .B(n37), .Y(ab_15__0_) );
  NOR2X1 U187 ( .A(n24), .B(n38), .Y(ab_14__0_) );
  NOR2X1 U188 ( .A(n24), .B(n39), .Y(ab_13__0_) );
  NOR2X1 U189 ( .A(n24), .B(n40), .Y(ab_12__0_) );
  NOR2X1 U190 ( .A(n24), .B(n41), .Y(ab_11__0_) );
endmodule


module multi16_4 ( in_17bit, in_8bit, out );
  input [16:0] in_17bit;
  input [7:0] in_8bit;
  output [16:0] out;
  wire   N21, N33, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118;
  wire   [16:1] in_17bit_b;
  wire   [6:1] in_8bit_b;
  wire   [23:8] mul;
  wire   [16:12] sub_add_52_b0_carry;

  multi16_4_DW02_mult_0 mult_55 ( .A({in_17bit_b, in_17bit[0]}), .B({n10, 
        in_8bit_b, n26}), .PRODUCT_23_(mul[23]), .PRODUCT_22_(mul[22]), 
        .PRODUCT_21_(mul[21]), .PRODUCT_20_(mul[20]), .PRODUCT_19_(mul[19]), 
        .PRODUCT_18_(mul[18]), .PRODUCT_17_(mul[17]), .PRODUCT_16_(mul[16]), 
        .PRODUCT_15_(mul[15]), .PRODUCT_14_(mul[14]), .PRODUCT_13_(mul[13]), 
        .PRODUCT_12_(mul[12]), .PRODUCT_11_(mul[11]), .PRODUCT_10_(mul[10]), 
        .PRODUCT_9_(mul[9]), .PRODUCT_8_(mul[8]), .PRODUCT_7_(out[0]) );
  XOR2X2 U2 ( .A(mul[18]), .B(n102), .Y(out[11]) );
  INVX4 U3 ( .A(n25), .Y(n23) );
  XOR2X2 U4 ( .A(n34), .B(n33), .Y(in_8bit_b[1]) );
  OAI21X2 U5 ( .A0(mul[18]), .A1(n103), .B0(n106), .Y(n104) );
  NOR3X2 U6 ( .A(n41), .B(n28), .C(in_8bit[2]), .Y(n42) );
  NAND2BX4 U7 ( .AN(mul[17]), .B(n18), .Y(n103) );
  NAND2XL U8 ( .A(in_17bit[2]), .B(n2), .Y(n3) );
  NAND2XL U9 ( .A(n1), .B(n50), .Y(n4) );
  NAND2X2 U10 ( .A(n3), .B(n4), .Y(in_17bit_b[2]) );
  INVXL U11 ( .A(in_17bit[2]), .Y(n1) );
  INVX1 U12 ( .A(n50), .Y(n2) );
  NOR2X4 U13 ( .A(n14), .B(n105), .Y(n102) );
  INVX4 U14 ( .A(n103), .Y(n105) );
  NOR2X1 U15 ( .A(n32), .B(n52), .Y(n15) );
  OAI21X4 U16 ( .A0(in_8bit[2]), .A1(n37), .B0(n23), .Y(n38) );
  NOR2X2 U17 ( .A(n14), .B(n20), .Y(n100) );
  NOR2X1 U18 ( .A(n14), .B(n18), .Y(n101) );
  XOR2X1 U19 ( .A(n59), .B(n57), .Y(in_17bit_b[5]) );
  NAND2BX1 U20 ( .AN(in_8bit[1]), .B(n27), .Y(n44) );
  NAND2BX2 U21 ( .AN(n26), .B(n39), .Y(n41) );
  INVX1 U22 ( .A(n44), .Y(n39) );
  NOR2X1 U23 ( .A(mul[13]), .B(n93), .Y(n13) );
  NOR2X2 U24 ( .A(mul[15]), .B(n97), .Y(n20) );
  NOR2X2 U25 ( .A(mul[16]), .B(n19), .Y(n18) );
  INVX1 U26 ( .A(n20), .Y(n19) );
  INVX1 U27 ( .A(n53), .Y(n56) );
  XOR2X1 U28 ( .A(mul[14]), .B(n96), .Y(out[7]) );
  NOR2X1 U29 ( .A(n14), .B(n13), .Y(n96) );
  XNOR2X1 U30 ( .A(n54), .B(n55), .Y(in_17bit_b[4]) );
  NOR2X1 U31 ( .A(n31), .B(n56), .Y(n54) );
  INVX1 U32 ( .A(in_8bit[3]), .Y(n27) );
  INVX1 U33 ( .A(in_8bit[4]), .Y(n29) );
  INVX1 U34 ( .A(mul[21]), .Y(n12) );
  CLKINVX3 U35 ( .A(n8), .Y(n10) );
  INVXL U36 ( .A(in_17bit[16]), .Y(n32) );
  XNOR2X1 U37 ( .A(n116), .B(sub_add_52_b0_carry[13]), .Y(n5) );
  XNOR2X1 U38 ( .A(n118), .B(sub_add_52_b0_carry[15]), .Y(n6) );
  XNOR2X1 U39 ( .A(n117), .B(sub_add_52_b0_carry[14]), .Y(n7) );
  INVX1 U40 ( .A(n93), .Y(n95) );
  NAND2BX1 U41 ( .AN(mul[12]), .B(n92), .Y(n93) );
  OR3X2 U42 ( .A(in_8bit[6]), .B(n48), .C(n24), .Y(n8) );
  NAND2BX2 U43 ( .AN(mul[18]), .B(n105), .Y(n108) );
  INVX1 U44 ( .A(n97), .Y(n99) );
  NAND2BX1 U45 ( .AN(mul[14]), .B(n13), .Y(n97) );
  OR2X4 U46 ( .A(n108), .B(mul[19]), .Y(n9) );
  AOI21X1 U47 ( .A0(n16), .A1(n111), .B0(n14), .Y(n112) );
  NOR3X2 U48 ( .A(in_8bit[2]), .B(n26), .C(n44), .Y(n46) );
  NOR2X2 U49 ( .A(n14), .B(n17), .Y(n109) );
  INVX3 U50 ( .A(mul[22]), .Y(n111) );
  NOR2X4 U51 ( .A(n9), .B(mul[20]), .Y(n17) );
  OAI22X1 U52 ( .A0(in_17bit[0]), .A1(in_17bit[1]), .B0(in_17bit[16]), .B1(
        in_17bit[1]), .Y(n49) );
  BUFX8 U53 ( .A(in_8bit[0]), .Y(n26) );
  NAND2X2 U54 ( .A(n23), .B(n37), .Y(n35) );
  XOR2X4 U55 ( .A(n43), .B(in_8bit[5]), .Y(in_8bit_b[5]) );
  NOR2X2 U56 ( .A(n42), .B(n24), .Y(n43) );
  XOR2X2 U57 ( .A(n36), .B(n35), .Y(in_8bit_b[2]) );
  XOR2X4 U58 ( .A(n40), .B(n29), .Y(in_8bit_b[4]) );
  OAI21X2 U59 ( .A0(in_8bit[2]), .A1(n41), .B0(n23), .Y(n40) );
  NAND2X1 U60 ( .A(n46), .B(n45), .Y(n48) );
  XOR2X2 U61 ( .A(mul[17]), .B(n101), .Y(out[10]) );
  NAND2BX4 U62 ( .AN(n26), .B(n34), .Y(n37) );
  XOR2X2 U63 ( .A(n27), .B(n38), .Y(in_8bit_b[3]) );
  AND2X4 U64 ( .A(n12), .B(n17), .Y(n16) );
  XOR2X2 U65 ( .A(mul[21]), .B(n109), .Y(out[14]) );
  XNOR2X4 U66 ( .A(mul[20]), .B(n107), .Y(out[13]) );
  BUFX3 U67 ( .A(n104), .Y(n11) );
  INVXL U68 ( .A(in_8bit[2]), .Y(n36) );
  NOR2X1 U69 ( .A(in_8bit[5]), .B(n28), .Y(n45) );
  INVX1 U70 ( .A(n29), .Y(n28) );
  NOR2X2 U71 ( .A(n32), .B(n22), .Y(n50) );
  NOR2X2 U72 ( .A(in_17bit[1]), .B(in_17bit[0]), .Y(n22) );
  XNOR2X1 U73 ( .A(in_17bit[16]), .B(n23), .Y(n14) );
  AND3X1 U74 ( .A(in_17bit[16]), .B(in_17bit[0]), .C(in_17bit[1]), .Y(n21) );
  NOR2X1 U75 ( .A(n14), .B(n86), .Y(n85) );
  MX2XL U76 ( .A(mul[8]), .B(N33), .S0(n106), .Y(out[1]) );
  INVXL U77 ( .A(in_8bit[7]), .Y(n25) );
  INVXL U78 ( .A(in_8bit[7]), .Y(n24) );
  NAND2XL U79 ( .A(n56), .B(n55), .Y(n58) );
  NAND2BXL U80 ( .AN(n58), .B(n59), .Y(n60) );
  NOR2XL U81 ( .A(n31), .B(n70), .Y(n68) );
  NAND2XL U82 ( .A(n63), .B(n62), .Y(n65) );
  NAND2BXL U83 ( .AN(n65), .B(n66), .Y(n67) );
  NOR2XL U84 ( .A(n31), .B(n77), .Y(n75) );
  NAND2XL U85 ( .A(n77), .B(n76), .Y(n79) );
  NAND2XL U86 ( .A(n70), .B(n69), .Y(n72) );
  NAND2BXL U87 ( .AN(n72), .B(n73), .Y(n74) );
  NOR2X2 U88 ( .A(n21), .B(n49), .Y(in_17bit_b[1]) );
  INVXL U89 ( .A(in_17bit[4]), .Y(n55) );
  INVXL U90 ( .A(in_8bit[1]), .Y(n34) );
  NAND2BXL U91 ( .AN(in_17bit[2]), .B(n22), .Y(n51) );
  XOR2X1 U92 ( .A(in_17bit[3]), .B(n15), .Y(in_17bit_b[3]) );
  NAND2BXL U93 ( .AN(in_17bit[3]), .B(n52), .Y(n53) );
  INVXL U94 ( .A(in_17bit[5]), .Y(n59) );
  INVXL U95 ( .A(in_17bit[6]), .Y(n62) );
  INVXL U96 ( .A(in_17bit[8]), .Y(n69) );
  INVXL U97 ( .A(in_17bit[7]), .Y(n66) );
  INVXL U98 ( .A(in_17bit[9]), .Y(n73) );
  INVX1 U99 ( .A(n87), .Y(n89) );
  NAND2BX1 U100 ( .AN(mul[10]), .B(n86), .Y(n87) );
  INVX1 U101 ( .A(n81), .Y(n83) );
  NAND2BX1 U102 ( .AN(mul[8]), .B(n113), .Y(n81) );
  INVX1 U103 ( .A(n84), .Y(n86) );
  NAND2BX1 U104 ( .AN(mul[9]), .B(n83), .Y(n84) );
  INVX1 U105 ( .A(out[0]), .Y(n113) );
  XNOR2X1 U106 ( .A(mul[8]), .B(n113), .Y(N33) );
  XOR2X1 U107 ( .A(mul[23]), .B(n112), .Y(out[16]) );
  INVX1 U108 ( .A(n90), .Y(n92) );
  NAND2BX1 U109 ( .AN(mul[11]), .B(n89), .Y(n90) );
  XOR2X1 U110 ( .A(mul[15]), .B(n98), .Y(out[8]) );
  NOR2XL U111 ( .A(n14), .B(n99), .Y(n98) );
  XOR2X1 U112 ( .A(mul[9]), .B(n82), .Y(out[2]) );
  NOR2X1 U113 ( .A(n14), .B(n83), .Y(n82) );
  XOR2X1 U114 ( .A(mul[11]), .B(n88), .Y(out[4]) );
  NOR2X1 U115 ( .A(n14), .B(n89), .Y(n88) );
  XOR2X1 U116 ( .A(mul[12]), .B(n91), .Y(out[5]) );
  NOR2X1 U117 ( .A(n14), .B(n92), .Y(n91) );
  XOR2X1 U118 ( .A(mul[13]), .B(n94), .Y(out[6]) );
  NOR2X1 U119 ( .A(n14), .B(n95), .Y(n94) );
  XOR2X1 U120 ( .A(mul[10]), .B(n85), .Y(out[3]) );
  INVX1 U121 ( .A(n14), .Y(n106) );
  NAND2XL U122 ( .A(n26), .B(n23), .Y(n33) );
  NOR2X1 U123 ( .A(n79), .B(in_17bit[11]), .Y(sub_add_52_b0_carry[12]) );
  XNOR2X1 U124 ( .A(n61), .B(n62), .Y(in_17bit_b[6]) );
  NOR2X1 U125 ( .A(n31), .B(n63), .Y(n61) );
  XNOR2X1 U126 ( .A(n68), .B(n69), .Y(in_17bit_b[8]) );
  XOR2X1 U127 ( .A(n66), .B(n64), .Y(in_17bit_b[7]) );
  XOR2X1 U128 ( .A(n73), .B(n71), .Y(in_17bit_b[9]) );
  INVX1 U129 ( .A(n60), .Y(n63) );
  INVX1 U130 ( .A(n67), .Y(n70) );
  INVX1 U131 ( .A(n74), .Y(n77) );
  INVXL U132 ( .A(in_8bit[6]), .Y(n30) );
  NAND2X2 U133 ( .A(n48), .B(n23), .Y(n47) );
  XNOR2X1 U134 ( .A(n75), .B(n76), .Y(in_17bit_b[10]) );
  XOR2X1 U135 ( .A(n79), .B(n114), .Y(n78) );
  XNOR2X1 U136 ( .A(n115), .B(sub_add_52_b0_carry[12]), .Y(n80) );
  INVX1 U137 ( .A(n51), .Y(n52) );
  INVX1 U138 ( .A(in_17bit[10]), .Y(n76) );
  INVX1 U139 ( .A(in_17bit[11]), .Y(n114) );
  INVXL U140 ( .A(in_17bit[16]), .Y(n31) );
  INVX1 U141 ( .A(in_17bit[12]), .Y(n115) );
  INVX1 U142 ( .A(in_17bit[13]), .Y(n116) );
  INVX1 U143 ( .A(in_17bit[14]), .Y(n117) );
  INVX1 U144 ( .A(in_17bit[15]), .Y(n118) );
  AND2X1 U145 ( .A(N21), .B(in_17bit[16]), .Y(in_17bit_b[16]) );
  MXI2XL U146 ( .A(n118), .B(n6), .S0(in_17bit[16]), .Y(in_17bit_b[15]) );
  MXI2XL U147 ( .A(n117), .B(n7), .S0(in_17bit[16]), .Y(in_17bit_b[14]) );
  MXI2XL U148 ( .A(n116), .B(n5), .S0(in_17bit[16]), .Y(in_17bit_b[13]) );
  MXI2XL U149 ( .A(n115), .B(n80), .S0(in_17bit[16]), .Y(in_17bit_b[12]) );
  MXI2XL U150 ( .A(n114), .B(n78), .S0(in_17bit[16]), .Y(in_17bit_b[11]) );
  NAND2XL U151 ( .A(n72), .B(in_17bit[16]), .Y(n71) );
  NAND2XL U152 ( .A(n65), .B(in_17bit[16]), .Y(n64) );
  NAND2XL U153 ( .A(n58), .B(in_17bit[16]), .Y(n57) );
  XOR2X4 U154 ( .A(n47), .B(n30), .Y(in_8bit_b[6]) );
  XOR2X4 U155 ( .A(mul[16]), .B(n100), .Y(out[9]) );
  XNOR2X4 U156 ( .A(mul[19]), .B(n11), .Y(out[12]) );
  OAI21X4 U157 ( .A0(mul[19]), .A1(n108), .B0(n106), .Y(n107) );
  NOR2X4 U158 ( .A(n14), .B(n16), .Y(n110) );
  XNOR2X4 U159 ( .A(n110), .B(n111), .Y(out[15]) );
  XOR2X1 U160 ( .A(n31), .B(sub_add_52_b0_carry[16]), .Y(N21) );
  AND2X1 U161 ( .A(sub_add_52_b0_carry[15]), .B(n118), .Y(
        sub_add_52_b0_carry[16]) );
  AND2X1 U162 ( .A(sub_add_52_b0_carry[14]), .B(n117), .Y(
        sub_add_52_b0_carry[15]) );
  AND2X1 U163 ( .A(sub_add_52_b0_carry[13]), .B(n116), .Y(
        sub_add_52_b0_carry[14]) );
  AND2X1 U164 ( .A(sub_add_52_b0_carry[12]), .B(n115), .Y(
        sub_add_52_b0_carry[13]) );
endmodule


module multi16_3_DW01_add_0 ( A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, 
        A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, 
        B_20_, B_19_, B_18_, B_17_, B_16_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, 
        SUM_17_, SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, 
        SUM_9_, SUM_8_, SUM_7_, SUM_6_, SUM_5_ );
  input A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_,
         A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, B_20_, B_19_,
         B_18_, B_17_, B_16_;
  output SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, SUM_15_,
         SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, SUM_7_,
         SUM_6_, SUM_5_;
  wire   n1, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39;

  INVX4 U2 ( .A(n29), .Y(n17) );
  OAI21X2 U3 ( .A0(n26), .A1(n27), .B0(n28), .Y(n22) );
  INVX4 U4 ( .A(n34), .Y(n16) );
  INVX2 U5 ( .A(n19), .Y(SUM_15_) );
  OAI21X2 U6 ( .A0(n37), .A1(n30), .B0(n32), .Y(n35) );
  NOR2X2 U7 ( .A(B_18_), .B(A_18_), .Y(n30) );
  INVX2 U8 ( .A(n30), .Y(n14) );
  BUFX3 U9 ( .A(A_14_), .Y(SUM_14_) );
  INVXL U10 ( .A(n32), .Y(n15) );
  INVX1 U11 ( .A(A_15_), .Y(n19) );
  NAND2X1 U12 ( .A(n24), .B(n23), .Y(n25) );
  XOR2X2 U13 ( .A(n35), .B(n36), .Y(SUM_19_) );
  CLKINVX4 U14 ( .A(n33), .Y(n18) );
  NAND2X2 U15 ( .A(B_16_), .B(A_16_), .Y(n33) );
  AND2X4 U16 ( .A(n33), .B(n1), .Y(SUM_16_) );
  NOR2BX2 U17 ( .AN(n28), .B(n27), .Y(n36) );
  NOR2X1 U18 ( .A(B_19_), .B(A_19_), .Y(n27) );
  XOR2X4 U19 ( .A(n38), .B(n37), .Y(SUM_18_) );
  OR2X2 U20 ( .A(B_16_), .B(A_16_), .Y(n1) );
  OR2X4 U21 ( .A(B_20_), .B(A_20_), .Y(n23) );
  NAND2X2 U22 ( .A(n32), .B(n14), .Y(n38) );
  NOR2X4 U23 ( .A(B_17_), .B(A_17_), .Y(n29) );
  NAND2X1 U24 ( .A(B_18_), .B(A_18_), .Y(n32) );
  NAND2X2 U25 ( .A(B_17_), .B(A_17_), .Y(n34) );
  NOR2X4 U26 ( .A(n29), .B(n16), .Y(n39) );
  XOR2X4 U27 ( .A(n18), .B(n39), .Y(SUM_17_) );
  INVXL U28 ( .A(n24), .Y(n13) );
  BUFX4 U29 ( .A(A_13_), .Y(SUM_13_) );
  BUFX3 U30 ( .A(A_5_), .Y(SUM_5_) );
  BUFX3 U31 ( .A(A_6_), .Y(SUM_6_) );
  BUFX3 U32 ( .A(A_7_), .Y(SUM_7_) );
  BUFX3 U33 ( .A(A_8_), .Y(SUM_8_) );
  BUFX3 U34 ( .A(A_10_), .Y(SUM_10_) );
  BUFX3 U35 ( .A(A_12_), .Y(SUM_12_) );
  BUFX3 U36 ( .A(A_11_), .Y(SUM_11_) );
  BUFX3 U37 ( .A(A_9_), .Y(SUM_9_) );
  AOI21X4 U38 ( .A0(n18), .A1(n17), .B0(n16), .Y(n37) );
  XOR2X1 U39 ( .A(n20), .B(n21), .Y(SUM_21_) );
  AOI21X1 U40 ( .A0(n22), .A1(n23), .B0(n13), .Y(n21) );
  XNOR2X1 U41 ( .A(B_21_), .B(A_21_), .Y(n20) );
  XNOR2X1 U42 ( .A(n25), .B(n22), .Y(SUM_20_) );
  AOI21X1 U43 ( .A0(n14), .A1(n31), .B0(n15), .Y(n26) );
  OAI21XL U44 ( .A0(n29), .A1(n33), .B0(n34), .Y(n31) );
  NAND2X1 U45 ( .A(B_20_), .B(A_20_), .Y(n24) );
  NAND2X1 U46 ( .A(B_19_), .B(A_19_), .Y(n28) );
endmodule


module multi16_3_DW02_mult_0 ( A, B, PRODUCT_23_, PRODUCT_22_, PRODUCT_21_, 
        PRODUCT_20_, PRODUCT_19_, PRODUCT_18_, PRODUCT_17_, PRODUCT_16_, 
        PRODUCT_15_, PRODUCT_14_, PRODUCT_13_, PRODUCT_12_, PRODUCT_11_, 
        PRODUCT_10_, PRODUCT_9_, PRODUCT_8_, PRODUCT_7_ );
  input [16:0] A;
  input [7:0] B;
  output PRODUCT_23_, PRODUCT_22_, PRODUCT_21_, PRODUCT_20_, PRODUCT_19_,
         PRODUCT_18_, PRODUCT_17_, PRODUCT_16_, PRODUCT_15_, PRODUCT_14_,
         PRODUCT_13_, PRODUCT_12_, PRODUCT_11_, PRODUCT_10_, PRODUCT_9_,
         PRODUCT_8_, PRODUCT_7_;
  wire   ab_16__7_, ab_16__6_, ab_16__5_, ab_16__4_, ab_16__3_, ab_16__2_,
         ab_16__1_, ab_16__0_, ab_15__7_, ab_15__6_, ab_15__5_, ab_15__4_,
         ab_15__3_, ab_15__2_, ab_15__1_, ab_15__0_, ab_14__7_, ab_14__6_,
         ab_14__5_, ab_14__4_, ab_14__3_, ab_14__2_, ab_14__1_, ab_14__0_,
         ab_13__7_, ab_13__6_, ab_13__5_, ab_13__4_, ab_13__3_, ab_13__2_,
         ab_13__1_, ab_13__0_, ab_12__7_, ab_12__6_, ab_12__5_, ab_12__4_,
         ab_12__3_, ab_12__2_, ab_12__1_, ab_12__0_, ab_11__7_, ab_11__6_,
         ab_11__5_, ab_11__4_, ab_11__3_, ab_11__2_, ab_11__1_, ab_11__0_,
         ab_10__7_, ab_10__6_, ab_10__5_, ab_10__4_, ab_10__3_, ab_10__2_,
         ab_10__1_, ab_10__0_, ab_9__7_, ab_9__6_, ab_9__5_, ab_9__4_,
         ab_9__3_, ab_9__2_, ab_9__1_, ab_9__0_, ab_8__7_, ab_8__6_, ab_8__5_,
         ab_8__4_, ab_8__3_, ab_8__2_, ab_8__1_, ab_8__0_, ab_7__7_, ab_7__6_,
         ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_, ab_7__0_, ab_6__7_,
         ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_, ab_6__1_, ab_6__0_,
         ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_, ab_5__2_, ab_5__1_,
         ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_, ab_4__3_, ab_4__2_,
         ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_, ab_3__4_, ab_3__3_,
         ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_, ab_2__5_, ab_2__4_,
         ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_, ab_1__6_, ab_1__5_,
         ab_1__4_, ab_1__3_, ab_1__2_, ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_,
         ab_0__3_, ab_0__2_, CARRYB_16__6_, CARRYB_16__5_, CARRYB_16__4_,
         CARRYB_16__3_, CARRYB_16__2_, CARRYB_16__1_, CARRYB_16__0_,
         CARRYB_15__6_, CARRYB_15__5_, CARRYB_15__4_, CARRYB_15__3_,
         CARRYB_15__2_, CARRYB_15__1_, CARRYB_15__0_, CARRYB_14__6_,
         CARRYB_14__5_, CARRYB_14__4_, CARRYB_14__3_, CARRYB_14__2_,
         CARRYB_14__1_, CARRYB_14__0_, CARRYB_13__6_, CARRYB_13__5_,
         CARRYB_13__4_, CARRYB_13__3_, CARRYB_13__2_, CARRYB_13__1_,
         CARRYB_13__0_, CARRYB_12__6_, CARRYB_12__5_, CARRYB_12__4_,
         CARRYB_12__3_, CARRYB_12__2_, CARRYB_12__1_, CARRYB_12__0_,
         CARRYB_11__6_, CARRYB_11__5_, CARRYB_11__4_, CARRYB_11__3_,
         CARRYB_11__2_, CARRYB_11__1_, CARRYB_11__0_, CARRYB_10__6_,
         CARRYB_10__5_, CARRYB_10__4_, CARRYB_10__3_, CARRYB_10__2_,
         CARRYB_10__1_, CARRYB_10__0_, CARRYB_9__6_, CARRYB_9__5_,
         CARRYB_9__4_, CARRYB_9__3_, CARRYB_9__2_, CARRYB_9__1_, CARRYB_9__0_,
         CARRYB_8__6_, CARRYB_8__5_, CARRYB_8__4_, CARRYB_8__3_, CARRYB_8__2_,
         CARRYB_8__1_, CARRYB_8__0_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_,
         CARRYB_7__3_, CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_,
         CARRYB_6__5_, CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_,
         CARRYB_6__0_, CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_,
         CARRYB_5__2_, CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_,
         CARRYB_4__4_, CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_,
         CARRYB_3__6_, CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_,
         CARRYB_3__1_, CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_,
         CARRYB_2__3_, CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__0_,
         SUMB_16__6_, SUMB_16__5_, SUMB_16__4_, SUMB_16__3_, SUMB_16__2_,
         SUMB_16__1_, SUMB_16__0_, SUMB_15__6_, SUMB_15__5_, SUMB_15__4_,
         SUMB_15__3_, SUMB_15__2_, SUMB_15__1_, SUMB_14__6_, SUMB_14__5_,
         SUMB_14__4_, SUMB_14__3_, SUMB_14__2_, SUMB_14__1_, SUMB_13__6_,
         SUMB_13__5_, SUMB_13__4_, SUMB_13__3_, SUMB_13__2_, SUMB_13__1_,
         SUMB_12__6_, SUMB_12__5_, SUMB_12__4_, SUMB_12__3_, SUMB_12__2_,
         SUMB_12__1_, SUMB_11__6_, SUMB_11__5_, SUMB_11__4_, SUMB_11__3_,
         SUMB_11__2_, SUMB_11__1_, SUMB_10__6_, SUMB_10__5_, SUMB_10__4_,
         SUMB_10__3_, SUMB_10__2_, SUMB_10__1_, SUMB_9__6_, SUMB_9__5_,
         SUMB_9__4_, SUMB_9__3_, SUMB_9__2_, SUMB_9__1_, SUMB_8__6_,
         SUMB_8__5_, SUMB_8__4_, SUMB_8__3_, SUMB_8__2_, SUMB_8__1_,
         SUMB_7__6_, SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_,
         SUMB_7__1_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, PROD1_7_, A1_21_, A1_20_, A1_19_, A1_18_,
         A1_17_, A1_16_, A1_15_, A1_13_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_,
         A1_7_, A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61;

  ADDFHX4 S1_14_0 ( .A(ab_14__0_), .B(CARRYB_13__0_), .CI(SUMB_13__1_), .CO(
        CARRYB_14__0_), .S(A1_12_) );
  ADDFHX4 S2_14_1 ( .A(ab_14__1_), .B(CARRYB_13__1_), .CI(SUMB_13__2_), .CO(
        CARRYB_14__1_), .S(SUMB_14__1_) );
  ADDFHX4 S2_14_2 ( .A(ab_14__2_), .B(CARRYB_13__2_), .CI(SUMB_13__3_), .CO(
        CARRYB_14__2_), .S(SUMB_14__2_) );
  ADDFHX4 S1_13_0 ( .A(ab_13__0_), .B(CARRYB_12__0_), .CI(SUMB_12__1_), .CO(
        CARRYB_13__0_), .S(A1_11_) );
  ADDFHX4 S2_13_1 ( .A(ab_13__1_), .B(CARRYB_12__1_), .CI(SUMB_12__2_), .CO(
        CARRYB_13__1_), .S(SUMB_13__1_) );
  ADDFHX4 S2_12_2 ( .A(ab_12__2_), .B(CARRYB_11__2_), .CI(SUMB_11__3_), .CO(
        CARRYB_12__2_), .S(SUMB_12__2_) );
  ADDFHX4 S2_11_1 ( .A(ab_11__1_), .B(CARRYB_10__1_), .CI(SUMB_10__2_), .CO(
        CARRYB_11__1_), .S(SUMB_11__1_) );
  ADDFHX4 S2_11_2 ( .A(ab_11__2_), .B(CARRYB_10__2_), .CI(SUMB_10__3_), .CO(
        CARRYB_11__2_), .S(SUMB_11__2_) );
  multi16_3_DW01_add_0 FS_1 ( .A_21_(A1_21_), .A_20_(A1_20_), .A_19_(A1_19_), 
        .A_18_(A1_18_), .A_17_(A1_17_), .A_16_(A1_16_), .A_15_(A1_15_), 
        .A_14_(SUMB_16__0_), .A_13_(A1_13_), .A_12_(A1_12_), .A_11_(A1_11_), 
        .A_10_(A1_10_), .A_9_(A1_9_), .A_8_(A1_8_), .A_7_(A1_7_), .A_6_(A1_6_), 
        .A_5_(PROD1_7_), .B_21_(n43), .B_20_(n42), .B_19_(n40), .B_18_(n38), 
        .B_17_(n39), .B_16_(n41), .SUM_21_(PRODUCT_23_), .SUM_20_(PRODUCT_22_), 
        .SUM_19_(PRODUCT_21_), .SUM_18_(PRODUCT_20_), .SUM_17_(PRODUCT_19_), 
        .SUM_16_(PRODUCT_18_), .SUM_15_(PRODUCT_17_), .SUM_14_(PRODUCT_16_), 
        .SUM_13_(PRODUCT_15_), .SUM_12_(PRODUCT_14_), .SUM_11_(PRODUCT_13_), 
        .SUM_10_(PRODUCT_12_), .SUM_9_(PRODUCT_11_), .SUM_8_(PRODUCT_10_), 
        .SUM_7_(PRODUCT_9_), .SUM_6_(PRODUCT_8_), .SUM_5_(PRODUCT_7_) );
  ADDFHX1 S3_13_6 ( .A(ab_13__6_), .B(CARRYB_12__6_), .CI(ab_12__7_), .CO(
        CARRYB_13__6_), .S(SUMB_13__6_) );
  ADDFHX2 S2_11_5 ( .A(ab_11__5_), .B(CARRYB_10__5_), .CI(SUMB_10__6_), .CO(
        CARRYB_11__5_), .S(SUMB_11__5_) );
  ADDFHX2 S2_9_4 ( .A(ab_9__4_), .B(CARRYB_8__4_), .CI(SUMB_8__5_), .CO(
        CARRYB_9__4_), .S(SUMB_9__4_) );
  ADDFHX2 S4_5 ( .A(ab_16__5_), .B(CARRYB_15__5_), .CI(SUMB_15__6_), .CO(
        CARRYB_16__5_), .S(SUMB_16__5_) );
  ADDFHX4 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  ADDFHX4 S2_12_3 ( .A(ab_12__3_), .B(CARRYB_11__3_), .CI(SUMB_11__4_), .CO(
        CARRYB_12__3_), .S(SUMB_12__3_) );
  ADDFHX4 S2_13_3 ( .A(ab_13__3_), .B(CARRYB_12__3_), .CI(SUMB_12__4_), .CO(
        CARRYB_13__3_), .S(SUMB_13__3_) );
  ADDFHX4 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  ADDFHX4 S2_15_3 ( .A(ab_15__3_), .B(CARRYB_14__3_), .CI(SUMB_14__4_), .CO(
        CARRYB_15__3_), .S(SUMB_15__3_) );
  ADDFHX4 S2_8_1 ( .A(ab_8__1_), .B(CARRYB_7__1_), .CI(SUMB_7__2_), .CO(
        CARRYB_8__1_), .S(SUMB_8__1_) );
  ADDFHX2 S2_14_4 ( .A(ab_14__4_), .B(CARRYB_13__4_), .CI(SUMB_13__5_), .CO(
        CARRYB_14__4_), .S(SUMB_14__4_) );
  ADDFHX2 S3_10_6 ( .A(ab_10__6_), .B(CARRYB_9__6_), .CI(ab_9__7_), .CO(
        CARRYB_10__6_), .S(SUMB_10__6_) );
  ADDFHX4 S2_8_2 ( .A(ab_8__2_), .B(CARRYB_7__2_), .CI(SUMB_7__3_), .CO(
        CARRYB_8__2_), .S(SUMB_8__2_) );
  ADDFHX4 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  ADDFHX4 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  ADDFHX4 S2_7_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  ADDFHX2 S4_2 ( .A(ab_16__2_), .B(CARRYB_15__2_), .CI(SUMB_15__3_), .CO(
        CARRYB_16__2_), .S(SUMB_16__2_) );
  ADDFHX4 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  ADDFHX4 S4_3 ( .A(ab_16__3_), .B(CARRYB_15__3_), .CI(SUMB_15__4_), .CO(
        CARRYB_16__3_), .S(SUMB_16__3_) );
  ADDFHX4 S1_11_0 ( .A(ab_11__0_), .B(CARRYB_10__0_), .CI(SUMB_10__1_), .CO(
        CARRYB_11__0_), .S(A1_9_) );
  ADDFHX4 S1_8_0 ( .A(ab_8__0_), .B(CARRYB_7__0_), .CI(SUMB_7__1_), .CO(
        CARRYB_8__0_), .S(A1_6_) );
  ADDFHX4 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  ADDFHX4 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  ADDFHX4 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  ADDFHX2 S2_14_5 ( .A(ab_14__5_), .B(CARRYB_13__5_), .CI(SUMB_13__6_), .CO(
        CARRYB_14__5_), .S(SUMB_14__5_) );
  ADDFHX2 S2_15_4 ( .A(ab_15__4_), .B(CARRYB_14__4_), .CI(SUMB_14__5_), .CO(
        CARRYB_15__4_), .S(SUMB_15__4_) );
  ADDFHX4 S2_11_4 ( .A(ab_11__4_), .B(CARRYB_10__4_), .CI(SUMB_10__5_), .CO(
        CARRYB_11__4_), .S(SUMB_11__4_) );
  ADDFHX4 S2_12_4 ( .A(ab_12__4_), .B(CARRYB_11__4_), .CI(SUMB_11__5_), .CO(
        CARRYB_12__4_), .S(SUMB_12__4_) );
  ADDFHX4 S2_7_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  ADDFHX4 S2_8_3 ( .A(ab_8__3_), .B(CARRYB_7__3_), .CI(SUMB_7__4_), .CO(
        CARRYB_8__3_), .S(SUMB_8__3_) );
  ADDFHX4 S3_7_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(
        CARRYB_7__6_), .S(SUMB_7__6_) );
  ADDFHX2 S3_15_6 ( .A(ab_15__6_), .B(CARRYB_14__6_), .CI(ab_14__7_), .CO(
        CARRYB_15__6_), .S(SUMB_15__6_) );
  ADDFHX4 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  ADDFHX4 S2_7_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  ADDFHX4 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  ADDFHX4 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  ADDFHX4 S1_10_0 ( .A(ab_10__0_), .B(CARRYB_9__0_), .CI(SUMB_9__1_), .CO(
        CARRYB_10__0_), .S(A1_8_) );
  ADDFHX4 S2_12_5 ( .A(ab_12__5_), .B(CARRYB_11__5_), .CI(SUMB_11__6_), .CO(
        CARRYB_12__5_), .S(SUMB_12__5_) );
  ADDFHX2 S2_13_5 ( .A(ab_13__5_), .B(CARRYB_12__5_), .CI(SUMB_12__6_), .CO(
        CARRYB_13__5_), .S(SUMB_13__5_) );
  ADDFHX2 S3_12_6 ( .A(ab_12__6_), .B(CARRYB_11__6_), .CI(ab_11__7_), .CO(
        CARRYB_12__6_), .S(SUMB_12__6_) );
  ADDFHX4 S2_11_3 ( .A(ab_11__3_), .B(CARRYB_10__3_), .CI(SUMB_10__4_), .CO(
        CARRYB_11__3_), .S(SUMB_11__3_) );
  ADDFHX4 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  ADDFHX4 S2_10_3 ( .A(ab_10__3_), .B(CARRYB_9__3_), .CI(SUMB_9__4_), .CO(
        CARRYB_10__3_), .S(SUMB_10__3_) );
  ADDFHX4 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  ADDFHX4 S2_14_3 ( .A(ab_14__3_), .B(CARRYB_13__3_), .CI(SUMB_13__4_), .CO(
        CARRYB_14__3_), .S(SUMB_14__3_) );
  ADDFHX4 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  ADDFHX4 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  ADDFHX4 S2_10_1 ( .A(ab_10__1_), .B(CARRYB_9__1_), .CI(SUMB_9__2_), .CO(
        CARRYB_10__1_), .S(SUMB_10__1_) );
  ADDFHX4 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  ADDFHX4 S2_10_2 ( .A(ab_10__2_), .B(CARRYB_9__2_), .CI(SUMB_9__3_), .CO(
        CARRYB_10__2_), .S(SUMB_10__2_) );
  ADDFX2 S5_6 ( .A(ab_16__6_), .B(CARRYB_15__6_), .CI(ab_15__7_), .CO(
        CARRYB_16__6_), .S(SUMB_16__6_) );
  ADDFHX2 S2_15_5 ( .A(ab_15__5_), .B(CARRYB_14__5_), .CI(SUMB_14__6_), .CO(
        CARRYB_15__5_), .S(SUMB_15__5_) );
  ADDFHX1 S4_1 ( .A(ab_16__1_), .B(CARRYB_15__1_), .CI(SUMB_15__2_), .CO(
        CARRYB_16__1_), .S(SUMB_16__1_) );
  ADDFHX2 S1_9_0 ( .A(ab_9__0_), .B(CARRYB_8__0_), .CI(SUMB_8__1_), .CO(
        CARRYB_9__0_), .S(A1_7_) );
  ADDFHX2 S3_8_6 ( .A(ab_8__6_), .B(CARRYB_7__6_), .CI(ab_7__7_), .CO(
        CARRYB_8__6_), .S(SUMB_8__6_) );
  ADDFHX2 S2_13_4 ( .A(ab_13__4_), .B(CARRYB_12__4_), .CI(SUMB_12__5_), .CO(
        CARRYB_13__4_), .S(SUMB_13__4_) );
  ADDFHX2 S2_9_2 ( .A(ab_9__2_), .B(CARRYB_8__2_), .CI(SUMB_8__3_), .CO(
        CARRYB_9__2_), .S(SUMB_9__2_) );
  ADDFHX2 S2_2_4 ( .A(ab_2__4_), .B(n24), .CI(SUMB_1__5_), .CO(CARRYB_2__4_), 
        .S(SUMB_2__4_) );
  ADDFHX2 S2_2_5 ( .A(ab_2__5_), .B(n29), .CI(SUMB_1__6_), .CO(CARRYB_2__5_), 
        .S(SUMB_2__5_) );
  ADDFHX2 S3_2_6 ( .A(ab_2__6_), .B(n27), .CI(ab_1__7_), .CO(CARRYB_2__6_), 
        .S(SUMB_2__6_) );
  ADDFHX2 S4_4 ( .A(ab_16__4_), .B(CARRYB_15__4_), .CI(SUMB_15__5_), .CO(
        CARRYB_16__4_), .S(SUMB_16__4_) );
  ADDFHX2 S3_9_6 ( .A(ab_9__6_), .B(CARRYB_8__6_), .CI(ab_8__7_), .CO(
        CARRYB_9__6_), .S(SUMB_9__6_) );
  ADDFHX2 S2_15_1 ( .A(ab_15__1_), .B(CARRYB_14__1_), .CI(SUMB_14__2_), .CO(
        CARRYB_15__1_), .S(SUMB_15__1_) );
  ADDFHX2 S2_7_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  ADDFHX4 S2_2_1 ( .A(ab_2__1_), .B(n28), .CI(SUMB_1__2_), .CO(CARRYB_2__1_), 
        .S(SUMB_2__1_) );
  ADDFHX2 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  ADDFHX4 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  ADDFHX4 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  ADDFHX4 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  ADDFHX4 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  ADDFHX4 S2_2_2 ( .A(ab_2__2_), .B(n26), .CI(SUMB_1__3_), .CO(CARRYB_2__2_), 
        .S(SUMB_2__2_) );
  ADDFHX4 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  ADDFHX1 S2_9_5 ( .A(ab_9__5_), .B(CARRYB_8__5_), .CI(SUMB_8__6_), .CO(
        CARRYB_9__5_), .S(SUMB_9__5_) );
  ADDFHX4 S2_7_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  ADDFHX4 S2_9_3 ( .A(ab_9__3_), .B(CARRYB_8__3_), .CI(SUMB_8__4_), .CO(
        CARRYB_9__3_), .S(SUMB_9__3_) );
  ADDFHX4 S2_9_1 ( .A(ab_9__1_), .B(CARRYB_8__1_), .CI(SUMB_8__2_), .CO(
        CARRYB_9__1_), .S(SUMB_9__1_) );
  ADDFHX4 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  ADDFHX4 S1_7_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(PROD1_7_) );
  ADDFHX4 S1_12_0 ( .A(ab_12__0_), .B(CARRYB_11__0_), .CI(SUMB_11__1_), .CO(
        CARRYB_12__0_), .S(A1_10_) );
  ADDFHX4 S1_15_0 ( .A(ab_15__0_), .B(CARRYB_14__0_), .CI(SUMB_14__1_), .CO(
        CARRYB_15__0_), .S(A1_13_) );
  ADDFHX2 S4_0 ( .A(ab_16__0_), .B(CARRYB_15__0_), .CI(SUMB_15__1_), .CO(
        CARRYB_16__0_), .S(SUMB_16__0_) );
  ADDFHX4 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  ADDFHX4 S2_13_2 ( .A(ab_13__2_), .B(CARRYB_12__2_), .CI(SUMB_12__3_), .CO(
        CARRYB_13__2_), .S(SUMB_13__2_) );
  ADDFHX4 S2_15_2 ( .A(ab_15__2_), .B(CARRYB_14__2_), .CI(SUMB_14__3_), .CO(
        CARRYB_15__2_), .S(SUMB_15__2_) );
  ADDFHX4 S3_11_6 ( .A(ab_11__6_), .B(CARRYB_10__6_), .CI(ab_10__7_), .CO(
        CARRYB_11__6_), .S(SUMB_11__6_) );
  ADDFHX1 S3_14_6 ( .A(ab_14__6_), .B(CARRYB_13__6_), .CI(ab_13__7_), .CO(
        CARRYB_14__6_), .S(SUMB_14__6_) );
  ADDFHX2 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  ADDFHX4 S2_2_3 ( .A(ab_2__3_), .B(n25), .CI(SUMB_1__4_), .CO(CARRYB_2__3_), 
        .S(SUMB_2__3_) );
  ADDFHX2 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  AND2X4 U2 ( .A(ab_0__5_), .B(ab_1__4_), .Y(n24) );
  NAND3X2 U3 ( .A(n20), .B(n21), .C(n22), .Y(CARRYB_5__6_) );
  NAND2X2 U4 ( .A(A[1]), .B(B[1]), .Y(n46) );
  NOR2X1 U5 ( .A(n46), .B(n45), .Y(CARRYB_1__0_) );
  INVX2 U6 ( .A(n46), .Y(n54) );
  AND2X4 U7 ( .A(ab_0__4_), .B(ab_1__3_), .Y(n25) );
  XOR3X4 U8 ( .A(CARRYB_7__4_), .B(ab_8__4_), .C(SUMB_7__5_), .Y(SUMB_8__4_)
         );
  NAND2X1 U9 ( .A(SUMB_7__5_), .B(CARRYB_7__4_), .Y(n3) );
  NAND2X1 U10 ( .A(ab_8__4_), .B(CARRYB_7__4_), .Y(n4) );
  NAND2X1 U11 ( .A(ab_8__4_), .B(SUMB_7__5_), .Y(n5) );
  NAND3X2 U12 ( .A(n5), .B(n3), .C(n4), .Y(CARRYB_8__4_) );
  XOR2X4 U13 ( .A(SUMB_7__6_), .B(ab_8__5_), .Y(n6) );
  XOR2X2 U14 ( .A(CARRYB_7__5_), .B(n6), .Y(SUMB_8__5_) );
  NAND2XL U15 ( .A(SUMB_7__6_), .B(CARRYB_7__5_), .Y(n7) );
  NAND2X1 U16 ( .A(ab_8__5_), .B(CARRYB_7__5_), .Y(n8) );
  NAND2XL U17 ( .A(ab_8__5_), .B(SUMB_7__6_), .Y(n9) );
  NAND3X2 U18 ( .A(n9), .B(n7), .C(n8), .Y(CARRYB_8__5_) );
  XOR3X4 U19 ( .A(CARRYB_4__2_), .B(ab_5__2_), .C(SUMB_4__3_), .Y(SUMB_5__2_)
         );
  NAND2X2 U20 ( .A(SUMB_4__3_), .B(CARRYB_4__2_), .Y(n10) );
  NAND2X2 U21 ( .A(ab_5__2_), .B(CARRYB_4__2_), .Y(n11) );
  NAND2X2 U22 ( .A(ab_5__2_), .B(SUMB_4__3_), .Y(n12) );
  NAND3X4 U23 ( .A(n12), .B(n10), .C(n11), .Y(CARRYB_5__2_) );
  AND2X2 U24 ( .A(A[5]), .B(B[2]), .Y(ab_5__2_) );
  XOR3X4 U25 ( .A(CARRYB_11__1_), .B(ab_12__1_), .C(SUMB_11__2_), .Y(
        SUMB_12__1_) );
  NAND2X2 U26 ( .A(SUMB_11__2_), .B(CARRYB_11__1_), .Y(n13) );
  NAND2X2 U27 ( .A(ab_12__1_), .B(CARRYB_11__1_), .Y(n14) );
  NAND2X2 U28 ( .A(ab_12__1_), .B(SUMB_11__2_), .Y(n15) );
  NAND3X4 U29 ( .A(n15), .B(n13), .C(n14), .Y(CARRYB_12__1_) );
  XOR3X2 U30 ( .A(ab_4__6_), .B(CARRYB_3__6_), .C(ab_3__7_), .Y(SUMB_4__6_) );
  NAND2XL U31 ( .A(ab_4__6_), .B(CARRYB_3__6_), .Y(n16) );
  NAND2XL U32 ( .A(ab_4__6_), .B(ab_3__7_), .Y(n17) );
  NAND2X1 U33 ( .A(CARRYB_3__6_), .B(ab_3__7_), .Y(n18) );
  NAND3X2 U34 ( .A(n16), .B(n17), .C(n18), .Y(CARRYB_4__6_) );
  XOR2X1 U35 ( .A(ab_5__6_), .B(ab_4__7_), .Y(n19) );
  XOR2X1 U36 ( .A(n19), .B(CARRYB_4__6_), .Y(SUMB_5__6_) );
  NAND2X1 U37 ( .A(ab_5__6_), .B(ab_4__7_), .Y(n20) );
  NAND2X1 U38 ( .A(ab_5__6_), .B(CARRYB_4__6_), .Y(n21) );
  NAND2X1 U39 ( .A(ab_4__7_), .B(CARRYB_4__6_), .Y(n22) );
  AND2X2 U40 ( .A(A[2]), .B(B[2]), .Y(ab_2__2_) );
  NOR2X4 U41 ( .A(n49), .B(n37), .Y(ab_0__4_) );
  INVX3 U42 ( .A(B[4]), .Y(n49) );
  AND2X2 U43 ( .A(A[1]), .B(B[4]), .Y(ab_1__4_) );
  AND2X2 U44 ( .A(A[1]), .B(B[5]), .Y(ab_1__5_) );
  AND2X2 U45 ( .A(A[1]), .B(B[3]), .Y(ab_1__3_) );
  NOR2X2 U46 ( .A(n47), .B(n37), .Y(ab_0__6_) );
  NOR2X1 U47 ( .A(n51), .B(n37), .Y(ab_0__2_) );
  INVX1 U48 ( .A(B[3]), .Y(n50) );
  INVX1 U49 ( .A(B[2]), .Y(n51) );
  XOR2X1 U50 ( .A(CARRYB_16__4_), .B(SUMB_16__5_), .Y(A1_19_) );
  XOR2X2 U51 ( .A(CARRYB_16__3_), .B(SUMB_16__4_), .Y(A1_18_) );
  XOR2X1 U52 ( .A(CARRYB_16__0_), .B(SUMB_16__1_), .Y(A1_15_) );
  AND2X2 U54 ( .A(ab_0__3_), .B(ab_1__2_), .Y(n26) );
  AND2X4 U55 ( .A(ab_0__7_), .B(ab_1__6_), .Y(n27) );
  AND2X2 U56 ( .A(ab_0__2_), .B(n54), .Y(n28) );
  AND2X2 U57 ( .A(ab_0__6_), .B(ab_1__5_), .Y(n29) );
  AND2X2 U58 ( .A(A[2]), .B(B[6]), .Y(ab_2__6_) );
  AND2X2 U59 ( .A(A[2]), .B(B[3]), .Y(ab_2__3_) );
  XOR2X2 U60 ( .A(CARRYB_16__5_), .B(SUMB_16__6_), .Y(A1_20_) );
  AND2X2 U61 ( .A(A[2]), .B(B[4]), .Y(ab_2__4_) );
  XOR2X4 U62 ( .A(CARRYB_16__2_), .B(SUMB_16__3_), .Y(A1_17_) );
  AND2X2 U63 ( .A(CARRYB_16__1_), .B(SUMB_16__2_), .Y(n39) );
  AND2X2 U64 ( .A(CARRYB_16__0_), .B(SUMB_16__1_), .Y(n41) );
  AND2X2 U65 ( .A(A[2]), .B(B[5]), .Y(ab_2__5_) );
  AND2XL U66 ( .A(A[7]), .B(B[3]), .Y(ab_7__3_) );
  AND2XL U67 ( .A(A[5]), .B(B[3]), .Y(ab_5__3_) );
  AND2XL U68 ( .A(A[4]), .B(B[3]), .Y(ab_4__3_) );
  AND2X2 U69 ( .A(A[3]), .B(B[3]), .Y(ab_3__3_) );
  XOR3X2 U70 ( .A(CARRYB_9__4_), .B(ab_10__4_), .C(SUMB_9__5_), .Y(SUMB_10__4_) );
  NAND2XL U71 ( .A(SUMB_9__5_), .B(CARRYB_9__4_), .Y(n30) );
  NAND2XL U72 ( .A(ab_10__4_), .B(CARRYB_9__4_), .Y(n31) );
  NAND2XL U73 ( .A(ab_10__4_), .B(SUMB_9__5_), .Y(n32) );
  NAND3X2 U74 ( .A(n32), .B(n30), .C(n31), .Y(CARRYB_10__4_) );
  XOR2X4 U75 ( .A(SUMB_9__6_), .B(ab_10__5_), .Y(n33) );
  XOR2X1 U76 ( .A(CARRYB_9__5_), .B(n33), .Y(SUMB_10__5_) );
  NAND2XL U77 ( .A(SUMB_9__6_), .B(CARRYB_9__5_), .Y(n34) );
  NAND2X1 U78 ( .A(ab_10__5_), .B(CARRYB_9__5_), .Y(n35) );
  NAND2XL U79 ( .A(ab_10__5_), .B(SUMB_9__6_), .Y(n36) );
  NAND3X2 U80 ( .A(n36), .B(n34), .C(n35), .Y(CARRYB_10__5_) );
  BUFX4 U81 ( .A(n44), .Y(n37) );
  INVX4 U82 ( .A(B[6]), .Y(n47) );
  INVX2 U83 ( .A(B[7]), .Y(n53) );
  XOR2X1 U84 ( .A(ab_1__5_), .B(ab_0__6_), .Y(SUMB_1__5_) );
  INVX4 U85 ( .A(B[5]), .Y(n48) );
  AND2X1 U86 ( .A(CARRYB_16__2_), .B(SUMB_16__3_), .Y(n38) );
  AND2X1 U87 ( .A(A[10]), .B(B[1]), .Y(ab_10__1_) );
  AND2X1 U88 ( .A(A[8]), .B(B[1]), .Y(ab_8__1_) );
  AND2X1 U89 ( .A(A[8]), .B(B[0]), .Y(ab_8__0_) );
  AND2X1 U90 ( .A(A[5]), .B(B[1]), .Y(ab_5__1_) );
  XOR2X1 U91 ( .A(n54), .B(ab_0__2_), .Y(SUMB_1__1_) );
  INVXL U92 ( .A(B[1]), .Y(n52) );
  NOR2X1 U93 ( .A(n53), .B(n37), .Y(ab_0__7_) );
  NOR2XL U94 ( .A(n60), .B(n52), .Y(ab_11__1_) );
  INVXL U95 ( .A(A[0]), .Y(n44) );
  NAND2XL U96 ( .A(A[0]), .B(B[0]), .Y(n45) );
  XOR2X2 U97 ( .A(CARRYB_16__1_), .B(SUMB_16__2_), .Y(A1_16_) );
  AND2X2 U98 ( .A(CARRYB_16__3_), .B(SUMB_16__4_), .Y(n40) );
  AND2X2 U99 ( .A(CARRYB_16__4_), .B(SUMB_16__5_), .Y(n42) );
  INVX1 U100 ( .A(B[0]), .Y(n61) );
  NOR2X1 U101 ( .A(n55), .B(n48), .Y(ab_16__5_) );
  NOR2XL U102 ( .A(n55), .B(n51), .Y(ab_16__2_) );
  NOR2X1 U103 ( .A(n55), .B(n49), .Y(ab_16__4_) );
  NOR2X1 U104 ( .A(n55), .B(n52), .Y(ab_16__1_) );
  AND2X1 U105 ( .A(A[10]), .B(B[2]), .Y(ab_10__2_) );
  AND2X1 U106 ( .A(A[9]), .B(B[2]), .Y(ab_9__2_) );
  AND2X2 U107 ( .A(A[9]), .B(B[1]), .Y(ab_9__1_) );
  AND2X1 U108 ( .A(A[8]), .B(B[2]), .Y(ab_8__2_) );
  AND2X2 U109 ( .A(A[10]), .B(B[0]), .Y(ab_10__0_) );
  AND2X1 U110 ( .A(A[7]), .B(B[2]), .Y(ab_7__2_) );
  AND2X1 U111 ( .A(A[10]), .B(B[5]), .Y(ab_10__5_) );
  AND2X1 U112 ( .A(A[9]), .B(B[5]), .Y(ab_9__5_) );
  AND2X1 U113 ( .A(A[8]), .B(B[5]), .Y(ab_8__5_) );
  AND2X1 U114 ( .A(A[7]), .B(B[5]), .Y(ab_7__5_) );
  AND2X2 U115 ( .A(A[7]), .B(B[1]), .Y(ab_7__1_) );
  AND2X1 U116 ( .A(A[6]), .B(B[2]), .Y(ab_6__2_) );
  AND2X1 U117 ( .A(A[6]), .B(B[5]), .Y(ab_6__5_) );
  AND2X1 U118 ( .A(A[4]), .B(B[5]), .Y(ab_4__5_) );
  AND2X1 U119 ( .A(A[5]), .B(B[5]), .Y(ab_5__5_) );
  AND2X2 U120 ( .A(A[9]), .B(B[0]), .Y(ab_9__0_) );
  AND2X1 U121 ( .A(A[10]), .B(B[6]), .Y(ab_10__6_) );
  AND2X1 U122 ( .A(A[9]), .B(B[6]), .Y(ab_9__6_) );
  AND2X1 U123 ( .A(A[8]), .B(B[6]), .Y(ab_8__6_) );
  AND2X1 U124 ( .A(A[7]), .B(B[6]), .Y(ab_7__6_) );
  AND2X1 U125 ( .A(A[6]), .B(B[6]), .Y(ab_6__6_) );
  AND2X1 U126 ( .A(A[5]), .B(B[6]), .Y(ab_5__6_) );
  AND2X2 U127 ( .A(A[6]), .B(B[1]), .Y(ab_6__1_) );
  AND2X1 U128 ( .A(A[4]), .B(B[2]), .Y(ab_4__2_) );
  AND2X2 U129 ( .A(A[4]), .B(B[1]), .Y(ab_4__1_) );
  AND2X2 U130 ( .A(A[5]), .B(B[0]), .Y(ab_5__0_) );
  AND2X2 U131 ( .A(A[4]), .B(B[0]), .Y(ab_4__0_) );
  AND2X2 U132 ( .A(A[7]), .B(B[0]), .Y(ab_7__0_) );
  AND2X2 U133 ( .A(A[6]), .B(B[0]), .Y(ab_6__0_) );
  XOR2X1 U134 ( .A(CARRYB_16__6_), .B(ab_16__7_), .Y(A1_21_) );
  AND2X2 U135 ( .A(CARRYB_16__5_), .B(SUMB_16__6_), .Y(n43) );
  NOR2X1 U136 ( .A(n55), .B(n53), .Y(ab_16__7_) );
  NOR2X1 U137 ( .A(n50), .B(n37), .Y(ab_0__3_) );
  NOR2XL U138 ( .A(n56), .B(n53), .Y(ab_15__7_) );
  NOR2XL U139 ( .A(n55), .B(n47), .Y(ab_16__6_) );
  AND2X1 U140 ( .A(A[3]), .B(B[4]), .Y(ab_3__4_) );
  NOR2X1 U141 ( .A(n57), .B(n52), .Y(ab_14__1_) );
  NOR2X1 U142 ( .A(n58), .B(n52), .Y(ab_13__1_) );
  NOR2X1 U143 ( .A(n56), .B(n52), .Y(ab_15__1_) );
  NOR2X1 U144 ( .A(n59), .B(n52), .Y(ab_12__1_) );
  NOR2XL U145 ( .A(n58), .B(n51), .Y(ab_13__2_) );
  NOR2XL U146 ( .A(n59), .B(n51), .Y(ab_12__2_) );
  NOR2XL U147 ( .A(n57), .B(n51), .Y(ab_14__2_) );
  NOR2XL U148 ( .A(n56), .B(n51), .Y(ab_15__2_) );
  NOR2XL U149 ( .A(n60), .B(n51), .Y(ab_11__2_) );
  AND2X1 U150 ( .A(A[10]), .B(B[4]), .Y(ab_10__4_) );
  NOR2XL U151 ( .A(n60), .B(n49), .Y(ab_11__4_) );
  NOR2XL U152 ( .A(n59), .B(n49), .Y(ab_12__4_) );
  NOR2XL U153 ( .A(n58), .B(n49), .Y(ab_13__4_) );
  NOR2XL U154 ( .A(n57), .B(n49), .Y(ab_14__4_) );
  AND2X1 U155 ( .A(A[9]), .B(B[4]), .Y(ab_9__4_) );
  AND2X1 U156 ( .A(A[8]), .B(B[4]), .Y(ab_8__4_) );
  AND2X1 U157 ( .A(A[7]), .B(B[4]), .Y(ab_7__4_) );
  AND2X1 U158 ( .A(A[6]), .B(B[4]), .Y(ab_6__4_) );
  NOR2XL U159 ( .A(n60), .B(n48), .Y(ab_11__5_) );
  NOR2XL U160 ( .A(n59), .B(n48), .Y(ab_12__5_) );
  NOR2XL U161 ( .A(n58), .B(n48), .Y(ab_13__5_) );
  AND2X1 U162 ( .A(A[4]), .B(B[4]), .Y(ab_4__4_) );
  AND2X1 U163 ( .A(A[5]), .B(B[4]), .Y(ab_5__4_) );
  NOR2XL U164 ( .A(n56), .B(n48), .Y(ab_15__5_) );
  AND2X1 U165 ( .A(A[3]), .B(B[5]), .Y(ab_3__5_) );
  NOR2XL U166 ( .A(n60), .B(n53), .Y(ab_11__7_) );
  NOR2XL U167 ( .A(n59), .B(n47), .Y(ab_12__6_) );
  NOR2XL U168 ( .A(n60), .B(n47), .Y(ab_11__6_) );
  AND2X1 U169 ( .A(A[4]), .B(B[6]), .Y(ab_4__6_) );
  AND2X1 U170 ( .A(A[3]), .B(B[6]), .Y(ab_3__6_) );
  AND2X1 U171 ( .A(A[3]), .B(B[2]), .Y(ab_3__2_) );
  AND2X1 U172 ( .A(A[3]), .B(B[1]), .Y(ab_3__1_) );
  NOR2XL U173 ( .A(n58), .B(n53), .Y(ab_13__7_) );
  NOR2XL U174 ( .A(n57), .B(n47), .Y(ab_14__6_) );
  AND2X1 U175 ( .A(A[3]), .B(B[0]), .Y(ab_3__0_) );
  XOR2X1 U176 ( .A(ab_1__6_), .B(ab_0__7_), .Y(SUMB_1__6_) );
  XOR2X1 U177 ( .A(ab_1__3_), .B(ab_0__4_), .Y(SUMB_1__3_) );
  XOR2X1 U178 ( .A(ab_1__2_), .B(ab_0__3_), .Y(SUMB_1__2_) );
  AND2X2 U179 ( .A(A[2]), .B(B[1]), .Y(ab_2__1_) );
  XOR2X1 U180 ( .A(ab_1__4_), .B(ab_0__5_), .Y(SUMB_1__4_) );
  NOR2XL U181 ( .A(n57), .B(n48), .Y(ab_14__5_) );
  NOR2XL U182 ( .A(n57), .B(n53), .Y(ab_14__7_) );
  NOR2XL U183 ( .A(n56), .B(n47), .Y(ab_15__6_) );
  NOR2XL U184 ( .A(n59), .B(n53), .Y(ab_12__7_) );
  NOR2XL U185 ( .A(n58), .B(n47), .Y(ab_13__6_) );
  NOR2XL U186 ( .A(n56), .B(n49), .Y(ab_15__4_) );
  AND2X2 U187 ( .A(A[2]), .B(B[0]), .Y(ab_2__0_) );
  INVX1 U188 ( .A(A[16]), .Y(n55) );
  INVX1 U189 ( .A(A[11]), .Y(n60) );
  INVX1 U190 ( .A(A[12]), .Y(n59) );
  INVX1 U191 ( .A(A[13]), .Y(n58) );
  INVX1 U192 ( .A(A[14]), .Y(n57) );
  INVX1 U193 ( .A(A[15]), .Y(n56) );
  NOR2XL U194 ( .A(n55), .B(n50), .Y(ab_16__3_) );
  NOR2XL U195 ( .A(n56), .B(n50), .Y(ab_15__3_) );
  NOR2XL U196 ( .A(n57), .B(n50), .Y(ab_14__3_) );
  NOR2XL U197 ( .A(n58), .B(n50), .Y(ab_13__3_) );
  NOR2XL U198 ( .A(n59), .B(n50), .Y(ab_12__3_) );
  NOR2XL U199 ( .A(n60), .B(n50), .Y(ab_11__3_) );
  AND2X1 U200 ( .A(A[10]), .B(B[3]), .Y(ab_10__3_) );
  AND2X1 U201 ( .A(A[9]), .B(B[3]), .Y(ab_9__3_) );
  AND2X1 U202 ( .A(A[8]), .B(B[3]), .Y(ab_8__3_) );
  AND2X1 U203 ( .A(A[6]), .B(B[3]), .Y(ab_6__3_) );
  AND2X1 U204 ( .A(A[10]), .B(B[7]), .Y(ab_10__7_) );
  AND2X1 U205 ( .A(A[9]), .B(B[7]), .Y(ab_9__7_) );
  AND2X1 U206 ( .A(A[8]), .B(B[7]), .Y(ab_8__7_) );
  AND2X1 U207 ( .A(A[7]), .B(B[7]), .Y(ab_7__7_) );
  AND2X1 U208 ( .A(A[6]), .B(B[7]), .Y(ab_6__7_) );
  AND2X1 U209 ( .A(A[5]), .B(B[7]), .Y(ab_5__7_) );
  AND2X1 U210 ( .A(A[4]), .B(B[7]), .Y(ab_4__7_) );
  AND2X1 U211 ( .A(A[3]), .B(B[7]), .Y(ab_3__7_) );
  AND2X1 U212 ( .A(A[2]), .B(B[7]), .Y(ab_2__7_) );
  AND2X2 U213 ( .A(A[1]), .B(B[2]), .Y(ab_1__2_) );
  AND2X1 U214 ( .A(A[1]), .B(B[7]), .Y(ab_1__7_) );
  AND2X2 U215 ( .A(A[1]), .B(B[6]), .Y(ab_1__6_) );
  NOR2X4 U216 ( .A(n48), .B(n37), .Y(ab_0__5_) );
  NOR2X1 U218 ( .A(n61), .B(n55), .Y(ab_16__0_) );
  NOR2X1 U219 ( .A(n61), .B(n56), .Y(ab_15__0_) );
  NOR2X1 U220 ( .A(n61), .B(n57), .Y(ab_14__0_) );
  NOR2X1 U221 ( .A(n61), .B(n58), .Y(ab_13__0_) );
  NOR2X1 U222 ( .A(n61), .B(n59), .Y(ab_12__0_) );
  NOR2X1 U223 ( .A(n61), .B(n60), .Y(ab_11__0_) );
endmodule


module multi16_3 ( in_17bit, in_8bit, out );
  input [16:0] in_17bit;
  input [7:0] in_8bit;
  output [16:0] out;
  wire   N18, N19, N20, N21, N32, N33, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n55, n56, n57, n58, n59, n60, n61, n63, n64, n65, n66, n67, n68,
         n69, n71, n72, n73, n74, n75, n76, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n118, n119, n120, n121;
  wire   [16:1] in_17bit_b;
  wire   [7:0] in_8bit_b;
  wire   [23:8] mul;
  wire   [16:12] sub_add_52_b0_carry;

  multi16_3_DW02_mult_0 mult_55 ( .A({in_17bit_b, in_17bit[0]}), .B({
        in_8bit_b[7:5], n2, in_8bit_b[3:0]}), .PRODUCT_23_(mul[23]), 
        .PRODUCT_22_(mul[22]), .PRODUCT_21_(mul[21]), .PRODUCT_20_(mul[20]), 
        .PRODUCT_19_(mul[19]), .PRODUCT_18_(mul[18]), .PRODUCT_17_(mul[17]), 
        .PRODUCT_16_(mul[16]), .PRODUCT_15_(mul[15]), .PRODUCT_14_(mul[14]), 
        .PRODUCT_13_(mul[13]), .PRODUCT_12_(mul[12]), .PRODUCT_11_(mul[11]), 
        .PRODUCT_10_(mul[10]), .PRODUCT_9_(mul[9]), .PRODUCT_8_(mul[8]), 
        .PRODUCT_7_(N32) );
  INVX3 U2 ( .A(mul[22]), .Y(n107) );
  CLKINVX2 U3 ( .A(in_8bit[5]), .Y(n33) );
  XOR2X2 U4 ( .A(n9), .B(n43), .Y(in_17bit_b[4]) );
  NOR2X2 U5 ( .A(in_17bit[1]), .B(in_17bit[0]), .Y(n15) );
  INVX4 U6 ( .A(n97), .Y(n99) );
  OR2X4 U7 ( .A(n23), .B(n15), .Y(n14) );
  CLKINVX2 U8 ( .A(in_17bit[16]), .Y(n23) );
  NAND3X1 U9 ( .A(in_17bit[0]), .B(n21), .C(in_17bit[1]), .Y(n38) );
  OAI21X4 U10 ( .A0(mul[18]), .A1(n97), .B0(n121), .Y(n98) );
  NAND2BX2 U11 ( .AN(mul[17]), .B(n8), .Y(n97) );
  NOR2XL U12 ( .A(in_17bit[1]), .B(in_17bit[0]), .Y(n36) );
  XNOR2X4 U13 ( .A(mul[19]), .B(n98), .Y(out[12]) );
  INVX2 U14 ( .A(in_8bit_b[4]), .Y(n1) );
  CLKINVX4 U15 ( .A(n1), .Y(n2) );
  XNOR2X2 U16 ( .A(in_17bit[2]), .B(n14), .Y(in_17bit_b[2]) );
  XOR2X1 U17 ( .A(n25), .B(n24), .Y(in_8bit_b[1]) );
  NOR2X1 U18 ( .A(n10), .B(n94), .Y(n93) );
  XOR2X2 U19 ( .A(in_17bit[3]), .B(n40), .Y(in_17bit_b[3]) );
  NOR2X2 U20 ( .A(n22), .B(n41), .Y(n40) );
  NOR2XL U21 ( .A(n22), .B(n51), .Y(n49) );
  INVX1 U22 ( .A(n118), .Y(in_8bit_b[0]) );
  XNOR2X2 U23 ( .A(n31), .B(n33), .Y(in_8bit_b[5]) );
  AOI21X1 U24 ( .A0(n30), .A1(n32), .B0(n17), .Y(n31) );
  NOR2X1 U25 ( .A(n10), .B(n88), .Y(n87) );
  CLKINVX3 U26 ( .A(n39), .Y(n41) );
  NAND2X1 U27 ( .A(n6), .B(n7), .Y(in_8bit_b[3]) );
  NAND2X1 U28 ( .A(n4), .B(n5), .Y(n7) );
  XOR2X1 U29 ( .A(n28), .B(n20), .Y(in_8bit_b[4]) );
  OAI21XL U30 ( .A0(in_8bit[3]), .A1(n29), .B0(in_8bit[7]), .Y(n28) );
  INVX1 U31 ( .A(n86), .Y(n88) );
  NAND2BX1 U32 ( .AN(mul[13]), .B(n85), .Y(n86) );
  INVX1 U33 ( .A(n83), .Y(n85) );
  NAND2BX1 U34 ( .AN(mul[12]), .B(n82), .Y(n83) );
  INVX1 U35 ( .A(in_8bit[0]), .Y(n19) );
  NOR2X1 U36 ( .A(mul[16]), .B(n92), .Y(n8) );
  NAND3BX2 U37 ( .AN(in_8bit[1]), .B(n27), .C(n19), .Y(n29) );
  XNOR2X1 U38 ( .A(n103), .B(n102), .Y(out[14]) );
  NOR2X1 U39 ( .A(n10), .B(n104), .Y(n103) );
  NOR3X2 U40 ( .A(mul[20]), .B(mul[19]), .C(n101), .Y(n104) );
  XOR2X1 U41 ( .A(mul[17]), .B(n95), .Y(out[10]) );
  NOR2X1 U42 ( .A(n10), .B(n8), .Y(n95) );
  XNOR2X2 U43 ( .A(mul[20]), .B(n100), .Y(out[13]) );
  CLKINVX4 U44 ( .A(n29), .Y(n32) );
  INVX4 U45 ( .A(n23), .Y(n21) );
  INVXL U46 ( .A(in_17bit[16]), .Y(n22) );
  OR2X2 U47 ( .A(in_8bit[6]), .B(n17), .Y(n3) );
  INVX1 U48 ( .A(n92), .Y(n94) );
  INVXL U49 ( .A(in_8bit[4]), .Y(n20) );
  CLKINVX3 U50 ( .A(n105), .Y(n108) );
  NAND2BXL U51 ( .AN(in_17bit[2]), .B(n15), .Y(n39) );
  NAND2X4 U52 ( .A(n35), .B(in_8bit[7]), .Y(n34) );
  XOR2X4 U53 ( .A(mul[18]), .B(n96), .Y(out[11]) );
  NAND2BX2 U54 ( .AN(mul[21]), .B(n104), .Y(n105) );
  OAI21X4 U55 ( .A0(mul[19]), .A1(n101), .B0(n121), .Y(n100) );
  NAND2BX4 U56 ( .AN(mul[18]), .B(n99), .Y(n101) );
  CLKINVX2 U57 ( .A(in_8bit[2]), .Y(n27) );
  NOR2X1 U58 ( .A(n21), .B(in_17bit[1]), .Y(n37) );
  NAND2XL U59 ( .A(in_8bit[3]), .B(n11), .Y(n6) );
  INVXL U60 ( .A(in_8bit[3]), .Y(n4) );
  CLKINVX1 U61 ( .A(n11), .Y(n5) );
  NAND2X1 U62 ( .A(n29), .B(in_8bit[7]), .Y(n11) );
  INVXL U63 ( .A(in_8bit[1]), .Y(n25) );
  NAND4BX2 U64 ( .AN(in_8bit[3]), .B(n33), .C(n32), .D(n20), .Y(n35) );
  XOR2X2 U65 ( .A(n27), .B(n26), .Y(in_8bit_b[2]) );
  NOR2X2 U66 ( .A(n3), .B(n35), .Y(in_8bit_b[7]) );
  NAND2X1 U67 ( .A(n53), .B(n21), .Y(n52) );
  INVX1 U68 ( .A(mul[21]), .Y(n102) );
  INVXL U69 ( .A(in_17bit[5]), .Y(n47) );
  INVXL U70 ( .A(in_17bit[6]), .Y(n50) );
  INVXL U71 ( .A(in_17bit[7]), .Y(n55) );
  NAND2BXL U72 ( .AN(mul[10]), .B(n75), .Y(n76) );
  INVXL U73 ( .A(n19), .Y(n18) );
  AOI22XL U74 ( .A0(n18), .A1(in_8bit[7]), .B0(n18), .B1(n17), .Y(n118) );
  XOR2X1 U75 ( .A(mul[16]), .B(n93), .Y(out[9]) );
  XOR2X1 U76 ( .A(mul[14]), .B(n87), .Y(out[7]) );
  XOR2X1 U77 ( .A(mul[23]), .B(n109), .Y(out[16]) );
  NOR2XL U78 ( .A(n10), .B(n82), .Y(n81) );
  NOR2XL U79 ( .A(n10), .B(n72), .Y(n71) );
  INVXL U80 ( .A(mul[8]), .Y(n110) );
  AOI22XL U81 ( .A0(mul[8]), .A1(n10), .B0(N33), .B1(n121), .Y(n120) );
  XOR2X1 U82 ( .A(mul[15]), .B(n90), .Y(out[8]) );
  NOR2XL U83 ( .A(n10), .B(n91), .Y(n90) );
  AOI22XL U84 ( .A0(N32), .A1(n10), .B0(N32), .B1(n121), .Y(n119) );
  INVXL U85 ( .A(in_8bit[7]), .Y(n17) );
  OR2X2 U86 ( .A(n22), .B(n44), .Y(n9) );
  INVXL U87 ( .A(in_8bit[6]), .Y(n16) );
  XNOR2X2 U88 ( .A(n49), .B(n50), .Y(in_17bit_b[6]) );
  NOR2XL U89 ( .A(n22), .B(n59), .Y(n57) );
  NAND2XL U90 ( .A(n51), .B(n50), .Y(n53) );
  NAND2BXL U91 ( .AN(n46), .B(n47), .Y(n48) );
  NAND2BXL U92 ( .AN(n53), .B(n55), .Y(n56) );
  NOR2XL U93 ( .A(n22), .B(n67), .Y(n65) );
  NAND2XL U94 ( .A(n61), .B(n21), .Y(n60) );
  NAND2XL U95 ( .A(n67), .B(n66), .Y(n68) );
  NAND2XL U96 ( .A(n59), .B(n58), .Y(n61) );
  NAND2BXL U97 ( .AN(n61), .B(n63), .Y(n64) );
  XNOR2X1 U98 ( .A(n21), .B(in_8bit[7]), .Y(n10) );
  AND2X1 U99 ( .A(N21), .B(n21), .Y(in_17bit_b[16]) );
  INVX1 U100 ( .A(n42), .Y(n44) );
  INVXL U101 ( .A(in_17bit[4]), .Y(n43) );
  MX2X1 U102 ( .A(in_17bit[11]), .B(n12), .S0(n21), .Y(in_17bit_b[11]) );
  XNOR2X1 U103 ( .A(n68), .B(n112), .Y(n12) );
  MX2X1 U104 ( .A(in_17bit[12]), .B(n13), .S0(n21), .Y(in_17bit_b[12]) );
  XOR2X1 U105 ( .A(n113), .B(sub_add_52_b0_carry[12]), .Y(n13) );
  MX2X1 U106 ( .A(in_17bit[13]), .B(N18), .S0(n21), .Y(in_17bit_b[13]) );
  MX2X1 U107 ( .A(in_17bit[14]), .B(N19), .S0(n21), .Y(in_17bit_b[14]) );
  MX2X1 U108 ( .A(in_17bit[15]), .B(N20), .S0(n21), .Y(in_17bit_b[15]) );
  INVXL U109 ( .A(in_17bit[8]), .Y(n58) );
  INVX1 U110 ( .A(n76), .Y(n79) );
  INVX1 U111 ( .A(n73), .Y(n75) );
  NAND2BX1 U112 ( .AN(mul[9]), .B(n72), .Y(n73) );
  INVX1 U113 ( .A(n69), .Y(n72) );
  NAND2BX1 U114 ( .AN(mul[8]), .B(n111), .Y(n69) );
  INVX1 U115 ( .A(N32), .Y(n111) );
  NAND2BX1 U116 ( .AN(mul[15]), .B(n91), .Y(n92) );
  INVX1 U117 ( .A(n89), .Y(n91) );
  NAND2BXL U118 ( .AN(mul[14]), .B(n88), .Y(n89) );
  INVX1 U119 ( .A(n80), .Y(n82) );
  NAND2BX1 U120 ( .AN(mul[11]), .B(n79), .Y(n80) );
  XOR2X1 U121 ( .A(mul[10]), .B(n74), .Y(out[3]) );
  NOR2X1 U122 ( .A(n10), .B(n75), .Y(n74) );
  XOR2X1 U123 ( .A(mul[9]), .B(n71), .Y(out[2]) );
  XOR2X1 U124 ( .A(mul[11]), .B(n78), .Y(out[4]) );
  NOR2X1 U125 ( .A(n10), .B(n79), .Y(n78) );
  XOR2X1 U126 ( .A(mul[12]), .B(n81), .Y(out[5]) );
  XOR2X1 U127 ( .A(mul[13]), .B(n84), .Y(out[6]) );
  NOR2X1 U128 ( .A(n10), .B(n85), .Y(n84) );
  AOI21XL U129 ( .A0(n108), .A1(n107), .B0(n10), .Y(n109) );
  INVX1 U130 ( .A(n120), .Y(out[1]) );
  INVX1 U131 ( .A(n119), .Y(out[0]) );
  INVXL U132 ( .A(n10), .Y(n121) );
  NAND2XL U133 ( .A(n18), .B(in_8bit[7]), .Y(n24) );
  OAI2BB1X1 U134 ( .A0N(n19), .A1N(n25), .B0(in_8bit[7]), .Y(n26) );
  XNOR2X1 U135 ( .A(n57), .B(n58), .Y(in_17bit_b[8]) );
  XNOR2X1 U136 ( .A(n65), .B(n66), .Y(in_17bit_b[10]) );
  XOR2X1 U137 ( .A(n47), .B(n45), .Y(in_17bit_b[5]) );
  NAND2X1 U138 ( .A(n46), .B(n21), .Y(n45) );
  XOR2X1 U139 ( .A(n55), .B(n52), .Y(in_17bit_b[7]) );
  XOR2X1 U140 ( .A(n63), .B(n60), .Y(in_17bit_b[9]) );
  NAND2X1 U141 ( .A(n44), .B(n43), .Y(n46) );
  INVX1 U142 ( .A(n48), .Y(n51) );
  INVX1 U143 ( .A(n56), .Y(n59) );
  INVX1 U144 ( .A(n64), .Y(n67) );
  NOR2X1 U145 ( .A(n68), .B(in_17bit[11]), .Y(sub_add_52_b0_carry[12]) );
  NAND2BXL U146 ( .AN(in_17bit[3]), .B(n41), .Y(n42) );
  INVX1 U147 ( .A(in_17bit[9]), .Y(n63) );
  INVX1 U148 ( .A(in_17bit[10]), .Y(n66) );
  INVX1 U149 ( .A(in_17bit[11]), .Y(n112) );
  INVX1 U150 ( .A(in_17bit[12]), .Y(n113) );
  INVX1 U151 ( .A(in_17bit[13]), .Y(n114) );
  INVX1 U152 ( .A(in_17bit[14]), .Y(n115) );
  INVX1 U153 ( .A(in_17bit[15]), .Y(n116) );
  NOR2XL U154 ( .A(in_8bit[4]), .B(in_8bit[3]), .Y(n30) );
  XOR2X4 U155 ( .A(n16), .B(n34), .Y(in_8bit_b[6]) );
  NOR3BX4 U156 ( .AN(n38), .B(n37), .C(n36), .Y(in_17bit_b[1]) );
  NOR2X4 U157 ( .A(n10), .B(n99), .Y(n96) );
  NOR2X4 U158 ( .A(n10), .B(n108), .Y(n106) );
  XNOR2X4 U159 ( .A(n106), .B(n107), .Y(out[15]) );
  XOR2X1 U160 ( .A(n110), .B(n111), .Y(N33) );
  XOR2X1 U161 ( .A(n22), .B(sub_add_52_b0_carry[16]), .Y(N21) );
  AND2X1 U162 ( .A(sub_add_52_b0_carry[15]), .B(n116), .Y(
        sub_add_52_b0_carry[16]) );
  XOR2X1 U163 ( .A(n116), .B(sub_add_52_b0_carry[15]), .Y(N20) );
  AND2X1 U164 ( .A(sub_add_52_b0_carry[14]), .B(n115), .Y(
        sub_add_52_b0_carry[15]) );
  XOR2X1 U165 ( .A(n115), .B(sub_add_52_b0_carry[14]), .Y(N19) );
  AND2X1 U166 ( .A(sub_add_52_b0_carry[13]), .B(n114), .Y(
        sub_add_52_b0_carry[14]) );
  XOR2X1 U167 ( .A(n114), .B(sub_add_52_b0_carry[13]), .Y(N18) );
  AND2X1 U168 ( .A(sub_add_52_b0_carry[12]), .B(n113), .Y(
        sub_add_52_b0_carry[13]) );
endmodule


module multi16_2_DW01_add_0 ( A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, 
        A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, 
        B_20_, B_19_, B_18_, B_17_, B_16_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, 
        SUM_17_, SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, 
        SUM_9_, SUM_8_, SUM_7_, SUM_6_, SUM_5_ );
  input A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_,
         A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, B_20_, B_19_,
         B_18_, B_17_, B_16_;
  output SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, SUM_15_,
         SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, SUM_7_,
         SUM_6_, SUM_5_;
  wire   n1, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39;

  INVX4 U2 ( .A(n33), .Y(n18) );
  INVX2 U3 ( .A(n19), .Y(SUM_15_) );
  OAI21X1 U4 ( .A0(n26), .A1(n27), .B0(n28), .Y(n22) );
  XOR2X2 U5 ( .A(n38), .B(n37), .Y(SUM_18_) );
  BUFX3 U6 ( .A(A_14_), .Y(SUM_14_) );
  INVX2 U7 ( .A(n29), .Y(n17) );
  INVX1 U8 ( .A(A_15_), .Y(n19) );
  OR2X4 U9 ( .A(B_16_), .B(A_16_), .Y(n1) );
  NAND2X1 U10 ( .A(B_19_), .B(A_19_), .Y(n28) );
  AOI21XL U11 ( .A0(n14), .A1(n31), .B0(n15), .Y(n26) );
  AND2X4 U12 ( .A(n33), .B(n1), .Y(SUM_16_) );
  NOR2BX2 U13 ( .AN(n28), .B(n27), .Y(n36) );
  NAND2X2 U14 ( .A(B_16_), .B(A_16_), .Y(n33) );
  XOR2X4 U15 ( .A(n35), .B(n36), .Y(SUM_19_) );
  AOI21X4 U16 ( .A0(n18), .A1(n17), .B0(n16), .Y(n37) );
  NOR2X2 U17 ( .A(B_18_), .B(A_18_), .Y(n30) );
  NOR2X4 U18 ( .A(B_17_), .B(A_17_), .Y(n29) );
  OAI21X2 U19 ( .A0(n37), .A1(n30), .B0(n32), .Y(n35) );
  XOR2X4 U20 ( .A(n18), .B(n39), .Y(SUM_17_) );
  NOR2X4 U21 ( .A(n29), .B(n16), .Y(n39) );
  INVX4 U22 ( .A(n34), .Y(n16) );
  NAND2X4 U23 ( .A(B_17_), .B(A_17_), .Y(n34) );
  NAND2X1 U24 ( .A(n32), .B(n14), .Y(n38) );
  INVXL U25 ( .A(n24), .Y(n13) );
  AOI21XL U26 ( .A0(n22), .A1(n23), .B0(n13), .Y(n21) );
  BUFX3 U27 ( .A(A_13_), .Y(SUM_13_) );
  INVXL U28 ( .A(n32), .Y(n15) );
  INVX1 U29 ( .A(n30), .Y(n14) );
  BUFX3 U30 ( .A(A_5_), .Y(SUM_5_) );
  BUFX3 U31 ( .A(A_6_), .Y(SUM_6_) );
  BUFX3 U32 ( .A(A_7_), .Y(SUM_7_) );
  BUFX3 U33 ( .A(A_8_), .Y(SUM_8_) );
  BUFX3 U34 ( .A(A_10_), .Y(SUM_10_) );
  BUFX4 U35 ( .A(A_12_), .Y(SUM_12_) );
  BUFX3 U36 ( .A(A_11_), .Y(SUM_11_) );
  BUFX3 U37 ( .A(A_9_), .Y(SUM_9_) );
  XOR2X1 U38 ( .A(n20), .B(n21), .Y(SUM_21_) );
  XNOR2X1 U39 ( .A(B_21_), .B(A_21_), .Y(n20) );
  XNOR2X1 U40 ( .A(n25), .B(n22), .Y(SUM_20_) );
  OAI21XL U41 ( .A0(n29), .A1(n33), .B0(n34), .Y(n31) );
  NAND2X1 U42 ( .A(n24), .B(n23), .Y(n25) );
  OR2X1 U43 ( .A(B_20_), .B(A_20_), .Y(n23) );
  NAND2X1 U44 ( .A(B_20_), .B(A_20_), .Y(n24) );
  NOR2X1 U45 ( .A(B_19_), .B(A_19_), .Y(n27) );
  NAND2X1 U46 ( .A(B_18_), .B(A_18_), .Y(n32) );
endmodule


module multi16_2_DW02_mult_0 ( A, B, PRODUCT_23_, PRODUCT_22_, PRODUCT_21_, 
        PRODUCT_20_, PRODUCT_19_, PRODUCT_18_, PRODUCT_17_, PRODUCT_16_, 
        PRODUCT_15_, PRODUCT_14_, PRODUCT_13_, PRODUCT_12_, PRODUCT_11_, 
        PRODUCT_10_, PRODUCT_9_, PRODUCT_8_, PRODUCT_7_ );
  input [16:0] A;
  input [7:0] B;
  output PRODUCT_23_, PRODUCT_22_, PRODUCT_21_, PRODUCT_20_, PRODUCT_19_,
         PRODUCT_18_, PRODUCT_17_, PRODUCT_16_, PRODUCT_15_, PRODUCT_14_,
         PRODUCT_13_, PRODUCT_12_, PRODUCT_11_, PRODUCT_10_, PRODUCT_9_,
         PRODUCT_8_, PRODUCT_7_;
  wire   ab_16__7_, ab_16__6_, ab_16__5_, ab_16__4_, ab_16__3_, ab_16__2_,
         ab_16__1_, ab_16__0_, ab_15__7_, ab_15__6_, ab_15__5_, ab_15__4_,
         ab_15__3_, ab_15__2_, ab_15__1_, ab_15__0_, ab_14__7_, ab_14__6_,
         ab_14__5_, ab_14__4_, ab_14__3_, ab_14__2_, ab_14__1_, ab_14__0_,
         ab_13__7_, ab_13__6_, ab_13__5_, ab_13__4_, ab_13__3_, ab_13__2_,
         ab_13__1_, ab_13__0_, ab_12__7_, ab_12__6_, ab_12__5_, ab_12__4_,
         ab_12__3_, ab_12__2_, ab_12__1_, ab_12__0_, ab_11__7_, ab_11__6_,
         ab_11__5_, ab_11__4_, ab_11__3_, ab_11__2_, ab_11__1_, ab_11__0_,
         ab_10__7_, ab_10__6_, ab_10__5_, ab_10__4_, ab_10__3_, ab_10__2_,
         ab_10__1_, ab_10__0_, ab_9__7_, ab_9__6_, ab_9__5_, ab_9__4_,
         ab_9__3_, ab_9__2_, ab_9__1_, ab_9__0_, ab_8__7_, ab_8__6_, ab_8__5_,
         ab_8__4_, ab_8__3_, ab_8__2_, ab_8__1_, ab_8__0_, ab_7__7_, ab_7__6_,
         ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_, ab_7__0_, ab_6__7_,
         ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_, ab_6__1_, ab_6__0_,
         ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_, ab_5__2_, ab_5__1_,
         ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_, ab_4__3_, ab_4__2_,
         ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_, ab_3__4_, ab_3__3_,
         ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_, ab_2__5_, ab_2__4_,
         ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_, ab_1__6_, ab_1__5_,
         ab_1__4_, ab_1__3_, ab_1__2_, ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_,
         ab_0__3_, ab_0__2_, CARRYB_16__6_, CARRYB_16__5_, CARRYB_16__4_,
         CARRYB_16__3_, CARRYB_16__2_, CARRYB_16__1_, CARRYB_16__0_,
         CARRYB_15__6_, CARRYB_15__5_, CARRYB_15__4_, CARRYB_15__3_,
         CARRYB_15__2_, CARRYB_15__1_, CARRYB_15__0_, CARRYB_14__6_,
         CARRYB_14__5_, CARRYB_14__4_, CARRYB_14__3_, CARRYB_14__2_,
         CARRYB_14__1_, CARRYB_14__0_, CARRYB_13__6_, CARRYB_13__5_,
         CARRYB_13__4_, CARRYB_13__3_, CARRYB_13__2_, CARRYB_13__1_,
         CARRYB_13__0_, CARRYB_12__6_, CARRYB_12__5_, CARRYB_12__4_,
         CARRYB_12__3_, CARRYB_12__2_, CARRYB_12__1_, CARRYB_12__0_,
         CARRYB_11__6_, CARRYB_11__5_, CARRYB_11__4_, CARRYB_11__3_,
         CARRYB_11__2_, CARRYB_11__1_, CARRYB_11__0_, CARRYB_10__6_,
         CARRYB_10__5_, CARRYB_10__4_, CARRYB_10__3_, CARRYB_10__2_,
         CARRYB_10__1_, CARRYB_10__0_, CARRYB_9__6_, CARRYB_9__5_,
         CARRYB_9__4_, CARRYB_9__3_, CARRYB_9__2_, CARRYB_9__1_, CARRYB_9__0_,
         CARRYB_8__6_, CARRYB_8__5_, CARRYB_8__4_, CARRYB_8__3_, CARRYB_8__2_,
         CARRYB_8__1_, CARRYB_8__0_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_,
         CARRYB_7__3_, CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_,
         CARRYB_6__5_, CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_,
         CARRYB_6__0_, CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_,
         CARRYB_5__2_, CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_,
         CARRYB_4__4_, CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_,
         CARRYB_3__6_, CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_,
         CARRYB_3__1_, CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_,
         CARRYB_2__3_, CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__0_,
         SUMB_16__6_, SUMB_16__5_, SUMB_16__4_, SUMB_16__3_, SUMB_16__2_,
         SUMB_16__1_, SUMB_16__0_, SUMB_15__6_, SUMB_15__5_, SUMB_15__4_,
         SUMB_15__3_, SUMB_15__2_, SUMB_15__1_, SUMB_14__6_, SUMB_14__5_,
         SUMB_14__4_, SUMB_14__3_, SUMB_14__2_, SUMB_14__1_, SUMB_13__6_,
         SUMB_13__5_, SUMB_13__4_, SUMB_13__3_, SUMB_13__2_, SUMB_13__1_,
         SUMB_12__6_, SUMB_12__5_, SUMB_12__4_, SUMB_12__3_, SUMB_12__2_,
         SUMB_12__1_, SUMB_11__6_, SUMB_11__5_, SUMB_11__4_, SUMB_11__3_,
         SUMB_11__2_, SUMB_11__1_, SUMB_10__6_, SUMB_10__5_, SUMB_10__4_,
         SUMB_10__3_, SUMB_10__2_, SUMB_10__1_, SUMB_9__6_, SUMB_9__5_,
         SUMB_9__4_, SUMB_9__3_, SUMB_9__2_, SUMB_9__1_, SUMB_8__6_,
         SUMB_8__5_, SUMB_8__4_, SUMB_8__3_, SUMB_8__2_, SUMB_8__1_,
         SUMB_7__6_, SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_,
         SUMB_7__1_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, PROD1_7_, A1_21_, A1_20_, A1_19_, A1_18_,
         A1_17_, A1_16_, A1_15_, A1_13_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_,
         A1_7_, A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66;

  ADDFHX4 S1_15_0 ( .A(ab_15__0_), .B(CARRYB_14__0_), .CI(SUMB_14__1_), .CO(
        CARRYB_15__0_), .S(A1_13_) );
  ADDFHX4 S1_14_0 ( .A(ab_14__0_), .B(CARRYB_13__0_), .CI(SUMB_13__1_), .CO(
        CARRYB_14__0_), .S(A1_12_) );
  ADDFHX4 S1_13_0 ( .A(ab_13__0_), .B(CARRYB_12__0_), .CI(SUMB_12__1_), .CO(
        CARRYB_13__0_), .S(A1_11_) );
  multi16_2_DW01_add_0 FS_1 ( .A_21_(A1_21_), .A_20_(A1_20_), .A_19_(A1_19_), 
        .A_18_(A1_18_), .A_17_(A1_17_), .A_16_(A1_16_), .A_15_(A1_15_), 
        .A_14_(SUMB_16__0_), .A_13_(A1_13_), .A_12_(A1_12_), .A_11_(A1_11_), 
        .A_10_(A1_10_), .A_9_(A1_9_), .A_8_(A1_8_), .A_7_(A1_7_), .A_6_(A1_6_), 
        .A_5_(PROD1_7_), .B_21_(n23), .B_20_(n48), .B_19_(n47), .B_18_(n46), 
        .B_17_(n45), .B_16_(n44), .SUM_21_(PRODUCT_23_), .SUM_20_(PRODUCT_22_), 
        .SUM_19_(PRODUCT_21_), .SUM_18_(PRODUCT_20_), .SUM_17_(PRODUCT_19_), 
        .SUM_16_(PRODUCT_18_), .SUM_15_(PRODUCT_17_), .SUM_14_(PRODUCT_16_), 
        .SUM_13_(PRODUCT_15_), .SUM_12_(PRODUCT_14_), .SUM_11_(PRODUCT_13_), 
        .SUM_10_(PRODUCT_12_), .SUM_9_(PRODUCT_11_), .SUM_8_(PRODUCT_10_), 
        .SUM_7_(PRODUCT_9_), .SUM_6_(PRODUCT_8_), .SUM_5_(PRODUCT_7_) );
  ADDFX2 S3_15_6 ( .A(ab_15__6_), .B(CARRYB_14__6_), .CI(ab_14__7_), .CO(
        CARRYB_15__6_), .S(SUMB_15__6_) );
  ADDFHX1 S2_15_5 ( .A(ab_15__5_), .B(CARRYB_14__5_), .CI(SUMB_14__6_), .CO(
        CARRYB_15__5_), .S(SUMB_15__5_) );
  ADDFHX4 S2_15_1 ( .A(ab_15__1_), .B(CARRYB_14__1_), .CI(SUMB_14__2_), .CO(
        CARRYB_15__1_), .S(SUMB_15__1_) );
  ADDFHX2 S2_2_5 ( .A(ab_2__5_), .B(n18), .CI(SUMB_1__6_), .CO(CARRYB_2__5_), 
        .S(SUMB_2__5_) );
  ADDFHX2 S3_13_6 ( .A(ab_13__6_), .B(CARRYB_12__6_), .CI(ab_12__7_), .CO(
        CARRYB_13__6_), .S(SUMB_13__6_) );
  ADDFHX4 S2_13_3 ( .A(ab_13__3_), .B(CARRYB_12__3_), .CI(SUMB_12__4_), .CO(
        CARRYB_13__3_), .S(SUMB_13__3_) );
  ADDFHX4 S3_9_6 ( .A(ab_9__6_), .B(CARRYB_8__6_), .CI(ab_8__7_), .CO(
        CARRYB_9__6_), .S(SUMB_9__6_) );
  ADDFHX4 S3_10_6 ( .A(ab_10__6_), .B(CARRYB_9__6_), .CI(ab_9__7_), .CO(
        CARRYB_10__6_), .S(SUMB_10__6_) );
  ADDFHX2 S2_10_5 ( .A(ab_10__5_), .B(CARRYB_9__5_), .CI(SUMB_9__6_), .CO(
        CARRYB_10__5_), .S(SUMB_10__5_) );
  ADDFHX4 S2_15_2 ( .A(ab_15__2_), .B(CARRYB_14__2_), .CI(SUMB_14__3_), .CO(
        CARRYB_15__2_), .S(SUMB_15__2_) );
  ADDFHX2 S2_9_3 ( .A(ab_9__3_), .B(CARRYB_8__3_), .CI(SUMB_8__4_), .CO(
        CARRYB_9__3_), .S(SUMB_9__3_) );
  ADDFHX4 S3_7_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(
        CARRYB_7__6_), .S(SUMB_7__6_) );
  ADDFHX4 S3_8_6 ( .A(ab_8__6_), .B(CARRYB_7__6_), .CI(ab_7__7_), .CO(
        CARRYB_8__6_), .S(SUMB_8__6_) );
  ADDFHX2 S2_8_3 ( .A(ab_8__3_), .B(CARRYB_7__3_), .CI(SUMB_7__4_), .CO(
        CARRYB_8__3_), .S(SUMB_8__3_) );
  ADDFHX4 S2_8_1 ( .A(ab_8__1_), .B(CARRYB_7__1_), .CI(SUMB_7__2_), .CO(
        CARRYB_8__1_), .S(SUMB_8__1_) );
  ADDFHX2 S2_15_3 ( .A(ab_15__3_), .B(CARRYB_14__3_), .CI(SUMB_14__4_), .CO(
        CARRYB_15__3_), .S(SUMB_15__3_) );
  ADDFHX4 S4_2 ( .A(ab_16__2_), .B(CARRYB_15__2_), .CI(SUMB_15__3_), .CO(
        CARRYB_16__2_), .S(SUMB_16__2_) );
  ADDFHX2 S2_9_5 ( .A(ab_9__5_), .B(CARRYB_8__5_), .CI(SUMB_8__6_), .CO(
        CARRYB_9__5_), .S(SUMB_9__5_) );
  ADDFHX4 S2_11_4 ( .A(ab_11__4_), .B(CARRYB_10__4_), .CI(SUMB_10__5_), .CO(
        CARRYB_11__4_), .S(SUMB_11__4_) );
  ADDFHX2 S2_11_5 ( .A(ab_11__5_), .B(CARRYB_10__5_), .CI(SUMB_10__6_), .CO(
        CARRYB_11__5_), .S(SUMB_11__5_) );
  ADDFHX4 S2_2_2 ( .A(ab_2__2_), .B(n21), .CI(SUMB_1__3_), .CO(CARRYB_2__2_), 
        .S(SUMB_2__2_) );
  ADDFHX4 S2_11_2 ( .A(ab_11__2_), .B(CARRYB_10__2_), .CI(SUMB_10__3_), .CO(
        CARRYB_11__2_), .S(SUMB_11__2_) );
  ADDFHX4 S3_2_6 ( .A(ab_2__6_), .B(n19), .CI(ab_1__7_), .CO(CARRYB_2__6_), 
        .S(SUMB_2__6_) );
  ADDFHX4 S3_12_6 ( .A(ab_12__6_), .B(CARRYB_11__6_), .CI(ab_11__7_), .CO(
        CARRYB_12__6_), .S(SUMB_12__6_) );
  ADDFHX4 S1_8_0 ( .A(ab_8__0_), .B(CARRYB_7__0_), .CI(SUMB_7__1_), .CO(
        CARRYB_8__0_), .S(A1_6_) );
  ADDFHX2 S2_9_2 ( .A(ab_9__2_), .B(CARRYB_8__2_), .CI(SUMB_8__3_), .CO(
        CARRYB_9__2_), .S(SUMB_9__2_) );
  ADDFHX4 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  ADDFHX4 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  ADDFHX4 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  ADDFHX4 S1_11_0 ( .A(ab_11__0_), .B(CARRYB_10__0_), .CI(SUMB_10__1_), .CO(
        CARRYB_11__0_), .S(A1_9_) );
  ADDFHX4 S2_10_1 ( .A(ab_10__1_), .B(CARRYB_9__1_), .CI(SUMB_9__2_), .CO(
        CARRYB_10__1_), .S(SUMB_10__1_) );
  ADDFHX4 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  ADDFHX4 S2_7_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  ADDFHX4 S2_9_4 ( .A(ab_9__4_), .B(CARRYB_8__4_), .CI(SUMB_8__5_), .CO(
        CARRYB_9__4_), .S(SUMB_9__4_) );
  ADDFHX4 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  ADDFHX2 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  ADDFHX2 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  ADDFHX4 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  ADDFHX2 S2_2_3 ( .A(ab_2__3_), .B(n22), .CI(SUMB_1__4_), .CO(CARRYB_2__3_), 
        .S(SUMB_2__3_) );
  ADDFHX4 S2_14_3 ( .A(ab_14__3_), .B(CARRYB_13__3_), .CI(SUMB_13__4_), .CO(
        CARRYB_14__3_), .S(SUMB_14__3_) );
  ADDFHX4 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  ADDFHX4 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  ADDFHX4 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  ADDFHX4 S2_7_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  ADDFHX4 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  ADDFHX4 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  ADDFHX4 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  ADDFHX4 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  ADDFHX4 S1_10_0 ( .A(ab_10__0_), .B(CARRYB_9__0_), .CI(SUMB_9__1_), .CO(
        CARRYB_10__0_), .S(A1_8_) );
  ADDFHX4 S2_7_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  ADDFHX4 S2_8_2 ( .A(ab_8__2_), .B(CARRYB_7__2_), .CI(SUMB_7__3_), .CO(
        CARRYB_8__2_), .S(SUMB_8__2_) );
  ADDFHX4 S3_11_6 ( .A(ab_11__6_), .B(CARRYB_10__6_), .CI(ab_10__7_), .CO(
        CARRYB_11__6_), .S(SUMB_11__6_) );
  ADDFHX2 S2_15_4 ( .A(ab_15__4_), .B(CARRYB_14__4_), .CI(SUMB_14__5_), .CO(
        CARRYB_15__4_), .S(SUMB_15__4_) );
  ADDFHX4 S2_10_4 ( .A(ab_10__4_), .B(CARRYB_9__4_), .CI(SUMB_9__5_), .CO(
        CARRYB_10__4_), .S(SUMB_10__4_) );
  ADDFHX4 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  ADDFHX4 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  ADDFHX4 S2_7_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  ADDFHX4 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  ADDFHX2 S2_13_2 ( .A(ab_13__2_), .B(CARRYB_12__2_), .CI(SUMB_12__3_), .CO(
        CARRYB_13__2_), .S(SUMB_13__2_) );
  ADDFHX4 S2_14_1 ( .A(ab_14__1_), .B(CARRYB_13__1_), .CI(SUMB_13__2_), .CO(
        CARRYB_14__1_), .S(SUMB_14__1_) );
  ADDFHX2 S2_10_2 ( .A(ab_10__2_), .B(CARRYB_9__2_), .CI(SUMB_9__3_), .CO(
        CARRYB_10__2_), .S(SUMB_10__2_) );
  ADDFHX4 S2_11_1 ( .A(ab_11__1_), .B(CARRYB_10__1_), .CI(SUMB_10__2_), .CO(
        CARRYB_11__1_), .S(SUMB_11__1_) );
  ADDFHX2 S2_12_2 ( .A(ab_12__2_), .B(CARRYB_11__2_), .CI(SUMB_11__3_), .CO(
        CARRYB_12__2_), .S(SUMB_12__2_) );
  ADDFHX4 S2_13_1 ( .A(ab_13__1_), .B(CARRYB_12__1_), .CI(SUMB_12__2_), .CO(
        CARRYB_13__1_), .S(SUMB_13__1_) );
  ADDFHX1 S3_14_6 ( .A(ab_14__6_), .B(CARRYB_13__6_), .CI(ab_13__7_), .CO(
        CARRYB_14__6_), .S(SUMB_14__6_) );
  ADDFX2 S4_5 ( .A(ab_16__5_), .B(CARRYB_15__5_), .CI(SUMB_15__6_), .CO(
        CARRYB_16__5_), .S(SUMB_16__5_) );
  ADDFHX1 S4_4 ( .A(ab_16__4_), .B(CARRYB_15__4_), .CI(SUMB_15__5_), .CO(
        CARRYB_16__4_), .S(SUMB_16__4_) );
  ADDFHX2 S4_0 ( .A(ab_16__0_), .B(CARRYB_15__0_), .CI(SUMB_15__1_), .CO(
        CARRYB_16__0_), .S(SUMB_16__0_) );
  ADDFHX2 S4_1 ( .A(ab_16__1_), .B(CARRYB_15__1_), .CI(SUMB_15__2_), .CO(
        CARRYB_16__1_), .S(SUMB_16__1_) );
  ADDFHX2 S4_3 ( .A(ab_16__3_), .B(CARRYB_15__3_), .CI(SUMB_15__4_), .CO(
        CARRYB_16__3_), .S(SUMB_16__3_) );
  ADDFHX2 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  ADDFHX2 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  ADDFHX2 S1_9_0 ( .A(ab_9__0_), .B(CARRYB_8__0_), .CI(SUMB_8__1_), .CO(
        CARRYB_9__0_), .S(A1_7_) );
  ADDFHX2 S2_9_1 ( .A(ab_9__1_), .B(CARRYB_8__1_), .CI(SUMB_8__2_), .CO(
        CARRYB_9__1_), .S(SUMB_9__1_) );
  ADDFHX2 S2_13_4 ( .A(ab_13__4_), .B(CARRYB_12__4_), .CI(SUMB_12__5_), .CO(
        CARRYB_13__4_), .S(SUMB_13__4_) );
  ADDFHX2 S2_8_5 ( .A(ab_8__5_), .B(CARRYB_7__5_), .CI(SUMB_7__6_), .CO(
        CARRYB_8__5_), .S(SUMB_8__5_) );
  ADDFHX2 S2_7_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  ADDFHX2 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  ADDFHX2 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  ADDFHX2 S2_2_4 ( .A(ab_2__4_), .B(n17), .CI(SUMB_1__5_), .CO(CARRYB_2__4_), 
        .S(SUMB_2__4_) );
  ADDFHX2 S2_12_4 ( .A(ab_12__4_), .B(CARRYB_11__4_), .CI(SUMB_11__5_), .CO(
        CARRYB_12__4_), .S(SUMB_12__4_) );
  ADDFHX2 S2_2_1 ( .A(ab_2__1_), .B(n20), .CI(SUMB_1__2_), .CO(CARRYB_2__1_), 
        .S(SUMB_2__1_) );
  ADDFHX4 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  ADDFHX4 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  ADDFHX4 S1_7_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(PROD1_7_) );
  ADDFHX2 S2_13_5 ( .A(ab_13__5_), .B(CARRYB_12__5_), .CI(SUMB_12__6_), .CO(
        CARRYB_13__5_), .S(SUMB_13__5_) );
  ADDFHX4 S2_10_3 ( .A(ab_10__3_), .B(CARRYB_9__3_), .CI(SUMB_9__4_), .CO(
        CARRYB_10__3_), .S(SUMB_10__3_) );
  ADDFHX2 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  ADDFHX4 S2_12_1 ( .A(ab_12__1_), .B(CARRYB_11__1_), .CI(SUMB_11__2_), .CO(
        CARRYB_12__1_), .S(SUMB_12__1_) );
  ADDFHX4 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  ADDFHX4 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  ADDFHX1 S5_6 ( .A(ab_16__6_), .B(CARRYB_15__6_), .CI(ab_15__7_), .CO(
        CARRYB_16__6_), .S(SUMB_16__6_) );
  ADDFHX4 S1_12_0 ( .A(ab_12__0_), .B(CARRYB_11__0_), .CI(SUMB_11__1_), .CO(
        CARRYB_12__0_), .S(A1_10_) );
  AND2X2 U2 ( .A(A[3]), .B(B[6]), .Y(ab_3__6_) );
  NAND3X4 U3 ( .A(n10), .B(n11), .C(n12), .Y(CARRYB_4__1_) );
  NAND2X2 U4 ( .A(ab_4__1_), .B(CARRYB_3__1_), .Y(n11) );
  NAND2X2 U5 ( .A(ab_4__1_), .B(SUMB_3__2_), .Y(n10) );
  NOR2X2 U6 ( .A(n56), .B(n50), .Y(ab_0__3_) );
  CLKINVX3 U7 ( .A(B[3]), .Y(n56) );
  INVX2 U8 ( .A(B[2]), .Y(n57) );
  XOR2X4 U9 ( .A(CARRYB_13__5_), .B(n35), .Y(SUMB_14__5_) );
  XOR2X4 U10 ( .A(SUMB_13__6_), .B(ab_14__5_), .Y(n35) );
  CLKINVX1 U11 ( .A(A[0]), .Y(n50) );
  AND2X4 U12 ( .A(ab_0__7_), .B(ab_1__6_), .Y(n19) );
  AND2X1 U13 ( .A(A[2]), .B(B[0]), .Y(ab_2__0_) );
  AND2X1 U14 ( .A(A[2]), .B(B[2]), .Y(ab_2__2_) );
  AND2X1 U15 ( .A(A[2]), .B(B[3]), .Y(ab_2__3_) );
  AND2X1 U16 ( .A(A[2]), .B(B[4]), .Y(ab_2__4_) );
  XOR3X2 U17 ( .A(CARRYB_7__4_), .B(ab_8__4_), .C(SUMB_7__5_), .Y(SUMB_8__4_)
         );
  NAND2X2 U18 ( .A(SUMB_7__5_), .B(CARRYB_7__4_), .Y(n3) );
  NAND2X1 U19 ( .A(ab_8__4_), .B(CARRYB_7__4_), .Y(n4) );
  NAND2X2 U20 ( .A(ab_8__4_), .B(SUMB_7__5_), .Y(n5) );
  NAND3X4 U21 ( .A(n5), .B(n3), .C(n4), .Y(CARRYB_8__4_) );
  XOR3X2 U22 ( .A(ab_3__1_), .B(CARRYB_2__1_), .C(SUMB_2__2_), .Y(SUMB_3__1_)
         );
  NAND2X1 U23 ( .A(ab_3__1_), .B(CARRYB_2__1_), .Y(n6) );
  NAND2X1 U24 ( .A(ab_3__1_), .B(SUMB_2__2_), .Y(n7) );
  NAND2X1 U25 ( .A(CARRYB_2__1_), .B(SUMB_2__2_), .Y(n8) );
  NAND3X4 U26 ( .A(n6), .B(n7), .C(n8), .Y(CARRYB_3__1_) );
  XOR2X4 U27 ( .A(ab_4__1_), .B(SUMB_3__2_), .Y(n9) );
  XOR2X4 U28 ( .A(n9), .B(CARRYB_3__1_), .Y(SUMB_4__1_) );
  NAND2X2 U29 ( .A(SUMB_3__2_), .B(CARRYB_3__1_), .Y(n12) );
  XOR3X4 U30 ( .A(CARRYB_10__3_), .B(ab_11__3_), .C(SUMB_10__4_), .Y(
        SUMB_11__3_) );
  NAND2X1 U31 ( .A(SUMB_10__4_), .B(CARRYB_10__3_), .Y(n13) );
  NAND2X1 U32 ( .A(ab_11__3_), .B(CARRYB_10__3_), .Y(n14) );
  NAND2X2 U33 ( .A(ab_11__3_), .B(SUMB_10__4_), .Y(n15) );
  NAND3X2 U34 ( .A(n15), .B(n13), .C(n14), .Y(CARRYB_11__3_) );
  NAND2X2 U35 ( .A(SUMB_11__4_), .B(CARRYB_11__3_), .Y(n39) );
  NAND3X4 U36 ( .A(n27), .B(n25), .C(n26), .Y(CARRYB_12__5_) );
  NOR2X4 U37 ( .A(n53), .B(n50), .Y(ab_0__6_) );
  INVX3 U38 ( .A(B[6]), .Y(n53) );
  NOR2X1 U39 ( .A(n65), .B(n42), .Y(ab_12__5_) );
  NAND2X1 U40 ( .A(ab_14__4_), .B(SUMB_13__5_), .Y(n30) );
  NAND2X1 U41 ( .A(SUMB_13__5_), .B(CARRYB_13__4_), .Y(n28) );
  NAND2X1 U42 ( .A(ab_12__5_), .B(CARRYB_11__5_), .Y(n26) );
  NOR2X1 U43 ( .A(n59), .B(n50), .Y(ab_0__7_) );
  NOR2X1 U44 ( .A(n54), .B(n50), .Y(ab_0__5_) );
  NOR2X1 U45 ( .A(n63), .B(n43), .Y(ab_14__4_) );
  NAND2X1 U46 ( .A(ab_14__2_), .B(CARRYB_13__2_), .Y(n33) );
  NAND2X1 U47 ( .A(SUMB_13__3_), .B(CARRYB_13__2_), .Y(n32) );
  NAND2X1 U48 ( .A(ab_14__4_), .B(CARRYB_13__4_), .Y(n29) );
  NOR2X1 U49 ( .A(n63), .B(n42), .Y(ab_14__5_) );
  NAND2X1 U50 ( .A(SUMB_11__6_), .B(CARRYB_11__5_), .Y(n25) );
  XOR2X1 U51 ( .A(CARRYB_16__0_), .B(SUMB_16__1_), .Y(A1_15_) );
  AND2X2 U53 ( .A(ab_0__5_), .B(ab_1__4_), .Y(n17) );
  AND2X2 U54 ( .A(ab_0__6_), .B(ab_1__5_), .Y(n18) );
  INVX1 U55 ( .A(B[0]), .Y(n49) );
  AND2X2 U56 ( .A(ab_0__2_), .B(n60), .Y(n20) );
  AND2X2 U57 ( .A(ab_0__3_), .B(ab_1__2_), .Y(n21) );
  AND2X2 U58 ( .A(ab_0__4_), .B(ab_1__3_), .Y(n22) );
  AND2X2 U59 ( .A(CARRYB_16__5_), .B(SUMB_16__6_), .Y(n23) );
  XOR2X1 U60 ( .A(ab_1__6_), .B(ab_0__7_), .Y(SUMB_1__6_) );
  XOR2X2 U61 ( .A(CARRYB_11__5_), .B(n24), .Y(SUMB_12__5_) );
  XOR2X4 U62 ( .A(SUMB_11__6_), .B(ab_12__5_), .Y(n24) );
  AND2X2 U63 ( .A(A[1]), .B(B[6]), .Y(ab_1__6_) );
  XOR2X4 U64 ( .A(CARRYB_16__1_), .B(SUMB_16__2_), .Y(A1_16_) );
  NAND3X4 U65 ( .A(n41), .B(n39), .C(n40), .Y(CARRYB_12__3_) );
  XOR3X2 U66 ( .A(CARRYB_11__3_), .B(ab_12__3_), .C(SUMB_11__4_), .Y(
        SUMB_12__3_) );
  NAND2X2 U67 ( .A(ab_14__2_), .B(SUMB_13__3_), .Y(n34) );
  NAND3X4 U68 ( .A(n34), .B(n32), .C(n33), .Y(CARRYB_14__2_) );
  XOR2XL U69 ( .A(n60), .B(ab_0__2_), .Y(SUMB_1__1_) );
  NAND2X1 U70 ( .A(ab_12__3_), .B(SUMB_11__4_), .Y(n41) );
  XOR2X2 U71 ( .A(CARRYB_16__3_), .B(SUMB_16__4_), .Y(A1_18_) );
  XOR3X4 U72 ( .A(CARRYB_13__4_), .B(ab_14__4_), .C(SUMB_13__5_), .Y(
        SUMB_14__4_) );
  AND2X2 U73 ( .A(A[1]), .B(B[3]), .Y(ab_1__3_) );
  AND2X4 U74 ( .A(CARRYB_16__1_), .B(SUMB_16__2_), .Y(n45) );
  XOR2X2 U75 ( .A(CARRYB_13__2_), .B(n31), .Y(SUMB_14__2_) );
  NAND2XL U76 ( .A(ab_12__5_), .B(SUMB_11__6_), .Y(n27) );
  NAND3X2 U77 ( .A(n30), .B(n28), .C(n29), .Y(CARRYB_14__4_) );
  XOR2X4 U78 ( .A(SUMB_13__3_), .B(ab_14__2_), .Y(n31) );
  NAND2X1 U79 ( .A(SUMB_13__6_), .B(CARRYB_13__5_), .Y(n36) );
  NAND2X1 U80 ( .A(ab_14__5_), .B(CARRYB_13__5_), .Y(n37) );
  NAND2XL U81 ( .A(ab_14__5_), .B(SUMB_13__6_), .Y(n38) );
  NAND3X2 U82 ( .A(n38), .B(n36), .C(n37), .Y(CARRYB_14__5_) );
  NAND2X1 U83 ( .A(ab_12__3_), .B(CARRYB_11__3_), .Y(n40) );
  NOR2X1 U84 ( .A(n65), .B(n56), .Y(ab_12__3_) );
  AND2X2 U85 ( .A(A[1]), .B(B[4]), .Y(ab_1__4_) );
  AND2X2 U86 ( .A(A[1]), .B(B[5]), .Y(ab_1__5_) );
  AND2X1 U87 ( .A(A[1]), .B(B[2]), .Y(ab_1__2_) );
  NAND2XL U88 ( .A(A[1]), .B(B[1]), .Y(n52) );
  XOR2X4 U89 ( .A(CARRYB_16__2_), .B(SUMB_16__3_), .Y(A1_17_) );
  INVX1 U90 ( .A(B[5]), .Y(n42) );
  INVX2 U91 ( .A(B[4]), .Y(n55) );
  INVX2 U92 ( .A(B[7]), .Y(n59) );
  INVX1 U93 ( .A(n52), .Y(n60) );
  AND2X1 U94 ( .A(A[10]), .B(B[2]), .Y(ab_10__2_) );
  NOR2XL U95 ( .A(n61), .B(n42), .Y(ab_16__5_) );
  AND2X1 U96 ( .A(A[4]), .B(B[1]), .Y(ab_4__1_) );
  AND2X1 U97 ( .A(A[7]), .B(B[0]), .Y(ab_7__0_) );
  AND2X1 U98 ( .A(A[6]), .B(B[0]), .Y(ab_6__0_) );
  AND2X1 U99 ( .A(A[6]), .B(B[1]), .Y(ab_6__1_) );
  INVXL U100 ( .A(B[1]), .Y(n58) );
  BUFX3 U101 ( .A(n55), .Y(n43) );
  NOR2X1 U102 ( .A(n55), .B(n50), .Y(ab_0__4_) );
  AND2X1 U103 ( .A(A[3]), .B(B[0]), .Y(ab_3__0_) );
  NOR2XL U104 ( .A(n52), .B(n51), .Y(CARRYB_1__0_) );
  NOR2XL U105 ( .A(n66), .B(n59), .Y(ab_11__7_) );
  NOR2XL U106 ( .A(n64), .B(n59), .Y(ab_13__7_) );
  NOR2XL U107 ( .A(n66), .B(n58), .Y(ab_11__1_) );
  NOR2XL U108 ( .A(n65), .B(n58), .Y(ab_12__1_) );
  NOR2XL U109 ( .A(n61), .B(n59), .Y(ab_16__7_) );
  AND2X1 U110 ( .A(A[4]), .B(B[6]), .Y(ab_4__6_) );
  AND2X1 U111 ( .A(A[5]), .B(B[6]), .Y(ab_5__6_) );
  AND2X2 U112 ( .A(CARRYB_16__0_), .B(SUMB_16__1_), .Y(n44) );
  XOR2X1 U113 ( .A(CARRYB_16__4_), .B(SUMB_16__5_), .Y(A1_19_) );
  AND2X1 U114 ( .A(CARRYB_16__2_), .B(SUMB_16__3_), .Y(n46) );
  AND2X2 U115 ( .A(CARRYB_16__3_), .B(SUMB_16__4_), .Y(n47) );
  AND2X2 U116 ( .A(CARRYB_16__4_), .B(SUMB_16__5_), .Y(n48) );
  AND2X2 U117 ( .A(A[4]), .B(B[2]), .Y(ab_4__2_) );
  NOR2X1 U118 ( .A(n61), .B(n58), .Y(ab_16__1_) );
  NOR2X1 U119 ( .A(n61), .B(n43), .Y(ab_16__4_) );
  NOR2BX1 U120 ( .AN(B[0]), .B(n61), .Y(ab_16__0_) );
  AND2X2 U121 ( .A(A[5]), .B(B[2]), .Y(ab_5__2_) );
  AND2X2 U122 ( .A(A[10]), .B(B[1]), .Y(ab_10__1_) );
  AND2X2 U123 ( .A(A[9]), .B(B[2]), .Y(ab_9__2_) );
  AND2X2 U124 ( .A(A[9]), .B(B[1]), .Y(ab_9__1_) );
  AND2X1 U125 ( .A(A[10]), .B(B[3]), .Y(ab_10__3_) );
  AND2X1 U126 ( .A(A[9]), .B(B[3]), .Y(ab_9__3_) );
  AND2X2 U127 ( .A(A[8]), .B(B[2]), .Y(ab_8__2_) );
  AND2X2 U128 ( .A(A[10]), .B(B[0]), .Y(ab_10__0_) );
  AND2X1 U129 ( .A(A[8]), .B(B[3]), .Y(ab_8__3_) );
  AND2X1 U130 ( .A(A[10]), .B(B[4]), .Y(ab_10__4_) );
  AND2X2 U131 ( .A(A[8]), .B(B[1]), .Y(ab_8__1_) );
  AND2X1 U132 ( .A(A[9]), .B(B[4]), .Y(ab_9__4_) );
  AND2X1 U133 ( .A(A[7]), .B(B[3]), .Y(ab_7__3_) );
  AND2X1 U134 ( .A(A[8]), .B(B[4]), .Y(ab_8__4_) );
  AND2X2 U135 ( .A(A[7]), .B(B[2]), .Y(ab_7__2_) );
  AND2X1 U136 ( .A(A[7]), .B(B[4]), .Y(ab_7__4_) );
  AND2X2 U137 ( .A(A[9]), .B(B[0]), .Y(ab_9__0_) );
  AND2X2 U138 ( .A(A[6]), .B(B[2]), .Y(ab_6__2_) );
  AND2X2 U139 ( .A(A[7]), .B(B[1]), .Y(ab_7__1_) );
  AND2X2 U140 ( .A(A[5]), .B(B[1]), .Y(ab_5__1_) );
  AND2X1 U141 ( .A(A[4]), .B(B[3]), .Y(ab_4__3_) );
  AND2X1 U142 ( .A(A[5]), .B(B[3]), .Y(ab_5__3_) );
  AND2X1 U143 ( .A(A[6]), .B(B[3]), .Y(ab_6__3_) );
  AND2X1 U144 ( .A(A[4]), .B(B[4]), .Y(ab_4__4_) );
  AND2X1 U145 ( .A(A[5]), .B(B[4]), .Y(ab_5__4_) );
  AND2X1 U146 ( .A(A[6]), .B(B[4]), .Y(ab_6__4_) );
  AND2X2 U147 ( .A(A[8]), .B(B[0]), .Y(ab_8__0_) );
  AND2X2 U148 ( .A(A[5]), .B(B[0]), .Y(ab_5__0_) );
  AND2X2 U149 ( .A(A[4]), .B(B[0]), .Y(ab_4__0_) );
  INVX1 U150 ( .A(B[5]), .Y(n54) );
  XOR2X1 U151 ( .A(CARRYB_16__5_), .B(SUMB_16__6_), .Y(A1_20_) );
  XOR2X1 U152 ( .A(CARRYB_16__6_), .B(ab_16__7_), .Y(A1_21_) );
  NOR2XL U153 ( .A(n61), .B(n53), .Y(ab_16__6_) );
  NOR2X1 U154 ( .A(n62), .B(n59), .Y(ab_15__7_) );
  NOR2XL U155 ( .A(n62), .B(n43), .Y(ab_15__4_) );
  NOR2X1 U156 ( .A(n63), .B(n58), .Y(ab_14__1_) );
  NOR2X1 U157 ( .A(n64), .B(n58), .Y(ab_13__1_) );
  NOR2XL U158 ( .A(n65), .B(n43), .Y(ab_12__4_) );
  NOR2XL U159 ( .A(n66), .B(n43), .Y(ab_11__4_) );
  AND2X1 U160 ( .A(A[3]), .B(B[1]), .Y(ab_3__1_) );
  AND2X1 U161 ( .A(A[3]), .B(B[4]), .Y(ab_3__4_) );
  AND2X1 U162 ( .A(A[10]), .B(B[5]), .Y(ab_10__5_) );
  AND2X1 U163 ( .A(A[9]), .B(B[5]), .Y(ab_9__5_) );
  AND2X1 U164 ( .A(A[4]), .B(B[5]), .Y(ab_4__5_) );
  AND2X1 U165 ( .A(A[8]), .B(B[5]), .Y(ab_8__5_) );
  AND2X1 U166 ( .A(A[5]), .B(B[5]), .Y(ab_5__5_) );
  AND2X1 U167 ( .A(A[7]), .B(B[5]), .Y(ab_7__5_) );
  AND2X1 U168 ( .A(A[6]), .B(B[5]), .Y(ab_6__5_) );
  NOR2X1 U169 ( .A(n65), .B(n59), .Y(ab_12__7_) );
  NOR2XL U170 ( .A(n64), .B(n53), .Y(ab_13__6_) );
  NOR2XL U171 ( .A(n65), .B(n53), .Y(ab_12__6_) );
  NOR2XL U172 ( .A(n64), .B(n43), .Y(ab_13__4_) );
  AND2X1 U173 ( .A(A[3]), .B(B[2]), .Y(ab_3__2_) );
  AND2X1 U174 ( .A(A[2]), .B(B[1]), .Y(ab_2__1_) );
  XOR2X1 U175 ( .A(ab_1__2_), .B(ab_0__3_), .Y(SUMB_1__2_) );
  XOR2X1 U176 ( .A(ab_1__3_), .B(ab_0__4_), .Y(SUMB_1__3_) );
  XOR2X1 U177 ( .A(ab_1__5_), .B(ab_0__6_), .Y(SUMB_1__5_) );
  XOR2X1 U178 ( .A(ab_1__4_), .B(ab_0__5_), .Y(SUMB_1__4_) );
  AND2X1 U179 ( .A(A[2]), .B(B[5]), .Y(ab_2__5_) );
  NOR2X1 U180 ( .A(n62), .B(n58), .Y(ab_15__1_) );
  NOR2XL U181 ( .A(n62), .B(n42), .Y(ab_15__5_) );
  AND2X1 U182 ( .A(A[3]), .B(B[5]), .Y(ab_3__5_) );
  NOR2X1 U183 ( .A(n63), .B(n59), .Y(ab_14__7_) );
  NOR2XL U184 ( .A(n62), .B(n53), .Y(ab_15__6_) );
  NOR2XL U185 ( .A(n63), .B(n53), .Y(ab_14__6_) );
  AND2X1 U186 ( .A(A[3]), .B(B[3]), .Y(ab_3__3_) );
  INVX1 U187 ( .A(A[16]), .Y(n61) );
  INVX1 U188 ( .A(A[14]), .Y(n63) );
  INVX1 U189 ( .A(A[15]), .Y(n62) );
  INVX1 U190 ( .A(A[11]), .Y(n66) );
  INVX1 U191 ( .A(A[12]), .Y(n65) );
  INVX1 U192 ( .A(A[13]), .Y(n64) );
  NAND2XL U193 ( .A(A[0]), .B(B[0]), .Y(n51) );
  AND2X1 U194 ( .A(A[9]), .B(B[6]), .Y(ab_9__6_) );
  AND2X1 U195 ( .A(A[8]), .B(B[6]), .Y(ab_8__6_) );
  AND2X1 U196 ( .A(A[7]), .B(B[6]), .Y(ab_7__6_) );
  AND2X1 U197 ( .A(A[6]), .B(B[6]), .Y(ab_6__6_) );
  NOR2XL U198 ( .A(n66), .B(n53), .Y(ab_11__6_) );
  AND2X1 U199 ( .A(A[10]), .B(B[6]), .Y(ab_10__6_) );
  NOR2XL U200 ( .A(n61), .B(n56), .Y(ab_16__3_) );
  NOR2XL U201 ( .A(n62), .B(n56), .Y(ab_15__3_) );
  NOR2XL U202 ( .A(n63), .B(n56), .Y(ab_14__3_) );
  NOR2XL U203 ( .A(n64), .B(n56), .Y(ab_13__3_) );
  NOR2XL U204 ( .A(n66), .B(n56), .Y(ab_11__3_) );
  NOR2XL U205 ( .A(n66), .B(n42), .Y(ab_11__5_) );
  NOR2XL U206 ( .A(n64), .B(n42), .Y(ab_13__5_) );
  AND2X1 U207 ( .A(A[10]), .B(B[7]), .Y(ab_10__7_) );
  AND2X1 U208 ( .A(A[9]), .B(B[7]), .Y(ab_9__7_) );
  AND2X1 U209 ( .A(A[8]), .B(B[7]), .Y(ab_8__7_) );
  AND2X1 U210 ( .A(A[7]), .B(B[7]), .Y(ab_7__7_) );
  AND2X1 U211 ( .A(A[6]), .B(B[7]), .Y(ab_6__7_) );
  AND2X1 U212 ( .A(A[5]), .B(B[7]), .Y(ab_5__7_) );
  AND2X1 U213 ( .A(A[4]), .B(B[7]), .Y(ab_4__7_) );
  AND2X1 U214 ( .A(A[3]), .B(B[7]), .Y(ab_3__7_) );
  AND2X1 U215 ( .A(A[2]), .B(B[7]), .Y(ab_2__7_) );
  AND2X2 U216 ( .A(A[2]), .B(B[6]), .Y(ab_2__6_) );
  NOR2XL U217 ( .A(n61), .B(n57), .Y(ab_16__2_) );
  NOR2XL U218 ( .A(n62), .B(n57), .Y(ab_15__2_) );
  NOR2XL U219 ( .A(n63), .B(n57), .Y(ab_14__2_) );
  NOR2XL U220 ( .A(n64), .B(n57), .Y(ab_13__2_) );
  NOR2XL U221 ( .A(n65), .B(n57), .Y(ab_12__2_) );
  NOR2XL U222 ( .A(n66), .B(n57), .Y(ab_11__2_) );
  NOR2X2 U223 ( .A(n57), .B(n50), .Y(ab_0__2_) );
  AND2X1 U224 ( .A(A[1]), .B(B[7]), .Y(ab_1__7_) );
  NOR2X1 U226 ( .A(n49), .B(n62), .Y(ab_15__0_) );
  NOR2X1 U227 ( .A(n49), .B(n63), .Y(ab_14__0_) );
  NOR2X1 U228 ( .A(n49), .B(n64), .Y(ab_13__0_) );
  NOR2X1 U229 ( .A(n49), .B(n65), .Y(ab_12__0_) );
  NOR2X1 U230 ( .A(n49), .B(n66), .Y(ab_11__0_) );
endmodule


module multi16_2 ( in_17bit, in_8bit, out );
  input [16:0] in_17bit;
  input [7:0] in_8bit;
  output [16:0] out;
  wire   N21, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126;
  wire   [16:1] in_17bit_b;
  wire   [6:1] in_8bit_b;
  wire   [23:8] mul;
  wire   [16:12] sub_add_52_b0_carry;

  multi16_2_DW02_mult_0 mult_55 ( .A({in_17bit_b, in_17bit[0]}), .B({n18, 
        in_8bit_b, n29}), .PRODUCT_23_(mul[23]), .PRODUCT_22_(mul[22]), 
        .PRODUCT_21_(mul[21]), .PRODUCT_20_(mul[20]), .PRODUCT_19_(mul[19]), 
        .PRODUCT_18_(mul[18]), .PRODUCT_17_(mul[17]), .PRODUCT_16_(mul[16]), 
        .PRODUCT_15_(mul[15]), .PRODUCT_14_(mul[14]), .PRODUCT_13_(mul[13]), 
        .PRODUCT_12_(mul[12]), .PRODUCT_11_(mul[11]), .PRODUCT_10_(mul[10]), 
        .PRODUCT_9_(mul[9]), .PRODUCT_8_(mul[8]), .PRODUCT_7_(out[0]) );
  CLKINVX3 U2 ( .A(n105), .Y(n107) );
  OAI21X2 U3 ( .A0(in_8bit[1]), .A1(n29), .B0(in_8bit[7]), .Y(n35) );
  NOR3X1 U4 ( .A(in_8bit[3]), .B(in_8bit[1]), .C(n44), .Y(n39) );
  INVX4 U5 ( .A(n25), .Y(n114) );
  NOR2X4 U6 ( .A(mul[18]), .B(n108), .Y(n25) );
  NAND2BX2 U7 ( .AN(n29), .B(n38), .Y(n41) );
  NAND2X2 U8 ( .A(in_17bit[2]), .B(n2), .Y(n3) );
  NAND2X2 U9 ( .A(n1), .B(n53), .Y(n4) );
  NAND2X4 U10 ( .A(n3), .B(n4), .Y(in_17bit_b[2]) );
  INVXL U11 ( .A(in_17bit[2]), .Y(n1) );
  INVX3 U12 ( .A(n53), .Y(n2) );
  NOR2X4 U13 ( .A(n33), .B(n28), .Y(n53) );
  NAND2XL U14 ( .A(n24), .B(n6), .Y(n7) );
  NAND2X1 U15 ( .A(n5), .B(in_17bit[3]), .Y(n8) );
  NAND2X2 U16 ( .A(n7), .B(n8), .Y(in_17bit_b[3]) );
  INVX1 U17 ( .A(n24), .Y(n5) );
  INVXL U18 ( .A(in_17bit[3]), .Y(n6) );
  NOR2X2 U19 ( .A(n32), .B(n55), .Y(n24) );
  NOR2X4 U20 ( .A(n15), .B(mul[20]), .Y(n116) );
  INVX4 U21 ( .A(in_17bit[16]), .Y(n33) );
  INVXL U22 ( .A(in_8bit[3]), .Y(n36) );
  XOR2X2 U23 ( .A(n35), .B(n38), .Y(in_8bit_b[2]) );
  INVX1 U24 ( .A(n23), .Y(n9) );
  INVX1 U25 ( .A(n54), .Y(n55) );
  XNOR2X1 U26 ( .A(n60), .B(n61), .Y(in_17bit_b[5]) );
  NOR2X1 U27 ( .A(mul[13]), .B(n95), .Y(n21) );
  INVX1 U28 ( .A(n102), .Y(n104) );
  NAND2BX1 U29 ( .AN(mul[16]), .B(n104), .Y(n105) );
  CLKINVX3 U30 ( .A(in_8bit[2]), .Y(n38) );
  NOR2X1 U31 ( .A(n23), .B(n25), .Y(n111) );
  NAND2BX2 U32 ( .AN(mul[17]), .B(n107), .Y(n108) );
  XOR2X2 U33 ( .A(mul[17]), .B(n106), .Y(out[10]) );
  NOR2X2 U34 ( .A(n23), .B(n107), .Y(n106) );
  CLKINVX3 U35 ( .A(n117), .Y(n120) );
  NOR2BX4 U36 ( .AN(n9), .B(n116), .Y(n115) );
  XNOR2X1 U37 ( .A(n125), .B(sub_add_52_b0_carry[14]), .Y(n10) );
  XNOR2X1 U38 ( .A(n124), .B(sub_add_52_b0_carry[13]), .Y(n11) );
  XNOR2X1 U39 ( .A(n126), .B(sub_add_52_b0_carry[15]), .Y(n12) );
  INVX1 U40 ( .A(n95), .Y(n97) );
  NAND2BX1 U41 ( .AN(mul[12]), .B(n94), .Y(n95) );
  OR2X2 U42 ( .A(n20), .B(n50), .Y(n13) );
  NAND2BX2 U43 ( .AN(mul[21]), .B(n116), .Y(n117) );
  CLKINVX3 U44 ( .A(n43), .Y(n46) );
  NOR2X4 U45 ( .A(in_17bit[1]), .B(in_17bit[0]), .Y(n28) );
  NOR3X1 U46 ( .A(n41), .B(in_8bit[1]), .C(n43), .Y(n42) );
  NAND2BX1 U47 ( .AN(in_17bit[2]), .B(n28), .Y(n54) );
  NOR2X1 U48 ( .A(in_17bit[16]), .B(in_17bit[1]), .Y(n51) );
  NAND3XL U49 ( .A(in_17bit[0]), .B(in_17bit[16]), .C(in_17bit[1]), .Y(n52) );
  INVX2 U50 ( .A(n44), .Y(n45) );
  XNOR2X4 U51 ( .A(n118), .B(n119), .Y(out[15]) );
  OAI21X4 U52 ( .A0(mul[19]), .A1(n114), .B0(n112), .Y(n113) );
  NOR2X4 U53 ( .A(n23), .B(n120), .Y(n118) );
  NOR2X1 U54 ( .A(n23), .B(n104), .Y(n103) );
  XNOR2X2 U55 ( .A(mul[20]), .B(n113), .Y(out[13]) );
  NAND2X1 U56 ( .A(n57), .B(in_17bit[16]), .Y(n56) );
  NOR2X2 U57 ( .A(mul[19]), .B(n114), .Y(n14) );
  INVX2 U58 ( .A(n14), .Y(n15) );
  OR2X2 U59 ( .A(in_8bit[4]), .B(in_8bit[3]), .Y(n43) );
  NAND2BX2 U60 ( .AN(n29), .B(n38), .Y(n44) );
  NAND2X1 U61 ( .A(n29), .B(in_8bit[7]), .Y(n34) );
  BUFX8 U62 ( .A(in_8bit[0]), .Y(n29) );
  INVX1 U63 ( .A(n37), .Y(n16) );
  CLKINVX3 U64 ( .A(n16), .Y(n17) );
  CLKINVX4 U65 ( .A(n13), .Y(n18) );
  NAND4BX2 U66 ( .AN(in_8bit[1]), .B(n31), .C(n46), .D(n45), .Y(n50) );
  XOR2X2 U67 ( .A(n111), .B(mul[19]), .Y(out[12]) );
  INVX2 U68 ( .A(mul[22]), .Y(n119) );
  NAND2BX1 U69 ( .AN(mul[14]), .B(n21), .Y(n99) );
  INVXL U70 ( .A(in_8bit[7]), .Y(n49) );
  XOR2X4 U71 ( .A(n27), .B(n31), .Y(in_8bit_b[5]) );
  OR2X2 U72 ( .A(n42), .B(n49), .Y(n27) );
  AND2X2 U73 ( .A(n59), .B(n58), .Y(n22) );
  NOR2XL U74 ( .A(in_8bit[6]), .B(n49), .Y(n19) );
  INVX1 U75 ( .A(n19), .Y(n20) );
  INVX4 U76 ( .A(n108), .Y(n110) );
  NAND2BXL U77 ( .AN(mul[10]), .B(n88), .Y(n89) );
  NAND2XL U78 ( .A(out[0]), .B(n112), .Y(n84) );
  AOI21XL U79 ( .A0(n120), .A1(n119), .B0(n23), .Y(n121) );
  NOR2XL U80 ( .A(n23), .B(n94), .Y(n93) );
  NOR2XL U81 ( .A(n23), .B(n101), .Y(n100) );
  NOR2XL U82 ( .A(n23), .B(n91), .Y(n90) );
  NOR2XL U83 ( .A(n23), .B(n26), .Y(n85) );
  OAI21XL U84 ( .A0(in_8bit[1]), .A1(n41), .B0(in_8bit[7]), .Y(n37) );
  INVXL U85 ( .A(in_8bit[5]), .Y(n31) );
  NAND2XL U86 ( .A(n63), .B(in_17bit[16]), .Y(n62) );
  NAND2XL U87 ( .A(n22), .B(n61), .Y(n63) );
  NOR2XL U88 ( .A(n33), .B(n68), .Y(n66) );
  NAND2XL U89 ( .A(n70), .B(in_17bit[16]), .Y(n69) );
  NAND2XL U90 ( .A(n68), .B(n67), .Y(n70) );
  NAND2BXL U91 ( .AN(n63), .B(n64), .Y(n65) );
  NAND2BXL U92 ( .AN(n70), .B(n71), .Y(n72) );
  INVXL U93 ( .A(n80), .Y(n81) );
  INVXL U94 ( .A(n83), .Y(sub_add_52_b0_carry[12]) );
  NAND2XL U95 ( .A(n75), .B(n74), .Y(n77) );
  XNOR2X1 U96 ( .A(in_17bit[16]), .B(in_8bit[7]), .Y(n23) );
  NAND2BXL U97 ( .AN(in_17bit[3]), .B(n55), .Y(n57) );
  INVX1 U98 ( .A(n89), .Y(n91) );
  INVX1 U99 ( .A(n86), .Y(n88) );
  NAND2BX1 U100 ( .AN(mul[9]), .B(n26), .Y(n86) );
  NOR2X1 U101 ( .A(mul[8]), .B(out[0]), .Y(n26) );
  XOR2X1 U102 ( .A(mul[23]), .B(n121), .Y(out[16]) );
  XNOR2X1 U103 ( .A(mul[8]), .B(n84), .Y(out[1]) );
  NAND2BX1 U104 ( .AN(mul[15]), .B(n101), .Y(n102) );
  INVX1 U105 ( .A(n99), .Y(n101) );
  INVX1 U106 ( .A(n92), .Y(n94) );
  NAND2BX1 U107 ( .AN(mul[11]), .B(n91), .Y(n92) );
  XOR2X1 U108 ( .A(mul[16]), .B(n103), .Y(out[9]) );
  XOR2X1 U109 ( .A(mul[15]), .B(n100), .Y(out[8]) );
  XOR2X1 U110 ( .A(mul[9]), .B(n85), .Y(out[2]) );
  XOR2X1 U111 ( .A(mul[10]), .B(n87), .Y(out[3]) );
  NOR2X1 U112 ( .A(n23), .B(n88), .Y(n87) );
  XOR2X1 U113 ( .A(mul[11]), .B(n90), .Y(out[4]) );
  XOR2X1 U114 ( .A(mul[12]), .B(n93), .Y(out[5]) );
  XOR2X1 U115 ( .A(mul[13]), .B(n96), .Y(out[6]) );
  NOR2X1 U116 ( .A(n23), .B(n97), .Y(n96) );
  INVX1 U117 ( .A(n23), .Y(n112) );
  INVX1 U118 ( .A(in_8bit[4]), .Y(n30) );
  NOR2X2 U119 ( .A(n39), .B(n49), .Y(n40) );
  XNOR2X1 U120 ( .A(in_8bit[1]), .B(n34), .Y(in_8bit_b[1]) );
  XNOR2X1 U121 ( .A(n66), .B(n67), .Y(in_17bit_b[7]) );
  XNOR2X1 U122 ( .A(n73), .B(n74), .Y(in_17bit_b[9]) );
  NOR2X1 U123 ( .A(n32), .B(n75), .Y(n73) );
  XOR2X1 U124 ( .A(n78), .B(n76), .Y(in_17bit_b[10]) );
  XOR2X1 U125 ( .A(n64), .B(n62), .Y(in_17bit_b[6]) );
  XOR2X1 U126 ( .A(n71), .B(n69), .Y(in_17bit_b[8]) );
  NOR2X1 U127 ( .A(n32), .B(n22), .Y(n60) );
  XOR2X1 U128 ( .A(n58), .B(n56), .Y(in_17bit_b[4]) );
  INVX1 U129 ( .A(n57), .Y(n59) );
  INVX1 U130 ( .A(n65), .Y(n68) );
  INVX1 U131 ( .A(n72), .Y(n75) );
  NAND2X1 U132 ( .A(n122), .B(n81), .Y(n83) );
  NAND2BX1 U133 ( .AN(n77), .B(n78), .Y(n80) );
  XOR2X1 U134 ( .A(n80), .B(n122), .Y(n79) );
  XOR2X1 U135 ( .A(n83), .B(n123), .Y(n82) );
  INVX1 U136 ( .A(in_17bit[5]), .Y(n61) );
  INVX1 U137 ( .A(in_17bit[4]), .Y(n58) );
  INVX1 U138 ( .A(in_17bit[16]), .Y(n32) );
  INVX1 U139 ( .A(in_17bit[7]), .Y(n67) );
  INVX1 U140 ( .A(in_17bit[9]), .Y(n74) );
  INVX1 U141 ( .A(in_17bit[6]), .Y(n64) );
  INVX1 U142 ( .A(in_17bit[8]), .Y(n71) );
  INVX1 U143 ( .A(in_17bit[10]), .Y(n78) );
  INVX1 U144 ( .A(in_17bit[11]), .Y(n122) );
  INVX1 U145 ( .A(in_17bit[12]), .Y(n123) );
  INVX1 U146 ( .A(in_17bit[13]), .Y(n124) );
  INVX1 U147 ( .A(in_17bit[14]), .Y(n125) );
  INVX1 U148 ( .A(in_17bit[15]), .Y(n126) );
  INVX1 U149 ( .A(in_8bit[6]), .Y(n47) );
  AND2X1 U150 ( .A(N21), .B(in_17bit[16]), .Y(in_17bit_b[16]) );
  MXI2XL U151 ( .A(n126), .B(n12), .S0(in_17bit[16]), .Y(in_17bit_b[15]) );
  MXI2XL U152 ( .A(n125), .B(n10), .S0(in_17bit[16]), .Y(in_17bit_b[14]) );
  MXI2XL U153 ( .A(n124), .B(n11), .S0(in_17bit[16]), .Y(in_17bit_b[13]) );
  MXI2XL U154 ( .A(n123), .B(n82), .S0(in_17bit[16]), .Y(in_17bit_b[12]) );
  MXI2XL U155 ( .A(n122), .B(n79), .S0(in_17bit[16]), .Y(in_17bit_b[11]) );
  NAND2XL U156 ( .A(n77), .B(in_17bit[16]), .Y(n76) );
  NAND2X2 U157 ( .A(n50), .B(in_8bit[7]), .Y(n48) );
  XOR2X4 U158 ( .A(n17), .B(n36), .Y(in_8bit_b[3]) );
  XNOR2X4 U159 ( .A(n40), .B(n30), .Y(in_8bit_b[4]) );
  XOR2X4 U160 ( .A(n48), .B(n47), .Y(in_8bit_b[6]) );
  NOR3BX4 U161 ( .AN(n52), .B(n28), .C(n51), .Y(in_17bit_b[1]) );
  NOR2X4 U162 ( .A(n23), .B(n21), .Y(n98) );
  XOR2X4 U163 ( .A(mul[14]), .B(n98), .Y(out[7]) );
  NOR2X4 U164 ( .A(n23), .B(n110), .Y(n109) );
  XOR2X4 U165 ( .A(mul[18]), .B(n109), .Y(out[11]) );
  XOR2X4 U166 ( .A(mul[21]), .B(n115), .Y(out[14]) );
  XOR2X1 U167 ( .A(n32), .B(sub_add_52_b0_carry[16]), .Y(N21) );
  AND2X1 U168 ( .A(sub_add_52_b0_carry[15]), .B(n126), .Y(
        sub_add_52_b0_carry[16]) );
  AND2X1 U169 ( .A(sub_add_52_b0_carry[14]), .B(n125), .Y(
        sub_add_52_b0_carry[15]) );
  AND2X1 U170 ( .A(sub_add_52_b0_carry[13]), .B(n124), .Y(
        sub_add_52_b0_carry[14]) );
  AND2X1 U171 ( .A(sub_add_52_b0_carry[12]), .B(n123), .Y(
        sub_add_52_b0_carry[13]) );
endmodule


module multi16_1_DW01_add_0 ( A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, 
        A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, 
        B_20_, B_19_, B_18_, B_17_, B_16_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, 
        SUM_17_, SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, 
        SUM_9_, SUM_8_, SUM_7_, SUM_6_, SUM_5_ );
  input A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_,
         A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, B_20_, B_19_,
         B_18_, B_17_, B_16_;
  output SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, SUM_15_,
         SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, SUM_7_,
         SUM_6_, SUM_5_;
  wire   n1, n2, n3, n5, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39;

  NAND2X2 U2 ( .A(n33), .B(n17), .Y(n39) );
  OAI21X1 U3 ( .A0(n38), .A1(n31), .B0(n33), .Y(n36) );
  NOR2X2 U4 ( .A(B_18_), .B(A_18_), .Y(n31) );
  BUFX3 U5 ( .A(A_12_), .Y(SUM_12_) );
  BUFX3 U6 ( .A(A_14_), .Y(SUM_14_) );
  CLKINVX3 U7 ( .A(n21), .Y(SUM_15_) );
  INVX1 U8 ( .A(A_15_), .Y(n21) );
  INVX2 U9 ( .A(n35), .Y(n19) );
  OAI21X1 U10 ( .A0(n27), .A1(n28), .B0(n29), .Y(n24) );
  AOI21XL U11 ( .A0(n17), .A1(n32), .B0(n18), .Y(n27) );
  INVX2 U12 ( .A(n30), .Y(n20) );
  AND2X4 U13 ( .A(B_16_), .B(A_16_), .Y(n1) );
  NAND2X2 U14 ( .A(B_17_), .B(A_17_), .Y(n35) );
  NOR2X2 U15 ( .A(B_17_), .B(A_17_), .Y(n30) );
  XOR2X2 U16 ( .A(n36), .B(n37), .Y(SUM_19_) );
  NOR2BX4 U17 ( .AN(n34), .B(n5), .Y(SUM_16_) );
  NOR2BX2 U18 ( .AN(n29), .B(n28), .Y(n37) );
  AOI21X2 U19 ( .A0(n1), .A1(n20), .B0(n19), .Y(n38) );
  NOR2X2 U20 ( .A(n30), .B(n19), .Y(n2) );
  XOR2X4 U21 ( .A(n1), .B(n2), .Y(SUM_17_) );
  XOR2X1 U22 ( .A(n3), .B(n24), .Y(SUM_20_) );
  INVXL U23 ( .A(n26), .Y(n16) );
  AOI21XL U24 ( .A0(n24), .A1(n25), .B0(n16), .Y(n23) );
  BUFX3 U25 ( .A(A_11_), .Y(SUM_11_) );
  INVXL U26 ( .A(n33), .Y(n18) );
  INVX1 U27 ( .A(n31), .Y(n17) );
  AND2X2 U28 ( .A(n26), .B(n25), .Y(n3) );
  NOR2X1 U29 ( .A(B_16_), .B(A_16_), .Y(n5) );
  BUFX3 U30 ( .A(A_5_), .Y(SUM_5_) );
  BUFX3 U31 ( .A(A_6_), .Y(SUM_6_) );
  BUFX3 U32 ( .A(A_7_), .Y(SUM_7_) );
  BUFX3 U33 ( .A(A_8_), .Y(SUM_8_) );
  BUFX3 U34 ( .A(A_9_), .Y(SUM_9_) );
  BUFX8 U35 ( .A(A_13_), .Y(SUM_13_) );
  BUFX3 U36 ( .A(A_10_), .Y(SUM_10_) );
  XOR2X2 U37 ( .A(n39), .B(n38), .Y(SUM_18_) );
  XOR2X1 U38 ( .A(n22), .B(n23), .Y(SUM_21_) );
  XNOR2X1 U39 ( .A(B_21_), .B(A_21_), .Y(n22) );
  OAI21XL U40 ( .A0(n30), .A1(n34), .B0(n35), .Y(n32) );
  OR2X1 U41 ( .A(B_20_), .B(A_20_), .Y(n25) );
  NAND2X1 U42 ( .A(B_20_), .B(A_20_), .Y(n26) );
  NOR2X1 U43 ( .A(B_19_), .B(A_19_), .Y(n28) );
  NAND2X1 U44 ( .A(B_19_), .B(A_19_), .Y(n29) );
  NAND2X1 U45 ( .A(B_18_), .B(A_18_), .Y(n33) );
  NAND2X1 U46 ( .A(B_16_), .B(A_16_), .Y(n34) );
endmodule


module multi16_1_DW02_mult_0 ( A, B, PRODUCT_23_, PRODUCT_22_, PRODUCT_21_, 
        PRODUCT_20_, PRODUCT_19_, PRODUCT_18_, PRODUCT_17_, PRODUCT_16_, 
        PRODUCT_15_, PRODUCT_14_, PRODUCT_13_, PRODUCT_12_, PRODUCT_11_, 
        PRODUCT_10_, PRODUCT_9_, PRODUCT_8_, PRODUCT_7_ );
  input [16:0] A;
  input [7:0] B;
  output PRODUCT_23_, PRODUCT_22_, PRODUCT_21_, PRODUCT_20_, PRODUCT_19_,
         PRODUCT_18_, PRODUCT_17_, PRODUCT_16_, PRODUCT_15_, PRODUCT_14_,
         PRODUCT_13_, PRODUCT_12_, PRODUCT_11_, PRODUCT_10_, PRODUCT_9_,
         PRODUCT_8_, PRODUCT_7_;
  wire   ab_16__7_, ab_16__6_, ab_16__5_, ab_16__4_, ab_16__3_, ab_16__2_,
         ab_16__1_, ab_16__0_, ab_15__7_, ab_15__6_, ab_15__5_, ab_15__4_,
         ab_15__3_, ab_15__2_, ab_15__1_, ab_15__0_, ab_14__7_, ab_14__6_,
         ab_14__5_, ab_14__4_, ab_14__3_, ab_14__2_, ab_14__1_, ab_14__0_,
         ab_13__7_, ab_13__6_, ab_13__5_, ab_13__4_, ab_13__3_, ab_13__2_,
         ab_13__1_, ab_13__0_, ab_12__7_, ab_12__6_, ab_12__5_, ab_12__4_,
         ab_12__3_, ab_12__2_, ab_12__1_, ab_12__0_, ab_11__7_, ab_11__6_,
         ab_11__5_, ab_11__4_, ab_11__3_, ab_11__2_, ab_11__1_, ab_11__0_,
         ab_10__7_, ab_10__6_, ab_10__5_, ab_10__4_, ab_10__3_, ab_10__2_,
         ab_10__1_, ab_10__0_, ab_9__7_, ab_9__6_, ab_9__5_, ab_9__4_,
         ab_9__3_, ab_9__2_, ab_9__1_, ab_9__0_, ab_8__7_, ab_8__6_, ab_8__5_,
         ab_8__4_, ab_8__3_, ab_8__2_, ab_8__1_, ab_8__0_, ab_7__7_, ab_7__6_,
         ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_, ab_7__0_, ab_6__7_,
         ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_, ab_6__1_, ab_6__0_,
         ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_, ab_5__2_, ab_5__1_,
         ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_, ab_4__3_, ab_4__2_,
         ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_, ab_3__4_, ab_3__3_,
         ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_, ab_2__5_, ab_2__4_,
         ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_, ab_1__6_, ab_1__5_,
         ab_1__4_, ab_1__3_, ab_1__2_, ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_,
         ab_0__3_, ab_0__2_, CARRYB_16__6_, CARRYB_16__5_, CARRYB_16__4_,
         CARRYB_16__3_, CARRYB_16__2_, CARRYB_16__1_, CARRYB_16__0_,
         CARRYB_15__6_, CARRYB_15__5_, CARRYB_15__4_, CARRYB_15__3_,
         CARRYB_15__2_, CARRYB_15__1_, CARRYB_15__0_, CARRYB_14__6_,
         CARRYB_14__5_, CARRYB_14__4_, CARRYB_14__3_, CARRYB_14__2_,
         CARRYB_14__1_, CARRYB_14__0_, CARRYB_13__6_, CARRYB_13__5_,
         CARRYB_13__4_, CARRYB_13__3_, CARRYB_13__2_, CARRYB_13__1_,
         CARRYB_13__0_, CARRYB_12__6_, CARRYB_12__5_, CARRYB_12__4_,
         CARRYB_12__3_, CARRYB_12__2_, CARRYB_12__1_, CARRYB_12__0_,
         CARRYB_11__6_, CARRYB_11__5_, CARRYB_11__4_, CARRYB_11__3_,
         CARRYB_11__2_, CARRYB_11__1_, CARRYB_11__0_, CARRYB_10__6_,
         CARRYB_10__5_, CARRYB_10__4_, CARRYB_10__3_, CARRYB_10__2_,
         CARRYB_10__1_, CARRYB_10__0_, CARRYB_9__6_, CARRYB_9__5_,
         CARRYB_9__4_, CARRYB_9__3_, CARRYB_9__2_, CARRYB_9__1_, CARRYB_9__0_,
         CARRYB_8__6_, CARRYB_8__5_, CARRYB_8__4_, CARRYB_8__3_, CARRYB_8__2_,
         CARRYB_8__1_, CARRYB_8__0_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_,
         CARRYB_7__3_, CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_,
         CARRYB_6__5_, CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_,
         CARRYB_6__0_, CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_,
         CARRYB_5__2_, CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_,
         CARRYB_4__4_, CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_,
         CARRYB_3__6_, CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_,
         CARRYB_3__1_, CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_,
         CARRYB_2__3_, CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__0_,
         SUMB_16__6_, SUMB_16__5_, SUMB_16__4_, SUMB_16__3_, SUMB_16__2_,
         SUMB_16__1_, SUMB_16__0_, SUMB_15__6_, SUMB_15__5_, SUMB_15__4_,
         SUMB_15__3_, SUMB_15__2_, SUMB_15__1_, SUMB_14__6_, SUMB_14__5_,
         SUMB_14__4_, SUMB_14__3_, SUMB_14__2_, SUMB_14__1_, SUMB_13__6_,
         SUMB_13__5_, SUMB_13__4_, SUMB_13__3_, SUMB_13__2_, SUMB_13__1_,
         SUMB_12__6_, SUMB_12__5_, SUMB_12__4_, SUMB_12__3_, SUMB_12__2_,
         SUMB_12__1_, SUMB_11__6_, SUMB_11__5_, SUMB_11__4_, SUMB_11__3_,
         SUMB_11__2_, SUMB_11__1_, SUMB_10__6_, SUMB_10__5_, SUMB_10__4_,
         SUMB_10__3_, SUMB_10__2_, SUMB_10__1_, SUMB_9__6_, SUMB_9__5_,
         SUMB_9__4_, SUMB_9__3_, SUMB_9__2_, SUMB_9__1_, SUMB_8__6_,
         SUMB_8__5_, SUMB_8__4_, SUMB_8__3_, SUMB_8__2_, SUMB_8__1_,
         SUMB_7__6_, SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_,
         SUMB_7__1_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, PROD1_7_, A1_21_, A1_20_, A1_19_, A1_18_,
         A1_17_, A1_16_, A1_15_, A1_13_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_,
         A1_7_, A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41;

  ADDFHX4 S1_14_0 ( .A(ab_14__0_), .B(CARRYB_13__0_), .CI(SUMB_13__1_), .CO(
        CARRYB_14__0_), .S(A1_12_) );
  ADDFHX4 S1_13_0 ( .A(ab_13__0_), .B(CARRYB_12__0_), .CI(SUMB_12__1_), .CO(
        CARRYB_13__0_), .S(A1_11_) );
  ADDFHX4 S2_13_1 ( .A(ab_13__1_), .B(CARRYB_12__1_), .CI(SUMB_12__2_), .CO(
        CARRYB_13__1_), .S(SUMB_13__1_) );
  ADDFHX4 S2_12_2 ( .A(ab_12__2_), .B(CARRYB_11__2_), .CI(SUMB_11__3_), .CO(
        CARRYB_12__2_), .S(SUMB_12__2_) );
  ADDFHX4 S1_11_0 ( .A(ab_11__0_), .B(CARRYB_10__0_), .CI(SUMB_10__1_), .CO(
        CARRYB_11__0_), .S(A1_9_) );
  ADDFHX4 S2_11_2 ( .A(ab_11__2_), .B(CARRYB_10__2_), .CI(SUMB_10__3_), .CO(
        CARRYB_11__2_), .S(SUMB_11__2_) );
  ADDFHX4 S2_10_2 ( .A(ab_10__2_), .B(CARRYB_9__2_), .CI(SUMB_9__3_), .CO(
        CARRYB_10__2_), .S(SUMB_10__2_) );
  multi16_1_DW01_add_0 FS_1 ( .A_21_(A1_21_), .A_20_(A1_20_), .A_19_(A1_19_), 
        .A_18_(A1_18_), .A_17_(A1_17_), .A_16_(A1_16_), .A_15_(A1_15_), 
        .A_14_(SUMB_16__0_), .A_13_(A1_13_), .A_12_(A1_12_), .A_11_(A1_11_), 
        .A_10_(A1_10_), .A_9_(A1_9_), .A_8_(A1_8_), .A_7_(A1_7_), .A_6_(A1_6_), 
        .A_5_(PROD1_7_), .B_21_(n10), .B_20_(n22), .B_19_(n20), .B_18_(n19), 
        .B_17_(n18), .B_16_(n21), .SUM_21_(PRODUCT_23_), .SUM_20_(PRODUCT_22_), 
        .SUM_19_(PRODUCT_21_), .SUM_18_(PRODUCT_20_), .SUM_17_(PRODUCT_19_), 
        .SUM_16_(PRODUCT_18_), .SUM_15_(PRODUCT_17_), .SUM_14_(PRODUCT_16_), 
        .SUM_13_(PRODUCT_15_), .SUM_12_(PRODUCT_14_), .SUM_11_(PRODUCT_13_), 
        .SUM_10_(PRODUCT_12_), .SUM_9_(PRODUCT_11_), .SUM_8_(PRODUCT_10_), 
        .SUM_7_(PRODUCT_9_), .SUM_6_(PRODUCT_8_), .SUM_5_(PRODUCT_7_) );
  ADDFHX1 S2_15_5 ( .A(ab_15__5_), .B(CARRYB_14__5_), .CI(SUMB_14__6_), .CO(
        CARRYB_15__5_), .S(SUMB_15__5_) );
  ADDFX2 S3_15_6 ( .A(ab_15__6_), .B(CARRYB_14__6_), .CI(ab_14__7_), .CO(
        CARRYB_15__6_), .S(SUMB_15__6_) );
  ADDFHX1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  ADDFHX1 S5_6 ( .A(ab_16__6_), .B(CARRYB_15__6_), .CI(ab_15__7_), .CO(
        CARRYB_16__6_), .S(SUMB_16__6_) );
  ADDFHX2 S2_9_3 ( .A(ab_9__3_), .B(CARRYB_8__3_), .CI(SUMB_8__4_), .CO(
        CARRYB_9__3_), .S(SUMB_9__3_) );
  ADDFHX2 S2_7_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  ADDFHX4 S2_11_5 ( .A(ab_11__5_), .B(CARRYB_10__5_), .CI(SUMB_10__6_), .CO(
        CARRYB_11__5_), .S(SUMB_11__5_) );
  ADDFHX4 S1_8_0 ( .A(ab_8__0_), .B(CARRYB_7__0_), .CI(SUMB_7__1_), .CO(
        CARRYB_8__0_), .S(A1_6_) );
  ADDFHX2 S2_2_1 ( .A(ab_2__1_), .B(n6), .CI(SUMB_1__2_), .CO(CARRYB_2__1_), 
        .S(SUMB_2__1_) );
  ADDFHX4 S2_7_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  ADDFHX4 S2_8_4 ( .A(ab_8__4_), .B(CARRYB_7__4_), .CI(SUMB_7__5_), .CO(
        CARRYB_8__4_), .S(SUMB_8__4_) );
  ADDFHX2 S3_11_6 ( .A(ab_11__6_), .B(CARRYB_10__6_), .CI(ab_10__7_), .CO(
        CARRYB_11__6_), .S(SUMB_11__6_) );
  ADDFHX4 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  ADDFHX4 S3_8_6 ( .A(ab_8__6_), .B(CARRYB_7__6_), .CI(ab_7__7_), .CO(
        CARRYB_8__6_), .S(SUMB_8__6_) );
  ADDFHX4 S2_7_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  ADDFHX4 S2_13_2 ( .A(ab_13__2_), .B(CARRYB_12__2_), .CI(SUMB_12__3_), .CO(
        CARRYB_13__2_), .S(SUMB_13__2_) );
  ADDFHX4 S2_14_2 ( .A(ab_14__2_), .B(CARRYB_13__2_), .CI(SUMB_13__3_), .CO(
        CARRYB_14__2_), .S(SUMB_14__2_) );
  ADDFHX2 S4_2 ( .A(ab_16__2_), .B(CARRYB_15__2_), .CI(SUMB_15__3_), .CO(
        CARRYB_16__2_), .S(SUMB_16__2_) );
  ADDFHX2 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  ADDFHX2 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  ADDFHX2 S2_14_5 ( .A(ab_14__5_), .B(CARRYB_13__5_), .CI(SUMB_13__6_), .CO(
        CARRYB_14__5_), .S(SUMB_14__5_) );
  ADDFHX2 S2_13_5 ( .A(ab_13__5_), .B(CARRYB_12__5_), .CI(SUMB_12__6_), .CO(
        CARRYB_13__5_), .S(SUMB_13__5_) );
  ADDFHX4 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  ADDFHX4 S2_8_1 ( .A(ab_8__1_), .B(CARRYB_7__1_), .CI(SUMB_7__2_), .CO(
        CARRYB_8__1_), .S(SUMB_8__1_) );
  ADDFHX4 S2_14_4 ( .A(ab_14__4_), .B(CARRYB_13__4_), .CI(SUMB_13__5_), .CO(
        CARRYB_14__4_), .S(SUMB_14__4_) );
  ADDFHX4 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  ADDFHX2 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  ADDFHX2 S3_2_6 ( .A(ab_2__6_), .B(n9), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  ADDFHX2 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  ADDFHX2 S3_13_6 ( .A(ab_13__6_), .B(CARRYB_12__6_), .CI(ab_12__7_), .CO(
        CARRYB_13__6_), .S(SUMB_13__6_) );
  ADDFHX2 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  ADDFHX2 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  ADDFHX2 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  ADDFHX2 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  ADDFHX4 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  ADDFHX4 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  ADDFHX4 S1_10_0 ( .A(ab_10__0_), .B(CARRYB_9__0_), .CI(SUMB_9__1_), .CO(
        CARRYB_10__0_), .S(A1_8_) );
  ADDFHX4 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  ADDFHX4 S2_10_5 ( .A(ab_10__5_), .B(CARRYB_9__5_), .CI(SUMB_9__6_), .CO(
        CARRYB_10__5_), .S(SUMB_10__5_) );
  ADDFHX4 S2_11_3 ( .A(ab_11__3_), .B(CARRYB_10__3_), .CI(SUMB_10__4_), .CO(
        CARRYB_11__3_), .S(SUMB_11__3_) );
  ADDFHX4 S2_12_3 ( .A(ab_12__3_), .B(CARRYB_11__3_), .CI(SUMB_11__4_), .CO(
        CARRYB_12__3_), .S(SUMB_12__3_) );
  ADDFHX4 S4_3 ( .A(ab_16__3_), .B(CARRYB_15__3_), .CI(SUMB_15__4_), .CO(
        CARRYB_16__3_), .S(SUMB_16__3_) );
  ADDFHX4 S2_11_4 ( .A(ab_11__4_), .B(CARRYB_10__4_), .CI(SUMB_10__5_), .CO(
        CARRYB_11__4_), .S(SUMB_11__4_) );
  ADDFHX2 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  ADDFHX2 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  ADDFHX4 S2_9_2 ( .A(ab_9__2_), .B(CARRYB_8__2_), .CI(SUMB_8__3_), .CO(
        CARRYB_9__2_), .S(SUMB_9__2_) );
  ADDFHX4 S2_13_3 ( .A(ab_13__3_), .B(CARRYB_12__3_), .CI(SUMB_12__4_), .CO(
        CARRYB_13__3_), .S(SUMB_13__3_) );
  ADDFHX4 S2_15_3 ( .A(ab_15__3_), .B(CARRYB_14__3_), .CI(SUMB_14__4_), .CO(
        CARRYB_15__3_), .S(SUMB_15__3_) );
  ADDFHX2 S2_15_4 ( .A(ab_15__4_), .B(CARRYB_14__4_), .CI(SUMB_14__5_), .CO(
        CARRYB_15__4_), .S(SUMB_15__4_) );
  ADDFHX2 S2_2_3 ( .A(ab_2__3_), .B(n7), .CI(SUMB_1__4_), .CO(CARRYB_2__3_), 
        .S(SUMB_2__3_) );
  ADDFHX4 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  ADDFHX4 S2_14_3 ( .A(ab_14__3_), .B(CARRYB_13__3_), .CI(SUMB_13__4_), .CO(
        CARRYB_14__3_), .S(SUMB_14__3_) );
  ADDFHX2 S2_2_2 ( .A(ab_2__2_), .B(n4), .CI(SUMB_1__3_), .CO(CARRYB_2__2_), 
        .S(SUMB_2__2_) );
  ADDFHX4 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  ADDFHX1 S3_14_6 ( .A(ab_14__6_), .B(CARRYB_13__6_), .CI(ab_13__7_), .CO(
        CARRYB_14__6_), .S(SUMB_14__6_) );
  ADDFX2 S4_5 ( .A(ab_16__5_), .B(CARRYB_15__5_), .CI(SUMB_15__6_), .CO(
        CARRYB_16__5_), .S(SUMB_16__5_) );
  ADDFHX2 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  ADDFHX2 S3_10_6 ( .A(ab_10__6_), .B(CARRYB_9__6_), .CI(ab_9__7_), .CO(
        CARRYB_10__6_), .S(SUMB_10__6_) );
  ADDFX2 S4_4 ( .A(ab_16__4_), .B(CARRYB_15__4_), .CI(SUMB_15__5_), .CO(
        CARRYB_16__4_), .S(SUMB_16__4_) );
  ADDFHX2 S2_9_1 ( .A(ab_9__1_), .B(CARRYB_8__1_), .CI(SUMB_8__2_), .CO(
        CARRYB_9__1_), .S(SUMB_9__1_) );
  ADDFHX2 S3_7_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(
        CARRYB_7__6_), .S(SUMB_7__6_) );
  ADDFHX2 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  ADDFHX2 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  ADDFHX2 S1_15_0 ( .A(ab_15__0_), .B(CARRYB_14__0_), .CI(SUMB_14__1_), .CO(
        CARRYB_15__0_), .S(A1_13_) );
  ADDFHX2 S2_7_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  ADDFHX2 S3_9_6 ( .A(ab_9__6_), .B(CARRYB_8__6_), .CI(ab_8__7_), .CO(
        CARRYB_9__6_), .S(SUMB_9__6_) );
  ADDFHX2 S2_10_1 ( .A(ab_10__1_), .B(CARRYB_9__1_), .CI(SUMB_9__2_), .CO(
        CARRYB_10__1_), .S(SUMB_10__1_) );
  ADDFHX4 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  ADDFHX4 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  ADDFHX4 S2_2_4 ( .A(ab_2__4_), .B(n8), .CI(SUMB_1__5_), .CO(CARRYB_2__4_), 
        .S(SUMB_2__4_) );
  ADDFHX4 S2_2_5 ( .A(ab_2__5_), .B(n5), .CI(SUMB_1__6_), .CO(CARRYB_2__5_), 
        .S(SUMB_2__5_) );
  ADDFHX4 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  ADDFHX4 S2_12_1 ( .A(ab_12__1_), .B(CARRYB_11__1_), .CI(SUMB_11__2_), .CO(
        CARRYB_12__1_), .S(SUMB_12__1_) );
  ADDFHX4 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  ADDFHX4 S2_14_1 ( .A(ab_14__1_), .B(CARRYB_13__1_), .CI(SUMB_13__2_), .CO(
        CARRYB_14__1_), .S(SUMB_14__1_) );
  ADDFHX4 S2_15_1 ( .A(ab_15__1_), .B(CARRYB_14__1_), .CI(SUMB_14__2_), .CO(
        CARRYB_15__1_), .S(SUMB_15__1_) );
  ADDFHX2 S4_1 ( .A(ab_16__1_), .B(CARRYB_15__1_), .CI(SUMB_15__2_), .CO(
        CARRYB_16__1_), .S(SUMB_16__1_) );
  ADDFHX4 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  ADDFHX4 S1_7_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(PROD1_7_) );
  ADDFHX4 S1_9_0 ( .A(ab_9__0_), .B(CARRYB_8__0_), .CI(SUMB_8__1_), .CO(
        CARRYB_9__0_), .S(A1_7_) );
  ADDFHX4 S1_12_0 ( .A(ab_12__0_), .B(CARRYB_11__0_), .CI(SUMB_11__1_), .CO(
        CARRYB_12__0_), .S(A1_10_) );
  ADDFHX4 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  ADDFHX4 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  ADDFHX4 S2_9_4 ( .A(ab_9__4_), .B(CARRYB_8__4_), .CI(SUMB_8__5_), .CO(
        CARRYB_9__4_), .S(SUMB_9__4_) );
  ADDFHX4 S2_12_4 ( .A(ab_12__4_), .B(CARRYB_11__4_), .CI(SUMB_11__5_), .CO(
        CARRYB_12__4_), .S(SUMB_12__4_) );
  ADDFHX4 S2_11_1 ( .A(ab_11__1_), .B(CARRYB_10__1_), .CI(SUMB_10__2_), .CO(
        CARRYB_11__1_), .S(SUMB_11__1_) );
  ADDFHX4 S2_8_5 ( .A(ab_8__5_), .B(CARRYB_7__5_), .CI(SUMB_7__6_), .CO(
        CARRYB_8__5_), .S(SUMB_8__5_) );
  ADDFHX4 S2_9_5 ( .A(ab_9__5_), .B(CARRYB_8__5_), .CI(SUMB_8__6_), .CO(
        CARRYB_9__5_), .S(SUMB_9__5_) );
  ADDFHX2 S3_12_6 ( .A(ab_12__6_), .B(CARRYB_11__6_), .CI(ab_11__7_), .CO(
        CARRYB_12__6_), .S(SUMB_12__6_) );
  ADDFHX4 S2_7_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  ADDFHX4 S2_8_2 ( .A(ab_8__2_), .B(CARRYB_7__2_), .CI(SUMB_7__3_), .CO(
        CARRYB_8__2_), .S(SUMB_8__2_) );
  ADDFHX4 S2_15_2 ( .A(ab_15__2_), .B(CARRYB_14__2_), .CI(SUMB_14__3_), .CO(
        CARRYB_15__2_), .S(SUMB_15__2_) );
  ADDFHX2 S2_12_5 ( .A(ab_12__5_), .B(CARRYB_11__5_), .CI(SUMB_11__6_), .CO(
        CARRYB_12__5_), .S(SUMB_12__5_) );
  ADDFHX4 S2_13_4 ( .A(ab_13__4_), .B(CARRYB_12__4_), .CI(SUMB_12__5_), .CO(
        CARRYB_13__4_), .S(SUMB_13__4_) );
  ADDFHX4 S2_10_4 ( .A(ab_10__4_), .B(CARRYB_9__4_), .CI(SUMB_9__5_), .CO(
        CARRYB_10__4_), .S(SUMB_10__4_) );
  ADDFXL S4_0 ( .A(ab_16__0_), .B(CARRYB_15__0_), .CI(SUMB_15__1_), .CO(
        CARRYB_16__0_), .S(SUMB_16__0_) );
  AND2X2 U2 ( .A(A[1]), .B(B[2]), .Y(ab_1__2_) );
  AND2XL U3 ( .A(A[1]), .B(B[5]), .Y(ab_1__5_) );
  XOR2X2 U4 ( .A(CARRYB_16__3_), .B(SUMB_16__4_), .Y(A1_18_) );
  XOR2X2 U5 ( .A(ab_1__2_), .B(ab_0__3_), .Y(SUMB_1__2_) );
  INVX1 U6 ( .A(A[0]), .Y(n26) );
  NOR2X2 U7 ( .A(n29), .B(n26), .Y(ab_0__6_) );
  NOR2X2 U8 ( .A(n33), .B(n26), .Y(ab_0__2_) );
  BUFX3 U9 ( .A(B[7]), .Y(n23) );
  INVX1 U10 ( .A(B[2]), .Y(n33) );
  XOR2X1 U11 ( .A(ab_1__5_), .B(ab_0__6_), .Y(SUMB_1__5_) );
  XOR2X1 U12 ( .A(CARRYB_16__0_), .B(SUMB_16__1_), .Y(A1_15_) );
  CLKINVX3 U13 ( .A(B[6]), .Y(n29) );
  CLKINVX3 U14 ( .A(n23), .Y(n35) );
  AND2X2 U16 ( .A(ab_0__3_), .B(ab_1__2_), .Y(n4) );
  AND2X2 U17 ( .A(ab_0__6_), .B(ab_1__5_), .Y(n5) );
  AND2X2 U18 ( .A(ab_0__2_), .B(n36), .Y(n6) );
  AND2X2 U19 ( .A(ab_0__4_), .B(ab_1__3_), .Y(n7) );
  AND2X2 U20 ( .A(ab_0__5_), .B(ab_1__4_), .Y(n8) );
  AND2X2 U21 ( .A(ab_0__7_), .B(ab_1__6_), .Y(n9) );
  AND2X2 U22 ( .A(CARRYB_16__5_), .B(SUMB_16__6_), .Y(n10) );
  AND2X2 U23 ( .A(A[2]), .B(B[4]), .Y(ab_2__4_) );
  NAND2X2 U24 ( .A(ab_8__3_), .B(CARRYB_7__3_), .Y(n14) );
  AND2X2 U25 ( .A(A[1]), .B(B[4]), .Y(ab_1__4_) );
  XOR2X4 U26 ( .A(CARRYB_16__2_), .B(SUMB_16__3_), .Y(A1_17_) );
  XOR2X2 U27 ( .A(SUMB_7__4_), .B(n11), .Y(SUMB_8__3_) );
  AND2X2 U28 ( .A(A[1]), .B(B[3]), .Y(ab_1__3_) );
  AND2X2 U29 ( .A(CARRYB_16__1_), .B(SUMB_16__2_), .Y(n18) );
  AND2X2 U30 ( .A(CARRYB_16__0_), .B(SUMB_16__1_), .Y(n21) );
  NOR2X2 U31 ( .A(n32), .B(n26), .Y(ab_0__3_) );
  NOR2X2 U32 ( .A(n31), .B(n26), .Y(ab_0__4_) );
  INVX2 U33 ( .A(B[4]), .Y(n31) );
  NOR2X2 U34 ( .A(n35), .B(n26), .Y(ab_0__7_) );
  INVX2 U35 ( .A(B[3]), .Y(n32) );
  XOR2X4 U36 ( .A(CARRYB_7__3_), .B(ab_8__3_), .Y(n11) );
  NAND2X2 U37 ( .A(CARRYB_7__3_), .B(SUMB_7__4_), .Y(n12) );
  NAND2X2 U38 ( .A(ab_8__3_), .B(SUMB_7__4_), .Y(n13) );
  NAND3X4 U39 ( .A(n14), .B(n12), .C(n13), .Y(CARRYB_8__3_) );
  XOR3X2 U40 ( .A(CARRYB_9__3_), .B(ab_10__3_), .C(SUMB_9__4_), .Y(SUMB_10__3_) );
  NAND2XL U41 ( .A(SUMB_9__4_), .B(CARRYB_9__3_), .Y(n15) );
  NAND2XL U42 ( .A(ab_10__3_), .B(CARRYB_9__3_), .Y(n16) );
  NAND2XL U43 ( .A(ab_10__3_), .B(SUMB_9__4_), .Y(n17) );
  NAND3X2 U44 ( .A(n17), .B(n15), .C(n16), .Y(CARRYB_10__3_) );
  NOR2XL U45 ( .A(n38), .B(n29), .Y(ab_15__6_) );
  NOR2XL U46 ( .A(n40), .B(n29), .Y(ab_13__6_) );
  INVX4 U47 ( .A(n25), .Y(n24) );
  XOR2X2 U48 ( .A(CARRYB_16__1_), .B(SUMB_16__2_), .Y(A1_16_) );
  XOR2X1 U49 ( .A(ab_1__3_), .B(ab_0__4_), .Y(SUMB_1__3_) );
  INVX2 U50 ( .A(B[5]), .Y(n30) );
  AND2X1 U51 ( .A(CARRYB_16__3_), .B(SUMB_16__4_), .Y(n20) );
  AND2X1 U52 ( .A(A[6]), .B(B[2]), .Y(ab_6__2_) );
  AND2X1 U53 ( .A(A[9]), .B(B[1]), .Y(ab_9__1_) );
  AND2X1 U54 ( .A(A[7]), .B(B[2]), .Y(ab_7__2_) );
  AND2X1 U55 ( .A(A[11]), .B(B[2]), .Y(ab_11__2_) );
  AND2X1 U56 ( .A(A[11]), .B(B[1]), .Y(ab_11__1_) );
  AND2X1 U57 ( .A(A[10]), .B(B[2]), .Y(ab_10__2_) );
  AND2X1 U58 ( .A(A[9]), .B(B[2]), .Y(ab_9__2_) );
  AND2X1 U59 ( .A(A[10]), .B(B[1]), .Y(ab_10__1_) );
  AND2X1 U60 ( .A(A[8]), .B(B[2]), .Y(ab_8__2_) );
  AND2X1 U61 ( .A(A[7]), .B(B[1]), .Y(ab_7__1_) );
  AND2X1 U62 ( .A(A[5]), .B(B[2]), .Y(ab_5__2_) );
  AND2X1 U63 ( .A(A[8]), .B(n24), .Y(ab_8__0_) );
  AND2X1 U64 ( .A(A[5]), .B(B[1]), .Y(ab_5__1_) );
  AND2X1 U65 ( .A(A[10]), .B(n24), .Y(ab_10__0_) );
  AND2X1 U66 ( .A(A[11]), .B(n24), .Y(ab_11__0_) );
  INVXL U67 ( .A(B[1]), .Y(n34) );
  NOR2XL U68 ( .A(n38), .B(n35), .Y(ab_15__7_) );
  NOR2XL U69 ( .A(n37), .B(n29), .Y(ab_16__6_) );
  NOR2XL U70 ( .A(n40), .B(n35), .Y(ab_13__7_) );
  NOR2XL U71 ( .A(n39), .B(n29), .Y(ab_14__6_) );
  NOR2XL U72 ( .A(n41), .B(n34), .Y(ab_12__1_) );
  NAND2XL U73 ( .A(A[1]), .B(B[1]), .Y(n28) );
  AND2X1 U74 ( .A(A[3]), .B(n24), .Y(ab_3__0_) );
  NOR2XL U75 ( .A(n28), .B(n27), .Y(CARRYB_1__0_) );
  AND2X1 U76 ( .A(A[2]), .B(B[1]), .Y(ab_2__1_) );
  AND2X1 U77 ( .A(A[2]), .B(n24), .Y(ab_2__0_) );
  NOR2XL U78 ( .A(n37), .B(n35), .Y(ab_16__7_) );
  AND2X1 U79 ( .A(A[6]), .B(n23), .Y(ab_6__7_) );
  AND2X1 U80 ( .A(A[4]), .B(n23), .Y(ab_4__7_) );
  AND2X1 U81 ( .A(A[7]), .B(n23), .Y(ab_7__7_) );
  AND2X1 U82 ( .A(A[10]), .B(n23), .Y(ab_10__7_) );
  AND2X1 U83 ( .A(A[9]), .B(n23), .Y(ab_9__7_) );
  AND2X1 U84 ( .A(A[11]), .B(n23), .Y(ab_11__7_) );
  NAND2XL U85 ( .A(A[0]), .B(n24), .Y(n27) );
  XOR2X1 U86 ( .A(CARRYB_16__4_), .B(SUMB_16__5_), .Y(A1_19_) );
  AND2X2 U87 ( .A(CARRYB_16__2_), .B(SUMB_16__3_), .Y(n19) );
  AND2X2 U88 ( .A(CARRYB_16__4_), .B(SUMB_16__5_), .Y(n22) );
  NOR2X1 U89 ( .A(n37), .B(n34), .Y(ab_16__1_) );
  NOR2X1 U90 ( .A(n37), .B(n32), .Y(ab_16__3_) );
  NOR2X1 U91 ( .A(n37), .B(n30), .Y(ab_16__5_) );
  INVX1 U92 ( .A(n28), .Y(n36) );
  AND2X2 U93 ( .A(A[4]), .B(B[2]), .Y(ab_4__2_) );
  AND2X1 U94 ( .A(A[11]), .B(B[3]), .Y(ab_11__3_) );
  AND2X1 U95 ( .A(A[10]), .B(B[3]), .Y(ab_10__3_) );
  AND2X1 U96 ( .A(A[9]), .B(B[3]), .Y(ab_9__3_) );
  AND2X1 U97 ( .A(A[11]), .B(B[4]), .Y(ab_11__4_) );
  AND2X1 U98 ( .A(A[10]), .B(B[4]), .Y(ab_10__4_) );
  AND2X1 U99 ( .A(A[9]), .B(B[4]), .Y(ab_9__4_) );
  AND2X1 U100 ( .A(A[8]), .B(B[3]), .Y(ab_8__3_) );
  AND2X1 U101 ( .A(A[8]), .B(B[4]), .Y(ab_8__4_) );
  AND2X1 U102 ( .A(A[7]), .B(B[3]), .Y(ab_7__3_) );
  AND2X1 U103 ( .A(A[7]), .B(B[4]), .Y(ab_7__4_) );
  AND2X1 U104 ( .A(A[6]), .B(B[4]), .Y(ab_6__4_) );
  AND2X1 U105 ( .A(A[6]), .B(B[3]), .Y(ab_6__3_) );
  AND2X1 U106 ( .A(A[5]), .B(B[4]), .Y(ab_5__4_) );
  AND2X2 U107 ( .A(A[8]), .B(B[1]), .Y(ab_8__1_) );
  AND2X1 U108 ( .A(A[5]), .B(B[3]), .Y(ab_5__3_) );
  AND2X1 U109 ( .A(A[4]), .B(B[4]), .Y(ab_4__4_) );
  AND2X1 U110 ( .A(A[4]), .B(B[3]), .Y(ab_4__3_) );
  AND2X2 U111 ( .A(A[9]), .B(n24), .Y(ab_9__0_) );
  AND2X2 U112 ( .A(A[4]), .B(B[1]), .Y(ab_4__1_) );
  AND2X2 U113 ( .A(A[6]), .B(B[1]), .Y(ab_6__1_) );
  AND2X2 U114 ( .A(A[5]), .B(n24), .Y(ab_5__0_) );
  AND2X2 U115 ( .A(A[4]), .B(n24), .Y(ab_4__0_) );
  AND2X2 U116 ( .A(A[7]), .B(n24), .Y(ab_7__0_) );
  AND2X2 U117 ( .A(A[6]), .B(n24), .Y(ab_6__0_) );
  XOR2X1 U118 ( .A(n36), .B(ab_0__2_), .Y(SUMB_1__1_) );
  XOR2X1 U119 ( .A(CARRYB_16__5_), .B(SUMB_16__6_), .Y(A1_20_) );
  XOR2X1 U120 ( .A(CARRYB_16__6_), .B(ab_16__7_), .Y(A1_21_) );
  INVX1 U121 ( .A(B[0]), .Y(n25) );
  NOR2X2 U122 ( .A(n30), .B(n26), .Y(ab_0__5_) );
  AND2X1 U123 ( .A(A[3]), .B(B[2]), .Y(ab_3__2_) );
  NOR2X1 U124 ( .A(n39), .B(n34), .Y(ab_14__1_) );
  NOR2X1 U125 ( .A(n40), .B(n34), .Y(ab_13__1_) );
  NOR2XL U126 ( .A(n39), .B(n32), .Y(ab_14__3_) );
  NOR2XL U127 ( .A(n41), .B(n32), .Y(ab_12__3_) );
  AND2X1 U128 ( .A(A[10]), .B(B[5]), .Y(ab_10__5_) );
  NOR2XL U129 ( .A(n41), .B(n30), .Y(ab_12__5_) );
  AND2X1 U130 ( .A(A[9]), .B(B[5]), .Y(ab_9__5_) );
  NOR2XL U131 ( .A(n39), .B(n30), .Y(ab_14__5_) );
  AND2X1 U132 ( .A(A[8]), .B(B[5]), .Y(ab_8__5_) );
  AND2X1 U133 ( .A(A[7]), .B(B[5]), .Y(ab_7__5_) );
  AND2X1 U134 ( .A(A[6]), .B(B[5]), .Y(ab_6__5_) );
  AND2X1 U135 ( .A(A[5]), .B(B[5]), .Y(ab_5__5_) );
  NOR2X1 U136 ( .A(n41), .B(n35), .Y(ab_12__7_) );
  AND2X1 U137 ( .A(A[4]), .B(B[5]), .Y(ab_4__5_) );
  AND2X1 U138 ( .A(A[3]), .B(B[4]), .Y(ab_3__4_) );
  AND2X1 U139 ( .A(A[3]), .B(B[3]), .Y(ab_3__3_) );
  AND2X1 U140 ( .A(A[3]), .B(B[1]), .Y(ab_3__1_) );
  AND2X1 U141 ( .A(A[3]), .B(B[5]), .Y(ab_3__5_) );
  AND2X1 U142 ( .A(A[2]), .B(B[2]), .Y(ab_2__2_) );
  NOR2X1 U143 ( .A(n39), .B(n35), .Y(ab_14__7_) );
  AND2X1 U144 ( .A(A[2]), .B(B[5]), .Y(ab_2__5_) );
  XOR2X1 U145 ( .A(ab_1__6_), .B(ab_0__7_), .Y(SUMB_1__6_) );
  NOR2X1 U146 ( .A(n38), .B(n34), .Y(ab_15__1_) );
  NOR2XL U147 ( .A(n40), .B(n32), .Y(ab_13__3_) );
  NOR2XL U148 ( .A(n38), .B(n32), .Y(ab_15__3_) );
  AND2X1 U149 ( .A(A[11]), .B(B[5]), .Y(ab_11__5_) );
  NOR2XL U150 ( .A(n40), .B(n30), .Y(ab_13__5_) );
  NOR2XL U151 ( .A(n38), .B(n30), .Y(ab_15__5_) );
  AND2X1 U152 ( .A(A[2]), .B(B[3]), .Y(ab_2__3_) );
  XOR2X1 U153 ( .A(ab_1__4_), .B(ab_0__5_), .Y(SUMB_1__4_) );
  INVX1 U154 ( .A(A[16]), .Y(n37) );
  AND2X2 U155 ( .A(A[8]), .B(n23), .Y(ab_8__7_) );
  AND2X2 U156 ( .A(A[5]), .B(n23), .Y(ab_5__7_) );
  AND2X1 U157 ( .A(A[3]), .B(n23), .Y(ab_3__7_) );
  AND2X1 U158 ( .A(A[2]), .B(n23), .Y(ab_2__7_) );
  AND2X1 U159 ( .A(A[1]), .B(n23), .Y(ab_1__7_) );
  NOR2XL U160 ( .A(n41), .B(n29), .Y(ab_12__6_) );
  INVX1 U161 ( .A(A[12]), .Y(n41) );
  INVX1 U162 ( .A(A[13]), .Y(n40) );
  INVX1 U163 ( .A(A[14]), .Y(n39) );
  INVX1 U164 ( .A(A[15]), .Y(n38) );
  NOR2XL U165 ( .A(n37), .B(n31), .Y(ab_16__4_) );
  NOR2XL U166 ( .A(n38), .B(n31), .Y(ab_15__4_) );
  NOR2XL U167 ( .A(n39), .B(n31), .Y(ab_14__4_) );
  NOR2XL U168 ( .A(n40), .B(n31), .Y(ab_13__4_) );
  NOR2XL U169 ( .A(n41), .B(n31), .Y(ab_12__4_) );
  AND2X2 U170 ( .A(A[1]), .B(B[6]), .Y(ab_1__6_) );
  AND2X1 U171 ( .A(A[11]), .B(B[6]), .Y(ab_11__6_) );
  AND2X1 U172 ( .A(A[10]), .B(B[6]), .Y(ab_10__6_) );
  AND2X1 U173 ( .A(A[9]), .B(B[6]), .Y(ab_9__6_) );
  AND2X1 U174 ( .A(A[8]), .B(B[6]), .Y(ab_8__6_) );
  AND2X1 U175 ( .A(A[7]), .B(B[6]), .Y(ab_7__6_) );
  AND2X1 U176 ( .A(A[6]), .B(B[6]), .Y(ab_6__6_) );
  AND2X1 U177 ( .A(A[5]), .B(B[6]), .Y(ab_5__6_) );
  AND2X1 U178 ( .A(A[4]), .B(B[6]), .Y(ab_4__6_) );
  AND2X1 U179 ( .A(A[3]), .B(B[6]), .Y(ab_3__6_) );
  AND2X1 U180 ( .A(A[2]), .B(B[6]), .Y(ab_2__6_) );
  NOR2XL U181 ( .A(n37), .B(n33), .Y(ab_16__2_) );
  NOR2XL U182 ( .A(n38), .B(n33), .Y(ab_15__2_) );
  NOR2XL U183 ( .A(n39), .B(n33), .Y(ab_14__2_) );
  NOR2XL U184 ( .A(n40), .B(n33), .Y(ab_13__2_) );
  NOR2XL U185 ( .A(n41), .B(n33), .Y(ab_12__2_) );
  NOR2X1 U187 ( .A(n25), .B(n37), .Y(ab_16__0_) );
  NOR2X1 U188 ( .A(n25), .B(n38), .Y(ab_15__0_) );
  NOR2X1 U189 ( .A(n25), .B(n39), .Y(ab_14__0_) );
  NOR2X1 U190 ( .A(n25), .B(n40), .Y(ab_13__0_) );
  NOR2X1 U191 ( .A(n25), .B(n41), .Y(ab_12__0_) );
endmodule


module multi16_1 ( in_17bit, in_8bit, out );
  input [16:0] in_17bit;
  input [7:0] in_8bit;
  output [16:0] out;
  wire   N19, N20, N21, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112;
  wire   [16:1] in_17bit_b;
  wire   [7:1] in_8bit_b;
  wire   [23:8] mul;
  wire   [16:13] sub_add_52_b0_carry;

  multi16_1_DW02_mult_0 mult_55 ( .A({in_17bit_b, in_17bit[0]}), .B({in_8bit_b, 
        n19}), .PRODUCT_23_(mul[23]), .PRODUCT_22_(mul[22]), .PRODUCT_21_(
        mul[21]), .PRODUCT_20_(mul[20]), .PRODUCT_19_(mul[19]), .PRODUCT_18_(
        mul[18]), .PRODUCT_17_(mul[17]), .PRODUCT_16_(mul[16]), .PRODUCT_15_(
        mul[15]), .PRODUCT_14_(mul[14]), .PRODUCT_13_(mul[13]), .PRODUCT_12_(
        mul[12]), .PRODUCT_11_(mul[11]), .PRODUCT_10_(mul[10]), .PRODUCT_9_(
        mul[9]), .PRODUCT_8_(mul[8]), .PRODUCT_7_(out[0]) );
  NOR2X2 U2 ( .A(in_8bit[1]), .B(n33), .Y(n31) );
  INVX4 U3 ( .A(n104), .Y(n107) );
  CLKINVX4 U4 ( .A(n95), .Y(n97) );
  NAND2BX1 U5 ( .AN(mul[17]), .B(n94), .Y(n95) );
  AOI21X2 U6 ( .A0(n31), .A1(n30), .B0(n6), .Y(n32) );
  INVX4 U7 ( .A(n96), .Y(n2) );
  NOR2X4 U8 ( .A(n11), .B(n97), .Y(n96) );
  XOR2X2 U9 ( .A(mul[17]), .B(n93), .Y(out[10]) );
  NOR2X2 U10 ( .A(n11), .B(n94), .Y(n93) );
  AOI21X1 U11 ( .A0(n107), .A1(n106), .B0(n11), .Y(n108) );
  CLKINVX2 U12 ( .A(n92), .Y(n94) );
  NOR2X2 U13 ( .A(n22), .B(n43), .Y(n42) );
  CLKINVX2 U14 ( .A(n41), .Y(n43) );
  XOR2X2 U15 ( .A(in_17bit[3]), .B(n42), .Y(in_17bit_b[3]) );
  INVX8 U16 ( .A(n23), .Y(n21) );
  XOR2X2 U17 ( .A(n32), .B(in_8bit[5]), .Y(in_8bit_b[5]) );
  INVX1 U18 ( .A(n87), .Y(n88) );
  NOR2X1 U19 ( .A(in_8bit[1]), .B(n33), .Y(n5) );
  XOR2X1 U20 ( .A(mul[14]), .B(n85), .Y(out[7]) );
  INVX1 U21 ( .A(n89), .Y(n91) );
  NAND2BX1 U22 ( .AN(mul[15]), .B(n88), .Y(n89) );
  NOR2X1 U23 ( .A(mul[12]), .B(n81), .Y(n7) );
  NAND2BX1 U24 ( .AN(mul[16]), .B(n91), .Y(n92) );
  XOR2X1 U25 ( .A(mul[15]), .B(n9), .Y(out[8]) );
  XOR2X1 U26 ( .A(n10), .B(n45), .Y(in_17bit_b[4]) );
  OR2X2 U27 ( .A(n22), .B(n46), .Y(n10) );
  CLKINVX3 U28 ( .A(in_8bit[2]), .Y(n26) );
  INVX2 U29 ( .A(mul[22]), .Y(n106) );
  NOR3X1 U30 ( .A(in_8bit[6]), .B(n37), .C(n6), .Y(in_8bit_b[7]) );
  OR2X2 U31 ( .A(n5), .B(n6), .Y(n27) );
  XOR2X2 U32 ( .A(mul[21]), .B(n103), .Y(out[14]) );
  CLKINVX3 U33 ( .A(in_17bit[16]), .Y(n23) );
  INVX1 U34 ( .A(in_8bit[4]), .Y(n20) );
  NOR2X2 U35 ( .A(n11), .B(n15), .Y(n103) );
  NOR2X2 U36 ( .A(n11), .B(n102), .Y(n98) );
  NOR2X1 U37 ( .A(n11), .B(n91), .Y(n90) );
  NOR2X1 U38 ( .A(n11), .B(n88), .Y(n9) );
  NOR2X1 U39 ( .A(n11), .B(n86), .Y(n85) );
  NOR2X1 U40 ( .A(n11), .B(n7), .Y(n8) );
  INVXL U41 ( .A(in_8bit[3]), .Y(n36) );
  NOR3XL U42 ( .A(n33), .B(in_8bit[3]), .C(in_8bit[1]), .Y(n28) );
  INVX4 U43 ( .A(n33), .Y(n34) );
  NAND2BXL U44 ( .AN(in_17bit[2]), .B(n18), .Y(n41) );
  INVX4 U45 ( .A(n100), .Y(n102) );
  NOR3BX4 U46 ( .AN(n39), .B(n38), .C(n18), .Y(in_17bit_b[1]) );
  XOR2X4 U47 ( .A(n25), .B(n26), .Y(in_8bit_b[2]) );
  OAI21X4 U48 ( .A0(in_8bit[1]), .A1(n19), .B0(in_8bit[7]), .Y(n25) );
  NAND2X4 U49 ( .A(mul[18]), .B(n2), .Y(n3) );
  NAND3X1 U50 ( .A(in_17bit[1]), .B(n21), .C(in_17bit[0]), .Y(n39) );
  NOR2X1 U51 ( .A(n21), .B(in_17bit[1]), .Y(n38) );
  NAND2X2 U52 ( .A(n37), .B(in_8bit[7]), .Y(n14) );
  NAND2X2 U53 ( .A(n1), .B(n96), .Y(n4) );
  NAND2X4 U54 ( .A(n3), .B(n4), .Y(out[11]) );
  INVXL U55 ( .A(mul[18]), .Y(n1) );
  INVX1 U56 ( .A(in_8bit[7]), .Y(n6) );
  NOR2X4 U57 ( .A(in_17bit[1]), .B(in_17bit[0]), .Y(n18) );
  NOR2X2 U58 ( .A(n23), .B(n18), .Y(n40) );
  NOR2X1 U59 ( .A(in_8bit[5]), .B(in_8bit[4]), .Y(n35) );
  NAND4BX2 U60 ( .AN(in_8bit[1]), .B(n36), .C(n35), .D(n34), .Y(n37) );
  NAND2X1 U61 ( .A(n48), .B(n21), .Y(n47) );
  NAND2X1 U62 ( .A(n55), .B(n21), .Y(n54) );
  NAND2XL U63 ( .A(n62), .B(n21), .Y(n61) );
  NOR2XL U64 ( .A(in_8bit[4]), .B(in_8bit[3]), .Y(n30) );
  XNOR2XL U65 ( .A(n21), .B(in_8bit[7]), .Y(n11) );
  NAND2BX4 U66 ( .AN(n19), .B(n26), .Y(n33) );
  BUFX8 U67 ( .A(in_8bit[0]), .Y(n19) );
  NAND2BX2 U68 ( .AN(mul[21]), .B(n15), .Y(n104) );
  XOR2X1 U69 ( .A(mul[13]), .B(n8), .Y(out[6]) );
  NOR2X1 U70 ( .A(n11), .B(n77), .Y(n76) );
  INVXL U71 ( .A(n102), .Y(n16) );
  NAND2BXL U72 ( .AN(mul[9]), .B(n17), .Y(n75) );
  NAND2BXL U73 ( .AN(mul[10]), .B(n77), .Y(n78) );
  NAND2BXL U74 ( .AN(mul[11]), .B(n80), .Y(n81) );
  NAND2XL U75 ( .A(out[0]), .B(n99), .Y(n73) );
  XOR2X1 U76 ( .A(mul[16]), .B(n90), .Y(out[9]) );
  NOR2XL U77 ( .A(n11), .B(n83), .Y(n82) );
  NOR2XL U78 ( .A(n11), .B(n17), .Y(n74) );
  NOR2X2 U79 ( .A(n28), .B(n6), .Y(n29) );
  NAND2XL U80 ( .A(n46), .B(n45), .Y(n48) );
  NAND2BXL U81 ( .AN(n48), .B(n49), .Y(n50) );
  NOR2XL U82 ( .A(n22), .B(n60), .Y(n58) );
  NAND2XL U83 ( .A(n53), .B(n52), .Y(n55) );
  NAND2XL U84 ( .A(n60), .B(n59), .Y(n62) );
  NAND2BXL U85 ( .AN(n55), .B(n56), .Y(n57) );
  NAND2XL U86 ( .A(n71), .B(n21), .Y(n68) );
  NAND3BXL U87 ( .AN(n71), .B(n109), .C(n70), .Y(n72) );
  NOR2XL U88 ( .A(n22), .B(n67), .Y(n65) );
  NAND2BXL U89 ( .AN(n62), .B(n63), .Y(n64) );
  AND2X1 U90 ( .A(N21), .B(n21), .Y(in_17bit_b[16]) );
  INVX1 U91 ( .A(n44), .Y(n46) );
  MX2X1 U92 ( .A(in_17bit[14]), .B(N19), .S0(n21), .Y(in_17bit_b[14]) );
  MX2X1 U93 ( .A(in_17bit[12]), .B(n12), .S0(n21), .Y(in_17bit_b[12]) );
  XNOR2X1 U94 ( .A(in_17bit[12]), .B(n69), .Y(n12) );
  MX2X1 U95 ( .A(in_17bit[13]), .B(n13), .S0(n21), .Y(in_17bit_b[13]) );
  XNOR2X1 U96 ( .A(n72), .B(n110), .Y(n13) );
  MX2X1 U97 ( .A(in_17bit[15]), .B(N20), .S0(n21), .Y(in_17bit_b[15]) );
  NOR2XL U98 ( .A(in_17bit[11]), .B(n71), .Y(n69) );
  XNOR2X4 U99 ( .A(n14), .B(in_8bit[6]), .Y(in_8bit_b[6]) );
  NAND2BX4 U100 ( .AN(mul[18]), .B(n97), .Y(n100) );
  NOR3X4 U101 ( .A(mul[20]), .B(n16), .C(mul[19]), .Y(n15) );
  INVX1 U102 ( .A(n78), .Y(n80) );
  INVX1 U103 ( .A(n81), .Y(n83) );
  NOR2X1 U104 ( .A(mul[8]), .B(out[0]), .Y(n17) );
  INVX1 U105 ( .A(n75), .Y(n77) );
  XOR2X1 U106 ( .A(mul[23]), .B(n108), .Y(out[16]) );
  XNOR2X1 U107 ( .A(mul[8]), .B(n73), .Y(out[1]) );
  NAND2BX1 U108 ( .AN(mul[14]), .B(n86), .Y(n87) );
  INVX1 U109 ( .A(n84), .Y(n86) );
  NAND2BX1 U110 ( .AN(mul[13]), .B(n7), .Y(n84) );
  XOR2X1 U111 ( .A(mul[11]), .B(n79), .Y(out[4]) );
  NOR2X1 U112 ( .A(n11), .B(n80), .Y(n79) );
  XOR2X1 U113 ( .A(mul[12]), .B(n82), .Y(out[5]) );
  XOR2X1 U114 ( .A(mul[10]), .B(n76), .Y(out[3]) );
  XOR2X1 U115 ( .A(mul[9]), .B(n74), .Y(out[2]) );
  XOR2X4 U116 ( .A(n98), .B(mul[19]), .Y(out[12]) );
  INVX1 U117 ( .A(n11), .Y(n99) );
  XNOR2X1 U118 ( .A(in_8bit[1]), .B(n24), .Y(in_8bit_b[1]) );
  XNOR2X1 U119 ( .A(n51), .B(n52), .Y(in_17bit_b[6]) );
  NOR2X1 U120 ( .A(n22), .B(n53), .Y(n51) );
  XNOR2X1 U121 ( .A(n58), .B(n59), .Y(in_17bit_b[8]) );
  XOR2X1 U122 ( .A(n49), .B(n47), .Y(in_17bit_b[5]) );
  XOR2X1 U123 ( .A(n63), .B(n61), .Y(in_17bit_b[9]) );
  XOR2X1 U124 ( .A(n56), .B(n54), .Y(in_17bit_b[7]) );
  INVX1 U125 ( .A(n50), .Y(n53) );
  INVX1 U126 ( .A(n57), .Y(n60) );
  NAND2X1 U127 ( .A(n67), .B(n66), .Y(n71) );
  XNOR2X1 U128 ( .A(n65), .B(n66), .Y(in_17bit_b[10]) );
  XOR2X1 U129 ( .A(n70), .B(n68), .Y(in_17bit_b[11]) );
  INVX1 U130 ( .A(n72), .Y(sub_add_52_b0_carry[13]) );
  INVX1 U131 ( .A(n64), .Y(n67) );
  XOR2X2 U132 ( .A(in_17bit[2]), .B(n40), .Y(in_17bit_b[2]) );
  INVX1 U133 ( .A(in_17bit[4]), .Y(n45) );
  INVX1 U134 ( .A(in_17bit[5]), .Y(n49) );
  NAND2BXL U135 ( .AN(in_17bit[3]), .B(n43), .Y(n44) );
  INVX1 U136 ( .A(in_17bit[16]), .Y(n22) );
  INVX1 U137 ( .A(in_17bit[6]), .Y(n52) );
  INVX1 U138 ( .A(in_17bit[8]), .Y(n59) );
  INVX1 U139 ( .A(in_17bit[7]), .Y(n56) );
  INVX1 U140 ( .A(in_17bit[10]), .Y(n66) );
  INVX1 U141 ( .A(in_17bit[11]), .Y(n70) );
  INVX1 U142 ( .A(in_17bit[9]), .Y(n63) );
  INVX1 U143 ( .A(in_17bit[12]), .Y(n109) );
  INVX1 U144 ( .A(in_17bit[13]), .Y(n110) );
  INVX1 U145 ( .A(in_17bit[14]), .Y(n111) );
  INVX1 U146 ( .A(in_17bit[15]), .Y(n112) );
  NAND2XL U147 ( .A(n19), .B(in_8bit[7]), .Y(n24) );
  XOR2X4 U148 ( .A(n27), .B(n36), .Y(in_8bit_b[3]) );
  XNOR2X4 U149 ( .A(n29), .B(n20), .Y(in_8bit_b[4]) );
  OAI21X4 U150 ( .A0(mul[19]), .A1(n100), .B0(n99), .Y(n101) );
  XNOR2X4 U151 ( .A(mul[20]), .B(n101), .Y(out[13]) );
  NOR2X4 U152 ( .A(n11), .B(n107), .Y(n105) );
  XNOR2X4 U153 ( .A(n105), .B(n106), .Y(out[15]) );
  XOR2X1 U154 ( .A(n22), .B(sub_add_52_b0_carry[16]), .Y(N21) );
  AND2X1 U155 ( .A(sub_add_52_b0_carry[15]), .B(n112), .Y(
        sub_add_52_b0_carry[16]) );
  XOR2X1 U156 ( .A(n112), .B(sub_add_52_b0_carry[15]), .Y(N20) );
  AND2X1 U157 ( .A(sub_add_52_b0_carry[14]), .B(n111), .Y(
        sub_add_52_b0_carry[15]) );
  XOR2X1 U158 ( .A(n111), .B(sub_add_52_b0_carry[14]), .Y(N19) );
  AND2X1 U159 ( .A(sub_add_52_b0_carry[13]), .B(n110), .Y(
        sub_add_52_b0_carry[14]) );
endmodule


module multi16_0_DW01_add_0 ( A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, 
        A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, 
        B_20_, B_19_, B_18_, B_17_, B_16_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, 
        SUM_17_, SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, 
        SUM_9_, SUM_8_, SUM_7_, SUM_6_, SUM_5_ );
  input A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_,
         A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, B_21_, B_20_, B_19_,
         B_18_, B_17_, B_16_;
  output SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, SUM_15_,
         SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, SUM_7_,
         SUM_6_, SUM_5_;
  wire   n1, n3, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39;

  INVX2 U2 ( .A(n20), .Y(SUM_15_) );
  XOR2X2 U3 ( .A(n38), .B(n37), .Y(SUM_18_) );
  NOR2X4 U4 ( .A(n29), .B(n17), .Y(n39) );
  NOR2X1 U5 ( .A(B_16_), .B(A_16_), .Y(n3) );
  XOR2X2 U6 ( .A(n1), .B(n23), .Y(SUM_20_) );
  NOR2BX2 U7 ( .AN(n33), .B(n3), .Y(SUM_16_) );
  AOI21X2 U8 ( .A0(n19), .A1(n18), .B0(n17), .Y(n37) );
  INVX2 U9 ( .A(n29), .Y(n18) );
  BUFX3 U10 ( .A(A_12_), .Y(SUM_12_) );
  INVX2 U11 ( .A(n34), .Y(n17) );
  BUFX3 U12 ( .A(A_13_), .Y(SUM_13_) );
  BUFX3 U13 ( .A(A_14_), .Y(SUM_14_) );
  INVX1 U14 ( .A(A_15_), .Y(n20) );
  NOR2X1 U15 ( .A(B_18_), .B(A_18_), .Y(n30) );
  XOR2X2 U16 ( .A(n19), .B(n39), .Y(SUM_17_) );
  NAND2X2 U17 ( .A(B_16_), .B(A_16_), .Y(n33) );
  NAND2X1 U18 ( .A(B_17_), .B(A_17_), .Y(n34) );
  AOI21XL U19 ( .A0(n15), .A1(n31), .B0(n16), .Y(n26) );
  OAI21X1 U20 ( .A0(n37), .A1(n30), .B0(n32), .Y(n35) );
  NOR2X4 U21 ( .A(B_17_), .B(A_17_), .Y(n29) );
  AND2X2 U22 ( .A(n25), .B(n24), .Y(n1) );
  INVXL U23 ( .A(n25), .Y(n14) );
  OR2X2 U24 ( .A(B_20_), .B(A_20_), .Y(n24) );
  OAI21XL U25 ( .A0(n26), .A1(n27), .B0(n28), .Y(n23) );
  INVXL U26 ( .A(n32), .Y(n16) );
  INVX2 U27 ( .A(n33), .Y(n19) );
  INVX1 U28 ( .A(n30), .Y(n15) );
  BUFX3 U29 ( .A(A_5_), .Y(SUM_5_) );
  BUFX3 U30 ( .A(A_6_), .Y(SUM_6_) );
  BUFX3 U31 ( .A(A_7_), .Y(SUM_7_) );
  BUFX3 U32 ( .A(A_8_), .Y(SUM_8_) );
  BUFX3 U33 ( .A(A_10_), .Y(SUM_10_) );
  BUFX3 U34 ( .A(A_11_), .Y(SUM_11_) );
  BUFX3 U35 ( .A(A_9_), .Y(SUM_9_) );
  XOR2X1 U36 ( .A(n21), .B(n22), .Y(SUM_21_) );
  AOI21X1 U37 ( .A0(n23), .A1(n24), .B0(n14), .Y(n22) );
  XNOR2X1 U38 ( .A(B_21_), .B(A_21_), .Y(n21) );
  OAI21XL U39 ( .A0(n29), .A1(n33), .B0(n34), .Y(n31) );
  NAND2X1 U40 ( .A(B_20_), .B(A_20_), .Y(n25) );
  XOR2X1 U41 ( .A(n35), .B(n36), .Y(SUM_19_) );
  NOR2BX1 U42 ( .AN(n28), .B(n27), .Y(n36) );
  NOR2X1 U43 ( .A(B_19_), .B(A_19_), .Y(n27) );
  NAND2X1 U44 ( .A(B_19_), .B(A_19_), .Y(n28) );
  NAND2X1 U45 ( .A(n32), .B(n15), .Y(n38) );
  NAND2X1 U46 ( .A(B_18_), .B(A_18_), .Y(n32) );
endmodule


module multi16_0_DW02_mult_0 ( A, B, PRODUCT_23_, PRODUCT_22_, PRODUCT_21_, 
        PRODUCT_20_, PRODUCT_19_, PRODUCT_18_, PRODUCT_17_, PRODUCT_16_, 
        PRODUCT_15_, PRODUCT_14_, PRODUCT_13_, PRODUCT_12_, PRODUCT_11_, 
        PRODUCT_10_, PRODUCT_9_, PRODUCT_8_, PRODUCT_7_ );
  input [16:0] A;
  input [7:0] B;
  output PRODUCT_23_, PRODUCT_22_, PRODUCT_21_, PRODUCT_20_, PRODUCT_19_,
         PRODUCT_18_, PRODUCT_17_, PRODUCT_16_, PRODUCT_15_, PRODUCT_14_,
         PRODUCT_13_, PRODUCT_12_, PRODUCT_11_, PRODUCT_10_, PRODUCT_9_,
         PRODUCT_8_, PRODUCT_7_;
  wire   ab_16__7_, ab_16__6_, ab_16__5_, ab_16__4_, ab_16__3_, ab_16__2_,
         ab_16__1_, ab_16__0_, ab_15__7_, ab_15__6_, ab_15__5_, ab_15__4_,
         ab_15__3_, ab_15__2_, ab_15__1_, ab_15__0_, ab_14__7_, ab_14__6_,
         ab_14__5_, ab_14__4_, ab_14__3_, ab_14__2_, ab_14__1_, ab_14__0_,
         ab_13__7_, ab_13__6_, ab_13__5_, ab_13__4_, ab_13__3_, ab_13__2_,
         ab_13__1_, ab_13__0_, ab_12__7_, ab_12__6_, ab_12__5_, ab_12__4_,
         ab_12__3_, ab_12__2_, ab_12__1_, ab_12__0_, ab_11__7_, ab_11__6_,
         ab_11__5_, ab_11__4_, ab_11__3_, ab_11__2_, ab_11__1_, ab_11__0_,
         ab_10__7_, ab_10__6_, ab_10__5_, ab_10__4_, ab_10__3_, ab_10__2_,
         ab_10__1_, ab_10__0_, ab_9__7_, ab_9__6_, ab_9__5_, ab_9__4_,
         ab_9__3_, ab_9__2_, ab_9__1_, ab_9__0_, ab_8__7_, ab_8__6_, ab_8__5_,
         ab_8__4_, ab_8__3_, ab_8__2_, ab_8__1_, ab_8__0_, ab_7__7_, ab_7__6_,
         ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_, ab_7__0_, ab_6__7_,
         ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_, ab_6__1_, ab_6__0_,
         ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_, ab_5__2_, ab_5__1_,
         ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_, ab_4__3_, ab_4__2_,
         ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_, ab_3__4_, ab_3__3_,
         ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_, ab_2__5_, ab_2__4_,
         ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_, ab_1__6_, ab_1__5_,
         ab_1__4_, ab_1__3_, ab_1__2_, ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_,
         ab_0__3_, ab_0__2_, CARRYB_16__6_, CARRYB_16__5_, CARRYB_16__4_,
         CARRYB_16__3_, CARRYB_16__2_, CARRYB_16__1_, CARRYB_16__0_,
         CARRYB_15__6_, CARRYB_15__5_, CARRYB_15__4_, CARRYB_15__3_,
         CARRYB_15__2_, CARRYB_15__1_, CARRYB_15__0_, CARRYB_14__6_,
         CARRYB_14__5_, CARRYB_14__4_, CARRYB_14__3_, CARRYB_14__2_,
         CARRYB_14__1_, CARRYB_14__0_, CARRYB_13__6_, CARRYB_13__5_,
         CARRYB_13__4_, CARRYB_13__3_, CARRYB_13__2_, CARRYB_13__1_,
         CARRYB_13__0_, CARRYB_12__6_, CARRYB_12__5_, CARRYB_12__4_,
         CARRYB_12__3_, CARRYB_12__2_, CARRYB_12__1_, CARRYB_12__0_,
         CARRYB_11__6_, CARRYB_11__5_, CARRYB_11__4_, CARRYB_11__3_,
         CARRYB_11__2_, CARRYB_11__1_, CARRYB_11__0_, CARRYB_10__6_,
         CARRYB_10__5_, CARRYB_10__4_, CARRYB_10__3_, CARRYB_10__2_,
         CARRYB_10__1_, CARRYB_10__0_, CARRYB_9__6_, CARRYB_9__5_,
         CARRYB_9__4_, CARRYB_9__3_, CARRYB_9__2_, CARRYB_9__1_, CARRYB_9__0_,
         CARRYB_8__6_, CARRYB_8__5_, CARRYB_8__4_, CARRYB_8__3_, CARRYB_8__2_,
         CARRYB_8__1_, CARRYB_8__0_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_,
         CARRYB_7__3_, CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_,
         CARRYB_6__5_, CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_,
         CARRYB_6__0_, CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_,
         CARRYB_5__2_, CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_,
         CARRYB_4__4_, CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_,
         CARRYB_3__6_, CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_,
         CARRYB_3__1_, CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_,
         CARRYB_2__3_, CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__6_,
         CARRYB_1__2_, CARRYB_1__0_, SUMB_16__6_, SUMB_16__5_, SUMB_16__4_,
         SUMB_16__3_, SUMB_16__2_, SUMB_16__1_, SUMB_16__0_, SUMB_15__6_,
         SUMB_15__5_, SUMB_15__4_, SUMB_15__3_, SUMB_15__2_, SUMB_15__1_,
         SUMB_14__6_, SUMB_14__5_, SUMB_14__4_, SUMB_14__3_, SUMB_14__2_,
         SUMB_14__1_, SUMB_13__6_, SUMB_13__5_, SUMB_13__4_, SUMB_13__3_,
         SUMB_13__2_, SUMB_13__1_, SUMB_12__6_, SUMB_12__5_, SUMB_12__4_,
         SUMB_12__3_, SUMB_12__2_, SUMB_12__1_, SUMB_11__6_, SUMB_11__5_,
         SUMB_11__4_, SUMB_11__3_, SUMB_11__2_, SUMB_11__1_, SUMB_10__6_,
         SUMB_10__5_, SUMB_10__4_, SUMB_10__3_, SUMB_10__2_, SUMB_10__1_,
         SUMB_9__6_, SUMB_9__5_, SUMB_9__4_, SUMB_9__3_, SUMB_9__2_,
         SUMB_9__1_, SUMB_8__6_, SUMB_8__5_, SUMB_8__4_, SUMB_8__3_,
         SUMB_8__2_, SUMB_8__1_, SUMB_7__6_, SUMB_7__5_, SUMB_7__4_,
         SUMB_7__3_, SUMB_7__2_, SUMB_7__1_, SUMB_6__6_, SUMB_6__5_,
         SUMB_6__4_, SUMB_6__3_, SUMB_6__2_, SUMB_6__1_, SUMB_5__6_,
         SUMB_5__5_, SUMB_5__4_, SUMB_5__3_, SUMB_5__2_, SUMB_5__1_,
         SUMB_4__6_, SUMB_4__5_, SUMB_4__4_, SUMB_4__3_, SUMB_4__2_,
         SUMB_4__1_, SUMB_3__6_, SUMB_3__5_, SUMB_3__4_, SUMB_3__3_,
         SUMB_3__2_, SUMB_3__1_, SUMB_2__6_, SUMB_2__5_, SUMB_2__4_,
         SUMB_2__3_, SUMB_2__2_, SUMB_2__1_, SUMB_1__6_, SUMB_1__5_,
         SUMB_1__4_, SUMB_1__3_, SUMB_1__2_, SUMB_1__1_, PROD1_7_, A1_21_,
         A1_20_, A1_19_, A1_18_, A1_17_, A1_16_, A1_15_, A1_13_, A1_12_,
         A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, A1_4_, A1_3_, A1_2_,
         A1_1_, A1_0_, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51;

  ADDFHX4 S1_15_0 ( .A(ab_15__0_), .B(CARRYB_14__0_), .CI(SUMB_14__1_), .CO(
        CARRYB_15__0_), .S(A1_13_) );
  ADDFHX4 S1_13_0 ( .A(ab_13__0_), .B(CARRYB_12__0_), .CI(SUMB_12__1_), .CO(
        CARRYB_13__0_), .S(A1_11_) );
  ADDFHX4 S2_13_1 ( .A(ab_13__1_), .B(CARRYB_12__1_), .CI(SUMB_12__2_), .CO(
        CARRYB_13__1_), .S(SUMB_13__1_) );
  ADDFHX4 S2_12_2 ( .A(ab_12__2_), .B(CARRYB_11__2_), .CI(SUMB_11__3_), .CO(
        CARRYB_12__2_), .S(SUMB_12__2_) );
  ADDFHX4 S2_11_1 ( .A(ab_11__1_), .B(CARRYB_10__1_), .CI(SUMB_10__2_), .CO(
        CARRYB_11__1_), .S(SUMB_11__1_) );
  ADDFHX4 S2_11_2 ( .A(ab_11__2_), .B(CARRYB_10__2_), .CI(SUMB_10__3_), .CO(
        CARRYB_11__2_), .S(SUMB_11__2_) );
  ADDFHX4 S2_11_3 ( .A(ab_11__3_), .B(CARRYB_10__3_), .CI(SUMB_10__4_), .CO(
        CARRYB_11__3_), .S(SUMB_11__3_) );
  ADDFHX4 S2_10_1 ( .A(ab_10__1_), .B(CARRYB_9__1_), .CI(SUMB_9__2_), .CO(
        CARRYB_10__1_), .S(SUMB_10__1_) );
  ADDFHX4 S2_10_2 ( .A(ab_10__2_), .B(CARRYB_9__2_), .CI(SUMB_9__3_), .CO(
        CARRYB_10__2_), .S(SUMB_10__2_) );
  ADDFHX4 S2_10_3 ( .A(ab_10__3_), .B(CARRYB_9__3_), .CI(SUMB_9__4_), .CO(
        CARRYB_10__3_), .S(SUMB_10__3_) );
  ADDFHX4 S2_10_4 ( .A(ab_10__4_), .B(CARRYB_9__4_), .CI(SUMB_9__5_), .CO(
        CARRYB_10__4_), .S(SUMB_10__4_) );
  ADDFHX4 S2_8_1 ( .A(ab_8__1_), .B(CARRYB_7__1_), .CI(SUMB_7__2_), .CO(
        CARRYB_8__1_), .S(SUMB_8__1_) );
  ADDFHX4 S2_8_3 ( .A(ab_8__3_), .B(CARRYB_7__3_), .CI(SUMB_7__4_), .CO(
        CARRYB_8__3_), .S(SUMB_8__3_) );
  ADDFHX4 S2_7_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  ADDFHX4 S2_7_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  ADDFHX4 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  ADDFHX4 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  multi16_0_DW01_add_0 FS_1 ( .A_21_(A1_21_), .A_20_(A1_20_), .A_19_(A1_19_), 
        .A_18_(A1_18_), .A_17_(A1_17_), .A_16_(A1_16_), .A_15_(A1_15_), 
        .A_14_(SUMB_16__0_), .A_13_(A1_13_), .A_12_(A1_12_), .A_11_(A1_11_), 
        .A_10_(A1_10_), .A_9_(A1_9_), .A_8_(A1_8_), .A_7_(A1_7_), .A_6_(A1_6_), 
        .A_5_(PROD1_7_), .B_21_(n31), .B_20_(n30), .B_19_(n28), .B_18_(n27), 
        .B_17_(n26), .B_16_(n29), .SUM_21_(PRODUCT_23_), .SUM_20_(PRODUCT_22_), 
        .SUM_19_(PRODUCT_21_), .SUM_18_(PRODUCT_20_), .SUM_17_(PRODUCT_19_), 
        .SUM_16_(PRODUCT_18_), .SUM_15_(PRODUCT_17_), .SUM_14_(PRODUCT_16_), 
        .SUM_13_(PRODUCT_15_), .SUM_12_(PRODUCT_14_), .SUM_11_(PRODUCT_13_), 
        .SUM_10_(PRODUCT_12_), .SUM_9_(PRODUCT_11_), .SUM_8_(PRODUCT_10_), 
        .SUM_7_(PRODUCT_9_), .SUM_6_(PRODUCT_8_), .SUM_5_(PRODUCT_7_) );
  ADDFHX1 S2_15_5 ( .A(ab_15__5_), .B(CARRYB_14__5_), .CI(SUMB_14__6_), .CO(
        CARRYB_15__5_), .S(SUMB_15__5_) );
  ADDFHX2 S2_7_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  ADDFX2 S5_6 ( .A(ab_16__6_), .B(CARRYB_15__6_), .CI(ab_15__7_), .CO(
        CARRYB_16__6_), .S(SUMB_16__6_) );
  ADDFHX1 S4_5 ( .A(ab_16__5_), .B(CARRYB_15__5_), .CI(SUMB_15__6_), .CO(
        CARRYB_16__5_), .S(SUMB_16__5_) );
  ADDFHX2 S4_1 ( .A(ab_16__1_), .B(CARRYB_15__1_), .CI(SUMB_15__2_), .CO(
        CARRYB_16__1_), .S(SUMB_16__1_) );
  ADDFHX2 S2_9_5 ( .A(ab_9__5_), .B(CARRYB_8__5_), .CI(SUMB_8__6_), .CO(
        CARRYB_9__5_), .S(SUMB_9__5_) );
  ADDFHX4 S3_7_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(
        CARRYB_7__6_), .S(SUMB_7__6_) );
  ADDFHX4 S2_13_2 ( .A(ab_13__2_), .B(CARRYB_12__2_), .CI(SUMB_12__3_), .CO(
        CARRYB_13__2_), .S(SUMB_13__2_) );
  ADDFHX2 S4_2 ( .A(ab_16__2_), .B(CARRYB_15__2_), .CI(SUMB_15__3_), .CO(
        CARRYB_16__2_), .S(SUMB_16__2_) );
  ADDFHX4 S1_8_0 ( .A(ab_8__0_), .B(CARRYB_7__0_), .CI(SUMB_7__1_), .CO(
        CARRYB_8__0_), .S(A1_6_) );
  ADDFHX2 S2_14_4 ( .A(ab_14__4_), .B(CARRYB_13__4_), .CI(SUMB_13__5_), .CO(
        CARRYB_14__4_), .S(SUMB_14__4_) );
  ADDFHX4 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  ADDFHX4 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  ADDFHX2 S2_14_5 ( .A(ab_14__5_), .B(CARRYB_13__5_), .CI(SUMB_13__6_), .CO(
        CARRYB_14__5_), .S(SUMB_14__5_) );
  ADDFHX2 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  ADDFHX4 S1_10_0 ( .A(ab_10__0_), .B(CARRYB_9__0_), .CI(SUMB_9__1_), .CO(
        CARRYB_10__0_), .S(A1_8_) );
  ADDFHX4 S1_11_0 ( .A(ab_11__0_), .B(CARRYB_10__0_), .CI(SUMB_10__1_), .CO(
        CARRYB_11__0_), .S(A1_9_) );
  ADDFHX2 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  ADDFHX4 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  ADDFHX4 S2_13_4 ( .A(ab_13__4_), .B(CARRYB_12__4_), .CI(SUMB_12__5_), .CO(
        CARRYB_13__4_), .S(SUMB_13__4_) );
  ADDFHX4 S2_13_3 ( .A(ab_13__3_), .B(CARRYB_12__3_), .CI(SUMB_12__4_), .CO(
        CARRYB_13__3_), .S(SUMB_13__3_) );
  ADDFHX2 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  ADDFHX2 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  ADDFHX4 S2_14_2 ( .A(ab_14__2_), .B(CARRYB_13__2_), .CI(SUMB_13__3_), .CO(
        CARRYB_14__2_), .S(SUMB_14__2_) );
  ADDFHX2 S3_14_6 ( .A(ab_14__6_), .B(CARRYB_13__6_), .CI(ab_13__7_), .CO(
        CARRYB_14__6_), .S(SUMB_14__6_) );
  ADDFHX2 S2_2_1 ( .A(ab_2__1_), .B(n16), .CI(SUMB_1__2_), .CO(CARRYB_2__1_), 
        .S(SUMB_2__1_) );
  ADDFHX4 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  ADDFHX2 S2_2_5 ( .A(ab_2__5_), .B(n15), .CI(SUMB_1__6_), .CO(CARRYB_2__5_), 
        .S(SUMB_2__5_) );
  ADDFHX2 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  ADDFHX4 S2_14_3 ( .A(ab_14__3_), .B(CARRYB_13__3_), .CI(SUMB_13__4_), .CO(
        CARRYB_14__3_), .S(SUMB_14__3_) );
  ADDFHX2 S2_15_4 ( .A(ab_15__4_), .B(CARRYB_14__4_), .CI(SUMB_14__5_), .CO(
        CARRYB_15__4_), .S(SUMB_15__4_) );
  ADDFHX2 S2_13_5 ( .A(ab_13__5_), .B(CARRYB_12__5_), .CI(SUMB_12__6_), .CO(
        CARRYB_13__5_), .S(SUMB_13__5_) );
  ADDFHX4 S2_8_2 ( .A(ab_8__2_), .B(CARRYB_7__2_), .CI(SUMB_7__3_), .CO(
        CARRYB_8__2_), .S(SUMB_8__2_) );
  ADDFHX2 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  ADDFHX4 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  ADDFHX4 S3_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(ab_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  ADDFHX4 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  ADDFHX2 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  ADDFHX2 S3_10_6 ( .A(ab_10__6_), .B(CARRYB_9__6_), .CI(ab_9__7_), .CO(
        CARRYB_10__6_), .S(SUMB_10__6_) );
  ADDFHX4 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  ADDFHX4 S2_7_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  ADDFHX4 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  ADDFHX2 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  ADDFHX4 S2_2_4 ( .A(ab_2__4_), .B(n14), .CI(SUMB_1__5_), .CO(CARRYB_2__4_), 
        .S(SUMB_2__4_) );
  ADDFX2 S3_15_6 ( .A(ab_15__6_), .B(CARRYB_14__6_), .CI(ab_14__7_), .CO(
        CARRYB_15__6_), .S(SUMB_15__6_) );
  ADDFHX1 S4_4 ( .A(ab_16__4_), .B(CARRYB_15__4_), .CI(SUMB_15__5_), .CO(
        CARRYB_16__4_), .S(SUMB_16__4_) );
  ADDFHX2 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  ADDFHX2 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  ADDFHX2 S1_9_0 ( .A(ab_9__0_), .B(CARRYB_8__0_), .CI(SUMB_8__1_), .CO(
        CARRYB_9__0_), .S(A1_7_) );
  ADDFHX2 S1_12_0 ( .A(ab_12__0_), .B(CARRYB_11__0_), .CI(SUMB_11__1_), .CO(
        CARRYB_12__0_), .S(A1_10_) );
  ADDFHX2 S3_8_6 ( .A(ab_8__6_), .B(CARRYB_7__6_), .CI(ab_7__7_), .CO(
        CARRYB_8__6_), .S(SUMB_8__6_) );
  ADDFHX2 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  ADDFHX2 S2_2_3 ( .A(ab_2__3_), .B(n17), .CI(SUMB_1__4_), .CO(CARRYB_2__3_), 
        .S(SUMB_2__3_) );
  ADDFHX2 S2_9_1 ( .A(ab_9__1_), .B(CARRYB_8__1_), .CI(SUMB_8__2_), .CO(
        CARRYB_9__1_), .S(SUMB_9__1_) );
  ADDFHX2 S1_14_0 ( .A(ab_14__0_), .B(CARRYB_13__0_), .CI(SUMB_13__1_), .CO(
        CARRYB_14__0_), .S(A1_12_) );
  ADDFHX2 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  ADDFHX2 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  ADDFHX2 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  ADDFHX2 S2_12_3 ( .A(ab_12__3_), .B(CARRYB_11__3_), .CI(SUMB_11__4_), .CO(
        CARRYB_12__3_), .S(SUMB_12__3_) );
  ADDFHX2 S2_15_1 ( .A(ab_15__1_), .B(CARRYB_14__1_), .CI(SUMB_14__2_), .CO(
        CARRYB_15__1_), .S(SUMB_15__1_) );
  ADDFHX2 S3_11_6 ( .A(ab_11__6_), .B(CARRYB_10__6_), .CI(ab_10__7_), .CO(
        CARRYB_11__6_), .S(SUMB_11__6_) );
  ADDFHX2 S4_0 ( .A(ab_16__0_), .B(CARRYB_15__0_), .CI(SUMB_15__1_), .CO(
        CARRYB_16__0_), .S(SUMB_16__0_) );
  ADDFHX2 S2_8_5 ( .A(ab_8__5_), .B(CARRYB_7__5_), .CI(SUMB_7__6_), .CO(
        CARRYB_8__5_), .S(SUMB_8__5_) );
  ADDFHX4 S2_11_4 ( .A(ab_11__4_), .B(CARRYB_10__4_), .CI(SUMB_10__5_), .CO(
        CARRYB_11__4_), .S(SUMB_11__4_) );
  ADDFHX4 S2_12_4 ( .A(ab_12__4_), .B(CARRYB_11__4_), .CI(SUMB_11__5_), .CO(
        CARRYB_12__4_), .S(SUMB_12__4_) );
  ADDFHX4 S2_8_4 ( .A(ab_8__4_), .B(CARRYB_7__4_), .CI(SUMB_7__5_), .CO(
        CARRYB_8__4_), .S(SUMB_8__4_) );
  ADDFHX4 S2_9_4 ( .A(ab_9__4_), .B(CARRYB_8__4_), .CI(SUMB_8__5_), .CO(
        CARRYB_9__4_), .S(SUMB_9__4_) );
  ADDFHX4 S2_11_5 ( .A(ab_11__5_), .B(CARRYB_10__5_), .CI(SUMB_10__6_), .CO(
        CARRYB_11__5_), .S(SUMB_11__5_) );
  ADDFHX4 S2_12_5 ( .A(ab_12__5_), .B(CARRYB_11__5_), .CI(SUMB_11__6_), .CO(
        CARRYB_12__5_), .S(SUMB_12__5_) );
  ADDFHX4 S3_12_6 ( .A(ab_12__6_), .B(CARRYB_11__6_), .CI(ab_11__7_), .CO(
        CARRYB_12__6_), .S(SUMB_12__6_) );
  ADDFHX2 S3_13_6 ( .A(ab_13__6_), .B(CARRYB_12__6_), .CI(ab_12__7_), .CO(
        CARRYB_13__6_), .S(SUMB_13__6_) );
  ADDFHX2 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  ADDFHX4 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  ADDFHX4 S2_15_3 ( .A(ab_15__3_), .B(CARRYB_14__3_), .CI(SUMB_14__4_), .CO(
        CARRYB_15__3_), .S(SUMB_15__3_) );
  ADDFHX2 S4_3 ( .A(ab_16__3_), .B(CARRYB_15__3_), .CI(SUMB_15__4_), .CO(
        CARRYB_16__3_), .S(SUMB_16__3_) );
  ADDFHX4 S2_15_2 ( .A(ab_15__2_), .B(CARRYB_14__2_), .CI(SUMB_14__3_), .CO(
        CARRYB_15__2_), .S(SUMB_15__2_) );
  ADDFHX4 S2_9_2 ( .A(ab_9__2_), .B(CARRYB_8__2_), .CI(SUMB_8__3_), .CO(
        CARRYB_9__2_), .S(SUMB_9__2_) );
  ADDFHX4 S2_9_3 ( .A(ab_9__3_), .B(CARRYB_8__3_), .CI(SUMB_8__4_), .CO(
        CARRYB_9__3_), .S(SUMB_9__3_) );
  ADDFHX4 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  ADDFHX4 S2_12_1 ( .A(ab_12__1_), .B(CARRYB_11__1_), .CI(SUMB_11__2_), .CO(
        CARRYB_12__1_), .S(SUMB_12__1_) );
  ADDFHX4 S2_14_1 ( .A(ab_14__1_), .B(CARRYB_13__1_), .CI(SUMB_13__2_), .CO(
        CARRYB_14__1_), .S(SUMB_14__1_) );
  ADDFHX4 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  ADDFHX4 S1_7_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(PROD1_7_) );
  ADDFHX4 S3_9_6 ( .A(ab_9__6_), .B(CARRYB_8__6_), .CI(ab_8__7_), .CO(
        CARRYB_9__6_), .S(SUMB_9__6_) );
  AND2X2 U2 ( .A(A[1]), .B(B[6]), .Y(ab_1__6_) );
  INVX2 U3 ( .A(n32), .Y(CARRYB_1__2_) );
  AND2X4 U4 ( .A(ab_0__4_), .B(ab_1__3_), .Y(n17) );
  AND2X2 U5 ( .A(A[1]), .B(B[3]), .Y(ab_1__3_) );
  XOR3X2 U6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .C(ab_4__7_), .Y(SUMB_5__6_) );
  NAND2X1 U7 ( .A(ab_5__6_), .B(CARRYB_4__6_), .Y(n3) );
  NAND2X1 U8 ( .A(ab_5__6_), .B(ab_4__7_), .Y(n4) );
  NAND2X1 U9 ( .A(CARRYB_4__6_), .B(ab_4__7_), .Y(n5) );
  NAND3X1 U10 ( .A(n3), .B(n4), .C(n5), .Y(CARRYB_5__6_) );
  XOR2X1 U11 ( .A(ab_6__6_), .B(ab_5__7_), .Y(n6) );
  XOR2X1 U12 ( .A(n6), .B(CARRYB_5__6_), .Y(SUMB_6__6_) );
  NAND2X1 U13 ( .A(ab_6__6_), .B(ab_5__7_), .Y(n7) );
  NAND2X1 U14 ( .A(ab_6__6_), .B(CARRYB_5__6_), .Y(n8) );
  NAND2X1 U15 ( .A(ab_5__7_), .B(CARRYB_5__6_), .Y(n9) );
  NAND3X1 U16 ( .A(n7), .B(n8), .C(n9), .Y(CARRYB_6__6_) );
  INVX4 U17 ( .A(B[6]), .Y(n37) );
  NAND3X4 U18 ( .A(n21), .B(n19), .C(n20), .Y(CARRYB_7__3_) );
  AND2X1 U19 ( .A(A[10]), .B(B[6]), .Y(ab_10__6_) );
  AND2X1 U20 ( .A(A[9]), .B(B[6]), .Y(ab_9__6_) );
  AND2X2 U21 ( .A(A[2]), .B(B[6]), .Y(ab_2__6_) );
  CLKINVX2 U22 ( .A(n38), .Y(n10) );
  INVX2 U23 ( .A(n10), .Y(n11) );
  INVXL U24 ( .A(n10), .Y(n12) );
  NAND2X1 U25 ( .A(ab_7__3_), .B(SUMB_6__4_), .Y(n20) );
  XOR2X2 U26 ( .A(CARRYB_9__5_), .B(n22), .Y(SUMB_10__5_) );
  XOR2X2 U27 ( .A(SUMB_6__4_), .B(n18), .Y(SUMB_7__3_) );
  NAND3X2 U28 ( .A(n25), .B(n23), .C(n24), .Y(CARRYB_10__5_) );
  XOR2X1 U29 ( .A(CARRYB_16__3_), .B(SUMB_16__4_), .Y(A1_18_) );
  NAND2X1 U30 ( .A(ab_0__7_), .B(ab_1__6_), .Y(n33) );
  NOR2X1 U31 ( .A(n42), .B(n34), .Y(ab_0__7_) );
  AND2X2 U32 ( .A(A[5]), .B(B[3]), .Y(ab_5__3_) );
  XOR2X2 U33 ( .A(CARRYB_16__2_), .B(SUMB_16__3_), .Y(A1_17_) );
  INVX1 U34 ( .A(B[5]), .Y(n38) );
  AND2X2 U36 ( .A(ab_0__5_), .B(ab_1__4_), .Y(n14) );
  AND2X2 U37 ( .A(ab_0__6_), .B(ab_1__5_), .Y(n15) );
  AND2X2 U38 ( .A(ab_0__2_), .B(n43), .Y(n16) );
  AND2X1 U39 ( .A(CARRYB_16__2_), .B(SUMB_16__3_), .Y(n27) );
  CLKINVX2 U40 ( .A(n36), .Y(n43) );
  XOR2X2 U41 ( .A(ab_1__5_), .B(ab_0__6_), .Y(SUMB_1__5_) );
  AND2X2 U42 ( .A(A[3]), .B(B[0]), .Y(ab_3__0_) );
  XOR2X4 U43 ( .A(SUMB_9__6_), .B(ab_10__5_), .Y(n22) );
  INVX2 U44 ( .A(n33), .Y(CARRYB_1__6_) );
  NAND2XL U45 ( .A(ab_0__3_), .B(ab_1__2_), .Y(n32) );
  NOR2X2 U46 ( .A(n39), .B(n34), .Y(ab_0__4_) );
  AND2X1 U47 ( .A(A[1]), .B(B[5]), .Y(ab_1__5_) );
  NAND2X1 U48 ( .A(A[1]), .B(B[1]), .Y(n36) );
  NOR2X1 U49 ( .A(n36), .B(n35), .Y(CARRYB_1__0_) );
  AND2X2 U50 ( .A(A[2]), .B(B[2]), .Y(ab_2__2_) );
  XOR2X2 U51 ( .A(n43), .B(ab_0__2_), .Y(SUMB_1__1_) );
  AND2X2 U52 ( .A(A[2]), .B(B[3]), .Y(ab_2__3_) );
  AND2X2 U53 ( .A(A[3]), .B(B[3]), .Y(ab_3__3_) );
  INVX2 U54 ( .A(B[7]), .Y(n42) );
  AND2X2 U55 ( .A(CARRYB_16__1_), .B(SUMB_16__2_), .Y(n26) );
  INVX4 U56 ( .A(A[0]), .Y(n34) );
  NAND2X1 U57 ( .A(ab_7__3_), .B(CARRYB_6__3_), .Y(n21) );
  NOR2X2 U58 ( .A(n37), .B(n34), .Y(ab_0__6_) );
  INVX2 U59 ( .A(B[4]), .Y(n39) );
  NAND2X1 U60 ( .A(CARRYB_6__3_), .B(SUMB_6__4_), .Y(n19) );
  XOR2X4 U61 ( .A(CARRYB_6__3_), .B(ab_7__3_), .Y(n18) );
  AND2X1 U62 ( .A(A[7]), .B(B[3]), .Y(ab_7__3_) );
  NAND2X1 U63 ( .A(SUMB_9__6_), .B(CARRYB_9__5_), .Y(n23) );
  NAND2X1 U64 ( .A(ab_10__5_), .B(CARRYB_9__5_), .Y(n24) );
  NAND2XL U65 ( .A(ab_10__5_), .B(SUMB_9__6_), .Y(n25) );
  CLKINVX2 U66 ( .A(B[2]), .Y(n41) );
  INVX2 U67 ( .A(B[3]), .Y(n40) );
  XOR2X1 U68 ( .A(CARRYB_16__0_), .B(SUMB_16__1_), .Y(A1_15_) );
  AND2X2 U69 ( .A(A[2]), .B(B[5]), .Y(ab_2__5_) );
  AND2X1 U70 ( .A(A[7]), .B(B[6]), .Y(ab_7__6_) );
  AND2X1 U71 ( .A(A[6]), .B(B[6]), .Y(ab_6__6_) );
  AND2X1 U72 ( .A(A[5]), .B(B[6]), .Y(ab_5__6_) );
  AND2X1 U73 ( .A(A[8]), .B(B[6]), .Y(ab_8__6_) );
  AND2X1 U74 ( .A(A[4]), .B(B[6]), .Y(ab_4__6_) );
  XOR2X1 U75 ( .A(ab_1__6_), .B(ab_0__7_), .Y(SUMB_1__6_) );
  XOR2X2 U76 ( .A(CARRYB_16__1_), .B(SUMB_16__2_), .Y(A1_16_) );
  AND2X1 U77 ( .A(A[7]), .B(B[0]), .Y(ab_7__0_) );
  AND2X1 U78 ( .A(A[6]), .B(B[0]), .Y(ab_6__0_) );
  AND2X1 U79 ( .A(A[9]), .B(B[0]), .Y(ab_9__0_) );
  AND2X1 U80 ( .A(A[10]), .B(B[1]), .Y(ab_10__1_) );
  AND2X1 U81 ( .A(A[9]), .B(B[1]), .Y(ab_9__1_) );
  AND2X1 U82 ( .A(A[8]), .B(B[1]), .Y(ab_8__1_) );
  AND2X1 U83 ( .A(A[10]), .B(B[0]), .Y(ab_10__0_) );
  AND2X1 U84 ( .A(A[7]), .B(B[1]), .Y(ab_7__1_) );
  AND2X1 U85 ( .A(A[6]), .B(B[1]), .Y(ab_6__1_) );
  AND2X1 U86 ( .A(A[6]), .B(B[3]), .Y(ab_6__3_) );
  AND2X1 U87 ( .A(A[8]), .B(B[3]), .Y(ab_8__3_) );
  AND2X1 U88 ( .A(A[7]), .B(B[4]), .Y(ab_7__4_) );
  AND2X1 U89 ( .A(A[10]), .B(B[3]), .Y(ab_10__3_) );
  AND2X1 U90 ( .A(A[9]), .B(B[3]), .Y(ab_9__3_) );
  AND2X1 U91 ( .A(A[9]), .B(B[4]), .Y(ab_9__4_) );
  AND2X1 U92 ( .A(A[8]), .B(B[4]), .Y(ab_8__4_) );
  AND2X1 U93 ( .A(A[10]), .B(B[4]), .Y(ab_10__4_) );
  XOR2X1 U94 ( .A(CARRYB_16__4_), .B(SUMB_16__5_), .Y(A1_19_) );
  AND2X2 U95 ( .A(CARRYB_16__3_), .B(SUMB_16__4_), .Y(n28) );
  AND2X2 U96 ( .A(CARRYB_16__0_), .B(SUMB_16__1_), .Y(n29) );
  AND2X2 U97 ( .A(CARRYB_16__4_), .B(SUMB_16__5_), .Y(n30) );
  INVX1 U98 ( .A(B[0]), .Y(n51) );
  NOR2XL U99 ( .A(n44), .B(n41), .Y(ab_16__2_) );
  NOR2X1 U100 ( .A(n44), .B(n40), .Y(ab_16__3_) );
  NOR2X1 U101 ( .A(n44), .B(n12), .Y(ab_16__5_) );
  AND2X1 U102 ( .A(A[10]), .B(B[2]), .Y(ab_10__2_) );
  AND2X1 U103 ( .A(A[9]), .B(B[2]), .Y(ab_9__2_) );
  AND2X1 U104 ( .A(A[8]), .B(B[2]), .Y(ab_8__2_) );
  AND2X1 U105 ( .A(A[7]), .B(B[2]), .Y(ab_7__2_) );
  AND2X1 U106 ( .A(A[6]), .B(B[2]), .Y(ab_6__2_) );
  AND2X1 U107 ( .A(A[5]), .B(B[2]), .Y(ab_5__2_) );
  AND2X1 U108 ( .A(A[4]), .B(B[2]), .Y(ab_4__2_) );
  AND2X2 U109 ( .A(A[5]), .B(B[1]), .Y(ab_5__1_) );
  AND2X2 U110 ( .A(A[8]), .B(B[0]), .Y(ab_8__0_) );
  AND2X2 U111 ( .A(A[4]), .B(B[1]), .Y(ab_4__1_) );
  AND2X2 U112 ( .A(A[5]), .B(B[0]), .Y(ab_5__0_) );
  AND2X2 U113 ( .A(A[4]), .B(B[0]), .Y(ab_4__0_) );
  XOR2X1 U114 ( .A(CARRYB_16__5_), .B(SUMB_16__6_), .Y(A1_20_) );
  XOR2X1 U115 ( .A(CARRYB_16__6_), .B(ab_16__7_), .Y(A1_21_) );
  AND2X2 U116 ( .A(CARRYB_16__5_), .B(SUMB_16__6_), .Y(n31) );
  NOR2X1 U117 ( .A(n44), .B(n42), .Y(ab_16__7_) );
  INVX1 U118 ( .A(B[1]), .Y(n50) );
  NOR2X2 U119 ( .A(n40), .B(n34), .Y(ab_0__3_) );
  NOR2X2 U120 ( .A(n11), .B(n34), .Y(ab_0__5_) );
  NOR2XL U121 ( .A(n45), .B(n42), .Y(ab_15__7_) );
  AND2X1 U122 ( .A(A[1]), .B(B[2]), .Y(ab_1__2_) );
  NOR2XL U123 ( .A(n45), .B(n41), .Y(ab_15__2_) );
  NOR2XL U124 ( .A(n47), .B(n41), .Y(ab_13__2_) );
  NOR2XL U125 ( .A(n48), .B(n41), .Y(ab_12__2_) );
  NOR2XL U126 ( .A(n49), .B(n41), .Y(ab_11__2_) );
  NOR2XL U127 ( .A(n45), .B(n40), .Y(ab_15__3_) );
  NOR2XL U128 ( .A(n46), .B(n40), .Y(ab_14__3_) );
  NOR2XL U129 ( .A(n48), .B(n40), .Y(ab_12__3_) );
  NOR2XL U130 ( .A(n49), .B(n40), .Y(ab_11__3_) );
  AND2X2 U131 ( .A(A[6]), .B(B[4]), .Y(ab_6__4_) );
  AND2X2 U132 ( .A(A[5]), .B(B[4]), .Y(ab_5__4_) );
  AND2X1 U133 ( .A(A[10]), .B(B[5]), .Y(ab_10__5_) );
  NOR2XL U134 ( .A(n47), .B(n12), .Y(ab_13__5_) );
  AND2X1 U135 ( .A(A[9]), .B(B[5]), .Y(ab_9__5_) );
  NOR2XL U136 ( .A(n48), .B(n12), .Y(ab_12__5_) );
  AND2X1 U137 ( .A(A[4]), .B(B[3]), .Y(ab_4__3_) );
  AND2X1 U138 ( .A(A[8]), .B(B[5]), .Y(ab_8__5_) );
  AND2X1 U139 ( .A(A[7]), .B(B[5]), .Y(ab_7__5_) );
  AND2X2 U140 ( .A(A[4]), .B(B[4]), .Y(ab_4__4_) );
  AND2X1 U141 ( .A(A[6]), .B(B[5]), .Y(ab_6__5_) );
  AND2X1 U142 ( .A(A[5]), .B(B[5]), .Y(ab_5__5_) );
  AND2X1 U143 ( .A(A[4]), .B(B[5]), .Y(ab_4__5_) );
  AND2X1 U144 ( .A(A[3]), .B(B[2]), .Y(ab_3__2_) );
  NOR2XL U145 ( .A(n49), .B(n42), .Y(ab_11__7_) );
  AND2X1 U146 ( .A(A[3]), .B(B[5]), .Y(ab_3__5_) );
  AND2X1 U147 ( .A(A[3]), .B(B[1]), .Y(ab_3__1_) );
  AND2X1 U148 ( .A(A[3]), .B(B[6]), .Y(ab_3__6_) );
  XOR2X1 U149 ( .A(ab_1__4_), .B(ab_0__5_), .Y(SUMB_1__4_) );
  XOR2X1 U150 ( .A(ab_1__3_), .B(ab_0__4_), .Y(SUMB_1__3_) );
  XOR2X1 U151 ( .A(ab_1__2_), .B(ab_0__3_), .Y(SUMB_1__2_) );
  AND2X2 U152 ( .A(A[2]), .B(B[1]), .Y(ab_2__1_) );
  AND2X2 U153 ( .A(A[2]), .B(B[4]), .Y(ab_2__4_) );
  NOR2XL U154 ( .A(n46), .B(n41), .Y(ab_14__2_) );
  NOR2XL U155 ( .A(n47), .B(n40), .Y(ab_13__3_) );
  NOR2XL U156 ( .A(n49), .B(n12), .Y(ab_11__5_) );
  NOR2XL U157 ( .A(n46), .B(n12), .Y(ab_14__5_) );
  NOR2XL U158 ( .A(n45), .B(n12), .Y(ab_15__5_) );
  AND2X2 U159 ( .A(A[3]), .B(B[4]), .Y(ab_3__4_) );
  NOR2XL U160 ( .A(n48), .B(n42), .Y(ab_12__7_) );
  NOR2XL U161 ( .A(n47), .B(n42), .Y(ab_13__7_) );
  NOR2XL U162 ( .A(n46), .B(n42), .Y(ab_14__7_) );
  AND2X2 U163 ( .A(A[2]), .B(B[0]), .Y(ab_2__0_) );
  INVX1 U164 ( .A(A[16]), .Y(n44) );
  NAND2XL U165 ( .A(A[0]), .B(B[0]), .Y(n35) );
  INVX1 U166 ( .A(A[11]), .Y(n49) );
  INVX1 U167 ( .A(A[12]), .Y(n48) );
  INVX1 U168 ( .A(A[13]), .Y(n47) );
  INVX1 U169 ( .A(A[14]), .Y(n46) );
  INVX1 U170 ( .A(A[15]), .Y(n45) );
  AND2X2 U171 ( .A(A[1]), .B(B[4]), .Y(ab_1__4_) );
  NOR2XL U172 ( .A(n44), .B(n39), .Y(ab_16__4_) );
  NOR2XL U173 ( .A(n45), .B(n39), .Y(ab_15__4_) );
  NOR2XL U174 ( .A(n46), .B(n39), .Y(ab_14__4_) );
  NOR2XL U175 ( .A(n47), .B(n39), .Y(ab_13__4_) );
  NOR2XL U176 ( .A(n48), .B(n39), .Y(ab_12__4_) );
  NOR2XL U177 ( .A(n49), .B(n39), .Y(ab_11__4_) );
  NOR2XL U178 ( .A(n44), .B(n37), .Y(ab_16__6_) );
  NOR2XL U179 ( .A(n45), .B(n37), .Y(ab_15__6_) );
  NOR2XL U180 ( .A(n46), .B(n37), .Y(ab_14__6_) );
  NOR2XL U181 ( .A(n47), .B(n37), .Y(ab_13__6_) );
  NOR2XL U182 ( .A(n48), .B(n37), .Y(ab_12__6_) );
  NOR2XL U183 ( .A(n49), .B(n37), .Y(ab_11__6_) );
  AND2X1 U184 ( .A(A[10]), .B(B[7]), .Y(ab_10__7_) );
  AND2X1 U185 ( .A(A[9]), .B(B[7]), .Y(ab_9__7_) );
  AND2X1 U186 ( .A(A[8]), .B(B[7]), .Y(ab_8__7_) );
  AND2X1 U187 ( .A(A[7]), .B(B[7]), .Y(ab_7__7_) );
  AND2X1 U188 ( .A(A[6]), .B(B[7]), .Y(ab_6__7_) );
  AND2X1 U189 ( .A(A[5]), .B(B[7]), .Y(ab_5__7_) );
  AND2X1 U190 ( .A(A[4]), .B(B[7]), .Y(ab_4__7_) );
  AND2X1 U191 ( .A(A[3]), .B(B[7]), .Y(ab_3__7_) );
  AND2X1 U192 ( .A(A[2]), .B(B[7]), .Y(ab_2__7_) );
  AND2X1 U193 ( .A(A[1]), .B(B[7]), .Y(ab_1__7_) );
  NOR2X4 U194 ( .A(n41), .B(n34), .Y(ab_0__2_) );
  NOR2X1 U196 ( .A(n50), .B(n44), .Y(ab_16__1_) );
  NOR2X1 U197 ( .A(n51), .B(n44), .Y(ab_16__0_) );
  NOR2X1 U198 ( .A(n50), .B(n45), .Y(ab_15__1_) );
  NOR2X1 U199 ( .A(n51), .B(n45), .Y(ab_15__0_) );
  NOR2X1 U200 ( .A(n50), .B(n46), .Y(ab_14__1_) );
  NOR2X1 U201 ( .A(n51), .B(n46), .Y(ab_14__0_) );
  NOR2X1 U202 ( .A(n50), .B(n47), .Y(ab_13__1_) );
  NOR2X1 U203 ( .A(n51), .B(n47), .Y(ab_13__0_) );
  NOR2X1 U204 ( .A(n50), .B(n48), .Y(ab_12__1_) );
  NOR2X1 U205 ( .A(n51), .B(n48), .Y(ab_12__0_) );
  NOR2X1 U206 ( .A(n50), .B(n49), .Y(ab_11__1_) );
  NOR2X1 U207 ( .A(n51), .B(n49), .Y(ab_11__0_) );
endmodule


module multi16_0 ( in_17bit, in_8bit, out );
  input [16:0] in_17bit;
  input [7:0] in_8bit;
  output [16:0] out;
  wire   N18, N19, N20, N21, N32, N33, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n55, n56, n57, n58, n59, n60, n61, n63, n64, n65, n66, n67, n68,
         n69, n71, n72, n73, n74, n75, n76, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n126, n127, n128, n129;
  wire   [16:1] in_17bit_b;
  wire   [6:0] in_8bit_b;
  wire   [23:8] mul;
  wire   [16:12] sub_add_52_b0_carry;

  multi16_0_DW02_mult_0 mult_55 ( .A({in_17bit_b, in_17bit[0]}), .B({n8, 
        in_8bit_b}), .PRODUCT_23_(mul[23]), .PRODUCT_22_(mul[22]), 
        .PRODUCT_21_(mul[21]), .PRODUCT_20_(mul[20]), .PRODUCT_19_(mul[19]), 
        .PRODUCT_18_(mul[18]), .PRODUCT_17_(mul[17]), .PRODUCT_16_(mul[16]), 
        .PRODUCT_15_(mul[15]), .PRODUCT_14_(mul[14]), .PRODUCT_13_(mul[13]), 
        .PRODUCT_12_(mul[12]), .PRODUCT_11_(mul[11]), .PRODUCT_10_(mul[10]), 
        .PRODUCT_9_(mul[9]), .PRODUCT_8_(mul[8]), .PRODUCT_7_(N32) );
  INVX2 U2 ( .A(n113), .Y(n116) );
  NAND2X2 U3 ( .A(n4), .B(n5), .Y(in_8bit_b[6]) );
  CLKINVX3 U4 ( .A(n6), .Y(n7) );
  INVX1 U5 ( .A(n40), .Y(n6) );
  CLKINVX3 U6 ( .A(n98), .Y(n100) );
  NAND3BX2 U7 ( .AN(mul[20]), .B(n109), .C(n108), .Y(n110) );
  OAI21X2 U8 ( .A0(mul[19]), .A1(n106), .B0(n129), .Y(n107) );
  AND2X2 U9 ( .A(n37), .B(n39), .Y(n1) );
  NOR2X4 U10 ( .A(n1), .B(n25), .Y(n38) );
  INVX3 U11 ( .A(n36), .Y(n39) );
  INVX8 U12 ( .A(in_8bit[7]), .Y(n25) );
  XNOR2X4 U13 ( .A(n38), .B(n7), .Y(in_8bit_b[5]) );
  NAND2X2 U14 ( .A(in_8bit[6]), .B(n3), .Y(n4) );
  NAND2X2 U15 ( .A(n2), .B(n22), .Y(n5) );
  INVXL U16 ( .A(in_8bit[6]), .Y(n2) );
  CLKINVX4 U17 ( .A(n22), .Y(n3) );
  NOR2XL U18 ( .A(in_17bit[1]), .B(in_17bit[0]), .Y(n43) );
  XOR2X2 U19 ( .A(mul[19]), .B(n105), .Y(out[12]) );
  NAND4BX4 U20 ( .AN(in_8bit[3]), .B(n7), .C(n39), .D(n28), .Y(n41) );
  NAND3BX2 U21 ( .AN(in_8bit[1]), .B(n33), .C(n27), .Y(n36) );
  CLKINVX1 U22 ( .A(in_8bit[5]), .Y(n40) );
  INVX4 U23 ( .A(in_17bit[16]), .Y(n29) );
  NAND3XL U24 ( .A(in_17bit[0]), .B(in_17bit[16]), .C(in_17bit[1]), .Y(n44) );
  INVXL U25 ( .A(n107), .Y(n10) );
  INVX4 U26 ( .A(mul[22]), .Y(n115) );
  XNOR2X1 U27 ( .A(in_8bit[3]), .B(n34), .Y(in_8bit_b[3]) );
  NAND2XL U28 ( .A(n36), .B(n24), .Y(n34) );
  INVX1 U29 ( .A(n92), .Y(n94) );
  NOR2X1 U30 ( .A(n30), .B(n47), .Y(n17) );
  INVX1 U31 ( .A(n126), .Y(in_8bit_b[0]) );
  NAND2X2 U32 ( .A(n11), .B(n12), .Y(out[13]) );
  NAND2X1 U33 ( .A(n9), .B(n10), .Y(n12) );
  INVX2 U34 ( .A(n110), .Y(n112) );
  NOR2X2 U35 ( .A(in_17bit[1]), .B(in_17bit[0]), .Y(n23) );
  INVX1 U36 ( .A(n46), .Y(n47) );
  NAND2BX1 U37 ( .AN(in_17bit[2]), .B(n23), .Y(n46) );
  NOR2X1 U38 ( .A(n14), .B(n94), .Y(n93) );
  INVX1 U39 ( .A(n95), .Y(n97) );
  NAND2BX1 U40 ( .AN(mul[14]), .B(n94), .Y(n95) );
  NAND2BX1 U41 ( .AN(mul[15]), .B(n97), .Y(n98) );
  INVX1 U42 ( .A(n90), .Y(n91) );
  NAND2BX1 U43 ( .AN(mul[12]), .B(n89), .Y(n90) );
  INVX1 U44 ( .A(in_8bit[0]), .Y(n27) );
  NAND2BX2 U45 ( .AN(mul[18]), .B(n20), .Y(n106) );
  XOR2X1 U46 ( .A(mul[16]), .B(n99), .Y(out[9]) );
  NOR2X1 U47 ( .A(n14), .B(n100), .Y(n99) );
  XOR2X2 U48 ( .A(mul[18]), .B(n104), .Y(out[11]) );
  NOR2X2 U49 ( .A(n14), .B(n20), .Y(n104) );
  XOR2X1 U50 ( .A(mul[17]), .B(n102), .Y(out[10]) );
  NOR2X1 U51 ( .A(n14), .B(n103), .Y(n102) );
  NOR2X2 U52 ( .A(n14), .B(n112), .Y(n111) );
  NAND2BX2 U53 ( .AN(mul[21]), .B(n112), .Y(n113) );
  INVX4 U54 ( .A(n25), .Y(n24) );
  INVX1 U55 ( .A(in_17bit[16]), .Y(n30) );
  NOR3X2 U56 ( .A(in_8bit[6]), .B(n25), .C(n41), .Y(n8) );
  INVX1 U57 ( .A(mul[19]), .Y(n108) );
  XOR2X2 U58 ( .A(mul[21]), .B(n111), .Y(out[14]) );
  XOR2X1 U59 ( .A(mul[23]), .B(n117), .Y(out[16]) );
  AOI21X1 U60 ( .A0(n116), .A1(n115), .B0(n14), .Y(n117) );
  XOR2X4 U61 ( .A(in_17bit[2]), .B(n45), .Y(in_17bit_b[2]) );
  OAI21X1 U62 ( .A0(in_8bit[3]), .A1(n36), .B0(n24), .Y(n35) );
  AND2X4 U63 ( .A(n41), .B(n24), .Y(n22) );
  CLKINVX8 U64 ( .A(n101), .Y(n103) );
  XOR2X2 U65 ( .A(n17), .B(in_17bit[3]), .Y(in_17bit_b[3]) );
  INVX2 U66 ( .A(n103), .Y(n21) );
  INVX4 U67 ( .A(n106), .Y(n109) );
  NAND2BX1 U68 ( .AN(in_17bit[3]), .B(n47), .Y(n49) );
  NOR3BX2 U69 ( .AN(n44), .B(n43), .C(n42), .Y(in_17bit_b[1]) );
  NOR2X4 U70 ( .A(mul[17]), .B(n21), .Y(n20) );
  NOR2X4 U71 ( .A(n29), .B(n23), .Y(n45) );
  NAND2BX4 U72 ( .AN(mul[16]), .B(n100), .Y(n101) );
  XNOR2X2 U73 ( .A(n31), .B(n16), .Y(in_8bit_b[1]) );
  AND2X2 U74 ( .A(n26), .B(n24), .Y(n16) );
  XOR2X2 U75 ( .A(n35), .B(n28), .Y(in_8bit_b[4]) );
  NAND2XL U76 ( .A(mul[20]), .B(n107), .Y(n11) );
  INVXL U77 ( .A(mul[20]), .Y(n9) );
  INVXL U78 ( .A(in_8bit[1]), .Y(n31) );
  INVXL U79 ( .A(in_8bit[4]), .Y(n28) );
  NAND2BX2 U80 ( .AN(mul[13]), .B(n91), .Y(n92) );
  OR2X2 U81 ( .A(n14), .B(n91), .Y(n13) );
  XNOR2X1 U82 ( .A(mul[13]), .B(n13), .Y(out[6]) );
  XNOR2X1 U83 ( .A(n52), .B(n53), .Y(in_17bit_b[5]) );
  NAND2BXL U84 ( .AN(mul[8]), .B(n119), .Y(n78) );
  INVXL U85 ( .A(n27), .Y(n26) );
  NOR2XL U86 ( .A(n14), .B(n80), .Y(n79) );
  AOI22XL U87 ( .A0(n26), .A1(n24), .B0(n26), .B1(n25), .Y(n126) );
  XNOR2XL U88 ( .A(in_17bit[16]), .B(n24), .Y(n14) );
  AND2X2 U89 ( .A(n51), .B(n50), .Y(n15) );
  NOR2XL U90 ( .A(n30), .B(n61), .Y(n59) );
  NAND2XL U91 ( .A(n56), .B(in_17bit[16]), .Y(n55) );
  NAND2XL U92 ( .A(n15), .B(n53), .Y(n56) );
  NAND2BXL U93 ( .AN(n56), .B(n57), .Y(n58) );
  NAND2XL U94 ( .A(n72), .B(in_17bit[16]), .Y(n71) );
  NAND2XL U95 ( .A(n64), .B(in_17bit[16]), .Y(n63) );
  NAND2XL U96 ( .A(n61), .B(n60), .Y(n64) );
  INVXL U97 ( .A(n76), .Y(sub_add_52_b0_carry[12]) );
  NAND2XL U98 ( .A(n69), .B(n68), .Y(n72) );
  NAND2BXL U99 ( .AN(n64), .B(n65), .Y(n66) );
  AND2X1 U100 ( .A(N21), .B(in_17bit[16]), .Y(in_17bit_b[16]) );
  INVXL U101 ( .A(in_17bit[4]), .Y(n50) );
  INVXL U102 ( .A(in_17bit[5]), .Y(n53) );
  INVXL U103 ( .A(in_17bit[6]), .Y(n57) );
  MX2X1 U104 ( .A(in_17bit[11]), .B(n18), .S0(in_17bit[16]), .Y(in_17bit_b[11]) );
  XNOR2X1 U105 ( .A(n74), .B(n120), .Y(n18) );
  MX2X1 U106 ( .A(in_17bit[12]), .B(n19), .S0(in_17bit[16]), .Y(in_17bit_b[12]) );
  XNOR2X1 U107 ( .A(n76), .B(n121), .Y(n19) );
  MX2X1 U108 ( .A(in_17bit[13]), .B(N18), .S0(in_17bit[16]), .Y(in_17bit_b[13]) );
  MX2X1 U109 ( .A(in_17bit[14]), .B(N19), .S0(in_17bit[16]), .Y(in_17bit_b[14]) );
  MX2X1 U110 ( .A(in_17bit[15]), .B(N20), .S0(in_17bit[16]), .Y(in_17bit_b[15]) );
  INVXL U111 ( .A(in_17bit[7]), .Y(n60) );
  INVXL U112 ( .A(in_17bit[8]), .Y(n65) );
  INVX1 U113 ( .A(n84), .Y(n86) );
  NAND2BX1 U114 ( .AN(mul[10]), .B(n83), .Y(n84) );
  INVX1 U115 ( .A(n78), .Y(n80) );
  INVX1 U116 ( .A(n81), .Y(n83) );
  NAND2BX1 U117 ( .AN(mul[9]), .B(n80), .Y(n81) );
  INVX1 U118 ( .A(N32), .Y(n119) );
  XOR2X1 U119 ( .A(mul[11]), .B(n85), .Y(out[4]) );
  NOR2X1 U120 ( .A(n14), .B(n86), .Y(n85) );
  XOR2X1 U121 ( .A(mul[12]), .B(n88), .Y(out[5]) );
  NOR2X1 U122 ( .A(n14), .B(n89), .Y(n88) );
  XOR2X1 U123 ( .A(mul[15]), .B(n96), .Y(out[8]) );
  NOR2X1 U124 ( .A(n14), .B(n97), .Y(n96) );
  XOR2X1 U125 ( .A(mul[14]), .B(n93), .Y(out[7]) );
  XOR2X1 U126 ( .A(mul[10]), .B(n82), .Y(out[3]) );
  NOR2X1 U127 ( .A(n14), .B(n83), .Y(n82) );
  XOR2X1 U128 ( .A(mul[9]), .B(n79), .Y(out[2]) );
  INVX1 U129 ( .A(n87), .Y(n89) );
  NAND2BX1 U130 ( .AN(mul[11]), .B(n86), .Y(n87) );
  INVX1 U131 ( .A(n128), .Y(out[1]) );
  AOI22X1 U132 ( .A0(mul[8]), .A1(n14), .B0(N33), .B1(n129), .Y(n128) );
  INVX1 U133 ( .A(mul[8]), .Y(n118) );
  INVX1 U134 ( .A(n127), .Y(out[0]) );
  AOI22XL U135 ( .A0(N32), .A1(n14), .B0(N32), .B1(n129), .Y(n127) );
  INVXL U136 ( .A(n14), .Y(n129) );
  NOR2X1 U137 ( .A(n30), .B(n15), .Y(n52) );
  XNOR2X1 U138 ( .A(n59), .B(n60), .Y(in_17bit_b[7]) );
  XNOR2X1 U139 ( .A(n67), .B(n68), .Y(in_17bit_b[9]) );
  NOR2X1 U140 ( .A(n29), .B(n69), .Y(n67) );
  XOR2X1 U141 ( .A(n50), .B(n48), .Y(in_17bit_b[4]) );
  NAND2X1 U142 ( .A(n49), .B(in_17bit[16]), .Y(n48) );
  XOR2X1 U143 ( .A(n57), .B(n55), .Y(in_17bit_b[6]) );
  XOR2X1 U144 ( .A(n65), .B(n63), .Y(in_17bit_b[8]) );
  XOR2X1 U145 ( .A(n73), .B(n71), .Y(in_17bit_b[10]) );
  NAND2BX1 U146 ( .AN(n72), .B(n73), .Y(n74) );
  CLKINVX2 U147 ( .A(in_8bit[2]), .Y(n33) );
  INVX1 U148 ( .A(n49), .Y(n51) );
  INVX1 U149 ( .A(n58), .Y(n61) );
  INVX1 U150 ( .A(n66), .Y(n69) );
  NAND2X1 U151 ( .A(n120), .B(n75), .Y(n76) );
  INVX1 U152 ( .A(n74), .Y(n75) );
  NOR2X1 U153 ( .A(in_17bit[16]), .B(in_17bit[1]), .Y(n42) );
  INVX1 U154 ( .A(in_17bit[9]), .Y(n68) );
  INVX1 U155 ( .A(in_17bit[10]), .Y(n73) );
  INVX1 U156 ( .A(in_17bit[11]), .Y(n120) );
  INVX1 U157 ( .A(in_17bit[12]), .Y(n121) );
  INVX1 U158 ( .A(in_17bit[13]), .Y(n122) );
  INVX1 U159 ( .A(in_17bit[14]), .Y(n123) );
  INVX1 U160 ( .A(in_17bit[15]), .Y(n124) );
  NOR2XL U161 ( .A(in_8bit[4]), .B(in_8bit[3]), .Y(n37) );
  OAI2BB1X4 U162 ( .A0N(n27), .A1N(n31), .B0(n24), .Y(n32) );
  XOR2X4 U163 ( .A(n33), .B(n32), .Y(in_8bit_b[2]) );
  NOR2X4 U164 ( .A(n14), .B(n109), .Y(n105) );
  NOR2X4 U165 ( .A(n14), .B(n116), .Y(n114) );
  XNOR2X4 U166 ( .A(n114), .B(n115), .Y(out[15]) );
  XOR2X1 U167 ( .A(n118), .B(n119), .Y(N33) );
  XOR2X1 U168 ( .A(n29), .B(sub_add_52_b0_carry[16]), .Y(N21) );
  AND2X1 U169 ( .A(sub_add_52_b0_carry[15]), .B(n124), .Y(
        sub_add_52_b0_carry[16]) );
  XOR2X1 U170 ( .A(n124), .B(sub_add_52_b0_carry[15]), .Y(N20) );
  AND2X1 U171 ( .A(sub_add_52_b0_carry[14]), .B(n123), .Y(
        sub_add_52_b0_carry[15]) );
  XOR2X1 U172 ( .A(n123), .B(sub_add_52_b0_carry[14]), .Y(N19) );
  AND2X1 U173 ( .A(sub_add_52_b0_carry[13]), .B(n122), .Y(
        sub_add_52_b0_carry[14]) );
  XOR2X1 U174 ( .A(n122), .B(sub_add_52_b0_carry[13]), .Y(N18) );
  AND2X1 U175 ( .A(sub_add_52_b0_carry[12]), .B(n121), .Y(
        sub_add_52_b0_carry[13]) );
endmodule


module butterfly_DW01_sub_18 ( A, B, DIFF );
  input [16:0] A;
  input [16:0] B;
  output [16:0] DIFF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170;

  NAND2X2 U3 ( .A(n3), .B(n4), .Y(n64) );
  CLKINVX4 U4 ( .A(n88), .Y(n77) );
  NAND2BX2 U5 ( .AN(A[10]), .B(B[10]), .Y(n97) );
  NAND2X1 U6 ( .A(B[16]), .B(A[16]), .Y(n3) );
  NAND2X1 U7 ( .A(n1), .B(n2), .Y(n4) );
  INVX1 U8 ( .A(B[16]), .Y(n1) );
  INVX1 U9 ( .A(A[16]), .Y(n2) );
  NAND2X2 U10 ( .A(n115), .B(n6), .Y(n7) );
  NAND2X2 U11 ( .A(n5), .B(n116), .Y(n8) );
  NAND2X4 U12 ( .A(n7), .B(n8), .Y(DIFF[13]) );
  CLKINVX3 U13 ( .A(n115), .Y(n5) );
  INVX2 U14 ( .A(n116), .Y(n6) );
  NAND2X2 U15 ( .A(n97), .B(n129), .Y(n140) );
  NAND2BX4 U16 ( .AN(B[10]), .B(A[10]), .Y(n129) );
  NAND2X2 U17 ( .A(n88), .B(n76), .Y(n115) );
  INVX2 U18 ( .A(n82), .Y(n112) );
  CLKINVX3 U19 ( .A(n87), .Y(n113) );
  NAND3X2 U20 ( .A(n114), .B(n90), .C(n91), .Y(n118) );
  NAND2X2 U21 ( .A(n144), .B(n19), .Y(n14) );
  NAND2XL U22 ( .A(n21), .B(n20), .Y(n144) );
  NAND2X1 U23 ( .A(n78), .B(n87), .Y(n123) );
  NAND2X2 U24 ( .A(A[12]), .B(n135), .Y(n78) );
  INVX1 U25 ( .A(B[12]), .Y(n135) );
  NAND2X1 U26 ( .A(A[14]), .B(n107), .Y(n75) );
  INVX1 U27 ( .A(B[14]), .Y(n107) );
  NOR2X2 U28 ( .A(n16), .B(n17), .Y(n15) );
  INVXL U29 ( .A(n18), .Y(n16) );
  INVX2 U30 ( .A(A[14]), .Y(n106) );
  OAI21XL U31 ( .A0(n32), .A1(n33), .B0(n34), .Y(n28) );
  OAI21XL U32 ( .A0(n39), .A1(n40), .B0(n41), .Y(n35) );
  INVX1 U33 ( .A(n96), .Y(n17) );
  NAND2X1 U34 ( .A(A[9]), .B(n142), .Y(n18) );
  NAND2X1 U35 ( .A(A[8]), .B(n145), .Y(n19) );
  NAND2X1 U36 ( .A(B[7]), .B(n154), .Y(n23) );
  OAI21XL U37 ( .A0(n40), .A1(n85), .B0(n94), .Y(n21) );
  NAND2X2 U38 ( .A(B[12]), .B(n134), .Y(n87) );
  INVX2 U39 ( .A(A[12]), .Y(n134) );
  OAI21X1 U40 ( .A0(n141), .A1(n17), .B0(n18), .Y(n137) );
  INVX1 U41 ( .A(n14), .Y(n141) );
  XNOR2X1 U42 ( .A(n21), .B(n12), .Y(DIFF[8]) );
  NAND2X1 U43 ( .A(n19), .B(n20), .Y(n12) );
  INVX1 U44 ( .A(n120), .Y(n91) );
  NAND2BX2 U45 ( .AN(B[11]), .B(A[11]), .Y(n90) );
  NOR2BX1 U46 ( .AN(n79), .B(n68), .Y(n67) );
  AND2X2 U47 ( .A(n23), .B(n24), .Y(n9) );
  AND4X4 U48 ( .A(n87), .B(n88), .C(n71), .D(n72), .Y(n10) );
  NOR2XL U49 ( .A(n69), .B(n70), .Y(n68) );
  NAND3X1 U50 ( .A(n88), .B(n110), .C(n111), .Y(n109) );
  NOR2X1 U51 ( .A(n112), .B(n113), .Y(n111) );
  NAND2X2 U52 ( .A(B[9]), .B(n143), .Y(n96) );
  INVX4 U53 ( .A(A[15]), .Y(n102) );
  INVX3 U54 ( .A(n71), .Y(n105) );
  OAI21X2 U55 ( .A0(n77), .A1(n78), .B0(n76), .Y(n108) );
  NAND2X2 U56 ( .A(A[13]), .B(n121), .Y(n76) );
  NAND2X4 U57 ( .A(B[15]), .B(n102), .Y(n72) );
  NAND4X2 U58 ( .A(n80), .B(n81), .C(n82), .D(n10), .Y(n66) );
  NAND2X2 U59 ( .A(n127), .B(n90), .Y(n126) );
  NAND2X2 U60 ( .A(n120), .B(n82), .Y(n127) );
  NAND3X1 U61 ( .A(n86), .B(n82), .C(n10), .Y(n65) );
  INVX1 U62 ( .A(n75), .Y(n11) );
  NAND2X2 U63 ( .A(A[15]), .B(n103), .Y(n79) );
  NAND3X2 U64 ( .A(n65), .B(n66), .C(n67), .Y(n63) );
  INVX2 U65 ( .A(A[13]), .Y(n122) );
  INVXL U66 ( .A(A[10]), .Y(n132) );
  INVX2 U67 ( .A(n75), .Y(n101) );
  NAND2BXL U68 ( .AN(n83), .B(n92), .Y(n89) );
  INVX1 U69 ( .A(n137), .Y(n139) );
  INVX2 U70 ( .A(n129), .Y(n138) );
  INVXL U71 ( .A(B[5]), .Y(n153) );
  NAND2X1 U72 ( .A(n132), .B(B[10]), .Y(n130) );
  NAND2XL U73 ( .A(A[1]), .B(n167), .Y(n57) );
  INVX1 U74 ( .A(n42), .Y(n40) );
  NOR2X2 U75 ( .A(n112), .B(n114), .Y(n125) );
  INVX1 U76 ( .A(B[13]), .Y(n121) );
  NAND2X2 U77 ( .A(n79), .B(n72), .Y(n98) );
  NAND2XL U78 ( .A(n93), .B(n94), .Y(n92) );
  NOR2X1 U79 ( .A(n30), .B(n26), .Y(n29) );
  NAND4XL U80 ( .A(n45), .B(n38), .C(n31), .D(n23), .Y(n85) );
  OAI21XL U81 ( .A0(n25), .A1(n26), .B0(n27), .Y(n22) );
  NAND3XL U82 ( .A(n38), .B(n151), .C(n31), .Y(n148) );
  NAND2BX1 U83 ( .AN(n62), .B(n61), .Y(n58) );
  AOI21X2 U84 ( .A0(n97), .A1(n137), .B0(n138), .Y(n136) );
  NAND2X1 U85 ( .A(B[8]), .B(n146), .Y(n20) );
  INVX1 U86 ( .A(B[6]), .Y(n150) );
  INVX1 U87 ( .A(A[0]), .Y(n169) );
  NOR2X2 U88 ( .A(n112), .B(n113), .Y(n117) );
  NAND2BXL U89 ( .AN(n85), .B(n95), .Y(n93) );
  INVX2 U90 ( .A(n78), .Y(n119) );
  NAND2X2 U91 ( .A(B[13]), .B(n122), .Y(n88) );
  NAND3XL U92 ( .A(n114), .B(n90), .C(n91), .Y(n110) );
  NOR2X4 U93 ( .A(n125), .B(n126), .Y(n124) );
  NAND3XL U94 ( .A(n89), .B(n90), .C(n91), .Y(n86) );
  XOR2X2 U95 ( .A(n22), .B(n9), .Y(DIFF[7]) );
  NAND3XL U96 ( .A(n96), .B(n20), .C(n97), .Y(n83) );
  NAND2XL U97 ( .A(n23), .B(n147), .Y(n94) );
  NAND3BXL U98 ( .AN(n54), .B(n158), .C(n51), .Y(n84) );
  INVXL U99 ( .A(n55), .Y(n50) );
  NAND2XL U100 ( .A(n34), .B(n41), .Y(n151) );
  NAND2XL U101 ( .A(n61), .B(n62), .Y(DIFF[0]) );
  NOR2XL U102 ( .A(n60), .B(n13), .Y(n59) );
  NAND4X1 U103 ( .A(n20), .B(n21), .C(n96), .D(n133), .Y(n114) );
  NAND2X1 U104 ( .A(n128), .B(n129), .Y(n120) );
  NAND2BX4 U105 ( .AN(A[11]), .B(B[11]), .Y(n82) );
  NAND2X1 U106 ( .A(A[7]), .B(n149), .Y(n24) );
  NAND2XL U107 ( .A(B[2]), .B(n164), .Y(n48) );
  INVXL U108 ( .A(A[2]), .Y(n164) );
  INVXL U109 ( .A(B[4]), .Y(n152) );
  INVXL U110 ( .A(B[1]), .Y(n167) );
  INVXL U111 ( .A(B[3]), .Y(n162) );
  INVXL U112 ( .A(B[0]), .Y(n170) );
  NAND2XL U113 ( .A(B[0]), .B(n169), .Y(n62) );
  NAND2BX1 U114 ( .AN(n95), .B(n84), .Y(n42) );
  XOR2X1 U115 ( .A(n49), .B(n53), .Y(DIFF[2]) );
  NOR2X1 U116 ( .A(n50), .B(n54), .Y(n53) );
  XOR2X1 U117 ( .A(n35), .B(n36), .Y(DIFF[5]) );
  NOR2X1 U118 ( .A(n37), .B(n33), .Y(n36) );
  INVX1 U119 ( .A(n34), .Y(n37) );
  XOR2X1 U120 ( .A(n28), .B(n29), .Y(DIFF[6]) );
  INVX1 U121 ( .A(n27), .Y(n30) );
  INVX1 U122 ( .A(n28), .Y(n25) );
  XOR2X1 U123 ( .A(n42), .B(n43), .Y(DIFF[4]) );
  NOR2X1 U124 ( .A(n44), .B(n39), .Y(n43) );
  INVX1 U125 ( .A(n41), .Y(n44) );
  XOR2X1 U126 ( .A(n46), .B(n47), .Y(DIFF[3]) );
  AOI21X1 U127 ( .A0(n48), .A1(n49), .B0(n50), .Y(n47) );
  NAND2X1 U128 ( .A(n51), .B(n52), .Y(n46) );
  INVX1 U129 ( .A(n35), .Y(n32) );
  OAI21XL U130 ( .A0(n160), .A1(n161), .B0(n52), .Y(n95) );
  NOR2X1 U131 ( .A(n165), .B(n166), .Y(n160) );
  NAND2X1 U132 ( .A(n48), .B(n51), .Y(n161) );
  NAND2X1 U133 ( .A(n55), .B(n57), .Y(n166) );
  NOR2X1 U134 ( .A(n13), .B(n159), .Y(n158) );
  INVX1 U135 ( .A(n62), .Y(n159) );
  NOR2XL U136 ( .A(n84), .B(n85), .Y(n80) );
  INVX1 U137 ( .A(n83), .Y(n81) );
  NAND3X1 U138 ( .A(n148), .B(n27), .C(n24), .Y(n147) );
  INVX1 U139 ( .A(n48), .Y(n54) );
  NOR2X1 U140 ( .A(n13), .B(n61), .Y(n165) );
  INVX1 U141 ( .A(n31), .Y(n26) );
  INVX1 U142 ( .A(n38), .Y(n33) );
  INVX1 U143 ( .A(n45), .Y(n39) );
  NOR2X1 U144 ( .A(n73), .B(n74), .Y(n69) );
  XOR2X1 U145 ( .A(n58), .B(n59), .Y(DIFF[1]) );
  INVX1 U146 ( .A(n57), .Y(n60) );
  OAI21XL U147 ( .A0(n56), .A1(n13), .B0(n57), .Y(n49) );
  INVX1 U148 ( .A(n58), .Y(n56) );
  INVX1 U149 ( .A(A[8]), .Y(n146) );
  INVX1 U150 ( .A(A[9]), .Y(n143) );
  NOR2BX1 U151 ( .AN(B[1]), .B(A[1]), .Y(n13) );
  NAND2BXL U152 ( .AN(A[10]), .B(B[10]), .Y(n133) );
  INVX1 U153 ( .A(A[7]), .Y(n154) );
  INVX1 U154 ( .A(B[8]), .Y(n145) );
  NAND2X1 U155 ( .A(B[3]), .B(n163), .Y(n51) );
  INVX1 U156 ( .A(A[3]), .Y(n163) );
  NAND2X1 U157 ( .A(B[6]), .B(n155), .Y(n31) );
  INVX1 U158 ( .A(A[6]), .Y(n155) );
  NAND2X1 U159 ( .A(B[5]), .B(n156), .Y(n38) );
  INVX1 U160 ( .A(A[5]), .Y(n156) );
  INVX1 U161 ( .A(B[9]), .Y(n142) );
  NAND2X1 U162 ( .A(A[5]), .B(n153), .Y(n34) );
  NAND2X1 U163 ( .A(A[4]), .B(n152), .Y(n41) );
  NAND2X1 U164 ( .A(A[6]), .B(n150), .Y(n27) );
  NAND2X1 U165 ( .A(A[3]), .B(n162), .Y(n52) );
  NAND2X1 U166 ( .A(B[4]), .B(n157), .Y(n45) );
  INVX1 U167 ( .A(A[4]), .Y(n157) );
  NAND3X1 U168 ( .A(n96), .B(n130), .C(n131), .Y(n128) );
  NAND2XL U169 ( .A(n18), .B(n19), .Y(n131) );
  INVX1 U170 ( .A(B[15]), .Y(n103) );
  NAND2X1 U171 ( .A(A[2]), .B(n168), .Y(n55) );
  INVX1 U172 ( .A(B[2]), .Y(n168) );
  INVX1 U173 ( .A(B[7]), .Y(n149) );
  NAND2X1 U174 ( .A(A[0]), .B(n170), .Y(n61) );
  NAND2XL U175 ( .A(n75), .B(n76), .Y(n74) );
  AOI21X4 U176 ( .A0(n71), .A1(n100), .B0(n11), .Y(n99) );
  NAND2XL U177 ( .A(n71), .B(n72), .Y(n70) );
  NOR2XL U178 ( .A(n77), .B(n78), .Y(n73) );
  XOR2X4 U179 ( .A(n14), .B(n15), .Y(DIFF[9]) );
  XOR2X4 U180 ( .A(n63), .B(n64), .Y(DIFF[16]) );
  XOR2X4 U181 ( .A(n98), .B(n99), .Y(DIFF[15]) );
  XOR2X4 U182 ( .A(n100), .B(n104), .Y(DIFF[14]) );
  NOR2X4 U183 ( .A(n101), .B(n105), .Y(n104) );
  NAND2X4 U184 ( .A(B[14]), .B(n106), .Y(n71) );
  NAND2BX4 U185 ( .AN(n108), .B(n109), .Y(n100) );
  AOI21X4 U186 ( .A0(n117), .A1(n118), .B0(n119), .Y(n116) );
  XOR2X4 U187 ( .A(n123), .B(n124), .Y(DIFF[12]) );
  XOR3X4 U188 ( .A(B[11]), .B(A[11]), .C(n136), .Y(DIFF[11]) );
  XOR2X4 U189 ( .A(n139), .B(n140), .Y(DIFF[10]) );
endmodule


module butterfly_DW01_sub_26 ( A, B, DIFF );
  input [16:0] A;
  input [16:0] B;
  output [16:0] DIFF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163;

  NAND2X1 U3 ( .A(n101), .B(n2), .Y(n3) );
  NAND2X2 U4 ( .A(n1), .B(n102), .Y(n4) );
  NAND2X2 U5 ( .A(n3), .B(n4), .Y(DIFF[15]) );
  INVX1 U6 ( .A(n101), .Y(n1) );
  INVX1 U7 ( .A(n102), .Y(n2) );
  NAND2XL U8 ( .A(n105), .B(n93), .Y(n101) );
  NOR2X1 U9 ( .A(n94), .B(n103), .Y(n102) );
  NAND2X2 U10 ( .A(B[12]), .B(n118), .Y(n74) );
  NAND2X2 U11 ( .A(A[12]), .B(n117), .Y(n100) );
  INVX1 U12 ( .A(B[12]), .Y(n117) );
  NAND2X1 U13 ( .A(A[11]), .B(n130), .Y(n67) );
  NAND2BX2 U14 ( .AN(B[13]), .B(A[13]), .Y(n99) );
  INVX1 U15 ( .A(A[12]), .Y(n118) );
  NAND2BXL U16 ( .AN(A[14]), .B(B[14]), .Y(n97) );
  NAND2BX1 U17 ( .AN(A[14]), .B(B[14]), .Y(n75) );
  NAND2X2 U18 ( .A(B[10]), .B(n135), .Y(n85) );
  OAI21X2 U19 ( .A0(n110), .A1(n111), .B0(n99), .Y(n107) );
  AOI21X2 U20 ( .A0(n112), .A1(n74), .B0(n113), .Y(n110) );
  NAND3X1 U21 ( .A(n119), .B(n67), .C(n68), .Y(n112) );
  NAND4X1 U22 ( .A(n124), .B(n83), .C(n85), .D(n86), .Y(n119) );
  CLKINVX3 U23 ( .A(n100), .Y(n113) );
  NOR2BX1 U24 ( .AN(n90), .B(n91), .Y(n56) );
  AOI21X1 U25 ( .A0(n92), .A1(n93), .B0(n94), .Y(n91) );
  NAND3BX1 U26 ( .AN(n59), .B(n60), .C(n61), .Y(n58) );
  NOR2X1 U27 ( .A(n106), .B(n109), .Y(n108) );
  INVX1 U28 ( .A(n93), .Y(n109) );
  XNOR2X1 U29 ( .A(n55), .B(n6), .Y(DIFF[16]) );
  XOR2X1 U30 ( .A(B[16]), .B(A[16]), .Y(n6) );
  NAND3X1 U31 ( .A(n56), .B(n57), .C(n58), .Y(n55) );
  NAND2BX2 U32 ( .AN(A[13]), .B(B[13]), .Y(n73) );
  NAND3X1 U33 ( .A(n95), .B(n96), .C(n97), .Y(n92) );
  NAND2X1 U34 ( .A(n99), .B(n100), .Y(n95) );
  NAND3XL U35 ( .A(n73), .B(n74), .C(n75), .Y(n59) );
  INVX1 U36 ( .A(n90), .Y(n103) );
  INVX2 U37 ( .A(n104), .Y(n94) );
  OAI21XL U38 ( .A0(n140), .A1(n72), .B0(n71), .Y(n13) );
  INVXL U39 ( .A(n71), .Y(n70) );
  NOR2XL U40 ( .A(n79), .B(n113), .Y(n116) );
  INVXL U41 ( .A(n72), .Y(n87) );
  AOI21XL U42 ( .A0(n87), .A1(n69), .B0(n70), .Y(n62) );
  INVXL U43 ( .A(n75), .Y(n106) );
  INVXL U44 ( .A(n74), .Y(n79) );
  INVXL U45 ( .A(n8), .Y(n136) );
  NOR2XL U46 ( .A(n10), .B(n11), .Y(n9) );
  INVXL U47 ( .A(n12), .Y(n10) );
  NAND2XL U48 ( .A(n23), .B(n141), .Y(n71) );
  NOR2XL U49 ( .A(n15), .B(n16), .Y(n14) );
  INVXL U50 ( .A(n17), .Y(n15) );
  INVXL U51 ( .A(n20), .Y(n26) );
  XNOR2X1 U52 ( .A(n37), .B(n5), .Y(DIFF[4]) );
  NAND2XL U53 ( .A(n38), .B(n36), .Y(n5) );
  AOI21XL U54 ( .A0(n20), .A1(n21), .B0(n22), .Y(n19) );
  NAND2XL U55 ( .A(n23), .B(n24), .Y(n18) );
  NOR2XL U56 ( .A(n33), .B(n29), .Y(n32) );
  INVXL U57 ( .A(n30), .Y(n33) );
  NAND2XL U58 ( .A(n35), .B(n36), .Y(n31) );
  NAND2XL U59 ( .A(n37), .B(n38), .Y(n35) );
  INVXL U60 ( .A(n27), .Y(n22) );
  NOR2XL U61 ( .A(n7), .B(n46), .Y(n45) );
  NAND2XL U62 ( .A(n43), .B(n44), .Y(n39) );
  AOI21XL U63 ( .A0(n41), .A1(n42), .B0(n7), .Y(n40) );
  NOR2XL U64 ( .A(n52), .B(n48), .Y(n51) );
  NAND2BX1 U65 ( .AN(B[15]), .B(A[15]), .Y(n90) );
  NAND2BX1 U66 ( .AN(A[15]), .B(B[15]), .Y(n104) );
  INVX1 U67 ( .A(B[11]), .Y(n130) );
  NAND2X1 U68 ( .A(A[10]), .B(n134), .Y(n122) );
  INVXL U69 ( .A(B[7]), .Y(n143) );
  NAND2XL U70 ( .A(B[9]), .B(n138), .Y(n83) );
  INVXL U71 ( .A(A[9]), .Y(n138) );
  NAND2XL U72 ( .A(B[8]), .B(n161), .Y(n84) );
  INVXL U73 ( .A(A[8]), .Y(n161) );
  INVXL U74 ( .A(A[15]), .Y(n78) );
  INVXL U75 ( .A(A[13]), .Y(n98) );
  NAND2XL U76 ( .A(B[5]), .B(n150), .Y(n34) );
  INVXL U77 ( .A(A[5]), .Y(n150) );
  INVXL U78 ( .A(B[6]), .Y(n144) );
  NAND2XL U79 ( .A(B[2]), .B(n160), .Y(n41) );
  NAND4XL U80 ( .A(n43), .B(n41), .C(n54), .D(n152), .Y(n89) );
  NAND2XL U81 ( .A(B[4]), .B(n151), .Y(n38) );
  INVXL U82 ( .A(B[1]), .Y(n158) );
  INVXL U83 ( .A(B[3]), .Y(n155) );
  INVX1 U84 ( .A(n13), .Y(n125) );
  INVX1 U85 ( .A(n37), .Y(n140) );
  XOR2X1 U86 ( .A(n112), .B(n116), .Y(DIFF[12]) );
  NAND2BX1 U87 ( .AN(n106), .B(n107), .Y(n105) );
  INVX1 U88 ( .A(n68), .Y(n65) );
  NAND4X1 U89 ( .A(n38), .B(n34), .C(n20), .D(n23), .Y(n72) );
  NOR2X1 U90 ( .A(n125), .B(n16), .Y(n124) );
  NAND4XL U91 ( .A(n83), .B(n84), .C(n85), .D(n86), .Y(n63) );
  OAI21XL U92 ( .A0(n136), .A1(n11), .B0(n12), .Y(n128) );
  INVX1 U93 ( .A(n73), .Y(n111) );
  NOR2X1 U94 ( .A(n80), .B(n81), .Y(n76) );
  NAND2X1 U95 ( .A(n87), .B(n88), .Y(n80) );
  OAI21XL U96 ( .A0(n16), .A1(n125), .B0(n17), .Y(n8) );
  XOR2X1 U97 ( .A(n114), .B(n115), .Y(DIFF[13]) );
  NAND2XL U98 ( .A(n73), .B(n99), .Y(n114) );
  AOI21XL U99 ( .A0(n112), .A1(n74), .B0(n113), .Y(n115) );
  INVX1 U100 ( .A(n84), .Y(n16) );
  NAND3X1 U101 ( .A(n142), .B(n27), .C(n24), .Y(n141) );
  NAND3X1 U102 ( .A(n34), .B(n145), .C(n20), .Y(n142) );
  OAI21XL U103 ( .A0(n62), .A1(n63), .B0(n64), .Y(n60) );
  NOR2X1 U104 ( .A(n65), .B(n66), .Y(n64) );
  NAND2X2 U105 ( .A(n121), .B(n122), .Y(n120) );
  NAND3X1 U106 ( .A(n123), .B(n83), .C(n85), .Y(n121) );
  NAND2X1 U107 ( .A(n12), .B(n17), .Y(n123) );
  INVX1 U108 ( .A(n83), .Y(n11) );
  NAND2XL U109 ( .A(B[13]), .B(n98), .Y(n96) );
  INVX1 U110 ( .A(n122), .Y(n129) );
  XOR2X1 U111 ( .A(n128), .B(n132), .Y(DIFF[10]) );
  NOR2X1 U112 ( .A(n133), .B(n129), .Y(n132) );
  INVXL U113 ( .A(n85), .Y(n133) );
  XOR2X1 U114 ( .A(n126), .B(n127), .Y(DIFF[11]) );
  AOI21XL U115 ( .A0(n85), .A1(n128), .B0(n129), .Y(n127) );
  NAND2XL U116 ( .A(n86), .B(n67), .Y(n126) );
  XOR2X1 U117 ( .A(n8), .B(n9), .Y(DIFF[9]) );
  XOR2X1 U118 ( .A(n107), .B(n108), .Y(DIFF[14]) );
  NAND2X1 U119 ( .A(n36), .B(n30), .Y(n145) );
  NAND2X1 U120 ( .A(n73), .B(n82), .Y(n81) );
  INVX1 U121 ( .A(n63), .Y(n82) );
  INVXL U122 ( .A(n67), .Y(n66) );
  OAI21XL U123 ( .A0(n28), .A1(n29), .B0(n30), .Y(n21) );
  INVX1 U124 ( .A(n31), .Y(n28) );
  NAND2BX1 U125 ( .AN(n69), .B(n89), .Y(n37) );
  INVX1 U126 ( .A(n152), .Y(n48) );
  INVX1 U127 ( .A(n41), .Y(n46) );
  INVX1 U128 ( .A(n34), .Y(n29) );
  XOR2X1 U129 ( .A(n21), .B(n25), .Y(DIFF[6]) );
  NOR2X1 U130 ( .A(n22), .B(n26), .Y(n25) );
  XOR2X1 U131 ( .A(n18), .B(n19), .Y(DIFF[7]) );
  XOR2X1 U132 ( .A(n13), .B(n14), .Y(DIFF[8]) );
  OAI21XL U133 ( .A0(n47), .A1(n48), .B0(n49), .Y(n42) );
  INVX1 U134 ( .A(n50), .Y(n47) );
  XOR2X1 U135 ( .A(n39), .B(n40), .Y(DIFF[3]) );
  XOR2X1 U136 ( .A(n31), .B(n32), .Y(DIFF[5]) );
  INVX1 U137 ( .A(n89), .Y(n88) );
  XOR2X1 U138 ( .A(n42), .B(n45), .Y(DIFF[2]) );
  XOR2X1 U139 ( .A(n50), .B(n51), .Y(DIFF[1]) );
  INVX1 U140 ( .A(n49), .Y(n52) );
  INVX1 U141 ( .A(A[10]), .Y(n135) );
  INVX1 U142 ( .A(A[11]), .Y(n131) );
  NAND2X1 U143 ( .A(B[6]), .B(n149), .Y(n20) );
  INVX1 U144 ( .A(A[6]), .Y(n149) );
  NAND2X1 U145 ( .A(B[7]), .B(n148), .Y(n23) );
  INVX1 U146 ( .A(A[7]), .Y(n148) );
  NAND2BX2 U147 ( .AN(B[14]), .B(A[14]), .Y(n93) );
  NAND2X1 U148 ( .A(A[9]), .B(n137), .Y(n12) );
  INVX1 U149 ( .A(B[9]), .Y(n137) );
  NAND2X1 U150 ( .A(A[8]), .B(n139), .Y(n17) );
  INVX1 U151 ( .A(B[8]), .Y(n139) );
  NAND2X1 U152 ( .A(A[5]), .B(n146), .Y(n30) );
  INVX1 U153 ( .A(B[5]), .Y(n146) );
  NAND2BXL U154 ( .AN(A[15]), .B(B[15]), .Y(n61) );
  INVXL U155 ( .A(B[10]), .Y(n134) );
  NAND2X1 U156 ( .A(A[7]), .B(n143), .Y(n24) );
  NAND2X1 U157 ( .A(A[6]), .B(n144), .Y(n27) );
  OAI21XL U158 ( .A0(n153), .A1(n154), .B0(n44), .Y(n69) );
  INVX1 U159 ( .A(n43), .Y(n154) );
  AOI21X1 U160 ( .A0(n41), .A1(n157), .B0(n7), .Y(n153) );
  OAI21XL U161 ( .A0(n48), .A1(n53), .B0(n49), .Y(n157) );
  INVX1 U162 ( .A(A[4]), .Y(n151) );
  NAND2X1 U163 ( .A(A[4]), .B(n147), .Y(n36) );
  INVX1 U164 ( .A(B[4]), .Y(n147) );
  INVX1 U165 ( .A(A[2]), .Y(n160) );
  NAND2X1 U166 ( .A(B[3]), .B(n156), .Y(n43) );
  INVX1 U167 ( .A(A[3]), .Y(n156) );
  NAND2X1 U168 ( .A(A[1]), .B(n158), .Y(n49) );
  NOR2BX1 U169 ( .AN(A[2]), .B(B[2]), .Y(n7) );
  NAND2X1 U170 ( .A(B[1]), .B(n159), .Y(n152) );
  INVX1 U171 ( .A(A[1]), .Y(n159) );
  NAND2X1 U172 ( .A(A[3]), .B(n155), .Y(n44) );
  NAND2X1 U173 ( .A(n53), .B(n54), .Y(DIFF[0]) );
  NAND2BX1 U174 ( .AN(n54), .B(n53), .Y(n50) );
  NAND2X1 U175 ( .A(A[0]), .B(n163), .Y(n53) );
  INVX1 U176 ( .A(B[0]), .Y(n163) );
  NAND2X1 U177 ( .A(B[0]), .B(n162), .Y(n54) );
  INVX1 U178 ( .A(A[0]), .Y(n162) );
  NAND3X1 U179 ( .A(n76), .B(n77), .C(n75), .Y(n57) );
  AOI21X1 U180 ( .A0(B[15]), .A1(n78), .B0(n79), .Y(n77) );
  NAND2X4 U181 ( .A(n86), .B(n120), .Y(n68) );
  NAND2X4 U182 ( .A(B[11]), .B(n131), .Y(n86) );
endmodule


module butterfly_DW01_add_36 ( A, B, SUM );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  wire   n1, n2, n4, n5, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123;

  NAND2XL U2 ( .A(B[11]), .B(A[11]), .Y(n65) );
  OR2X2 U3 ( .A(B[11]), .B(A[11]), .Y(n82) );
  NAND3X1 U4 ( .A(n102), .B(n81), .C(n83), .Y(n1) );
  NAND2XL U5 ( .A(n2), .B(n82), .Y(n99) );
  INVX1 U6 ( .A(n1), .Y(n2) );
  NAND3X2 U7 ( .A(n99), .B(n65), .C(n66), .Y(n96) );
  OAI21XL U8 ( .A0(n117), .A1(n71), .B0(n70), .Y(n13) );
  NAND2X1 U9 ( .A(n96), .B(n60), .Y(n95) );
  INVX1 U10 ( .A(n61), .Y(n88) );
  NAND2X1 U11 ( .A(B[14]), .B(A[14]), .Y(n80) );
  XOR2X1 U12 ( .A(B[16]), .B(A[16]), .Y(n8) );
  AND2X2 U13 ( .A(n52), .B(n118), .Y(SUM[0]) );
  OAI21X2 U14 ( .A0(n91), .A1(n5), .B0(n92), .Y(n89) );
  NAND2X2 U15 ( .A(n95), .B(n79), .Y(n93) );
  INVX2 U16 ( .A(n93), .Y(n91) );
  XOR2X4 U17 ( .A(n85), .B(n86), .Y(SUM[15]) );
  NAND2X2 U18 ( .A(n87), .B(n80), .Y(n85) );
  NAND2XL U19 ( .A(B[12]), .B(A[12]), .Y(n79) );
  OR2X2 U20 ( .A(B[12]), .B(A[12]), .Y(n60) );
  NOR2XL U21 ( .A(n19), .B(n20), .Y(n18) );
  INVXL U22 ( .A(n101), .Y(n106) );
  INVXL U23 ( .A(n71), .Y(n67) );
  INVXL U24 ( .A(n70), .Y(n69) );
  NOR2BXL U25 ( .AN(n24), .B(n23), .Y(n26) );
  NOR2BXL U26 ( .AN(n29), .B(n28), .Y(n31) );
  INVXL U27 ( .A(n25), .Y(n22) );
  INVXL U28 ( .A(n68), .Y(n117) );
  NOR2BX2 U29 ( .AN(n54), .B(n56), .Y(n86) );
  NOR2BXL U30 ( .AN(n80), .B(n88), .Y(n90) );
  NOR2BX1 U31 ( .AN(n13), .B(n16), .Y(n102) );
  INVXL U32 ( .A(n60), .Y(n98) );
  NAND2XL U33 ( .A(n60), .B(n61), .Y(n59) );
  NAND2XL U34 ( .A(n82), .B(n65), .Y(n103) );
  NAND2XL U35 ( .A(n110), .B(n15), .Y(n9) );
  NAND2XL U36 ( .A(n13), .B(n84), .Y(n110) );
  NAND4XL U37 ( .A(n81), .B(n82), .C(n83), .D(n84), .Y(n63) );
  INVXL U38 ( .A(n116), .Y(n20) );
  NAND2XL U39 ( .A(B[6]), .B(A[6]), .Y(n24) );
  NAND2XL U40 ( .A(B[5]), .B(A[5]), .Y(n29) );
  INVXL U41 ( .A(n39), .Y(n38) );
  NOR2BXL U42 ( .AN(n47), .B(n51), .Y(n50) );
  NAND2XL U43 ( .A(n48), .B(n49), .Y(n46) );
  INVXL U44 ( .A(n45), .Y(n41) );
  INVXL U45 ( .A(n79), .Y(n78) );
  NOR2X1 U46 ( .A(A[13]), .B(B[13]), .Y(n5) );
  NAND2X1 U47 ( .A(B[10]), .B(A[10]), .Y(n101) );
  OR2X2 U48 ( .A(B[9]), .B(A[9]), .Y(n83) );
  OR2X2 U49 ( .A(A[14]), .B(B[14]), .Y(n61) );
  NAND2XL U50 ( .A(B[7]), .B(A[7]), .Y(n21) );
  OR2X2 U51 ( .A(B[10]), .B(A[10]), .Y(n81) );
  NAND2XL U52 ( .A(B[1]), .B(A[1]), .Y(n47) );
  NOR2X1 U53 ( .A(B[3]), .B(A[3]), .Y(n4) );
  OR2XL U54 ( .A(B[4]), .B(A[4]), .Y(n35) );
  AND3X1 U55 ( .A(n54), .B(n55), .C(n53), .Y(n7) );
  INVX1 U56 ( .A(B[0]), .Y(n122) );
  INVX1 U57 ( .A(n114), .Y(n28) );
  NAND2BX1 U58 ( .AN(n88), .B(n89), .Y(n87) );
  INVX1 U59 ( .A(n115), .Y(n23) );
  OAI21XL U60 ( .A0(n27), .A1(n28), .B0(n29), .Y(n25) );
  INVX1 U61 ( .A(n30), .Y(n27) );
  AOI21X1 U62 ( .A0(n67), .A1(n68), .B0(n69), .Y(n62) );
  XOR2X1 U63 ( .A(n25), .B(n26), .Y(SUM[6]) );
  XOR2X1 U64 ( .A(n17), .B(n18), .Y(SUM[7]) );
  OAI21XL U65 ( .A0(n22), .A1(n23), .B0(n24), .Y(n17) );
  XOR2X1 U66 ( .A(n30), .B(n31), .Y(SUM[5]) );
  INVX1 U67 ( .A(n43), .Y(n40) );
  OAI21XL U68 ( .A0(n109), .A1(n12), .B0(n11), .Y(n105) );
  INVX1 U69 ( .A(n9), .Y(n109) );
  NAND4X1 U70 ( .A(n35), .B(n114), .C(n115), .D(n116), .Y(n71) );
  NAND3X1 U71 ( .A(n100), .B(n81), .C(n82), .Y(n66) );
  OAI211X1 U72 ( .A0(n12), .A1(n15), .B0(n11), .C0(n101), .Y(n100) );
  XOR2X1 U73 ( .A(n96), .B(n97), .Y(SUM[12]) );
  NOR2BX1 U74 ( .AN(n79), .B(n98), .Y(n97) );
  NAND2BX1 U75 ( .AN(n20), .B(n111), .Y(n70) );
  NAND3X1 U76 ( .A(n112), .B(n24), .C(n21), .Y(n111) );
  NAND2BX1 U77 ( .AN(n23), .B(n113), .Y(n112) );
  OAI21XL U78 ( .A0(n28), .A1(n33), .B0(n29), .Y(n113) );
  INVX1 U79 ( .A(n83), .Y(n12) );
  OR2X2 U80 ( .A(B[6]), .B(A[6]), .Y(n115) );
  OR2X2 U81 ( .A(B[5]), .B(A[5]), .Y(n114) );
  INVX1 U82 ( .A(n84), .Y(n16) );
  AND2X1 U83 ( .A(n66), .B(n65), .Y(n64) );
  XOR2X1 U84 ( .A(n105), .B(n107), .Y(SUM[10]) );
  NOR2BX1 U85 ( .AN(n101), .B(n108), .Y(n107) );
  INVX1 U86 ( .A(n81), .Y(n108) );
  XOR2X1 U87 ( .A(n103), .B(n104), .Y(SUM[11]) );
  AOI21X1 U88 ( .A0(n81), .A1(n105), .B0(n106), .Y(n104) );
  XOR2X1 U89 ( .A(n9), .B(n10), .Y(SUM[9]) );
  NOR2BXL U90 ( .AN(n11), .B(n12), .Y(n10) );
  OAI21XL U91 ( .A0(n119), .A1(n4), .B0(n39), .Y(n68) );
  AOI21X1 U92 ( .A0(n45), .A1(n120), .B0(n121), .Y(n119) );
  INVX1 U93 ( .A(n42), .Y(n121) );
  OAI21XL U94 ( .A0(n51), .A1(n52), .B0(n47), .Y(n120) );
  OAI21XL U95 ( .A0(n32), .A1(n117), .B0(n33), .Y(n30) );
  INVX1 U96 ( .A(n35), .Y(n32) );
  INVX1 U97 ( .A(n48), .Y(n51) );
  XOR2X1 U98 ( .A(n13), .B(n14), .Y(SUM[8]) );
  NOR2BX1 U99 ( .AN(n15), .B(n16), .Y(n14) );
  INVX1 U100 ( .A(n21), .Y(n19) );
  XOR2X1 U101 ( .A(n68), .B(n34), .Y(SUM[4]) );
  NOR2BX1 U102 ( .AN(n33), .B(n32), .Y(n34) );
  XOR2X1 U103 ( .A(n49), .B(n50), .Y(SUM[1]) );
  XOR2X1 U104 ( .A(n43), .B(n44), .Y(SUM[2]) );
  NOR2BX1 U105 ( .AN(n42), .B(n41), .Y(n44) );
  XOR2X1 U106 ( .A(n36), .B(n37), .Y(SUM[3]) );
  NOR2X1 U107 ( .A(n38), .B(n4), .Y(n37) );
  OAI21XL U108 ( .A0(n40), .A1(n41), .B0(n42), .Y(n36) );
  NAND2X1 U109 ( .A(n46), .B(n47), .Y(n43) );
  INVX1 U110 ( .A(n52), .Y(n49) );
  OAI21XL U111 ( .A0(n72), .A1(n73), .B0(n74), .Y(n53) );
  INVXL U112 ( .A(n80), .Y(n72) );
  OR2X2 U113 ( .A(B[8]), .B(A[8]), .Y(n84) );
  NAND2X1 U114 ( .A(B[8]), .B(A[8]), .Y(n15) );
  OR2X2 U115 ( .A(B[7]), .B(A[7]), .Y(n116) );
  NAND2XL U116 ( .A(B[9]), .B(A[9]), .Y(n11) );
  NAND3BX1 U117 ( .AN(n56), .B(n57), .C(n58), .Y(n55) );
  OAI21XL U118 ( .A0(n62), .A1(n63), .B0(n64), .Y(n57) );
  NOR2X1 U119 ( .A(n59), .B(n5), .Y(n58) );
  OR2X2 U120 ( .A(A[15]), .B(B[15]), .Y(n74) );
  NAND2X1 U121 ( .A(B[4]), .B(A[4]), .Y(n33) );
  NAND2X1 U122 ( .A(B[2]), .B(A[2]), .Y(n42) );
  OR2X2 U123 ( .A(B[2]), .B(A[2]), .Y(n45) );
  NAND2X1 U124 ( .A(B[3]), .B(A[3]), .Y(n39) );
  OR2X2 U125 ( .A(B[1]), .B(A[1]), .Y(n48) );
  NAND2X1 U126 ( .A(B[0]), .B(A[0]), .Y(n52) );
  NAND2X1 U127 ( .A(n122), .B(n123), .Y(n118) );
  INVX1 U128 ( .A(A[0]), .Y(n123) );
  XNOR2X2 U129 ( .A(n7), .B(n8), .Y(SUM[16]) );
  NAND2X1 U130 ( .A(B[15]), .B(A[15]), .Y(n54) );
  NOR2X1 U131 ( .A(A[15]), .B(B[15]), .Y(n56) );
  XOR2X1 U132 ( .A(n93), .B(n94), .Y(SUM[13]) );
  XOR2X1 U133 ( .A(n89), .B(n90), .Y(SUM[14]) );
  NAND2XL U134 ( .A(B[13]), .B(A[13]), .Y(n92) );
  NAND2XL U135 ( .A(B[13]), .B(A[13]), .Y(n75) );
  OAI21XL U136 ( .A0(A[13]), .A1(B[13]), .B0(n78), .Y(n76) );
  NOR2BX1 U137 ( .AN(n92), .B(n5), .Y(n94) );
  AOI21X1 U138 ( .A0(n75), .A1(n76), .B0(n77), .Y(n73) );
  NOR2XL U139 ( .A(B[14]), .B(A[14]), .Y(n77) );
endmodule


module butterfly_DW01_add_35 ( A, B, SUM );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  wire   n2, n3, n4, n5, n6, n7, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126;

  NAND2X2 U2 ( .A(n98), .B(n81), .Y(n96) );
  NAND2X2 U3 ( .A(n62), .B(n63), .Y(n61) );
  OR2X4 U4 ( .A(A[15]), .B(B[15]), .Y(n6) );
  OAI21X2 U5 ( .A0(n74), .A1(n75), .B0(n76), .Y(n56) );
  OR2X4 U6 ( .A(A[15]), .B(B[15]), .Y(n76) );
  OR2X2 U7 ( .A(A[14]), .B(B[14]), .Y(n63) );
  OAI21XL U8 ( .A0(n120), .A1(n73), .B0(n72), .Y(n16) );
  NOR2X1 U9 ( .A(n11), .B(n61), .Y(n60) );
  AND2X2 U10 ( .A(n55), .B(n121), .Y(SUM[0]) );
  OAI21X2 U11 ( .A0(n94), .A1(n11), .B0(n95), .Y(n92) );
  INVX2 U12 ( .A(n96), .Y(n94) );
  INVX1 U13 ( .A(A[16]), .Y(n3) );
  NOR2X1 U14 ( .A(A[13]), .B(B[13]), .Y(n11) );
  NAND2XL U15 ( .A(B[14]), .B(A[14]), .Y(n82) );
  NOR2XL U16 ( .A(B[14]), .B(A[14]), .Y(n79) );
  NAND2X1 U17 ( .A(B[16]), .B(n3), .Y(n4) );
  NAND2X1 U18 ( .A(n2), .B(A[16]), .Y(n5) );
  NAND2X2 U19 ( .A(n4), .B(n5), .Y(n10) );
  INVX1 U20 ( .A(B[16]), .Y(n2) );
  NOR2XL U21 ( .A(n22), .B(n23), .Y(n21) );
  NAND2XL U22 ( .A(B[12]), .B(A[12]), .Y(n81) );
  NAND2XL U23 ( .A(B[11]), .B(A[11]), .Y(n67) );
  XNOR2X4 U24 ( .A(n9), .B(n10), .Y(SUM[16]) );
  AOI21XL U25 ( .A0(n69), .A1(n70), .B0(n71), .Y(n64) );
  INVXL U26 ( .A(n73), .Y(n69) );
  INVXL U27 ( .A(n72), .Y(n71) );
  NOR2BXL U28 ( .AN(n27), .B(n26), .Y(n29) );
  NOR2BXL U29 ( .AN(n32), .B(n31), .Y(n34) );
  INVXL U30 ( .A(n28), .Y(n25) );
  INVXL U31 ( .A(n70), .Y(n120) );
  XOR2X2 U32 ( .A(n87), .B(n88), .Y(SUM[15]) );
  NOR2BX2 U33 ( .AN(n57), .B(n89), .Y(n88) );
  NOR2BX1 U34 ( .AN(n16), .B(n19), .Y(n105) );
  NAND4XL U35 ( .A(n83), .B(n84), .C(n85), .D(n86), .Y(n65) );
  INVXL U36 ( .A(n63), .Y(n91) );
  NOR2BXL U37 ( .AN(n14), .B(n15), .Y(n13) );
  NAND2XL U38 ( .A(n113), .B(n18), .Y(n12) );
  NAND2XL U39 ( .A(n16), .B(n86), .Y(n113) );
  INVXL U40 ( .A(n119), .Y(n23) );
  NAND2XL U41 ( .A(B[6]), .B(A[6]), .Y(n27) );
  NAND2XL U42 ( .A(B[5]), .B(A[5]), .Y(n32) );
  NOR2BXL U43 ( .AN(n50), .B(n54), .Y(n53) );
  NAND2XL U44 ( .A(n51), .B(n52), .Y(n49) );
  INVXL U45 ( .A(n48), .Y(n44) );
  INVXL U46 ( .A(n42), .Y(n41) );
  NAND3X1 U47 ( .A(n6), .B(n59), .C(n60), .Y(n58) );
  OR2X2 U48 ( .A(B[12]), .B(A[12]), .Y(n62) );
  NAND2X1 U49 ( .A(B[10]), .B(A[10]), .Y(n104) );
  OR2X2 U50 ( .A(B[11]), .B(A[11]), .Y(n84) );
  OR2X2 U51 ( .A(B[9]), .B(A[9]), .Y(n85) );
  NAND2XL U52 ( .A(B[9]), .B(A[9]), .Y(n14) );
  NAND2XL U53 ( .A(B[7]), .B(A[7]), .Y(n24) );
  OR2X2 U54 ( .A(B[10]), .B(A[10]), .Y(n83) );
  NAND2XL U55 ( .A(B[1]), .B(A[1]), .Y(n50) );
  NOR2X1 U56 ( .A(B[3]), .B(A[3]), .Y(n7) );
  OR2XL U57 ( .A(B[4]), .B(A[4]), .Y(n38) );
  AND3X4 U58 ( .A(n57), .B(n58), .C(n56), .Y(n9) );
  INVX1 U59 ( .A(n117), .Y(n31) );
  NAND2BX1 U60 ( .AN(n91), .B(n92), .Y(n90) );
  INVX1 U61 ( .A(n118), .Y(n26) );
  OAI21XL U62 ( .A0(n30), .A1(n31), .B0(n32), .Y(n28) );
  INVX1 U63 ( .A(n33), .Y(n30) );
  XOR2X1 U64 ( .A(n28), .B(n29), .Y(SUM[6]) );
  XOR2X1 U65 ( .A(n20), .B(n21), .Y(SUM[7]) );
  OAI21XL U66 ( .A0(n25), .A1(n26), .B0(n27), .Y(n20) );
  XOR2X1 U67 ( .A(n33), .B(n34), .Y(SUM[5]) );
  NOR2BX1 U68 ( .AN(n82), .B(n91), .Y(n93) );
  OAI21XL U69 ( .A0(n112), .A1(n15), .B0(n14), .Y(n108) );
  INVX1 U70 ( .A(n12), .Y(n112) );
  NAND4X1 U71 ( .A(n38), .B(n117), .C(n118), .D(n119), .Y(n73) );
  NAND3X1 U72 ( .A(n102), .B(n67), .C(n68), .Y(n99) );
  NAND4X1 U73 ( .A(n105), .B(n85), .C(n83), .D(n84), .Y(n102) );
  XOR2X1 U74 ( .A(n12), .B(n13), .Y(SUM[9]) );
  XOR2X1 U75 ( .A(n108), .B(n110), .Y(SUM[10]) );
  NOR2BX1 U76 ( .AN(n104), .B(n111), .Y(n110) );
  INVX1 U77 ( .A(n83), .Y(n111) );
  XOR2X1 U78 ( .A(n99), .B(n100), .Y(SUM[12]) );
  NOR2BX1 U79 ( .AN(n81), .B(n101), .Y(n100) );
  INVX1 U80 ( .A(n62), .Y(n101) );
  NAND2BX1 U81 ( .AN(n23), .B(n114), .Y(n72) );
  NAND3X1 U82 ( .A(n115), .B(n27), .C(n24), .Y(n114) );
  NAND2BX1 U83 ( .AN(n26), .B(n116), .Y(n115) );
  OAI21XL U84 ( .A0(n31), .A1(n36), .B0(n32), .Y(n116) );
  NAND3X1 U85 ( .A(n103), .B(n83), .C(n84), .Y(n68) );
  OAI211X1 U86 ( .A0(n15), .A1(n18), .B0(n14), .C0(n104), .Y(n103) );
  INVX1 U87 ( .A(n85), .Y(n15) );
  OR2X2 U88 ( .A(B[6]), .B(A[6]), .Y(n118) );
  OR2X2 U89 ( .A(B[5]), .B(A[5]), .Y(n117) );
  INVX1 U90 ( .A(n86), .Y(n19) );
  XOR2X1 U91 ( .A(n106), .B(n107), .Y(SUM[11]) );
  AOI21X1 U92 ( .A0(n83), .A1(n108), .B0(n109), .Y(n107) );
  INVX1 U93 ( .A(n104), .Y(n109) );
  AND2X1 U94 ( .A(n68), .B(n67), .Y(n66) );
  NAND2X1 U95 ( .A(n90), .B(n82), .Y(n87) );
  INVX1 U96 ( .A(n76), .Y(n89) );
  NAND2X1 U97 ( .A(n99), .B(n62), .Y(n98) );
  OAI21XL U98 ( .A0(n122), .A1(n7), .B0(n42), .Y(n70) );
  AOI21X1 U99 ( .A0(n48), .A1(n123), .B0(n124), .Y(n122) );
  INVX1 U100 ( .A(n45), .Y(n124) );
  OAI21XL U101 ( .A0(n54), .A1(n55), .B0(n50), .Y(n123) );
  XOR2X1 U102 ( .A(n16), .B(n17), .Y(SUM[8]) );
  NOR2BX1 U103 ( .AN(n18), .B(n19), .Y(n17) );
  INVX1 U104 ( .A(n51), .Y(n54) );
  INVX1 U105 ( .A(n24), .Y(n22) );
  OAI21XL U106 ( .A0(n35), .A1(n120), .B0(n36), .Y(n33) );
  INVX1 U107 ( .A(n38), .Y(n35) );
  XOR2X1 U108 ( .A(n70), .B(n37), .Y(SUM[4]) );
  NOR2BX1 U109 ( .AN(n36), .B(n35), .Y(n37) );
  XOR2X1 U110 ( .A(n52), .B(n53), .Y(SUM[1]) );
  XOR2X1 U111 ( .A(n46), .B(n47), .Y(SUM[2]) );
  NOR2BX1 U112 ( .AN(n45), .B(n44), .Y(n47) );
  XOR2X1 U113 ( .A(n39), .B(n40), .Y(SUM[3]) );
  OAI21XL U114 ( .A0(n43), .A1(n44), .B0(n45), .Y(n39) );
  NOR2X1 U115 ( .A(n41), .B(n7), .Y(n40) );
  INVX1 U116 ( .A(n46), .Y(n43) );
  NAND2X1 U117 ( .A(n49), .B(n50), .Y(n46) );
  INVX1 U118 ( .A(n55), .Y(n52) );
  NAND2X1 U119 ( .A(n125), .B(n126), .Y(n121) );
  INVX1 U120 ( .A(B[0]), .Y(n125) );
  INVXL U121 ( .A(n82), .Y(n74) );
  AOI21X1 U122 ( .A0(n77), .A1(n78), .B0(n79), .Y(n75) );
  OR2X2 U123 ( .A(B[8]), .B(A[8]), .Y(n86) );
  NAND2X1 U124 ( .A(B[8]), .B(A[8]), .Y(n18) );
  OR2X2 U125 ( .A(B[7]), .B(A[7]), .Y(n119) );
  OAI21XL U126 ( .A0(n64), .A1(n65), .B0(n66), .Y(n59) );
  OAI21X1 U127 ( .A0(A[13]), .A1(B[13]), .B0(n80), .Y(n78) );
  INVX1 U128 ( .A(n81), .Y(n80) );
  NAND2XL U129 ( .A(B[15]), .B(A[15]), .Y(n57) );
  NAND2X1 U130 ( .A(B[4]), .B(A[4]), .Y(n36) );
  NAND2X1 U131 ( .A(B[2]), .B(A[2]), .Y(n45) );
  OR2X2 U132 ( .A(B[2]), .B(A[2]), .Y(n48) );
  NAND2X1 U133 ( .A(B[3]), .B(A[3]), .Y(n42) );
  OR2X2 U134 ( .A(B[1]), .B(A[1]), .Y(n51) );
  NAND2X1 U135 ( .A(B[0]), .B(A[0]), .Y(n55) );
  INVX1 U136 ( .A(A[0]), .Y(n126) );
  XOR2X1 U137 ( .A(n96), .B(n97), .Y(SUM[13]) );
  XOR2X1 U138 ( .A(n92), .B(n93), .Y(SUM[14]) );
  NAND2XL U139 ( .A(n84), .B(n67), .Y(n106) );
  NAND2XL U140 ( .A(B[13]), .B(A[13]), .Y(n95) );
  NAND2X1 U141 ( .A(B[13]), .B(A[13]), .Y(n77) );
  NOR2BX1 U142 ( .AN(n95), .B(n11), .Y(n97) );
endmodule


module butterfly_DW01_add_37 ( A, B, SUM );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n14, n15, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145;

  NAND2X2 U2 ( .A(n17), .B(n18), .Y(n3) );
  NAND2X4 U3 ( .A(n1), .B(n2), .Y(n4) );
  NAND2X4 U4 ( .A(n3), .B(n4), .Y(SUM[16]) );
  INVX4 U5 ( .A(n17), .Y(n1) );
  INVX8 U6 ( .A(n18), .Y(n2) );
  NAND2X2 U7 ( .A(n101), .B(n6), .Y(n7) );
  NAND2X4 U8 ( .A(n5), .B(n102), .Y(n8) );
  NAND2X4 U9 ( .A(n7), .B(n8), .Y(SUM[15]) );
  INVX4 U10 ( .A(n101), .Y(n5) );
  INVX1 U11 ( .A(n102), .Y(n6) );
  NAND2X4 U12 ( .A(n105), .B(n95), .Y(n101) );
  NAND2X1 U13 ( .A(n112), .B(n10), .Y(n11) );
  NAND2XL U14 ( .A(n9), .B(n113), .Y(n12) );
  NAND2X2 U15 ( .A(n11), .B(n12), .Y(SUM[13]) );
  INVXL U16 ( .A(n112), .Y(n9) );
  INVXL U17 ( .A(n113), .Y(n10) );
  NOR2BXL U18 ( .AN(n111), .B(n73), .Y(n113) );
  NAND2BX2 U19 ( .AN(n106), .B(n107), .Y(n105) );
  NAND2X2 U20 ( .A(n119), .B(n120), .Y(n75) );
  INVX2 U21 ( .A(A[12]), .Y(n120) );
  AOI21X1 U22 ( .A0(n90), .A1(n91), .B0(n92), .Y(n88) );
  OAI21X2 U23 ( .A0(n87), .A1(n88), .B0(n89), .Y(n68) );
  NAND3X1 U24 ( .A(n122), .B(n97), .C(n98), .Y(n81) );
  OAI211X1 U25 ( .A0(n26), .A1(n29), .B0(n25), .C0(n123), .Y(n122) );
  NAND2XL U26 ( .A(B[11]), .B(A[11]), .Y(n80) );
  NAND2X2 U27 ( .A(n115), .B(n94), .Y(n112) );
  NAND2X1 U28 ( .A(n116), .B(n75), .Y(n115) );
  INVXL U29 ( .A(B[13]), .Y(n114) );
  INVX2 U30 ( .A(B[15]), .Y(n104) );
  OAI21X2 U31 ( .A0(n110), .A1(n73), .B0(n111), .Y(n107) );
  CLKINVX3 U32 ( .A(n112), .Y(n110) );
  OAI21XL U33 ( .A0(n139), .A1(n86), .B0(n85), .Y(n27) );
  NAND2X1 U34 ( .A(B[10]), .B(A[10]), .Y(n123) );
  NAND3X1 U35 ( .A(n14), .B(n71), .C(n72), .Y(n70) );
  OR2X2 U36 ( .A(A[15]), .B(B[15]), .Y(n14) );
  AND2X2 U37 ( .A(n67), .B(n140), .Y(SUM[0]) );
  NAND2BX1 U38 ( .AN(A[13]), .B(n114), .Y(n96) );
  CLKINVX2 U39 ( .A(B[16]), .Y(n19) );
  NAND2X2 U40 ( .A(n19), .B(n20), .Y(n22) );
  NAND2X1 U41 ( .A(B[16]), .B(A[16]), .Y(n21) );
  NAND3X2 U42 ( .A(n121), .B(n80), .C(n81), .Y(n116) );
  NOR2X2 U43 ( .A(n74), .B(n73), .Y(n72) );
  NAND2X2 U44 ( .A(n75), .B(n76), .Y(n74) );
  INVX2 U45 ( .A(n89), .Y(n103) );
  NAND2X2 U46 ( .A(B[13]), .B(A[13]), .Y(n111) );
  NAND2X4 U47 ( .A(n21), .B(n22), .Y(n18) );
  NAND2X1 U48 ( .A(B[15]), .B(A[15]), .Y(n69) );
  NAND4X1 U49 ( .A(n124), .B(n99), .C(n97), .D(n98), .Y(n121) );
  NAND2XL U50 ( .A(n136), .B(n41), .Y(n135) );
  INVX2 U51 ( .A(A[16]), .Y(n20) );
  AND2X1 U52 ( .A(n81), .B(n80), .Y(n79) );
  NAND3X2 U53 ( .A(n69), .B(n70), .C(n68), .Y(n17) );
  OR2X2 U54 ( .A(B[8]), .B(A[8]), .Y(n100) );
  NAND4XL U55 ( .A(n97), .B(n98), .C(n99), .D(n100), .Y(n78) );
  INVXL U56 ( .A(n76), .Y(n106) );
  INVXL U57 ( .A(n97), .Y(n131) );
  NAND2XL U58 ( .A(n133), .B(n29), .Y(n23) );
  NAND2XL U59 ( .A(n27), .B(n100), .Y(n133) );
  INVXL U60 ( .A(n138), .Y(n34) );
  NOR2XL U61 ( .A(n33), .B(n34), .Y(n32) );
  INVXL U62 ( .A(n39), .Y(n36) );
  INVXL U63 ( .A(n86), .Y(n82) );
  INVXL U64 ( .A(n85), .Y(n84) );
  NOR2BXL U65 ( .AN(n44), .B(n43), .Y(n46) );
  INVXL U66 ( .A(n83), .Y(n139) );
  INVXL U67 ( .A(n41), .Y(n37) );
  INVXL U68 ( .A(n60), .Y(n56) );
  INVXL U69 ( .A(n54), .Y(n53) );
  NAND2X2 U70 ( .A(B[14]), .B(A[14]), .Y(n95) );
  NAND2X2 U71 ( .A(B[12]), .B(A[12]), .Y(n94) );
  INVX1 U72 ( .A(n94), .Y(n93) );
  INVXL U73 ( .A(B[12]), .Y(n119) );
  NOR2XL U74 ( .A(B[14]), .B(A[14]), .Y(n92) );
  OR2X2 U75 ( .A(B[9]), .B(A[9]), .Y(n99) );
  NAND2XL U76 ( .A(B[9]), .B(A[9]), .Y(n25) );
  NAND2XL U77 ( .A(B[6]), .B(A[6]), .Y(n38) );
  NAND2XL U78 ( .A(B[5]), .B(A[5]), .Y(n44) );
  NAND2XL U79 ( .A(B[7]), .B(A[7]), .Y(n35) );
  NOR2X1 U80 ( .A(B[3]), .B(A[3]), .Y(n15) );
  OR2XL U81 ( .A(B[4]), .B(A[4]), .Y(n50) );
  INVX1 U82 ( .A(B[0]), .Y(n144) );
  XOR2X1 U83 ( .A(n126), .B(n127), .Y(SUM[11]) );
  AOI21X1 U84 ( .A0(n97), .A1(n128), .B0(n129), .Y(n127) );
  INVXL U85 ( .A(n123), .Y(n129) );
  XOR2X1 U86 ( .A(n116), .B(n117), .Y(SUM[12]) );
  NOR2BX1 U87 ( .AN(n94), .B(n118), .Y(n117) );
  INVXL U88 ( .A(n75), .Y(n118) );
  OAI21XL U89 ( .A0(n132), .A1(n26), .B0(n25), .Y(n128) );
  INVX1 U90 ( .A(n23), .Y(n132) );
  XOR2X1 U91 ( .A(n107), .B(n108), .Y(SUM[14]) );
  NOR2BX1 U92 ( .AN(n95), .B(n106), .Y(n108) );
  NAND4X1 U93 ( .A(n50), .B(n137), .C(n41), .D(n138), .Y(n86) );
  NOR2X1 U94 ( .A(n125), .B(n30), .Y(n124) );
  INVX1 U95 ( .A(n27), .Y(n125) );
  INVX1 U96 ( .A(n137), .Y(n43) );
  XOR2X1 U97 ( .A(n23), .B(n24), .Y(SUM[9]) );
  NOR2BX1 U98 ( .AN(n25), .B(n26), .Y(n24) );
  XOR2X1 U99 ( .A(n27), .B(n28), .Y(SUM[8]) );
  NOR2BX1 U100 ( .AN(n29), .B(n30), .Y(n28) );
  XOR2X1 U101 ( .A(n128), .B(n130), .Y(SUM[10]) );
  NOR2BX1 U102 ( .AN(n123), .B(n131), .Y(n130) );
  NAND2BX1 U103 ( .AN(n34), .B(n134), .Y(n85) );
  NAND3X1 U104 ( .A(n135), .B(n38), .C(n35), .Y(n134) );
  OAI21XL U105 ( .A0(n43), .A1(n48), .B0(n44), .Y(n136) );
  AOI21X1 U106 ( .A0(n82), .A1(n83), .B0(n84), .Y(n77) );
  INVX1 U107 ( .A(n99), .Y(n26) );
  INVX1 U108 ( .A(n100), .Y(n30) );
  XOR2X1 U109 ( .A(n39), .B(n40), .Y(SUM[6]) );
  NOR2BX1 U110 ( .AN(n38), .B(n37), .Y(n40) );
  XOR2X1 U111 ( .A(n45), .B(n46), .Y(SUM[5]) );
  XOR2X1 U112 ( .A(n31), .B(n32), .Y(SUM[7]) );
  OAI21XL U113 ( .A0(n36), .A1(n37), .B0(n38), .Y(n31) );
  OAI21XL U114 ( .A0(n42), .A1(n43), .B0(n44), .Y(n39) );
  INVX1 U115 ( .A(n45), .Y(n42) );
  OAI21XL U116 ( .A0(n47), .A1(n139), .B0(n48), .Y(n45) );
  INVX1 U117 ( .A(n50), .Y(n47) );
  INVX1 U118 ( .A(n63), .Y(n66) );
  INVX1 U119 ( .A(n35), .Y(n33) );
  XOR2X1 U120 ( .A(n83), .B(n49), .Y(SUM[4]) );
  NOR2BX1 U121 ( .AN(n48), .B(n47), .Y(n49) );
  XOR2X1 U122 ( .A(n51), .B(n52), .Y(SUM[3]) );
  OAI21XL U123 ( .A0(n55), .A1(n56), .B0(n57), .Y(n51) );
  NOR2X1 U124 ( .A(n53), .B(n15), .Y(n52) );
  INVX1 U125 ( .A(n58), .Y(n55) );
  XOR2X1 U126 ( .A(n64), .B(n65), .Y(SUM[1]) );
  NOR2BX1 U127 ( .AN(n62), .B(n66), .Y(n65) );
  XOR2X1 U128 ( .A(n58), .B(n59), .Y(SUM[2]) );
  NOR2BX1 U129 ( .AN(n57), .B(n56), .Y(n59) );
  NAND2X1 U130 ( .A(n61), .B(n62), .Y(n58) );
  NAND2X1 U131 ( .A(n63), .B(n64), .Y(n61) );
  OR2X4 U132 ( .A(B[10]), .B(A[10]), .Y(n97) );
  OR2X2 U133 ( .A(B[6]), .B(A[6]), .Y(n41) );
  OAI21XL U134 ( .A0(A[13]), .A1(B[13]), .B0(n93), .Y(n91) );
  INVXL U135 ( .A(n95), .Y(n87) );
  NAND2XL U136 ( .A(B[13]), .B(A[13]), .Y(n90) );
  OR2X4 U137 ( .A(B[11]), .B(A[11]), .Y(n98) );
  NAND2X1 U138 ( .A(B[8]), .B(A[8]), .Y(n29) );
  OR2X2 U139 ( .A(B[7]), .B(A[7]), .Y(n138) );
  OAI21XL U140 ( .A0(n77), .A1(n78), .B0(n79), .Y(n71) );
  OR2X2 U141 ( .A(B[5]), .B(A[5]), .Y(n137) );
  OAI21XL U142 ( .A0(n141), .A1(n15), .B0(n54), .Y(n83) );
  AOI21X1 U143 ( .A0(n60), .A1(n142), .B0(n143), .Y(n141) );
  INVX1 U144 ( .A(n57), .Y(n143) );
  OAI21XL U145 ( .A0(n66), .A1(n67), .B0(n62), .Y(n142) );
  NAND2X1 U146 ( .A(B[4]), .B(A[4]), .Y(n48) );
  NAND2X1 U147 ( .A(B[1]), .B(A[1]), .Y(n62) );
  NAND2X1 U148 ( .A(B[2]), .B(A[2]), .Y(n57) );
  OR2X2 U149 ( .A(B[2]), .B(A[2]), .Y(n60) );
  NAND2X1 U150 ( .A(B[3]), .B(A[3]), .Y(n54) );
  OR2X2 U151 ( .A(B[1]), .B(A[1]), .Y(n63) );
  INVX1 U152 ( .A(n67), .Y(n64) );
  NAND2X1 U153 ( .A(B[0]), .B(A[0]), .Y(n67) );
  NAND2X1 U154 ( .A(n144), .B(n145), .Y(n140) );
  INVX1 U155 ( .A(A[0]), .Y(n145) );
  INVX4 U156 ( .A(B[14]), .Y(n109) );
  INVX2 U157 ( .A(n96), .Y(n73) );
  NAND2XL U158 ( .A(n98), .B(n80), .Y(n126) );
  NOR2BX4 U159 ( .AN(n69), .B(n103), .Y(n102) );
  NAND2BX4 U160 ( .AN(A[15]), .B(n104), .Y(n89) );
  NAND2BX4 U161 ( .AN(A[14]), .B(n109), .Y(n76) );
endmodule


module butterfly_DW01_add_34 ( A, B, SUM );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  wire   n2, n3, n4, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124;

  NAND2X2 U2 ( .A(n95), .B(n79), .Y(n93) );
  NAND3X2 U3 ( .A(n54), .B(n55), .C(n53), .Y(n52) );
  NAND2X2 U4 ( .A(n96), .B(n60), .Y(n95) );
  NAND3X2 U5 ( .A(n99), .B(n65), .C(n66), .Y(n96) );
  OAI21X1 U6 ( .A0(A[13]), .A1(B[13]), .B0(n78), .Y(n76) );
  NOR2BX2 U7 ( .AN(n54), .B(n87), .Y(n86) );
  OR2X2 U8 ( .A(B[11]), .B(A[11]), .Y(n82) );
  NAND2X1 U9 ( .A(n3), .B(n92), .Y(n90) );
  NAND2X1 U10 ( .A(n93), .B(n2), .Y(n3) );
  INVX1 U11 ( .A(n7), .Y(n2) );
  NAND2X1 U12 ( .A(n60), .B(n61), .Y(n59) );
  XOR2X2 U13 ( .A(n85), .B(n86), .Y(SUM[15]) );
  NAND2X1 U14 ( .A(n88), .B(n80), .Y(n85) );
  NAND2BX1 U15 ( .AN(n89), .B(n90), .Y(n88) );
  AND2X2 U16 ( .A(n51), .B(n119), .Y(SUM[0]) );
  AOI21XL U17 ( .A0(n75), .A1(n76), .B0(n77), .Y(n73) );
  NAND2XL U18 ( .A(B[14]), .B(A[14]), .Y(n80) );
  OR2X4 U19 ( .A(A[14]), .B(B[14]), .Y(n61) );
  NAND2X1 U20 ( .A(B[12]), .B(A[12]), .Y(n79) );
  NOR2X1 U21 ( .A(n59), .B(n7), .Y(n58) );
  NOR2X2 U22 ( .A(A[13]), .B(B[13]), .Y(n7) );
  NAND4X1 U23 ( .A(n102), .B(n83), .C(n81), .D(n82), .Y(n99) );
  NOR2X1 U24 ( .A(n103), .B(n15), .Y(n102) );
  INVX1 U25 ( .A(n12), .Y(n103) );
  XOR2X1 U26 ( .A(n96), .B(n97), .Y(SUM[12]) );
  INVXL U27 ( .A(n60), .Y(n98) );
  INVXL U28 ( .A(n101), .Y(n107) );
  INVXL U29 ( .A(n61), .Y(n89) );
  NAND2XL U30 ( .A(n111), .B(n14), .Y(n8) );
  NAND2XL U31 ( .A(n12), .B(n84), .Y(n111) );
  INVXL U32 ( .A(n71), .Y(n67) );
  INVXL U33 ( .A(n70), .Y(n69) );
  INVXL U34 ( .A(n68), .Y(n118) );
  INVXL U35 ( .A(n24), .Y(n21) );
  NAND2XL U36 ( .A(n82), .B(n65), .Y(n104) );
  NAND4XL U37 ( .A(n81), .B(n82), .C(n83), .D(n84), .Y(n63) );
  INVXL U38 ( .A(n117), .Y(n19) );
  NOR2BXL U39 ( .AN(n23), .B(n22), .Y(n25) );
  NOR2BXL U40 ( .AN(n28), .B(n27), .Y(n30) );
  NOR2BXL U41 ( .AN(n46), .B(n50), .Y(n49) );
  NAND2XL U42 ( .A(n47), .B(n48), .Y(n45) );
  INVXL U43 ( .A(n44), .Y(n40) );
  INVXL U44 ( .A(n38), .Y(n37) );
  NAND2XL U45 ( .A(B[13]), .B(A[13]), .Y(n75) );
  OAI21X1 U46 ( .A0(n72), .A1(n73), .B0(n74), .Y(n53) );
  NAND2XL U47 ( .A(B[11]), .B(A[11]), .Y(n65) );
  OR2X2 U48 ( .A(B[12]), .B(A[12]), .Y(n60) );
  OR2X2 U49 ( .A(B[9]), .B(A[9]), .Y(n83) );
  NAND2X1 U50 ( .A(B[10]), .B(A[10]), .Y(n101) );
  OR2X2 U51 ( .A(B[10]), .B(A[10]), .Y(n81) );
  NAND2XL U52 ( .A(B[6]), .B(A[6]), .Y(n23) );
  NAND2XL U53 ( .A(B[5]), .B(A[5]), .Y(n28) );
  NAND2XL U54 ( .A(B[7]), .B(A[7]), .Y(n20) );
  NAND2XL U55 ( .A(B[1]), .B(A[1]), .Y(n46) );
  NOR2X1 U56 ( .A(B[3]), .B(A[3]), .Y(n4) );
  OR2XL U57 ( .A(B[4]), .B(A[4]), .Y(n34) );
  XOR2X2 U58 ( .A(n52), .B(n6), .Y(SUM[16]) );
  XOR2X2 U59 ( .A(B[16]), .B(A[16]), .Y(n6) );
  OR2X2 U60 ( .A(A[15]), .B(B[15]), .Y(n74) );
  INVX1 U61 ( .A(B[0]), .Y(n123) );
  OAI21XL U62 ( .A0(n118), .A1(n71), .B0(n70), .Y(n12) );
  AOI21X1 U63 ( .A0(n67), .A1(n68), .B0(n69), .Y(n62) );
  INVX1 U64 ( .A(n84), .Y(n15) );
  XOR2X1 U65 ( .A(n12), .B(n13), .Y(SUM[8]) );
  NOR2BX1 U66 ( .AN(n14), .B(n15), .Y(n13) );
  OAI21XL U67 ( .A0(n110), .A1(n11), .B0(n10), .Y(n106) );
  INVX1 U68 ( .A(n8), .Y(n110) );
  NAND4X1 U69 ( .A(n34), .B(n115), .C(n116), .D(n117), .Y(n71) );
  NAND3X1 U70 ( .A(n100), .B(n81), .C(n82), .Y(n66) );
  OAI211X1 U71 ( .A0(n11), .A1(n14), .B0(n10), .C0(n101), .Y(n100) );
  OR2X2 U72 ( .A(B[8]), .B(A[8]), .Y(n84) );
  INVX1 U73 ( .A(n115), .Y(n27) );
  NOR2BX1 U74 ( .AN(n79), .B(n98), .Y(n97) );
  NAND2BX1 U75 ( .AN(n19), .B(n112), .Y(n70) );
  NAND3X1 U76 ( .A(n113), .B(n23), .C(n20), .Y(n112) );
  NAND2BX1 U77 ( .AN(n22), .B(n114), .Y(n113) );
  OAI21XL U78 ( .A0(n27), .A1(n32), .B0(n28), .Y(n114) );
  INVX1 U79 ( .A(n83), .Y(n11) );
  INVX1 U80 ( .A(n116), .Y(n22) );
  NAND2X1 U81 ( .A(B[8]), .B(A[8]), .Y(n14) );
  AND2X1 U82 ( .A(n66), .B(n65), .Y(n64) );
  XOR2X1 U83 ( .A(n93), .B(n94), .Y(SUM[13]) );
  XOR2X1 U84 ( .A(n106), .B(n108), .Y(SUM[10]) );
  NOR2BX1 U85 ( .AN(n101), .B(n109), .Y(n108) );
  INVX1 U86 ( .A(n81), .Y(n109) );
  XOR2X1 U87 ( .A(n104), .B(n105), .Y(SUM[11]) );
  AOI21X1 U88 ( .A0(n81), .A1(n106), .B0(n107), .Y(n105) );
  XOR2X1 U89 ( .A(n8), .B(n9), .Y(SUM[9]) );
  NOR2BXL U90 ( .AN(n10), .B(n11), .Y(n9) );
  OAI21XL U91 ( .A0(n120), .A1(n4), .B0(n38), .Y(n68) );
  AOI21X1 U92 ( .A0(n44), .A1(n121), .B0(n122), .Y(n120) );
  INVX1 U93 ( .A(n41), .Y(n122) );
  OAI21XL U94 ( .A0(n50), .A1(n51), .B0(n46), .Y(n121) );
  OAI21XL U95 ( .A0(n26), .A1(n27), .B0(n28), .Y(n24) );
  INVX1 U96 ( .A(n29), .Y(n26) );
  OAI21XL U97 ( .A0(n31), .A1(n118), .B0(n32), .Y(n29) );
  INVX1 U98 ( .A(n47), .Y(n50) );
  XOR2X1 U99 ( .A(n24), .B(n25), .Y(SUM[6]) );
  XOR2X1 U100 ( .A(n16), .B(n17), .Y(SUM[7]) );
  NOR2X1 U101 ( .A(n18), .B(n19), .Y(n17) );
  OAI21XL U102 ( .A0(n21), .A1(n22), .B0(n23), .Y(n16) );
  INVX1 U103 ( .A(n20), .Y(n18) );
  XOR2X1 U104 ( .A(n35), .B(n36), .Y(SUM[3]) );
  OAI21XL U105 ( .A0(n39), .A1(n40), .B0(n41), .Y(n35) );
  NOR2X1 U106 ( .A(n37), .B(n4), .Y(n36) );
  INVX1 U107 ( .A(n42), .Y(n39) );
  NAND2X1 U108 ( .A(n45), .B(n46), .Y(n42) );
  INVX1 U109 ( .A(n34), .Y(n31) );
  XOR2X1 U110 ( .A(n29), .B(n30), .Y(SUM[5]) );
  XOR2X1 U111 ( .A(n68), .B(n33), .Y(SUM[4]) );
  NOR2BX1 U112 ( .AN(n32), .B(n31), .Y(n33) );
  XOR2X1 U113 ( .A(n48), .B(n49), .Y(SUM[1]) );
  XOR2X1 U114 ( .A(n42), .B(n43), .Y(SUM[2]) );
  NOR2BX1 U115 ( .AN(n41), .B(n40), .Y(n43) );
  INVX1 U116 ( .A(n51), .Y(n48) );
  INVXL U117 ( .A(n79), .Y(n78) );
  OR2X2 U118 ( .A(B[7]), .B(A[7]), .Y(n117) );
  NAND2XL U119 ( .A(B[9]), .B(A[9]), .Y(n10) );
  OR2X2 U120 ( .A(B[6]), .B(A[6]), .Y(n116) );
  OR2X2 U121 ( .A(B[5]), .B(A[5]), .Y(n115) );
  INVX1 U122 ( .A(n74), .Y(n87) );
  XOR2X1 U123 ( .A(n90), .B(n91), .Y(SUM[14]) );
  NOR2BX1 U124 ( .AN(n80), .B(n89), .Y(n91) );
  NAND2XL U125 ( .A(B[13]), .B(A[13]), .Y(n92) );
  NAND2X1 U126 ( .A(B[4]), .B(A[4]), .Y(n32) );
  NAND2X1 U127 ( .A(B[2]), .B(A[2]), .Y(n41) );
  OR2X2 U128 ( .A(B[2]), .B(A[2]), .Y(n44) );
  NAND2X1 U129 ( .A(B[3]), .B(A[3]), .Y(n38) );
  OR2X2 U130 ( .A(B[1]), .B(A[1]), .Y(n47) );
  NAND2X1 U131 ( .A(B[0]), .B(A[0]), .Y(n51) );
  NAND2X1 U132 ( .A(n123), .B(n124), .Y(n119) );
  INVX1 U133 ( .A(A[0]), .Y(n124) );
  NAND2XL U134 ( .A(B[15]), .B(A[15]), .Y(n54) );
  NAND3BX1 U135 ( .AN(n56), .B(n57), .C(n58), .Y(n55) );
  OAI21XL U136 ( .A0(n62), .A1(n63), .B0(n64), .Y(n57) );
  INVX1 U137 ( .A(n80), .Y(n72) );
  NOR2XL U138 ( .A(B[14]), .B(A[14]), .Y(n77) );
  NOR2X1 U139 ( .A(A[15]), .B(B[15]), .Y(n56) );
  NOR2BX1 U140 ( .AN(n92), .B(n7), .Y(n94) );
endmodule


module butterfly_DW01_add_38 ( A, B, SUM );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  wire   n2, n3, n4, n5, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127;

  NAND2X4 U2 ( .A(n94), .B(n77), .Y(n92) );
  NAND2X4 U3 ( .A(n95), .B(n58), .Y(n94) );
  OAI21X4 U4 ( .A0(n90), .A1(n5), .B0(n91), .Y(n88) );
  INVX4 U5 ( .A(n92), .Y(n90) );
  NAND3X2 U6 ( .A(n98), .B(n63), .C(n64), .Y(n95) );
  NAND2X2 U7 ( .A(n80), .B(n99), .Y(n64) );
  NAND2BX1 U8 ( .AN(A[11]), .B(n105), .Y(n80) );
  NAND2X1 U9 ( .A(B[14]), .B(A[14]), .Y(n78) );
  NAND4X1 U10 ( .A(n103), .B(n81), .C(n79), .D(n104), .Y(n98) );
  NAND2BX1 U11 ( .AN(A[11]), .B(n105), .Y(n104) );
  NAND2X1 U12 ( .A(B[12]), .B(A[12]), .Y(n77) );
  OR2X2 U13 ( .A(B[12]), .B(A[12]), .Y(n58) );
  XOR2X2 U14 ( .A(n83), .B(n84), .Y(SUM[15]) );
  NOR2BX1 U15 ( .AN(n52), .B(n85), .Y(n84) );
  AND2X2 U16 ( .A(n50), .B(n122), .Y(SUM[0]) );
  XOR2X2 U17 ( .A(n88), .B(n89), .Y(SUM[14]) );
  NOR2BX2 U18 ( .AN(n91), .B(n5), .Y(n93) );
  NAND2X1 U19 ( .A(B[13]), .B(A[13]), .Y(n91) );
  XNOR2X4 U20 ( .A(B[16]), .B(A[16]), .Y(n4) );
  NAND2XL U21 ( .A(n58), .B(n59), .Y(n57) );
  INVX4 U22 ( .A(n59), .Y(n87) );
  INVX1 U23 ( .A(n72), .Y(n85) );
  OAI21XL U24 ( .A0(n121), .A1(n69), .B0(n68), .Y(n11) );
  XOR2X2 U25 ( .A(n92), .B(n93), .Y(SUM[13]) );
  NOR2BX4 U26 ( .AN(n78), .B(n87), .Y(n89) );
  OAI21XL U27 ( .A0(n113), .A1(n10), .B0(n9), .Y(n109) );
  XOR2X1 U28 ( .A(n7), .B(n8), .Y(SUM[9]) );
  NOR2X2 U29 ( .A(A[13]), .B(B[13]), .Y(n5) );
  AOI21XL U30 ( .A0(n73), .A1(n74), .B0(n75), .Y(n71) );
  NAND2X1 U31 ( .A(B[8]), .B(A[8]), .Y(n13) );
  XNOR2X4 U32 ( .A(n3), .B(n4), .Y(SUM[16]) );
  NAND2BXL U33 ( .AN(n87), .B(n88), .Y(n86) );
  NAND2XL U34 ( .A(n86), .B(n78), .Y(n83) );
  NAND2XL U35 ( .A(n11), .B(n82), .Y(n114) );
  INVXL U36 ( .A(n81), .Y(n10) );
  INVXL U37 ( .A(n120), .Y(n18) );
  NOR2BXL U38 ( .AN(n13), .B(n14), .Y(n12) );
  INVXL U39 ( .A(n69), .Y(n65) );
  INVXL U40 ( .A(n68), .Y(n67) );
  NOR2BXL U41 ( .AN(n22), .B(n21), .Y(n24) );
  NOR2BXL U42 ( .AN(n27), .B(n26), .Y(n29) );
  INVXL U43 ( .A(n37), .Y(n36) );
  NOR2XL U44 ( .A(n17), .B(n18), .Y(n16) );
  INVXL U45 ( .A(n23), .Y(n20) );
  INVXL U46 ( .A(n66), .Y(n121) );
  NOR2BXL U47 ( .AN(n45), .B(n49), .Y(n48) );
  NAND2XL U48 ( .A(n46), .B(n47), .Y(n44) );
  INVXL U49 ( .A(n43), .Y(n39) );
  NAND2XL U50 ( .A(B[13]), .B(A[13]), .Y(n73) );
  NOR2XL U51 ( .A(n5), .B(n57), .Y(n56) );
  OR2X4 U52 ( .A(B[10]), .B(A[10]), .Y(n79) );
  OR2X2 U53 ( .A(A[15]), .B(B[15]), .Y(n72) );
  NAND2XL U54 ( .A(n80), .B(n63), .Y(n107) );
  AOI21XL U55 ( .A0(n79), .A1(n109), .B0(n110), .Y(n108) );
  INVXL U56 ( .A(n101), .Y(n110) );
  NAND2X1 U57 ( .A(B[9]), .B(A[9]), .Y(n9) );
  NAND4XL U58 ( .A(n79), .B(n80), .C(n81), .D(n82), .Y(n61) );
  NAND2XL U59 ( .A(B[6]), .B(A[6]), .Y(n22) );
  NAND2XL U60 ( .A(B[5]), .B(A[5]), .Y(n27) );
  NAND2XL U61 ( .A(B[7]), .B(A[7]), .Y(n19) );
  NAND2XL U62 ( .A(B[1]), .B(A[1]), .Y(n45) );
  NOR2X1 U63 ( .A(B[3]), .B(A[3]), .Y(n2) );
  OR2XL U64 ( .A(B[4]), .B(A[4]), .Y(n33) );
  NAND3X1 U65 ( .A(n52), .B(n53), .C(n51), .Y(n3) );
  NAND2XL U66 ( .A(B[11]), .B(A[11]), .Y(n63) );
  INVX1 U67 ( .A(n11), .Y(n106) );
  INVX1 U68 ( .A(n41), .Y(n38) );
  XOR2X1 U69 ( .A(n11), .B(n12), .Y(SUM[8]) );
  XOR2X1 U70 ( .A(n109), .B(n111), .Y(SUM[10]) );
  NOR2BX1 U71 ( .AN(n101), .B(n112), .Y(n111) );
  INVX1 U72 ( .A(n79), .Y(n112) );
  NOR2BX1 U73 ( .AN(n9), .B(n10), .Y(n8) );
  INVX1 U74 ( .A(n7), .Y(n113) );
  NAND4X1 U75 ( .A(n33), .B(n118), .C(n119), .D(n120), .Y(n69) );
  INVX1 U76 ( .A(n118), .Y(n26) );
  NAND2BX1 U77 ( .AN(n18), .B(n115), .Y(n68) );
  NAND3X1 U78 ( .A(n116), .B(n22), .C(n19), .Y(n115) );
  NAND2BX1 U79 ( .AN(n21), .B(n117), .Y(n116) );
  OAI21XL U80 ( .A0(n26), .A1(n31), .B0(n27), .Y(n117) );
  INVX1 U81 ( .A(n119), .Y(n21) );
  INVX1 U82 ( .A(n82), .Y(n14) );
  NAND2X1 U83 ( .A(n114), .B(n13), .Y(n7) );
  INVX1 U84 ( .A(B[11]), .Y(n105) );
  XOR2X1 U85 ( .A(n23), .B(n24), .Y(SUM[6]) );
  XOR2X1 U86 ( .A(n28), .B(n29), .Y(SUM[5]) );
  XOR2X1 U87 ( .A(n15), .B(n16), .Y(SUM[7]) );
  OAI21XL U88 ( .A0(n20), .A1(n21), .B0(n22), .Y(n15) );
  OAI21XL U89 ( .A0(n25), .A1(n26), .B0(n27), .Y(n23) );
  INVX1 U90 ( .A(n28), .Y(n25) );
  OAI21XL U91 ( .A0(n30), .A1(n121), .B0(n31), .Y(n28) );
  AOI21X1 U92 ( .A0(n65), .A1(n66), .B0(n67), .Y(n60) );
  INVX1 U93 ( .A(n33), .Y(n30) );
  INVX1 U94 ( .A(n46), .Y(n49) );
  INVX1 U95 ( .A(n19), .Y(n17) );
  XOR2X1 U96 ( .A(n66), .B(n32), .Y(SUM[4]) );
  NOR2BX1 U97 ( .AN(n31), .B(n30), .Y(n32) );
  XOR2X1 U98 ( .A(n41), .B(n42), .Y(SUM[2]) );
  NOR2BX1 U99 ( .AN(n40), .B(n39), .Y(n42) );
  XOR2X1 U100 ( .A(n34), .B(n35), .Y(SUM[3]) );
  NOR2X1 U101 ( .A(n36), .B(n2), .Y(n35) );
  OAI21XL U102 ( .A0(n38), .A1(n39), .B0(n40), .Y(n34) );
  NAND2X1 U103 ( .A(n44), .B(n45), .Y(n41) );
  XOR2X1 U104 ( .A(n47), .B(n48), .Y(SUM[1]) );
  XOR2X1 U105 ( .A(n107), .B(n108), .Y(SUM[11]) );
  OR2X2 U106 ( .A(B[9]), .B(A[9]), .Y(n81) );
  OR2X2 U107 ( .A(B[8]), .B(A[8]), .Y(n82) );
  OAI21XL U108 ( .A0(A[13]), .A1(B[13]), .B0(n76), .Y(n74) );
  INVXL U109 ( .A(n77), .Y(n76) );
  NAND3BX1 U110 ( .AN(n54), .B(n55), .C(n56), .Y(n53) );
  OAI21XL U111 ( .A0(n60), .A1(n61), .B0(n62), .Y(n55) );
  XOR2X1 U112 ( .A(n95), .B(n96), .Y(SUM[12]) );
  NOR2BX1 U113 ( .AN(n77), .B(n97), .Y(n96) );
  INVXL U114 ( .A(n58), .Y(n97) );
  NAND2X1 U115 ( .A(n100), .B(n101), .Y(n99) );
  NAND3X1 U116 ( .A(n102), .B(n81), .C(n79), .Y(n100) );
  NAND2X1 U117 ( .A(n9), .B(n13), .Y(n102) );
  OAI21XL U118 ( .A0(n70), .A1(n71), .B0(n72), .Y(n51) );
  INVXL U119 ( .A(n78), .Y(n70) );
  NAND2XL U120 ( .A(B[10]), .B(A[10]), .Y(n101) );
  OR2X2 U121 ( .A(B[7]), .B(A[7]), .Y(n120) );
  OR2X2 U122 ( .A(B[6]), .B(A[6]), .Y(n119) );
  OR2X2 U123 ( .A(B[5]), .B(A[5]), .Y(n118) );
  OR2X4 U124 ( .A(A[14]), .B(B[14]), .Y(n59) );
  NOR2XL U125 ( .A(B[14]), .B(A[14]), .Y(n75) );
  AND2X1 U126 ( .A(n64), .B(n63), .Y(n62) );
  OAI21XL U127 ( .A0(n123), .A1(n2), .B0(n37), .Y(n66) );
  AOI21X1 U128 ( .A0(n43), .A1(n124), .B0(n125), .Y(n123) );
  INVX1 U129 ( .A(n40), .Y(n125) );
  OAI21XL U130 ( .A0(n49), .A1(n50), .B0(n45), .Y(n124) );
  NAND2X1 U131 ( .A(B[4]), .B(A[4]), .Y(n31) );
  NAND2X1 U132 ( .A(B[2]), .B(A[2]), .Y(n40) );
  OR2X2 U133 ( .A(B[2]), .B(A[2]), .Y(n43) );
  NAND2X1 U134 ( .A(B[3]), .B(A[3]), .Y(n37) );
  OR2X2 U135 ( .A(B[1]), .B(A[1]), .Y(n46) );
  NAND2X1 U136 ( .A(n126), .B(n127), .Y(n122) );
  INVX1 U137 ( .A(B[0]), .Y(n126) );
  INVX1 U138 ( .A(n50), .Y(n47) );
  NOR2X1 U139 ( .A(n106), .B(n14), .Y(n103) );
  NAND2X1 U140 ( .A(B[0]), .B(A[0]), .Y(n50) );
  INVX1 U141 ( .A(A[0]), .Y(n127) );
  NAND2X1 U142 ( .A(B[15]), .B(A[15]), .Y(n52) );
  NOR2XL U143 ( .A(A[15]), .B(B[15]), .Y(n54) );
endmodule


module butterfly_DW01_add_48 ( A, B, SUM );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  wire   n1, n2, n3, n4, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142;

  OR2XL U2 ( .A(n96), .B(n97), .Y(n1) );
  NAND2XL U3 ( .A(n1), .B(n98), .Y(n92) );
  AOI21XL U4 ( .A0(n80), .A1(n99), .B0(n76), .Y(n98) );
  NAND2X1 U5 ( .A(n71), .B(n113), .Y(n2) );
  INVX1 U6 ( .A(n114), .Y(n3) );
  AND2X4 U7 ( .A(n2), .B(n3), .Y(n112) );
  XOR2X4 U8 ( .A(n111), .B(n112), .Y(SUM[13]) );
  OR2X2 U9 ( .A(A[12]), .B(B[12]), .Y(n71) );
  INVX1 U10 ( .A(n79), .Y(n119) );
  INVX2 U11 ( .A(n80), .Y(n96) );
  XOR2X1 U12 ( .A(n122), .B(n123), .Y(SUM[11]) );
  OR2X2 U13 ( .A(B[15]), .B(A[15]), .Y(n66) );
  INVX1 U14 ( .A(A[13]), .Y(n101) );
  CLKINVX3 U15 ( .A(n71), .Y(n67) );
  OR2X2 U16 ( .A(B[14]), .B(A[14]), .Y(n90) );
  NAND2X1 U17 ( .A(n116), .B(n78), .Y(n113) );
  NAND2X1 U18 ( .A(n127), .B(n128), .Y(n79) );
  INVX1 U19 ( .A(n66), .Y(n64) );
  XNOR2X1 U20 ( .A(n54), .B(n7), .Y(SUM[16]) );
  NAND2X1 U21 ( .A(B[14]), .B(A[14]), .Y(n4) );
  AND2X2 U22 ( .A(n53), .B(n137), .Y(SUM[0]) );
  NAND2X1 U23 ( .A(n73), .B(n63), .Y(n111) );
  NAND2X1 U24 ( .A(n55), .B(n56), .Y(n54) );
  AOI21X1 U25 ( .A0(n100), .A1(n101), .B0(n67), .Y(n104) );
  XNOR2X1 U26 ( .A(B[16]), .B(A[16]), .Y(n7) );
  AOI21X1 U27 ( .A0(n57), .A1(n58), .B0(n59), .Y(n56) );
  NOR2X1 U28 ( .A(n64), .B(n65), .Y(n57) );
  INVX1 U29 ( .A(n73), .Y(n61) );
  NOR2X1 U30 ( .A(A[13]), .B(B[13]), .Y(n94) );
  NAND2X2 U31 ( .A(B[13]), .B(A[13]), .Y(n63) );
  OR2X2 U32 ( .A(B[11]), .B(A[11]), .Y(n80) );
  AOI21X1 U33 ( .A0(n91), .A1(n92), .B0(n93), .Y(n89) );
  INVX2 U34 ( .A(n90), .Y(n65) );
  INVX2 U35 ( .A(B[13]), .Y(n100) );
  OAI21XL U36 ( .A0(n107), .A1(n108), .B0(n63), .Y(n106) );
  OAI21X1 U37 ( .A0(n94), .A1(n95), .B0(n63), .Y(n93) );
  OAI211XL U38 ( .A0(n61), .A1(n62), .B0(n63), .C0(n4), .Y(n58) );
  INVX1 U39 ( .A(A[10]), .Y(n128) );
  INVX1 U40 ( .A(B[10]), .Y(n127) );
  OR2XL U41 ( .A(B[2]), .B(A[2]), .Y(n46) );
  NAND4XL U42 ( .A(n79), .B(n80), .C(n81), .D(n16), .Y(n68) );
  INVX1 U43 ( .A(n110), .Y(n76) );
  INVXL U44 ( .A(n78), .Y(n77) );
  NOR2XL U45 ( .A(n61), .B(n65), .Y(n72) );
  OAI21X1 U46 ( .A0(n136), .A1(n69), .B0(n85), .Y(n12) );
  INVXL U47 ( .A(n83), .Y(n136) );
  INVXL U48 ( .A(n69), .Y(n82) );
  INVXL U49 ( .A(n85), .Y(n84) );
  XOR2X1 U50 ( .A(n113), .B(n115), .Y(SUM[12]) );
  AOI21XL U51 ( .A0(n82), .A1(n83), .B0(n84), .Y(n74) );
  NOR2X1 U52 ( .A(n76), .B(n77), .Y(n75) );
  NOR2BX1 U53 ( .AN(n110), .B(n121), .Y(n116) );
  XOR2X1 U54 ( .A(n125), .B(n126), .Y(SUM[10]) );
  NOR2BX1 U55 ( .AN(n118), .B(n119), .Y(n126) );
  NAND4XL U56 ( .A(n16), .B(n12), .C(n81), .D(n79), .Y(n97) );
  NOR2XL U57 ( .A(n19), .B(n20), .Y(n18) );
  INVXL U58 ( .A(n25), .Y(n22) );
  INVXL U59 ( .A(n31), .Y(n28) );
  AOI21XL U60 ( .A0(n46), .A1(n139), .B0(n140), .Y(n138) );
  NOR2BXL U61 ( .AN(n30), .B(n29), .Y(n32) );
  NAND2XL U62 ( .A(n49), .B(n50), .Y(n47) );
  NOR2BXL U63 ( .AN(n34), .B(n33), .Y(n35) );
  NOR2BXL U64 ( .AN(n48), .B(n52), .Y(n51) );
  OR2XL U65 ( .A(B[8]), .B(A[8]), .Y(n16) );
  OR2XL U66 ( .A(B[9]), .B(A[9]), .Y(n81) );
  NAND2XL U67 ( .A(B[10]), .B(A[10]), .Y(n118) );
  NAND2XL U68 ( .A(B[6]), .B(A[6]), .Y(n24) );
  NAND2XL U69 ( .A(B[8]), .B(A[8]), .Y(n14) );
  NAND2XL U70 ( .A(B[7]), .B(A[7]), .Y(n21) );
  OR2XL U71 ( .A(B[6]), .B(A[6]), .Y(n27) );
  OR2XL U72 ( .A(B[7]), .B(A[7]), .Y(n135) );
  NAND2XL U73 ( .A(B[2]), .B(A[2]), .Y(n43) );
  NAND2XL U74 ( .A(B[4]), .B(A[4]), .Y(n34) );
  NAND2XL U75 ( .A(B[5]), .B(A[5]), .Y(n30) );
  NAND2XL U76 ( .A(B[3]), .B(A[3]), .Y(n40) );
  NOR2XL U77 ( .A(B[3]), .B(A[3]), .Y(n6) );
  OR2XL U78 ( .A(B[4]), .B(A[4]), .Y(n36) );
  OR2XL U79 ( .A(B[5]), .B(A[5]), .Y(n134) );
  NAND2XL U80 ( .A(B[1]), .B(A[1]), .Y(n48) );
  NAND2BX1 U81 ( .AN(n96), .B(n99), .Y(n78) );
  OAI21XL U82 ( .A0(n138), .A1(n6), .B0(n40), .Y(n83) );
  INVX1 U83 ( .A(n43), .Y(n140) );
  OAI21XL U84 ( .A0(n52), .A1(n53), .B0(n48), .Y(n139) );
  OAI21XL U85 ( .A0(n11), .A1(n129), .B0(n10), .Y(n125) );
  INVX1 U86 ( .A(n8), .Y(n129) );
  OAI21XL U87 ( .A0(n28), .A1(n29), .B0(n30), .Y(n25) );
  OAI21XL U88 ( .A0(n33), .A1(n136), .B0(n34), .Y(n31) );
  NAND2X1 U89 ( .A(n117), .B(n118), .Y(n99) );
  NAND2BX1 U90 ( .AN(n119), .B(n120), .Y(n117) );
  OAI21XL U91 ( .A0(n11), .A1(n14), .B0(n10), .Y(n120) );
  NAND4X1 U92 ( .A(n36), .B(n134), .C(n27), .D(n135), .Y(n69) );
  INVX1 U93 ( .A(n81), .Y(n11) );
  OAI21XL U94 ( .A0(n96), .A1(n97), .B0(n109), .Y(n105) );
  AOI21XL U95 ( .A0(n80), .A1(n99), .B0(n76), .Y(n109) );
  INVX1 U96 ( .A(n134), .Y(n29) );
  OAI21X1 U97 ( .A0(n124), .A1(n119), .B0(n118), .Y(n122) );
  NOR2BX1 U98 ( .AN(n110), .B(n96), .Y(n123) );
  INVX1 U99 ( .A(n125), .Y(n124) );
  AOI21X1 U100 ( .A0(n100), .A1(n101), .B0(n67), .Y(n91) );
  XOR2X1 U101 ( .A(n12), .B(n13), .Y(SUM[8]) );
  NOR2BX1 U102 ( .AN(n14), .B(n15), .Y(n13) );
  INVX1 U103 ( .A(n16), .Y(n15) );
  NOR2BX1 U104 ( .AN(n62), .B(n67), .Y(n115) );
  XOR2X1 U105 ( .A(n8), .B(n9), .Y(SUM[9]) );
  NOR2BXL U106 ( .AN(n10), .B(n11), .Y(n9) );
  XOR2X1 U107 ( .A(n31), .B(n32), .Y(SUM[5]) );
  XOR2X1 U108 ( .A(n17), .B(n18), .Y(SUM[7]) );
  OAI21XL U109 ( .A0(n22), .A1(n23), .B0(n24), .Y(n17) );
  XOR2X1 U110 ( .A(n25), .B(n26), .Y(SUM[6]) );
  NOR2BX1 U111 ( .AN(n24), .B(n23), .Y(n26) );
  XOR2X2 U112 ( .A(n102), .B(n103), .Y(SUM[14]) );
  NAND2X1 U113 ( .A(n90), .B(n4), .Y(n102) );
  AOI21X2 U114 ( .A0(n104), .A1(n105), .B0(n106), .Y(n103) );
  OAI21XL U115 ( .A0(n74), .A1(n68), .B0(n75), .Y(n70) );
  NAND2BX1 U116 ( .AN(n20), .B(n131), .Y(n85) );
  NAND3X1 U117 ( .A(n132), .B(n24), .C(n21), .Y(n131) );
  NAND2X1 U118 ( .A(n133), .B(n27), .Y(n132) );
  OAI21XL U119 ( .A0(n29), .A1(n34), .B0(n30), .Y(n133) );
  INVX1 U120 ( .A(n27), .Y(n23) );
  INVX1 U121 ( .A(n36), .Y(n33) );
  INVX1 U122 ( .A(n49), .Y(n52) );
  NOR2X1 U123 ( .A(n96), .B(n97), .Y(n121) );
  NAND2X1 U124 ( .A(n130), .B(n14), .Y(n8) );
  NAND2X1 U125 ( .A(n12), .B(n16), .Y(n130) );
  INVX1 U126 ( .A(n135), .Y(n20) );
  INVX1 U127 ( .A(n21), .Y(n19) );
  XOR2X1 U128 ( .A(n50), .B(n51), .Y(SUM[1]) );
  XOR2X1 U129 ( .A(n37), .B(n38), .Y(SUM[3]) );
  OAI21XL U130 ( .A0(n41), .A1(n42), .B0(n43), .Y(n37) );
  NOR2X1 U131 ( .A(n39), .B(n6), .Y(n38) );
  INVX1 U132 ( .A(n44), .Y(n41) );
  XOR2X1 U133 ( .A(n44), .B(n45), .Y(SUM[2]) );
  NOR2BX1 U134 ( .AN(n43), .B(n42), .Y(n45) );
  XOR2X1 U135 ( .A(n83), .B(n35), .Y(SUM[4]) );
  NAND2X1 U136 ( .A(n47), .B(n48), .Y(n44) );
  INVX1 U137 ( .A(n46), .Y(n42) );
  INVX1 U138 ( .A(n40), .Y(n39) );
  INVX1 U139 ( .A(n53), .Y(n50) );
  NAND2XL U140 ( .A(B[9]), .B(A[9]), .Y(n10) );
  XOR2X2 U141 ( .A(n86), .B(n87), .Y(SUM[15]) );
  NOR2X2 U142 ( .A(n89), .B(n65), .Y(n88) );
  OR2X2 U143 ( .A(B[1]), .B(A[1]), .Y(n49) );
  NAND2X1 U144 ( .A(B[0]), .B(A[0]), .Y(n53) );
  NAND2X1 U145 ( .A(n141), .B(n142), .Y(n137) );
  INVX1 U146 ( .A(A[0]), .Y(n142) );
  INVX1 U147 ( .A(B[0]), .Y(n141) );
  NAND4XL U148 ( .A(n70), .B(n71), .C(n66), .D(n72), .Y(n55) );
  INVX1 U149 ( .A(n60), .Y(n59) );
  NAND2X1 U150 ( .A(n60), .B(n66), .Y(n86) );
  NAND2XL U151 ( .A(B[15]), .B(A[15]), .Y(n60) );
  INVXL U152 ( .A(n62), .Y(n114) );
  NAND2XL U153 ( .A(A[12]), .B(B[12]), .Y(n108) );
  NAND2XL U154 ( .A(A[12]), .B(B[12]), .Y(n95) );
  NAND2XL U155 ( .A(B[12]), .B(A[12]), .Y(n62) );
  NAND2XL U156 ( .A(B[11]), .B(A[11]), .Y(n110) );
  NOR2XL U157 ( .A(A[13]), .B(B[13]), .Y(n107) );
  NAND2BX1 U158 ( .AN(A[13]), .B(n100), .Y(n73) );
  NOR2BX4 U159 ( .AN(n4), .B(n88), .Y(n87) );
endmodule


module butterfly_DW01_sub_37 ( A, B, DIFF );
  input [16:0] A;
  input [16:0] B;
  output [16:0] DIFF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n11, n12, n13, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176;

  INVX1 U3 ( .A(n117), .Y(n2) );
  NAND2BX2 U4 ( .AN(B[15]), .B(A[15]), .Y(n101) );
  NAND2X1 U5 ( .A(B[9]), .B(n151), .Y(n94) );
  XOR2X2 U6 ( .A(B[16]), .B(A[16]), .Y(n13) );
  NOR2BX2 U7 ( .AN(B[13]), .B(A[13]), .Y(n128) );
  INVX2 U8 ( .A(n92), .Y(n103) );
  NAND3X2 U9 ( .A(n120), .B(n75), .C(n76), .Y(n125) );
  NAND2X2 U10 ( .A(n97), .B(n121), .Y(n76) );
  NAND2X2 U11 ( .A(n1), .B(n2), .Y(n3) );
  NAND2X2 U12 ( .A(n3), .B(n105), .Y(n126) );
  INVX2 U13 ( .A(n127), .Y(n1) );
  NOR2BX4 U14 ( .AN(B[13]), .B(A[13]), .Y(n127) );
  AOI21X2 U15 ( .A0(n124), .A1(n125), .B0(n126), .Y(n122) );
  NAND2X2 U16 ( .A(B[12]), .B(n133), .Y(n85) );
  INVX2 U17 ( .A(n85), .Y(n129) );
  OAI21X1 U18 ( .A0(n112), .A1(n113), .B0(n106), .Y(n109) );
  INVX1 U19 ( .A(n92), .Y(n91) );
  OAI21X1 U20 ( .A0(n153), .A1(n81), .B0(n80), .Y(n23) );
  NAND2BX1 U21 ( .AN(A[10]), .B(B[10]), .Y(n96) );
  INVX1 U22 ( .A(A[12]), .Y(n133) );
  INVX1 U23 ( .A(B[14]), .Y(n114) );
  NAND2BX1 U24 ( .AN(A[11]), .B(B[11]), .Y(n97) );
  OAI2BB2X1 U25 ( .B0(n114), .B1(A[14]), .A0N(n17), .A1N(B[13]), .Y(n113) );
  NAND2BXL U26 ( .AN(A[14]), .B(B[14]), .Y(n86) );
  NAND2BX2 U27 ( .AN(A[15]), .B(B[15]), .Y(n92) );
  NAND2XL U28 ( .A(n131), .B(n117), .Y(n9) );
  NAND2XL U29 ( .A(n117), .B(n118), .Y(n116) );
  INVX2 U30 ( .A(n117), .Y(n108) );
  NAND2BXL U31 ( .AN(A[11]), .B(B[11]), .Y(n141) );
  NAND2BX1 U32 ( .AN(B[11]), .B(A[11]), .Y(n75) );
  AOI21X1 U33 ( .A0(n96), .A1(n145), .B0(n139), .Y(n144) );
  XNOR2X2 U34 ( .A(n9), .B(n130), .Y(DIFF[13]) );
  NAND2X1 U35 ( .A(n122), .B(n5), .Y(n6) );
  XOR2X2 U36 ( .A(n109), .B(n11), .Y(DIFF[15]) );
  NAND2BX2 U37 ( .AN(B[13]), .B(A[13]), .Y(n105) );
  NOR2X2 U38 ( .A(n108), .B(n129), .Y(n132) );
  NAND2X2 U39 ( .A(n4), .B(n123), .Y(n7) );
  NAND2X2 U40 ( .A(n6), .B(n7), .Y(DIFF[14]) );
  INVX1 U41 ( .A(n122), .Y(n4) );
  INVXL U42 ( .A(n123), .Y(n5) );
  XOR2X1 U43 ( .A(B[14]), .B(A[14]), .Y(n123) );
  AND2X1 U44 ( .A(B[14]), .B(n102), .Y(n8) );
  NOR2X1 U45 ( .A(n8), .B(n103), .Y(n99) );
  NOR2BXL U46 ( .AN(A[2]), .B(B[2]), .Y(n16) );
  NAND2XL U47 ( .A(n33), .B(n154), .Y(n80) );
  NAND3BXL U48 ( .AN(n56), .B(n165), .C(n53), .Y(n93) );
  NAND2X2 U49 ( .A(A[12]), .B(n134), .Y(n117) );
  NAND2BXL U50 ( .AN(B[10]), .B(A[10]), .Y(n148) );
  NOR2XL U51 ( .A(B[10]), .B(n21), .Y(n138) );
  NAND2X1 U52 ( .A(A[5]), .B(n159), .Y(n40) );
  INVXL U53 ( .A(n76), .Y(n73) );
  INVXL U54 ( .A(n47), .Y(n153) );
  NAND4XL U55 ( .A(n94), .B(n95), .C(n96), .D(n97), .Y(n71) );
  NAND3XL U56 ( .A(n75), .B(n119), .C(n120), .Y(n115) );
  AND2X2 U57 ( .A(n101), .B(n110), .Y(n11) );
  INVXL U58 ( .A(n22), .Y(n20) );
  NAND2XL U59 ( .A(n88), .B(n89), .Y(n66) );
  NOR3XL U60 ( .A(n71), .B(n81), .C(n93), .Y(n88) );
  INVXL U61 ( .A(n37), .Y(n32) );
  AOI21XL U62 ( .A0(n30), .A1(n31), .B0(n32), .Y(n29) );
  NAND2XL U63 ( .A(n33), .B(n34), .Y(n28) );
  NOR2XL U64 ( .A(n25), .B(n26), .Y(n24) );
  INVXL U65 ( .A(n27), .Y(n25) );
  INVXL U66 ( .A(n44), .Y(n39) );
  NOR2XL U67 ( .A(n43), .B(n39), .Y(n42) );
  NOR2XL U68 ( .A(n16), .B(n56), .Y(n55) );
  NAND2XL U69 ( .A(n53), .B(n54), .Y(n49) );
  AOI21XL U70 ( .A0(n51), .A1(n52), .B0(n16), .Y(n50) );
  NOR2XL U71 ( .A(n61), .B(n15), .Y(n60) );
  INVXL U72 ( .A(n58), .Y(n61) );
  XNOR2X1 U73 ( .A(n47), .B(n12), .Y(DIFF[4]) );
  NAND2XL U74 ( .A(n46), .B(n48), .Y(n12) );
  NOR2XL U75 ( .A(n142), .B(n26), .Y(n140) );
  NOR2XL U76 ( .A(n82), .B(n83), .Y(n68) );
  NAND2X1 U77 ( .A(n135), .B(n136), .Y(n121) );
  NAND2XL U78 ( .A(n22), .B(n27), .Y(n137) );
  INVXL U79 ( .A(A[9]), .Y(n151) );
  INVX1 U80 ( .A(n148), .Y(n139) );
  NAND2XL U81 ( .A(B[6]), .B(n162), .Y(n30) );
  INVXL U82 ( .A(A[6]), .Y(n162) );
  NAND2XL U83 ( .A(B[7]), .B(n161), .Y(n33) );
  INVXL U84 ( .A(B[8]), .Y(n152) );
  INVXL U85 ( .A(B[7]), .Y(n156) );
  INVXL U86 ( .A(B[6]), .Y(n157) );
  NAND2XL U87 ( .A(B[8]), .B(n174), .Y(n95) );
  INVXL U88 ( .A(A[8]), .Y(n174) );
  INVXL U89 ( .A(A[5]), .Y(n163) );
  NAND2XL U90 ( .A(B[2]), .B(n173), .Y(n51) );
  INVXL U91 ( .A(A[2]), .Y(n173) );
  NAND2XL U92 ( .A(B[3]), .B(n170), .Y(n53) );
  NAND2XL U93 ( .A(B[4]), .B(n164), .Y(n48) );
  INVXL U94 ( .A(A[4]), .Y(n164) );
  INVXL U95 ( .A(B[4]), .Y(n160) );
  INVXL U96 ( .A(B[3]), .Y(n169) );
  INVXL U97 ( .A(B[1]), .Y(n172) );
  XNOR2X1 U98 ( .A(n64), .B(n13), .Y(DIFF[16]) );
  INVX1 U99 ( .A(n23), .Y(n142) );
  NAND2BX1 U100 ( .AN(n78), .B(n93), .Y(n47) );
  OAI21XL U101 ( .A0(n70), .A1(n71), .B0(n72), .Y(n69) );
  AOI21X1 U102 ( .A0(n77), .A1(n78), .B0(n79), .Y(n70) );
  NOR2X1 U103 ( .A(n73), .B(n74), .Y(n72) );
  INVX1 U104 ( .A(n81), .Y(n77) );
  XOR2X1 U105 ( .A(n125), .B(n132), .Y(DIFF[12]) );
  INVX1 U106 ( .A(n80), .Y(n79) );
  NAND4X1 U107 ( .A(n48), .B(n44), .C(n30), .D(n33), .Y(n81) );
  OAI21XL U108 ( .A0(n149), .A1(n21), .B0(n22), .Y(n145) );
  INVX1 U109 ( .A(n18), .Y(n149) );
  OAI21XL U110 ( .A0(n38), .A1(n39), .B0(n40), .Y(n31) );
  INVX1 U111 ( .A(n41), .Y(n38) );
  OAI21XL U112 ( .A0(n167), .A1(n168), .B0(n54), .Y(n78) );
  AOI21X1 U113 ( .A0(n51), .A1(n171), .B0(n16), .Y(n167) );
  INVX1 U114 ( .A(n53), .Y(n168) );
  OAI21XL U115 ( .A0(n15), .A1(n62), .B0(n58), .Y(n171) );
  OAI21X1 U116 ( .A0(n26), .A1(n142), .B0(n27), .Y(n18) );
  INVX1 U117 ( .A(n94), .Y(n21) );
  XOR2X1 U118 ( .A(n18), .B(n19), .Y(DIFF[9]) );
  NOR2XL U119 ( .A(n20), .B(n21), .Y(n19) );
  XOR2X1 U120 ( .A(n23), .B(n24), .Y(DIFF[8]) );
  INVX1 U121 ( .A(n95), .Y(n26) );
  NAND3X1 U122 ( .A(n155), .B(n37), .C(n34), .Y(n154) );
  NAND3X1 U123 ( .A(n44), .B(n158), .C(n30), .Y(n155) );
  NAND2XL U124 ( .A(n85), .B(n125), .Y(n131) );
  XOR2X1 U125 ( .A(n143), .B(n144), .Y(DIFF[11]) );
  XOR2X1 U126 ( .A(n145), .B(n146), .Y(DIFF[10]) );
  NOR2X1 U127 ( .A(n147), .B(n139), .Y(n146) );
  INVX1 U128 ( .A(n96), .Y(n147) );
  XOR2X1 U129 ( .A(n31), .B(n35), .Y(DIFF[6]) );
  NOR2X1 U130 ( .A(n32), .B(n36), .Y(n35) );
  INVX1 U131 ( .A(n30), .Y(n36) );
  XOR2X1 U132 ( .A(n28), .B(n29), .Y(DIFF[7]) );
  XOR2X1 U133 ( .A(n41), .B(n42), .Y(DIFF[5]) );
  INVX1 U134 ( .A(n40), .Y(n43) );
  NOR2X1 U135 ( .A(n90), .B(n91), .Y(n89) );
  NAND2X1 U136 ( .A(n45), .B(n46), .Y(n41) );
  NAND2X1 U137 ( .A(n47), .B(n48), .Y(n45) );
  AOI21XL U138 ( .A0(n115), .A1(n85), .B0(n116), .Y(n112) );
  NAND2X1 U139 ( .A(n46), .B(n40), .Y(n158) );
  INVX1 U140 ( .A(n75), .Y(n74) );
  OAI21XL U141 ( .A0(n57), .A1(n15), .B0(n58), .Y(n52) );
  INVX1 U142 ( .A(n59), .Y(n57) );
  NOR2X1 U143 ( .A(n15), .B(n166), .Y(n165) );
  INVX1 U144 ( .A(n63), .Y(n166) );
  INVX1 U145 ( .A(n51), .Y(n56) );
  XOR2X1 U146 ( .A(n52), .B(n55), .Y(DIFF[2]) );
  XOR2X1 U147 ( .A(n49), .B(n50), .Y(DIFF[3]) );
  XOR2X1 U148 ( .A(n59), .B(n60), .Y(DIFF[1]) );
  NAND2BX1 U149 ( .AN(n63), .B(n62), .Y(n59) );
  NAND2X1 U150 ( .A(n62), .B(n63), .Y(DIFF[0]) );
  INVX1 U151 ( .A(B[12]), .Y(n134) );
  NOR2BX1 U152 ( .AN(B[1]), .B(A[1]), .Y(n15) );
  NAND4X1 U153 ( .A(n140), .B(n94), .C(n96), .D(n141), .Y(n120) );
  INVXL U154 ( .A(B[13]), .Y(n107) );
  INVX1 U155 ( .A(A[7]), .Y(n161) );
  NAND2X1 U156 ( .A(B[5]), .B(n163), .Y(n44) );
  NAND2X1 U157 ( .A(A[9]), .B(n150), .Y(n22) );
  INVXL U158 ( .A(B[9]), .Y(n150) );
  INVX1 U159 ( .A(B[5]), .Y(n159) );
  NAND2X1 U160 ( .A(A[8]), .B(n152), .Y(n27) );
  INVX1 U161 ( .A(A[3]), .Y(n170) );
  AOI21X1 U162 ( .A0(n98), .A1(n99), .B0(n100), .Y(n65) );
  INVXL U163 ( .A(n101), .Y(n100) );
  INVXL U164 ( .A(B[15]), .Y(n87) );
  NAND2X1 U165 ( .A(A[7]), .B(n156), .Y(n34) );
  NAND2XL U166 ( .A(B[15]), .B(n111), .Y(n110) );
  NAND2X1 U167 ( .A(A[6]), .B(n157), .Y(n37) );
  NAND3XL U168 ( .A(n137), .B(n94), .C(A[10]), .Y(n136) );
  AOI21X1 U169 ( .A0(n138), .A1(n137), .B0(n139), .Y(n135) );
  NAND2X1 U170 ( .A(A[4]), .B(n160), .Y(n46) );
  NAND2X1 U171 ( .A(A[1]), .B(n172), .Y(n58) );
  NAND2X1 U172 ( .A(A[3]), .B(n169), .Y(n54) );
  NAND2X1 U173 ( .A(B[0]), .B(n175), .Y(n63) );
  INVX1 U174 ( .A(A[0]), .Y(n175) );
  NAND2X1 U175 ( .A(A[0]), .B(n176), .Y(n62) );
  INVX1 U176 ( .A(B[0]), .Y(n176) );
  NAND3X1 U177 ( .A(n65), .B(n66), .C(n67), .Y(n64) );
  NAND2X1 U178 ( .A(n68), .B(n69), .Y(n67) );
  INVXL U179 ( .A(A[14]), .Y(n102) );
  NAND2BXL U180 ( .AN(B[14]), .B(A[14]), .Y(n106) );
  NAND2X1 U181 ( .A(n97), .B(n121), .Y(n119) );
  NAND2X1 U182 ( .A(n97), .B(n75), .Y(n143) );
  INVXL U183 ( .A(A[13]), .Y(n17) );
  INVXL U184 ( .A(A[15]), .Y(n111) );
  NAND2X1 U185 ( .A(n105), .B(n84), .Y(n130) );
  NOR2X1 U186 ( .A(n128), .B(n129), .Y(n124) );
  NAND3XL U187 ( .A(n104), .B(n105), .C(n106), .Y(n98) );
  NAND3XL U188 ( .A(n85), .B(n84), .C(n86), .Y(n90) );
  NAND3XL U189 ( .A(n84), .B(n85), .C(n86), .Y(n83) );
  NAND2BXL U190 ( .AN(A[13]), .B(B[13]), .Y(n84) );
  NOR2XL U191 ( .A(A[15]), .B(n87), .Y(n82) );
  OAI21XL U192 ( .A0(n107), .A1(A[13]), .B0(n108), .Y(n104) );
  NAND2XL U193 ( .A(A[13]), .B(n107), .Y(n118) );
endmodule


module butterfly_DW01_sub_38 ( A, B, DIFF );
  input [16:0] A;
  input [16:0] B;
  output [16:0] DIFF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159;

  INVX2 U3 ( .A(n63), .Y(n72) );
  NAND4X1 U4 ( .A(n68), .B(n69), .C(n70), .D(n71), .Y(n57) );
  AOI21X2 U5 ( .A0(n66), .A1(n98), .B0(n6), .Y(n97) );
  NAND2X1 U6 ( .A(B[13]), .B(n109), .Y(n66) );
  NOR2BX4 U7 ( .AN(A[13]), .B(B[13]), .Y(n6) );
  NAND2BX2 U8 ( .AN(A[15]), .B(B[15]), .Y(n64) );
  AOI21XL U9 ( .A0(n65), .A1(n66), .B0(n6), .Y(n60) );
  NOR2X2 U10 ( .A(n65), .B(n6), .Y(n93) );
  OAI21XL U11 ( .A0(n119), .A1(n75), .B0(n82), .Y(n116) );
  NAND3X1 U12 ( .A(n101), .B(n100), .C(n99), .Y(n98) );
  NAND2X1 U13 ( .A(B[9]), .B(n134), .Y(n114) );
  OAI21XL U14 ( .A0(n136), .A1(n73), .B0(n86), .Y(n13) );
  OAI21XL U15 ( .A0(n16), .A1(n119), .B0(n17), .Y(n8) );
  INVX1 U16 ( .A(n114), .Y(n11) );
  NAND2BX1 U17 ( .AN(n102), .B(n103), .Y(n101) );
  NAND2X2 U18 ( .A(B[14]), .B(n107), .Y(n63) );
  INVX2 U19 ( .A(A[14]), .Y(n107) );
  NAND2X1 U20 ( .A(A[14]), .B(n106), .Y(n61) );
  INVX1 U21 ( .A(B[14]), .Y(n106) );
  AND2X2 U22 ( .A(n121), .B(n122), .Y(n1) );
  NAND2BX2 U23 ( .AN(A[11]), .B(B[11]), .Y(n105) );
  NAND2BX4 U24 ( .AN(A[12]), .B(B[12]), .Y(n111) );
  NAND2BXL U25 ( .AN(B[15]), .B(A[15]), .Y(n67) );
  INVX1 U26 ( .A(A[13]), .Y(n109) );
  NAND3X1 U27 ( .A(n92), .B(n93), .C(n94), .Y(n90) );
  NAND2BXL U28 ( .AN(A[12]), .B(B[12]), .Y(n112) );
  NAND2BX2 U29 ( .AN(B[12]), .B(A[12]), .Y(n100) );
  NOR2BXL U30 ( .AN(n67), .B(n59), .Y(n58) );
  NAND2X1 U31 ( .A(n63), .B(n64), .Y(n62) );
  NAND2X1 U32 ( .A(n104), .B(n103), .Y(n82) );
  AOI21XL U33 ( .A0(n60), .A1(n61), .B0(n62), .Y(n59) );
  XNOR2X2 U34 ( .A(n2), .B(n108), .Y(DIFF[13]) );
  AND3X2 U35 ( .A(n92), .B(n100), .C(n94), .Y(n2) );
  NOR2X2 U36 ( .A(n6), .B(n95), .Y(n108) );
  NOR2X2 U37 ( .A(n65), .B(n118), .Y(n117) );
  INVX2 U38 ( .A(n100), .Y(n65) );
  NAND2X2 U39 ( .A(n1), .B(n120), .Y(n103) );
  NAND2BX1 U40 ( .AN(n110), .B(n103), .Y(n94) );
  NAND2X2 U41 ( .A(B[6]), .B(n145), .Y(n20) );
  INVXL U42 ( .A(A[8]), .Y(n157) );
  NAND2XL U43 ( .A(A[7]), .B(n139), .Y(n24) );
  INVXL U44 ( .A(A[1]), .Y(n155) );
  NOR2X1 U45 ( .A(n72), .B(n95), .Y(n89) );
  INVX1 U46 ( .A(n80), .Y(n118) );
  OAI21XL U47 ( .A0(n132), .A1(n11), .B0(n12), .Y(n126) );
  INVX1 U48 ( .A(n121), .Y(n127) );
  INVXL U49 ( .A(n17), .Y(n15) );
  NAND2XL U50 ( .A(n36), .B(n38), .Y(n3) );
  INVXL U51 ( .A(n49), .Y(n52) );
  NAND2X1 U52 ( .A(B[7]), .B(n144), .Y(n23) );
  NAND2X1 U53 ( .A(B[8]), .B(n157), .Y(n113) );
  INVX1 U54 ( .A(A[9]), .Y(n134) );
  NOR2BX1 U55 ( .AN(A[2]), .B(B[2]), .Y(n7) );
  NAND2X1 U56 ( .A(B[4]), .B(n147), .Y(n38) );
  NAND2X1 U57 ( .A(B[2]), .B(n156), .Y(n41) );
  NAND2X1 U58 ( .A(B[3]), .B(n152), .Y(n43) );
  NOR2XL U59 ( .A(n72), .B(n73), .Y(n70) );
  INVXL U60 ( .A(n37), .Y(n136) );
  INVXL U61 ( .A(n27), .Y(n22) );
  NOR2XL U62 ( .A(n33), .B(n29), .Y(n32) );
  INVXL U63 ( .A(n30), .Y(n33) );
  INVXL U64 ( .A(n73), .Y(n83) );
  NOR2X1 U65 ( .A(n79), .B(n74), .Y(n78) );
  AOI21XL U66 ( .A0(n83), .A1(n84), .B0(n85), .Y(n81) );
  NAND2XL U67 ( .A(n80), .B(n66), .Y(n74) );
  XOR2X1 U68 ( .A(n87), .B(n88), .Y(DIFF[15]) );
  NAND2XL U69 ( .A(n67), .B(n64), .Y(n87) );
  AOI21X1 U70 ( .A0(n89), .A1(n90), .B0(n91), .Y(n88) );
  INVXL U71 ( .A(B[6]), .Y(n140) );
  NAND2X1 U72 ( .A(n23), .B(n137), .Y(n86) );
  NOR2XL U73 ( .A(n75), .B(n76), .Y(n68) );
  NOR2XL U74 ( .A(n15), .B(n16), .Y(n14) );
  AOI21XL U75 ( .A0(n20), .A1(n21), .B0(n22), .Y(n19) );
  AOI21XL U76 ( .A0(n41), .A1(n153), .B0(n7), .Y(n149) );
  NAND4XL U77 ( .A(n43), .B(n41), .C(n54), .D(n148), .Y(n76) );
  NAND2XL U78 ( .A(B[5]), .B(n146), .Y(n34) );
  INVXL U79 ( .A(B[5]), .Y(n142) );
  XNOR2X1 U80 ( .A(n37), .B(n3), .Y(DIFF[4]) );
  NOR2XL U81 ( .A(n7), .B(n46), .Y(n45) );
  NOR2XL U82 ( .A(n52), .B(n48), .Y(n51) );
  NAND2X1 U83 ( .A(B[10]), .B(n130), .Y(n115) );
  NAND2X1 U84 ( .A(A[9]), .B(n133), .Y(n12) );
  INVXL U85 ( .A(B[9]), .Y(n133) );
  NAND2X1 U86 ( .A(A[8]), .B(n135), .Y(n17) );
  INVXL U87 ( .A(B[8]), .Y(n135) );
  INVXL U88 ( .A(B[7]), .Y(n139) );
  INVXL U89 ( .A(A[4]), .Y(n147) );
  NAND2XL U90 ( .A(A[4]), .B(n143), .Y(n36) );
  INVXL U91 ( .A(B[4]), .Y(n143) );
  NAND2XL U92 ( .A(A[3]), .B(n151), .Y(n44) );
  INVXL U93 ( .A(B[3]), .Y(n151) );
  INVXL U94 ( .A(A[2]), .Y(n156) );
  NAND2XL U95 ( .A(A[1]), .B(n154), .Y(n49) );
  INVXL U96 ( .A(B[1]), .Y(n154) );
  XNOR2X1 U97 ( .A(n55), .B(n4), .Y(DIFF[16]) );
  XOR2X1 U98 ( .A(B[16]), .B(A[16]), .Y(n4) );
  NAND2BXL U99 ( .AN(B[11]), .B(A[11]), .Y(n122) );
  INVX1 U100 ( .A(n13), .Y(n119) );
  OAI21XL U101 ( .A0(n28), .A1(n29), .B0(n30), .Y(n21) );
  INVX1 U102 ( .A(n31), .Y(n28) );
  NAND2BX1 U103 ( .AN(n84), .B(n76), .Y(n37) );
  XOR2X1 U104 ( .A(n21), .B(n25), .Y(DIFF[6]) );
  NOR2X1 U105 ( .A(n22), .B(n26), .Y(n25) );
  INVX1 U106 ( .A(n20), .Y(n26) );
  XOR2X1 U107 ( .A(n31), .B(n32), .Y(DIFF[5]) );
  INVX1 U108 ( .A(n34), .Y(n29) );
  INVX1 U109 ( .A(n74), .Y(n69) );
  INVX1 U110 ( .A(n86), .Y(n85) );
  NAND4X1 U111 ( .A(n38), .B(n34), .C(n20), .D(n23), .Y(n73) );
  INVX1 U112 ( .A(n8), .Y(n132) );
  INVX1 U113 ( .A(A[6]), .Y(n145) );
  OAI21XL U114 ( .A0(n149), .A1(n150), .B0(n44), .Y(n84) );
  INVX1 U115 ( .A(n43), .Y(n150) );
  OAI21XL U116 ( .A0(n48), .A1(n53), .B0(n49), .Y(n153) );
  INVX1 U117 ( .A(A[5]), .Y(n146) );
  INVX1 U118 ( .A(n148), .Y(n48) );
  NAND2X1 U119 ( .A(A[5]), .B(n142), .Y(n30) );
  XOR2X1 U120 ( .A(n13), .B(n14), .Y(DIFF[8]) );
  XOR2X1 U121 ( .A(n126), .B(n128), .Y(DIFF[10]) );
  NOR2X1 U122 ( .A(n127), .B(n129), .Y(n128) );
  INVX1 U123 ( .A(n115), .Y(n129) );
  XOR2X1 U124 ( .A(n18), .B(n19), .Y(DIFF[7]) );
  NAND2X1 U125 ( .A(n23), .B(n24), .Y(n18) );
  XOR2X1 U126 ( .A(n116), .B(n117), .Y(DIFF[12]) );
  XOR2X1 U127 ( .A(n8), .B(n9), .Y(DIFF[9]) );
  NOR2X1 U128 ( .A(n10), .B(n11), .Y(n9) );
  INVX1 U129 ( .A(n12), .Y(n10) );
  NAND2X1 U130 ( .A(n35), .B(n36), .Y(n31) );
  NAND2X1 U131 ( .A(n37), .B(n38), .Y(n35) );
  NAND3X1 U132 ( .A(n138), .B(n27), .C(n24), .Y(n137) );
  NAND3X1 U133 ( .A(n34), .B(n141), .C(n20), .Y(n138) );
  INVX1 U134 ( .A(n113), .Y(n16) );
  NAND3X1 U135 ( .A(n77), .B(n63), .C(n78), .Y(n56) );
  OAI21XL U136 ( .A0(n81), .A1(n75), .B0(n82), .Y(n77) );
  NAND2X1 U137 ( .A(A[6]), .B(n140), .Y(n27) );
  INVX1 U138 ( .A(n66), .Y(n95) );
  AND4X1 U139 ( .A(n113), .B(n13), .C(n114), .D(n115), .Y(n5) );
  INVX1 U140 ( .A(n61), .Y(n91) );
  NAND2X1 U141 ( .A(n36), .B(n30), .Y(n141) );
  INVX1 U142 ( .A(n71), .Y(n79) );
  XOR2X1 U143 ( .A(n96), .B(n97), .Y(DIFF[14]) );
  OAI21XL U144 ( .A0(n47), .A1(n48), .B0(n49), .Y(n42) );
  INVX1 U145 ( .A(n50), .Y(n47) );
  INVX1 U146 ( .A(n41), .Y(n46) );
  XOR2X1 U147 ( .A(n42), .B(n45), .Y(DIFF[2]) );
  XOR2X1 U148 ( .A(n39), .B(n40), .Y(DIFF[3]) );
  NAND2X1 U149 ( .A(n43), .B(n44), .Y(n39) );
  AOI21X1 U150 ( .A0(n41), .A1(n42), .B0(n7), .Y(n40) );
  XOR2X1 U151 ( .A(n50), .B(n51), .Y(DIFF[1]) );
  NAND2BX1 U152 ( .AN(n54), .B(n53), .Y(n50) );
  NAND2X1 U153 ( .A(n53), .B(n54), .Y(DIFF[0]) );
  INVXL U154 ( .A(B[10]), .Y(n131) );
  NAND4X1 U155 ( .A(n114), .B(n113), .C(n115), .D(n105), .Y(n75) );
  NAND3XL U156 ( .A(n123), .B(n114), .C(n115), .Y(n120) );
  NAND2X1 U157 ( .A(n12), .B(n17), .Y(n123) );
  INVX1 U158 ( .A(A[7]), .Y(n144) );
  INVX1 U159 ( .A(A[3]), .Y(n152) );
  NAND3X1 U160 ( .A(n5), .B(n105), .C(n112), .Y(n92) );
  NAND2X1 U161 ( .A(B[1]), .B(n155), .Y(n148) );
  XOR2X1 U162 ( .A(n124), .B(n125), .Y(DIFF[11]) );
  NAND2XL U163 ( .A(n105), .B(n122), .Y(n124) );
  AOI21XL U164 ( .A0(n115), .A1(n126), .B0(n127), .Y(n125) );
  NAND3X1 U165 ( .A(n5), .B(n105), .C(n111), .Y(n99) );
  NAND2X1 U166 ( .A(n104), .B(n111), .Y(n110) );
  NAND2X1 U167 ( .A(n111), .B(n104), .Y(n102) );
  NAND2X1 U168 ( .A(B[0]), .B(n158), .Y(n54) );
  INVX1 U169 ( .A(A[0]), .Y(n158) );
  NAND2X1 U170 ( .A(A[0]), .B(n159), .Y(n53) );
  INVX1 U171 ( .A(B[0]), .Y(n159) );
  NAND2BXL U172 ( .AN(A[11]), .B(B[11]), .Y(n104) );
  NAND3X1 U173 ( .A(n56), .B(n57), .C(n58), .Y(n55) );
  NAND2BXL U174 ( .AN(A[12]), .B(B[12]), .Y(n80) );
  NAND2XL U175 ( .A(A[10]), .B(n131), .Y(n121) );
  INVXL U176 ( .A(A[10]), .Y(n130) );
  NAND2X1 U177 ( .A(n63), .B(n61), .Y(n96) );
  NAND2BX1 U178 ( .AN(A[15]), .B(B[15]), .Y(n71) );
endmodule


module butterfly_DW01_sub_39 ( A, B, DIFF );
  input [16:0] A;
  input [16:0] B;
  output [16:0] DIFF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173;

  OAI21X2 U3 ( .A0(A[14]), .A1(n63), .B0(n64), .Y(n62) );
  NAND2BX1 U4 ( .AN(A[15]), .B(B[15]), .Y(n64) );
  NOR2BX2 U5 ( .AN(B[15]), .B(A[15]), .Y(n76) );
  NAND2X1 U6 ( .A(n91), .B(n127), .Y(n88) );
  OAI21X1 U7 ( .A0(n128), .A1(n129), .B0(n130), .Y(n127) );
  NAND3XL U8 ( .A(n105), .B(n109), .C(n88), .Y(n122) );
  INVX2 U9 ( .A(n109), .Y(n86) );
  NAND2X2 U10 ( .A(A[11]), .B(n139), .Y(n109) );
  INVXL U11 ( .A(n88), .Y(n87) );
  INVX1 U12 ( .A(n90), .Y(n129) );
  NAND2X1 U13 ( .A(A[10]), .B(n144), .Y(n130) );
  NOR2X2 U14 ( .A(n124), .B(n75), .Y(n123) );
  XOR2X1 U15 ( .A(n118), .B(n119), .Y(DIFF[13]) );
  INVX1 U16 ( .A(B[11]), .Y(n139) );
  OAI21XL U17 ( .A0(n151), .A1(n78), .B0(n95), .Y(n14) );
  OAI21XL U18 ( .A0(n134), .A1(n17), .B0(n132), .Y(n9) );
  OAI21XL U19 ( .A0(n114), .A1(n70), .B0(n68), .Y(n113) );
  NAND2X1 U20 ( .A(A[12]), .B(n126), .Y(n70) );
  INVX1 U21 ( .A(B[12]), .Y(n126) );
  NAND2X1 U22 ( .A(B[12]), .B(n125), .Y(n83) );
  XOR2X1 U23 ( .A(n141), .B(n142), .Y(DIFF[10]) );
  XOR2X1 U24 ( .A(n110), .B(n111), .Y(DIFF[14]) );
  NOR2X1 U25 ( .A(n107), .B(n108), .Y(n106) );
  XOR2X1 U26 ( .A(n122), .B(n123), .Y(DIFF[12]) );
  NAND2X1 U27 ( .A(n122), .B(n83), .Y(n121) );
  AOI31X1 U28 ( .A0(n105), .A1(n109), .A2(n88), .B0(n115), .Y(n112) );
  NOR2BX2 U29 ( .AN(B[13]), .B(A[13]), .Y(n114) );
  NAND2XL U30 ( .A(n54), .B(n2), .Y(n3) );
  OAI2BB1X2 U31 ( .A0N(B[13]), .A1N(n116), .B0(n83), .Y(n115) );
  NAND2BXL U32 ( .AN(A[14]), .B(B[14]), .Y(n73) );
  NOR2BX2 U33 ( .AN(B[14]), .B(A[14]), .Y(n104) );
  INVX2 U34 ( .A(n70), .Y(n124) );
  NAND2X2 U35 ( .A(n3), .B(n4), .Y(DIFF[16]) );
  NOR2X1 U36 ( .A(n112), .B(n113), .Y(n111) );
  NAND2X1 U37 ( .A(n100), .B(n67), .Y(n96) );
  NAND3X1 U38 ( .A(n101), .B(n102), .C(n103), .Y(n100) );
  NAND2BX4 U39 ( .AN(B[13]), .B(A[13]), .Y(n68) );
  NAND2X1 U40 ( .A(n1), .B(n55), .Y(n4) );
  INVX1 U41 ( .A(n54), .Y(n1) );
  INVXL U42 ( .A(n55), .Y(n2) );
  NAND2X1 U43 ( .A(n67), .B(n68), .Y(n66) );
  INVX2 U44 ( .A(n68), .Y(n107) );
  NAND2XL U45 ( .A(B[3]), .B(n168), .Y(n43) );
  NAND3BX1 U46 ( .AN(n46), .B(n163), .C(n43), .Y(n79) );
  XNOR2X1 U47 ( .A(B[16]), .B(A[16]), .Y(n55) );
  NAND2XL U48 ( .A(B[9]), .B(n148), .Y(n13) );
  NAND2XL U49 ( .A(B[6]), .B(n160), .Y(n20) );
  INVXL U50 ( .A(B[5]), .Y(n157) );
  NAND2XL U51 ( .A(B[7]), .B(n159), .Y(n23) );
  INVX2 U52 ( .A(n83), .Y(n75) );
  NOR2X1 U53 ( .A(n86), .B(n137), .Y(n136) );
  NAND4XL U54 ( .A(n133), .B(n13), .C(n90), .D(n91), .Y(n105) );
  NAND2X1 U55 ( .A(B[8]), .B(n150), .Y(n89) );
  NOR2BX1 U56 ( .AN(A[2]), .B(B[2]), .Y(n8) );
  INVXL U57 ( .A(n37), .Y(n151) );
  AOI21XL U58 ( .A0(n92), .A1(n93), .B0(n94), .Y(n84) );
  INVXL U59 ( .A(n78), .Y(n92) );
  NAND2XL U60 ( .A(n121), .B(n70), .Y(n118) );
  AOI21XL U61 ( .A0(n16), .A1(n13), .B0(n11), .Y(n128) );
  NOR2XL U62 ( .A(n134), .B(n17), .Y(n133) );
  XOR2X1 U63 ( .A(n135), .B(n136), .Y(DIFF[11]) );
  OAI21XL U64 ( .A0(n140), .A1(n129), .B0(n130), .Y(n135) );
  INVXL U65 ( .A(n132), .Y(n16) );
  NAND2X1 U66 ( .A(n23), .B(n152), .Y(n95) );
  NOR2X1 U67 ( .A(n129), .B(n143), .Y(n142) );
  INVX1 U68 ( .A(n130), .Y(n143) );
  XOR2X1 U69 ( .A(n9), .B(n10), .Y(DIFF[9]) );
  INVXL U70 ( .A(n91), .Y(n137) );
  INVXL U71 ( .A(n27), .Y(n22) );
  NOR2XL U72 ( .A(n8), .B(n46), .Y(n45) );
  AOI21XL U73 ( .A0(n20), .A1(n21), .B0(n22), .Y(n19) );
  NAND2XL U74 ( .A(n23), .B(n24), .Y(n18) );
  NOR2XL U75 ( .A(n51), .B(n7), .Y(n50) );
  INVXL U76 ( .A(n48), .Y(n51) );
  NOR2XL U77 ( .A(n33), .B(n29), .Y(n32) );
  INVXL U78 ( .A(n30), .Y(n33) );
  XNOR2X1 U79 ( .A(n37), .B(n5), .Y(DIFF[4]) );
  NAND2XL U80 ( .A(n36), .B(n38), .Y(n5) );
  NAND2XL U81 ( .A(n43), .B(n44), .Y(n39) );
  NOR2X1 U82 ( .A(n75), .B(n76), .Y(n74) );
  NAND4X1 U83 ( .A(n71), .B(n72), .C(n73), .D(n74), .Y(n57) );
  NOR3X1 U84 ( .A(n77), .B(n78), .C(n79), .Y(n72) );
  INVX1 U85 ( .A(n99), .Y(n59) );
  NAND3X1 U86 ( .A(n106), .B(n88), .C(n105), .Y(n101) );
  NAND2XL U87 ( .A(B[10]), .B(n145), .Y(n90) );
  NAND2BXL U88 ( .AN(A[13]), .B(B[13]), .Y(n71) );
  INVXL U89 ( .A(B[7]), .Y(n154) );
  INVXL U90 ( .A(B[6]), .Y(n155) );
  INVXL U91 ( .A(B[8]), .Y(n149) );
  NAND2X1 U92 ( .A(A[9]), .B(n147), .Y(n131) );
  NAND2XL U93 ( .A(B[5]), .B(n161), .Y(n34) );
  NAND2XL U94 ( .A(B[2]), .B(n171), .Y(n41) );
  INVXL U95 ( .A(B[4]), .Y(n158) );
  NAND2XL U96 ( .A(B[4]), .B(n162), .Y(n38) );
  INVXL U97 ( .A(B[1]), .Y(n170) );
  INVXL U98 ( .A(B[3]), .Y(n167) );
  INVX1 U99 ( .A(n14), .Y(n134) );
  OAI21XL U100 ( .A0(n84), .A1(n77), .B0(n85), .Y(n81) );
  NOR2X1 U101 ( .A(n86), .B(n87), .Y(n85) );
  XOR2X1 U102 ( .A(n14), .B(n15), .Y(DIFF[8]) );
  NOR2X1 U103 ( .A(n16), .B(n17), .Y(n15) );
  NAND2BX1 U104 ( .AN(n93), .B(n79), .Y(n37) );
  INVX1 U105 ( .A(n95), .Y(n94) );
  NAND4X1 U106 ( .A(n38), .B(n34), .C(n20), .D(n23), .Y(n78) );
  OAI21XL U107 ( .A0(n28), .A1(n29), .B0(n30), .Y(n21) );
  INVX1 U108 ( .A(n31), .Y(n28) );
  NOR2X1 U109 ( .A(n107), .B(n120), .Y(n119) );
  INVX1 U110 ( .A(n89), .Y(n17) );
  XOR2X1 U111 ( .A(n21), .B(n25), .Y(DIFF[6]) );
  NOR2X1 U112 ( .A(n22), .B(n26), .Y(n25) );
  INVX1 U113 ( .A(n20), .Y(n26) );
  NOR2X1 U114 ( .A(n11), .B(n12), .Y(n10) );
  INVX1 U115 ( .A(n13), .Y(n12) );
  XOR2X1 U116 ( .A(n18), .B(n19), .Y(DIFF[7]) );
  INVX1 U117 ( .A(n141), .Y(n140) );
  XOR2X1 U118 ( .A(n31), .B(n32), .Y(DIFF[5]) );
  NAND2X1 U119 ( .A(n146), .B(n131), .Y(n141) );
  NAND2X1 U120 ( .A(n9), .B(n13), .Y(n146) );
  NAND3X1 U121 ( .A(n153), .B(n27), .C(n24), .Y(n152) );
  NAND3X1 U122 ( .A(n34), .B(n156), .C(n20), .Y(n153) );
  INVX1 U123 ( .A(n34), .Y(n29) );
  INVX1 U124 ( .A(n131), .Y(n11) );
  AND2X2 U125 ( .A(n73), .B(n6), .Y(n82) );
  AND2X1 U126 ( .A(n71), .B(n83), .Y(n6) );
  NAND2X1 U127 ( .A(n36), .B(n30), .Y(n156) );
  NAND2XL U128 ( .A(n70), .B(n109), .Y(n108) );
  INVX1 U129 ( .A(n71), .Y(n120) );
  OAI21XL U130 ( .A0(n47), .A1(n7), .B0(n48), .Y(n42) );
  INVX1 U131 ( .A(n49), .Y(n47) );
  OAI21XL U132 ( .A0(n165), .A1(n166), .B0(n44), .Y(n93) );
  AOI21X1 U133 ( .A0(n41), .A1(n169), .B0(n8), .Y(n165) );
  INVX1 U134 ( .A(n43), .Y(n166) );
  OAI21XL U135 ( .A0(n7), .A1(n52), .B0(n48), .Y(n169) );
  NOR2X1 U136 ( .A(n7), .B(n164), .Y(n163) );
  INVX1 U137 ( .A(n53), .Y(n164) );
  INVX1 U138 ( .A(n41), .Y(n46) );
  XOR2X1 U139 ( .A(n42), .B(n45), .Y(DIFF[2]) );
  XOR2X1 U140 ( .A(n39), .B(n40), .Y(DIFF[3]) );
  AOI21X1 U141 ( .A0(n41), .A1(n42), .B0(n8), .Y(n40) );
  XOR2X1 U142 ( .A(n49), .B(n50), .Y(DIFF[1]) );
  NAND2X1 U143 ( .A(n35), .B(n36), .Y(n31) );
  NAND2X1 U144 ( .A(n37), .B(n38), .Y(n35) );
  NAND2BX1 U145 ( .AN(n53), .B(n52), .Y(n49) );
  NAND2X1 U146 ( .A(n52), .B(n53), .Y(DIFF[0]) );
  INVX1 U147 ( .A(A[11]), .Y(n138) );
  INVX1 U148 ( .A(A[13]), .Y(n116) );
  INVX1 U149 ( .A(A[12]), .Y(n125) );
  INVX1 U150 ( .A(A[6]), .Y(n160) );
  INVX1 U151 ( .A(A[9]), .Y(n148) );
  NAND2X1 U152 ( .A(A[5]), .B(n157), .Y(n30) );
  INVXL U153 ( .A(B[10]), .Y(n144) );
  INVX1 U154 ( .A(A[7]), .Y(n159) );
  INVX1 U155 ( .A(A[5]), .Y(n161) );
  INVXL U156 ( .A(B[9]), .Y(n147) );
  NAND2X1 U157 ( .A(A[8]), .B(n149), .Y(n132) );
  NAND2X1 U158 ( .A(A[7]), .B(n154), .Y(n24) );
  NAND2X1 U159 ( .A(A[6]), .B(n155), .Y(n27) );
  NOR2X1 U160 ( .A(n59), .B(n60), .Y(n58) );
  NOR2X1 U161 ( .A(n61), .B(n62), .Y(n60) );
  NOR2X1 U162 ( .A(n65), .B(n66), .Y(n61) );
  INVX1 U163 ( .A(A[10]), .Y(n145) );
  INVX1 U164 ( .A(A[8]), .Y(n150) );
  NAND2XL U165 ( .A(n67), .B(n117), .Y(n110) );
  NAND3X1 U166 ( .A(n56), .B(n57), .C(n58), .Y(n54) );
  NAND3X1 U167 ( .A(n80), .B(n81), .C(n82), .Y(n56) );
  NOR2X1 U168 ( .A(n69), .B(n70), .Y(n65) );
  NAND2BXL U169 ( .AN(B[15]), .B(A[15]), .Y(n99) );
  XOR2X2 U170 ( .A(n96), .B(n97), .Y(DIFF[15]) );
  NOR2X2 U171 ( .A(n59), .B(n98), .Y(n97) );
  NOR2BX1 U172 ( .AN(B[1]), .B(A[1]), .Y(n7) );
  NAND2X1 U173 ( .A(A[4]), .B(n158), .Y(n36) );
  NAND2X1 U174 ( .A(A[1]), .B(n170), .Y(n48) );
  INVX1 U175 ( .A(A[4]), .Y(n162) );
  INVX1 U176 ( .A(A[2]), .Y(n171) );
  NAND2X1 U177 ( .A(A[3]), .B(n167), .Y(n44) );
  INVX1 U178 ( .A(A[3]), .Y(n168) );
  NAND2X1 U179 ( .A(A[0]), .B(n173), .Y(n52) );
  INVX1 U180 ( .A(B[0]), .Y(n173) );
  NAND2X1 U181 ( .A(B[0]), .B(n172), .Y(n53) );
  INVX1 U182 ( .A(A[0]), .Y(n172) );
  NAND2X1 U183 ( .A(B[11]), .B(n138), .Y(n91) );
  INVXL U184 ( .A(B[14]), .Y(n63) );
  NAND4XL U185 ( .A(n13), .B(n89), .C(n90), .D(n91), .Y(n77) );
  NAND2BXL U186 ( .AN(A[14]), .B(B[14]), .Y(n117) );
  NAND2BX2 U187 ( .AN(B[14]), .B(A[14]), .Y(n67) );
  NAND2BXL U188 ( .AN(A[15]), .B(B[15]), .Y(n80) );
  NOR2BX1 U189 ( .AN(B[15]), .B(A[15]), .Y(n98) );
  NAND2BXL U190 ( .AN(A[13]), .B(B[13]), .Y(n102) );
  AOI21XL U191 ( .A0(n75), .A1(n68), .B0(n104), .Y(n103) );
  NOR2BX1 U192 ( .AN(B[13]), .B(A[13]), .Y(n69) );
endmodule


module butterfly_DW01_add_47 ( A, B, SUM );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  wire   n1, n2, n3, n4, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140;

  AND2X2 U2 ( .A(B[15]), .B(A[15]), .Y(n8) );
  XOR2X4 U3 ( .A(n89), .B(n90), .Y(SUM[15]) );
  NAND2X2 U4 ( .A(n100), .B(n2), .Y(n3) );
  NAND2X2 U5 ( .A(n1), .B(n101), .Y(n4) );
  NAND2X4 U6 ( .A(n3), .B(n4), .Y(SUM[14]) );
  CLKINVX2 U7 ( .A(n100), .Y(n1) );
  INVX1 U8 ( .A(n101), .Y(n2) );
  NAND2X1 U9 ( .A(n73), .B(n106), .Y(n100) );
  NAND2X1 U10 ( .A(B[13]), .B(A[13]), .Y(n63) );
  AOI31X2 U11 ( .A0(n96), .A1(n79), .A2(n104), .B0(n105), .Y(n102) );
  NAND2X2 U12 ( .A(n71), .B(n93), .Y(n105) );
  OAI21X2 U13 ( .A0(n59), .A1(n60), .B0(n63), .Y(n103) );
  NOR2X2 U14 ( .A(n102), .B(n103), .Y(n101) );
  NAND4X1 U15 ( .A(n118), .B(n80), .C(n82), .D(n119), .Y(n96) );
  INVX1 U16 ( .A(B[11]), .Y(n84) );
  INVX1 U17 ( .A(n71), .Y(n67) );
  XOR2X1 U18 ( .A(n122), .B(n125), .Y(SUM[10]) );
  NOR2BX1 U19 ( .AN(n124), .B(n126), .Y(n125) );
  XOR2X1 U20 ( .A(n107), .B(n108), .Y(SUM[13]) );
  NAND2X1 U21 ( .A(n110), .B(n71), .Y(n109) );
  OR2X2 U22 ( .A(B[12]), .B(A[12]), .Y(n71) );
  CLKINVX3 U23 ( .A(B[14]), .Y(n62) );
  AND2X2 U24 ( .A(n53), .B(n135), .Y(SUM[0]) );
  XOR2X1 U25 ( .A(n110), .B(n111), .Y(SUM[12]) );
  NAND2BXL U26 ( .AN(A[11]), .B(n84), .Y(n83) );
  NAND2BX1 U27 ( .AN(A[11]), .B(n84), .Y(n119) );
  AOI31XL U28 ( .A0(n96), .A1(n79), .A2(n97), .B0(n67), .Y(n94) );
  NAND3X2 U29 ( .A(n96), .B(n79), .C(n78), .Y(n110) );
  OAI21X1 U30 ( .A0(n127), .A1(n12), .B0(n11), .Y(n122) );
  CLKINVX1 U31 ( .A(n80), .Y(n12) );
  NAND2X1 U32 ( .A(n109), .B(n60), .Y(n107) );
  OAI22X2 U33 ( .A0(n91), .A1(n92), .B0(n61), .B1(n62), .Y(n89) );
  NAND2X1 U34 ( .A(n93), .B(n73), .Y(n92) );
  CLKINVX4 U35 ( .A(n93), .Y(n59) );
  XNOR2X2 U36 ( .A(n54), .B(n7), .Y(SUM[16]) );
  NOR2X2 U37 ( .A(n64), .B(n8), .Y(n90) );
  INVX2 U38 ( .A(n66), .Y(n64) );
  NAND2BX2 U39 ( .AN(n98), .B(n99), .Y(n78) );
  NAND2BX2 U40 ( .AN(A[14]), .B(n62), .Y(n73) );
  INVX1 U41 ( .A(B[10]), .Y(n113) );
  INVXL U42 ( .A(n82), .Y(n126) );
  NAND2XL U43 ( .A(n63), .B(n60), .Y(n95) );
  NOR2XL U44 ( .A(n76), .B(n77), .Y(n75) );
  NOR2BX1 U45 ( .AN(n60), .B(n67), .Y(n111) );
  INVX1 U46 ( .A(n9), .Y(n127) );
  NOR2BX1 U47 ( .AN(n34), .B(n33), .Y(n35) );
  OR2X2 U48 ( .A(B[9]), .B(A[9]), .Y(n80) );
  XNOR2X1 U49 ( .A(B[16]), .B(A[16]), .Y(n7) );
  INVXL U50 ( .A(n31), .Y(n28) );
  NOR2BXL U51 ( .AN(n30), .B(n29), .Y(n32) );
  NOR2XL U52 ( .A(n19), .B(n20), .Y(n18) );
  INVXL U53 ( .A(n25), .Y(n22) );
  INVXL U54 ( .A(n69), .Y(n85) );
  INVXL U55 ( .A(n88), .Y(n87) );
  INVXL U56 ( .A(n86), .Y(n134) );
  AOI21XL U57 ( .A0(n57), .A1(n58), .B0(n8), .Y(n56) );
  NAND2BXL U58 ( .AN(n98), .B(n99), .Y(n104) );
  NAND2XL U59 ( .A(B[6]), .B(A[6]), .Y(n24) );
  NOR2BXL U60 ( .AN(n11), .B(n12), .Y(n10) );
  INVXL U61 ( .A(n81), .Y(n16) );
  OR2XL U62 ( .A(B[6]), .B(A[6]), .Y(n27) );
  NAND2XL U63 ( .A(B[5]), .B(A[5]), .Y(n30) );
  OR2XL U64 ( .A(B[5]), .B(A[5]), .Y(n132) );
  AOI21XL U65 ( .A0(n46), .A1(n137), .B0(n138), .Y(n136) );
  NOR2BXL U66 ( .AN(n48), .B(n52), .Y(n51) );
  AOI21XL U67 ( .A0(n85), .A1(n86), .B0(n87), .Y(n74) );
  NAND2BXL U68 ( .AN(n98), .B(n99), .Y(n97) );
  XOR2X1 U69 ( .A(n120), .B(n121), .Y(SUM[11]) );
  NAND2XL U70 ( .A(n117), .B(n79), .Y(n120) );
  AOI21X1 U71 ( .A0(n82), .A1(n122), .B0(n123), .Y(n121) );
  NAND2XL U72 ( .A(B[7]), .B(A[7]), .Y(n21) );
  OR2XL U73 ( .A(B[7]), .B(A[7]), .Y(n133) );
  NAND2XL U74 ( .A(B[4]), .B(A[4]), .Y(n34) );
  OR2XL U75 ( .A(B[4]), .B(A[4]), .Y(n36) );
  NAND2XL U76 ( .A(B[1]), .B(A[1]), .Y(n48) );
  NAND2XL U77 ( .A(B[2]), .B(A[2]), .Y(n43) );
  NAND2XL U78 ( .A(B[3]), .B(A[3]), .Y(n40) );
  NOR2XL U79 ( .A(B[3]), .B(A[3]), .Y(n6) );
  OR2XL U80 ( .A(B[2]), .B(A[2]), .Y(n46) );
  OR2XL U81 ( .A(B[1]), .B(A[1]), .Y(n49) );
  NOR2BX1 U82 ( .AN(n13), .B(n16), .Y(n118) );
  OAI21XL U83 ( .A0(n134), .A1(n69), .B0(n88), .Y(n13) );
  OAI21XL U84 ( .A0(n28), .A1(n29), .B0(n30), .Y(n25) );
  INVX1 U85 ( .A(n132), .Y(n29) );
  NOR2X1 U86 ( .A(n59), .B(n65), .Y(n72) );
  XOR2X1 U87 ( .A(n31), .B(n32), .Y(SUM[5]) );
  XOR2X1 U88 ( .A(n25), .B(n26), .Y(SUM[6]) );
  NOR2BX1 U89 ( .AN(n24), .B(n23), .Y(n26) );
  XOR2X1 U90 ( .A(n17), .B(n18), .Y(SUM[7]) );
  OAI21XL U91 ( .A0(n22), .A1(n23), .B0(n24), .Y(n17) );
  INVX1 U92 ( .A(n27), .Y(n23) );
  INVX1 U93 ( .A(n78), .Y(n77) );
  NOR2X1 U94 ( .A(n94), .B(n95), .Y(n91) );
  NAND4X1 U95 ( .A(n36), .B(n132), .C(n27), .D(n133), .Y(n69) );
  NOR2XL U96 ( .A(n64), .B(n65), .Y(n57) );
  XOR2X1 U97 ( .A(n13), .B(n14), .Y(SUM[8]) );
  NOR2BX1 U98 ( .AN(n15), .B(n16), .Y(n14) );
  XOR2X1 U99 ( .A(n9), .B(n10), .Y(SUM[9]) );
  NAND2BX1 U100 ( .AN(n20), .B(n129), .Y(n88) );
  NAND3X1 U101 ( .A(n130), .B(n24), .C(n21), .Y(n129) );
  NAND2X1 U102 ( .A(n131), .B(n27), .Y(n130) );
  OAI21XL U103 ( .A0(n29), .A1(n34), .B0(n30), .Y(n131) );
  NAND2X1 U104 ( .A(n128), .B(n15), .Y(n9) );
  NAND2X1 U105 ( .A(n13), .B(n81), .Y(n128) );
  INVX1 U106 ( .A(n133), .Y(n20) );
  INVX1 U107 ( .A(n21), .Y(n19) );
  OAI21XL U108 ( .A0(n136), .A1(n6), .B0(n40), .Y(n86) );
  INVX1 U109 ( .A(n43), .Y(n138) );
  OAI21XL U110 ( .A0(n52), .A1(n53), .B0(n48), .Y(n137) );
  OAI21XL U111 ( .A0(n33), .A1(n134), .B0(n34), .Y(n31) );
  XOR2X1 U112 ( .A(n50), .B(n51), .Y(SUM[1]) );
  XOR2X1 U113 ( .A(n37), .B(n38), .Y(SUM[3]) );
  OAI21XL U114 ( .A0(n41), .A1(n42), .B0(n43), .Y(n37) );
  NOR2X1 U115 ( .A(n39), .B(n6), .Y(n38) );
  INVX1 U116 ( .A(n44), .Y(n41) );
  XOR2X1 U117 ( .A(n44), .B(n45), .Y(SUM[2]) );
  NOR2BX1 U118 ( .AN(n43), .B(n42), .Y(n45) );
  XOR2X1 U119 ( .A(n86), .B(n35), .Y(SUM[4]) );
  NAND2X1 U120 ( .A(n47), .B(n48), .Y(n44) );
  NAND2X1 U121 ( .A(n49), .B(n50), .Y(n47) );
  INVX1 U122 ( .A(n36), .Y(n33) );
  INVX1 U123 ( .A(n49), .Y(n52) );
  INVX1 U124 ( .A(n46), .Y(n42) );
  INVX1 U125 ( .A(n53), .Y(n50) );
  INVX1 U126 ( .A(n40), .Y(n39) );
  NAND2X1 U127 ( .A(n139), .B(n140), .Y(n135) );
  INVX1 U128 ( .A(B[0]), .Y(n139) );
  OAI21XL U129 ( .A0(n112), .A1(n113), .B0(n114), .Y(n99) );
  NAND3X1 U130 ( .A(n115), .B(n80), .C(n116), .Y(n114) );
  NAND2X1 U131 ( .A(n11), .B(n15), .Y(n115) );
  OR2XL U132 ( .A(B[8]), .B(A[8]), .Y(n81) );
  NAND2XL U133 ( .A(B[9]), .B(A[9]), .Y(n11) );
  NAND2XL U134 ( .A(B[8]), .B(A[8]), .Y(n15) );
  INVX1 U135 ( .A(n124), .Y(n123) );
  INVXL U136 ( .A(n79), .Y(n76) );
  OAI21XL U137 ( .A0(n74), .A1(n68), .B0(n75), .Y(n70) );
  NAND4XL U138 ( .A(n80), .B(n81), .C(n82), .D(n83), .Y(n68) );
  OR2X4 U139 ( .A(B[13]), .B(A[13]), .Y(n93) );
  OR2X2 U140 ( .A(B[15]), .B(A[15]), .Y(n66) );
  INVX1 U141 ( .A(n117), .Y(n98) );
  NAND2X1 U142 ( .A(B[0]), .B(A[0]), .Y(n53) );
  INVX1 U143 ( .A(A[0]), .Y(n140) );
  NAND2BX1 U144 ( .AN(A[11]), .B(n84), .Y(n117) );
  NAND2X1 U145 ( .A(n55), .B(n56), .Y(n54) );
  NAND4XL U146 ( .A(n70), .B(n71), .C(n66), .D(n72), .Y(n55) );
  NAND2X1 U147 ( .A(B[11]), .B(A[11]), .Y(n79) );
  NAND2X1 U148 ( .A(B[12]), .B(A[12]), .Y(n60) );
  NAND2XL U149 ( .A(B[10]), .B(A[10]), .Y(n124) );
  INVXL U150 ( .A(A[10]), .Y(n112) );
  NAND2BX1 U151 ( .AN(A[10]), .B(n113), .Y(n82) );
  NAND2BX1 U152 ( .AN(A[10]), .B(n113), .Y(n116) );
  INVX1 U153 ( .A(n73), .Y(n65) );
  NOR2BX2 U154 ( .AN(n63), .B(n59), .Y(n108) );
  OAI221XL U155 ( .A0(n59), .A1(n60), .B0(n61), .B1(n62), .C0(n63), .Y(n58) );
  INVX1 U156 ( .A(A[14]), .Y(n61) );
  NAND2XL U157 ( .A(B[14]), .B(A[14]), .Y(n106) );
endmodule


module butterfly_DW01_add_52 ( A, B, SUM );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143;

  OR2X4 U2 ( .A(A[12]), .B(B[12]), .Y(n76) );
  NAND3BXL U3 ( .AN(n9), .B(n112), .C(B[12]), .Y(n96) );
  NAND2BX1 U4 ( .AN(n10), .B(n109), .Y(n100) );
  CLKINVX2 U5 ( .A(B[13]), .Y(n109) );
  NAND3X2 U6 ( .A(n95), .B(n104), .C(n105), .Y(n101) );
  INVX1 U7 ( .A(n78), .Y(n66) );
  NAND2X1 U8 ( .A(n113), .B(n114), .Y(n110) );
  NAND2X2 U9 ( .A(n128), .B(n129), .Y(n83) );
  INVXL U10 ( .A(B[10]), .Y(n128) );
  INVXL U11 ( .A(A[10]), .Y(n129) );
  INVXL U12 ( .A(A[9]), .Y(n141) );
  INVXL U13 ( .A(B[9]), .Y(n140) );
  INVX1 U14 ( .A(n83), .Y(n120) );
  INVX4 U15 ( .A(n100), .Y(n71) );
  OAI21X1 U16 ( .A0(n65), .A1(n66), .B0(n67), .Y(n62) );
  NOR2X1 U17 ( .A(n3), .B(n68), .Y(n65) );
  NAND2BX1 U18 ( .AN(n117), .B(n108), .Y(n81) );
  NAND2X1 U19 ( .A(n118), .B(n119), .Y(n108) );
  NAND2BX1 U20 ( .AN(n120), .B(n121), .Y(n118) );
  OAI21XL U21 ( .A0(n14), .A1(n17), .B0(n13), .Y(n121) );
  NAND4X1 U22 ( .A(n122), .B(n85), .C(n83), .D(n84), .Y(n107) );
  NAND2BX1 U23 ( .AN(n10), .B(n109), .Y(n98) );
  BUFX8 U24 ( .A(A[13]), .Y(n10) );
  OAI21XL U25 ( .A0(n37), .A1(n74), .B0(n90), .Y(n15) );
  NAND2BX2 U26 ( .AN(n10), .B(n109), .Y(n112) );
  NAND2X2 U27 ( .A(n102), .B(n103), .Y(n78) );
  INVX1 U28 ( .A(B[14]), .Y(n102) );
  NAND2X1 U29 ( .A(B[13]), .B(n10), .Y(n95) );
  XOR2X1 U30 ( .A(n123), .B(n124), .Y(SUM[11]) );
  OAI21XL U31 ( .A0(n125), .A1(n120), .B0(n119), .Y(n123) );
  INVX1 U32 ( .A(n126), .Y(n125) );
  XOR2X1 U33 ( .A(n126), .B(n127), .Y(SUM[10]) );
  NOR2BX1 U34 ( .AN(n119), .B(n120), .Y(n127) );
  XNOR2X1 U35 ( .A(n58), .B(n8), .Y(SUM[16]) );
  XNOR2X4 U36 ( .A(n91), .B(n4), .Y(SUM[15]) );
  AND2X2 U37 ( .A(n57), .B(n136), .Y(SUM[0]) );
  AND2X2 U38 ( .A(B[13]), .B(n10), .Y(n3) );
  AND2X2 U39 ( .A(n61), .B(n64), .Y(n4) );
  AND2X2 U40 ( .A(n67), .B(n78), .Y(n5) );
  NAND2X1 U41 ( .A(B[14]), .B(A[14]), .Y(n67) );
  NAND2X1 U42 ( .A(B[10]), .B(A[10]), .Y(n119) );
  NAND2X1 U43 ( .A(n59), .B(n60), .Y(n58) );
  NAND4XL U44 ( .A(n75), .B(n76), .C(n61), .D(n77), .Y(n59) );
  AOI21X1 U45 ( .A0(n61), .A1(n62), .B0(n63), .Y(n60) );
  NAND2X1 U46 ( .A(B[15]), .B(A[15]), .Y(n64) );
  NAND3X1 U47 ( .A(n107), .B(n82), .C(n81), .Y(n115) );
  INVX2 U48 ( .A(n84), .Y(n117) );
  NAND3XL U49 ( .A(n112), .B(n76), .C(n99), .Y(n105) );
  INVX1 U50 ( .A(B[15]), .Y(n92) );
  NAND3XL U51 ( .A(A[12]), .B(B[12]), .C(n98), .Y(n104) );
  NAND2XL U52 ( .A(B[11]), .B(A[11]), .Y(n82) );
  OR2X2 U53 ( .A(B[11]), .B(A[11]), .Y(n84) );
  NAND2X2 U54 ( .A(n92), .B(n93), .Y(n61) );
  NAND3X1 U55 ( .A(n82), .B(n106), .C(n107), .Y(n99) );
  NAND2X1 U56 ( .A(n108), .B(n84), .Y(n106) );
  NAND3X1 U57 ( .A(n95), .B(n96), .C(n97), .Y(n94) );
  AND2X4 U58 ( .A(n6), .B(n67), .Y(n91) );
  NAND2X1 U59 ( .A(n78), .B(n94), .Y(n6) );
  NAND3XL U60 ( .A(n98), .B(n76), .C(n99), .Y(n97) );
  OAI21X2 U61 ( .A0(n14), .A1(n130), .B0(n13), .Y(n126) );
  NAND2X1 U62 ( .A(n115), .B(n76), .Y(n113) );
  INVX4 U63 ( .A(n76), .Y(n72) );
  OR2X1 U64 ( .A(B[5]), .B(A[5]), .Y(n35) );
  XOR2X2 U65 ( .A(n115), .B(n116), .Y(SUM[12]) );
  NOR2BX2 U66 ( .AN(n82), .B(n117), .Y(n124) );
  NOR2XL U67 ( .A(n21), .B(n22), .Y(n20) );
  INVXL U68 ( .A(A[15]), .Y(n93) );
  NAND2X1 U69 ( .A(B[2]), .B(A[2]), .Y(n47) );
  OR2X2 U70 ( .A(B[4]), .B(A[4]), .Y(n40) );
  OR2X2 U71 ( .A(B[1]), .B(A[1]), .Y(n53) );
  OR2X2 U72 ( .A(B[2]), .B(A[2]), .Y(n50) );
  INVXL U73 ( .A(n74), .Y(n87) );
  INVXL U74 ( .A(n90), .Y(n89) );
  AOI21XL U75 ( .A0(n87), .A1(n88), .B0(n89), .Y(n79) );
  OAI21X1 U76 ( .A0(n79), .A1(n73), .B0(n80), .Y(n75) );
  INVX4 U77 ( .A(n85), .Y(n14) );
  NAND2X1 U78 ( .A(n131), .B(n17), .Y(n11) );
  INVXL U79 ( .A(n86), .Y(n18) );
  INVXL U80 ( .A(n27), .Y(n24) );
  INVXL U81 ( .A(n135), .Y(n22) );
  INVXL U82 ( .A(n23), .Y(n21) );
  INVXL U83 ( .A(n33), .Y(n30) );
  INVXL U84 ( .A(n29), .Y(n25) );
  NOR2BXL U85 ( .AN(n47), .B(n46), .Y(n49) );
  NOR2BXL U86 ( .AN(n52), .B(n56), .Y(n55) );
  NAND2X1 U87 ( .A(B[8]), .B(A[8]), .Y(n17) );
  NAND2XL U88 ( .A(B[9]), .B(A[9]), .Y(n13) );
  NAND2XL U89 ( .A(B[6]), .B(A[6]), .Y(n26) );
  AOI21XL U90 ( .A0(n50), .A1(n138), .B0(n139), .Y(n137) );
  NAND2XL U91 ( .A(B[3]), .B(A[3]), .Y(n44) );
  NOR2XL U92 ( .A(B[3]), .B(A[3]), .Y(n7) );
  NAND2XL U93 ( .A(B[1]), .B(A[1]), .Y(n52) );
  XNOR2X1 U94 ( .A(B[16]), .B(A[16]), .Y(n8) );
  INVX1 U95 ( .A(n88), .Y(n37) );
  NOR2BX1 U96 ( .AN(n15), .B(n18), .Y(n122) );
  INVX1 U97 ( .A(n11), .Y(n130) );
  OAI21XL U98 ( .A0(n30), .A1(n31), .B0(n32), .Y(n27) );
  OAI21XL U99 ( .A0(n36), .A1(n37), .B0(n38), .Y(n33) );
  NAND4X1 U100 ( .A(n40), .B(n35), .C(n29), .D(n135), .Y(n74) );
  XOR2X1 U101 ( .A(n15), .B(n16), .Y(SUM[8]) );
  NOR2BX1 U102 ( .AN(n17), .B(n18), .Y(n16) );
  XOR2X1 U103 ( .A(n11), .B(n12), .Y(SUM[9]) );
  NOR2BXL U104 ( .AN(n13), .B(n14), .Y(n12) );
  XOR2X1 U105 ( .A(n33), .B(n34), .Y(SUM[5]) );
  NOR2BX1 U106 ( .AN(n32), .B(n31), .Y(n34) );
  XOR2X1 U107 ( .A(n27), .B(n28), .Y(SUM[6]) );
  NOR2BX1 U108 ( .AN(n26), .B(n25), .Y(n28) );
  XOR2X1 U109 ( .A(n19), .B(n20), .Y(SUM[7]) );
  OAI21XL U110 ( .A0(n24), .A1(n25), .B0(n26), .Y(n19) );
  NAND2X1 U111 ( .A(n15), .B(n86), .Y(n131) );
  NAND2BX1 U112 ( .AN(n22), .B(n132), .Y(n90) );
  NAND3X1 U113 ( .A(n133), .B(n26), .C(n23), .Y(n132) );
  NAND3X1 U114 ( .A(n35), .B(n134), .C(n29), .Y(n133) );
  NAND2X1 U115 ( .A(n38), .B(n32), .Y(n134) );
  INVX1 U116 ( .A(n35), .Y(n31) );
  INVX1 U117 ( .A(n40), .Y(n36) );
  INVX1 U118 ( .A(n53), .Y(n56) );
  AND2X1 U119 ( .A(n82), .B(n81), .Y(n80) );
  INVX1 U120 ( .A(n64), .Y(n63) );
  XOR2X1 U121 ( .A(n54), .B(n55), .Y(SUM[1]) );
  XOR2X1 U122 ( .A(n48), .B(n49), .Y(SUM[2]) );
  XOR2X1 U123 ( .A(n88), .B(n39), .Y(SUM[4]) );
  NOR2BX1 U124 ( .AN(n38), .B(n36), .Y(n39) );
  XOR2X1 U125 ( .A(n41), .B(n42), .Y(SUM[3]) );
  OAI21XL U126 ( .A0(n45), .A1(n46), .B0(n47), .Y(n41) );
  NOR2X1 U127 ( .A(n43), .B(n7), .Y(n42) );
  INVX1 U128 ( .A(n48), .Y(n45) );
  NAND2X1 U129 ( .A(n51), .B(n52), .Y(n48) );
  NAND2X1 U130 ( .A(n53), .B(n54), .Y(n51) );
  INVX1 U131 ( .A(n50), .Y(n46) );
  INVX1 U132 ( .A(n44), .Y(n43) );
  OAI21XL U133 ( .A0(n137), .A1(n7), .B0(n44), .Y(n88) );
  INVX1 U134 ( .A(n47), .Y(n139) );
  OAI21XL U135 ( .A0(n56), .A1(n57), .B0(n52), .Y(n138) );
  NAND2X1 U136 ( .A(B[4]), .B(A[4]), .Y(n38) );
  NAND2X1 U137 ( .A(B[5]), .B(A[5]), .Y(n32) );
  INVX1 U138 ( .A(A[14]), .Y(n103) );
  OR2X2 U139 ( .A(B[6]), .B(A[6]), .Y(n29) );
  OR2X2 U140 ( .A(B[7]), .B(A[7]), .Y(n135) );
  OR2X2 U141 ( .A(B[8]), .B(A[8]), .Y(n86) );
  NAND2XL U142 ( .A(B[7]), .B(A[7]), .Y(n23) );
  INVX1 U143 ( .A(n57), .Y(n54) );
  NAND2X1 U144 ( .A(n142), .B(n143), .Y(n136) );
  INVX1 U145 ( .A(B[0]), .Y(n142) );
  NAND2X1 U146 ( .A(B[0]), .B(A[0]), .Y(n57) );
  INVX1 U147 ( .A(A[0]), .Y(n143) );
  INVXL U148 ( .A(A[12]), .Y(n9) );
  NOR2X1 U149 ( .A(n69), .B(n70), .Y(n68) );
  NOR2X2 U150 ( .A(n71), .B(n66), .Y(n77) );
  NAND4XL U151 ( .A(n83), .B(n84), .C(n85), .D(n86), .Y(n73) );
  NAND2XL U152 ( .A(A[12]), .B(B[12]), .Y(n70) );
  NAND2XL U153 ( .A(B[12]), .B(A[12]), .Y(n114) );
  NOR2XL U154 ( .A(n10), .B(B[13]), .Y(n69) );
  XOR2X4 U155 ( .A(n101), .B(n5), .Y(SUM[14]) );
  XOR2X4 U156 ( .A(n110), .B(n111), .Y(SUM[13]) );
  NOR2BX4 U157 ( .AN(n95), .B(n71), .Y(n111) );
  NOR2BX4 U158 ( .AN(n114), .B(n72), .Y(n116) );
  NAND2X4 U159 ( .A(n140), .B(n141), .Y(n85) );
endmodule


module butterfly_DW01_add_50 ( A, B, SUM );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  wire   n1, n2, n3, n4, n6, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146;

  NAND2X2 U2 ( .A(n1), .B(n2), .Y(n3) );
  NAND2X2 U3 ( .A(n3), .B(n107), .Y(n103) );
  INVX1 U4 ( .A(n105), .Y(n1) );
  INVX2 U5 ( .A(n106), .Y(n2) );
  XOR2X1 U6 ( .A(n91), .B(n8), .Y(SUM[15]) );
  NOR2BX2 U7 ( .AN(n121), .B(n73), .Y(n122) );
  INVX4 U8 ( .A(B[13]), .Y(n11) );
  INVX2 U9 ( .A(B[10]), .Y(n127) );
  XOR2X2 U10 ( .A(n103), .B(n104), .Y(SUM[14]) );
  NOR3X1 U11 ( .A(n112), .B(n113), .C(n114), .Y(n105) );
  AND2X2 U12 ( .A(n63), .B(n66), .Y(n8) );
  OAI21XL U13 ( .A0(n140), .A1(n75), .B0(n90), .Y(n16) );
  NOR2X1 U14 ( .A(A[13]), .B(n10), .Y(n100) );
  OAI21XL U15 ( .A0(n97), .A1(n98), .B0(n99), .Y(n96) );
  NOR2X1 U16 ( .A(A[13]), .B(n10), .Y(n97) );
  NOR2BX1 U17 ( .AN(n124), .B(n133), .Y(n132) );
  NAND2X1 U18 ( .A(n61), .B(n62), .Y(n59) );
  XOR2X1 U19 ( .A(B[16]), .B(A[16]), .Y(n60) );
  XOR2X1 U20 ( .A(n59), .B(n60), .Y(SUM[16]) );
  OAI21X1 U21 ( .A0(n92), .A1(n68), .B0(n69), .Y(n91) );
  CLKINVX3 U22 ( .A(n93), .Y(n68) );
  AND4X2 U23 ( .A(n20), .B(n16), .C(n86), .D(n84), .Y(n4) );
  OR2X2 U24 ( .A(A[12]), .B(B[12]), .Y(n77) );
  AND2X2 U25 ( .A(n58), .B(n141), .Y(SUM[0]) );
  NOR2X1 U26 ( .A(A[13]), .B(n10), .Y(n110) );
  XOR2X2 U27 ( .A(n128), .B(n129), .Y(SUM[11]) );
  OAI21X2 U28 ( .A0(n134), .A1(n15), .B0(n14), .Y(n130) );
  CLKINVX2 U29 ( .A(n12), .Y(n134) );
  AOI21X1 U30 ( .A0(n63), .A1(n64), .B0(n65), .Y(n62) );
  OAI21XL U31 ( .A0(n67), .A1(n68), .B0(n69), .Y(n64) );
  NAND2X1 U32 ( .A(B[14]), .B(A[14]), .Y(n69) );
  INVX8 U33 ( .A(n11), .Y(n10) );
  NOR2BX2 U34 ( .AN(n108), .B(n109), .Y(n107) );
  NOR2X1 U35 ( .A(n110), .B(n98), .Y(n109) );
  OR2X2 U36 ( .A(B[11]), .B(A[11]), .Y(n85) );
  NAND2XL U37 ( .A(n14), .B(n18), .Y(n125) );
  OR2XL U38 ( .A(B[6]), .B(A[6]), .Y(n31) );
  NAND4X1 U39 ( .A(n41), .B(n37), .C(n31), .D(n139), .Y(n75) );
  INVXL U40 ( .A(n84), .Y(n133) );
  NOR2BX2 U41 ( .AN(n69), .B(n68), .Y(n104) );
  NOR2BX1 U42 ( .AN(n28), .B(n27), .Y(n30) );
  NOR2BX1 U43 ( .AN(n34), .B(n33), .Y(n36) );
  OR2X2 U44 ( .A(B[15]), .B(A[15]), .Y(n63) );
  NAND2X1 U45 ( .A(n123), .B(n124), .Y(n116) );
  NOR2XL U46 ( .A(B[3]), .B(A[3]), .Y(n6) );
  INVXL U47 ( .A(n102), .Y(n112) );
  INVXL U48 ( .A(n88), .Y(n140) );
  INVXL U49 ( .A(n90), .Y(n89) );
  INVXL U50 ( .A(n66), .Y(n65) );
  NOR2XL U51 ( .A(n9), .B(n70), .Y(n67) );
  AOI21XL U52 ( .A0(n87), .A1(n88), .B0(n89), .Y(n80) );
  AOI21X1 U53 ( .A0(n84), .A1(n130), .B0(n131), .Y(n129) );
  INVXL U54 ( .A(n124), .Y(n131) );
  NOR2BXL U55 ( .AN(n14), .B(n15), .Y(n13) );
  NOR2BXL U56 ( .AN(n79), .B(n68), .Y(n78) );
  XOR2X1 U57 ( .A(n130), .B(n132), .Y(SUM[10]) );
  NAND2X1 U58 ( .A(n4), .B(n85), .Y(n115) );
  INVXL U59 ( .A(n35), .Y(n32) );
  AOI21XL U60 ( .A0(n51), .A1(n143), .B0(n144), .Y(n142) );
  NAND2XL U61 ( .A(n54), .B(n55), .Y(n52) );
  NOR2XL U62 ( .A(n23), .B(n24), .Y(n22) );
  INVXL U63 ( .A(n29), .Y(n26) );
  NOR2BXL U64 ( .AN(n53), .B(n57), .Y(n56) );
  NOR2BXL U65 ( .AN(n39), .B(n38), .Y(n40) );
  INVXL U66 ( .A(n51), .Y(n47) );
  INVXL U67 ( .A(n25), .Y(n23) );
  OAI2BB1X1 U68 ( .A0N(n11), .A1N(n111), .B0(n77), .Y(n106) );
  NOR2XL U69 ( .A(A[13]), .B(n10), .Y(n71) );
  OR2X2 U70 ( .A(B[14]), .B(A[14]), .Y(n93) );
  NAND2XL U71 ( .A(B[11]), .B(A[11]), .Y(n82) );
  OR2X2 U72 ( .A(B[9]), .B(A[9]), .Y(n86) );
  NAND2XL U73 ( .A(B[8]), .B(A[8]), .Y(n18) );
  NAND2XL U74 ( .A(B[6]), .B(A[6]), .Y(n28) );
  OR2XL U75 ( .A(B[8]), .B(A[8]), .Y(n20) );
  OR2XL U76 ( .A(B[7]), .B(A[7]), .Y(n139) );
  NAND2XL U77 ( .A(B[4]), .B(A[4]), .Y(n39) );
  NAND2XL U78 ( .A(B[1]), .B(A[1]), .Y(n53) );
  NAND2XL U79 ( .A(B[5]), .B(A[5]), .Y(n34) );
  NAND2XL U80 ( .A(B[3]), .B(A[3]), .Y(n45) );
  OR2XL U81 ( .A(B[5]), .B(A[5]), .Y(n37) );
  INVX1 U82 ( .A(n115), .Y(n114) );
  INVX1 U83 ( .A(n75), .Y(n87) );
  INVX1 U84 ( .A(B[0]), .Y(n145) );
  OAI21XL U85 ( .A0(n142), .A1(n6), .B0(n45), .Y(n88) );
  INVX1 U86 ( .A(n48), .Y(n144) );
  OAI21XL U87 ( .A0(n57), .A1(n58), .B0(n53), .Y(n143) );
  OAI21XL U88 ( .A0(n32), .A1(n33), .B0(n34), .Y(n29) );
  OAI21XL U89 ( .A0(n38), .A1(n140), .B0(n39), .Y(n35) );
  NAND3X1 U90 ( .A(n115), .B(n82), .C(n83), .Y(n119) );
  XOR2X2 U91 ( .A(n119), .B(n122), .Y(SUM[12]) );
  INVX1 U92 ( .A(n77), .Y(n73) );
  XOR2X1 U93 ( .A(n35), .B(n36), .Y(SUM[5]) );
  XOR2X1 U94 ( .A(n16), .B(n17), .Y(SUM[8]) );
  NOR2BX1 U95 ( .AN(n18), .B(n19), .Y(n17) );
  INVX1 U96 ( .A(n20), .Y(n19) );
  NAND2X1 U97 ( .A(n85), .B(n82), .Y(n128) );
  XOR2X1 U98 ( .A(n12), .B(n13), .Y(SUM[9]) );
  XOR2X1 U99 ( .A(n29), .B(n30), .Y(SUM[6]) );
  XOR2X1 U100 ( .A(n21), .B(n22), .Y(SUM[7]) );
  OAI21XL U101 ( .A0(n26), .A1(n27), .B0(n28), .Y(n21) );
  AOI21X1 U102 ( .A0(n94), .A1(n95), .B0(n96), .Y(n92) );
  NAND3X1 U103 ( .A(n82), .B(n101), .C(n102), .Y(n94) );
  NOR2X1 U104 ( .A(n100), .B(n73), .Y(n95) );
  OAI21XL U105 ( .A0(n80), .A1(n74), .B0(n81), .Y(n76) );
  NAND4XL U106 ( .A(n84), .B(n85), .C(n86), .D(n20), .Y(n74) );
  NOR2BX1 U107 ( .AN(n82), .B(n112), .Y(n81) );
  INVX1 U108 ( .A(n86), .Y(n15) );
  NAND2BX1 U109 ( .AN(n24), .B(n136), .Y(n90) );
  NAND3X1 U110 ( .A(n137), .B(n28), .C(n25), .Y(n136) );
  NAND3X1 U111 ( .A(n37), .B(n138), .C(n31), .Y(n137) );
  NAND2X1 U112 ( .A(n39), .B(n34), .Y(n138) );
  INVX1 U113 ( .A(n31), .Y(n27) );
  INVX1 U114 ( .A(n37), .Y(n33) );
  NAND2X1 U115 ( .A(n85), .B(n116), .Y(n83) );
  NAND2X1 U116 ( .A(n85), .B(n116), .Y(n102) );
  INVX1 U117 ( .A(n41), .Y(n38) );
  INVX1 U118 ( .A(n54), .Y(n57) );
  NAND2X1 U119 ( .A(n135), .B(n18), .Y(n12) );
  NAND2X1 U120 ( .A(n16), .B(n20), .Y(n135) );
  XOR2X2 U121 ( .A(n117), .B(n118), .Y(SUM[13]) );
  NAND2X1 U122 ( .A(n108), .B(n79), .Y(n117) );
  AOI21X2 U123 ( .A0(n119), .A1(n77), .B0(n120), .Y(n118) );
  INVX1 U124 ( .A(n121), .Y(n120) );
  INVX1 U125 ( .A(n139), .Y(n24) );
  INVX1 U126 ( .A(n82), .Y(n113) );
  NAND2X1 U127 ( .A(n85), .B(n4), .Y(n101) );
  XOR2X1 U128 ( .A(n55), .B(n56), .Y(SUM[1]) );
  XOR2X1 U129 ( .A(n42), .B(n43), .Y(SUM[3]) );
  OAI21XL U130 ( .A0(n46), .A1(n47), .B0(n48), .Y(n42) );
  NOR2X1 U131 ( .A(n44), .B(n6), .Y(n43) );
  INVX1 U132 ( .A(n49), .Y(n46) );
  XOR2X1 U133 ( .A(n49), .B(n50), .Y(SUM[2]) );
  NOR2BX1 U134 ( .AN(n48), .B(n47), .Y(n50) );
  XOR2X1 U135 ( .A(n88), .B(n40), .Y(SUM[4]) );
  NAND2X1 U136 ( .A(n52), .B(n53), .Y(n49) );
  INVX1 U137 ( .A(n45), .Y(n44) );
  INVX1 U138 ( .A(n58), .Y(n55) );
  NAND2XL U139 ( .A(B[9]), .B(A[9]), .Y(n14) );
  NAND2XL U140 ( .A(B[10]), .B(A[10]), .Y(n124) );
  NAND2XL U141 ( .A(B[7]), .B(A[7]), .Y(n25) );
  NAND3X1 U142 ( .A(n125), .B(n86), .C(n126), .Y(n123) );
  NAND2BXL U143 ( .AN(A[10]), .B(n127), .Y(n126) );
  OR2X2 U144 ( .A(B[4]), .B(A[4]), .Y(n41) );
  NOR2X1 U145 ( .A(n71), .B(n72), .Y(n70) );
  NAND2BXL U146 ( .AN(A[13]), .B(n11), .Y(n79) );
  OR2X2 U147 ( .A(B[1]), .B(A[1]), .Y(n54) );
  INVX1 U148 ( .A(A[13]), .Y(n111) );
  NAND4XL U149 ( .A(n76), .B(n77), .C(n63), .D(n78), .Y(n61) );
  AND2X1 U150 ( .A(n10), .B(A[13]), .Y(n9) );
  NAND2X1 U151 ( .A(B[2]), .B(A[2]), .Y(n48) );
  OR2X2 U152 ( .A(B[2]), .B(A[2]), .Y(n51) );
  NAND2X1 U153 ( .A(B[0]), .B(A[0]), .Y(n58) );
  NAND2X1 U154 ( .A(n145), .B(n146), .Y(n141) );
  INVX1 U155 ( .A(A[0]), .Y(n146) );
  NAND2X1 U156 ( .A(B[15]), .B(A[15]), .Y(n66) );
  NAND2XL U157 ( .A(A[12]), .B(B[12]), .Y(n72) );
  NAND2XL U158 ( .A(B[12]), .B(A[12]), .Y(n121) );
  NAND2XL U159 ( .A(B[12]), .B(A[12]), .Y(n98) );
  NAND2X1 U160 ( .A(n10), .B(A[13]), .Y(n108) );
  NAND2XL U161 ( .A(n10), .B(A[13]), .Y(n99) );
  NAND2BX4 U162 ( .AN(A[10]), .B(n127), .Y(n84) );
endmodule


module butterfly_DW01_add_51 ( A, B, SUM );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  wire   n1, n2, n3, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142;

  OAI21X4 U2 ( .A0(n90), .A1(n91), .B0(n92), .Y(n89) );
  NOR2X2 U3 ( .A(n93), .B(n94), .Y(n92) );
  INVX1 U4 ( .A(n110), .Y(n1) );
  CLKINVX3 U5 ( .A(n1), .Y(n2) );
  INVX2 U6 ( .A(n83), .Y(n107) );
  XOR2X2 U7 ( .A(n109), .B(n2), .Y(SUM[13]) );
  AOI21XL U8 ( .A0(n96), .A1(n97), .B0(n111), .Y(n110) );
  NAND2X1 U9 ( .A(n130), .B(n131), .Y(n84) );
  INVX1 U10 ( .A(B[9]), .Y(n130) );
  OAI21XL U11 ( .A0(n34), .A1(n73), .B0(n88), .Y(n11) );
  INVX1 U12 ( .A(n84), .Y(n10) );
  NAND2X2 U13 ( .A(n126), .B(n127), .Y(n83) );
  NAND2BX1 U14 ( .AN(A[10]), .B(n119), .Y(n82) );
  INVX1 U15 ( .A(n136), .Y(n19) );
  INVX1 U16 ( .A(n69), .Y(n77) );
  INVX1 U17 ( .A(n96), .Y(n71) );
  NAND2BX2 U18 ( .AN(A[12]), .B(n113), .Y(n96) );
  INVX1 U19 ( .A(B[12]), .Y(n113) );
  NAND2X1 U20 ( .A(B[12]), .B(A[12]), .Y(n98) );
  NAND2X1 U21 ( .A(n114), .B(n81), .Y(n97) );
  NAND2BX1 U22 ( .AN(A[15]), .B(n70), .Y(n67) );
  OR2X2 U23 ( .A(A[14]), .B(B[14]), .Y(n69) );
  NOR2X1 U24 ( .A(n63), .B(n71), .Y(n104) );
  NAND2X1 U25 ( .A(B[13]), .B(A[13]), .Y(n95) );
  NAND2X1 U26 ( .A(n83), .B(n80), .Y(n122) );
  XOR2X1 U27 ( .A(n124), .B(n128), .Y(SUM[10]) );
  XOR2X1 U28 ( .A(n97), .B(n112), .Y(SUM[12]) );
  NOR2BX1 U29 ( .AN(n98), .B(n71), .Y(n112) );
  XOR2X1 U30 ( .A(n122), .B(n123), .Y(SUM[11]) );
  AND2X2 U31 ( .A(n62), .B(n67), .Y(n3) );
  OR2X2 U32 ( .A(A[13]), .B(B[13]), .Y(n68) );
  AND2X2 U33 ( .A(n54), .B(n137), .Y(SUM[0]) );
  NAND2XL U34 ( .A(B[14]), .B(A[14]), .Y(n66) );
  OAI21X2 U35 ( .A0(n102), .A1(n103), .B0(n104), .Y(n101) );
  NAND2X1 U36 ( .A(n108), .B(n83), .Y(n81) );
  NAND2XL U37 ( .A(n115), .B(n116), .Y(n108) );
  INVX4 U38 ( .A(B[10]), .Y(n119) );
  OAI21X1 U39 ( .A0(n129), .A1(n10), .B0(n9), .Y(n124) );
  NOR2BX2 U40 ( .AN(n80), .B(n120), .Y(n114) );
  INVXL U41 ( .A(n108), .Y(n105) );
  INVXL U42 ( .A(B[15]), .Y(n70) );
  OR2X4 U43 ( .A(B[8]), .B(A[8]), .Y(n15) );
  INVX1 U44 ( .A(n62), .Y(n61) );
  NOR2X2 U45 ( .A(n107), .B(n106), .Y(n120) );
  NAND4X1 U46 ( .A(n15), .B(n11), .C(n84), .D(n121), .Y(n106) );
  NAND2BXL U47 ( .AN(A[10]), .B(n119), .Y(n121) );
  INVXL U48 ( .A(B[11]), .Y(n126) );
  NAND3X1 U49 ( .A(n117), .B(n84), .C(n118), .Y(n115) );
  NAND2BXL U50 ( .AN(A[10]), .B(n119), .Y(n118) );
  AOI21XL U51 ( .A0(n85), .A1(n86), .B0(n87), .Y(n78) );
  INVXL U52 ( .A(n73), .Y(n85) );
  INVXL U53 ( .A(n88), .Y(n87) );
  NAND2X2 U54 ( .A(n68), .B(n95), .Y(n109) );
  NOR2BX1 U55 ( .AN(n98), .B(n97), .Y(n90) );
  NOR2BXL U56 ( .AN(n9), .B(n10), .Y(n8) );
  AND2X1 U57 ( .A(n116), .B(n82), .Y(n128) );
  INVXL U58 ( .A(n30), .Y(n27) );
  AOI21XL U59 ( .A0(n47), .A1(n139), .B0(n140), .Y(n138) );
  NOR2XL U60 ( .A(n18), .B(n19), .Y(n17) );
  INVXL U61 ( .A(n24), .Y(n21) );
  NOR2BXL U62 ( .AN(n49), .B(n53), .Y(n52) );
  INVXL U63 ( .A(n32), .Y(n28) );
  INVXL U64 ( .A(n26), .Y(n22) );
  NAND2XL U65 ( .A(B[10]), .B(A[10]), .Y(n116) );
  NAND2XL U66 ( .A(B[11]), .B(A[11]), .Y(n80) );
  NAND2XL U67 ( .A(B[6]), .B(A[6]), .Y(n23) );
  NAND2XL U68 ( .A(B[7]), .B(A[7]), .Y(n20) );
  NAND2XL U69 ( .A(B[1]), .B(A[1]), .Y(n49) );
  NAND2XL U70 ( .A(B[2]), .B(A[2]), .Y(n44) );
  NAND2XL U71 ( .A(B[3]), .B(A[3]), .Y(n41) );
  NOR2XL U72 ( .A(B[3]), .B(A[3]), .Y(n5) );
  OR2XL U73 ( .A(B[4]), .B(A[4]), .Y(n37) );
  OR2XL U74 ( .A(B[2]), .B(A[2]), .Y(n47) );
  OR2XL U75 ( .A(B[1]), .B(A[1]), .Y(n50) );
  INVX1 U76 ( .A(B[0]), .Y(n141) );
  INVX1 U77 ( .A(n86), .Y(n34) );
  INVX1 U78 ( .A(n7), .Y(n129) );
  OAI21XL U79 ( .A0(n138), .A1(n5), .B0(n41), .Y(n86) );
  INVX1 U80 ( .A(n44), .Y(n140) );
  OAI21XL U81 ( .A0(n53), .A1(n54), .B0(n49), .Y(n139) );
  OAI21XL U82 ( .A0(n27), .A1(n28), .B0(n29), .Y(n24) );
  OAI21XL U83 ( .A0(n33), .A1(n34), .B0(n35), .Y(n30) );
  NAND4X1 U84 ( .A(n37), .B(n32), .C(n26), .D(n136), .Y(n73) );
  INVXL U85 ( .A(n98), .Y(n111) );
  NAND4XL U86 ( .A(n82), .B(n83), .C(n84), .D(n15), .Y(n72) );
  AOI21X1 U87 ( .A0(n105), .A1(n106), .B0(n107), .Y(n102) );
  XOR2X1 U88 ( .A(n11), .B(n12), .Y(SUM[8]) );
  NOR2BX1 U89 ( .AN(n13), .B(n14), .Y(n12) );
  INVX1 U90 ( .A(n15), .Y(n14) );
  AOI21X1 U91 ( .A0(n82), .A1(n124), .B0(n125), .Y(n123) );
  INVX1 U92 ( .A(n116), .Y(n125) );
  XOR2X1 U93 ( .A(n7), .B(n8), .Y(SUM[9]) );
  XOR2X1 U94 ( .A(n30), .B(n31), .Y(SUM[5]) );
  NOR2BX1 U95 ( .AN(n29), .B(n28), .Y(n31) );
  XOR2X1 U96 ( .A(n24), .B(n25), .Y(SUM[6]) );
  NOR2BX1 U97 ( .AN(n23), .B(n22), .Y(n25) );
  XOR2X1 U98 ( .A(n16), .B(n17), .Y(SUM[7]) );
  OAI21XL U99 ( .A0(n21), .A1(n22), .B0(n23), .Y(n16) );
  XNOR2X4 U100 ( .A(n99), .B(n100), .Y(SUM[14]) );
  NAND2X1 U101 ( .A(n132), .B(n13), .Y(n7) );
  NAND2X1 U102 ( .A(n11), .B(n15), .Y(n132) );
  NAND2BX1 U103 ( .AN(n19), .B(n133), .Y(n88) );
  NAND3X1 U104 ( .A(n134), .B(n23), .C(n20), .Y(n133) );
  NAND3X1 U105 ( .A(n32), .B(n135), .C(n26), .Y(n134) );
  NAND2X1 U106 ( .A(n29), .B(n35), .Y(n135) );
  NAND3X1 U107 ( .A(n68), .B(n69), .C(n96), .Y(n91) );
  INVX1 U108 ( .A(n37), .Y(n33) );
  INVX1 U109 ( .A(n50), .Y(n53) );
  NAND2XL U110 ( .A(n98), .B(n80), .Y(n103) );
  AND2X1 U111 ( .A(n80), .B(n81), .Y(n79) );
  INVXL U112 ( .A(n66), .Y(n94) );
  NOR2XL U113 ( .A(n77), .B(n95), .Y(n93) );
  INVX1 U114 ( .A(n20), .Y(n18) );
  XOR2X1 U115 ( .A(n51), .B(n52), .Y(SUM[1]) );
  XOR2X1 U116 ( .A(n45), .B(n46), .Y(SUM[2]) );
  NOR2BX1 U117 ( .AN(n44), .B(n43), .Y(n46) );
  XOR2X1 U118 ( .A(n86), .B(n36), .Y(SUM[4]) );
  NOR2BX1 U119 ( .AN(n35), .B(n33), .Y(n36) );
  XOR2X1 U120 ( .A(n38), .B(n39), .Y(SUM[3]) );
  OAI21XL U121 ( .A0(n42), .A1(n43), .B0(n44), .Y(n38) );
  NOR2X1 U122 ( .A(n40), .B(n5), .Y(n39) );
  INVX1 U123 ( .A(n45), .Y(n42) );
  NAND2X1 U124 ( .A(n48), .B(n49), .Y(n45) );
  NAND2X1 U125 ( .A(n50), .B(n51), .Y(n48) );
  INVX1 U126 ( .A(n47), .Y(n43) );
  INVX1 U127 ( .A(n41), .Y(n40) );
  INVX1 U128 ( .A(n54), .Y(n51) );
  OAI21XL U129 ( .A0(n78), .A1(n72), .B0(n79), .Y(n75) );
  OAI211XL U130 ( .A0(n63), .A1(n64), .B0(n65), .C0(n66), .Y(n60) );
  INVX1 U131 ( .A(A[11]), .Y(n127) );
  INVX1 U132 ( .A(A[9]), .Y(n131) );
  NAND2XL U133 ( .A(B[9]), .B(A[9]), .Y(n9) );
  NAND2X1 U134 ( .A(B[5]), .B(A[5]), .Y(n29) );
  NAND2X1 U135 ( .A(B[8]), .B(A[8]), .Y(n13) );
  OR2X2 U136 ( .A(B[6]), .B(A[6]), .Y(n26) );
  NAND2XL U137 ( .A(n9), .B(n13), .Y(n117) );
  OR2X2 U138 ( .A(B[5]), .B(A[5]), .Y(n32) );
  OR2X2 U139 ( .A(B[7]), .B(A[7]), .Y(n136) );
  AND2X2 U140 ( .A(n67), .B(n6), .Y(n59) );
  OR2XL U141 ( .A(A[14]), .B(B[14]), .Y(n6) );
  NAND2X2 U142 ( .A(n57), .B(n58), .Y(n55) );
  NAND2X1 U143 ( .A(B[4]), .B(A[4]), .Y(n35) );
  NAND2X1 U144 ( .A(B[0]), .B(A[0]), .Y(n54) );
  NAND2X1 U145 ( .A(n141), .B(n142), .Y(n137) );
  INVX1 U146 ( .A(A[0]), .Y(n142) );
  AOI21X2 U147 ( .A0(n59), .A1(n60), .B0(n61), .Y(n58) );
  XOR2X2 U148 ( .A(n55), .B(n56), .Y(SUM[16]) );
  NAND3BX1 U149 ( .AN(n74), .B(n75), .C(n76), .Y(n57) );
  NOR3XL U150 ( .A(n77), .B(n71), .C(n63), .Y(n76) );
  NAND2XL U151 ( .A(A[12]), .B(B[12]), .Y(n64) );
  NOR2XL U152 ( .A(A[15]), .B(B[15]), .Y(n74) );
  NAND2X1 U153 ( .A(B[15]), .B(A[15]), .Y(n62) );
  NAND2XL U154 ( .A(B[13]), .B(A[13]), .Y(n65) );
  NOR2XL U155 ( .A(A[13]), .B(B[13]), .Y(n63) );
  XOR2X4 U156 ( .A(B[16]), .B(A[16]), .Y(n56) );
  XOR2X4 U157 ( .A(n89), .B(n3), .Y(SUM[15]) );
  NAND2X4 U158 ( .A(n66), .B(n69), .Y(n100) );
  NAND2X4 U159 ( .A(n101), .B(n95), .Y(n99) );
endmodule


module butterfly_DW01_add_68 ( A, B, SUM );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154;

  NAND2X2 U2 ( .A(n129), .B(n130), .Y(n101) );
  NOR2X2 U3 ( .A(n64), .B(n65), .Y(n63) );
  NAND2X2 U4 ( .A(n74), .B(n67), .Y(n90) );
  NAND2BX2 U5 ( .AN(n104), .B(n83), .Y(n124) );
  NAND3X1 U6 ( .A(n80), .B(n123), .C(n124), .Y(n120) );
  NAND2X1 U7 ( .A(n70), .B(n71), .Y(n69) );
  NAND2BX4 U8 ( .AN(A[10]), .B(n128), .Y(n82) );
  INVX3 U9 ( .A(B[10]), .Y(n128) );
  CLKINVX3 U10 ( .A(n80), .Y(n113) );
  CLKINVX2 U11 ( .A(n83), .Y(n103) );
  NAND2X2 U12 ( .A(n8), .B(n2), .Y(n3) );
  NAND2X2 U13 ( .A(n1), .B(n125), .Y(n4) );
  NAND2X4 U14 ( .A(n3), .B(n4), .Y(SUM[12]) );
  INVX2 U15 ( .A(n8), .Y(n1) );
  INVX4 U16 ( .A(n125), .Y(n2) );
  NAND2X2 U17 ( .A(n122), .B(n89), .Y(n8) );
  CLKINVX4 U18 ( .A(B[13]), .Y(n99) );
  NAND2BX2 U19 ( .AN(A[10]), .B(n128), .Y(n127) );
  INVX1 U20 ( .A(n95), .Y(n6) );
  NAND2X2 U21 ( .A(n16), .B(n19), .Y(n141) );
  OR2X2 U22 ( .A(n23), .B(n9), .Y(n87) );
  OR2X2 U23 ( .A(B[8]), .B(A[8]), .Y(n19) );
  CLKINVX3 U24 ( .A(B[11]), .Y(n137) );
  OAI21X2 U25 ( .A0(n140), .A1(n15), .B0(n14), .Y(n135) );
  INVX2 U26 ( .A(n12), .Y(n140) );
  NAND2X1 U27 ( .A(n83), .B(n101), .Y(n123) );
  XOR2X1 U28 ( .A(n20), .B(n21), .Y(SUM[7]) );
  OAI21X1 U29 ( .A0(n36), .A1(n88), .B0(n87), .Y(n16) );
  NAND2X1 U30 ( .A(B[8]), .B(A[8]), .Y(n18) );
  CLKINVX3 U31 ( .A(n84), .Y(n15) );
  NAND2X1 U32 ( .A(B[9]), .B(A[9]), .Y(n14) );
  INVX1 U33 ( .A(n145), .Y(n26) );
  NAND2X1 U34 ( .A(B[10]), .B(A[10]), .Y(n130) );
  INVX1 U35 ( .A(n144), .Y(n31) );
  NAND4X1 U36 ( .A(n19), .B(n16), .C(n84), .D(n127), .Y(n104) );
  NAND2X2 U37 ( .A(n7), .B(n96), .Y(n92) );
  NAND2X1 U38 ( .A(n5), .B(n6), .Y(n7) );
  NAND2BX2 U39 ( .AN(n11), .B(n77), .Y(n60) );
  OAI21XL U40 ( .A0(n78), .A1(n76), .B0(n79), .Y(n77) );
  NAND2X2 U41 ( .A(B[13]), .B(A[13]), .Y(n71) );
  AOI21X2 U42 ( .A0(n82), .A1(n135), .B0(n136), .Y(n134) );
  OAI21X1 U43 ( .A0(n103), .A1(n104), .B0(n112), .Y(n110) );
  INVX1 U44 ( .A(n130), .Y(n136) );
  NOR2X2 U45 ( .A(n62), .B(n63), .Y(n61) );
  AND2X4 U46 ( .A(n130), .B(n82), .Y(n139) );
  NAND4X1 U47 ( .A(n89), .B(n73), .C(n67), .D(n66), .Y(n11) );
  AND2X2 U48 ( .A(n18), .B(n19), .Y(n17) );
  NOR2X2 U49 ( .A(n98), .B(n72), .Y(n97) );
  CLKINVX4 U50 ( .A(A[11]), .Y(n138) );
  XOR2X4 U51 ( .A(n133), .B(n134), .Y(SUM[11]) );
  OAI21X2 U52 ( .A0(n98), .A1(n72), .B0(n71), .Y(n111) );
  CLKINVX2 U53 ( .A(n89), .Y(n114) );
  NAND2X2 U54 ( .A(n83), .B(n80), .Y(n133) );
  NAND2X1 U55 ( .A(n66), .B(n67), .Y(n65) );
  CLKINVX3 U56 ( .A(A[13]), .Y(n100) );
  NOR2BX4 U57 ( .AN(n14), .B(n15), .Y(n13) );
  NOR2X2 U58 ( .A(A[13]), .B(B[13]), .Y(n98) );
  INVX1 U59 ( .A(n94), .Y(n5) );
  OAI2BB1X2 U60 ( .A0N(n99), .A1N(n100), .B0(n89), .Y(n95) );
  NOR2BX2 U61 ( .AN(n71), .B(n97), .Y(n96) );
  INVX2 U62 ( .A(n124), .Y(n126) );
  INVX2 U63 ( .A(n123), .Y(n81) );
  NAND2X2 U64 ( .A(B[12]), .B(A[12]), .Y(n72) );
  AOI21X2 U65 ( .A0(n120), .A1(n89), .B0(n121), .Y(n118) );
  NAND2X4 U66 ( .A(n71), .B(n73), .Y(n119) );
  INVXL U67 ( .A(n72), .Y(n121) );
  NAND3X1 U68 ( .A(n131), .B(n84), .C(n132), .Y(n129) );
  NAND2XL U69 ( .A(B[7]), .B(A[7]), .Y(n24) );
  AOI21X2 U70 ( .A0(n99), .A1(n100), .B0(n114), .Y(n109) );
  NOR2X1 U71 ( .A(n68), .B(n69), .Y(n64) );
  XOR2X1 U72 ( .A(n33), .B(n34), .Y(SUM[5]) );
  INVXL U73 ( .A(A[0]), .Y(n154) );
  INVX4 U74 ( .A(B[14]), .Y(n115) );
  INVX4 U75 ( .A(A[14]), .Y(n116) );
  INVXL U76 ( .A(n88), .Y(n75) );
  NOR2BXL U77 ( .AN(n52), .B(n56), .Y(n55) );
  NAND2XL U78 ( .A(n53), .B(n54), .Y(n51) );
  AOI21XL U79 ( .A0(n75), .A1(n85), .B0(n86), .Y(n78) );
  NOR2BX1 U80 ( .AN(n80), .B(n81), .Y(n79) );
  AND3X2 U81 ( .A(n142), .B(n27), .C(n24), .Y(n9) );
  INVXL U82 ( .A(n33), .Y(n30) );
  NOR2XL U83 ( .A(n42), .B(n43), .Y(n41) );
  NAND2XL U84 ( .A(B[1]), .B(A[1]), .Y(n52) );
  INVXL U85 ( .A(n50), .Y(n46) );
  AND2X1 U86 ( .A(n57), .B(n148), .Y(SUM[0]) );
  NAND2XL U87 ( .A(B[0]), .B(A[0]), .Y(n57) );
  INVXL U88 ( .A(B[0]), .Y(n153) );
  OR2X4 U89 ( .A(A[12]), .B(B[12]), .Y(n89) );
  NAND2XL U90 ( .A(B[12]), .B(A[12]), .Y(n122) );
  OR2X4 U91 ( .A(B[9]), .B(A[9]), .Y(n84) );
  OR2X2 U92 ( .A(B[7]), .B(A[7]), .Y(n146) );
  NAND2XL U93 ( .A(B[5]), .B(A[5]), .Y(n32) );
  NAND2BX1 U94 ( .AN(B[3]), .B(n150), .Y(n147) );
  NAND2XL U95 ( .A(B[4]), .B(A[4]), .Y(n37) );
  NAND2XL U96 ( .A(B[3]), .B(A[3]), .Y(n44) );
  INVX1 U97 ( .A(n85), .Y(n36) );
  XOR2X1 U98 ( .A(n54), .B(n55), .Y(SUM[1]) );
  INVX1 U99 ( .A(n53), .Y(n56) );
  NAND2X1 U100 ( .A(n51), .B(n52), .Y(n48) );
  INVX1 U101 ( .A(n57), .Y(n54) );
  INVX1 U102 ( .A(n87), .Y(n86) );
  XOR2X1 U103 ( .A(n28), .B(n29), .Y(SUM[6]) );
  NOR2BX1 U104 ( .AN(n27), .B(n26), .Y(n29) );
  NOR2BX1 U105 ( .AN(n32), .B(n31), .Y(n34) );
  OAI21XL U106 ( .A0(n25), .A1(n26), .B0(n27), .Y(n20) );
  NOR2X1 U107 ( .A(n22), .B(n23), .Y(n21) );
  INVX1 U108 ( .A(n28), .Y(n25) );
  XOR2X1 U109 ( .A(n40), .B(n41), .Y(SUM[3]) );
  OAI21XL U110 ( .A0(n45), .A1(n46), .B0(n47), .Y(n40) );
  INVX1 U111 ( .A(n48), .Y(n45) );
  XOR2X1 U112 ( .A(n85), .B(n38), .Y(SUM[4]) );
  NOR2BX1 U113 ( .AN(n37), .B(n35), .Y(n38) );
  INVX2 U114 ( .A(n70), .Y(n93) );
  OAI21XL U115 ( .A0(n149), .A1(n43), .B0(n44), .Y(n85) );
  AOI21X1 U116 ( .A0(n50), .A1(n151), .B0(n152), .Y(n149) );
  INVX1 U117 ( .A(n47), .Y(n152) );
  OAI21XL U118 ( .A0(n56), .A1(n57), .B0(n52), .Y(n151) );
  OAI21XL U119 ( .A0(n30), .A1(n31), .B0(n32), .Y(n28) );
  OAI21XL U120 ( .A0(n35), .A1(n36), .B0(n37), .Y(n33) );
  NAND4X1 U121 ( .A(n39), .B(n144), .C(n145), .D(n146), .Y(n88) );
  NAND2BX1 U122 ( .AN(n26), .B(n143), .Y(n142) );
  OAI21XL U123 ( .A0(n31), .A1(n37), .B0(n32), .Y(n143) );
  INVX1 U124 ( .A(n39), .Y(n35) );
  OR2X2 U125 ( .A(B[1]), .B(A[1]), .Y(n53) );
  NOR2BX1 U126 ( .AN(n73), .B(n72), .Y(n68) );
  OAI21XL U127 ( .A0(n103), .A1(n104), .B0(n80), .Y(n102) );
  INVX1 U128 ( .A(n146), .Y(n23) );
  INVX1 U129 ( .A(n44), .Y(n42) );
  INVX1 U130 ( .A(n24), .Y(n22) );
  XOR2X1 U131 ( .A(n48), .B(n49), .Y(SUM[2]) );
  NOR2BX1 U132 ( .AN(n47), .B(n46), .Y(n49) );
  NAND2X1 U133 ( .A(n153), .B(n154), .Y(n148) );
  NAND2X1 U134 ( .A(B[2]), .B(A[2]), .Y(n47) );
  NAND2X1 U135 ( .A(B[6]), .B(A[6]), .Y(n27) );
  OR2X2 U136 ( .A(B[6]), .B(A[6]), .Y(n145) );
  OR2X2 U137 ( .A(B[5]), .B(A[5]), .Y(n144) );
  OR2X2 U138 ( .A(B[4]), .B(A[4]), .Y(n39) );
  OR2X2 U139 ( .A(B[2]), .B(A[2]), .Y(n50) );
  INVX1 U140 ( .A(n147), .Y(n43) );
  INVX1 U141 ( .A(A[3]), .Y(n150) );
  NAND2XL U142 ( .A(n14), .B(n18), .Y(n131) );
  NAND2BXL U143 ( .AN(A[10]), .B(n128), .Y(n132) );
  NAND2X4 U144 ( .A(n60), .B(n61), .Y(n58) );
  XNOR2X4 U145 ( .A(n118), .B(n119), .Y(n117) );
  INVX8 U146 ( .A(n117), .Y(SUM[13]) );
  INVXL U147 ( .A(n74), .Y(n62) );
  NAND2X1 U148 ( .A(B[15]), .B(A[15]), .Y(n74) );
  NAND2X2 U149 ( .A(B[14]), .B(A[14]), .Y(n70) );
  INVX4 U150 ( .A(B[15]), .Y(n105) );
  INVX4 U151 ( .A(A[15]), .Y(n106) );
  NAND4XL U152 ( .A(n82), .B(n83), .C(n84), .D(n19), .Y(n76) );
  AOI21XL U153 ( .A0(n83), .A1(n101), .B0(n102), .Y(n94) );
  AOI21XL U154 ( .A0(n83), .A1(n101), .B0(n113), .Y(n112) );
  XOR2X4 U155 ( .A(n12), .B(n13), .Y(SUM[9]) );
  XOR2X4 U156 ( .A(n16), .B(n17), .Y(SUM[8]) );
  XOR2X4 U157 ( .A(n58), .B(n59), .Y(SUM[16]) );
  XOR2X4 U158 ( .A(B[16]), .B(A[16]), .Y(n59) );
  XOR2X4 U159 ( .A(n90), .B(n91), .Y(SUM[15]) );
  AOI21X4 U160 ( .A0(n92), .A1(n66), .B0(n93), .Y(n91) );
  NAND2X4 U161 ( .A(n105), .B(n106), .Y(n67) );
  XOR2X4 U162 ( .A(n107), .B(n108), .Y(SUM[14]) );
  AOI21X4 U163 ( .A0(n109), .A1(n110), .B0(n111), .Y(n108) );
  NAND2X4 U164 ( .A(n66), .B(n70), .Y(n107) );
  NAND2X4 U165 ( .A(n115), .B(n116), .Y(n66) );
  NAND2BX4 U166 ( .AN(A[13]), .B(n99), .Y(n73) );
  NOR3X4 U167 ( .A(n81), .B(n113), .C(n126), .Y(n125) );
  NAND2X4 U168 ( .A(B[11]), .B(A[11]), .Y(n80) );
  NAND2X4 U169 ( .A(n137), .B(n138), .Y(n83) );
  XOR2X4 U170 ( .A(n135), .B(n139), .Y(SUM[10]) );
  NAND2X4 U171 ( .A(n141), .B(n18), .Y(n12) );
endmodule


module butterfly_DW01_sub_42 ( A, B, DIFF );
  input [16:0] A;
  input [16:0] B;
  output [16:0] DIFF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157;

  NOR2X2 U3 ( .A(n75), .B(n76), .Y(n73) );
  AOI21X1 U4 ( .A0(B[15]), .A1(n68), .B0(n69), .Y(n67) );
  NAND2BX4 U5 ( .AN(A[14]), .B(B[14]), .Y(n65) );
  NAND2X1 U6 ( .A(B[9]), .B(n130), .Y(n116) );
  NAND2XL U7 ( .A(A[10]), .B(n127), .Y(n115) );
  NAND2X1 U8 ( .A(B[10]), .B(n126), .Y(n118) );
  NAND2X1 U9 ( .A(A[11]), .B(n123), .Y(n112) );
  INVX1 U10 ( .A(B[11]), .Y(n123) );
  AND2X2 U11 ( .A(n82), .B(n81), .Y(n80) );
  OAI21XL U12 ( .A0(n9), .A1(n15), .B0(n112), .Y(n109) );
  NAND2BX1 U13 ( .AN(A[13]), .B(B[13]), .Y(n63) );
  NAND2BX2 U14 ( .AN(A[12]), .B(B[12]), .Y(n64) );
  NAND2BX2 U15 ( .AN(B[14]), .B(A[14]), .Y(n82) );
  INVX1 U16 ( .A(A[15]), .Y(n68) );
  NAND2X1 U17 ( .A(B[11]), .B(n124), .Y(n114) );
  NAND2BX2 U18 ( .AN(B[13]), .B(A[13]), .Y(n81) );
  AOI21XL U19 ( .A0(n111), .A1(n112), .B0(n113), .Y(n110) );
  AOI21X1 U20 ( .A0(n92), .A1(n64), .B0(n93), .Y(n89) );
  NAND2XL U21 ( .A(n56), .B(B[15]), .Y(n55) );
  NOR2BXL U22 ( .AN(B[15]), .B(A[15]), .Y(n87) );
  NAND2BXL U23 ( .AN(B[15]), .B(A[15]), .Y(n88) );
  NAND3BX1 U24 ( .AN(n66), .B(n67), .C(n65), .Y(n52) );
  INVX2 U25 ( .A(n88), .Y(n74) );
  NOR2X2 U26 ( .A(n74), .B(n87), .Y(n86) );
  NAND3X2 U27 ( .A(n1), .B(n54), .C(n55), .Y(n53) );
  AOI21X2 U28 ( .A0(n72), .A1(n73), .B0(n74), .Y(n51) );
  OAI21X2 U29 ( .A0(n78), .A1(n79), .B0(n80), .Y(n72) );
  NOR2BX2 U30 ( .AN(B[15]), .B(A[15]), .Y(n76) );
  OAI21X1 U31 ( .A0(n89), .A1(n90), .B0(n82), .Y(n85) );
  XOR2X2 U32 ( .A(n85), .B(n86), .Y(DIFF[15]) );
  XOR2X4 U33 ( .A(B[16]), .B(A[16]), .Y(n3) );
  XNOR2X4 U34 ( .A(n50), .B(n3), .Y(DIFF[16]) );
  NAND3X2 U35 ( .A(n51), .B(n52), .C(n53), .Y(n50) );
  XOR2X1 U36 ( .A(n102), .B(n103), .Y(DIFF[13]) );
  AND3X2 U37 ( .A(n63), .B(n64), .C(n65), .Y(n1) );
  INVXL U38 ( .A(n118), .Y(n111) );
  INVX1 U39 ( .A(n116), .Y(n9) );
  INVX1 U40 ( .A(n20), .Y(n136) );
  NOR2XL U41 ( .A(n8), .B(n9), .Y(n7) );
  NAND2XL U42 ( .A(A[12]), .B(n83), .Y(n79) );
  CLKINVX3 U43 ( .A(n107), .Y(n99) );
  INVX1 U44 ( .A(A[6]), .Y(n143) );
  INVXL U45 ( .A(B[12]), .Y(n83) );
  NOR2XL U46 ( .A(n122), .B(n111), .Y(n125) );
  INVXL U47 ( .A(n61), .Y(n134) );
  AOI21X1 U48 ( .A0(n97), .A1(n92), .B0(n98), .Y(n96) );
  INVX2 U49 ( .A(n64), .Y(n69) );
  OAI21X1 U50 ( .A0(n108), .A1(n109), .B0(n110), .Y(n59) );
  NAND4BBX1 U51 ( .AN(n58), .BN(n71), .C(n70), .D(n63), .Y(n66) );
  NAND4X1 U52 ( .A(n116), .B(n117), .C(n114), .D(n118), .Y(n58) );
  AOI21XL U53 ( .A0(n92), .A1(n64), .B0(n99), .Y(n103) );
  INVXL U54 ( .A(n114), .Y(n113) );
  INVXL U55 ( .A(n6), .Y(n128) );
  INVXL U56 ( .A(n10), .Y(n8) );
  INVXL U57 ( .A(n11), .Y(n131) );
  AOI21XL U58 ( .A0(n18), .A1(n138), .B0(n4), .Y(n135) );
  NOR2XL U59 ( .A(n13), .B(n14), .Y(n12) );
  INVXL U60 ( .A(n15), .Y(n14) );
  AOI21XL U61 ( .A0(n70), .A1(n60), .B0(n61), .Y(n57) );
  NOR2XL U62 ( .A(n4), .B(n23), .Y(n22) );
  INVXL U63 ( .A(n18), .Y(n23) );
  XNOR2X1 U64 ( .A(n32), .B(n2), .Y(DIFF[4]) );
  NAND2XL U65 ( .A(n33), .B(n31), .Y(n2) );
  NAND2XL U66 ( .A(n20), .B(n21), .Y(n16) );
  AOI21XL U67 ( .A0(n18), .A1(n19), .B0(n4), .Y(n17) );
  NOR2XL U68 ( .A(n29), .B(n25), .Y(n28) );
  INVXL U69 ( .A(n26), .Y(n29) );
  NAND2XL U70 ( .A(n30), .B(n31), .Y(n27) );
  NAND2XL U71 ( .A(n32), .B(n33), .Y(n30) );
  NAND2XL U72 ( .A(n38), .B(n39), .Y(n34) );
  NAND2BX2 U73 ( .AN(B[12]), .B(A[12]), .Y(n107) );
  INVX2 U74 ( .A(A[11]), .Y(n124) );
  NOR2X1 U75 ( .A(A[14]), .B(n77), .Y(n75) );
  INVXL U76 ( .A(B[14]), .Y(n77) );
  NOR2XL U77 ( .A(A[13]), .B(n84), .Y(n78) );
  INVX1 U78 ( .A(B[10]), .Y(n127) );
  NAND2XL U79 ( .A(B[8]), .B(n155), .Y(n117) );
  INVXL U80 ( .A(A[8]), .Y(n155) );
  INVXL U81 ( .A(B[9]), .Y(n129) );
  INVXL U82 ( .A(B[5]), .Y(n139) );
  INVXL U83 ( .A(B[7]), .Y(n137) );
  NAND4XL U84 ( .A(n38), .B(n36), .C(n49), .D(n146), .Y(n71) );
  NAND2XL U85 ( .A(B[4]), .B(n145), .Y(n33) );
  INVXL U86 ( .A(A[4]), .Y(n145) );
  INVXL U87 ( .A(B[3]), .Y(n149) );
  OAI21XL U88 ( .A0(n133), .A1(n62), .B0(n134), .Y(n11) );
  INVX1 U89 ( .A(n32), .Y(n133) );
  NAND2X1 U90 ( .A(n104), .B(n59), .Y(n92) );
  NAND2BX1 U91 ( .AN(n58), .B(n11), .Y(n104) );
  XOR2X1 U92 ( .A(n121), .B(n125), .Y(DIFF[10]) );
  NAND4X1 U93 ( .A(n33), .B(n141), .C(n18), .D(n20), .Y(n62) );
  NAND2X1 U94 ( .A(n10), .B(n115), .Y(n108) );
  OAI21XL U95 ( .A0(n128), .A1(n9), .B0(n10), .Y(n121) );
  OAI21XL U96 ( .A0(n13), .A1(n131), .B0(n15), .Y(n6) );
  OAI21XL U97 ( .A0(n135), .A1(n136), .B0(n21), .Y(n61) );
  OAI21XL U98 ( .A0(n25), .A1(n31), .B0(n26), .Y(n138) );
  INVX1 U99 ( .A(n141), .Y(n25) );
  XOR2X1 U100 ( .A(n105), .B(n106), .Y(DIFF[12]) );
  NAND2XL U101 ( .A(n104), .B(n59), .Y(n105) );
  NOR2X1 U102 ( .A(n69), .B(n99), .Y(n106) );
  OAI21XL U103 ( .A0(n57), .A1(n58), .B0(n59), .Y(n54) );
  INVX1 U104 ( .A(n62), .Y(n70) );
  INVX1 U105 ( .A(n117), .Y(n13) );
  INVXL U106 ( .A(n115), .Y(n122) );
  XOR2X1 U107 ( .A(n95), .B(n96), .Y(DIFF[14]) );
  NOR2XL U108 ( .A(n69), .B(n101), .Y(n97) );
  XOR2X1 U109 ( .A(n11), .B(n12), .Y(DIFF[8]) );
  XOR2X1 U110 ( .A(n119), .B(n120), .Y(DIFF[11]) );
  NAND2XL U111 ( .A(n114), .B(n112), .Y(n119) );
  AOI21XL U112 ( .A0(n118), .A1(n121), .B0(n122), .Y(n120) );
  XOR2X1 U113 ( .A(n6), .B(n7), .Y(DIFF[9]) );
  INVX1 U114 ( .A(n91), .Y(n101) );
  OAI21XL U115 ( .A0(n24), .A1(n25), .B0(n26), .Y(n19) );
  INVX1 U116 ( .A(n27), .Y(n24) );
  NAND2BX1 U117 ( .AN(n60), .B(n71), .Y(n32) );
  INVX1 U118 ( .A(n146), .Y(n43) );
  INVX1 U119 ( .A(n36), .Y(n41) );
  XOR2X1 U120 ( .A(n19), .B(n22), .Y(DIFF[6]) );
  XOR2X1 U121 ( .A(n16), .B(n17), .Y(DIFF[7]) );
  XOR2X1 U122 ( .A(n27), .B(n28), .Y(DIFF[5]) );
  OAI21XL U123 ( .A0(n42), .A1(n43), .B0(n44), .Y(n37) );
  INVX1 U124 ( .A(n45), .Y(n42) );
  XOR2X1 U125 ( .A(n37), .B(n40), .Y(DIFF[2]) );
  NOR2X1 U126 ( .A(n5), .B(n41), .Y(n40) );
  XOR2X1 U127 ( .A(n34), .B(n35), .Y(DIFF[3]) );
  AOI21X1 U128 ( .A0(n36), .A1(n37), .B0(n5), .Y(n35) );
  XOR2X1 U129 ( .A(n45), .B(n46), .Y(DIFF[1]) );
  NOR2X1 U130 ( .A(n47), .B(n43), .Y(n46) );
  INVX1 U131 ( .A(n44), .Y(n47) );
  NAND2X1 U132 ( .A(B[6]), .B(n143), .Y(n18) );
  INVX1 U133 ( .A(A[10]), .Y(n126) );
  NAND2X1 U134 ( .A(B[7]), .B(n142), .Y(n20) );
  INVX1 U135 ( .A(A[7]), .Y(n142) );
  NAND2X1 U136 ( .A(A[9]), .B(n129), .Y(n10) );
  NOR2BX1 U137 ( .AN(A[6]), .B(B[6]), .Y(n4) );
  INVXL U138 ( .A(B[13]), .Y(n84) );
  NAND2X1 U139 ( .A(A[7]), .B(n137), .Y(n21) );
  NAND2X1 U140 ( .A(B[5]), .B(n144), .Y(n141) );
  INVX1 U141 ( .A(A[5]), .Y(n144) );
  INVX1 U142 ( .A(A[9]), .Y(n130) );
  NAND2BXL U143 ( .AN(A[13]), .B(B[13]), .Y(n91) );
  NAND2X1 U144 ( .A(n99), .B(n100), .Y(n94) );
  NAND2BXL U145 ( .AN(A[13]), .B(B[13]), .Y(n100) );
  INVX1 U146 ( .A(A[15]), .Y(n56) );
  NAND2X1 U147 ( .A(A[8]), .B(n132), .Y(n15) );
  INVX1 U148 ( .A(B[8]), .Y(n132) );
  OAI21XL U149 ( .A0(n147), .A1(n148), .B0(n39), .Y(n60) );
  INVX1 U150 ( .A(n38), .Y(n148) );
  AOI21X1 U151 ( .A0(n36), .A1(n151), .B0(n5), .Y(n147) );
  OAI21XL U152 ( .A0(n43), .A1(n48), .B0(n44), .Y(n151) );
  NAND2X1 U153 ( .A(A[4]), .B(n140), .Y(n31) );
  INVX1 U154 ( .A(B[4]), .Y(n140) );
  NAND2X1 U155 ( .A(B[2]), .B(n154), .Y(n36) );
  INVX1 U156 ( .A(A[2]), .Y(n154) );
  NAND2X1 U157 ( .A(B[3]), .B(n150), .Y(n38) );
  INVX1 U158 ( .A(A[3]), .Y(n150) );
  NAND2X1 U159 ( .A(A[1]), .B(n152), .Y(n44) );
  INVX1 U160 ( .A(B[1]), .Y(n152) );
  NAND2X1 U161 ( .A(A[5]), .B(n139), .Y(n26) );
  NOR2BX1 U162 ( .AN(A[2]), .B(B[2]), .Y(n5) );
  NAND2X1 U163 ( .A(B[1]), .B(n153), .Y(n146) );
  INVX1 U164 ( .A(A[1]), .Y(n153) );
  NAND2X1 U165 ( .A(A[3]), .B(n149), .Y(n39) );
  NAND2X1 U166 ( .A(n48), .B(n49), .Y(DIFF[0]) );
  NAND2BX1 U167 ( .AN(n49), .B(n48), .Y(n45) );
  NAND2X1 U168 ( .A(A[0]), .B(n157), .Y(n48) );
  INVX1 U169 ( .A(B[0]), .Y(n157) );
  NAND2X1 U170 ( .A(B[0]), .B(n156), .Y(n49) );
  INVX1 U171 ( .A(A[0]), .Y(n156) );
  NAND2XL U172 ( .A(n91), .B(n65), .Y(n90) );
  NAND2XL U173 ( .A(n82), .B(n65), .Y(n95) );
  NAND2XL U174 ( .A(n63), .B(n81), .Y(n102) );
  NAND2XL U175 ( .A(n94), .B(n81), .Y(n98) );
  NAND2XL U176 ( .A(n94), .B(n81), .Y(n93) );
endmodule


module butterfly_DW01_add_72 ( A, B, SUM );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132;

  NAND2X2 U2 ( .A(n51), .B(n52), .Y(n50) );
  NAND3BX2 U3 ( .AN(n53), .B(n54), .C(n55), .Y(n52) );
  AOI21X2 U4 ( .A0(n74), .A1(n75), .B0(n76), .Y(n51) );
  NAND2X2 U5 ( .A(n113), .B(n114), .Y(n71) );
  XOR2X2 U6 ( .A(n91), .B(n92), .Y(SUM[14]) );
  NOR2X2 U7 ( .A(n56), .B(n57), .Y(n55) );
  OAI21X1 U8 ( .A0(B[14]), .A1(A[14]), .B0(n60), .Y(n79) );
  NAND2X2 U9 ( .A(n58), .B(n59), .Y(n57) );
  INVX1 U10 ( .A(B[11]), .Y(n113) );
  NAND2BX1 U11 ( .AN(A[15]), .B(n90), .Y(n74) );
  NAND2X1 U12 ( .A(B[12]), .B(A[12]), .Y(n81) );
  AND2X2 U13 ( .A(n49), .B(n126), .Y(SUM[0]) );
  NAND2X1 U14 ( .A(n96), .B(n58), .Y(n87) );
  NAND2X1 U15 ( .A(n60), .B(n59), .Y(n88) );
  NAND2XL U16 ( .A(B[14]), .B(A[14]), .Y(n80) );
  NAND2XL U17 ( .A(n94), .B(n89), .Y(n91) );
  OAI21X1 U18 ( .A0(n78), .A1(n79), .B0(n80), .Y(n75) );
  OR2X4 U19 ( .A(A[14]), .B(B[14]), .Y(n59) );
  XOR2X2 U20 ( .A(n82), .B(n83), .Y(SUM[15]) );
  NOR2X2 U21 ( .A(n84), .B(n85), .Y(n83) );
  NAND3XL U22 ( .A(n103), .B(n70), .C(n71), .Y(n65) );
  NAND2XL U23 ( .A(B[6]), .B(A[6]), .Y(n20) );
  NAND2X1 U24 ( .A(n11), .B(n7), .Y(n106) );
  NAND2X1 U25 ( .A(n104), .B(n105), .Y(n103) );
  NAND4XL U26 ( .A(n107), .B(n72), .C(n70), .D(n71), .Y(n102) );
  AOI21X1 U27 ( .A0(n86), .A1(n87), .B0(n88), .Y(n85) );
  AND2X1 U28 ( .A(n65), .B(n64), .Y(n63) );
  NOR2BXL U29 ( .AN(n44), .B(n48), .Y(n47) );
  NAND2XL U30 ( .A(n45), .B(n46), .Y(n43) );
  NAND2XL U31 ( .A(B[9]), .B(A[9]), .Y(n7) );
  NAND2XL U32 ( .A(B[1]), .B(A[1]), .Y(n44) );
  INVXL U33 ( .A(n68), .Y(n119) );
  AOI21XL U34 ( .A0(n66), .A1(n67), .B0(n68), .Y(n61) );
  INVXL U35 ( .A(n67), .Y(n125) );
  NAND2XL U36 ( .A(n60), .B(n89), .Y(n97) );
  NAND3X1 U37 ( .A(n102), .B(n64), .C(n65), .Y(n96) );
  INVXL U38 ( .A(n60), .Y(n56) );
  NAND2XL U39 ( .A(n95), .B(n60), .Y(n94) );
  NAND2XL U40 ( .A(n87), .B(n81), .Y(n95) );
  INVXL U41 ( .A(n105), .Y(n112) );
  NOR2BXL U42 ( .AN(n7), .B(n8), .Y(n6) );
  NAND4XL U43 ( .A(n32), .B(n124), .C(n23), .D(n121), .Y(n69) );
  NAND2XL U44 ( .A(n118), .B(n11), .Y(n5) );
  NAND2XL U45 ( .A(n9), .B(n73), .Y(n118) );
  NOR2BXL U46 ( .AN(n26), .B(n25), .Y(n28) );
  NOR2XL U47 ( .A(n15), .B(n16), .Y(n14) );
  INVXL U48 ( .A(n21), .Y(n18) );
  INVXL U49 ( .A(n23), .Y(n19) );
  INVXL U50 ( .A(n42), .Y(n38) );
  NAND2XL U51 ( .A(B[13]), .B(A[13]), .Y(n89) );
  INVXL U52 ( .A(B[15]), .Y(n90) );
  NAND2XL U53 ( .A(B[15]), .B(A[15]), .Y(n77) );
  OR2X2 U54 ( .A(B[10]), .B(A[10]), .Y(n70) );
  OR2X2 U55 ( .A(B[9]), .B(A[9]), .Y(n72) );
  NAND2XL U56 ( .A(B[5]), .B(A[5]), .Y(n26) );
  NAND2XL U57 ( .A(B[7]), .B(A[7]), .Y(n17) );
  NAND2XL U58 ( .A(B[3]), .B(A[3]), .Y(n36) );
  NOR2BXL U59 ( .AN(n128), .B(A[3]), .Y(n2) );
  OR2XL U60 ( .A(B[4]), .B(A[4]), .Y(n32) );
  XOR2X2 U61 ( .A(n50), .B(n4), .Y(SUM[16]) );
  XOR2X2 U62 ( .A(B[16]), .B(A[16]), .Y(n4) );
  OAI21XL U63 ( .A0(n125), .A1(n69), .B0(n119), .Y(n9) );
  XOR2X1 U64 ( .A(n96), .B(n100), .Y(SUM[12]) );
  NOR2BX1 U65 ( .AN(n81), .B(n101), .Y(n100) );
  INVX1 U66 ( .A(n58), .Y(n101) );
  INVX1 U67 ( .A(n69), .Y(n66) );
  NOR2X1 U68 ( .A(n108), .B(n12), .Y(n107) );
  INVX1 U69 ( .A(n9), .Y(n108) );
  OAI21XL U70 ( .A0(n117), .A1(n8), .B0(n7), .Y(n111) );
  INVX1 U71 ( .A(n5), .Y(n117) );
  NAND2X1 U72 ( .A(n106), .B(n72), .Y(n104) );
  OR2X2 U73 ( .A(B[12]), .B(A[12]), .Y(n58) );
  OAI21XL U74 ( .A0(n120), .A1(n16), .B0(n17), .Y(n68) );
  AOI21X1 U75 ( .A0(n23), .A1(n122), .B0(n123), .Y(n120) );
  INVX1 U76 ( .A(n20), .Y(n123) );
  OAI21XL U77 ( .A0(n25), .A1(n30), .B0(n26), .Y(n122) );
  INVX1 U78 ( .A(n124), .Y(n25) );
  NAND4XL U79 ( .A(n70), .B(n71), .C(n72), .D(n73), .Y(n62) );
  AND2X1 U80 ( .A(n89), .B(n81), .Y(n86) );
  INVX1 U81 ( .A(n72), .Y(n8) );
  INVX1 U82 ( .A(n73), .Y(n12) );
  INVX1 U83 ( .A(n121), .Y(n16) );
  XOR2X1 U84 ( .A(n9), .B(n10), .Y(SUM[8]) );
  NOR2BX1 U85 ( .AN(n11), .B(n12), .Y(n10) );
  XOR2X1 U86 ( .A(n111), .B(n115), .Y(SUM[10]) );
  NOR2BX1 U87 ( .AN(n105), .B(n116), .Y(n115) );
  INVX1 U88 ( .A(n70), .Y(n116) );
  XOR2X1 U89 ( .A(n97), .B(n98), .Y(SUM[13]) );
  AOI21XL U90 ( .A0(n96), .A1(n58), .B0(n99), .Y(n98) );
  INVXL U91 ( .A(n81), .Y(n99) );
  XOR2X1 U92 ( .A(n109), .B(n110), .Y(SUM[11]) );
  AOI21X1 U93 ( .A0(n70), .A1(n111), .B0(n112), .Y(n110) );
  NAND2XL U94 ( .A(n71), .B(n64), .Y(n109) );
  NAND2X1 U95 ( .A(n77), .B(n74), .Y(n82) );
  INVX1 U96 ( .A(n80), .Y(n84) );
  NOR2BX1 U97 ( .AN(n80), .B(n93), .Y(n92) );
  INVX1 U98 ( .A(n59), .Y(n93) );
  XOR2X1 U99 ( .A(n5), .B(n6), .Y(SUM[9]) );
  OAI21XL U100 ( .A0(n127), .A1(n2), .B0(n36), .Y(n67) );
  AOI21X1 U101 ( .A0(n42), .A1(n129), .B0(n130), .Y(n127) );
  INVX1 U102 ( .A(n39), .Y(n130) );
  OAI21XL U103 ( .A0(n48), .A1(n49), .B0(n44), .Y(n129) );
  OAI21XL U104 ( .A0(n24), .A1(n25), .B0(n26), .Y(n21) );
  INVX1 U105 ( .A(n27), .Y(n24) );
  OAI21XL U106 ( .A0(n29), .A1(n125), .B0(n30), .Y(n27) );
  INVX1 U107 ( .A(n45), .Y(n48) );
  XOR2X1 U108 ( .A(n21), .B(n22), .Y(SUM[6]) );
  NOR2BX1 U109 ( .AN(n20), .B(n19), .Y(n22) );
  XOR2X1 U110 ( .A(n13), .B(n14), .Y(SUM[7]) );
  OAI21XL U111 ( .A0(n18), .A1(n19), .B0(n20), .Y(n13) );
  INVX1 U112 ( .A(n17), .Y(n15) );
  INVX1 U113 ( .A(n32), .Y(n29) );
  XOR2X1 U114 ( .A(n27), .B(n28), .Y(SUM[5]) );
  XOR2X1 U115 ( .A(n67), .B(n31), .Y(SUM[4]) );
  NOR2BX1 U116 ( .AN(n30), .B(n29), .Y(n31) );
  XOR2X1 U117 ( .A(n46), .B(n47), .Y(SUM[1]) );
  XOR2X1 U118 ( .A(n40), .B(n41), .Y(SUM[2]) );
  NOR2BX1 U119 ( .AN(n39), .B(n38), .Y(n41) );
  XOR2X1 U120 ( .A(n33), .B(n34), .Y(SUM[3]) );
  OAI21XL U121 ( .A0(n37), .A1(n38), .B0(n39), .Y(n33) );
  NOR2X1 U122 ( .A(n35), .B(n2), .Y(n34) );
  INVX1 U123 ( .A(n40), .Y(n37) );
  NAND2X1 U124 ( .A(n43), .B(n44), .Y(n40) );
  INVX1 U125 ( .A(n36), .Y(n35) );
  INVX1 U126 ( .A(n49), .Y(n46) );
  NAND2X1 U127 ( .A(n131), .B(n132), .Y(n126) );
  INVX1 U128 ( .A(B[0]), .Y(n131) );
  OR2X4 U129 ( .A(A[13]), .B(B[13]), .Y(n60) );
  INVX1 U130 ( .A(A[11]), .Y(n114) );
  INVX1 U131 ( .A(n77), .Y(n76) );
  AOI21XL U132 ( .A0(B[13]), .A1(A[13]), .B0(n99), .Y(n78) );
  NAND2X1 U133 ( .A(B[11]), .B(A[11]), .Y(n64) );
  OR2X2 U134 ( .A(B[6]), .B(A[6]), .Y(n23) );
  OR2X2 U135 ( .A(B[8]), .B(A[8]), .Y(n73) );
  OAI21XL U136 ( .A0(n61), .A1(n62), .B0(n63), .Y(n54) );
  NAND2X1 U137 ( .A(B[8]), .B(A[8]), .Y(n11) );
  NAND2X1 U138 ( .A(B[10]), .B(A[10]), .Y(n105) );
  OR2X2 U139 ( .A(B[7]), .B(A[7]), .Y(n121) );
  OR2X2 U140 ( .A(B[5]), .B(A[5]), .Y(n124) );
  NAND2X1 U141 ( .A(B[4]), .B(A[4]), .Y(n30) );
  NAND2X1 U142 ( .A(B[2]), .B(A[2]), .Y(n39) );
  OR2X2 U143 ( .A(B[2]), .B(A[2]), .Y(n42) );
  OR2X2 U144 ( .A(B[1]), .B(A[1]), .Y(n45) );
  INVX1 U145 ( .A(B[3]), .Y(n128) );
  NAND2X1 U146 ( .A(B[0]), .B(A[0]), .Y(n49) );
  INVX1 U147 ( .A(A[0]), .Y(n132) );
  NOR2XL U148 ( .A(A[15]), .B(B[15]), .Y(n53) );
endmodule


module butterfly_DW01_sub_57 ( A, B, DIFF );
  input [16:0] A;
  input [16:0] B;
  output [16:0] DIFF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172;

  NOR2X1 U3 ( .A(n13), .B(n63), .Y(n62) );
  AOI21X2 U4 ( .A0(n64), .A1(n65), .B0(n66), .Y(n63) );
  OAI21X1 U5 ( .A0(n101), .A1(n102), .B0(n103), .Y(n100) );
  NOR2BX2 U6 ( .AN(B[13]), .B(A[13]), .Y(n116) );
  NAND4X1 U7 ( .A(n90), .B(n21), .C(n20), .D(n132), .Y(n107) );
  NAND2XL U8 ( .A(n78), .B(n83), .Y(n1) );
  NAND3XL U9 ( .A(n2), .B(n84), .C(n68), .Y(n60) );
  INVX1 U10 ( .A(n1), .Y(n2) );
  NOR2BXL U11 ( .AN(n79), .B(n77), .Y(n84) );
  NAND3XL U12 ( .A(n73), .B(n68), .C(n74), .Y(n3) );
  NAND2X1 U13 ( .A(n4), .B(n75), .Y(n61) );
  INVX1 U14 ( .A(n3), .Y(n4) );
  NOR2XL U15 ( .A(n76), .B(n77), .Y(n75) );
  NOR2BX1 U16 ( .AN(B[13]), .B(A[13]), .Y(n104) );
  NOR2BX2 U17 ( .AN(B[13]), .B(A[13]), .Y(n119) );
  INVX2 U18 ( .A(A[15]), .Y(n99) );
  NAND2BXL U19 ( .AN(A[13]), .B(B[13]), .Y(n70) );
  INVX1 U20 ( .A(n65), .Y(n5) );
  NAND2BX1 U21 ( .AN(B[14]), .B(A[14]), .Y(n65) );
  INVXL U22 ( .A(B[12]), .Y(n125) );
  OAI21XL U23 ( .A0(n127), .A1(n128), .B0(n129), .Y(n111) );
  NAND2X1 U24 ( .A(B[11]), .B(n136), .Y(n92) );
  NAND2X1 U25 ( .A(n111), .B(n92), .Y(n89) );
  OAI21XL U26 ( .A0(n148), .A1(n81), .B0(n149), .Y(n21) );
  INVX1 U27 ( .A(n78), .Y(n118) );
  INVX1 U28 ( .A(n116), .Y(n8) );
  XOR2X1 U29 ( .A(n58), .B(n59), .Y(DIFF[16]) );
  NAND2BX1 U30 ( .AN(A[14]), .B(n7), .Y(n105) );
  INVX2 U31 ( .A(n106), .Y(n69) );
  INVX1 U32 ( .A(n5), .Y(n6) );
  BUFX3 U33 ( .A(B[14]), .Y(n7) );
  NAND2X2 U34 ( .A(n100), .B(n6), .Y(n96) );
  NAND2BX2 U35 ( .AN(B[13]), .B(A[13]), .Y(n72) );
  NAND2BXL U36 ( .AN(A[14]), .B(n7), .Y(n120) );
  OAI2BB1X2 U37 ( .A0N(n7), .A1N(n67), .B0(n68), .Y(n66) );
  AOI21X1 U38 ( .A0(n69), .A1(n70), .B0(n71), .Y(n64) );
  INVX2 U39 ( .A(n105), .Y(n77) );
  NOR2X2 U40 ( .A(n77), .B(n104), .Y(n103) );
  NAND2X2 U41 ( .A(n8), .B(n69), .Y(n9) );
  NAND2X2 U42 ( .A(n9), .B(n72), .Y(n115) );
  NAND2X1 U43 ( .A(A[12]), .B(n125), .Y(n106) );
  AOI21X4 U44 ( .A0(n113), .A1(n114), .B0(n115), .Y(n112) );
  INVXL U45 ( .A(n129), .Y(n142) );
  XNOR2X2 U46 ( .A(n11), .B(n112), .Y(DIFF[14]) );
  INVXL U47 ( .A(n92), .Y(n135) );
  INVXL U48 ( .A(A[6]), .Y(n158) );
  INVXL U49 ( .A(A[5]), .Y(n159) );
  NAND2XL U50 ( .A(A[4]), .B(n155), .Y(n40) );
  INVXL U51 ( .A(B[4]), .Y(n155) );
  NOR2X1 U52 ( .A(n18), .B(n19), .Y(n17) );
  NOR2X1 U53 ( .A(n139), .B(n142), .Y(n141) );
  NAND2X1 U54 ( .A(n41), .B(n42), .Y(n39) );
  INVXL U55 ( .A(n35), .Y(n38) );
  NAND3XL U56 ( .A(n117), .B(n108), .C(n89), .Y(n114) );
  NAND2X1 U57 ( .A(B[8]), .B(n170), .Y(n90) );
  INVXL U58 ( .A(n95), .Y(n149) );
  NOR2XL U59 ( .A(n23), .B(n24), .Y(n22) );
  NOR2XL U60 ( .A(n81), .B(n82), .Y(n73) );
  INVXL U61 ( .A(n80), .Y(n74) );
  XOR2X1 U62 ( .A(n96), .B(n97), .Y(DIFF[15]) );
  XOR2X1 U63 ( .A(n123), .B(n124), .Y(DIFF[12]) );
  NAND2XL U64 ( .A(n78), .B(n79), .Y(n76) );
  AOI21XL U65 ( .A0(n93), .A1(n94), .B0(n95), .Y(n85) );
  NOR2XL U66 ( .A(n87), .B(n88), .Y(n86) );
  INVXL U67 ( .A(n81), .Y(n93) );
  INVXL U68 ( .A(n20), .Y(n19) );
  NAND2XL U69 ( .A(n16), .B(n20), .Y(n143) );
  NOR2XL U70 ( .A(n12), .B(n32), .Y(n31) );
  INVXL U71 ( .A(n27), .Y(n32) );
  AOI21XL U72 ( .A0(n27), .A1(n28), .B0(n12), .Y(n26) );
  NAND2XL U73 ( .A(n29), .B(n30), .Y(n25) );
  NOR2XL U74 ( .A(n38), .B(n34), .Y(n37) );
  NAND3BXL U75 ( .AN(n50), .B(n161), .C(n47), .Y(n82) );
  NOR2XL U76 ( .A(n15), .B(n50), .Y(n49) );
  INVXL U77 ( .A(n45), .Y(n50) );
  NAND2XL U78 ( .A(n47), .B(n48), .Y(n43) );
  AOI21XL U79 ( .A0(n45), .A1(n46), .B0(n15), .Y(n44) );
  XNOR2X1 U80 ( .A(n41), .B(n10), .Y(DIFF[4]) );
  NAND2XL U81 ( .A(n42), .B(n40), .Y(n10) );
  NOR2BXL U82 ( .AN(B[10]), .B(A[10]), .Y(n128) );
  INVXL U83 ( .A(n111), .Y(n109) );
  NAND2XL U84 ( .A(n78), .B(n92), .Y(n110) );
  NAND2BXL U85 ( .AN(A[13]), .B(B[13]), .Y(n79) );
  NAND3X1 U86 ( .A(n117), .B(n108), .C(n89), .Y(n123) );
  NAND2BX1 U87 ( .AN(n107), .B(n92), .Y(n117) );
  AND2X2 U88 ( .A(n65), .B(n120), .Y(n11) );
  NAND2XL U89 ( .A(A[9]), .B(n144), .Y(n130) );
  INVXL U90 ( .A(B[8]), .Y(n147) );
  INVXL U91 ( .A(A[3]), .Y(n166) );
  INVXL U92 ( .A(A[4]), .Y(n160) );
  NAND2XL U93 ( .A(A[5]), .B(n154), .Y(n35) );
  INVXL U94 ( .A(B[5]), .Y(n154) );
  NOR2BXL U95 ( .AN(B[1]), .B(A[1]), .Y(n14) );
  INVXL U96 ( .A(A[2]), .Y(n169) );
  NAND2XL U97 ( .A(A[1]), .B(n168), .Y(n52) );
  INVXL U98 ( .A(B[1]), .Y(n168) );
  NAND2XL U99 ( .A(A[3]), .B(n165), .Y(n48) );
  INVXL U100 ( .A(B[3]), .Y(n165) );
  NAND2XL U101 ( .A(A[11]), .B(n137), .Y(n108) );
  INVX1 U102 ( .A(n41), .Y(n148) );
  XOR2X1 U103 ( .A(n21), .B(n22), .Y(DIFF[8]) );
  NAND2BX1 U104 ( .AN(n94), .B(n82), .Y(n41) );
  NAND4X1 U105 ( .A(n42), .B(n156), .C(n27), .D(n29), .Y(n81) );
  OAI21XL U106 ( .A0(n33), .A1(n34), .B0(n35), .Y(n28) );
  INVX1 U107 ( .A(n36), .Y(n33) );
  OAI21XL U108 ( .A0(n23), .A1(n146), .B0(n131), .Y(n16) );
  INVX1 U109 ( .A(n21), .Y(n146) );
  OAI21XL U110 ( .A0(n150), .A1(n151), .B0(n30), .Y(n95) );
  AOI21X1 U111 ( .A0(n27), .A1(n153), .B0(n12), .Y(n150) );
  INVX1 U112 ( .A(n29), .Y(n151) );
  OAI21XL U113 ( .A0(n34), .A1(n40), .B0(n35), .Y(n153) );
  XOR2X1 U114 ( .A(n121), .B(n122), .Y(DIFF[13]) );
  AOI21X1 U115 ( .A0(n123), .A1(n78), .B0(n69), .Y(n122) );
  NAND2X1 U116 ( .A(n79), .B(n72), .Y(n121) );
  INVX1 U117 ( .A(n156), .Y(n34) );
  XOR2X1 U118 ( .A(n133), .B(n134), .Y(DIFF[11]) );
  OAI21XL U119 ( .A0(n138), .A1(n139), .B0(n129), .Y(n133) );
  NOR2X1 U120 ( .A(n87), .B(n135), .Y(n134) );
  INVX1 U121 ( .A(n140), .Y(n138) );
  NOR2X1 U122 ( .A(n98), .B(n13), .Y(n97) );
  XOR2X1 U123 ( .A(n28), .B(n31), .Y(DIFF[6]) );
  XOR2X1 U124 ( .A(n16), .B(n17), .Y(DIFF[9]) );
  XOR2X1 U125 ( .A(n25), .B(n26), .Y(DIFF[7]) );
  NOR2X1 U126 ( .A(n118), .B(n69), .Y(n124) );
  XOR2X1 U127 ( .A(n140), .B(n141), .Y(DIFF[10]) );
  XOR2X1 U128 ( .A(n36), .B(n37), .Y(DIFF[5]) );
  INVX1 U129 ( .A(n90), .Y(n23) );
  NAND2X1 U130 ( .A(n143), .B(n130), .Y(n140) );
  INVX1 U131 ( .A(n91), .Y(n139) );
  INVXL U132 ( .A(n68), .Y(n98) );
  OAI21XL U133 ( .A0(n85), .A1(n80), .B0(n86), .Y(n83) );
  INVX1 U134 ( .A(n131), .Y(n24) );
  INVX1 U135 ( .A(n130), .Y(n18) );
  INVX1 U136 ( .A(n89), .Y(n88) );
  OAI21XL U137 ( .A0(n51), .A1(n14), .B0(n52), .Y(n46) );
  INVX1 U138 ( .A(n53), .Y(n51) );
  OAI21XL U139 ( .A0(n163), .A1(n164), .B0(n48), .Y(n94) );
  AOI21X1 U140 ( .A0(n45), .A1(n167), .B0(n15), .Y(n163) );
  INVX1 U141 ( .A(n47), .Y(n164) );
  OAI21XL U142 ( .A0(n14), .A1(n56), .B0(n52), .Y(n167) );
  NOR2X1 U143 ( .A(n14), .B(n162), .Y(n161) );
  INVX1 U144 ( .A(n57), .Y(n162) );
  XOR2X1 U145 ( .A(n46), .B(n49), .Y(DIFF[2]) );
  XOR2X1 U146 ( .A(n43), .B(n44), .Y(DIFF[3]) );
  XOR2X1 U147 ( .A(n53), .B(n54), .Y(DIFF[1]) );
  NOR2X1 U148 ( .A(n55), .B(n14), .Y(n54) );
  INVX1 U149 ( .A(n52), .Y(n55) );
  NAND2X1 U150 ( .A(n39), .B(n40), .Y(n36) );
  NAND2BX1 U151 ( .AN(n57), .B(n56), .Y(n53) );
  NAND2X1 U152 ( .A(n56), .B(n57), .Y(DIFF[0]) );
  NAND2X1 U153 ( .A(B[9]), .B(n145), .Y(n20) );
  INVXL U154 ( .A(A[9]), .Y(n145) );
  AOI31X1 U155 ( .A0(n107), .A1(n108), .A2(n109), .B0(n110), .Y(n101) );
  NAND2X2 U156 ( .A(B[12]), .B(n126), .Y(n78) );
  INVXL U157 ( .A(A[12]), .Y(n126) );
  NAND2X1 U158 ( .A(B[6]), .B(n158), .Y(n27) );
  AOI21X1 U159 ( .A0(n24), .A1(n20), .B0(n18), .Y(n127) );
  NAND4XL U160 ( .A(n20), .B(n90), .C(n91), .D(n92), .Y(n80) );
  INVX1 U161 ( .A(A[8]), .Y(n170) );
  NAND2X1 U162 ( .A(B[7]), .B(n157), .Y(n29) );
  INVX1 U163 ( .A(A[7]), .Y(n157) );
  NAND2BXL U164 ( .AN(B[10]), .B(A[10]), .Y(n129) );
  NAND2BXL U165 ( .AN(A[10]), .B(B[10]), .Y(n132) );
  NAND2BXL U166 ( .AN(A[10]), .B(B[10]), .Y(n91) );
  NOR2BX1 U167 ( .AN(A[6]), .B(B[6]), .Y(n12) );
  NAND2X1 U168 ( .A(A[7]), .B(n152), .Y(n30) );
  INVX1 U169 ( .A(B[7]), .Y(n152) );
  NAND2X1 U170 ( .A(B[5]), .B(n159), .Y(n156) );
  INVXL U171 ( .A(B[9]), .Y(n144) );
  NAND2X1 U172 ( .A(A[8]), .B(n147), .Y(n131) );
  NOR2X2 U173 ( .A(n118), .B(n119), .Y(n113) );
  INVX1 U174 ( .A(n108), .Y(n87) );
  NOR2BX1 U175 ( .AN(A[15]), .B(B[15]), .Y(n13) );
  NAND2X1 U176 ( .A(B[4]), .B(n160), .Y(n42) );
  NAND2X1 U177 ( .A(B[2]), .B(n169), .Y(n45) );
  NAND2X1 U178 ( .A(B[3]), .B(n166), .Y(n47) );
  NOR2BX1 U179 ( .AN(A[2]), .B(B[2]), .Y(n15) );
  NAND2X1 U180 ( .A(A[0]), .B(n172), .Y(n56) );
  INVX1 U181 ( .A(B[0]), .Y(n172) );
  NAND2X1 U182 ( .A(B[0]), .B(n171), .Y(n57) );
  INVX1 U183 ( .A(A[0]), .Y(n171) );
  INVXL U184 ( .A(A[11]), .Y(n136) );
  XNOR2X1 U185 ( .A(B[16]), .B(A[16]), .Y(n59) );
  NAND3X1 U186 ( .A(n60), .B(n61), .C(n62), .Y(n58) );
  NAND2X2 U187 ( .A(B[15]), .B(n99), .Y(n68) );
  INVXL U188 ( .A(A[14]), .Y(n67) );
  INVXL U189 ( .A(n72), .Y(n71) );
  NAND2XL U190 ( .A(n72), .B(n106), .Y(n102) );
  INVXL U191 ( .A(B[11]), .Y(n137) );
endmodule


module butterfly_DW01_sub_61 ( A, B, DIFF );
  input [16:0] A;
  input [16:0] B;
  output [16:0] DIFF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157;

  XOR2X1 U3 ( .A(n95), .B(n96), .Y(DIFF[15]) );
  NAND2X1 U4 ( .A(A[14]), .B(n107), .Y(n69) );
  NAND2X1 U5 ( .A(A[9]), .B(n132), .Y(n12) );
  OAI21XL U6 ( .A0(n126), .A1(n15), .B0(n17), .Y(n7) );
  AOI31X1 U7 ( .A0(n97), .A1(n85), .A2(n98), .B0(n99), .Y(n96) );
  OAI21XL U8 ( .A0(n68), .A1(n71), .B0(n69), .Y(n99) );
  OAI21XL U9 ( .A0(n135), .A1(n79), .B0(n94), .Y(n13) );
  NOR2X1 U10 ( .A(n100), .B(n101), .Y(n98) );
  NOR2X1 U11 ( .A(n9), .B(n10), .Y(n8) );
  INVX1 U12 ( .A(n12), .Y(n9) );
  XOR2X1 U13 ( .A(n113), .B(n114), .Y(DIFF[13]) );
  AOI21X1 U14 ( .A0(n115), .A1(n73), .B0(n116), .Y(n114) );
  XOR2X1 U15 ( .A(n103), .B(n104), .Y(DIFF[14]) );
  NOR2X1 U16 ( .A(n105), .B(n68), .Y(n104) );
  XOR2X1 U17 ( .A(n57), .B(n58), .Y(DIFF[16]) );
  BUFX8 U18 ( .A(B[13]), .Y(n6) );
  NAND2XL U19 ( .A(n73), .B(n85), .Y(n84) );
  CLKINVX3 U20 ( .A(n85), .Y(n68) );
  NAND2BX1 U21 ( .AN(B[12]), .B(A[12]), .Y(n70) );
  NAND2X1 U22 ( .A(B[14]), .B(n106), .Y(n85) );
  INVX1 U23 ( .A(n77), .Y(n67) );
  NAND2XL U24 ( .A(n89), .B(n124), .Y(n3) );
  NAND2X1 U25 ( .A(n108), .B(n71), .Y(n103) );
  INVXL U26 ( .A(n38), .Y(n40) );
  INVXL U27 ( .A(n37), .Y(n135) );
  AOI21XL U28 ( .A0(n91), .A1(n92), .B0(n93), .Y(n86) );
  INVXL U29 ( .A(n79), .Y(n91) );
  INVXL U30 ( .A(n94), .Y(n93) );
  NOR2XL U31 ( .A(n67), .B(n68), .Y(n64) );
  NOR2XL U32 ( .A(n22), .B(n26), .Y(n25) );
  NOR2XL U33 ( .A(n33), .B(n29), .Y(n32) );
  NAND2X1 U34 ( .A(n66), .B(n77), .Y(n95) );
  INVX1 U35 ( .A(n69), .Y(n105) );
  NAND2X1 U36 ( .A(n75), .B(n71), .Y(n113) );
  NAND2XL U37 ( .A(n110), .B(n111), .Y(n115) );
  NOR2XL U38 ( .A(n126), .B(n15), .Y(n125) );
  NAND2X1 U39 ( .A(n1), .B(n120), .Y(n118) );
  AND2X2 U40 ( .A(n123), .B(n124), .Y(n1) );
  NOR3XL U41 ( .A(n78), .B(n79), .C(n80), .Y(n74) );
  NOR2XL U42 ( .A(n67), .B(n68), .Y(n76) );
  XOR2X2 U43 ( .A(n2), .B(n119), .Y(DIFF[12]) );
  AND2X2 U44 ( .A(n73), .B(n70), .Y(n2) );
  NAND2XL U45 ( .A(n72), .B(n69), .Y(n62) );
  NAND3XL U46 ( .A(n69), .B(n70), .C(n71), .Y(n63) );
  INVXL U47 ( .A(n66), .Y(n65) );
  NOR2BX1 U48 ( .AN(n75), .B(n84), .Y(n83) );
  AOI21XL U49 ( .A0(n41), .A1(n34), .B0(n33), .Y(n137) );
  NAND2X1 U50 ( .A(n117), .B(n118), .Y(n87) );
  XNOR2X1 U51 ( .A(n130), .B(n3), .Y(DIFF[10]) );
  XNOR2X1 U52 ( .A(n127), .B(n128), .Y(DIFF[11]) );
  XOR2X1 U53 ( .A(n7), .B(n8), .Y(DIFF[9]) );
  NAND3BXL U54 ( .AN(n49), .B(n146), .C(n46), .Y(n80) );
  INVXL U55 ( .A(n27), .Y(n22) );
  NOR2XL U56 ( .A(n5), .B(n49), .Y(n48) );
  AOI21XL U57 ( .A0(n20), .A1(n21), .B0(n22), .Y(n19) );
  NAND2XL U58 ( .A(n23), .B(n24), .Y(n18) );
  NOR2XL U59 ( .A(n54), .B(n4), .Y(n53) );
  INVXL U60 ( .A(n51), .Y(n54) );
  NOR2XL U61 ( .A(n40), .B(n41), .Y(n39) );
  NAND2XL U62 ( .A(n46), .B(n47), .Y(n42) );
  NAND2BXL U63 ( .AN(A[13]), .B(n6), .Y(n75) );
  NAND2XL U64 ( .A(n102), .B(n112), .Y(n109) );
  NAND2BX1 U65 ( .AN(A[13]), .B(n6), .Y(n112) );
  NAND2BXL U66 ( .AN(A[12]), .B(B[12]), .Y(n73) );
  NAND2XL U67 ( .A(B[9]), .B(n155), .Y(n11) );
  NAND2BXL U68 ( .AN(A[10]), .B(B[10]), .Y(n89) );
  NAND2XL U69 ( .A(B[6]), .B(n143), .Y(n20) );
  NAND2XL U70 ( .A(B[7]), .B(n142), .Y(n23) );
  NAND2BXL U71 ( .AN(B[11]), .B(A[11]), .Y(n123) );
  INVXL U72 ( .A(B[8]), .Y(n133) );
  NAND2XL U73 ( .A(B[8]), .B(n134), .Y(n88) );
  NAND2BXL U74 ( .AN(A[11]), .B(B[11]), .Y(n90) );
  NOR2BXL U75 ( .AN(A[2]), .B(B[2]), .Y(n5) );
  NAND2XL U76 ( .A(B[2]), .B(n154), .Y(n44) );
  NAND2XL U77 ( .A(B[5]), .B(n144), .Y(n34) );
  NAND2XL U78 ( .A(B[4]), .B(n145), .Y(n38) );
  INVXL U79 ( .A(B[1]), .Y(n153) );
  INVXL U80 ( .A(B[6]), .Y(n139) );
  INVXL U81 ( .A(B[4]), .Y(n141) );
  INVXL U82 ( .A(B[3]), .Y(n150) );
  INVXL U83 ( .A(B[5]), .Y(n140) );
  INVX1 U84 ( .A(n13), .Y(n126) );
  XOR2X1 U85 ( .A(n21), .B(n25), .Y(DIFF[6]) );
  XOR2X1 U86 ( .A(n31), .B(n32), .Y(DIFF[5]) );
  OAI21XL U87 ( .A0(n86), .A1(n78), .B0(n87), .Y(n82) );
  NAND2BX1 U88 ( .AN(n92), .B(n80), .Y(n37) );
  NAND4X1 U89 ( .A(n125), .B(n11), .C(n89), .D(n90), .Y(n110) );
  NAND4X1 U90 ( .A(n38), .B(n34), .C(n20), .D(n23), .Y(n79) );
  OAI21XL U91 ( .A0(n28), .A1(n29), .B0(n30), .Y(n21) );
  INVX1 U92 ( .A(n31), .Y(n28) );
  NAND4X1 U93 ( .A(n11), .B(n88), .C(n89), .D(n90), .Y(n78) );
  AOI31X1 U94 ( .A0(n62), .A1(n63), .A2(n64), .B0(n65), .Y(n61) );
  NAND3X1 U95 ( .A(n110), .B(n70), .C(n111), .Y(n97) );
  NAND4X1 U96 ( .A(n73), .B(n74), .C(n75), .D(n76), .Y(n60) );
  INVX1 U97 ( .A(n88), .Y(n15) );
  NAND2X1 U98 ( .A(n131), .B(n12), .Y(n130) );
  NAND2X1 U99 ( .A(n11), .B(n7), .Y(n131) );
  NAND3X1 U100 ( .A(n121), .B(n11), .C(n122), .Y(n120) );
  NAND2X1 U101 ( .A(n17), .B(n12), .Y(n121) );
  NAND2X2 U102 ( .A(n110), .B(n87), .Y(n119) );
  INVX1 U103 ( .A(n11), .Y(n10) );
  XOR2X1 U104 ( .A(n18), .B(n19), .Y(DIFF[7]) );
  XOR2X1 U105 ( .A(n13), .B(n14), .Y(DIFF[8]) );
  NOR2X1 U106 ( .A(n15), .B(n16), .Y(n14) );
  INVX1 U107 ( .A(n17), .Y(n16) );
  NAND2X1 U108 ( .A(n117), .B(n118), .Y(n111) );
  NAND2X1 U109 ( .A(n23), .B(n136), .Y(n94) );
  OAI211X1 U110 ( .A0(n137), .A1(n26), .B0(n27), .C0(n24), .Y(n136) );
  INVX1 U111 ( .A(n34), .Y(n29) );
  INVX1 U112 ( .A(n36), .Y(n41) );
  NAND2X1 U113 ( .A(n123), .B(n90), .Y(n128) );
  INVX1 U114 ( .A(n30), .Y(n33) );
  INVX1 U115 ( .A(n102), .Y(n100) );
  INVX1 U116 ( .A(n20), .Y(n26) );
  INVX1 U117 ( .A(n70), .Y(n116) );
  NAND2BX1 U118 ( .AN(n109), .B(n97), .Y(n108) );
  NAND2X1 U119 ( .A(n124), .B(n129), .Y(n127) );
  NAND2X1 U120 ( .A(n130), .B(n89), .Y(n129) );
  OAI21XL U121 ( .A0(n50), .A1(n4), .B0(n51), .Y(n45) );
  INVX1 U122 ( .A(n52), .Y(n50) );
  OAI21XL U123 ( .A0(n148), .A1(n149), .B0(n47), .Y(n92) );
  AOI21X1 U124 ( .A0(n44), .A1(n152), .B0(n5), .Y(n148) );
  INVX1 U125 ( .A(n46), .Y(n149) );
  OAI21XL U126 ( .A0(n4), .A1(n55), .B0(n51), .Y(n152) );
  NOR2X1 U127 ( .A(n4), .B(n147), .Y(n146) );
  INVX1 U128 ( .A(n56), .Y(n147) );
  INVX1 U129 ( .A(n44), .Y(n49) );
  XOR2X1 U130 ( .A(n45), .B(n48), .Y(DIFF[2]) );
  XOR2X1 U131 ( .A(n42), .B(n43), .Y(DIFF[3]) );
  AOI21X1 U132 ( .A0(n44), .A1(n45), .B0(n5), .Y(n43) );
  XOR2X1 U133 ( .A(n52), .B(n53), .Y(DIFF[1]) );
  XOR2X1 U134 ( .A(n37), .B(n39), .Y(DIFF[4]) );
  NAND2X1 U135 ( .A(n35), .B(n36), .Y(n31) );
  NAND2X1 U136 ( .A(n37), .B(n38), .Y(n35) );
  NAND2BX1 U137 ( .AN(n56), .B(n55), .Y(n52) );
  NAND2X1 U138 ( .A(n55), .B(n56), .Y(DIFF[0]) );
  INVX1 U139 ( .A(A[9]), .Y(n155) );
  INVXL U140 ( .A(B[14]), .Y(n107) );
  NAND2BXL U141 ( .AN(B[10]), .B(A[10]), .Y(n124) );
  NAND2X1 U142 ( .A(A[8]), .B(n133), .Y(n17) );
  INVXL U143 ( .A(B[9]), .Y(n132) );
  INVX1 U144 ( .A(A[7]), .Y(n142) );
  INVX1 U145 ( .A(A[6]), .Y(n143) );
  INVX1 U146 ( .A(A[5]), .Y(n144) );
  INVX1 U147 ( .A(A[14]), .Y(n106) );
  NAND2X1 U148 ( .A(A[4]), .B(n141), .Y(n36) );
  NAND2X1 U149 ( .A(A[5]), .B(n140), .Y(n30) );
  NAND2BXL U150 ( .AN(A[11]), .B(B[11]), .Y(n117) );
  NAND2X1 U151 ( .A(A[7]), .B(n138), .Y(n24) );
  INVXL U152 ( .A(B[7]), .Y(n138) );
  INVX1 U153 ( .A(A[8]), .Y(n134) );
  NOR2BX1 U154 ( .AN(n6), .B(A[13]), .Y(n72) );
  NOR2BX1 U155 ( .AN(n6), .B(A[13]), .Y(n101) );
  NAND2X1 U156 ( .A(A[6]), .B(n139), .Y(n27) );
  XNOR2X1 U157 ( .A(B[16]), .B(A[16]), .Y(n58) );
  NAND3X1 U158 ( .A(n59), .B(n60), .C(n61), .Y(n57) );
  NAND3X1 U159 ( .A(n81), .B(n82), .C(n83), .Y(n59) );
  NAND2BXL U160 ( .AN(A[10]), .B(B[10]), .Y(n122) );
  NOR2BX1 U161 ( .AN(B[1]), .B(A[1]), .Y(n4) );
  NAND2X1 U162 ( .A(A[1]), .B(n153), .Y(n51) );
  INVX1 U163 ( .A(A[2]), .Y(n154) );
  INVX1 U164 ( .A(A[4]), .Y(n145) );
  NAND2X1 U165 ( .A(A[3]), .B(n150), .Y(n47) );
  NAND2X1 U166 ( .A(B[3]), .B(n151), .Y(n46) );
  INVX1 U167 ( .A(A[3]), .Y(n151) );
  NAND2X1 U168 ( .A(A[0]), .B(n157), .Y(n55) );
  INVX1 U169 ( .A(B[0]), .Y(n157) );
  NAND2X1 U170 ( .A(B[0]), .B(n156), .Y(n56) );
  INVX1 U171 ( .A(A[0]), .Y(n156) );
  NAND2BXL U172 ( .AN(A[15]), .B(B[15]), .Y(n81) );
  NAND2BX1 U173 ( .AN(B[15]), .B(A[15]), .Y(n66) );
  NAND2BX1 U174 ( .AN(A[15]), .B(B[15]), .Y(n77) );
  NAND2BXL U175 ( .AN(A[12]), .B(B[12]), .Y(n102) );
  NAND2BX4 U176 ( .AN(n6), .B(A[13]), .Y(n71) );
endmodule


module butterfly_DW01_sub_62 ( A, B, DIFF );
  input [16:0] A;
  input [16:0] B;
  output [16:0] DIFF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156;

  NAND2BX1 U3 ( .AN(A[15]), .B(B[15]), .Y(n78) );
  XNOR2X2 U4 ( .A(B[16]), .B(A[16]), .Y(n59) );
  NAND2BX4 U5 ( .AN(B[14]), .B(A[14]), .Y(n70) );
  OAI21X2 U6 ( .A0(n69), .A1(n72), .B0(n70), .Y(n99) );
  NAND4X1 U7 ( .A(n74), .B(n75), .C(n76), .D(n77), .Y(n61) );
  INVX4 U8 ( .A(n85), .Y(n69) );
  NAND2X2 U9 ( .A(B[14]), .B(n106), .Y(n85) );
  NAND2XL U10 ( .A(n73), .B(n70), .Y(n63) );
  INVX2 U11 ( .A(n70), .Y(n105) );
  NAND2X1 U12 ( .A(A[9]), .B(n131), .Y(n13) );
  XOR2X1 U13 ( .A(n103), .B(n104), .Y(DIFF[14]) );
  XOR2X1 U14 ( .A(n112), .B(n113), .Y(DIFF[13]) );
  AOI21XL U15 ( .A0(n114), .A1(n74), .B0(n115), .Y(n113) );
  XOR2X1 U16 ( .A(n95), .B(n96), .Y(DIFF[15]) );
  AOI31X1 U17 ( .A0(n97), .A1(n85), .A2(n98), .B0(n99), .Y(n96) );
  NOR2X1 U18 ( .A(n100), .B(n101), .Y(n98) );
  OAI21XL U19 ( .A0(n134), .A1(n80), .B0(n94), .Y(n14) );
  NAND2BX2 U20 ( .AN(A[13]), .B(n7), .Y(n111) );
  INVX1 U21 ( .A(n71), .Y(n115) );
  NOR2BX2 U22 ( .AN(n7), .B(A[13]), .Y(n101) );
  NOR2X1 U23 ( .A(n10), .B(n11), .Y(n9) );
  INVX1 U24 ( .A(n13), .Y(n10) );
  NAND2X1 U25 ( .A(n109), .B(n87), .Y(n118) );
  NAND2X1 U26 ( .A(n116), .B(n117), .Y(n110) );
  NAND2BX2 U27 ( .AN(n108), .B(n97), .Y(n107) );
  BUFX8 U28 ( .A(B[13]), .Y(n7) );
  NAND2X1 U29 ( .A(n102), .B(n111), .Y(n108) );
  NAND2BX2 U30 ( .AN(B[12]), .B(A[12]), .Y(n71) );
  NAND2X1 U31 ( .A(n116), .B(n117), .Y(n87) );
  NAND2XL U32 ( .A(n122), .B(n90), .Y(n127) );
  NAND2BX2 U33 ( .AN(B[11]), .B(A[11]), .Y(n122) );
  NAND2BX2 U34 ( .AN(A[12]), .B(B[12]), .Y(n74) );
  AND2X2 U35 ( .A(n122), .B(n123), .Y(n2) );
  XOR2X1 U36 ( .A(n3), .B(n118), .Y(DIFF[12]) );
  AOI21XL U37 ( .A0(n45), .A1(n46), .B0(n6), .Y(n44) );
  INVXL U38 ( .A(n39), .Y(n41) );
  NAND2X1 U39 ( .A(n36), .B(n37), .Y(n32) );
  INVXL U40 ( .A(n38), .Y(n134) );
  AOI21XL U41 ( .A0(n91), .A1(n92), .B0(n93), .Y(n86) );
  INVXL U42 ( .A(n80), .Y(n91) );
  INVXL U43 ( .A(n94), .Y(n93) );
  NOR2XL U44 ( .A(n23), .B(n27), .Y(n26) );
  NOR2XL U45 ( .A(n34), .B(n30), .Y(n33) );
  NAND2XL U46 ( .A(n67), .B(n78), .Y(n95) );
  NAND3XL U47 ( .A(n70), .B(n71), .C(n72), .Y(n64) );
  NOR3XL U48 ( .A(n79), .B(n80), .C(n81), .Y(n75) );
  NOR2BX1 U49 ( .AN(n76), .B(n1), .Y(n84) );
  NAND2XL U50 ( .A(n74), .B(n85), .Y(n1) );
  OAI21X1 U51 ( .A0(n125), .A1(n16), .B0(n18), .Y(n8) );
  NOR2XL U52 ( .A(n125), .B(n16), .Y(n124) );
  NAND2X1 U53 ( .A(n2), .B(n119), .Y(n117) );
  AOI21XL U54 ( .A0(n42), .A1(n35), .B0(n34), .Y(n136) );
  AND2X2 U55 ( .A(n74), .B(n71), .Y(n3) );
  XNOR2X1 U56 ( .A(n129), .B(n4), .Y(DIFF[10]) );
  NAND2XL U57 ( .A(n89), .B(n123), .Y(n4) );
  XNOR2X1 U58 ( .A(n126), .B(n127), .Y(DIFF[11]) );
  XOR2X1 U59 ( .A(n8), .B(n9), .Y(DIFF[9]) );
  INVXL U60 ( .A(n102), .Y(n100) );
  NAND3BXL U61 ( .AN(n50), .B(n145), .C(n47), .Y(n81) );
  INVXL U62 ( .A(n28), .Y(n23) );
  NOR2XL U63 ( .A(n6), .B(n50), .Y(n49) );
  AOI21XL U64 ( .A0(n21), .A1(n22), .B0(n23), .Y(n20) );
  NAND2XL U65 ( .A(n24), .B(n25), .Y(n19) );
  NOR2XL U66 ( .A(n55), .B(n5), .Y(n54) );
  INVXL U67 ( .A(n52), .Y(n55) );
  NOR2XL U68 ( .A(n41), .B(n42), .Y(n40) );
  NAND2XL U69 ( .A(n47), .B(n48), .Y(n43) );
  NAND2BXL U70 ( .AN(A[13]), .B(n7), .Y(n76) );
  XOR2X1 U71 ( .A(n58), .B(n59), .Y(DIFF[16]) );
  NAND2XL U72 ( .A(B[9]), .B(n154), .Y(n12) );
  NAND2BXL U73 ( .AN(A[10]), .B(B[10]), .Y(n89) );
  NAND2BXL U74 ( .AN(A[11]), .B(B[11]), .Y(n90) );
  NAND2XL U75 ( .A(B[6]), .B(n142), .Y(n21) );
  NAND2XL U76 ( .A(B[7]), .B(n141), .Y(n24) );
  INVXL U77 ( .A(B[8]), .Y(n132) );
  NAND2XL U78 ( .A(B[8]), .B(n133), .Y(n88) );
  NOR2BXL U79 ( .AN(A[2]), .B(B[2]), .Y(n6) );
  NAND2XL U80 ( .A(B[2]), .B(n153), .Y(n45) );
  NAND2XL U81 ( .A(B[5]), .B(n143), .Y(n35) );
  NAND2XL U82 ( .A(B[4]), .B(n144), .Y(n39) );
  INVXL U83 ( .A(B[1]), .Y(n152) );
  INVXL U84 ( .A(B[6]), .Y(n138) );
  INVXL U85 ( .A(B[4]), .Y(n140) );
  INVXL U86 ( .A(B[3]), .Y(n149) );
  INVXL U87 ( .A(B[5]), .Y(n139) );
  INVX1 U88 ( .A(n14), .Y(n125) );
  XOR2X1 U89 ( .A(n22), .B(n26), .Y(DIFF[6]) );
  XOR2X1 U90 ( .A(n32), .B(n33), .Y(DIFF[5]) );
  OAI21XL U91 ( .A0(n86), .A1(n79), .B0(n87), .Y(n83) );
  NAND2BX1 U92 ( .AN(n92), .B(n81), .Y(n38) );
  NAND4X1 U93 ( .A(n124), .B(n12), .C(n89), .D(n90), .Y(n109) );
  NAND4X1 U94 ( .A(n39), .B(n35), .C(n21), .D(n24), .Y(n80) );
  OAI21XL U95 ( .A0(n29), .A1(n30), .B0(n31), .Y(n22) );
  INVX1 U96 ( .A(n32), .Y(n29) );
  NAND4X1 U97 ( .A(n12), .B(n88), .C(n89), .D(n90), .Y(n79) );
  AOI31X1 U98 ( .A0(n63), .A1(n64), .A2(n65), .B0(n66), .Y(n62) );
  INVX1 U99 ( .A(n67), .Y(n66) );
  NAND3X1 U100 ( .A(n109), .B(n71), .C(n110), .Y(n97) );
  INVX1 U101 ( .A(n88), .Y(n16) );
  NAND2X1 U102 ( .A(n130), .B(n13), .Y(n129) );
  NAND2X1 U103 ( .A(n12), .B(n8), .Y(n130) );
  NAND3X1 U104 ( .A(n120), .B(n12), .C(n121), .Y(n119) );
  NAND2X1 U105 ( .A(n18), .B(n13), .Y(n120) );
  INVX1 U106 ( .A(n12), .Y(n11) );
  XOR2X1 U107 ( .A(n19), .B(n20), .Y(DIFF[7]) );
  XOR2X1 U108 ( .A(n14), .B(n15), .Y(DIFF[8]) );
  NOR2X1 U109 ( .A(n16), .B(n17), .Y(n15) );
  INVX1 U110 ( .A(n18), .Y(n17) );
  NAND2X1 U111 ( .A(n123), .B(n128), .Y(n126) );
  NAND2X1 U112 ( .A(n129), .B(n89), .Y(n128) );
  NAND2X1 U113 ( .A(n24), .B(n135), .Y(n94) );
  OAI211X1 U114 ( .A0(n136), .A1(n27), .B0(n28), .C0(n25), .Y(n135) );
  INVX1 U115 ( .A(n35), .Y(n30) );
  INVX1 U116 ( .A(n31), .Y(n34) );
  NAND2X1 U117 ( .A(n76), .B(n72), .Y(n112) );
  NAND2X1 U118 ( .A(n109), .B(n110), .Y(n114) );
  INVX1 U119 ( .A(n21), .Y(n27) );
  NAND2X2 U120 ( .A(n107), .B(n72), .Y(n103) );
  NOR2X2 U121 ( .A(n105), .B(n69), .Y(n104) );
  INVX1 U122 ( .A(n78), .Y(n68) );
  OAI21XL U123 ( .A0(n51), .A1(n5), .B0(n52), .Y(n46) );
  INVX1 U124 ( .A(n53), .Y(n51) );
  OAI21XL U125 ( .A0(n147), .A1(n148), .B0(n48), .Y(n92) );
  AOI21X1 U126 ( .A0(n45), .A1(n151), .B0(n6), .Y(n147) );
  INVX1 U127 ( .A(n47), .Y(n148) );
  OAI21XL U128 ( .A0(n5), .A1(n56), .B0(n52), .Y(n151) );
  NOR2X1 U129 ( .A(n5), .B(n146), .Y(n145) );
  INVX1 U130 ( .A(n57), .Y(n146) );
  INVX1 U131 ( .A(n45), .Y(n50) );
  XOR2X1 U132 ( .A(n46), .B(n49), .Y(DIFF[2]) );
  XOR2X1 U133 ( .A(n43), .B(n44), .Y(DIFF[3]) );
  XOR2X1 U134 ( .A(n53), .B(n54), .Y(DIFF[1]) );
  XOR2X1 U135 ( .A(n38), .B(n40), .Y(DIFF[4]) );
  NAND2X1 U136 ( .A(n38), .B(n39), .Y(n36) );
  INVX1 U137 ( .A(n37), .Y(n42) );
  NAND2BX1 U138 ( .AN(n57), .B(n56), .Y(n53) );
  NAND2X1 U139 ( .A(n56), .B(n57), .Y(DIFF[0]) );
  INVX1 U140 ( .A(A[9]), .Y(n154) );
  NAND2BXL U141 ( .AN(B[10]), .B(A[10]), .Y(n123) );
  NAND2X1 U142 ( .A(A[8]), .B(n132), .Y(n18) );
  INVXL U143 ( .A(B[9]), .Y(n131) );
  INVX1 U144 ( .A(A[7]), .Y(n141) );
  INVX1 U145 ( .A(A[6]), .Y(n142) );
  INVX1 U146 ( .A(A[5]), .Y(n143) );
  INVX1 U147 ( .A(A[14]), .Y(n106) );
  NOR2BX1 U148 ( .AN(n7), .B(A[13]), .Y(n73) );
  NAND2X1 U149 ( .A(A[5]), .B(n139), .Y(n31) );
  NAND2BXL U150 ( .AN(A[11]), .B(B[11]), .Y(n116) );
  NAND2X1 U151 ( .A(A[7]), .B(n137), .Y(n25) );
  INVXL U152 ( .A(B[7]), .Y(n137) );
  INVX1 U153 ( .A(A[8]), .Y(n133) );
  NAND2X1 U154 ( .A(A[6]), .B(n138), .Y(n28) );
  NAND3X1 U155 ( .A(n60), .B(n61), .C(n62), .Y(n58) );
  NAND3X1 U156 ( .A(n82), .B(n83), .C(n84), .Y(n60) );
  NAND2BXL U157 ( .AN(A[10]), .B(B[10]), .Y(n121) );
  NOR2BX1 U158 ( .AN(B[1]), .B(A[1]), .Y(n5) );
  NAND2X1 U159 ( .A(A[1]), .B(n152), .Y(n52) );
  INVX1 U160 ( .A(A[2]), .Y(n153) );
  INVX1 U161 ( .A(A[4]), .Y(n144) );
  NAND2X1 U162 ( .A(A[3]), .B(n149), .Y(n48) );
  NAND2X1 U163 ( .A(B[3]), .B(n150), .Y(n47) );
  INVX1 U164 ( .A(A[3]), .Y(n150) );
  NAND2X1 U165 ( .A(A[4]), .B(n140), .Y(n37) );
  NAND2X1 U166 ( .A(A[0]), .B(n156), .Y(n56) );
  INVX1 U167 ( .A(B[0]), .Y(n156) );
  NAND2X1 U168 ( .A(B[0]), .B(n155), .Y(n57) );
  INVX1 U169 ( .A(A[0]), .Y(n155) );
  NAND2BXL U170 ( .AN(A[15]), .B(B[15]), .Y(n82) );
  NAND2BX1 U171 ( .AN(B[15]), .B(A[15]), .Y(n67) );
  NOR2XL U172 ( .A(n68), .B(n69), .Y(n65) );
  NOR2XL U173 ( .A(n68), .B(n69), .Y(n77) );
  NAND2BXL U174 ( .AN(A[12]), .B(B[12]), .Y(n102) );
  NAND2BX4 U175 ( .AN(n7), .B(A[13]), .Y(n72) );
endmodule


module butterfly_DW01_add_81 ( A, B, SUM );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131;

  AOI21X1 U2 ( .A0(B[11]), .A1(A[11]), .B0(n102), .Y(n113) );
  INVX2 U3 ( .A(n75), .Y(n102) );
  XOR2X1 U4 ( .A(n115), .B(n116), .Y(SUM[10]) );
  NAND2X1 U5 ( .A(n58), .B(n60), .Y(n92) );
  NOR2BX1 U6 ( .AN(n63), .B(n5), .Y(n82) );
  INVX1 U7 ( .A(B[12]), .Y(n99) );
  OAI21XL U8 ( .A0(n10), .A1(n117), .B0(n9), .Y(n115) );
  NAND2BX1 U9 ( .AN(A[12]), .B(n99), .Y(n90) );
  NAND2X1 U10 ( .A(B[13]), .B(A[13]), .Y(n91) );
  NAND2BX1 U11 ( .AN(A[11]), .B(n110), .Y(n75) );
  OR2X2 U12 ( .A(B[9]), .B(A[9]), .Y(n76) );
  OAI21XL U13 ( .A0(n120), .A1(n18), .B0(n19), .Y(n80) );
  OAI21XL U14 ( .A0(n27), .A1(n32), .B0(n28), .Y(n122) );
  NAND2X1 U15 ( .A(B[14]), .B(A[14]), .Y(n58) );
  OR2X2 U16 ( .A(A[13]), .B(B[13]), .Y(n71) );
  AND2X2 U17 ( .A(n51), .B(n126), .Y(SUM[0]) );
  XOR2X1 U18 ( .A(n112), .B(n113), .Y(SUM[11]) );
  NAND2XL U19 ( .A(B[15]), .B(A[15]), .Y(n63) );
  NAND2X1 U20 ( .A(n91), .B(n71), .Y(n95) );
  NAND2XL U21 ( .A(n71), .B(n60), .Y(n84) );
  NAND2XL U22 ( .A(n71), .B(n94), .Y(n93) );
  NOR2X1 U23 ( .A(B[3]), .B(A[3]), .Y(n4) );
  AOI21XL U24 ( .A0(n44), .A1(n128), .B0(n129), .Y(n127) );
  OAI21X1 U25 ( .A0(n83), .A1(n84), .B0(n58), .Y(n81) );
  NAND2XL U26 ( .A(n87), .B(n73), .Y(n101) );
  NAND2X1 U27 ( .A(n91), .B(n93), .Y(n2) );
  AOI21X1 U28 ( .A0(n57), .A1(n58), .B0(n5), .Y(n56) );
  NAND4X1 U29 ( .A(n34), .B(n124), .C(n25), .D(n121), .Y(n67) );
  NAND2BXL U30 ( .AN(A[11]), .B(n110), .Y(n109) );
  NAND2XL U31 ( .A(n115), .B(n74), .Y(n114) );
  NAND2XL U32 ( .A(B[10]), .B(A[10]), .Y(n104) );
  OR2XL U33 ( .A(B[8]), .B(A[8]), .Y(n77) );
  INVXL U34 ( .A(n79), .Y(n125) );
  XOR2X1 U35 ( .A(n81), .B(n82), .Y(SUM[15]) );
  NOR2XL U36 ( .A(n85), .B(n86), .Y(n83) );
  NOR2BXL U37 ( .AN(n63), .B(n56), .Y(n55) );
  NAND3X1 U38 ( .A(n62), .B(n96), .C(n97), .Y(n94) );
  NAND2X1 U39 ( .A(n98), .B(n90), .Y(n97) );
  XNOR2X1 U40 ( .A(n100), .B(n101), .Y(SUM[12]) );
  NAND2XL U41 ( .A(n62), .B(n90), .Y(n100) );
  XNOR2X1 U42 ( .A(n94), .B(n95), .Y(SUM[13]) );
  XNOR2X2 U43 ( .A(n2), .B(n92), .Y(SUM[14]) );
  OAI2BB2X1 U44 ( .B0(n65), .B1(n87), .A0N(n89), .A1N(n3), .Y(n86) );
  AND2X1 U45 ( .A(n88), .B(n75), .Y(n3) );
  AOI21XL U46 ( .A0(n78), .A1(n79), .B0(n80), .Y(n72) );
  INVX2 U47 ( .A(n76), .Y(n10) );
  INVXL U48 ( .A(n90), .Y(n65) );
  NAND2X1 U49 ( .A(n118), .B(n13), .Y(n7) );
  XOR2X1 U50 ( .A(n7), .B(n8), .Y(SUM[9]) );
  NOR2BXL U51 ( .AN(n9), .B(n10), .Y(n8) );
  INVXL U52 ( .A(n29), .Y(n26) );
  NOR2BXL U53 ( .AN(n28), .B(n27), .Y(n30) );
  NOR2XL U54 ( .A(n17), .B(n18), .Y(n16) );
  INVXL U55 ( .A(n23), .Y(n20) );
  INVXL U56 ( .A(n25), .Y(n21) );
  NAND2XL U57 ( .A(n47), .B(n48), .Y(n45) );
  NOR2BXL U58 ( .AN(n46), .B(n50), .Y(n49) );
  INVXL U59 ( .A(n44), .Y(n40) );
  NAND2XL U60 ( .A(B[12]), .B(A[12]), .Y(n62) );
  NOR2XL U61 ( .A(A[15]), .B(B[15]), .Y(n5) );
  OR2XL U62 ( .A(B[14]), .B(A[14]), .Y(n60) );
  NAND2BX1 U63 ( .AN(A[12]), .B(n99), .Y(n88) );
  NAND3X1 U64 ( .A(n103), .B(n104), .C(n105), .Y(n89) );
  NAND2XL U65 ( .A(B[8]), .B(A[8]), .Y(n13) );
  NAND2X1 U66 ( .A(n104), .B(n114), .Y(n112) );
  NAND4X1 U67 ( .A(n108), .B(n76), .C(n74), .D(n109), .Y(n87) );
  INVXL U68 ( .A(n11), .Y(n111) );
  NAND2XL U69 ( .A(B[6]), .B(A[6]), .Y(n22) );
  NAND2XL U70 ( .A(B[7]), .B(A[7]), .Y(n19) );
  OR2X2 U71 ( .A(B[10]), .B(A[10]), .Y(n74) );
  NAND2XL U72 ( .A(B[5]), .B(A[5]), .Y(n28) );
  OR2XL U73 ( .A(B[4]), .B(A[4]), .Y(n34) );
  NAND2XL U74 ( .A(B[1]), .B(A[1]), .Y(n46) );
  NAND2XL U75 ( .A(B[3]), .B(A[3]), .Y(n38) );
  INVX1 U76 ( .A(B[11]), .Y(n110) );
  INVX1 U77 ( .A(B[0]), .Y(n130) );
  OAI21XL U78 ( .A0(n125), .A1(n67), .B0(n119), .Y(n11) );
  INVX1 U79 ( .A(n80), .Y(n119) );
  INVX1 U80 ( .A(n7), .Y(n117) );
  OAI21XL U81 ( .A0(n127), .A1(n4), .B0(n38), .Y(n79) );
  INVX1 U82 ( .A(n41), .Y(n129) );
  OAI21XL U83 ( .A0(n50), .A1(n51), .B0(n46), .Y(n128) );
  OAI21XL U84 ( .A0(n26), .A1(n27), .B0(n28), .Y(n23) );
  OAI21XL U85 ( .A0(n31), .A1(n125), .B0(n32), .Y(n29) );
  AOI21X1 U86 ( .A0(n25), .A1(n122), .B0(n123), .Y(n120) );
  INVX1 U87 ( .A(n22), .Y(n123) );
  NOR3X1 U88 ( .A(n64), .B(n65), .C(n61), .Y(n70) );
  INVX1 U89 ( .A(n60), .Y(n64) );
  NAND3X1 U90 ( .A(n88), .B(n75), .C(n89), .Y(n96) );
  INVX1 U91 ( .A(n87), .Y(n98) );
  INVX1 U92 ( .A(n124), .Y(n27) );
  XOR2X1 U93 ( .A(n11), .B(n12), .Y(SUM[8]) );
  NOR2BX1 U94 ( .AN(n13), .B(n14), .Y(n12) );
  OAI21XL U95 ( .A0(n72), .A1(n66), .B0(n73), .Y(n69) );
  NAND4XL U96 ( .A(n74), .B(n75), .C(n76), .D(n77), .Y(n66) );
  INVX1 U97 ( .A(n67), .Y(n78) );
  NAND2BX1 U98 ( .AN(n102), .B(n89), .Y(n73) );
  NOR2BX1 U99 ( .AN(n104), .B(n106), .Y(n116) );
  XOR2X1 U100 ( .A(n29), .B(n30), .Y(SUM[5]) );
  XOR2X1 U101 ( .A(n23), .B(n24), .Y(SUM[6]) );
  NOR2BX1 U102 ( .AN(n22), .B(n21), .Y(n24) );
  XOR2X1 U103 ( .A(n15), .B(n16), .Y(SUM[7]) );
  OAI21XL U104 ( .A0(n20), .A1(n21), .B0(n22), .Y(n15) );
  NAND2X1 U105 ( .A(n11), .B(n77), .Y(n118) );
  INVX1 U106 ( .A(n34), .Y(n31) );
  INVX1 U107 ( .A(n47), .Y(n50) );
  INVX1 U108 ( .A(n77), .Y(n14) );
  INVX1 U109 ( .A(n121), .Y(n18) );
  NAND2XL U110 ( .A(n91), .B(n62), .Y(n85) );
  INVX1 U111 ( .A(n74), .Y(n106) );
  INVX1 U112 ( .A(n19), .Y(n17) );
  XOR2X1 U113 ( .A(n48), .B(n49), .Y(SUM[1]) );
  XOR2X1 U114 ( .A(n42), .B(n43), .Y(SUM[2]) );
  NOR2BX1 U115 ( .AN(n41), .B(n40), .Y(n43) );
  XOR2X1 U116 ( .A(n79), .B(n33), .Y(SUM[4]) );
  NOR2BX1 U117 ( .AN(n32), .B(n31), .Y(n33) );
  XOR2X1 U118 ( .A(n35), .B(n36), .Y(SUM[3]) );
  OAI21XL U119 ( .A0(n39), .A1(n40), .B0(n41), .Y(n35) );
  NOR2X1 U120 ( .A(n37), .B(n4), .Y(n36) );
  INVX1 U121 ( .A(n42), .Y(n39) );
  NAND2X1 U122 ( .A(n45), .B(n46), .Y(n42) );
  INVX1 U123 ( .A(n38), .Y(n37) );
  INVX1 U124 ( .A(n51), .Y(n48) );
  NOR2X1 U125 ( .A(n111), .B(n14), .Y(n108) );
  NAND2BXL U126 ( .AN(n106), .B(n107), .Y(n103) );
  OAI21XL U127 ( .A0(n10), .A1(n13), .B0(n9), .Y(n107) );
  NAND2X1 U128 ( .A(B[4]), .B(A[4]), .Y(n32) );
  NAND2XL U129 ( .A(B[9]), .B(A[9]), .Y(n9) );
  NAND2X1 U130 ( .A(B[2]), .B(A[2]), .Y(n41) );
  OR2X2 U131 ( .A(B[6]), .B(A[6]), .Y(n25) );
  OR2X2 U132 ( .A(B[7]), .B(A[7]), .Y(n121) );
  OR2X2 U133 ( .A(B[5]), .B(A[5]), .Y(n124) );
  OR2X2 U134 ( .A(B[2]), .B(A[2]), .Y(n44) );
  OR2X2 U135 ( .A(B[1]), .B(A[1]), .Y(n47) );
  XOR2X2 U136 ( .A(n52), .B(n53), .Y(SUM[16]) );
  XOR2X1 U137 ( .A(B[16]), .B(A[16]), .Y(n53) );
  NAND2X1 U138 ( .A(n54), .B(n55), .Y(n52) );
  NAND3BX1 U139 ( .AN(n68), .B(n69), .C(n70), .Y(n54) );
  AND2X1 U140 ( .A(B[13]), .B(A[13]), .Y(n6) );
  NAND2X1 U141 ( .A(B[0]), .B(A[0]), .Y(n51) );
  NAND2X1 U142 ( .A(n130), .B(n131), .Y(n126) );
  INVX1 U143 ( .A(A[0]), .Y(n131) );
  NAND2XL U144 ( .A(B[11]), .B(A[11]), .Y(n105) );
  NOR2XL U145 ( .A(n61), .B(n62), .Y(n59) );
  OAI21XL U146 ( .A0(n6), .A1(n59), .B0(n60), .Y(n57) );
  NOR2XL U147 ( .A(A[13]), .B(B[13]), .Y(n61) );
  NOR2XL U148 ( .A(A[15]), .B(B[15]), .Y(n68) );
endmodule


module butterfly_DW01_add_86 ( A, B, SUM );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  wire   n1, n2, n3, n4, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149;

  NAND2X4 U2 ( .A(n103), .B(n7), .Y(n8) );
  NAND2X2 U3 ( .A(n80), .B(n87), .Y(n116) );
  NAND2BX2 U4 ( .AN(A[10]), .B(n123), .Y(n86) );
  INVX2 U5 ( .A(B[10]), .Y(n123) );
  NOR3X2 U6 ( .A(n1), .B(n2), .C(n3), .Y(n4) );
  NOR2X2 U7 ( .A(n4), .B(n116), .Y(n115) );
  INVX1 U8 ( .A(n109), .Y(n1) );
  INVX1 U9 ( .A(n110), .Y(n2) );
  INVX1 U10 ( .A(n111), .Y(n3) );
  NAND2X4 U11 ( .A(n131), .B(n132), .Y(n87) );
  INVX2 U12 ( .A(A[11]), .Y(n132) );
  NOR2X2 U13 ( .A(n102), .B(n109), .Y(n121) );
  INVX3 U14 ( .A(n110), .Y(n85) );
  NAND2X2 U15 ( .A(B[11]), .B(A[11]), .Y(n110) );
  XOR2X2 U16 ( .A(n11), .B(n114), .Y(SUM[13]) );
  INVX2 U17 ( .A(n104), .Y(n7) );
  OAI21X1 U18 ( .A0(n133), .A1(n134), .B0(n125), .Y(n129) );
  XOR2X2 U19 ( .A(n135), .B(n136), .Y(SUM[10]) );
  OAI21XL U20 ( .A0(n35), .A1(n36), .B0(n37), .Y(n32) );
  NAND2X1 U21 ( .A(n100), .B(n73), .Y(n106) );
  AND3X2 U22 ( .A(n10), .B(n87), .C(n80), .Y(n105) );
  OR2XL U23 ( .A(A[13]), .B(B[13]), .Y(n10) );
  NAND2X1 U24 ( .A(n124), .B(n125), .Y(n117) );
  OAI21XL U25 ( .A0(n19), .A1(n22), .B0(n18), .Y(n126) );
  INVX2 U26 ( .A(B[11]), .Y(n131) );
  NAND2BX1 U27 ( .AN(n72), .B(n107), .Y(n100) );
  OAI21XL U28 ( .A0(n19), .A1(n137), .B0(n18), .Y(n135) );
  INVX1 U29 ( .A(n16), .Y(n137) );
  CLKINVX3 U30 ( .A(n86), .Y(n134) );
  NAND2X1 U31 ( .A(B[10]), .B(A[10]), .Y(n125) );
  OAI21XL U32 ( .A0(n40), .A1(n41), .B0(n42), .Y(n38) );
  NAND2BX1 U33 ( .AN(A[13]), .B(n108), .Y(n82) );
  NAND4X1 U34 ( .A(n24), .B(n20), .C(n88), .D(n122), .Y(n109) );
  NAND2X1 U35 ( .A(B[12]), .B(A[12]), .Y(n72) );
  NAND2X1 U36 ( .A(B[13]), .B(A[13]), .Y(n73) );
  XNOR2X2 U37 ( .A(n25), .B(n12), .Y(SUM[7]) );
  OR2X2 U38 ( .A(n26), .B(n27), .Y(n12) );
  NAND2X1 U39 ( .A(n100), .B(n73), .Y(n99) );
  XOR2X2 U40 ( .A(n16), .B(n17), .Y(SUM[9]) );
  INVX1 U41 ( .A(n103), .Y(n6) );
  AND2X2 U42 ( .A(n61), .B(n145), .Y(SUM[0]) );
  INVX2 U43 ( .A(B[14]), .Y(n112) );
  AOI21X1 U44 ( .A0(n97), .A1(n98), .B0(n99), .Y(n95) );
  NAND2X1 U45 ( .A(n72), .B(n80), .Y(n119) );
  AOI21XL U46 ( .A0(n68), .A1(n69), .B0(n15), .Y(n67) );
  CLKINVX4 U47 ( .A(A[12]), .Y(n128) );
  NOR2X2 U48 ( .A(n74), .B(n75), .Y(n70) );
  NOR2BX4 U49 ( .AN(n110), .B(n102), .Y(n130) );
  AND2X2 U50 ( .A(n117), .B(n87), .Y(n14) );
  INVX4 U51 ( .A(n87), .Y(n102) );
  NOR2BX2 U52 ( .AN(n72), .B(n115), .Y(n114) );
  INVX4 U53 ( .A(A[14]), .Y(n113) );
  INVX4 U54 ( .A(B[13]), .Y(n108) );
  NAND2X2 U55 ( .A(n6), .B(n104), .Y(n9) );
  NAND2X4 U56 ( .A(n8), .B(n9), .Y(SUM[14]) );
  NAND2X2 U57 ( .A(B[14]), .B(A[14]), .Y(n69) );
  NOR3XL U58 ( .A(n15), .B(n75), .C(n74), .Y(n81) );
  INVX2 U59 ( .A(n94), .Y(n66) );
  XOR2X4 U60 ( .A(n92), .B(n93), .Y(SUM[15]) );
  NOR2X2 U61 ( .A(n15), .B(n66), .Y(n93) );
  INVXL U62 ( .A(n80), .Y(n76) );
  NOR2X1 U63 ( .A(B[15]), .B(A[15]), .Y(n15) );
  INVX1 U64 ( .A(n135), .Y(n133) );
  NOR2BX1 U65 ( .AN(n31), .B(n30), .Y(n33) );
  NOR2BX2 U66 ( .AN(n18), .B(n19), .Y(n17) );
  INVX1 U67 ( .A(n117), .Y(n111) );
  INVX1 U68 ( .A(n90), .Y(n41) );
  OAI21XL U69 ( .A0(n83), .A1(n77), .B0(n84), .Y(n79) );
  NAND3XL U70 ( .A(n79), .B(n80), .C(n81), .Y(n64) );
  NAND3XL U71 ( .A(n109), .B(n110), .C(n111), .Y(n98) );
  OAI21XL U72 ( .A0(A[10]), .A1(B[10]), .B0(n126), .Y(n124) );
  OAI21X2 U73 ( .A0(n41), .A1(n78), .B0(n139), .Y(n20) );
  NOR2XL U74 ( .A(n85), .B(n14), .Y(n84) );
  INVXL U75 ( .A(n78), .Y(n89) );
  OAI21X2 U76 ( .A0(n95), .A1(n74), .B0(n69), .Y(n92) );
  INVX4 U77 ( .A(n88), .Y(n19) );
  NOR2BX4 U78 ( .AN(n125), .B(n134), .Y(n136) );
  NAND2X2 U79 ( .A(n82), .B(n118), .Y(n11) );
  INVX4 U80 ( .A(n96), .Y(n74) );
  AOI21XL U81 ( .A0(n34), .A1(n142), .B0(n143), .Y(n140) );
  NOR2BXL U82 ( .AN(n56), .B(n60), .Y(n59) );
  NAND2XL U83 ( .A(n57), .B(n58), .Y(n55) );
  INVXL U84 ( .A(n54), .Y(n50) );
  INVXL U85 ( .A(n48), .Y(n47) );
  NAND2BXL U86 ( .AN(B[0]), .B(n149), .Y(n145) );
  NAND2BXL U87 ( .AN(A[10]), .B(n123), .Y(n122) );
  XOR2X2 U88 ( .A(B[16]), .B(A[16]), .Y(n63) );
  NAND2XL U89 ( .A(B[6]), .B(A[6]), .Y(n31) );
  NAND2XL U90 ( .A(B[4]), .B(A[4]), .Y(n42) );
  NAND2XL U91 ( .A(B[5]), .B(A[5]), .Y(n37) );
  NAND2XL U92 ( .A(B[7]), .B(A[7]), .Y(n28) );
  NOR2X1 U93 ( .A(B[3]), .B(A[3]), .Y(n13) );
  NAND2XL U94 ( .A(B[0]), .B(A[0]), .Y(n61) );
  NAND2XL U95 ( .A(B[1]), .B(A[1]), .Y(n56) );
  INVXL U96 ( .A(A[0]), .Y(n149) );
  INVX1 U97 ( .A(n91), .Y(n139) );
  XOR2X2 U98 ( .A(n20), .B(n21), .Y(SUM[8]) );
  NOR2BX1 U99 ( .AN(n22), .B(n23), .Y(n21) );
  INVX1 U100 ( .A(n24), .Y(n23) );
  XOR2X1 U101 ( .A(n32), .B(n33), .Y(SUM[6]) );
  XOR2X1 U102 ( .A(n38), .B(n39), .Y(SUM[5]) );
  NOR2BX1 U103 ( .AN(n37), .B(n36), .Y(n39) );
  OAI21XL U104 ( .A0(n29), .A1(n30), .B0(n31), .Y(n25) );
  INVX1 U105 ( .A(n32), .Y(n29) );
  XOR2X1 U106 ( .A(n45), .B(n46), .Y(SUM[3]) );
  OAI21XL U107 ( .A0(n49), .A1(n50), .B0(n51), .Y(n45) );
  NOR2X1 U108 ( .A(n47), .B(n13), .Y(n46) );
  INVX1 U109 ( .A(n52), .Y(n49) );
  XOR2X1 U110 ( .A(n90), .B(n43), .Y(SUM[4]) );
  NOR2BX1 U111 ( .AN(n42), .B(n40), .Y(n43) );
  XOR2X1 U112 ( .A(n58), .B(n59), .Y(SUM[1]) );
  NAND2X1 U113 ( .A(n70), .B(n71), .Y(n68) );
  NAND2XL U114 ( .A(n72), .B(n73), .Y(n71) );
  OAI21XL U115 ( .A0(n146), .A1(n13), .B0(n48), .Y(n90) );
  AOI21X1 U116 ( .A0(n54), .A1(n147), .B0(n148), .Y(n146) );
  INVX1 U117 ( .A(n51), .Y(n148) );
  OAI21XL U118 ( .A0(n60), .A1(n61), .B0(n56), .Y(n147) );
  INVX1 U119 ( .A(n38), .Y(n35) );
  OAI21XL U120 ( .A0(n140), .A1(n27), .B0(n28), .Y(n91) );
  INVX1 U121 ( .A(n31), .Y(n143) );
  OAI21XL U122 ( .A0(n36), .A1(n42), .B0(n37), .Y(n142) );
  NAND4X1 U123 ( .A(n44), .B(n144), .C(n34), .D(n141), .Y(n78) );
  INVX1 U124 ( .A(n144), .Y(n36) );
  NAND4XL U125 ( .A(n86), .B(n87), .C(n88), .D(n24), .Y(n77) );
  AOI21XL U126 ( .A0(n89), .A1(n90), .B0(n91), .Y(n83) );
  INVX1 U127 ( .A(n34), .Y(n30) );
  INVX1 U128 ( .A(n44), .Y(n40) );
  INVX1 U129 ( .A(n57), .Y(n60) );
  INVX1 U130 ( .A(n141), .Y(n27) );
  INVX1 U131 ( .A(n82), .Y(n75) );
  INVX1 U132 ( .A(n28), .Y(n26) );
  XOR2X1 U133 ( .A(n52), .B(n53), .Y(SUM[2]) );
  NOR2BX1 U134 ( .AN(n51), .B(n50), .Y(n53) );
  NAND2X1 U135 ( .A(n55), .B(n56), .Y(n52) );
  INVX1 U136 ( .A(n61), .Y(n58) );
  OR2X2 U137 ( .A(B[8]), .B(A[8]), .Y(n24) );
  NOR3X1 U138 ( .A(n101), .B(n102), .C(n76), .Y(n97) );
  NOR2XL U139 ( .A(A[13]), .B(B[13]), .Y(n101) );
  NAND2X2 U140 ( .A(n64), .B(n65), .Y(n62) );
  INVX4 U141 ( .A(B[12]), .Y(n127) );
  OR2X4 U142 ( .A(B[9]), .B(A[9]), .Y(n88) );
  OR2X2 U143 ( .A(B[6]), .B(A[6]), .Y(n34) );
  NAND2X1 U144 ( .A(B[8]), .B(A[8]), .Y(n22) );
  NAND2XL U145 ( .A(B[9]), .B(A[9]), .Y(n18) );
  NAND2X1 U146 ( .A(B[2]), .B(A[2]), .Y(n51) );
  OR2X2 U147 ( .A(B[7]), .B(A[7]), .Y(n141) );
  OR2X2 U148 ( .A(B[5]), .B(A[5]), .Y(n144) );
  OR2X2 U149 ( .A(B[4]), .B(A[4]), .Y(n44) );
  OR2X2 U150 ( .A(B[2]), .B(A[2]), .Y(n54) );
  NAND2X1 U151 ( .A(B[3]), .B(A[3]), .Y(n48) );
  OR2X2 U152 ( .A(B[1]), .B(A[1]), .Y(n57) );
  NAND2XL U153 ( .A(B[13]), .B(A[13]), .Y(n118) );
  NOR2X1 U154 ( .A(n67), .B(n66), .Y(n65) );
  NAND2X1 U155 ( .A(B[15]), .B(A[15]), .Y(n94) );
  XOR2X4 U156 ( .A(n62), .B(n63), .Y(SUM[16]) );
  AOI21X4 U157 ( .A0(n105), .A1(n98), .B0(n106), .Y(n104) );
  NAND2BX4 U158 ( .AN(A[13]), .B(n108), .Y(n107) );
  NAND2X4 U159 ( .A(n69), .B(n96), .Y(n103) );
  NAND2X4 U160 ( .A(n112), .B(n113), .Y(n96) );
  XOR2X4 U161 ( .A(n119), .B(n120), .Y(SUM[12]) );
  NOR3X4 U162 ( .A(n14), .B(n85), .C(n121), .Y(n120) );
  NAND2X4 U163 ( .A(n127), .B(n128), .Y(n80) );
  XOR2X4 U164 ( .A(n129), .B(n130), .Y(SUM[11]) );
  NAND2X4 U165 ( .A(n138), .B(n22), .Y(n16) );
  NAND2X4 U166 ( .A(n20), .B(n24), .Y(n138) );
endmodule


module butterfly_DW01_add_85 ( A, B, SUM );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  wire   n1, n2, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147;

  CLKINVX3 U2 ( .A(n65), .Y(n92) );
  NAND2X4 U3 ( .A(n117), .B(n118), .Y(n116) );
  NOR2X1 U4 ( .A(n59), .B(n60), .Y(n58) );
  NAND2X1 U5 ( .A(n61), .B(n62), .Y(n60) );
  NAND2X2 U6 ( .A(n85), .B(n86), .Y(n71) );
  OR2X4 U7 ( .A(B[12]), .B(A[12]), .Y(n118) );
  NAND2X2 U8 ( .A(B[12]), .B(A[12]), .Y(n68) );
  NAND2BX2 U9 ( .AN(n101), .B(n103), .Y(n78) );
  INVX8 U10 ( .A(n80), .Y(n101) );
  OAI21X2 U11 ( .A0(n112), .A1(n68), .B0(n66), .Y(n111) );
  NAND2X2 U12 ( .A(B[13]), .B(A[13]), .Y(n66) );
  NAND2X1 U13 ( .A(n9), .B(n13), .Y(n131) );
  NAND2X1 U14 ( .A(n144), .B(n145), .Y(n81) );
  INVX1 U15 ( .A(A[9]), .Y(n145) );
  INVX2 U16 ( .A(n81), .Y(n8) );
  NAND2X2 U17 ( .A(n88), .B(n66), .Y(n115) );
  OAI21XL U18 ( .A0(n26), .A1(n32), .B0(n27), .Y(n135) );
  NAND2X1 U19 ( .A(n121), .B(n122), .Y(n103) );
  OAI21XL U20 ( .A0(n8), .A1(n11), .B0(n7), .Y(n123) );
  INVX2 U21 ( .A(B[13]), .Y(n98) );
  NAND2BX2 U22 ( .AN(A[13]), .B(n98), .Y(n88) );
  OAI21X1 U23 ( .A0(n31), .A1(n84), .B0(n132), .Y(n9) );
  NAND2X1 U24 ( .A(B[10]), .B(A[10]), .Y(n122) );
  INVX1 U25 ( .A(n5), .Y(n130) );
  OAI21XL U26 ( .A0(n30), .A1(n31), .B0(n32), .Y(n28) );
  NOR2X1 U27 ( .A(A[13]), .B(B[13]), .Y(n112) );
  NOR2X1 U28 ( .A(n57), .B(n58), .Y(n56) );
  OAI21XL U29 ( .A0(n74), .A1(n72), .B0(n75), .Y(n73) );
  OAI21XL U30 ( .A0(n140), .A1(n38), .B0(n39), .Y(n82) );
  INVX3 U31 ( .A(n118), .Y(n87) );
  AND2X4 U32 ( .A(n62), .B(n61), .Y(n86) );
  OAI21X1 U33 ( .A0(n126), .A1(n127), .B0(n122), .Y(n124) );
  CLKINVX3 U34 ( .A(n79), .Y(n127) );
  NAND2X2 U35 ( .A(B[14]), .B(A[14]), .Y(n65) );
  XOR2X2 U36 ( .A(B[16]), .B(A[16]), .Y(n54) );
  NOR2X1 U37 ( .A(A[13]), .B(B[13]), .Y(n105) );
  NAND2X4 U38 ( .A(n68), .B(n116), .Y(n2) );
  OAI21XL U39 ( .A0(n101), .A1(n104), .B0(n113), .Y(n110) );
  NOR2BX2 U40 ( .AN(n102), .B(n101), .Y(n125) );
  OAI21X1 U41 ( .A0(n105), .A1(n68), .B0(n66), .Y(n93) );
  OAI21X2 U42 ( .A0(n95), .A1(n96), .B0(n97), .Y(n94) );
  INVX2 U43 ( .A(A[13]), .Y(n99) );
  AOI21X2 U44 ( .A0(n98), .A1(n99), .B0(n87), .Y(n97) );
  XOR2X2 U45 ( .A(n124), .B(n125), .Y(SUM[11]) );
  NAND2X4 U46 ( .A(n120), .B(n78), .Y(n117) );
  NOR2BX4 U47 ( .AN(n102), .B(n1), .Y(n120) );
  NOR2BX4 U48 ( .AN(n122), .B(n127), .Y(n129) );
  NOR2X2 U49 ( .A(n101), .B(n104), .Y(n1) );
  AOI21X2 U50 ( .A0(n98), .A1(n99), .B0(n87), .Y(n109) );
  NAND4X2 U51 ( .A(n13), .B(n9), .C(n81), .D(n79), .Y(n104) );
  XOR2X2 U52 ( .A(n128), .B(n129), .Y(SUM[10]) );
  NAND2X2 U53 ( .A(B[8]), .B(A[8]), .Y(n11) );
  INVX1 U54 ( .A(n18), .Y(n16) );
  OAI21X1 U55 ( .A0(n8), .A1(n130), .B0(n7), .Y(n128) );
  XNOR2X4 U56 ( .A(n115), .B(n2), .Y(SUM[13]) );
  INVX1 U57 ( .A(n82), .Y(n31) );
  NAND2BX4 U58 ( .AN(n71), .B(n73), .Y(n55) );
  NOR2XL U59 ( .A(n16), .B(n17), .Y(n15) );
  XOR2X1 U60 ( .A(n14), .B(n15), .Y(SUM[7]) );
  OAI21XL U61 ( .A0(n19), .A1(n20), .B0(n21), .Y(n14) );
  OAI21XL U62 ( .A0(n25), .A1(n26), .B0(n27), .Y(n22) );
  NAND2XL U63 ( .A(B[9]), .B(A[9]), .Y(n7) );
  NAND2BX4 U64 ( .AN(B[15]), .B(n106), .Y(n62) );
  NOR2XL U65 ( .A(n67), .B(n87), .Y(n85) );
  INVXL U66 ( .A(n84), .Y(n70) );
  INVXL U67 ( .A(A[0]), .Y(n147) );
  NAND2X2 U68 ( .A(n69), .B(n62), .Y(n89) );
  AOI21XL U69 ( .A0(n45), .A1(n142), .B0(n143), .Y(n140) );
  OAI21X2 U70 ( .A0(n133), .A1(n17), .B0(n18), .Y(n83) );
  AOI21XL U71 ( .A0(n24), .A1(n135), .B0(n136), .Y(n133) );
  XOR2X1 U72 ( .A(n9), .B(n10), .Y(SUM[8]) );
  INVXL U73 ( .A(n13), .Y(n12) );
  AOI21XL U74 ( .A0(n80), .A1(n103), .B0(n76), .Y(n113) );
  INVXL U75 ( .A(n69), .Y(n57) );
  INVXL U76 ( .A(n24), .Y(n20) );
  NOR2BXL U77 ( .AN(n27), .B(n26), .Y(n29) );
  NOR2XL U78 ( .A(n37), .B(n38), .Y(n36) );
  NOR2BXL U79 ( .AN(n47), .B(n51), .Y(n50) );
  NAND2XL U80 ( .A(n48), .B(n49), .Y(n46) );
  INVXL U81 ( .A(n52), .Y(n49) );
  INVXL U82 ( .A(n45), .Y(n41) );
  NAND2XL U83 ( .A(B[1]), .B(A[1]), .Y(n47) );
  NAND2XL U84 ( .A(B[6]), .B(A[6]), .Y(n21) );
  NAND2XL U85 ( .A(B[4]), .B(A[4]), .Y(n32) );
  NAND2XL U86 ( .A(B[5]), .B(A[5]), .Y(n27) );
  NAND2XL U87 ( .A(B[3]), .B(A[3]), .Y(n39) );
  NAND2BX1 U88 ( .AN(B[3]), .B(n141), .Y(n138) );
  OR2X2 U89 ( .A(B[7]), .B(A[7]), .Y(n134) );
  AND2X1 U90 ( .A(n52), .B(n139), .Y(SUM[0]) );
  INVX1 U91 ( .A(n83), .Y(n132) );
  AOI21X1 U92 ( .A0(n70), .A1(n82), .B0(n83), .Y(n74) );
  NOR2X1 U93 ( .A(n76), .B(n77), .Y(n75) );
  INVX1 U94 ( .A(n78), .Y(n77) );
  INVX1 U95 ( .A(n88), .Y(n67) );
  INVX1 U96 ( .A(n103), .Y(n100) );
  NOR2BX1 U97 ( .AN(n11), .B(n12), .Y(n10) );
  XOR2X1 U98 ( .A(n22), .B(n23), .Y(SUM[6]) );
  NOR2BX1 U99 ( .AN(n21), .B(n20), .Y(n23) );
  XOR2X1 U100 ( .A(n28), .B(n29), .Y(SUM[5]) );
  INVX1 U101 ( .A(n22), .Y(n19) );
  XOR2X1 U102 ( .A(n35), .B(n36), .Y(SUM[3]) );
  OAI21XL U103 ( .A0(n40), .A1(n41), .B0(n42), .Y(n35) );
  INVX1 U104 ( .A(n43), .Y(n40) );
  XOR2X1 U105 ( .A(n82), .B(n33), .Y(SUM[4]) );
  NOR2BX1 U106 ( .AN(n32), .B(n30), .Y(n33) );
  XOR2X1 U107 ( .A(n49), .B(n50), .Y(SUM[1]) );
  INVX1 U108 ( .A(n128), .Y(n126) );
  INVX1 U109 ( .A(n42), .Y(n143) );
  OAI21XL U110 ( .A0(n51), .A1(n52), .B0(n47), .Y(n142) );
  INVX1 U111 ( .A(n28), .Y(n25) );
  INVX1 U112 ( .A(n21), .Y(n136) );
  NAND4X1 U113 ( .A(n34), .B(n137), .C(n24), .D(n134), .Y(n84) );
  INVX1 U114 ( .A(n137), .Y(n26) );
  NAND4XL U115 ( .A(n79), .B(n80), .C(n81), .D(n13), .Y(n72) );
  INVXL U116 ( .A(n102), .Y(n76) );
  NOR2XL U117 ( .A(n67), .B(n68), .Y(n63) );
  NOR2X1 U118 ( .A(n63), .B(n64), .Y(n59) );
  NAND2XL U119 ( .A(n65), .B(n66), .Y(n64) );
  INVX1 U120 ( .A(n34), .Y(n30) );
  INVX1 U121 ( .A(n48), .Y(n51) );
  INVX1 U122 ( .A(n134), .Y(n17) );
  NOR2XL U123 ( .A(n101), .B(n104), .Y(n95) );
  INVX1 U124 ( .A(n39), .Y(n37) );
  XOR2X1 U125 ( .A(n43), .B(n44), .Y(SUM[2]) );
  NOR2BX1 U126 ( .AN(n42), .B(n41), .Y(n44) );
  NAND2X1 U127 ( .A(n46), .B(n47), .Y(n43) );
  OR2X4 U128 ( .A(B[8]), .B(A[8]), .Y(n13) );
  OR2X4 U129 ( .A(B[11]), .B(A[11]), .Y(n80) );
  OR2X4 U130 ( .A(A[10]), .B(B[10]), .Y(n79) );
  INVX1 U131 ( .A(B[9]), .Y(n144) );
  OR2X2 U132 ( .A(B[6]), .B(A[6]), .Y(n24) );
  NAND2BX4 U133 ( .AN(B[14]), .B(n114), .Y(n61) );
  OAI21XL U134 ( .A0(A[10]), .A1(B[10]), .B0(n123), .Y(n121) );
  NAND2X1 U135 ( .A(B[2]), .B(A[2]), .Y(n42) );
  OR2X2 U136 ( .A(B[5]), .B(A[5]), .Y(n137) );
  OR2X2 U137 ( .A(B[4]), .B(A[4]), .Y(n34) );
  OR2X2 U138 ( .A(B[2]), .B(A[2]), .Y(n45) );
  NAND2X1 U139 ( .A(B[15]), .B(A[15]), .Y(n69) );
  NAND2X1 U140 ( .A(B[7]), .B(A[7]), .Y(n18) );
  OR2X2 U141 ( .A(B[1]), .B(A[1]), .Y(n48) );
  INVX1 U142 ( .A(n138), .Y(n38) );
  INVX1 U143 ( .A(A[3]), .Y(n141) );
  NAND2X1 U144 ( .A(B[0]), .B(A[0]), .Y(n52) );
  NAND2X1 U145 ( .A(n146), .B(n147), .Y(n139) );
  INVX1 U146 ( .A(B[0]), .Y(n146) );
  NAND2X4 U147 ( .A(n55), .B(n56), .Y(n53) );
  OAI21XL U148 ( .A0(n100), .A1(n101), .B0(n102), .Y(n96) );
  INVX4 U149 ( .A(A[15]), .Y(n106) );
  INVX4 U150 ( .A(A[14]), .Y(n114) );
  NAND2X1 U151 ( .A(B[11]), .B(A[11]), .Y(n102) );
  AOI21X4 U152 ( .A0(n91), .A1(n61), .B0(n92), .Y(n90) );
  XOR2X4 U153 ( .A(n5), .B(n6), .Y(SUM[9]) );
  NOR2BX4 U154 ( .AN(n7), .B(n8), .Y(n6) );
  XOR2X4 U155 ( .A(n53), .B(n54), .Y(SUM[16]) );
  XOR2X4 U156 ( .A(n89), .B(n90), .Y(SUM[15]) );
  NAND2BX4 U157 ( .AN(n93), .B(n94), .Y(n91) );
  XOR2X4 U158 ( .A(n107), .B(n108), .Y(SUM[14]) );
  AOI21X4 U159 ( .A0(n109), .A1(n110), .B0(n111), .Y(n108) );
  NAND2X4 U160 ( .A(n61), .B(n65), .Y(n107) );
  XOR2X4 U161 ( .A(n117), .B(n119), .Y(SUM[12]) );
  NOR2BX4 U162 ( .AN(n68), .B(n87), .Y(n119) );
  NAND2X4 U163 ( .A(n131), .B(n11), .Y(n5) );
endmodule


module butterfly_DW01_sub_72 ( A, B, DIFF );
  input [16:0] A;
  input [16:0] B;
  output [16:0] DIFF;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175;

  CLKINVX2 U3 ( .A(n110), .Y(n138) );
  NAND2X2 U4 ( .A(A[9]), .B(n149), .Y(n16) );
  NAND2X2 U5 ( .A(n85), .B(n84), .Y(n4) );
  AOI2BB1X2 U6 ( .A0N(n12), .A1N(n109), .B0(n110), .Y(n108) );
  NAND2X2 U7 ( .A(n74), .B(n75), .Y(n101) );
  NOR2BX4 U8 ( .AN(n69), .B(n103), .Y(n102) );
  INVX2 U9 ( .A(n70), .Y(n97) );
  NAND2X2 U10 ( .A(n69), .B(n73), .Y(n114) );
  NAND2X1 U11 ( .A(A[14]), .B(n122), .Y(n73) );
  INVX2 U12 ( .A(A[14]), .Y(n123) );
  NAND4X1 U13 ( .A(n88), .B(n17), .C(n87), .D(n89), .Y(n110) );
  NAND2X2 U14 ( .A(A[10]), .B(n146), .Y(n136) );
  OAI21X2 U15 ( .A0(n148), .A1(n15), .B0(n16), .Y(n143) );
  NAND2X1 U16 ( .A(n75), .B(n83), .Y(n132) );
  INVX1 U17 ( .A(A[7]), .Y(n160) );
  INVX1 U18 ( .A(n17), .Y(n151) );
  INVX1 U19 ( .A(n12), .Y(n134) );
  NAND2X2 U20 ( .A(n135), .B(n136), .Y(n113) );
  XOR2X1 U21 ( .A(n35), .B(n36), .Y(DIFF[5]) );
  NOR2BX2 U22 ( .AN(n89), .B(n144), .Y(n145) );
  NAND3X2 U23 ( .A(n65), .B(n64), .C(n63), .Y(n61) );
  INVX1 U24 ( .A(n24), .Y(n30) );
  INVX1 U25 ( .A(n34), .Y(n37) );
  INVX1 U26 ( .A(B[9]), .Y(n149) );
  NAND2X1 U27 ( .A(A[8]), .B(n152), .Y(n21) );
  OAI21XL U28 ( .A0(n153), .A1(n94), .B0(n93), .Y(n17) );
  NAND4X1 U29 ( .A(n42), .B(n38), .C(n24), .D(n27), .Y(n94) );
  NAND2X1 U30 ( .A(B[8]), .B(n173), .Y(n88) );
  NAND2X2 U31 ( .A(B[9]), .B(n150), .Y(n87) );
  INVX1 U32 ( .A(A[10]), .Y(n147) );
  INVX1 U33 ( .A(n136), .Y(n144) );
  INVX2 U34 ( .A(B[11]), .Y(n109) );
  OAI2BB1X2 U35 ( .A0N(B[11]), .A1N(n134), .B0(n113), .Y(n84) );
  CLKINVX3 U36 ( .A(B[12]), .Y(n140) );
  AOI21X2 U37 ( .A0(n128), .A1(n129), .B0(n105), .Y(n126) );
  NAND2X1 U38 ( .A(n138), .B(n130), .Y(n129) );
  AOI21X2 U39 ( .A0(n131), .A1(n113), .B0(n107), .Y(n128) );
  XOR2X4 U40 ( .A(n125), .B(n124), .Y(DIFF[13]) );
  XNOR2X4 U41 ( .A(n132), .B(n8), .Y(DIFF[12]) );
  CLKINVX3 U42 ( .A(n83), .Y(n105) );
  BUFX8 U43 ( .A(A[11]), .Y(n12) );
  NAND2X2 U44 ( .A(B[10]), .B(n147), .Y(n89) );
  NAND2BX2 U45 ( .AN(n3), .B(n102), .Y(n99) );
  NOR2X1 U46 ( .A(n100), .B(n101), .Y(n3) );
  NOR2BX1 U47 ( .AN(B[11]), .B(n12), .Y(n119) );
  NAND2BXL U48 ( .AN(n12), .B(B[11]), .Y(n121) );
  OAI21X1 U49 ( .A0(n81), .A1(n82), .B0(n7), .Y(n63) );
  NAND2X2 U50 ( .A(B[7]), .B(n160), .Y(n27) );
  INVX2 U51 ( .A(B[14]), .Y(n122) );
  NAND2X4 U52 ( .A(B[14]), .B(n123), .Y(n69) );
  NAND2X2 U53 ( .A(n76), .B(n74), .Y(n125) );
  OAI21X2 U54 ( .A0(n103), .A1(n75), .B0(n74), .Y(n118) );
  NAND2XL U55 ( .A(n84), .B(n85), .Y(n82) );
  NOR2X2 U56 ( .A(n105), .B(n103), .Y(n116) );
  NOR3X1 U57 ( .A(n106), .B(n107), .C(n108), .Y(n104) );
  INVX4 U58 ( .A(n85), .Y(n107) );
  OAI21X1 U59 ( .A0(n109), .A1(n12), .B0(n138), .Y(n133) );
  NAND2BX1 U60 ( .AN(n12), .B(B[11]), .Y(n131) );
  NOR2XL U61 ( .A(n104), .B(n105), .Y(n100) );
  INVX4 U62 ( .A(A[15]), .Y(n98) );
  NOR2BX1 U63 ( .AN(n76), .B(n75), .Y(n71) );
  XOR2X4 U64 ( .A(n143), .B(n145), .Y(DIFF[10]) );
  INVX2 U65 ( .A(n4), .Y(n5) );
  AOI21XL U66 ( .A0(n89), .A1(n143), .B0(n144), .Y(n142) );
  INVX2 U67 ( .A(n13), .Y(n148) );
  AND4X4 U68 ( .A(n83), .B(n76), .C(n69), .D(n70), .Y(n7) );
  OAI21X1 U69 ( .A0(n119), .A1(n110), .B0(n120), .Y(n117) );
  NAND3X2 U70 ( .A(n137), .B(n87), .C(n89), .Y(n135) );
  NAND2X1 U71 ( .A(n27), .B(n154), .Y(n93) );
  NAND2BX2 U72 ( .AN(A[13]), .B(B[13]), .Y(n76) );
  NOR2BX4 U73 ( .AN(B[13]), .B(A[13]), .Y(n103) );
  NAND2X4 U74 ( .A(n5), .B(n133), .Y(n8) );
  BUFX3 U75 ( .A(n142), .Y(n6) );
  XOR2X1 U76 ( .A(n17), .B(n18), .Y(DIFF[8]) );
  NAND4BX2 U77 ( .AN(n80), .B(n77), .C(n78), .D(n7), .Y(n64) );
  NAND2X2 U78 ( .A(B[12]), .B(n139), .Y(n83) );
  NOR2X4 U79 ( .A(n97), .B(n11), .Y(n96) );
  NOR2BX2 U80 ( .AN(A[15]), .B(B[15]), .Y(n11) );
  OAI21X2 U81 ( .A0(n12), .A1(n109), .B0(n85), .Y(n141) );
  NOR2XL U82 ( .A(n67), .B(n68), .Y(n66) );
  NOR2BX2 U83 ( .AN(n16), .B(n15), .Y(n14) );
  NOR2BX1 U84 ( .AN(B[11]), .B(n12), .Y(n112) );
  INVXL U85 ( .A(n21), .Y(n20) );
  NOR2X1 U86 ( .A(n19), .B(n20), .Y(n18) );
  INVX2 U87 ( .A(n75), .Y(n127) );
  NOR2XL U88 ( .A(n111), .B(n112), .Y(n106) );
  INVX1 U89 ( .A(B[8]), .Y(n152) );
  NOR2XL U90 ( .A(n37), .B(n33), .Y(n36) );
  NAND2X2 U91 ( .A(n99), .B(n73), .Y(n95) );
  AOI21X1 U92 ( .A0(n45), .A1(n38), .B0(n37), .Y(n155) );
  NAND2X1 U93 ( .A(n21), .B(n16), .Y(n137) );
  INVX2 U94 ( .A(n87), .Y(n15) );
  AOI21X1 U95 ( .A0(n48), .A1(n170), .B0(n10), .Y(n166) );
  INVXL U96 ( .A(n60), .Y(n165) );
  NAND2X1 U97 ( .A(n39), .B(n40), .Y(n35) );
  NAND2X1 U98 ( .A(B[4]), .B(n163), .Y(n42) );
  INVX1 U99 ( .A(A[4]), .Y(n163) );
  NAND2X1 U100 ( .A(B[2]), .B(n172), .Y(n48) );
  XOR2X2 U101 ( .A(n25), .B(n29), .Y(DIFF[6]) );
  INVXL U102 ( .A(n113), .Y(n111) );
  AOI21XL U103 ( .A0(n77), .A1(n91), .B0(n92), .Y(n86) );
  NOR2XL U104 ( .A(n86), .B(n79), .Y(n81) );
  INVX2 U105 ( .A(n88), .Y(n19) );
  AOI21XL U106 ( .A0(n24), .A1(n25), .B0(n26), .Y(n23) );
  NAND2XL U107 ( .A(n27), .B(n28), .Y(n22) );
  INVXL U108 ( .A(n31), .Y(n26) );
  NOR2XL U109 ( .A(n44), .B(n45), .Y(n43) );
  NAND3BXL U110 ( .AN(n53), .B(n164), .C(n50), .Y(n80) );
  NAND2XL U111 ( .A(n59), .B(n60), .Y(DIFF[0]) );
  NOR2XL U112 ( .A(n58), .B(n9), .Y(n57) );
  INVXL U113 ( .A(n55), .Y(n58) );
  NOR2XL U114 ( .A(n10), .B(n53), .Y(n52) );
  NAND2BXL U115 ( .AN(n60), .B(n59), .Y(n56) );
  NAND2BX4 U116 ( .AN(B[11]), .B(n12), .Y(n85) );
  INVXL U117 ( .A(B[7]), .Y(n156) );
  INVX2 U118 ( .A(B[10]), .Y(n146) );
  NAND2XL U119 ( .A(B[5]), .B(n162), .Y(n38) );
  INVXL U120 ( .A(A[5]), .Y(n162) );
  INVXL U121 ( .A(B[6]), .Y(n157) );
  INVXL U122 ( .A(A[2]), .Y(n172) );
  INVXL U123 ( .A(B[1]), .Y(n171) );
  INVXL U124 ( .A(B[3]), .Y(n168) );
  NAND2XL U125 ( .A(B[0]), .B(n174), .Y(n60) );
  NOR2X1 U126 ( .A(n26), .B(n30), .Y(n29) );
  INVX1 U127 ( .A(n41), .Y(n153) );
  NAND2BX1 U128 ( .AN(n91), .B(n80), .Y(n41) );
  INVX1 U129 ( .A(n94), .Y(n77) );
  INVX1 U130 ( .A(n93), .Y(n92) );
  XOR2X1 U131 ( .A(n49), .B(n52), .Y(DIFF[2]) );
  XOR2X2 U132 ( .A(n22), .B(n23), .Y(DIFF[7]) );
  XOR2X1 U133 ( .A(n56), .B(n57), .Y(DIFF[1]) );
  XOR2X1 U134 ( .A(n46), .B(n47), .Y(DIFF[3]) );
  AOI21X1 U135 ( .A0(n48), .A1(n49), .B0(n10), .Y(n47) );
  NAND2X1 U136 ( .A(n50), .B(n51), .Y(n46) );
  OAI21XL U137 ( .A0(n54), .A1(n9), .B0(n55), .Y(n49) );
  INVX1 U138 ( .A(n56), .Y(n54) );
  OAI21XL U139 ( .A0(n32), .A1(n33), .B0(n34), .Y(n25) );
  INVX1 U140 ( .A(n35), .Y(n32) );
  INVX2 U141 ( .A(A[12]), .Y(n139) );
  OAI21XL U142 ( .A0(n166), .A1(n167), .B0(n51), .Y(n91) );
  INVX1 U143 ( .A(n50), .Y(n167) );
  OAI21XL U144 ( .A0(n9), .A1(n59), .B0(n55), .Y(n170) );
  OAI21X2 U145 ( .A0(n19), .A1(n151), .B0(n21), .Y(n13) );
  NOR2X1 U146 ( .A(n9), .B(n165), .Y(n164) );
  INVX1 U147 ( .A(n79), .Y(n78) );
  XOR2X1 U148 ( .A(n41), .B(n43), .Y(DIFF[4]) );
  INVX1 U149 ( .A(n42), .Y(n44) );
  INVX1 U150 ( .A(n48), .Y(n53) );
  OAI211X1 U151 ( .A0(n155), .A1(n30), .B0(n31), .C0(n28), .Y(n154) );
  NAND2X1 U152 ( .A(n41), .B(n42), .Y(n39) );
  INVX1 U153 ( .A(n38), .Y(n33) );
  INVX1 U154 ( .A(n40), .Y(n45) );
  NAND2XL U155 ( .A(n73), .B(n74), .Y(n72) );
  NOR2X1 U156 ( .A(n11), .B(n66), .Y(n65) );
  NAND2XL U157 ( .A(n69), .B(n70), .Y(n68) );
  NOR2X1 U158 ( .A(n71), .B(n72), .Y(n67) );
  NAND4XL U159 ( .A(n87), .B(n88), .C(n89), .D(n90), .Y(n79) );
  NAND2BXL U160 ( .AN(n12), .B(B[11]), .Y(n90) );
  XNOR2X2 U161 ( .A(B[16]), .B(A[16]), .Y(n62) );
  NOR2BX1 U162 ( .AN(B[1]), .B(A[1]), .Y(n9) );
  INVX1 U163 ( .A(A[9]), .Y(n150) );
  NAND2X2 U164 ( .A(B[6]), .B(n161), .Y(n24) );
  INVX1 U165 ( .A(A[6]), .Y(n161) );
  NAND2X1 U166 ( .A(B[3]), .B(n169), .Y(n50) );
  INVX1 U167 ( .A(A[3]), .Y(n169) );
  NAND2X1 U168 ( .A(A[1]), .B(n171), .Y(n55) );
  INVX1 U169 ( .A(A[8]), .Y(n173) );
  NOR2BX1 U170 ( .AN(A[2]), .B(B[2]), .Y(n10) );
  AOI21XL U171 ( .A0(n121), .A1(n113), .B0(n107), .Y(n120) );
  NAND2X1 U172 ( .A(A[3]), .B(n168), .Y(n51) );
  NAND2X1 U173 ( .A(A[4]), .B(n159), .Y(n40) );
  INVX1 U174 ( .A(B[4]), .Y(n159) );
  NAND2X1 U175 ( .A(A[5]), .B(n158), .Y(n34) );
  INVX1 U176 ( .A(B[5]), .Y(n158) );
  NAND2X1 U177 ( .A(A[7]), .B(n156), .Y(n28) );
  NAND2X1 U178 ( .A(A[6]), .B(n157), .Y(n31) );
  NAND2XL U179 ( .A(B[11]), .B(n134), .Y(n130) );
  INVX1 U180 ( .A(A[0]), .Y(n174) );
  NAND2X1 U181 ( .A(A[0]), .B(n175), .Y(n59) );
  INVX1 U182 ( .A(B[0]), .Y(n175) );
  AOI21X4 U183 ( .A0(n116), .A1(n117), .B0(n118), .Y(n115) );
  XOR2X4 U184 ( .A(n13), .B(n14), .Y(DIFF[9]) );
  XOR2X4 U185 ( .A(n61), .B(n62), .Y(DIFF[16]) );
  XOR2X4 U186 ( .A(n95), .B(n96), .Y(DIFF[15]) );
  NAND2X4 U187 ( .A(n98), .B(B[15]), .Y(n70) );
  XOR2X4 U188 ( .A(n114), .B(n115), .Y(DIFF[14]) );
  NAND2BX4 U189 ( .AN(B[13]), .B(A[13]), .Y(n74) );
  NOR2X4 U190 ( .A(n126), .B(n127), .Y(n124) );
  NAND2X4 U191 ( .A(A[12]), .B(n140), .Y(n75) );
  XOR2X4 U192 ( .A(n141), .B(n6), .Y(DIFF[11]) );
endmodule


module butterfly_DW01_add_97 ( A, B, SUM );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138;

  INVX2 U2 ( .A(n94), .Y(n62) );
  NOR2BX1 U3 ( .AN(n66), .B(n9), .Y(n90) );
  OAI21XL U4 ( .A0(n13), .A1(n123), .B0(n12), .Y(n120) );
  OAI21XL U5 ( .A0(n126), .A1(n21), .B0(n22), .Y(n88) );
  OAI21XL U6 ( .A0(n30), .A1(n35), .B0(n31), .Y(n128) );
  OR2X2 U7 ( .A(B[10]), .B(A[10]), .Y(n83) );
  OAI21XL U8 ( .A0(n62), .A1(n63), .B0(n64), .Y(n61) );
  XOR2X1 U9 ( .A(n108), .B(n4), .Y(SUM[13]) );
  XNOR2X1 U10 ( .A(n55), .B(n6), .Y(SUM[16]) );
  OR2X2 U11 ( .A(B[14]), .B(A[14]), .Y(n94) );
  AND2X2 U12 ( .A(n54), .B(n132), .Y(SUM[0]) );
  AND2X2 U13 ( .A(n64), .B(n94), .Y(n2) );
  NAND2BXL U14 ( .AN(A[11]), .B(n85), .Y(n84) );
  NAND2BXL U15 ( .AN(A[11]), .B(n85), .Y(n113) );
  NAND2BXL U16 ( .AN(A[11]), .B(n85), .Y(n116) );
  NAND2X1 U17 ( .A(B[11]), .B(A[11]), .Y(n80) );
  NOR2XL U18 ( .A(n20), .B(n21), .Y(n19) );
  NOR2BX1 U19 ( .AN(n66), .B(n58), .Y(n57) );
  NAND4X1 U20 ( .A(n37), .B(n130), .C(n28), .D(n127), .Y(n70) );
  OR2XL U21 ( .A(B[8]), .B(A[8]), .Y(n82) );
  OR2XL U22 ( .A(B[4]), .B(A[4]), .Y(n37) );
  NOR2XL U23 ( .A(n62), .B(n74), .Y(n98) );
  INVXL U24 ( .A(n26), .Y(n23) );
  INVXL U25 ( .A(n32), .Y(n29) );
  INVXL U26 ( .A(n87), .Y(n131) );
  NOR2BXL U27 ( .AN(n31), .B(n30), .Y(n33) );
  INVXL U28 ( .A(n28), .Y(n24) );
  OAI21X1 U29 ( .A0(n103), .A1(n104), .B0(n105), .Y(n102) );
  AND2X1 U30 ( .A(n106), .B(n68), .Y(n4) );
  NAND2XL U31 ( .A(B[6]), .B(A[6]), .Y(n25) );
  NAND2XL U32 ( .A(B[5]), .B(A[5]), .Y(n31) );
  NAND2XL U33 ( .A(n50), .B(n51), .Y(n48) );
  NOR2BXL U34 ( .AN(n49), .B(n53), .Y(n52) );
  INVXL U35 ( .A(n47), .Y(n43) );
  NAND3X1 U36 ( .A(n99), .B(n80), .C(n79), .Y(n110) );
  NOR2XL U37 ( .A(A[15]), .B(B[15]), .Y(n9) );
  NAND2XL U38 ( .A(B[12]), .B(A[12]), .Y(n65) );
  OR2XL U39 ( .A(B[12]), .B(A[12]), .Y(n67) );
  INVXL U40 ( .A(n99), .Y(n103) );
  NAND2XL U41 ( .A(B[7]), .B(A[7]), .Y(n22) );
  INVXL U42 ( .A(n79), .Y(n78) );
  NAND2XL U43 ( .A(B[3]), .B(A[3]), .Y(n41) );
  NOR2BXL U44 ( .AN(n134), .B(A[3]), .Y(n5) );
  NAND2XL U45 ( .A(B[1]), .B(A[1]), .Y(n49) );
  XNOR2X1 U46 ( .A(n117), .B(n118), .Y(SUM[11]) );
  NOR2BX1 U47 ( .AN(n14), .B(n17), .Y(n115) );
  OAI211XL U48 ( .A0(n13), .A1(n16), .B0(n12), .C0(n114), .Y(n112) );
  XNOR2XL U49 ( .A(B[16]), .B(A[16]), .Y(n6) );
  OAI21XL U50 ( .A0(n131), .A1(n70), .B0(n125), .Y(n14) );
  INVX1 U51 ( .A(n88), .Y(n125) );
  OAI21XL U52 ( .A0(n29), .A1(n30), .B0(n31), .Y(n26) );
  INVX1 U53 ( .A(n130), .Y(n30) );
  XOR2X1 U54 ( .A(n32), .B(n33), .Y(SUM[5]) );
  XOR2X1 U55 ( .A(n26), .B(n27), .Y(SUM[6]) );
  NOR2BX1 U56 ( .AN(n25), .B(n24), .Y(n27) );
  XOR2X1 U57 ( .A(n18), .B(n19), .Y(SUM[7]) );
  OAI21XL U58 ( .A0(n23), .A1(n24), .B0(n25), .Y(n18) );
  INVX1 U59 ( .A(n70), .Y(n86) );
  NOR3X1 U60 ( .A(n62), .B(n65), .C(n96), .Y(n60) );
  INVX1 U61 ( .A(n10), .Y(n123) );
  OAI21XL U62 ( .A0(n133), .A1(n5), .B0(n41), .Y(n87) );
  AOI21X1 U63 ( .A0(n47), .A1(n135), .B0(n136), .Y(n133) );
  INVX1 U64 ( .A(n44), .Y(n136) );
  OAI21XL U65 ( .A0(n53), .A1(n54), .B0(n49), .Y(n135) );
  OAI21XL U66 ( .A0(n34), .A1(n131), .B0(n35), .Y(n32) );
  AOI21X1 U67 ( .A0(n28), .A1(n128), .B0(n129), .Y(n126) );
  INVX1 U68 ( .A(n25), .Y(n129) );
  XOR2X2 U69 ( .A(n100), .B(n2), .Y(SUM[14]) );
  NAND2X1 U70 ( .A(n101), .B(n102), .Y(n100) );
  OR2X2 U71 ( .A(B[6]), .B(A[6]), .Y(n28) );
  INVX1 U72 ( .A(n81), .Y(n13) );
  XOR2X1 U73 ( .A(n14), .B(n15), .Y(SUM[8]) );
  NOR2BX1 U74 ( .AN(n16), .B(n17), .Y(n15) );
  XOR2X1 U75 ( .A(n110), .B(n111), .Y(SUM[12]) );
  NOR2BX1 U76 ( .AN(n65), .B(n74), .Y(n111) );
  XOR2X1 U77 ( .A(n10), .B(n11), .Y(SUM[9]) );
  NOR2BXL U78 ( .AN(n12), .B(n13), .Y(n11) );
  OR2X2 U79 ( .A(B[5]), .B(A[5]), .Y(n130) );
  NAND2X1 U80 ( .A(n124), .B(n16), .Y(n10) );
  NAND2X1 U81 ( .A(n14), .B(n82), .Y(n124) );
  INVX1 U82 ( .A(n37), .Y(n34) );
  NAND2X1 U83 ( .A(n109), .B(n65), .Y(n108) );
  INVX1 U84 ( .A(n50), .Y(n53) );
  INVX1 U85 ( .A(n127), .Y(n21) );
  INVX1 U86 ( .A(n82), .Y(n17) );
  NOR2X1 U87 ( .A(n59), .B(n9), .Y(n58) );
  NOR2X1 U88 ( .A(n60), .B(n61), .Y(n59) );
  XOR2X1 U89 ( .A(n120), .B(n121), .Y(SUM[10]) );
  NOR2BX1 U90 ( .AN(n114), .B(n122), .Y(n121) );
  INVX1 U91 ( .A(n83), .Y(n122) );
  INVX1 U92 ( .A(n67), .Y(n74) );
  NAND2X1 U93 ( .A(n110), .B(n67), .Y(n109) );
  INVXL U94 ( .A(B[11]), .Y(n85) );
  INVX1 U95 ( .A(n22), .Y(n20) );
  XOR2X1 U96 ( .A(n51), .B(n52), .Y(SUM[1]) );
  XOR2X1 U97 ( .A(n45), .B(n46), .Y(SUM[2]) );
  NOR2BX1 U98 ( .AN(n44), .B(n43), .Y(n46) );
  XOR2X1 U99 ( .A(n87), .B(n36), .Y(SUM[4]) );
  NOR2BX1 U100 ( .AN(n35), .B(n34), .Y(n36) );
  XOR2X1 U101 ( .A(n38), .B(n39), .Y(SUM[3]) );
  OAI21XL U102 ( .A0(n42), .A1(n43), .B0(n44), .Y(n38) );
  NOR2X1 U103 ( .A(n40), .B(n5), .Y(n39) );
  INVX1 U104 ( .A(n45), .Y(n42) );
  NAND2X1 U105 ( .A(n48), .B(n49), .Y(n45) );
  INVX1 U106 ( .A(n41), .Y(n40) );
  INVX1 U107 ( .A(n54), .Y(n51) );
  NAND2X1 U108 ( .A(n137), .B(n138), .Y(n132) );
  INVX1 U109 ( .A(B[0]), .Y(n137) );
  NOR2XL U110 ( .A(n65), .B(n96), .Y(n93) );
  OR2XL U111 ( .A(B[9]), .B(A[9]), .Y(n81) );
  NAND2X1 U112 ( .A(B[4]), .B(A[4]), .Y(n35) );
  NAND2XL U113 ( .A(B[8]), .B(A[8]), .Y(n16) );
  NAND2XL U114 ( .A(B[9]), .B(A[9]), .Y(n12) );
  OAI21XL U115 ( .A0(n75), .A1(n69), .B0(n76), .Y(n72) );
  AOI21X1 U116 ( .A0(n86), .A1(n87), .B0(n88), .Y(n75) );
  NAND4XL U117 ( .A(n81), .B(n82), .C(n83), .D(n84), .Y(n69) );
  NOR2X1 U118 ( .A(n77), .B(n78), .Y(n76) );
  OR2X2 U119 ( .A(B[7]), .B(A[7]), .Y(n127) );
  AND2X2 U120 ( .A(n7), .B(n67), .Y(n105) );
  OR2XL U121 ( .A(A[13]), .B(B[13]), .Y(n7) );
  OR2X2 U122 ( .A(B[2]), .B(A[2]), .Y(n47) );
  OR2X2 U123 ( .A(B[1]), .B(A[1]), .Y(n50) );
  AND2X2 U124 ( .A(n8), .B(n106), .Y(n101) );
  OR2X2 U125 ( .A(n107), .B(n65), .Y(n8) );
  OR2XL U126 ( .A(A[13]), .B(B[13]), .Y(n68) );
  NAND2XL U127 ( .A(n80), .B(n79), .Y(n104) );
  INVX1 U128 ( .A(B[3]), .Y(n134) );
  NAND3XL U129 ( .A(n99), .B(n80), .C(n79), .Y(n97) );
  INVXL U130 ( .A(n80), .Y(n77) );
  XOR2X1 U131 ( .A(n89), .B(n90), .Y(SUM[15]) );
  NAND2X1 U132 ( .A(B[0]), .B(A[0]), .Y(n54) );
  NAND2X1 U133 ( .A(B[2]), .B(A[2]), .Y(n44) );
  INVX1 U134 ( .A(A[0]), .Y(n138) );
  NAND3X1 U135 ( .A(n112), .B(n83), .C(n113), .Y(n79) );
  NAND4X1 U136 ( .A(n115), .B(n81), .C(n83), .D(n116), .Y(n99) );
  NAND2X1 U137 ( .A(n114), .B(n119), .Y(n118) );
  NAND2XL U138 ( .A(n120), .B(n83), .Y(n119) );
  NAND2X1 U139 ( .A(n56), .B(n57), .Y(n55) );
  NAND3BX1 U140 ( .AN(n71), .B(n72), .C(n73), .Y(n56) );
  NAND2XL U141 ( .A(B[13]), .B(A[13]), .Y(n106) );
  NAND2XL U142 ( .A(B[14]), .B(A[14]), .Y(n64) );
  OAI21XL U143 ( .A0(A[11]), .A1(B[11]), .B0(n80), .Y(n117) );
  NAND2X1 U144 ( .A(B[10]), .B(A[10]), .Y(n114) );
  NAND3X1 U145 ( .A(n91), .B(n64), .C(n92), .Y(n89) );
  OAI211XL U146 ( .A0(A[13]), .A1(B[13]), .B0(n97), .C0(n98), .Y(n91) );
  NAND2XL U147 ( .A(A[13]), .B(B[13]), .Y(n63) );
  NOR2XL U148 ( .A(A[13]), .B(B[13]), .Y(n107) );
  NAND2XL U149 ( .A(A[13]), .B(B[13]), .Y(n95) );
  NOR2XL U150 ( .A(A[13]), .B(B[13]), .Y(n96) );
  NOR2XL U151 ( .A(A[15]), .B(B[15]), .Y(n71) );
  NAND2XL U152 ( .A(B[15]), .B(A[15]), .Y(n66) );
  NOR3XL U153 ( .A(n62), .B(n74), .C(n96), .Y(n73) );
  AOI2BB2XL U154 ( .B0(n93), .B1(n94), .A0N(n62), .A1N(n95), .Y(n92) );
endmodule


module butterfly_DW01_sub_70 ( A, B, DIFF );
  input [16:0] A;
  input [16:0] B;
  output [16:0] DIFF;
  wire   n1, n2, n3, n4, n5, n7, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164;

  NAND2X2 U3 ( .A(n111), .B(n73), .Y(n106) );
  INVX8 U4 ( .A(n101), .Y(n64) );
  OAI2BB1X2 U5 ( .A0N(B[13]), .A1N(n118), .B0(n68), .Y(n103) );
  NAND2X2 U6 ( .A(A[14]), .B(n110), .Y(n72) );
  INVX4 U7 ( .A(B[14]), .Y(n110) );
  NAND2XL U8 ( .A(n113), .B(n114), .Y(n1) );
  NAND2X2 U9 ( .A(n2), .B(n7), .Y(n104) );
  INVX1 U10 ( .A(n1), .Y(n2) );
  NAND2BX4 U11 ( .AN(B[12]), .B(A[12]), .Y(n114) );
  NAND3X1 U12 ( .A(n113), .B(n90), .C(n91), .Y(n120) );
  NAND4X2 U13 ( .A(n128), .B(n13), .C(n93), .D(n129), .Y(n113) );
  INVXL U14 ( .A(n133), .Y(n134) );
  NAND2X2 U15 ( .A(n126), .B(n93), .Y(n135) );
  NAND2X1 U16 ( .A(n119), .B(n114), .Y(n4) );
  NAND2BX2 U17 ( .AN(A[15]), .B(B[15]), .Y(n69) );
  OAI21X1 U18 ( .A0(n130), .A1(n17), .B0(n19), .Y(n11) );
  INVX1 U19 ( .A(A[7]), .Y(n149) );
  NOR2X1 U20 ( .A(n24), .B(n28), .Y(n27) );
  NOR2BXL U21 ( .AN(n74), .B(n114), .Y(n70) );
  INVX1 U22 ( .A(B[6]), .Y(n146) );
  OAI21XL U23 ( .A0(n142), .A1(n80), .B0(n97), .Y(n15) );
  INVX1 U24 ( .A(A[13]), .Y(n118) );
  NAND2X2 U25 ( .A(n123), .B(n124), .Y(n91) );
  NAND2X1 U26 ( .A(n125), .B(n126), .Y(n123) );
  NAND3X1 U27 ( .A(n127), .B(n13), .C(n93), .Y(n125) );
  NAND2X1 U28 ( .A(n138), .B(n14), .Y(n133) );
  NAND2X1 U29 ( .A(n13), .B(n11), .Y(n138) );
  NAND2X1 U30 ( .A(A[10]), .B(n137), .Y(n126) );
  INVX1 U31 ( .A(B[10]), .Y(n137) );
  NAND2BX2 U32 ( .AN(B[11]), .B(A[11]), .Y(n90) );
  INVX1 U33 ( .A(n73), .Y(n105) );
  NOR2X1 U34 ( .A(n66), .B(n67), .Y(n65) );
  NOR2X1 U35 ( .A(n77), .B(n78), .Y(n76) );
  NOR2BX1 U36 ( .AN(B[15]), .B(A[15]), .Y(n78) );
  INVX4 U37 ( .A(n69), .Y(n100) );
  NAND2X1 U38 ( .A(n68), .B(n69), .Y(n67) );
  NAND2BX2 U39 ( .AN(B[13]), .B(A[13]), .Y(n73) );
  OAI21XL U40 ( .A0(A[13]), .A1(n115), .B0(n87), .Y(n112) );
  NAND2X2 U41 ( .A(n117), .B(n73), .Y(n116) );
  NAND2XL U42 ( .A(B[13]), .B(n118), .Y(n117) );
  NAND2X1 U43 ( .A(n120), .B(n87), .Y(n119) );
  AND2X1 U44 ( .A(n91), .B(n90), .Y(n7) );
  INVX4 U45 ( .A(A[14]), .Y(n109) );
  XNOR2X2 U46 ( .A(B[16]), .B(A[16]), .Y(n60) );
  INVX4 U47 ( .A(n68), .Y(n85) );
  NOR2X1 U48 ( .A(n64), .B(n65), .Y(n63) );
  NAND2X4 U49 ( .A(B[14]), .B(n109), .Y(n68) );
  NAND4X1 U50 ( .A(n74), .B(n75), .C(n68), .D(n76), .Y(n62) );
  NAND2BX4 U51 ( .AN(B[15]), .B(A[15]), .Y(n101) );
  BUFX3 U52 ( .A(n98), .Y(n3) );
  OAI21X1 U53 ( .A0(n102), .A1(n103), .B0(n72), .Y(n98) );
  INVX4 U54 ( .A(n87), .Y(n77) );
  NAND2BX4 U55 ( .AN(A[11]), .B(B[11]), .Y(n129) );
  NAND2BX2 U56 ( .AN(A[11]), .B(B[11]), .Y(n124) );
  XOR2X4 U57 ( .A(n59), .B(n60), .Y(DIFF[16]) );
  NAND3X2 U58 ( .A(n61), .B(n62), .C(n63), .Y(n59) );
  INVX2 U59 ( .A(n72), .Y(n108) );
  XOR2X1 U60 ( .A(n20), .B(n21), .Y(DIFF[7]) );
  NAND2X2 U61 ( .A(A[9]), .B(n139), .Y(n14) );
  AOI21XL U62 ( .A0(n22), .A1(n23), .B0(n24), .Y(n21) );
  OAI211X1 U63 ( .A0(n144), .A1(n28), .B0(n29), .C0(n26), .Y(n143) );
  NOR2X1 U64 ( .A(n17), .B(n18), .Y(n16) );
  INVX1 U65 ( .A(n19), .Y(n18) );
  NAND4X2 U66 ( .A(n40), .B(n36), .C(n22), .D(n25), .Y(n80) );
  AND2X4 U67 ( .A(n14), .B(n13), .Y(n12) );
  INVXL U68 ( .A(n39), .Y(n142) );
  XOR2X2 U69 ( .A(n23), .B(n27), .Y(DIFF[6]) );
  AOI21XL U70 ( .A0(n94), .A1(n95), .B0(n96), .Y(n88) );
  INVXL U71 ( .A(n97), .Y(n96) );
  NOR2X4 U72 ( .A(n108), .B(n85), .Y(n107) );
  XNOR2X4 U73 ( .A(n4), .B(n116), .Y(DIFF[13]) );
  INVX2 U74 ( .A(n92), .Y(n17) );
  XOR2X1 U75 ( .A(n15), .B(n16), .Y(DIFF[8]) );
  AOI21XL U76 ( .A0(n43), .A1(n36), .B0(n35), .Y(n144) );
  XNOR2X4 U77 ( .A(n5), .B(n131), .Y(DIFF[11]) );
  NAND2XL U78 ( .A(n126), .B(n132), .Y(n5) );
  NAND2XL U79 ( .A(n19), .B(n14), .Y(n127) );
  NAND2X1 U80 ( .A(n133), .B(n93), .Y(n132) );
  INVXL U81 ( .A(n40), .Y(n42) );
  NAND3BXL U82 ( .AN(n51), .B(n153), .C(n48), .Y(n81) );
  NOR2XL U83 ( .A(n9), .B(n51), .Y(n50) );
  NAND2XL U84 ( .A(n48), .B(n49), .Y(n44) );
  AOI21XL U85 ( .A0(n46), .A1(n47), .B0(n9), .Y(n45) );
  NOR2XL U86 ( .A(n56), .B(n10), .Y(n55) );
  INVXL U87 ( .A(n53), .Y(n56) );
  INVXL U88 ( .A(n46), .Y(n51) );
  NOR3X1 U89 ( .A(n79), .B(n80), .C(n81), .Y(n75) );
  NAND2BX4 U90 ( .AN(A[12]), .B(B[12]), .Y(n87) );
  NAND2X2 U91 ( .A(B[9]), .B(n162), .Y(n13) );
  NAND2X2 U92 ( .A(B[7]), .B(n149), .Y(n25) );
  NAND2XL U93 ( .A(A[7]), .B(n145), .Y(n26) );
  INVX4 U94 ( .A(A[10]), .Y(n136) );
  NAND2XL U95 ( .A(A[4]), .B(n148), .Y(n38) );
  INVXL U96 ( .A(B[4]), .Y(n148) );
  NAND2XL U97 ( .A(A[3]), .B(n157), .Y(n49) );
  INVXL U98 ( .A(B[3]), .Y(n157) );
  NAND2XL U99 ( .A(A[5]), .B(n147), .Y(n32) );
  INVXL U100 ( .A(B[5]), .Y(n147) );
  INVXL U101 ( .A(A[2]), .Y(n161) );
  NAND2XL U102 ( .A(A[0]), .B(n164), .Y(n57) );
  INVXL U103 ( .A(B[1]), .Y(n160) );
  NAND2XL U104 ( .A(B[0]), .B(n163), .Y(n58) );
  INVXL U105 ( .A(A[0]), .Y(n163) );
  INVX1 U106 ( .A(n15), .Y(n130) );
  NAND2BX1 U107 ( .AN(n95), .B(n81), .Y(n39) );
  XOR2X1 U108 ( .A(n33), .B(n34), .Y(DIFF[5]) );
  NOR2X1 U109 ( .A(n35), .B(n31), .Y(n34) );
  INVX1 U110 ( .A(n80), .Y(n94) );
  XOR2X1 U111 ( .A(n47), .B(n50), .Y(DIFF[2]) );
  XOR2X1 U112 ( .A(n39), .B(n41), .Y(DIFF[4]) );
  NOR2X1 U113 ( .A(n42), .B(n43), .Y(n41) );
  NAND2X1 U114 ( .A(n25), .B(n26), .Y(n20) );
  XOR2X1 U115 ( .A(n54), .B(n55), .Y(DIFF[1]) );
  XOR2X1 U116 ( .A(n44), .B(n45), .Y(DIFF[3]) );
  INVX2 U117 ( .A(n114), .Y(n122) );
  OAI21XL U118 ( .A0(n52), .A1(n10), .B0(n53), .Y(n47) );
  INVX1 U119 ( .A(n54), .Y(n52) );
  OAI21XL U120 ( .A0(n30), .A1(n31), .B0(n32), .Y(n23) );
  INVX1 U121 ( .A(n33), .Y(n30) );
  NAND4XL U122 ( .A(n13), .B(n92), .C(n93), .D(n124), .Y(n79) );
  OAI21XL U123 ( .A0(n155), .A1(n156), .B0(n49), .Y(n95) );
  AOI21X1 U124 ( .A0(n46), .A1(n159), .B0(n9), .Y(n155) );
  INVX1 U125 ( .A(n48), .Y(n156) );
  OAI21XL U126 ( .A0(n10), .A1(n57), .B0(n53), .Y(n159) );
  NOR2X1 U127 ( .A(n10), .B(n154), .Y(n153) );
  INVX1 U128 ( .A(n58), .Y(n154) );
  NAND2X1 U129 ( .A(n25), .B(n143), .Y(n97) );
  NAND2X1 U130 ( .A(n37), .B(n38), .Y(n33) );
  NAND2X1 U131 ( .A(n39), .B(n40), .Y(n37) );
  INVX1 U132 ( .A(n36), .Y(n31) );
  INVX1 U133 ( .A(n38), .Y(n43) );
  AND2X1 U134 ( .A(n90), .B(n91), .Y(n89) );
  INVX1 U135 ( .A(n32), .Y(n35) );
  INVX1 U136 ( .A(n29), .Y(n24) );
  INVX1 U137 ( .A(n22), .Y(n28) );
  NOR2X1 U138 ( .A(n70), .B(n71), .Y(n66) );
  NAND2X1 U139 ( .A(n57), .B(n58), .Y(DIFF[0]) );
  NAND2BX1 U140 ( .AN(n58), .B(n57), .Y(n54) );
  INVX1 U141 ( .A(A[9]), .Y(n162) );
  NOR2XL U142 ( .A(n130), .B(n17), .Y(n128) );
  NAND2X1 U143 ( .A(B[6]), .B(n150), .Y(n22) );
  INVX1 U144 ( .A(A[6]), .Y(n150) );
  NAND2X1 U145 ( .A(B[5]), .B(n151), .Y(n36) );
  INVX1 U146 ( .A(A[5]), .Y(n151) );
  NAND2X1 U147 ( .A(B[2]), .B(n161), .Y(n46) );
  NAND2X1 U148 ( .A(B[4]), .B(n152), .Y(n40) );
  INVX1 U149 ( .A(A[4]), .Y(n152) );
  NAND2X1 U150 ( .A(A[8]), .B(n140), .Y(n19) );
  INVX1 U151 ( .A(B[8]), .Y(n140) );
  INVX1 U152 ( .A(B[9]), .Y(n139) );
  NAND2X1 U153 ( .A(B[3]), .B(n158), .Y(n48) );
  INVX1 U154 ( .A(A[3]), .Y(n158) );
  NAND2X1 U155 ( .A(A[1]), .B(n160), .Y(n53) );
  NOR2BX1 U156 ( .AN(A[2]), .B(B[2]), .Y(n9) );
  NAND2X1 U157 ( .A(B[8]), .B(n141), .Y(n92) );
  INVX1 U158 ( .A(A[8]), .Y(n141) );
  NAND3X1 U159 ( .A(n82), .B(n83), .C(n84), .Y(n61) );
  OAI21XL U160 ( .A0(n88), .A1(n79), .B0(n89), .Y(n83) );
  NOR2XL U161 ( .A(n85), .B(n86), .Y(n84) );
  INVX1 U162 ( .A(B[7]), .Y(n145) );
  NAND2X1 U163 ( .A(A[6]), .B(n146), .Y(n29) );
  NOR2BX1 U164 ( .AN(B[1]), .B(A[1]), .Y(n10) );
  INVX1 U165 ( .A(B[0]), .Y(n164) );
  NAND2BX2 U166 ( .AN(n112), .B(n104), .Y(n111) );
  INVXL U167 ( .A(B[13]), .Y(n115) );
  NAND2BX1 U168 ( .AN(A[13]), .B(B[13]), .Y(n74) );
  NAND2XL U169 ( .A(n72), .B(n73), .Y(n71) );
  NAND2XL U170 ( .A(n74), .B(n87), .Y(n86) );
  AOI21XL U171 ( .A0(n104), .A1(n87), .B0(n105), .Y(n102) );
  NAND2BXL U172 ( .AN(A[15]), .B(B[15]), .Y(n82) );
  XOR2X4 U173 ( .A(n11), .B(n12), .Y(DIFF[9]) );
  XOR2X4 U174 ( .A(n3), .B(n99), .Y(DIFF[15]) );
  NOR2X4 U175 ( .A(n100), .B(n64), .Y(n99) );
  XOR2X4 U176 ( .A(n106), .B(n107), .Y(DIFF[14]) );
  XOR2X4 U177 ( .A(n120), .B(n121), .Y(DIFF[12]) );
  NOR2X4 U178 ( .A(n122), .B(n77), .Y(n121) );
  NAND2X4 U179 ( .A(n90), .B(n129), .Y(n131) );
  XOR2X4 U180 ( .A(n134), .B(n135), .Y(DIFF[10]) );
  NAND2X4 U181 ( .A(B[10]), .B(n136), .Y(n93) );
endmodule


module butterfly_DW01_sub_69 ( A, B, DIFF );
  input [16:0] A;
  input [16:0] B;
  output [16:0] DIFF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156;

  NAND2X1 U3 ( .A(A[12]), .B(n110), .Y(n87) );
  NAND2X1 U4 ( .A(A[9]), .B(n129), .Y(n12) );
  OAI21XL U5 ( .A0(n15), .A1(n119), .B0(n17), .Y(n8) );
  NAND2X1 U6 ( .A(B[10]), .B(n127), .Y(n76) );
  INVX1 U7 ( .A(n87), .Y(n108) );
  NAND2BX1 U8 ( .AN(B[13]), .B(A[13]), .Y(n86) );
  NAND3X1 U9 ( .A(n94), .B(n60), .C(n61), .Y(n102) );
  NAND2X1 U10 ( .A(A[14]), .B(n97), .Y(n83) );
  INVX1 U11 ( .A(B[14]), .Y(n97) );
  OAI2BB1X1 U12 ( .A0N(B[11]), .A1N(n112), .B0(n113), .Y(n61) );
  XNOR2X2 U13 ( .A(n95), .B(n96), .Y(DIFF[14]) );
  NOR2X1 U14 ( .A(n103), .B(n104), .Y(n99) );
  INVX1 U15 ( .A(n86), .Y(n104) );
  NAND2X1 U16 ( .A(n66), .B(n83), .Y(n96) );
  NAND2X2 U17 ( .A(B[14]), .B(n98), .Y(n66) );
  OR2XL U18 ( .A(n84), .B(n4), .Y(n1) );
  NOR2XL U19 ( .A(n79), .B(n80), .Y(n71) );
  INVXL U20 ( .A(n115), .Y(n123) );
  XOR2X2 U21 ( .A(n6), .B(n7), .Y(DIFF[16]) );
  NAND2XL U22 ( .A(B[5]), .B(n143), .Y(n140) );
  INVX1 U23 ( .A(n13), .Y(n119) );
  AOI21XL U24 ( .A0(n20), .A1(n21), .B0(n3), .Y(n19) );
  AOI21XL U25 ( .A0(n38), .A1(n39), .B0(n5), .Y(n37) );
  NOR2XL U26 ( .A(n65), .B(n78), .Y(n72) );
  INVXL U27 ( .A(n34), .Y(n132) );
  INVXL U28 ( .A(n64), .Y(n133) );
  INVXL U29 ( .A(n65), .Y(n62) );
  NAND2XL U30 ( .A(n86), .B(n87), .Y(n85) );
  INVXL U31 ( .A(n68), .Y(n84) );
  NOR2XL U32 ( .A(n92), .B(n93), .Y(n90) );
  XNOR2X1 U33 ( .A(n88), .B(n1), .Y(DIFF[15]) );
  XOR2X1 U34 ( .A(n120), .B(n121), .Y(DIFF[11]) );
  AOI21XL U35 ( .A0(n76), .A1(n122), .B0(n123), .Y(n121) );
  NAND4XL U36 ( .A(n74), .B(n75), .C(n76), .D(n77), .Y(n58) );
  XOR2X1 U37 ( .A(n8), .B(n9), .Y(DIFF[9]) );
  NOR2XL U38 ( .A(n10), .B(n11), .Y(n9) );
  XOR2X1 U39 ( .A(n122), .B(n124), .Y(DIFF[10]) );
  INVXL U40 ( .A(n76), .Y(n125) );
  NAND2XL U41 ( .A(n32), .B(n33), .Y(n29) );
  NOR2XL U42 ( .A(n15), .B(n16), .Y(n14) );
  INVXL U43 ( .A(n17), .Y(n16) );
  NAND2XL U44 ( .A(n22), .B(n23), .Y(n18) );
  NOR2XL U45 ( .A(n31), .B(n27), .Y(n30) );
  INVXL U46 ( .A(n28), .Y(n31) );
  NOR2XL U47 ( .A(n5), .B(n43), .Y(n42) );
  NOR2XL U48 ( .A(n49), .B(n45), .Y(n48) );
  INVXL U49 ( .A(n46), .Y(n49) );
  XNOR2X1 U50 ( .A(n34), .B(n2), .Y(DIFF[4]) );
  NAND2XL U51 ( .A(n35), .B(n33), .Y(n2) );
  NAND2XL U52 ( .A(n40), .B(n41), .Y(n36) );
  XOR2X1 U53 ( .A(B[16]), .B(A[16]), .Y(n7) );
  NAND2BXL U54 ( .AN(A[13]), .B(B[13]), .Y(n67) );
  NAND2XL U55 ( .A(B[12]), .B(n111), .Y(n69) );
  NAND2BXL U56 ( .AN(B[11]), .B(A[11]), .Y(n60) );
  NOR2XL U57 ( .A(n119), .B(n15), .Y(n117) );
  NOR2BXL U58 ( .AN(A[6]), .B(B[6]), .Y(n3) );
  NAND2XL U59 ( .A(B[6]), .B(n142), .Y(n20) );
  NAND2XL U60 ( .A(B[7]), .B(n141), .Y(n22) );
  INVXL U61 ( .A(B[7]), .Y(n136) );
  NAND2XL U62 ( .A(B[4]), .B(n144), .Y(n35) );
  INVXL U63 ( .A(B[5]), .Y(n138) );
  NOR2BXL U64 ( .AN(A[2]), .B(B[2]), .Y(n5) );
  NAND2XL U65 ( .A(B[2]), .B(n153), .Y(n38) );
  NAND2XL U66 ( .A(B[3]), .B(n149), .Y(n40) );
  INVXL U67 ( .A(B[1]), .Y(n151) );
  INVXL U68 ( .A(B[3]), .Y(n148) );
  NAND2XL U69 ( .A(B[1]), .B(n152), .Y(n145) );
  OAI21XL U70 ( .A0(n132), .A1(n65), .B0(n133), .Y(n13) );
  NAND4BXL U71 ( .AN(n70), .B(n71), .C(n72), .D(n73), .Y(n53) );
  INVX1 U72 ( .A(n58), .Y(n73) );
  XOR2X1 U73 ( .A(n102), .B(n109), .Y(DIFF[12]) );
  NOR2X1 U74 ( .A(n80), .B(n108), .Y(n109) );
  NAND2BX1 U75 ( .AN(n63), .B(n78), .Y(n34) );
  NAND4X1 U76 ( .A(n35), .B(n140), .C(n20), .D(n22), .Y(n65) );
  OAI21XL U77 ( .A0(n26), .A1(n27), .B0(n28), .Y(n21) );
  INVX1 U78 ( .A(n29), .Y(n26) );
  OAI21XL U79 ( .A0(n128), .A1(n11), .B0(n12), .Y(n122) );
  INVX1 U80 ( .A(n8), .Y(n128) );
  NAND2BX1 U81 ( .AN(n55), .B(n56), .Y(n54) );
  OAI21XL U82 ( .A0(n57), .A1(n58), .B0(n59), .Y(n56) );
  AOI21X1 U83 ( .A0(n62), .A1(n63), .B0(n64), .Y(n57) );
  OAI21XL U84 ( .A0(n134), .A1(n135), .B0(n23), .Y(n64) );
  AOI21X1 U85 ( .A0(n20), .A1(n137), .B0(n3), .Y(n134) );
  INVX1 U86 ( .A(n22), .Y(n135) );
  OAI21XL U87 ( .A0(n27), .A1(n33), .B0(n28), .Y(n137) );
  INVX1 U88 ( .A(n140), .Y(n27) );
  INVX1 U89 ( .A(n75), .Y(n15) );
  NOR2X1 U90 ( .A(n125), .B(n123), .Y(n124) );
  AOI21XL U91 ( .A0(n82), .A1(n83), .B0(n84), .Y(n81) );
  INVX1 U92 ( .A(n69), .Y(n80) );
  XOR2X2 U93 ( .A(n106), .B(n107), .Y(DIFF[13]) );
  NAND2X1 U94 ( .A(n67), .B(n86), .Y(n106) );
  AOI21X2 U95 ( .A0(n102), .A1(n69), .B0(n108), .Y(n107) );
  XOR2X1 U96 ( .A(n21), .B(n24), .Y(DIFF[6]) );
  NOR2X1 U97 ( .A(n3), .B(n25), .Y(n24) );
  INVX1 U98 ( .A(n20), .Y(n25) );
  NAND2XL U99 ( .A(n86), .B(n87), .Y(n93) );
  AOI31XL U100 ( .A0(n94), .A1(n60), .A2(n61), .B0(n80), .Y(n92) );
  NAND2X1 U101 ( .A(n77), .B(n60), .Y(n120) );
  XOR2X1 U102 ( .A(n18), .B(n19), .Y(DIFF[7]) );
  XOR2X1 U103 ( .A(n29), .B(n30), .Y(DIFF[5]) );
  INVX1 U104 ( .A(n74), .Y(n11) );
  AND2X2 U105 ( .A(n61), .B(n60), .Y(n59) );
  OAI21X1 U106 ( .A0(n90), .A1(n91), .B0(n83), .Y(n88) );
  NAND2X1 U107 ( .A(n67), .B(n66), .Y(n91) );
  NAND2X1 U108 ( .A(n17), .B(n12), .Y(n116) );
  NAND2X1 U109 ( .A(n99), .B(n100), .Y(n95) );
  NAND3XL U110 ( .A(n69), .B(n101), .C(n102), .Y(n100) );
  INVXL U111 ( .A(n12), .Y(n10) );
  XOR2X1 U112 ( .A(n13), .B(n14), .Y(DIFF[8]) );
  INVX1 U113 ( .A(n67), .Y(n79) );
  OAI21XL U114 ( .A0(n44), .A1(n45), .B0(n46), .Y(n39) );
  INVX1 U115 ( .A(n47), .Y(n44) );
  OAI21XL U116 ( .A0(n146), .A1(n147), .B0(n41), .Y(n63) );
  INVX1 U117 ( .A(n40), .Y(n147) );
  AOI21X1 U118 ( .A0(n38), .A1(n150), .B0(n5), .Y(n146) );
  OAI21XL U119 ( .A0(n45), .A1(n50), .B0(n46), .Y(n150) );
  NAND4X1 U120 ( .A(n40), .B(n38), .C(n51), .D(n145), .Y(n78) );
  INVX1 U121 ( .A(n145), .Y(n45) );
  INVX1 U122 ( .A(n38), .Y(n43) );
  XOR2X1 U123 ( .A(n39), .B(n42), .Y(DIFF[2]) );
  XOR2X1 U124 ( .A(n36), .B(n37), .Y(DIFF[3]) );
  XOR2X1 U125 ( .A(n47), .B(n48), .Y(DIFF[1]) );
  NAND2X1 U126 ( .A(n34), .B(n35), .Y(n32) );
  NAND2BX1 U127 ( .AN(n51), .B(n50), .Y(n47) );
  NAND2X1 U128 ( .A(n50), .B(n51), .Y(DIFF[0]) );
  INVX1 U129 ( .A(A[10]), .Y(n127) );
  INVX1 U130 ( .A(A[6]), .Y(n142) );
  INVXL U131 ( .A(B[12]), .Y(n110) );
  NAND2XL U132 ( .A(B[9]), .B(n130), .Y(n74) );
  INVX1 U133 ( .A(A[9]), .Y(n130) );
  NAND2X1 U134 ( .A(A[8]), .B(n131), .Y(n17) );
  INVXL U135 ( .A(B[8]), .Y(n131) );
  INVXL U136 ( .A(B[9]), .Y(n129) );
  INVX1 U137 ( .A(A[14]), .Y(n98) );
  NAND2X1 U138 ( .A(A[5]), .B(n138), .Y(n28) );
  NAND4X1 U139 ( .A(n117), .B(n74), .C(n76), .D(n118), .Y(n94) );
  NAND2BXL U140 ( .AN(A[11]), .B(B[11]), .Y(n118) );
  INVX1 U141 ( .A(A[7]), .Y(n141) );
  INVX1 U142 ( .A(A[12]), .Y(n111) );
  INVX1 U143 ( .A(A[11]), .Y(n112) );
  NAND2X1 U144 ( .A(n114), .B(n115), .Y(n113) );
  NAND3X1 U145 ( .A(n116), .B(n74), .C(n76), .Y(n114) );
  NAND2X1 U146 ( .A(A[7]), .B(n136), .Y(n23) );
  NAND2X1 U147 ( .A(A[10]), .B(n126), .Y(n115) );
  NAND2X1 U148 ( .A(B[15]), .B(n89), .Y(n68) );
  INVX1 U149 ( .A(A[15]), .Y(n89) );
  NAND2XL U150 ( .A(B[8]), .B(n154), .Y(n75) );
  INVX1 U151 ( .A(A[8]), .Y(n154) );
  INVX1 U152 ( .A(A[5]), .Y(n143) );
  AOI21XL U153 ( .A0(n105), .A1(B[13]), .B0(n87), .Y(n103) );
  INVX1 U154 ( .A(A[13]), .Y(n105) );
  NOR2BXL U155 ( .AN(A[15]), .B(B[15]), .Y(n4) );
  NOR2X1 U156 ( .A(n4), .B(n81), .Y(n52) );
  NAND2XL U157 ( .A(B[13]), .B(n105), .Y(n101) );
  NAND2X1 U158 ( .A(A[4]), .B(n139), .Y(n33) );
  INVX1 U159 ( .A(B[4]), .Y(n139) );
  NAND2X1 U160 ( .A(A[1]), .B(n151), .Y(n46) );
  INVX1 U161 ( .A(A[4]), .Y(n144) );
  INVX1 U162 ( .A(A[2]), .Y(n153) );
  INVX1 U163 ( .A(A[3]), .Y(n149) );
  NAND2X1 U164 ( .A(A[3]), .B(n148), .Y(n41) );
  INVX1 U165 ( .A(A[1]), .Y(n152) );
  NAND2X1 U166 ( .A(B[0]), .B(n155), .Y(n51) );
  INVX1 U167 ( .A(A[0]), .Y(n155) );
  NAND2X1 U168 ( .A(A[0]), .B(n156), .Y(n50) );
  INVX1 U169 ( .A(B[0]), .Y(n156) );
  NAND2BXL U170 ( .AN(A[11]), .B(B[11]), .Y(n77) );
  INVXL U171 ( .A(B[10]), .Y(n126) );
  NAND4XL U172 ( .A(n66), .B(n67), .C(n68), .D(n69), .Y(n55) );
  NAND2X1 U173 ( .A(n66), .B(n68), .Y(n70) );
  NAND3X1 U174 ( .A(n85), .B(n67), .C(n66), .Y(n82) );
  AND3X4 U175 ( .A(n52), .B(n53), .C(n54), .Y(n6) );
endmodule


module butterfly_DW01_add_93 ( A, B, SUM );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134;

  XNOR2X4 U2 ( .A(n86), .B(n87), .Y(n85) );
  NAND2X2 U3 ( .A(n62), .B(n57), .Y(n87) );
  NAND2BX4 U4 ( .AN(A[15]), .B(n64), .Y(n57) );
  XOR2X4 U5 ( .A(n49), .B(n50), .Y(SUM[16]) );
  XOR2X4 U6 ( .A(B[16]), .B(A[16]), .Y(n50) );
  XOR2X4 U7 ( .A(n98), .B(n99), .Y(SUM[13]) );
  NOR2BX2 U8 ( .AN(n61), .B(n65), .Y(n102) );
  NAND2X2 U9 ( .A(B[12]), .B(A[12]), .Y(n61) );
  NAND3X2 U10 ( .A(n105), .B(n77), .C(n76), .Y(n97) );
  NAND4X1 U11 ( .A(n110), .B(n80), .C(n78), .D(n79), .Y(n105) );
  NAND2X1 U12 ( .A(n97), .B(n69), .Y(n92) );
  INVX1 U13 ( .A(n59), .Y(n71) );
  NAND3X1 U14 ( .A(n106), .B(n107), .C(n79), .Y(n76) );
  NAND2BX1 U15 ( .AN(A[10]), .B(n108), .Y(n78) );
  AND2X2 U16 ( .A(n59), .B(n63), .Y(n89) );
  XOR2X2 U17 ( .A(n93), .B(n94), .Y(SUM[14]) );
  NOR2BX2 U18 ( .AN(n55), .B(n71), .Y(n94) );
  AND2X2 U19 ( .A(n48), .B(n129), .Y(SUM[0]) );
  NAND3X1 U20 ( .A(n91), .B(n61), .C(n92), .Y(n88) );
  NAND2X1 U21 ( .A(B[11]), .B(A[11]), .Y(n77) );
  INVX2 U22 ( .A(B[11]), .Y(n114) );
  XOR2X1 U23 ( .A(n97), .B(n102), .Y(SUM[12]) );
  AOI21X2 U24 ( .A0(n97), .A1(n69), .B0(n100), .Y(n99) );
  AOI21X1 U25 ( .A0(n54), .A1(n55), .B0(n56), .Y(n53) );
  INVX1 U26 ( .A(n57), .Y(n56) );
  NAND2X2 U27 ( .A(n51), .B(n52), .Y(n49) );
  NOR2BX1 U28 ( .AN(n62), .B(n53), .Y(n52) );
  NAND2X2 U29 ( .A(n103), .B(n104), .Y(n69) );
  INVX1 U30 ( .A(B[12]), .Y(n103) );
  NAND2X1 U31 ( .A(n95), .B(n91), .Y(n93) );
  AOI21X4 U32 ( .A0(n89), .A1(n88), .B0(n90), .Y(n86) );
  NAND2X2 U33 ( .A(B[13]), .B(A[13]), .Y(n91) );
  OR2X4 U34 ( .A(B[14]), .B(A[14]), .Y(n59) );
  INVX4 U35 ( .A(n85), .Y(SUM[15]) );
  INVX1 U36 ( .A(B[10]), .Y(n108) );
  NAND2X1 U37 ( .A(n96), .B(n63), .Y(n95) );
  NOR2X1 U38 ( .A(n74), .B(n75), .Y(n73) );
  INVX1 U39 ( .A(n78), .Y(n117) );
  NAND2XL U40 ( .A(B[5]), .B(A[5]), .Y(n25) );
  NAND4XL U41 ( .A(n68), .B(n69), .C(n70), .D(n57), .Y(n51) );
  OR2X4 U42 ( .A(B[9]), .B(A[9]), .Y(n80) );
  OR2X2 U43 ( .A(B[7]), .B(A[7]), .Y(n124) );
  OR2X2 U44 ( .A(B[6]), .B(A[6]), .Y(n22) );
  OR2X2 U45 ( .A(B[5]), .B(A[5]), .Y(n127) );
  NAND2X1 U46 ( .A(B[4]), .B(A[4]), .Y(n29) );
  INVXL U47 ( .A(n84), .Y(n122) );
  INVXL U48 ( .A(n83), .Y(n128) );
  INVXL U49 ( .A(n67), .Y(n82) );
  NOR2BXL U50 ( .AN(n63), .B(n71), .Y(n70) );
  INVXL U51 ( .A(n55), .Y(n90) );
  INVXL U52 ( .A(n69), .Y(n65) );
  NOR2BX1 U53 ( .AN(n8), .B(n11), .Y(n110) );
  AOI21XL U54 ( .A0(n82), .A1(n83), .B0(n84), .Y(n72) );
  XOR2X1 U55 ( .A(n118), .B(n119), .Y(SUM[10]) );
  OAI21X1 U56 ( .A0(n116), .A1(n117), .B0(n109), .Y(n111) );
  INVX1 U57 ( .A(n118), .Y(n116) );
  XOR2X1 U58 ( .A(n4), .B(n5), .Y(SUM[9]) );
  NOR2BXL U59 ( .AN(n6), .B(n7), .Y(n5) );
  INVXL U60 ( .A(n26), .Y(n23) );
  NOR2XL U61 ( .A(n14), .B(n15), .Y(n13) );
  INVXL U62 ( .A(n20), .Y(n17) );
  INVXL U63 ( .A(n81), .Y(n11) );
  AOI21XL U64 ( .A0(n41), .A1(n131), .B0(n132), .Y(n130) );
  NOR2BXL U65 ( .AN(n25), .B(n24), .Y(n27) );
  NOR2BXL U66 ( .AN(n29), .B(n28), .Y(n30) );
  NOR2BXL U67 ( .AN(n43), .B(n47), .Y(n46) );
  NAND2XL U68 ( .A(B[15]), .B(A[15]), .Y(n62) );
  INVX2 U69 ( .A(B[15]), .Y(n64) );
  NAND2XL U70 ( .A(B[10]), .B(A[10]), .Y(n109) );
  NAND2XL U71 ( .A(B[8]), .B(A[8]), .Y(n10) );
  NAND2XL U72 ( .A(B[7]), .B(A[7]), .Y(n16) );
  NAND2XL U73 ( .A(B[6]), .B(A[6]), .Y(n19) );
  NAND2XL U74 ( .A(B[1]), .B(A[1]), .Y(n43) );
  NAND2XL U75 ( .A(B[2]), .B(A[2]), .Y(n38) );
  NAND2XL U76 ( .A(B[3]), .B(A[3]), .Y(n35) );
  NOR2XL U77 ( .A(B[3]), .B(A[3]), .Y(n2) );
  OR2XL U78 ( .A(B[4]), .B(A[4]), .Y(n31) );
  OR2XL U79 ( .A(B[2]), .B(A[2]), .Y(n41) );
  OR2XL U80 ( .A(B[1]), .B(A[1]), .Y(n44) );
  INVX1 U81 ( .A(B[0]), .Y(n133) );
  OAI21XL U82 ( .A0(n128), .A1(n67), .B0(n122), .Y(n8) );
  OAI21XL U83 ( .A0(n23), .A1(n24), .B0(n25), .Y(n20) );
  OAI21XL U84 ( .A0(n7), .A1(n120), .B0(n6), .Y(n118) );
  INVX1 U85 ( .A(n4), .Y(n120) );
  OAI21XL U86 ( .A0(n123), .A1(n15), .B0(n16), .Y(n84) );
  AOI21X1 U87 ( .A0(n22), .A1(n125), .B0(n126), .Y(n123) );
  INVX1 U88 ( .A(n19), .Y(n126) );
  OAI21XL U89 ( .A0(n24), .A1(n29), .B0(n25), .Y(n125) );
  NAND4X1 U90 ( .A(n31), .B(n127), .C(n22), .D(n124), .Y(n67) );
  OAI21XL U91 ( .A0(n3), .A1(n58), .B0(n59), .Y(n54) );
  INVX1 U92 ( .A(n61), .Y(n100) );
  INVX1 U93 ( .A(n127), .Y(n24) );
  INVX1 U94 ( .A(n80), .Y(n7) );
  XOR2X1 U95 ( .A(n8), .B(n9), .Y(SUM[8]) );
  NOR2BX1 U96 ( .AN(n10), .B(n11), .Y(n9) );
  XOR2X2 U97 ( .A(n111), .B(n112), .Y(SUM[11]) );
  NOR2BX2 U98 ( .AN(n77), .B(n113), .Y(n112) );
  NOR2BX1 U99 ( .AN(n109), .B(n117), .Y(n119) );
  XOR2X1 U100 ( .A(n26), .B(n27), .Y(SUM[5]) );
  XOR2X1 U101 ( .A(n12), .B(n13), .Y(SUM[7]) );
  OAI21XL U102 ( .A0(n17), .A1(n18), .B0(n19), .Y(n12) );
  XOR2X1 U103 ( .A(n20), .B(n21), .Y(SUM[6]) );
  NOR2BX1 U104 ( .AN(n19), .B(n18), .Y(n21) );
  OAI21XL U105 ( .A0(n72), .A1(n66), .B0(n73), .Y(n68) );
  NAND4XL U106 ( .A(n78), .B(n79), .C(n80), .D(n81), .Y(n66) );
  INVX1 U107 ( .A(n22), .Y(n18) );
  INVXL U108 ( .A(n77), .Y(n74) );
  INVX1 U109 ( .A(n124), .Y(n15) );
  NAND2X1 U110 ( .A(n92), .B(n61), .Y(n96) );
  NAND2X1 U111 ( .A(n121), .B(n10), .Y(n4) );
  NAND2X1 U112 ( .A(n8), .B(n81), .Y(n121) );
  INVXL U113 ( .A(n79), .Y(n113) );
  INVXL U114 ( .A(n76), .Y(n75) );
  INVX1 U115 ( .A(n16), .Y(n14) );
  OAI21XL U116 ( .A0(n130), .A1(n2), .B0(n35), .Y(n83) );
  INVX1 U117 ( .A(n38), .Y(n132) );
  OAI21XL U118 ( .A0(n47), .A1(n48), .B0(n43), .Y(n131) );
  OAI21XL U119 ( .A0(n28), .A1(n128), .B0(n29), .Y(n26) );
  XOR2X1 U120 ( .A(n32), .B(n33), .Y(SUM[3]) );
  OAI21XL U121 ( .A0(n36), .A1(n37), .B0(n38), .Y(n32) );
  NOR2X1 U122 ( .A(n34), .B(n2), .Y(n33) );
  INVX1 U123 ( .A(n39), .Y(n36) );
  XOR2X1 U124 ( .A(n45), .B(n46), .Y(SUM[1]) );
  XOR2X1 U125 ( .A(n39), .B(n40), .Y(SUM[2]) );
  NOR2BX1 U126 ( .AN(n38), .B(n37), .Y(n40) );
  XOR2X1 U127 ( .A(n83), .B(n30), .Y(SUM[4]) );
  NAND2X1 U128 ( .A(n42), .B(n43), .Y(n39) );
  NAND2X1 U129 ( .A(n44), .B(n45), .Y(n42) );
  INVX1 U130 ( .A(n31), .Y(n28) );
  INVX1 U131 ( .A(n44), .Y(n47) );
  INVX1 U132 ( .A(n41), .Y(n37) );
  INVX1 U133 ( .A(n35), .Y(n34) );
  INVX1 U134 ( .A(n48), .Y(n45) );
  NAND2BX1 U135 ( .AN(A[10]), .B(n108), .Y(n107) );
  OAI211X1 U136 ( .A0(n7), .A1(n10), .B0(n6), .C0(n109), .Y(n106) );
  INVX1 U137 ( .A(A[11]), .Y(n115) );
  INVX1 U138 ( .A(A[12]), .Y(n104) );
  NAND2XL U139 ( .A(B[9]), .B(A[9]), .Y(n6) );
  OR2X2 U140 ( .A(B[8]), .B(A[8]), .Y(n81) );
  AND2X1 U141 ( .A(B[13]), .B(A[13]), .Y(n3) );
  NAND2X1 U142 ( .A(B[0]), .B(A[0]), .Y(n48) );
  NAND2X1 U143 ( .A(n133), .B(n134), .Y(n129) );
  INVX1 U144 ( .A(A[0]), .Y(n134) );
  NAND2X1 U145 ( .A(n63), .B(n91), .Y(n98) );
  INVX2 U146 ( .A(B[13]), .Y(n101) );
  NOR2XL U147 ( .A(n60), .B(n61), .Y(n58) );
  NOR2XL U148 ( .A(A[13]), .B(B[13]), .Y(n60) );
  NAND2X2 U149 ( .A(B[14]), .B(A[14]), .Y(n55) );
  NAND2BX4 U150 ( .AN(A[13]), .B(n101), .Y(n63) );
  NAND2X4 U151 ( .A(n114), .B(n115), .Y(n79) );
endmodule


module butterfly_DW01_sub_67 ( A, B, DIFF );
  input [16:0] A;
  input [16:0] B;
  output [16:0] DIFF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172;

  NAND2X1 U3 ( .A(n135), .B(n2), .Y(n3) );
  NAND2XL U4 ( .A(n1), .B(n136), .Y(n4) );
  NAND2X1 U5 ( .A(n3), .B(n4), .Y(DIFF[11]) );
  INVXL U6 ( .A(n135), .Y(n1) );
  INVX1 U7 ( .A(n136), .Y(n2) );
  NOR2X2 U8 ( .A(n90), .B(n137), .Y(n136) );
  NOR2BXL U9 ( .AN(A[12]), .B(B[12]), .Y(n121) );
  NOR2BXL U10 ( .AN(A[12]), .B(B[12]), .Y(n109) );
  INVX2 U11 ( .A(n72), .Y(n79) );
  INVX1 U12 ( .A(A[14]), .Y(n116) );
  INVXL U13 ( .A(A[11]), .Y(n138) );
  NOR2X1 U14 ( .A(n79), .B(n112), .Y(n102) );
  OAI21XL U15 ( .A0(n147), .A1(n17), .B0(n19), .Y(n9) );
  NAND2X1 U16 ( .A(B[9]), .B(n170), .Y(n13) );
  OAI21XL U17 ( .A0(n105), .A1(n106), .B0(n107), .Y(n103) );
  OAI21XL U18 ( .A0(n140), .A1(n141), .B0(n132), .Y(n135) );
  NOR2X2 U19 ( .A(n104), .B(n79), .Y(n114) );
  NAND2BXL U20 ( .AN(B[15]), .B(A[15]), .Y(n67) );
  NAND2BX1 U21 ( .AN(A[15]), .B(B[15]), .Y(n64) );
  NAND2BX1 U22 ( .AN(A[12]), .B(B[12]), .Y(n87) );
  NAND2X2 U23 ( .A(A[11]), .B(n139), .Y(n110) );
  AOI21X2 U24 ( .A0(n102), .A1(n103), .B0(n104), .Y(n101) );
  NAND2X2 U25 ( .A(B[14]), .B(n116), .Y(n72) );
  INVXL U26 ( .A(n110), .Y(n90) );
  INVX2 U27 ( .A(B[11]), .Y(n139) );
  INVX2 U28 ( .A(n95), .Y(n137) );
  NAND2XL U29 ( .A(B[5]), .B(n159), .Y(n36) );
  INVXL U30 ( .A(A[6]), .Y(n158) );
  INVXL U31 ( .A(B[4]), .Y(n156) );
  NOR3XL U32 ( .A(n120), .B(n6), .C(n121), .Y(n117) );
  INVXL U33 ( .A(n19), .Y(n18) );
  INVX1 U34 ( .A(n78), .Y(n86) );
  NAND2BXL U35 ( .AN(A[10]), .B(B[10]), .Y(n94) );
  NAND2X1 U36 ( .A(A[4]), .B(n156), .Y(n38) );
  NOR2XL U37 ( .A(n79), .B(n80), .Y(n77) );
  OAI21X1 U38 ( .A0(n150), .A1(n80), .B0(n99), .Y(n15) );
  INVXL U39 ( .A(n39), .Y(n150) );
  NOR2XL U40 ( .A(n82), .B(n83), .Y(n75) );
  NOR2XL U41 ( .A(n24), .B(n28), .Y(n27) );
  NOR2XL U42 ( .A(n35), .B(n31), .Y(n34) );
  INVXL U43 ( .A(n80), .Y(n96) );
  XOR2X1 U44 ( .A(n124), .B(n125), .Y(DIFF[12]) );
  INVX2 U45 ( .A(n70), .Y(n104) );
  NOR2XL U46 ( .A(n141), .B(n144), .Y(n143) );
  INVXL U47 ( .A(n132), .Y(n144) );
  AOI21XL U48 ( .A0(n96), .A1(n97), .B0(n98), .Y(n88) );
  NOR2X1 U49 ( .A(n86), .B(n81), .Y(n85) );
  XOR2X1 U50 ( .A(n122), .B(n123), .Y(DIFF[13]) );
  AOI21XL U51 ( .A0(n124), .A1(n87), .B0(n74), .Y(n123) );
  NAND2XL U52 ( .A(n71), .B(n107), .Y(n122) );
  OAI21XL U53 ( .A0(n117), .A1(n118), .B0(n107), .Y(n113) );
  NAND2X1 U54 ( .A(n145), .B(n14), .Y(n142) );
  INVXL U55 ( .A(n111), .Y(n105) );
  NOR2XL U56 ( .A(n17), .B(n18), .Y(n16) );
  NAND2XL U57 ( .A(n25), .B(n151), .Y(n99) );
  AOI21XL U58 ( .A0(n43), .A1(n36), .B0(n35), .Y(n152) );
  AOI21XL U59 ( .A0(n22), .A1(n23), .B0(n24), .Y(n21) );
  NAND2XL U60 ( .A(n25), .B(n26), .Y(n20) );
  NAND3BXL U61 ( .AN(n51), .B(n161), .C(n48), .Y(n83) );
  INVXL U62 ( .A(n46), .Y(n51) );
  NOR2XL U63 ( .A(n8), .B(n51), .Y(n50) );
  NAND2XL U64 ( .A(n48), .B(n49), .Y(n44) );
  AOI21XL U65 ( .A0(n46), .A1(n47), .B0(n8), .Y(n45) );
  AOI21XL U66 ( .A0(n64), .A1(n65), .B0(n66), .Y(n63) );
  INVXL U67 ( .A(n67), .Y(n66) );
  INVX1 U68 ( .A(n127), .Y(n74) );
  INVXL U69 ( .A(A[8]), .Y(n149) );
  NOR3X1 U70 ( .A(n108), .B(n6), .C(n109), .Y(n106) );
  INVXL U71 ( .A(A[9]), .Y(n170) );
  INVXL U72 ( .A(A[7]), .Y(n157) );
  NAND2XL U73 ( .A(A[8]), .B(n148), .Y(n19) );
  NAND2XL U74 ( .A(A[7]), .B(n153), .Y(n26) );
  NAND2XL U75 ( .A(A[6]), .B(n154), .Y(n29) );
  INVXL U76 ( .A(B[6]), .Y(n154) );
  NAND2XL U77 ( .A(A[9]), .B(n146), .Y(n14) );
  INVXL U78 ( .A(B[9]), .Y(n146) );
  AND4X1 U79 ( .A(n93), .B(n15), .C(n13), .D(n134), .Y(n5) );
  INVXL U80 ( .A(A[2]), .Y(n169) );
  INVXL U81 ( .A(A[4]), .Y(n160) );
  NAND2XL U82 ( .A(A[3]), .B(n165), .Y(n49) );
  INVXL U83 ( .A(B[3]), .Y(n165) );
  INVXL U84 ( .A(B[5]), .Y(n155) );
  NOR2BXL U85 ( .AN(B[1]), .B(A[1]), .Y(n7) );
  NAND2XL U86 ( .A(A[1]), .B(n168), .Y(n53) );
  INVXL U87 ( .A(B[1]), .Y(n168) );
  NAND2BX1 U88 ( .AN(n97), .B(n83), .Y(n39) );
  XOR2X1 U89 ( .A(n23), .B(n27), .Y(DIFF[6]) );
  XOR2X1 U90 ( .A(n33), .B(n34), .Y(DIFF[5]) );
  INVX1 U91 ( .A(n81), .Y(n76) );
  INVX1 U92 ( .A(n99), .Y(n98) );
  NAND4X1 U93 ( .A(n40), .B(n36), .C(n22), .D(n25), .Y(n80) );
  OAI21XL U94 ( .A0(n30), .A1(n31), .B0(n32), .Y(n23) );
  INVX1 U95 ( .A(n33), .Y(n30) );
  NAND3X1 U96 ( .A(n128), .B(n110), .C(n92), .Y(n124) );
  INVX1 U97 ( .A(n15), .Y(n147) );
  OAI21XL U98 ( .A0(n163), .A1(n164), .B0(n49), .Y(n97) );
  AOI21X1 U99 ( .A0(n46), .A1(n167), .B0(n8), .Y(n163) );
  INVX1 U100 ( .A(n48), .Y(n164) );
  OAI21XL U101 ( .A0(n7), .A1(n57), .B0(n53), .Y(n167) );
  OAI21XL U102 ( .A0(n88), .A1(n82), .B0(n89), .Y(n84) );
  XOR2X1 U103 ( .A(n15), .B(n16), .Y(DIFF[8]) );
  NOR2X1 U104 ( .A(n74), .B(n126), .Y(n125) );
  INVX1 U105 ( .A(n87), .Y(n126) );
  XOR2X1 U106 ( .A(n9), .B(n10), .Y(DIFF[9]) );
  NOR2X1 U107 ( .A(n11), .B(n12), .Y(n10) );
  INVX1 U108 ( .A(n14), .Y(n11) );
  INVX1 U109 ( .A(n13), .Y(n12) );
  INVX1 U110 ( .A(n142), .Y(n140) );
  XOR2X1 U111 ( .A(n142), .B(n143), .Y(DIFF[10]) );
  NAND2XL U112 ( .A(n13), .B(n9), .Y(n145) );
  NAND2X1 U113 ( .A(n37), .B(n38), .Y(n33) );
  NAND2X1 U114 ( .A(n39), .B(n40), .Y(n37) );
  OAI211X1 U115 ( .A0(n152), .A1(n28), .B0(n29), .C0(n26), .Y(n151) );
  INVX1 U116 ( .A(n36), .Y(n31) );
  INVX1 U117 ( .A(n93), .Y(n17) );
  AND2X1 U118 ( .A(n5), .B(n95), .Y(n6) );
  INVX1 U119 ( .A(n94), .Y(n141) );
  NOR2XL U120 ( .A(n90), .B(n91), .Y(n89) );
  INVXL U121 ( .A(n92), .Y(n91) );
  INVX1 U122 ( .A(n38), .Y(n43) );
  INVX1 U123 ( .A(n32), .Y(n35) );
  INVX1 U124 ( .A(n29), .Y(n24) );
  NAND2XL U125 ( .A(n92), .B(n110), .Y(n120) );
  INVX1 U126 ( .A(n22), .Y(n28) );
  NAND2X1 U127 ( .A(n19), .B(n14), .Y(n133) );
  XOR2X2 U128 ( .A(n113), .B(n114), .Y(DIFF[14]) );
  XOR2X1 U129 ( .A(n20), .B(n21), .Y(DIFF[7]) );
  OAI21XL U130 ( .A0(n52), .A1(n7), .B0(n53), .Y(n47) );
  INVX1 U131 ( .A(n54), .Y(n52) );
  NOR2X1 U132 ( .A(n7), .B(n162), .Y(n161) );
  INVX1 U133 ( .A(n58), .Y(n162) );
  XOR2X1 U134 ( .A(n47), .B(n50), .Y(DIFF[2]) );
  XOR2X1 U135 ( .A(n44), .B(n45), .Y(DIFF[3]) );
  XOR2X1 U136 ( .A(n54), .B(n55), .Y(DIFF[1]) );
  NOR2X1 U137 ( .A(n56), .B(n7), .Y(n55) );
  INVX1 U138 ( .A(n53), .Y(n56) );
  XOR2X1 U139 ( .A(n39), .B(n41), .Y(DIFF[4]) );
  NOR2X1 U140 ( .A(n42), .B(n43), .Y(n41) );
  INVX1 U141 ( .A(n40), .Y(n42) );
  NAND2X1 U142 ( .A(n57), .B(n58), .Y(DIFF[0]) );
  NAND2BX1 U143 ( .AN(n58), .B(n57), .Y(n54) );
  OAI21XL U144 ( .A0(A[13]), .A1(n119), .B0(n111), .Y(n118) );
  NAND2BXL U145 ( .AN(A[10]), .B(B[10]), .Y(n130) );
  NAND2X1 U146 ( .A(n131), .B(n132), .Y(n129) );
  NAND2XL U147 ( .A(n133), .B(n13), .Y(n131) );
  NAND2BXL U148 ( .AN(B[13]), .B(A[13]), .Y(n107) );
  NAND2XL U149 ( .A(n92), .B(n110), .Y(n108) );
  NAND2X1 U150 ( .A(B[7]), .B(n157), .Y(n25) );
  NAND2X1 U151 ( .A(B[6]), .B(n158), .Y(n22) );
  NAND2BXL U152 ( .AN(B[10]), .B(A[10]), .Y(n132) );
  INVX1 U153 ( .A(A[5]), .Y(n159) );
  NAND2X1 U154 ( .A(B[4]), .B(n160), .Y(n40) );
  INVX1 U155 ( .A(B[8]), .Y(n148) );
  NAND2X1 U156 ( .A(B[3]), .B(n166), .Y(n48) );
  INVX1 U157 ( .A(A[3]), .Y(n166) );
  OAI21XL U158 ( .A0(n68), .A1(n69), .B0(n70), .Y(n65) );
  NAND2X1 U159 ( .A(B[8]), .B(n149), .Y(n93) );
  NAND2X1 U160 ( .A(A[5]), .B(n155), .Y(n32) );
  INVX1 U161 ( .A(B[7]), .Y(n153) );
  XOR2X2 U162 ( .A(n100), .B(n101), .Y(DIFF[15]) );
  NAND2X1 U163 ( .A(n67), .B(n64), .Y(n100) );
  NAND2XL U164 ( .A(A[14]), .B(n115), .Y(n70) );
  NAND2BXL U165 ( .AN(A[10]), .B(B[10]), .Y(n134) );
  NAND2X1 U166 ( .A(B[2]), .B(n169), .Y(n46) );
  NOR2BX1 U167 ( .AN(A[2]), .B(B[2]), .Y(n8) );
  NAND2X1 U168 ( .A(B[0]), .B(n171), .Y(n58) );
  INVX1 U169 ( .A(A[0]), .Y(n171) );
  NAND2X1 U170 ( .A(A[0]), .B(n172), .Y(n57) );
  INVX1 U171 ( .A(B[0]), .Y(n172) );
  XOR2X1 U172 ( .A(n59), .B(n60), .Y(DIFF[16]) );
  XNOR2XL U173 ( .A(B[16]), .B(A[16]), .Y(n60) );
  NAND3X1 U174 ( .A(n61), .B(n62), .C(n63), .Y(n59) );
  NAND2X2 U175 ( .A(B[11]), .B(n138), .Y(n95) );
  NAND2BXL U176 ( .AN(A[15]), .B(B[15]), .Y(n78) );
  INVXL U177 ( .A(B[14]), .Y(n115) );
  NOR2XL U178 ( .A(n73), .B(n74), .Y(n68) );
  INVX1 U179 ( .A(B[13]), .Y(n119) );
  NAND2BXL U180 ( .AN(A[12]), .B(B[12]), .Y(n111) );
  NAND3X1 U181 ( .A(n84), .B(n72), .C(n85), .Y(n61) );
  NAND4X1 U182 ( .A(n75), .B(n76), .C(n77), .D(n78), .Y(n62) );
  NAND2BXL U183 ( .AN(B[12]), .B(A[12]), .Y(n127) );
  NAND4XL U184 ( .A(n13), .B(n93), .C(n94), .D(n95), .Y(n82) );
  NAND2XL U185 ( .A(n5), .B(n95), .Y(n128) );
  NAND3X2 U186 ( .A(n129), .B(n130), .C(n95), .Y(n92) );
  NAND2X1 U187 ( .A(n87), .B(n71), .Y(n81) );
  NAND2XL U188 ( .A(n71), .B(n72), .Y(n69) );
  NOR2BXL U189 ( .AN(A[13]), .B(B[13]), .Y(n73) );
  NOR2BX1 U190 ( .AN(B[13]), .B(A[13]), .Y(n112) );
  NAND2BXL U191 ( .AN(A[13]), .B(B[13]), .Y(n71) );
endmodule


module butterfly ( calc_in, rotation, calc_out );
  input [135:0] calc_in;
  input [2:0] rotation;
  output [135:0] calc_out;
  wire   N5, N6, N42, n7, n13, N306, N305, N304, N303, N302, N301, N300, N299,
         N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288,
         N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277,
         N276, N275, N274, N273, N238, N237, N236, N235, N234, N233, N232,
         N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221,
         N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210,
         N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199,
         N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188,
         N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177,
         N176, N175, N174, N173, N172, N171, N136, N135, N134, N133, N132,
         N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121,
         N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110,
         N109, N108, N107, N106, N105, N104, N103, N340, N339, N338, N337,
         N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326,
         N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315,
         N314, N313, N312, N311, N310, N309, N308, N307, N272, N271, N270,
         N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259,
         N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248,
         N247, N246, N245, N244, N243, N242, N241, N240, N239, N170, N169,
         N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158,
         N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147,
         N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N99, N98,
         N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84,
         N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70,
         N69, N102, N101, N100, n8, n9, n10, n11, n12, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55;
  wire   [16:0] temp_2_1_real;
  wire   [16:0] temp_2_2_real;
  wire   [16:0] temp_2_1_imag;
  wire   [16:0] temp_2_2_imag;
  wire   [16:0] temp_3_1_real;
  wire   [16:0] temp_3_2_real;
  wire   [16:0] temp_3_1_imag;
  wire   [16:0] temp_3_2_imag;
  wire   [16:0] temp_4_1_real;
  wire   [16:0] temp_4_2_real;
  wire   [16:0] temp_4_1_imag;
  wire   [16:0] temp_4_2_imag;
  wire   [16:0] temp_1_real;
  wire   [16:0] temp_1_imag;
  wire   [16:0] temp_2_real;
  wire   [16:0] temp_2_imag;
  wire   [16:0] temp_3_real;
  wire   [16:0] temp_3_imag;

  multi16_11 multiBRR ( .in_17bit({n43, calc_in[66:51]}), .in_8bit({1'b0, n16, 
        n35, 1'b1, n30, n40, n16, n18}), .out(temp_2_1_real) );
  multi16_10 multiBII ( .in_17bit({n42, calc_in[49:34]}), .in_8bit({n39, n9, 
        n51, 1'b0, n55, n25, n39, n9}), .out(temp_2_2_real) );
  multi16_9 multiBRI ( .in_17bit({n43, calc_in[66:51]}), .in_8bit({n39, n9, 
        n51, 1'b0, n55, n25, n39, n54}), .out(temp_2_1_imag) );
  multi16_8 multiBIR ( .in_17bit({n42, calc_in[49:34]}), .in_8bit({1'b0, n16, 
        n35, 1'b1, n30, n40, n16, n50}), .out(temp_2_2_imag) );
  multi16_7 multiCRR ( .in_17bit({n45, calc_in[100:85]}), .in_8bit({n36, n40, 
        n18, n40, n40, n24, n35, n38}), .out(temp_3_1_real) );
  multi16_6 multiCII ( .in_17bit({n44, calc_in[83:68]}), .in_8bit({n39, 1'b0, 
        n55, 1'b0, 1'b0, n55, n55, n51}), .out(temp_3_2_real) );
  multi16_5 multiCRI ( .in_17bit({n45, calc_in[100:85]}), .in_8bit({n39, 1'b0, 
        n55, 1'b0, 1'b0, n55, n55, n51}), .out(temp_3_1_imag) );
  multi16_4 multiCIR ( .in_17bit({n44, calc_in[83:68]}), .in_8bit({n36, n40, 
        n18, n40, n40, n18, n35, n38}), .out(temp_3_2_imag) );
  multi16_3 multiDRR ( .in_17bit({n47, calc_in[134:119]}), .in_8bit({n15, n38, 
        n16, n40, n50, n30, n19, n40}), .out(temp_4_1_real) );
  multi16_2 multiDII ( .in_17bit({n46, calc_in[117:102]}), .in_8bit({n26, 1'b0, 
        n41, n36, n9, n51, n53, n36}), .out(temp_4_2_real) );
  multi16_1 multiDRI ( .in_17bit({n47, calc_in[134:119]}), .in_8bit({n52, 1'b0, 
        n15, n36, n54, n51, n21, n36}), .out(temp_4_1_imag) );
  multi16_0 multiDIR ( .in_17bit({n46, calc_in[117:102]}), .in_8bit({n15, n38, 
        n16, n40, n20, n30, n19, n40}), .out(temp_4_2_imag) );
  butterfly_DW01_sub_18 sub_281 ( .A(temp_4_1_real), .B(temp_4_2_real), .DIFF(
        temp_3_real) );
  butterfly_DW01_sub_26 sub_0_root_sub_0_root_sub_300_2 ( .A({N306, N305, N304, 
        N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, 
        N291, N290}), .B({N289, N288, N287, N286, N285, N284, N283, N282, N281, 
        N280, N279, N278, N277, N276, N275, N274, N273}), .DIFF(
        calc_out[67:51]) );
  butterfly_DW01_add_36 add_0_root_sub_0_root_add_298 ( .A({N238, N237, N236, 
        N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, 
        N223, N222}), .B({N221, N220, N219, N218, N217, N216, N215, N214, N213, 
        N212, N211, N210, N209, N208, N207, N206, N205}), .SUM(
        calc_out[135:119]) );
  butterfly_DW01_add_35 add_0_root_sub_0_root_sub_296_2 ( .A({N204, N203, N202, 
        N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, 
        N189, N188}), .B({N187, N186, N185, N184, N183, N182, N181, N180, N179, 
        N178, N177, N176, N175, N174, N173, N172, N171}), .SUM(calc_out[84:68]) );
  butterfly_DW01_add_37 add_0_root_add_0_root_add_293_3 ( .A({N136, N135, N134, 
        N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, 
        N121, N120}), .B({N119, N118, N117, N116, N115, N114, N113, N112, N111, 
        N110, N109, N108, N107, N106, N105, N104, N103}), .SUM(calc_out[16:0])
         );
  butterfly_DW01_add_34 add_0_root_sub_0_root_sub_299_2 ( .A({N272, N271, N270, 
        N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, 
        N257, N256}), .B({N255, N254, N253, N252, N251, N250, N249, N248, N247, 
        N246, N245, N244, N243, N242, N241, N240, N239}), .SUM(
        calc_out[118:102]) );
  butterfly_DW01_add_38 add_0_root_add_0_root_add_292_3 ( .A({N102, N101, N100, 
        N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86}), 
        .B({N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, 
        N72, N71, N70, N69}), .SUM(calc_out[33:17]) );
  butterfly_DW01_add_48 add_1_root_sub_0_root_sub_300_2 ( .A(temp_3_imag), .B(
        temp_2_real), .SUM({N289, N288, N287, N286, N285, N284, N283, N282, 
        N281, N280, N279, N278, N277, N276, N275, N274, N273}) );
  butterfly_DW01_sub_37 sub_1_root_sub_0_root_sub_296_2 ( .A({
        temp_2_imag[16:14], n28, temp_2_imag[12:0]}), .B(temp_3_imag), .DIFF({
        N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, 
        N175, N174, N173, N172, N171}) );
  butterfly_DW01_sub_38 sub_1_root_sub_0_root_sub_299_2 ( .A(temp_1_real), .B(
        temp_3_real), .DIFF({N255, N254, N253, N252, N251, N250, N249, N248, 
        N247, N246, N245, N244, N243, N242, N241, N240, N239}) );
  butterfly_DW01_sub_39 sub_2_root_sub_0_root_sub_299_2 ( .A(calc_in[16:0]), 
        .B({temp_2_imag[16:14], n28, temp_2_imag[12:0]}), .DIFF({N272, N271, 
        N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, 
        N258, N257, N256}) );
  butterfly_DW01_add_47 add_1_root_sub_0_root_sub_295_2 ( .A(temp_1_real), .B(
        temp_3_real), .SUM({N153, N152, N151, N150, N149, N148, N147, N146, 
        N145, N144, N143, N142, N141, N140, N139, N138, N137}) );
  butterfly_DW01_add_52 add_1_root_add_0_root_add_293_3 ( .A({
        temp_1_imag[16:14], n37, temp_1_imag[12:0]}), .B(temp_3_imag), .SUM({
        N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, 
        N107, N106, N105, N104, N103}) );
  butterfly_DW01_add_50 add_2_root_sub_0_root_sub_300_2 ( .A(calc_in[33:17]), 
        .B({temp_1_imag[16:14], n37, temp_1_imag[12:0]}), .SUM({N306, N305, 
        N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, 
        N292, N291, N290}) );
  butterfly_DW01_add_51 add_2_root_add_0_root_add_293_3 ( .A(calc_in[16:0]), 
        .B({n11, temp_2_imag[15:14], n28, temp_2_imag[12:0]}), .SUM({N136, 
        N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, 
        N123, N122, N121, N120}) );
  butterfly_DW01_add_68 add_282 ( .A(temp_4_1_imag), .B(temp_4_2_imag), .SUM(
        temp_3_imag) );
  butterfly_DW01_sub_42 sub_0_root_sub_0_root_sub_295_2 ( .A({N170, N169, N168, 
        N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, 
        N155, N154}), .B({N153, N152, N151, N150, N149, N148, N147, N146, N145, 
        N144, N143, N142, N141, N140, N139, N138, N137}), .DIFF(
        calc_out[101:85]) );
  butterfly_DW01_add_72 add_0_root_sub_0_root_add_301 ( .A({N340, N339, N338, 
        N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, 
        N325, N324}), .B({N323, N322, N321, N320, N319, N318, N317, N316, N315, 
        N314, N313, N312, N311, N310, N309, N308, N307}), .SUM(calc_out[50:34]) );
  butterfly_DW01_sub_57 sub_1_root_sub_0_root_add_301 ( .A(temp_3_real), .B({
        temp_2_imag[16:14], n28, temp_2_imag[12:0]}), .DIFF({N323, N322, N321, 
        N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, 
        N308, N307}) );
  butterfly_DW01_sub_61 sub_2_root_sub_0_root_add_298 ( .A(calc_in[33:17]), 
        .B({temp_1_imag[16:14], n37, temp_1_imag[12:0]}), .DIFF({N238, N237, 
        N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, 
        N224, N223, N222}) );
  butterfly_DW01_sub_62 sub_2_root_sub_0_root_sub_296_2 ( .A(calc_in[16:0]), 
        .B({temp_1_imag[16:14], n37, temp_1_imag[12:0]}), .DIFF({N204, N203, 
        N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, 
        N190, N189, N188}) );
  butterfly_DW01_add_81 add_2_root_add_0_root_add_292_3 ( .A(calc_in[33:17]), 
        .B(temp_2_real), .SUM({N102, N101, N100, N99, N98, N97, N96, N95, N94, 
        N93, N92, N91, N90, N89, N88, N87, N86}) );
  butterfly_DW01_add_86 add_279 ( .A(temp_3_1_imag), .B(temp_3_2_imag), .SUM(
        temp_2_imag) );
  butterfly_DW01_add_85 add_276 ( .A(temp_2_1_imag), .B(temp_2_2_imag), .SUM(
        temp_1_imag) );
  butterfly_DW01_sub_72 sub_275 ( .A(temp_2_1_real), .B(temp_2_2_real), .DIFF(
        temp_1_real) );
  butterfly_DW01_add_97 add_1_root_add_0_root_add_292_3 ( .A({
        temp_1_real[16:13], n14, temp_1_real[11:0]}), .B(temp_3_real), .SUM({
        N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, 
        N71, N70, N69}) );
  butterfly_DW01_sub_70 sub_278 ( .A(temp_3_1_real), .B(temp_3_2_real), .DIFF(
        temp_2_real) );
  butterfly_DW01_sub_69 sub_2_root_sub_0_root_add_301 ( .A(calc_in[16:0]), .B(
        temp_1_real), .DIFF({N340, N339, N338, N337, N336, N335, N334, N333, 
        N332, N331, N330, N329, N328, N327, N326, N325, N324}) );
  butterfly_DW01_add_93 add_2_root_sub_0_root_sub_295_2 ( .A(calc_in[33:17]), 
        .B(temp_2_real), .SUM({N170, N169, N168, N167, N166, N165, N164, N163, 
        N162, N161, N160, N159, N158, N157, N156, N155, N154}) );
  butterfly_DW01_sub_67 sub_1_root_sub_0_root_add_298 ( .A(temp_3_imag), .B(
        temp_2_real), .DIFF({N221, N220, N219, N218, N217, N216, N215, N214, 
        N213, N212, N211, N210, N209, N208, N207, N206, N205}) );
  AND3X2 U9 ( .A(rotation[0]), .B(rotation[2]), .C(rotation[1]), .Y(n23) );
  BUFX4 U10 ( .A(calc_in[67]), .Y(n43) );
  INVX1 U11 ( .A(rotation[1]), .Y(n49) );
  INVX8 U12 ( .A(n33), .Y(n17) );
  INVX2 U13 ( .A(n7), .Y(n34) );
  INVX16 U14 ( .A(N5), .Y(n55) );
  CLKINVX8 U15 ( .A(N42), .Y(n39) );
  INVXL U16 ( .A(N5), .Y(n29) );
  BUFX12 U17 ( .A(calc_in[84]), .Y(n44) );
  BUFX8 U18 ( .A(calc_in[50]), .Y(n42) );
  INVX4 U19 ( .A(n26), .Y(n20) );
  INVX2 U20 ( .A(n54), .Y(n19) );
  INVX8 U21 ( .A(n36), .Y(n16) );
  BUFX8 U22 ( .A(n23), .Y(n36) );
  BUFX8 U23 ( .A(calc_in[118]), .Y(n46) );
  CLKINVX3 U24 ( .A(n22), .Y(n8) );
  INVX4 U25 ( .A(n8), .Y(n9) );
  BUFX8 U26 ( .A(n50), .Y(n33) );
  INVX3 U27 ( .A(n50), .Y(n26) );
  INVX3 U28 ( .A(n50), .Y(n25) );
  CLKINVX3 U29 ( .A(n13), .Y(n54) );
  INVX2 U30 ( .A(n29), .Y(n30) );
  BUFX12 U31 ( .A(temp_2_imag[13]), .Y(n28) );
  BUFX8 U32 ( .A(temp_1_imag[13]), .Y(n37) );
  INVX1 U33 ( .A(n31), .Y(n32) );
  INVX4 U34 ( .A(n34), .Y(n35) );
  INVX1 U35 ( .A(n13), .Y(n22) );
  BUFX3 U36 ( .A(calc_in[135]), .Y(n47) );
  BUFX3 U37 ( .A(calc_in[101]), .Y(n45) );
  INVX1 U38 ( .A(temp_2_imag[16]), .Y(n10) );
  CLKINVX3 U39 ( .A(n10), .Y(n11) );
  INVXL U40 ( .A(temp_1_real[12]), .Y(n12) );
  INVX1 U41 ( .A(n12), .Y(n14) );
  OAI2BB1X2 U42 ( .A0N(n49), .A1N(n48), .B0(rotation[2]), .Y(N42) );
  INVX8 U43 ( .A(n41), .Y(n40) );
  NAND3BXL U44 ( .AN(rotation[0]), .B(rotation[2]), .C(rotation[1]), .Y(n7) );
  INVX2 U45 ( .A(n50), .Y(n52) );
  NAND3BX1 U46 ( .AN(rotation[1]), .B(rotation[2]), .C(rotation[0]), .Y(n13)
         );
  XOR2X2 U47 ( .A(rotation[0]), .B(rotation[1]), .Y(n27) );
  NAND2XL U48 ( .A(rotation[1]), .B(rotation[2]), .Y(N6) );
  NAND2XL U49 ( .A(rotation[0]), .B(rotation[2]), .Y(N5) );
  INVX4 U50 ( .A(n21), .Y(n24) );
  INVX4 U51 ( .A(n24), .Y(n53) );
  CLKINVX4 U52 ( .A(n40), .Y(n15) );
  CLKINVX3 U53 ( .A(N6), .Y(n41) );
  INVX8 U54 ( .A(n17), .Y(n18) );
  AND2X4 U55 ( .A(n27), .B(n32), .Y(n21) );
  INVX4 U56 ( .A(n39), .Y(n38) );
  INVX8 U57 ( .A(n35), .Y(n51) );
  NAND2X4 U58 ( .A(n27), .B(n32), .Y(n50) );
  INVXL U59 ( .A(rotation[0]), .Y(n48) );
  INVXL U60 ( .A(rotation[2]), .Y(n31) );
endmodule


module reg1 ( clk, rst_n, data_in_2, reg_datain_flag, data_out_2 );
  input [135:0] data_in_2;
  output [135:0] data_out_2;
  input clk, rst_n, reg_datain_flag;
  wire   reg_flag_mux, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62,
         N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76,
         N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90,
         N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, N124, N125,
         N126, N127, N128, N129, N130, N131, N132, N133, N134, N135, N136,
         N137, N138, N139, N140, N141, N142, N143, N144, N145, N146, N147,
         N148, N149, N150, N151, N152, N153, N154, N155, N156, N157, N158,
         N159, N160, N161, N162, N163, N164, N165, N166, N167, N168, N169,
         N170, N171, N172, N173, N174, N175, N176, N177, N178, N179, N180,
         N181, N182, N183, N184, N185, N186, N187, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n961, n962, n964, n965, n966, n969, n971,
         n973, n974, n975, n976, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
         n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
         n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
         n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
         n1116, n8, n9, n10, n11, n96, n97, n959, n960, n963, n967, n968, n970,
         n972, n977, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173;
  wire   [1:0] counter1;
  wire   [33:0] R0;
  wire   [33:0] R1;
  wire   [33:0] R4;
  wire   [33:0] R5;
  wire   [33:0] R8;
  wire   [33:0] R9;
  wire   [33:0] R12;
  wire   [33:0] R13;
  wire   [1:0] counter2;

  CLKINVX8 U302 ( .A(rst_n), .Y(n961) );
  EDFFXL R4_reg_33_ ( .D(data_in_2[33]), .E(n969), .CK(clk), .Q(R4[33]) );
  EDFFXL R0_reg_33_ ( .D(data_in_2[33]), .E(n1117), .CK(clk), .Q(R0[33]) );
  EDFFXL R12_reg_33_ ( .D(data_in_2[33]), .E(n1131), .CK(clk), .Q(R12[33]) );
  EDFFXL R8_reg_33_ ( .D(data_in_2[33]), .E(n959), .CK(clk), .Q(R8[33]) );
  EDFFXL R4_reg_14_ ( .D(data_in_2[14]), .E(n969), .CK(clk), .Q(R4[14]) );
  EDFFXL R0_reg_14_ ( .D(data_in_2[14]), .E(n1117), .CK(clk), .Q(R0[14]) );
  EDFFXL R12_reg_14_ ( .D(data_in_2[14]), .E(n1134), .CK(clk), .Q(R12[14]) );
  EDFFXL R8_reg_14_ ( .D(data_in_2[14]), .E(n960), .CK(clk), .Q(R8[14]) );
  EDFFXL R7_reg_33_ ( .D(data_in_2[135]), .E(n1138), .CK(clk), .QN(n924) );
  EDFFXL R3_reg_33_ ( .D(data_in_2[135]), .E(n97), .CK(clk), .QN(n856) );
  EDFFXL R15_reg_33_ ( .D(data_in_2[135]), .E(n1130), .CK(clk), .QN(n788) );
  EDFFXL R11_reg_33_ ( .D(data_in_2[135]), .E(n96), .CK(clk), .QN(n686) );
  EDFFX1 R13_reg_15_ ( .D(data_in_2[49]), .E(n1134), .CK(clk), .Q(R13[15]) );
  EDFFX1 R10_reg_33_ ( .D(data_in_2[101]), .E(n96), .CK(clk), .QN(n720) );
  EDFFX1 R10_reg_32_ ( .D(data_in_2[100]), .E(n96), .CK(clk), .QN(n721) );
  EDFFX1 R10_reg_31_ ( .D(data_in_2[99]), .E(n96), .CK(clk), .QN(n722) );
  EDFFX1 R10_reg_30_ ( .D(data_in_2[98]), .E(n96), .CK(clk), .QN(n723) );
  EDFFX1 R10_reg_29_ ( .D(data_in_2[97]), .E(n96), .CK(clk), .QN(n724) );
  EDFFXL R10_reg_28_ ( .D(data_in_2[96]), .E(n96), .CK(clk), .QN(n725) );
  EDFFXL R10_reg_27_ ( .D(data_in_2[95]), .E(n96), .CK(clk), .QN(n726) );
  EDFFX1 R10_reg_22_ ( .D(data_in_2[90]), .E(n968), .CK(clk), .QN(n731) );
  EDFFX1 R10_reg_21_ ( .D(data_in_2[89]), .E(n968), .CK(clk), .QN(n732) );
  EDFFX1 R10_reg_20_ ( .D(data_in_2[88]), .E(n968), .CK(clk), .QN(n733) );
  EDFFX1 R10_reg_19_ ( .D(data_in_2[87]), .E(n968), .CK(clk), .QN(n734) );
  EDFFX1 R10_reg_18_ ( .D(data_in_2[86]), .E(n968), .CK(clk), .QN(n735) );
  EDFFX1 R10_reg_17_ ( .D(data_in_2[85]), .E(n968), .CK(clk), .QN(n736) );
  EDFFX1 R10_reg_16_ ( .D(data_in_2[84]), .E(n968), .CK(clk), .QN(n737) );
  EDFFX1 R10_reg_15_ ( .D(data_in_2[83]), .E(n968), .CK(clk), .QN(n738) );
  EDFFX1 R10_reg_14_ ( .D(data_in_2[82]), .E(n968), .CK(clk), .QN(n739) );
  EDFFX1 R10_reg_13_ ( .D(data_in_2[81]), .E(n968), .CK(clk), .QN(n740) );
  EDFFX1 R10_reg_12_ ( .D(data_in_2[80]), .E(n968), .CK(clk), .QN(n741) );
  EDFFX1 R10_reg_5_ ( .D(data_in_2[73]), .E(n970), .CK(clk), .QN(n748) );
  EDFFX1 R10_reg_4_ ( .D(data_in_2[72]), .E(n970), .CK(clk), .QN(n749) );
  EDFFX1 R10_reg_3_ ( .D(data_in_2[71]), .E(n970), .CK(clk), .QN(n750) );
  EDFFX1 R10_reg_2_ ( .D(data_in_2[70]), .E(n970), .CK(clk), .QN(n751) );
  EDFFX1 R10_reg_1_ ( .D(data_in_2[69]), .E(n970), .CK(clk), .QN(n752) );
  EDFFX1 R10_reg_0_ ( .D(data_in_2[68]), .E(n970), .CK(clk), .QN(n753) );
  EDFFX1 R14_reg_33_ ( .D(data_in_2[101]), .E(n1133), .CK(clk), .QN(n754) );
  EDFFX1 R14_reg_32_ ( .D(data_in_2[100]), .E(n1133), .CK(clk), .QN(n755) );
  EDFFX1 R14_reg_31_ ( .D(data_in_2[99]), .E(n1133), .CK(clk), .QN(n756) );
  EDFFX1 R14_reg_30_ ( .D(data_in_2[98]), .E(n1132), .CK(clk), .QN(n757) );
  EDFFX1 R14_reg_29_ ( .D(data_in_2[97]), .E(n1132), .CK(clk), .QN(n758) );
  EDFFXL R14_reg_28_ ( .D(data_in_2[96]), .E(n1132), .CK(clk), .QN(n759) );
  EDFFXL R14_reg_27_ ( .D(data_in_2[95]), .E(n1132), .CK(clk), .QN(n760) );
  EDFFX1 R14_reg_26_ ( .D(data_in_2[94]), .E(n1132), .CK(clk), .QN(n761) );
  EDFFX1 R14_reg_25_ ( .D(data_in_2[93]), .E(n1132), .CK(clk), .QN(n762) );
  EDFFX1 R14_reg_24_ ( .D(data_in_2[92]), .E(n1132), .CK(clk), .QN(n763) );
  EDFFX1 R14_reg_23_ ( .D(data_in_2[91]), .E(n1132), .CK(clk), .QN(n764) );
  EDFFX1 R14_reg_22_ ( .D(data_in_2[90]), .E(n1132), .CK(clk), .QN(n765) );
  EDFFX1 R14_reg_21_ ( .D(data_in_2[89]), .E(n1132), .CK(clk), .QN(n766) );
  EDFFX1 R14_reg_20_ ( .D(data_in_2[88]), .E(n1132), .CK(clk), .QN(n767) );
  EDFFX1 R14_reg_19_ ( .D(data_in_2[87]), .E(n1132), .CK(clk), .QN(n768) );
  EDFFX1 R14_reg_18_ ( .D(data_in_2[86]), .E(n1132), .CK(clk), .QN(n769) );
  EDFFX1 R14_reg_17_ ( .D(data_in_2[85]), .E(n1131), .CK(clk), .QN(n770) );
  EDFFX1 R14_reg_16_ ( .D(data_in_2[84]), .E(n1131), .CK(clk), .QN(n771) );
  EDFFX1 R14_reg_15_ ( .D(data_in_2[83]), .E(n1131), .CK(clk), .QN(n772) );
  EDFFX1 R14_reg_14_ ( .D(data_in_2[82]), .E(n1131), .CK(clk), .QN(n773) );
  EDFFX1 R14_reg_13_ ( .D(data_in_2[81]), .E(n1131), .CK(clk), .QN(n774) );
  EDFFX1 R14_reg_12_ ( .D(data_in_2[80]), .E(n1131), .CK(clk), .QN(n775) );
  EDFFX1 R14_reg_11_ ( .D(data_in_2[79]), .E(n1131), .CK(clk), .QN(n776) );
  EDFFX1 R14_reg_10_ ( .D(data_in_2[78]), .E(n1131), .CK(clk), .QN(n777) );
  EDFFX1 R14_reg_9_ ( .D(data_in_2[77]), .E(n1131), .CK(clk), .QN(n778) );
  EDFFX1 R14_reg_8_ ( .D(data_in_2[76]), .E(n1131), .CK(clk), .QN(n779) );
  EDFFX1 R14_reg_7_ ( .D(data_in_2[75]), .E(n1131), .CK(clk), .QN(n780) );
  EDFFX1 R14_reg_6_ ( .D(data_in_2[74]), .E(n1131), .CK(clk), .QN(n781) );
  EDFFX1 R14_reg_5_ ( .D(data_in_2[73]), .E(n1131), .CK(clk), .QN(n782) );
  EDFFX1 R14_reg_4_ ( .D(data_in_2[72]), .E(n1130), .CK(clk), .QN(n783) );
  EDFFX1 R14_reg_3_ ( .D(data_in_2[71]), .E(n1130), .CK(clk), .QN(n784) );
  EDFFX1 R14_reg_2_ ( .D(data_in_2[70]), .E(n1130), .CK(clk), .QN(n785) );
  EDFFX1 R14_reg_1_ ( .D(data_in_2[69]), .E(n1130), .CK(clk), .QN(n786) );
  EDFFX1 R14_reg_0_ ( .D(data_in_2[68]), .E(n1130), .CK(clk), .QN(n787) );
  EDFFX1 R2_reg_33_ ( .D(data_in_2[101]), .E(n97), .CK(clk), .QN(n822) );
  EDFFX1 R2_reg_32_ ( .D(data_in_2[100]), .E(n97), .CK(clk), .QN(n823) );
  EDFFX1 R2_reg_31_ ( .D(data_in_2[99]), .E(n97), .CK(clk), .QN(n824) );
  EDFFX1 R2_reg_30_ ( .D(data_in_2[98]), .E(n97), .CK(clk), .QN(n825) );
  EDFFX1 R2_reg_29_ ( .D(data_in_2[97]), .E(n97), .CK(clk), .QN(n826) );
  EDFFXL R2_reg_28_ ( .D(data_in_2[96]), .E(n97), .CK(clk), .QN(n827) );
  EDFFXL R2_reg_27_ ( .D(data_in_2[95]), .E(n97), .CK(clk), .QN(n828) );
  EDFFX1 R2_reg_26_ ( .D(data_in_2[94]), .E(n97), .CK(clk), .QN(n829) );
  EDFFX1 R2_reg_25_ ( .D(data_in_2[93]), .E(n97), .CK(clk), .QN(n830) );
  EDFFX1 R2_reg_24_ ( .D(data_in_2[92]), .E(n97), .CK(clk), .QN(n831) );
  EDFFX1 R2_reg_23_ ( .D(data_in_2[91]), .E(n97), .CK(clk), .QN(n832) );
  EDFFX1 R2_reg_22_ ( .D(data_in_2[90]), .E(n97), .CK(clk), .QN(n833) );
  EDFFX1 R2_reg_21_ ( .D(data_in_2[89]), .E(n97), .CK(clk), .QN(n834) );
  EDFFX1 R2_reg_20_ ( .D(data_in_2[88]), .E(n97), .CK(clk), .QN(n835) );
  EDFFX1 R2_reg_19_ ( .D(data_in_2[87]), .E(n97), .CK(clk), .QN(n836) );
  EDFFX1 R2_reg_18_ ( .D(data_in_2[86]), .E(n97), .CK(clk), .QN(n837) );
  EDFFX1 R2_reg_17_ ( .D(data_in_2[85]), .E(n97), .CK(clk), .QN(n838) );
  EDFFX1 R2_reg_16_ ( .D(data_in_2[84]), .E(n97), .CK(clk), .QN(n839) );
  EDFFX1 R2_reg_15_ ( .D(data_in_2[83]), .E(n97), .CK(clk), .QN(n840) );
  EDFFX1 R2_reg_14_ ( .D(data_in_2[82]), .E(n97), .CK(clk), .QN(n841) );
  EDFFX1 R2_reg_13_ ( .D(data_in_2[81]), .E(n97), .CK(clk), .QN(n842) );
  EDFFX1 R2_reg_12_ ( .D(data_in_2[80]), .E(n97), .CK(clk), .QN(n843) );
  EDFFX1 R2_reg_11_ ( .D(data_in_2[79]), .E(n97), .CK(clk), .QN(n844) );
  EDFFX1 R2_reg_10_ ( .D(data_in_2[78]), .E(n97), .CK(clk), .QN(n845) );
  EDFFX1 R2_reg_9_ ( .D(data_in_2[77]), .E(n97), .CK(clk), .QN(n846) );
  EDFFX1 R2_reg_8_ ( .D(data_in_2[76]), .E(n97), .CK(clk), .QN(n847) );
  EDFFX1 R2_reg_7_ ( .D(data_in_2[75]), .E(n97), .CK(clk), .QN(n848) );
  EDFFX1 R2_reg_6_ ( .D(data_in_2[74]), .E(n97), .CK(clk), .QN(n849) );
  EDFFX1 R2_reg_5_ ( .D(data_in_2[73]), .E(n97), .CK(clk), .QN(n850) );
  EDFFX1 R2_reg_4_ ( .D(data_in_2[72]), .E(n97), .CK(clk), .QN(n851) );
  EDFFX1 R2_reg_3_ ( .D(data_in_2[71]), .E(n97), .CK(clk), .QN(n852) );
  EDFFX1 R2_reg_2_ ( .D(data_in_2[70]), .E(n97), .CK(clk), .QN(n853) );
  EDFFX1 R2_reg_1_ ( .D(data_in_2[69]), .E(n97), .CK(clk), .QN(n854) );
  EDFFX1 R2_reg_0_ ( .D(data_in_2[68]), .E(n97), .CK(clk), .QN(n855) );
  EDFFXL R6_reg_33_ ( .D(data_in_2[101]), .E(n1137), .CK(clk), .QN(n890) );
  EDFFXL R6_reg_32_ ( .D(data_in_2[100]), .E(n1137), .CK(clk), .QN(n891) );
  EDFFXL R6_reg_31_ ( .D(data_in_2[99]), .E(n1137), .CK(clk), .QN(n892) );
  EDFFXL R6_reg_30_ ( .D(data_in_2[98]), .E(n1137), .CK(clk), .QN(n893) );
  EDFFXL R6_reg_29_ ( .D(data_in_2[97]), .E(n1137), .CK(clk), .QN(n894) );
  EDFFXL R6_reg_28_ ( .D(data_in_2[96]), .E(n1137), .CK(clk), .QN(n895) );
  EDFFXL R6_reg_27_ ( .D(data_in_2[95]), .E(n1137), .CK(clk), .QN(n896) );
  EDFFX1 R6_reg_26_ ( .D(data_in_2[94]), .E(n1137), .CK(clk), .QN(n897) );
  EDFFX1 R6_reg_25_ ( .D(data_in_2[93]), .E(n1137), .CK(clk), .QN(n898) );
  EDFFX1 R6_reg_24_ ( .D(data_in_2[92]), .E(n1137), .CK(clk), .QN(n899) );
  EDFFX1 R6_reg_23_ ( .D(data_in_2[91]), .E(n1137), .CK(clk), .QN(n900) );
  EDFFX1 R6_reg_22_ ( .D(data_in_2[90]), .E(n1137), .CK(clk), .QN(n901) );
  EDFFX1 R6_reg_21_ ( .D(data_in_2[89]), .E(n1137), .CK(clk), .QN(n902) );
  EDFFX1 R6_reg_20_ ( .D(data_in_2[88]), .E(n1137), .CK(clk), .QN(n903) );
  EDFFX1 R6_reg_19_ ( .D(data_in_2[87]), .E(n1137), .CK(clk), .QN(n904) );
  EDFFX1 R6_reg_18_ ( .D(data_in_2[86]), .E(n1137), .CK(clk), .QN(n905) );
  EDFFX1 R6_reg_17_ ( .D(data_in_2[85]), .E(n1137), .CK(clk), .QN(n906) );
  EDFFXL R6_reg_16_ ( .D(data_in_2[84]), .E(n1137), .CK(clk), .QN(n907) );
  EDFFXL R6_reg_15_ ( .D(data_in_2[83]), .E(n1137), .CK(clk), .QN(n908) );
  EDFFXL R6_reg_14_ ( .D(data_in_2[82]), .E(n1137), .CK(clk), .QN(n909) );
  EDFFXL R6_reg_13_ ( .D(data_in_2[81]), .E(n1137), .CK(clk), .QN(n910) );
  EDFFXL R6_reg_12_ ( .D(data_in_2[80]), .E(n1137), .CK(clk), .QN(n911) );
  EDFFX1 R6_reg_11_ ( .D(data_in_2[79]), .E(n1137), .CK(clk), .QN(n912) );
  EDFFX1 R6_reg_10_ ( .D(data_in_2[78]), .E(n1137), .CK(clk), .QN(n913) );
  EDFFX1 R6_reg_9_ ( .D(data_in_2[77]), .E(n1137), .CK(clk), .QN(n914) );
  EDFFX1 R6_reg_8_ ( .D(data_in_2[76]), .E(n1137), .CK(clk), .QN(n915) );
  EDFFX1 R6_reg_7_ ( .D(data_in_2[75]), .E(n1137), .CK(clk), .QN(n916) );
  EDFFX1 R6_reg_6_ ( .D(data_in_2[74]), .E(n1137), .CK(clk), .QN(n917) );
  EDFFX1 R6_reg_5_ ( .D(data_in_2[73]), .E(n1137), .CK(clk), .QN(n918) );
  EDFFX1 R6_reg_4_ ( .D(data_in_2[72]), .E(n1137), .CK(clk), .QN(n919) );
  EDFFX1 R6_reg_3_ ( .D(data_in_2[71]), .E(n1137), .CK(clk), .QN(n920) );
  EDFFX1 R6_reg_2_ ( .D(data_in_2[70]), .E(n1137), .CK(clk), .QN(n921) );
  EDFFX1 R6_reg_1_ ( .D(data_in_2[69]), .E(n1137), .CK(clk), .QN(n922) );
  EDFFX1 R6_reg_0_ ( .D(data_in_2[68]), .E(n1137), .CK(clk), .QN(n923) );
  EDFFX1 R11_reg_32_ ( .D(data_in_2[134]), .E(n96), .CK(clk), .QN(n687) );
  EDFFX1 R11_reg_31_ ( .D(data_in_2[133]), .E(n96), .CK(clk), .QN(n688) );
  EDFFX1 R11_reg_30_ ( .D(data_in_2[132]), .E(n96), .CK(clk), .QN(n689) );
  EDFFX1 R11_reg_29_ ( .D(data_in_2[131]), .E(n96), .CK(clk), .QN(n690) );
  EDFFX1 R11_reg_22_ ( .D(data_in_2[124]), .E(n963), .CK(clk), .QN(n697) );
  EDFFX1 R11_reg_21_ ( .D(data_in_2[123]), .E(n963), .CK(clk), .QN(n698) );
  EDFFX1 R11_reg_20_ ( .D(data_in_2[122]), .E(n963), .CK(clk), .QN(n699) );
  EDFFX1 R11_reg_19_ ( .D(data_in_2[121]), .E(n963), .CK(clk), .QN(n700) );
  EDFFX1 R11_reg_18_ ( .D(data_in_2[120]), .E(n963), .CK(clk), .QN(n701) );
  EDFFX1 R11_reg_17_ ( .D(data_in_2[119]), .E(n963), .CK(clk), .QN(n702) );
  EDFFX1 R11_reg_16_ ( .D(data_in_2[118]), .E(n963), .CK(clk), .QN(n703) );
  EDFFX1 R11_reg_15_ ( .D(data_in_2[117]), .E(n967), .CK(clk), .QN(n704) );
  EDFFX1 R11_reg_14_ ( .D(data_in_2[116]), .E(n967), .CK(clk), .QN(n705) );
  EDFFX1 R11_reg_13_ ( .D(data_in_2[115]), .E(n967), .CK(clk), .QN(n706) );
  EDFFX1 R11_reg_12_ ( .D(data_in_2[114]), .E(n967), .CK(clk), .QN(n707) );
  EDFFX1 R11_reg_5_ ( .D(data_in_2[107]), .E(n967), .CK(clk), .QN(n714) );
  EDFFX1 R11_reg_4_ ( .D(data_in_2[106]), .E(n967), .CK(clk), .QN(n715) );
  EDFFX1 R11_reg_3_ ( .D(data_in_2[105]), .E(n967), .CK(clk), .QN(n716) );
  EDFFX1 R11_reg_2_ ( .D(data_in_2[104]), .E(n96), .CK(clk), .QN(n717) );
  EDFFX1 R11_reg_1_ ( .D(data_in_2[103]), .E(n959), .CK(clk), .QN(n718) );
  EDFFX1 R11_reg_0_ ( .D(data_in_2[102]), .E(n970), .CK(clk), .QN(n719) );
  EDFFX1 R15_reg_32_ ( .D(data_in_2[134]), .E(n1130), .CK(clk), .QN(n789) );
  EDFFX1 R15_reg_31_ ( .D(data_in_2[133]), .E(n1130), .CK(clk), .QN(n790) );
  EDFFX1 R15_reg_30_ ( .D(data_in_2[132]), .E(n1130), .CK(clk), .QN(n791) );
  EDFFX1 R15_reg_29_ ( .D(data_in_2[131]), .E(n1130), .CK(clk), .QN(n792) );
  EDFFX1 R15_reg_28_ ( .D(data_in_2[130]), .E(n1130), .CK(clk), .QN(n793) );
  EDFFX1 R15_reg_27_ ( .D(data_in_2[129]), .E(n1130), .CK(clk), .QN(n794) );
  EDFFX1 R15_reg_26_ ( .D(data_in_2[128]), .E(n1130), .CK(clk), .QN(n795) );
  EDFFX1 R15_reg_25_ ( .D(data_in_2[127]), .E(n1129), .CK(clk), .QN(n796) );
  EDFFX1 R15_reg_24_ ( .D(data_in_2[126]), .E(n1129), .CK(clk), .QN(n797) );
  EDFFX1 R15_reg_23_ ( .D(data_in_2[125]), .E(n1129), .CK(clk), .QN(n798) );
  EDFFX1 R15_reg_22_ ( .D(data_in_2[124]), .E(n1129), .CK(clk), .QN(n799) );
  EDFFX1 R15_reg_21_ ( .D(data_in_2[123]), .E(n1129), .CK(clk), .QN(n800) );
  EDFFX1 R15_reg_20_ ( .D(data_in_2[122]), .E(n1129), .CK(clk), .QN(n801) );
  EDFFX1 R15_reg_19_ ( .D(data_in_2[121]), .E(n1129), .CK(clk), .QN(n802) );
  EDFFX1 R15_reg_18_ ( .D(data_in_2[120]), .E(n1129), .CK(clk), .QN(n803) );
  EDFFX1 R15_reg_17_ ( .D(data_in_2[119]), .E(n1129), .CK(clk), .QN(n804) );
  EDFFX1 R15_reg_16_ ( .D(data_in_2[118]), .E(n1129), .CK(clk), .QN(n805) );
  EDFFX1 R15_reg_15_ ( .D(data_in_2[117]), .E(n1129), .CK(clk), .QN(n806) );
  EDFFX1 R15_reg_14_ ( .D(data_in_2[116]), .E(n1129), .CK(clk), .QN(n807) );
  EDFFX1 R15_reg_13_ ( .D(data_in_2[115]), .E(n1129), .CK(clk), .QN(n808) );
  EDFFX1 R15_reg_12_ ( .D(data_in_2[114]), .E(n1128), .CK(clk), .QN(n809) );
  EDFFX1 R15_reg_11_ ( .D(data_in_2[113]), .E(n1128), .CK(clk), .QN(n810) );
  EDFFX1 R15_reg_10_ ( .D(data_in_2[112]), .E(n1128), .CK(clk), .QN(n811) );
  EDFFX1 R15_reg_9_ ( .D(data_in_2[111]), .E(n1128), .CK(clk), .QN(n812) );
  EDFFX1 R15_reg_8_ ( .D(data_in_2[110]), .E(n1128), .CK(clk), .QN(n813) );
  EDFFX1 R15_reg_7_ ( .D(data_in_2[109]), .E(n1128), .CK(clk), .QN(n814) );
  EDFFX1 R15_reg_6_ ( .D(data_in_2[108]), .E(n1128), .CK(clk), .QN(n815) );
  EDFFX1 R15_reg_5_ ( .D(data_in_2[107]), .E(n1128), .CK(clk), .QN(n816) );
  EDFFX1 R15_reg_4_ ( .D(data_in_2[106]), .E(n1128), .CK(clk), .QN(n817) );
  EDFFX1 R15_reg_3_ ( .D(data_in_2[105]), .E(n1128), .CK(clk), .QN(n818) );
  EDFFX1 R15_reg_2_ ( .D(data_in_2[104]), .E(n1128), .CK(clk), .QN(n819) );
  EDFFX1 R15_reg_1_ ( .D(data_in_2[103]), .E(n1128), .CK(clk), .QN(n820) );
  EDFFX1 R15_reg_0_ ( .D(data_in_2[102]), .E(n1128), .CK(clk), .QN(n821) );
  EDFFX1 R3_reg_32_ ( .D(data_in_2[134]), .E(n97), .CK(clk), .QN(n857) );
  EDFFX1 R3_reg_31_ ( .D(data_in_2[133]), .E(n97), .CK(clk), .QN(n858) );
  EDFFX1 R3_reg_30_ ( .D(data_in_2[132]), .E(n97), .CK(clk), .QN(n859) );
  EDFFX1 R3_reg_29_ ( .D(data_in_2[131]), .E(n97), .CK(clk), .QN(n860) );
  EDFFX1 R3_reg_28_ ( .D(data_in_2[130]), .E(n97), .CK(clk), .QN(n861) );
  EDFFX1 R3_reg_27_ ( .D(data_in_2[129]), .E(n97), .CK(clk), .QN(n862) );
  EDFFX1 R3_reg_26_ ( .D(data_in_2[128]), .E(n97), .CK(clk), .QN(n863) );
  EDFFX1 R3_reg_25_ ( .D(data_in_2[127]), .E(n97), .CK(clk), .QN(n864) );
  EDFFX1 R3_reg_24_ ( .D(data_in_2[126]), .E(n97), .CK(clk), .QN(n865) );
  EDFFX1 R3_reg_23_ ( .D(data_in_2[125]), .E(n97), .CK(clk), .QN(n866) );
  EDFFX1 R3_reg_22_ ( .D(data_in_2[124]), .E(n97), .CK(clk), .QN(n867) );
  EDFFX1 R3_reg_21_ ( .D(data_in_2[123]), .E(n97), .CK(clk), .QN(n868) );
  EDFFX1 R3_reg_20_ ( .D(data_in_2[122]), .E(n97), .CK(clk), .QN(n869) );
  EDFFX1 R3_reg_19_ ( .D(data_in_2[121]), .E(n97), .CK(clk), .QN(n870) );
  EDFFX1 R3_reg_18_ ( .D(data_in_2[120]), .E(n1117), .CK(clk), .QN(n871) );
  EDFFX1 R3_reg_17_ ( .D(data_in_2[119]), .E(n1117), .CK(clk), .QN(n872) );
  EDFFX1 R3_reg_16_ ( .D(data_in_2[118]), .E(n97), .CK(clk), .QN(n873) );
  EDFFX1 R3_reg_15_ ( .D(data_in_2[117]), .E(n97), .CK(clk), .QN(n874) );
  EDFFX1 R3_reg_14_ ( .D(data_in_2[116]), .E(n97), .CK(clk), .QN(n875) );
  EDFFX1 R3_reg_13_ ( .D(data_in_2[115]), .E(n97), .CK(clk), .QN(n876) );
  EDFFX1 R3_reg_12_ ( .D(data_in_2[114]), .E(n97), .CK(clk), .QN(n877) );
  EDFFX1 R3_reg_11_ ( .D(data_in_2[113]), .E(n97), .CK(clk), .QN(n878) );
  EDFFX1 R3_reg_10_ ( .D(data_in_2[112]), .E(n97), .CK(clk), .QN(n879) );
  EDFFX1 R3_reg_9_ ( .D(data_in_2[111]), .E(n1117), .CK(clk), .QN(n880) );
  EDFFX1 R3_reg_8_ ( .D(data_in_2[110]), .E(n1117), .CK(clk), .QN(n881) );
  EDFFX1 R3_reg_7_ ( .D(data_in_2[109]), .E(n1117), .CK(clk), .QN(n882) );
  EDFFX1 R3_reg_6_ ( .D(data_in_2[108]), .E(n1117), .CK(clk), .QN(n883) );
  EDFFX1 R3_reg_5_ ( .D(data_in_2[107]), .E(n1117), .CK(clk), .QN(n884) );
  EDFFX1 R3_reg_4_ ( .D(data_in_2[106]), .E(n1117), .CK(clk), .QN(n885) );
  EDFFX1 R3_reg_3_ ( .D(data_in_2[105]), .E(n1117), .CK(clk), .QN(n886) );
  EDFFX1 R3_reg_2_ ( .D(data_in_2[104]), .E(n1117), .CK(clk), .QN(n887) );
  EDFFX1 R3_reg_1_ ( .D(data_in_2[103]), .E(n1117), .CK(clk), .QN(n888) );
  EDFFX1 R3_reg_0_ ( .D(data_in_2[102]), .E(n1117), .CK(clk), .QN(n889) );
  EDFFXL R7_reg_32_ ( .D(data_in_2[134]), .E(n1138), .CK(clk), .QN(n925) );
  EDFFXL R7_reg_31_ ( .D(data_in_2[133]), .E(n1138), .CK(clk), .QN(n926) );
  EDFFXL R7_reg_30_ ( .D(data_in_2[132]), .E(n1138), .CK(clk), .QN(n927) );
  EDFFXL R7_reg_29_ ( .D(data_in_2[131]), .E(n1138), .CK(clk), .QN(n928) );
  EDFFX1 R7_reg_28_ ( .D(data_in_2[130]), .E(n1138), .CK(clk), .QN(n929) );
  EDFFX1 R7_reg_27_ ( .D(data_in_2[129]), .E(n1138), .CK(clk), .QN(n930) );
  EDFFX1 R7_reg_26_ ( .D(data_in_2[128]), .E(n1138), .CK(clk), .QN(n931) );
  EDFFX1 R7_reg_25_ ( .D(data_in_2[127]), .E(n1138), .CK(clk), .QN(n932) );
  EDFFX1 R7_reg_24_ ( .D(data_in_2[126]), .E(n1138), .CK(clk), .QN(n933) );
  EDFFX1 R7_reg_23_ ( .D(data_in_2[125]), .E(n1138), .CK(clk), .QN(n934) );
  EDFFX1 R7_reg_22_ ( .D(data_in_2[124]), .E(n1138), .CK(clk), .QN(n935) );
  EDFFX1 R7_reg_21_ ( .D(data_in_2[123]), .E(n1138), .CK(clk), .QN(n936) );
  EDFFX1 R7_reg_20_ ( .D(data_in_2[122]), .E(n1138), .CK(clk), .QN(n937) );
  EDFFX1 R7_reg_19_ ( .D(data_in_2[121]), .E(n1138), .CK(clk), .QN(n938) );
  EDFFX1 R7_reg_18_ ( .D(data_in_2[120]), .E(n1138), .CK(clk), .QN(n939) );
  EDFFX1 R7_reg_17_ ( .D(data_in_2[119]), .E(n1138), .CK(clk), .QN(n940) );
  EDFFXL R7_reg_15_ ( .D(data_in_2[117]), .E(n1138), .CK(clk), .QN(n942) );
  EDFFXL R7_reg_14_ ( .D(data_in_2[116]), .E(n1138), .CK(clk), .QN(n943) );
  EDFFXL R7_reg_13_ ( .D(data_in_2[115]), .E(n1138), .CK(clk), .QN(n944) );
  EDFFXL R7_reg_12_ ( .D(data_in_2[114]), .E(n1138), .CK(clk), .QN(n945) );
  EDFFX1 R7_reg_11_ ( .D(data_in_2[113]), .E(n1138), .CK(clk), .QN(n946) );
  EDFFX1 R7_reg_10_ ( .D(data_in_2[112]), .E(n1138), .CK(clk), .QN(n947) );
  EDFFX1 R7_reg_9_ ( .D(data_in_2[111]), .E(n1138), .CK(clk), .QN(n948) );
  EDFFX1 R7_reg_8_ ( .D(data_in_2[110]), .E(n1138), .CK(clk), .QN(n949) );
  EDFFX1 R7_reg_7_ ( .D(data_in_2[109]), .E(n1138), .CK(clk), .QN(n950) );
  EDFFX1 R7_reg_6_ ( .D(data_in_2[108]), .E(n1138), .CK(clk), .QN(n951) );
  EDFFX1 R7_reg_5_ ( .D(data_in_2[107]), .E(n1138), .CK(clk), .QN(n952) );
  EDFFX1 R7_reg_4_ ( .D(data_in_2[106]), .E(n1138), .CK(clk), .QN(n953) );
  EDFFX1 R7_reg_3_ ( .D(data_in_2[105]), .E(n1138), .CK(clk), .QN(n954) );
  EDFFX1 R7_reg_2_ ( .D(data_in_2[104]), .E(n1138), .CK(clk), .QN(n955) );
  EDFFX1 R7_reg_1_ ( .D(data_in_2[103]), .E(n1138), .CK(clk), .QN(n956) );
  EDFFX1 R7_reg_0_ ( .D(data_in_2[102]), .E(n1138), .CK(clk), .QN(n957) );
  EDFFX1 R8_reg_31_ ( .D(data_in_2[31]), .E(n959), .CK(clk), .Q(R8[31]) );
  EDFFX1 R8_reg_30_ ( .D(data_in_2[30]), .E(n959), .CK(clk), .Q(R8[30]) );
  EDFFX1 R8_reg_29_ ( .D(data_in_2[29]), .E(n959), .CK(clk), .Q(R8[29]) );
  EDFFX1 R8_reg_22_ ( .D(data_in_2[22]), .E(n959), .CK(clk), .Q(R8[22]) );
  EDFFX1 R8_reg_21_ ( .D(data_in_2[21]), .E(n959), .CK(clk), .Q(R8[21]) );
  EDFFX1 R8_reg_20_ ( .D(data_in_2[20]), .E(n960), .CK(clk), .Q(R8[20]) );
  EDFFX1 R8_reg_19_ ( .D(data_in_2[19]), .E(n960), .CK(clk), .Q(R8[19]) );
  EDFFX1 R8_reg_18_ ( .D(data_in_2[18]), .E(n960), .CK(clk), .Q(R8[18]) );
  EDFFX1 R8_reg_17_ ( .D(data_in_2[17]), .E(n960), .CK(clk), .Q(R8[17]) );
  EDFFX1 R8_reg_13_ ( .D(data_in_2[13]), .E(n960), .CK(clk), .Q(R8[13]) );
  EDFFX1 R8_reg_12_ ( .D(data_in_2[12]), .E(n960), .CK(clk), .Q(R8[12]) );
  EDFFX1 R8_reg_5_ ( .D(data_in_2[5]), .E(n96), .CK(clk), .Q(R8[5]) );
  EDFFX1 R8_reg_4_ ( .D(data_in_2[4]), .E(n96), .CK(clk), .Q(R8[4]) );
  EDFFX1 R8_reg_3_ ( .D(data_in_2[3]), .E(n963), .CK(clk), .Q(R8[3]) );
  EDFFX1 R8_reg_2_ ( .D(data_in_2[2]), .E(n967), .CK(clk), .Q(R8[2]) );
  EDFFX1 R8_reg_1_ ( .D(data_in_2[1]), .E(n968), .CK(clk), .Q(R8[1]) );
  EDFFX1 R8_reg_0_ ( .D(data_in_2[0]), .E(n960), .CK(clk), .Q(R8[0]) );
  EDFFX1 R12_reg_31_ ( .D(data_in_2[31]), .E(n1130), .CK(clk), .Q(R12[31]) );
  EDFFX1 R12_reg_30_ ( .D(data_in_2[30]), .E(n1129), .CK(clk), .Q(R12[30]) );
  EDFFX1 R12_reg_29_ ( .D(data_in_2[29]), .E(n1128), .CK(clk), .Q(R12[29]) );
  EDFFX1 R12_reg_22_ ( .D(data_in_2[22]), .E(n1134), .CK(clk), .Q(R12[22]) );
  EDFFX1 R12_reg_21_ ( .D(data_in_2[21]), .E(n1134), .CK(clk), .Q(R12[21]) );
  EDFFX1 R12_reg_20_ ( .D(data_in_2[20]), .E(n1134), .CK(clk), .Q(R12[20]) );
  EDFFX1 R12_reg_19_ ( .D(data_in_2[19]), .E(n1134), .CK(clk), .Q(R12[19]) );
  EDFFX1 R12_reg_18_ ( .D(data_in_2[18]), .E(n1134), .CK(clk), .Q(R12[18]) );
  EDFFX1 R12_reg_17_ ( .D(data_in_2[17]), .E(n1134), .CK(clk), .Q(R12[17]) );
  EDFFX1 R12_reg_13_ ( .D(data_in_2[13]), .E(n1134), .CK(clk), .Q(R12[13]) );
  EDFFX1 R12_reg_12_ ( .D(data_in_2[12]), .E(n1134), .CK(clk), .Q(R12[12]) );
  EDFFX1 R12_reg_5_ ( .D(data_in_2[5]), .E(n1133), .CK(clk), .Q(R12[5]) );
  EDFFX1 R12_reg_4_ ( .D(data_in_2[4]), .E(n1133), .CK(clk), .Q(R12[4]) );
  EDFFX1 R12_reg_3_ ( .D(data_in_2[3]), .E(n1133), .CK(clk), .Q(R12[3]) );
  EDFFX1 R12_reg_2_ ( .D(data_in_2[2]), .E(n1133), .CK(clk), .Q(R12[2]) );
  EDFFX1 R12_reg_1_ ( .D(data_in_2[1]), .E(n1133), .CK(clk), .Q(R12[1]) );
  EDFFX1 R12_reg_0_ ( .D(data_in_2[0]), .E(n1133), .CK(clk), .Q(R12[0]) );
  EDFFX1 R0_reg_31_ ( .D(data_in_2[31]), .E(n1117), .CK(clk), .Q(R0[31]) );
  EDFFX1 R0_reg_30_ ( .D(data_in_2[30]), .E(n1117), .CK(clk), .Q(R0[30]) );
  EDFFX1 R0_reg_29_ ( .D(data_in_2[29]), .E(n1117), .CK(clk), .Q(R0[29]) );
  EDFFX1 R0_reg_22_ ( .D(data_in_2[22]), .E(n1117), .CK(clk), .Q(R0[22]) );
  EDFFX1 R0_reg_21_ ( .D(data_in_2[21]), .E(n1117), .CK(clk), .Q(R0[21]) );
  EDFFX1 R0_reg_20_ ( .D(data_in_2[20]), .E(n1117), .CK(clk), .Q(R0[20]) );
  EDFFX1 R0_reg_19_ ( .D(data_in_2[19]), .E(n1117), .CK(clk), .Q(R0[19]) );
  EDFFX1 R0_reg_18_ ( .D(data_in_2[18]), .E(n1117), .CK(clk), .Q(R0[18]) );
  EDFFX1 R0_reg_17_ ( .D(data_in_2[17]), .E(n1117), .CK(clk), .Q(R0[17]) );
  EDFFX1 R0_reg_13_ ( .D(data_in_2[13]), .E(n1117), .CK(clk), .Q(R0[13]) );
  EDFFX1 R0_reg_12_ ( .D(data_in_2[12]), .E(n1117), .CK(clk), .Q(R0[12]) );
  EDFFX1 R0_reg_5_ ( .D(data_in_2[5]), .E(n1117), .CK(clk), .Q(R0[5]) );
  EDFFX1 R0_reg_4_ ( .D(data_in_2[4]), .E(n1117), .CK(clk), .Q(R0[4]) );
  EDFFX1 R0_reg_3_ ( .D(data_in_2[3]), .E(n1117), .CK(clk), .Q(R0[3]) );
  EDFFX1 R0_reg_2_ ( .D(data_in_2[2]), .E(n1117), .CK(clk), .Q(R0[2]) );
  EDFFX1 R0_reg_1_ ( .D(data_in_2[1]), .E(n1117), .CK(clk), .Q(R0[1]) );
  EDFFX1 R0_reg_0_ ( .D(data_in_2[0]), .E(n1117), .CK(clk), .Q(R0[0]) );
  EDFFXL R4_reg_31_ ( .D(data_in_2[31]), .E(n969), .CK(clk), .Q(R4[31]) );
  EDFFXL R4_reg_30_ ( .D(data_in_2[30]), .E(n969), .CK(clk), .Q(R4[30]) );
  EDFFXL R4_reg_29_ ( .D(data_in_2[29]), .E(n969), .CK(clk), .Q(R4[29]) );
  EDFFX1 R4_reg_22_ ( .D(data_in_2[22]), .E(n969), .CK(clk), .Q(R4[22]) );
  EDFFX1 R4_reg_21_ ( .D(data_in_2[21]), .E(n969), .CK(clk), .Q(R4[21]) );
  EDFFX1 R4_reg_20_ ( .D(data_in_2[20]), .E(n969), .CK(clk), .Q(R4[20]) );
  EDFFX1 R4_reg_19_ ( .D(data_in_2[19]), .E(n969), .CK(clk), .Q(R4[19]) );
  EDFFX1 R4_reg_18_ ( .D(data_in_2[18]), .E(n969), .CK(clk), .Q(R4[18]) );
  EDFFX1 R4_reg_17_ ( .D(data_in_2[17]), .E(n1136), .CK(clk), .Q(R4[17]) );
  EDFFXL R4_reg_16_ ( .D(data_in_2[16]), .E(n969), .CK(clk), .Q(R4[16]) );
  EDFFXL R4_reg_15_ ( .D(data_in_2[15]), .E(n969), .CK(clk), .Q(R4[15]) );
  EDFFXL R4_reg_13_ ( .D(data_in_2[13]), .E(n969), .CK(clk), .Q(R4[13]) );
  EDFFXL R4_reg_12_ ( .D(data_in_2[12]), .E(n969), .CK(clk), .Q(R4[12]) );
  EDFFX1 R4_reg_5_ ( .D(data_in_2[5]), .E(n1137), .CK(clk), .Q(R4[5]) );
  EDFFX1 R4_reg_4_ ( .D(data_in_2[4]), .E(n1138), .CK(clk), .Q(R4[4]) );
  EDFFX1 R4_reg_3_ ( .D(data_in_2[3]), .E(n1136), .CK(clk), .Q(R4[3]) );
  EDFFX1 R4_reg_2_ ( .D(data_in_2[2]), .E(n1138), .CK(clk), .Q(R4[2]) );
  EDFFX1 R4_reg_1_ ( .D(data_in_2[1]), .E(n1136), .CK(clk), .Q(R4[1]) );
  EDFFX1 R4_reg_0_ ( .D(data_in_2[0]), .E(n1136), .CK(clk), .Q(R4[0]) );
  EDFFXL R13_reg_33_ ( .D(data_in_2[67]), .E(n1133), .CK(clk), .Q(R13[33]) );
  EDFFXL R13_reg_32_ ( .D(data_in_2[66]), .E(n1133), .CK(clk), .Q(R13[32]) );
  EDFFXL R13_reg_31_ ( .D(data_in_2[65]), .E(n1133), .CK(clk), .Q(R13[31]) );
  EDFFXL R13_reg_30_ ( .D(data_in_2[64]), .E(n1132), .CK(clk), .Q(R13[30]) );
  EDFFXL R13_reg_29_ ( .D(data_in_2[63]), .E(n1133), .CK(clk), .Q(R13[29]) );
  EDFFX1 R13_reg_28_ ( .D(data_in_2[62]), .E(n1133), .CK(clk), .Q(R13[28]) );
  EDFFX1 R13_reg_27_ ( .D(data_in_2[61]), .E(n1133), .CK(clk), .Q(R13[27]) );
  EDFFX1 R13_reg_26_ ( .D(data_in_2[60]), .E(n1132), .CK(clk), .Q(R13[26]) );
  EDFFX1 R13_reg_25_ ( .D(data_in_2[59]), .E(n1131), .CK(clk), .Q(R13[25]) );
  EDFFX1 R13_reg_24_ ( .D(data_in_2[58]), .E(n1130), .CK(clk), .Q(R13[24]) );
  EDFFX1 R13_reg_23_ ( .D(data_in_2[57]), .E(n1129), .CK(clk), .Q(R13[23]) );
  EDFFX1 R13_reg_22_ ( .D(data_in_2[56]), .E(n1128), .CK(clk), .Q(R13[22]) );
  EDFFX1 R13_reg_21_ ( .D(data_in_2[55]), .E(n1128), .CK(clk), .Q(R13[21]) );
  EDFFX1 R13_reg_20_ ( .D(data_in_2[54]), .E(n1134), .CK(clk), .Q(R13[20]) );
  EDFFX1 R13_reg_19_ ( .D(data_in_2[53]), .E(n1133), .CK(clk), .Q(R13[19]) );
  EDFFX1 R13_reg_18_ ( .D(data_in_2[52]), .E(n1132), .CK(clk), .Q(R13[18]) );
  EDFFX1 R13_reg_17_ ( .D(data_in_2[51]), .E(n1130), .CK(clk), .Q(R13[17]) );
  EDFFXL R13_reg_14_ ( .D(data_in_2[48]), .E(n971), .CK(clk), .Q(R13[14]) );
  EDFFXL R13_reg_13_ ( .D(data_in_2[47]), .E(n971), .CK(clk), .Q(R13[13]) );
  EDFFXL R13_reg_12_ ( .D(data_in_2[46]), .E(n971), .CK(clk), .Q(R13[12]) );
  EDFFX1 R13_reg_11_ ( .D(data_in_2[45]), .E(n1130), .CK(clk), .Q(R13[11]) );
  EDFFX1 R13_reg_10_ ( .D(data_in_2[44]), .E(n1131), .CK(clk), .Q(R13[10]) );
  EDFFX1 R13_reg_9_ ( .D(data_in_2[43]), .E(n1129), .CK(clk), .Q(R13[9]) );
  EDFFX1 R13_reg_8_ ( .D(data_in_2[42]), .E(n1128), .CK(clk), .Q(R13[8]) );
  EDFFX1 R13_reg_7_ ( .D(data_in_2[41]), .E(n1134), .CK(clk), .Q(R13[7]) );
  EDFFX1 R13_reg_6_ ( .D(data_in_2[40]), .E(n1133), .CK(clk), .Q(R13[6]) );
  EDFFX1 R13_reg_5_ ( .D(data_in_2[39]), .E(n1132), .CK(clk), .Q(R13[5]) );
  EDFFX1 R13_reg_4_ ( .D(data_in_2[38]), .E(n1130), .CK(clk), .Q(R13[4]) );
  EDFFX1 R13_reg_3_ ( .D(data_in_2[37]), .E(n1131), .CK(clk), .Q(R13[3]) );
  EDFFX1 R13_reg_2_ ( .D(data_in_2[36]), .E(n1129), .CK(clk), .Q(R13[2]) );
  EDFFX1 R13_reg_1_ ( .D(data_in_2[35]), .E(n1128), .CK(clk), .Q(R13[1]) );
  EDFFX1 R13_reg_0_ ( .D(data_in_2[34]), .E(n1131), .CK(clk), .Q(R13[0]) );
  EDFFXL R9_reg_33_ ( .D(data_in_2[67]), .E(n970), .CK(clk), .Q(R9[33]) );
  EDFFXL R9_reg_32_ ( .D(data_in_2[66]), .E(n970), .CK(clk), .Q(R9[32]) );
  EDFFXL R9_reg_31_ ( .D(data_in_2[65]), .E(n972), .CK(clk), .Q(R9[31]) );
  EDFFXL R9_reg_30_ ( .D(data_in_2[64]), .E(n972), .CK(clk), .Q(R9[30]) );
  EDFFXL R9_reg_29_ ( .D(data_in_2[63]), .E(n972), .CK(clk), .Q(R9[29]) );
  EDFFX1 R9_reg_28_ ( .D(data_in_2[62]), .E(n972), .CK(clk), .Q(R9[28]) );
  EDFFX1 R9_reg_27_ ( .D(data_in_2[61]), .E(n972), .CK(clk), .Q(R9[27]) );
  EDFFX1 R9_reg_26_ ( .D(data_in_2[60]), .E(n972), .CK(clk), .Q(R9[26]) );
  EDFFX1 R9_reg_25_ ( .D(data_in_2[59]), .E(n972), .CK(clk), .Q(R9[25]) );
  EDFFX1 R9_reg_24_ ( .D(data_in_2[58]), .E(n972), .CK(clk), .Q(R9[24]) );
  EDFFX1 R9_reg_23_ ( .D(data_in_2[57]), .E(n972), .CK(clk), .Q(R9[23]) );
  EDFFX1 R9_reg_22_ ( .D(data_in_2[56]), .E(n972), .CK(clk), .Q(R9[22]) );
  EDFFX1 R9_reg_21_ ( .D(data_in_2[55]), .E(n972), .CK(clk), .Q(R9[21]) );
  EDFFX1 R9_reg_20_ ( .D(data_in_2[54]), .E(n972), .CK(clk), .Q(R9[20]) );
  EDFFX1 R9_reg_19_ ( .D(data_in_2[53]), .E(n972), .CK(clk), .Q(R9[19]) );
  EDFFX1 R9_reg_18_ ( .D(data_in_2[52]), .E(n96), .CK(clk), .Q(R9[18]) );
  EDFFX1 R9_reg_17_ ( .D(data_in_2[51]), .E(n96), .CK(clk), .Q(R9[17]) );
  EDFFXL R9_reg_15_ ( .D(data_in_2[49]), .E(n96), .CK(clk), .Q(R9[15]) );
  EDFFXL R9_reg_14_ ( .D(data_in_2[48]), .E(n96), .CK(clk), .Q(R9[14]) );
  EDFFXL R9_reg_13_ ( .D(data_in_2[47]), .E(n96), .CK(clk), .Q(R9[13]) );
  EDFFXL R9_reg_12_ ( .D(data_in_2[46]), .E(n96), .CK(clk), .Q(R9[12]) );
  EDFFX1 R9_reg_11_ ( .D(data_in_2[45]), .E(n96), .CK(clk), .Q(R9[11]) );
  EDFFX1 R9_reg_10_ ( .D(data_in_2[44]), .E(n96), .CK(clk), .Q(R9[10]) );
  EDFFX1 R9_reg_9_ ( .D(data_in_2[43]), .E(n96), .CK(clk), .Q(R9[9]) );
  EDFFX1 R9_reg_8_ ( .D(data_in_2[42]), .E(n96), .CK(clk), .Q(R9[8]) );
  EDFFX1 R9_reg_7_ ( .D(data_in_2[41]), .E(n963), .CK(clk), .Q(R9[7]) );
  EDFFX1 R9_reg_6_ ( .D(data_in_2[40]), .E(n967), .CK(clk), .Q(R9[6]) );
  EDFFX1 R9_reg_5_ ( .D(data_in_2[39]), .E(n960), .CK(clk), .Q(R9[5]) );
  EDFFX1 R9_reg_4_ ( .D(data_in_2[38]), .E(n959), .CK(clk), .Q(R9[4]) );
  EDFFX1 R9_reg_3_ ( .D(data_in_2[37]), .E(n959), .CK(clk), .Q(R9[3]) );
  EDFFX1 R9_reg_2_ ( .D(data_in_2[36]), .E(n959), .CK(clk), .Q(R9[2]) );
  EDFFX1 R9_reg_1_ ( .D(data_in_2[35]), .E(n959), .CK(clk), .Q(R9[1]) );
  EDFFX1 R9_reg_0_ ( .D(data_in_2[34]), .E(n959), .CK(clk), .Q(R9[0]) );
  EDFFXL R1_reg_33_ ( .D(data_in_2[67]), .E(n97), .CK(clk), .Q(R1[33]) );
  EDFFXL R1_reg_32_ ( .D(data_in_2[66]), .E(n97), .CK(clk), .Q(R1[32]) );
  EDFFXL R1_reg_31_ ( .D(data_in_2[65]), .E(n97), .CK(clk), .Q(R1[31]) );
  EDFFXL R1_reg_30_ ( .D(data_in_2[64]), .E(n97), .CK(clk), .Q(R1[30]) );
  EDFFXL R1_reg_29_ ( .D(data_in_2[63]), .E(n97), .CK(clk), .Q(R1[29]) );
  EDFFX1 R1_reg_28_ ( .D(data_in_2[62]), .E(n97), .CK(clk), .Q(R1[28]) );
  EDFFX1 R1_reg_27_ ( .D(data_in_2[61]), .E(n97), .CK(clk), .Q(R1[27]) );
  EDFFX1 R1_reg_26_ ( .D(data_in_2[60]), .E(n97), .CK(clk), .Q(R1[26]) );
  EDFFX1 R1_reg_25_ ( .D(data_in_2[59]), .E(n97), .CK(clk), .Q(R1[25]) );
  EDFFX1 R1_reg_24_ ( .D(data_in_2[58]), .E(n97), .CK(clk), .Q(R1[24]) );
  EDFFX1 R1_reg_23_ ( .D(data_in_2[57]), .E(n97), .CK(clk), .Q(R1[23]) );
  EDFFX1 R1_reg_22_ ( .D(data_in_2[56]), .E(n97), .CK(clk), .Q(R1[22]) );
  EDFFX1 R1_reg_21_ ( .D(data_in_2[55]), .E(n97), .CK(clk), .Q(R1[21]) );
  EDFFX1 R1_reg_20_ ( .D(data_in_2[54]), .E(n97), .CK(clk), .Q(R1[20]) );
  EDFFX1 R1_reg_19_ ( .D(data_in_2[53]), .E(n97), .CK(clk), .Q(R1[19]) );
  EDFFX1 R1_reg_18_ ( .D(data_in_2[52]), .E(n97), .CK(clk), .Q(R1[18]) );
  EDFFX1 R1_reg_17_ ( .D(data_in_2[51]), .E(n97), .CK(clk), .Q(R1[17]) );
  EDFFXL R1_reg_15_ ( .D(data_in_2[49]), .E(n97), .CK(clk), .Q(R1[15]) );
  EDFFXL R1_reg_14_ ( .D(data_in_2[48]), .E(n97), .CK(clk), .Q(R1[14]) );
  EDFFXL R1_reg_13_ ( .D(data_in_2[47]), .E(n97), .CK(clk), .Q(R1[13]) );
  EDFFXL R1_reg_12_ ( .D(data_in_2[46]), .E(n97), .CK(clk), .Q(R1[12]) );
  EDFFX1 R1_reg_11_ ( .D(data_in_2[45]), .E(n97), .CK(clk), .Q(R1[11]) );
  EDFFX1 R1_reg_10_ ( .D(data_in_2[44]), .E(n97), .CK(clk), .Q(R1[10]) );
  EDFFX1 R1_reg_9_ ( .D(data_in_2[43]), .E(n97), .CK(clk), .Q(R1[9]) );
  EDFFX1 R1_reg_8_ ( .D(data_in_2[42]), .E(n97), .CK(clk), .Q(R1[8]) );
  EDFFX1 R1_reg_7_ ( .D(data_in_2[41]), .E(n97), .CK(clk), .Q(R1[7]) );
  EDFFX1 R1_reg_6_ ( .D(data_in_2[40]), .E(n97), .CK(clk), .Q(R1[6]) );
  EDFFX1 R1_reg_5_ ( .D(data_in_2[39]), .E(n97), .CK(clk), .Q(R1[5]) );
  EDFFX1 R1_reg_4_ ( .D(data_in_2[38]), .E(n97), .CK(clk), .Q(R1[4]) );
  EDFFX1 R1_reg_3_ ( .D(data_in_2[37]), .E(n97), .CK(clk), .Q(R1[3]) );
  EDFFX1 R1_reg_2_ ( .D(data_in_2[36]), .E(n97), .CK(clk), .Q(R1[2]) );
  EDFFX1 R1_reg_1_ ( .D(data_in_2[35]), .E(n97), .CK(clk), .Q(R1[1]) );
  EDFFX1 R1_reg_0_ ( .D(data_in_2[34]), .E(n97), .CK(clk), .Q(R1[0]) );
  EDFFXL R5_reg_33_ ( .D(data_in_2[67]), .E(n1136), .CK(clk), .Q(R5[33]) );
  EDFFXL R5_reg_32_ ( .D(data_in_2[66]), .E(n1136), .CK(clk), .Q(R5[32]) );
  EDFFXL R5_reg_31_ ( .D(data_in_2[65]), .E(n1136), .CK(clk), .Q(R5[31]) );
  EDFFXL R5_reg_30_ ( .D(data_in_2[64]), .E(n1136), .CK(clk), .Q(R5[30]) );
  EDFFXL R5_reg_29_ ( .D(data_in_2[63]), .E(n1136), .CK(clk), .Q(R5[29]) );
  EDFFX1 R5_reg_28_ ( .D(data_in_2[62]), .E(n1136), .CK(clk), .Q(R5[28]) );
  EDFFX1 R5_reg_27_ ( .D(data_in_2[61]), .E(n1136), .CK(clk), .Q(R5[27]) );
  EDFFX1 R5_reg_26_ ( .D(data_in_2[60]), .E(n1136), .CK(clk), .Q(R5[26]) );
  EDFFX1 R5_reg_25_ ( .D(data_in_2[59]), .E(n1136), .CK(clk), .Q(R5[25]) );
  EDFFX1 R5_reg_24_ ( .D(data_in_2[58]), .E(n1136), .CK(clk), .Q(R5[24]) );
  EDFFX1 R5_reg_23_ ( .D(data_in_2[57]), .E(n1136), .CK(clk), .Q(R5[23]) );
  EDFFX1 R5_reg_22_ ( .D(data_in_2[56]), .E(n1136), .CK(clk), .Q(R5[22]) );
  EDFFX1 R5_reg_21_ ( .D(data_in_2[55]), .E(n1136), .CK(clk), .Q(R5[21]) );
  EDFFX1 R5_reg_20_ ( .D(data_in_2[54]), .E(n1136), .CK(clk), .Q(R5[20]) );
  EDFFX1 R5_reg_19_ ( .D(data_in_2[53]), .E(n1136), .CK(clk), .Q(R5[19]) );
  EDFFX1 R5_reg_18_ ( .D(data_in_2[52]), .E(n1136), .CK(clk), .Q(R5[18]) );
  EDFFX1 R5_reg_17_ ( .D(data_in_2[51]), .E(n1136), .CK(clk), .Q(R5[17]) );
  EDFFXL R5_reg_15_ ( .D(data_in_2[49]), .E(n1136), .CK(clk), .Q(R5[15]) );
  EDFFXL R5_reg_14_ ( .D(data_in_2[48]), .E(n1136), .CK(clk), .Q(R5[14]) );
  EDFFXL R5_reg_13_ ( .D(data_in_2[47]), .E(n1136), .CK(clk), .Q(R5[13]) );
  EDFFXL R5_reg_12_ ( .D(data_in_2[46]), .E(n1136), .CK(clk), .Q(R5[12]) );
  EDFFX1 R5_reg_11_ ( .D(data_in_2[45]), .E(n1136), .CK(clk), .Q(R5[11]) );
  EDFFX1 R5_reg_10_ ( .D(data_in_2[44]), .E(n1136), .CK(clk), .Q(R5[10]) );
  EDFFX1 R5_reg_9_ ( .D(data_in_2[43]), .E(n1136), .CK(clk), .Q(R5[9]) );
  EDFFX1 R5_reg_8_ ( .D(data_in_2[42]), .E(n1136), .CK(clk), .Q(R5[8]) );
  EDFFX1 R5_reg_7_ ( .D(data_in_2[41]), .E(n1136), .CK(clk), .Q(R5[7]) );
  EDFFX1 R5_reg_6_ ( .D(data_in_2[40]), .E(n1136), .CK(clk), .Q(R5[6]) );
  EDFFX1 R5_reg_5_ ( .D(data_in_2[39]), .E(n1136), .CK(clk), .Q(R5[5]) );
  EDFFX1 R5_reg_4_ ( .D(data_in_2[38]), .E(n1136), .CK(clk), .Q(R5[4]) );
  EDFFX1 R5_reg_3_ ( .D(data_in_2[37]), .E(n1136), .CK(clk), .Q(R5[3]) );
  EDFFX1 R5_reg_2_ ( .D(data_in_2[36]), .E(n1136), .CK(clk), .Q(R5[2]) );
  EDFFX1 R5_reg_1_ ( .D(data_in_2[35]), .E(n1136), .CK(clk), .Q(R5[1]) );
  EDFFX1 R5_reg_0_ ( .D(data_in_2[34]), .E(n1137), .CK(clk), .Q(R5[0]) );
  DFFHQX1 reg_flag_mux_reg ( .D(n1169), .CK(clk), .Q(reg_flag_mux) );
  EDFFX1 data_out_2_reg_33_ ( .D(N85), .E(n1166), .CK(clk), .Q(data_out_2[33])
         );
  EDFFX1 data_out_2_reg_32_ ( .D(N84), .E(n1166), .CK(clk), .Q(data_out_2[32])
         );
  EDFFX1 data_out_2_reg_16_ ( .D(N68), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[16]) );
  EDFFX1 data_out_2_reg_15_ ( .D(N67), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[15]) );
  DFFHQX1 counter1_reg_0_ ( .D(n1116), .CK(clk), .Q(counter1[0]) );
  DFFHQX1 counter1_reg_1_ ( .D(n1115), .CK(clk), .Q(counter1[1]) );
  DFFHQX1 counter2_reg_0_ ( .D(n1114), .CK(clk), .Q(counter2[0]) );
  DFFHQX1 counter2_reg_1_ ( .D(n1113), .CK(clk), .Q(counter2[1]) );
  EDFFX1 data_out_2_reg_30_ ( .D(N82), .E(n1166), .CK(clk), .Q(data_out_2[30])
         );
  EDFFX1 data_out_2_reg_31_ ( .D(N83), .E(n1166), .CK(clk), .Q(data_out_2[31])
         );
  EDFFX1 data_out_2_reg_29_ ( .D(N81), .E(n1166), .CK(clk), .Q(data_out_2[29])
         );
  EDFFX1 data_out_2_reg_28_ ( .D(N80), .E(n1166), .CK(clk), .Q(data_out_2[28])
         );
  EDFFX1 data_out_2_reg_27_ ( .D(N79), .E(n1166), .CK(clk), .Q(data_out_2[27])
         );
  EDFFX1 data_out_2_reg_14_ ( .D(N66), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[14]) );
  EDFFX1 data_out_2_reg_13_ ( .D(N65), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[13]) );
  EDFFX1 data_out_2_reg_12_ ( .D(N64), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[12]) );
  EDFFX1 data_out_2_reg_11_ ( .D(N63), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[11]) );
  EDFFX1 data_out_2_reg_10_ ( .D(N62), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[10]) );
  EDFFX1 data_out_2_reg_26_ ( .D(N78), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[26]) );
  EDFFX1 data_out_2_reg_25_ ( .D(N77), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[25]) );
  EDFFX1 data_out_2_reg_24_ ( .D(N76), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[24]) );
  EDFFX1 data_out_2_reg_23_ ( .D(N75), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[23]) );
  EDFFX1 data_out_2_reg_22_ ( .D(N74), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[22]) );
  EDFFX1 data_out_2_reg_21_ ( .D(N73), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[21]) );
  EDFFX1 data_out_2_reg_9_ ( .D(N61), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[9]) );
  EDFFX1 data_out_2_reg_8_ ( .D(N60), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[8]) );
  EDFFX1 data_out_2_reg_7_ ( .D(N59), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[7]) );
  EDFFX1 data_out_2_reg_6_ ( .D(N58), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[6]) );
  EDFFX1 data_out_2_reg_5_ ( .D(N57), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[5]) );
  EDFFX1 data_out_2_reg_4_ ( .D(N56), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[4]) );
  EDFFX1 data_out_2_reg_20_ ( .D(N72), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[20]) );
  EDFFX1 data_out_2_reg_19_ ( .D(N71), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[19]) );
  EDFFX1 data_out_2_reg_18_ ( .D(N70), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[18]) );
  EDFFX1 data_out_2_reg_17_ ( .D(N69), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[17]) );
  EDFFX1 data_out_2_reg_3_ ( .D(N55), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[3]) );
  EDFFX1 data_out_2_reg_2_ ( .D(N54), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[2]) );
  EDFFX1 data_out_2_reg_1_ ( .D(N53), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[1]) );
  EDFFX1 data_out_2_reg_0_ ( .D(N52), .E(n1166), .CK(clk), .Q(data_out_2[0])
         );
  EDFFX1 data_out_2_reg_134_ ( .D(N186), .E(n1167), .CK(clk), .Q(
        data_out_2[134]) );
  EDFFX1 data_out_2_reg_133_ ( .D(N185), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[133]) );
  EDFFX1 data_out_2_reg_132_ ( .D(N184), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[132]) );
  EDFFX1 data_out_2_reg_117_ ( .D(N169), .E(n1167), .CK(clk), .Q(
        data_out_2[117]) );
  EDFFX1 data_out_2_reg_116_ ( .D(N168), .E(n1167), .CK(clk), .Q(
        data_out_2[116]) );
  EDFFX1 data_out_2_reg_100_ ( .D(N152), .E(n1167), .CK(clk), .Q(
        data_out_2[100]) );
  EDFFX1 data_out_2_reg_99_ ( .D(N151), .E(n1167), .CK(clk), .Q(data_out_2[99]) );
  EDFFX1 data_out_2_reg_98_ ( .D(N150), .E(n1167), .CK(clk), .Q(data_out_2[98]) );
  EDFFX1 data_out_2_reg_83_ ( .D(N135), .E(n1167), .CK(clk), .Q(data_out_2[83]) );
  EDFFX1 data_out_2_reg_82_ ( .D(N134), .E(n1166), .CK(clk), .Q(data_out_2[82]) );
  EDFFX1 data_out_2_reg_66_ ( .D(N118), .E(n1167), .CK(clk), .Q(data_out_2[66]) );
  EDFFX1 data_out_2_reg_65_ ( .D(N117), .E(n1166), .CK(clk), .Q(data_out_2[65]) );
  EDFFX1 data_out_2_reg_64_ ( .D(N116), .E(n1167), .CK(clk), .Q(data_out_2[64]) );
  EDFFX1 data_out_2_reg_49_ ( .D(N101), .E(n1166), .CK(clk), .Q(data_out_2[49]) );
  EDFFX1 data_out_2_reg_48_ ( .D(N100), .E(n1166), .CK(clk), .Q(data_out_2[48]) );
  EDFFX1 data_out_2_reg_47_ ( .D(N99), .E(n1166), .CK(clk), .Q(data_out_2[47])
         );
  EDFFX1 data_out_2_reg_131_ ( .D(N183), .E(n1167), .CK(clk), .Q(
        data_out_2[131]) );
  EDFFX1 data_out_2_reg_130_ ( .D(N182), .E(n1166), .CK(clk), .Q(
        data_out_2[130]) );
  EDFFX1 data_out_2_reg_129_ ( .D(N181), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[129]) );
  EDFFX1 data_out_2_reg_128_ ( .D(N180), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[128]) );
  EDFFX1 data_out_2_reg_115_ ( .D(N167), .E(n1167), .CK(clk), .Q(
        data_out_2[115]) );
  EDFFX1 data_out_2_reg_114_ ( .D(N166), .E(n1167), .CK(clk), .Q(
        data_out_2[114]) );
  EDFFX1 data_out_2_reg_113_ ( .D(N165), .E(n1167), .CK(clk), .Q(
        data_out_2[113]) );
  EDFFX1 data_out_2_reg_112_ ( .D(N164), .E(n1167), .CK(clk), .Q(
        data_out_2[112]) );
  EDFFX1 data_out_2_reg_111_ ( .D(N163), .E(n1167), .CK(clk), .Q(
        data_out_2[111]) );
  EDFFX1 data_out_2_reg_97_ ( .D(N149), .E(n1167), .CK(clk), .Q(data_out_2[97]) );
  EDFFX1 data_out_2_reg_96_ ( .D(N148), .E(n1167), .CK(clk), .Q(data_out_2[96]) );
  EDFFX1 data_out_2_reg_95_ ( .D(N147), .E(n1167), .CK(clk), .Q(data_out_2[95]) );
  EDFFX1 data_out_2_reg_94_ ( .D(N146), .E(n1167), .CK(clk), .Q(data_out_2[94]) );
  EDFFX1 data_out_2_reg_81_ ( .D(N133), .E(n1166), .CK(clk), .Q(data_out_2[81]) );
  EDFFX1 data_out_2_reg_80_ ( .D(N132), .E(n1167), .CK(clk), .Q(data_out_2[80]) );
  EDFFX1 data_out_2_reg_79_ ( .D(N131), .E(n1166), .CK(clk), .Q(data_out_2[79]) );
  EDFFX1 data_out_2_reg_78_ ( .D(N130), .E(n1167), .CK(clk), .Q(data_out_2[78]) );
  EDFFX1 data_out_2_reg_63_ ( .D(N115), .E(n1166), .CK(clk), .Q(data_out_2[63]) );
  EDFFX1 data_out_2_reg_62_ ( .D(N114), .E(n1167), .CK(clk), .Q(data_out_2[62]) );
  EDFFX1 data_out_2_reg_61_ ( .D(N113), .E(n1166), .CK(clk), .Q(data_out_2[61]) );
  EDFFX1 data_out_2_reg_60_ ( .D(N112), .E(n1167), .CK(clk), .Q(data_out_2[60]) );
  EDFFX1 data_out_2_reg_46_ ( .D(N98), .E(n1166), .CK(clk), .Q(data_out_2[46])
         );
  EDFFX1 data_out_2_reg_45_ ( .D(N97), .E(n1166), .CK(clk), .Q(data_out_2[45])
         );
  EDFFX1 data_out_2_reg_44_ ( .D(N96), .E(n1166), .CK(clk), .Q(data_out_2[44])
         );
  EDFFX1 data_out_2_reg_43_ ( .D(N95), .E(n1166), .CK(clk), .Q(data_out_2[43])
         );
  EDFFX1 data_out_2_reg_127_ ( .D(N179), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[127]) );
  EDFFX1 data_out_2_reg_126_ ( .D(N178), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[126]) );
  EDFFX1 data_out_2_reg_125_ ( .D(N177), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[125]) );
  EDFFX1 data_out_2_reg_110_ ( .D(N162), .E(n1167), .CK(clk), .Q(
        data_out_2[110]) );
  EDFFX1 data_out_2_reg_109_ ( .D(N161), .E(n1167), .CK(clk), .Q(
        data_out_2[109]) );
  EDFFX1 data_out_2_reg_108_ ( .D(N160), .E(n1167), .CK(clk), .Q(
        data_out_2[108]) );
  EDFFX1 data_out_2_reg_93_ ( .D(N145), .E(n1167), .CK(clk), .Q(data_out_2[93]) );
  EDFFX1 data_out_2_reg_92_ ( .D(N144), .E(n1167), .CK(clk), .Q(data_out_2[92]) );
  EDFFX1 data_out_2_reg_91_ ( .D(N143), .E(n1167), .CK(clk), .Q(data_out_2[91]) );
  EDFFX1 data_out_2_reg_77_ ( .D(N129), .E(n1166), .CK(clk), .Q(data_out_2[77]) );
  EDFFX1 data_out_2_reg_76_ ( .D(N128), .E(n1167), .CK(clk), .Q(data_out_2[76]) );
  EDFFX1 data_out_2_reg_75_ ( .D(N127), .E(n1166), .CK(clk), .Q(data_out_2[75]) );
  EDFFX1 data_out_2_reg_74_ ( .D(N126), .E(n1167), .CK(clk), .Q(data_out_2[74]) );
  EDFFX1 data_out_2_reg_59_ ( .D(N111), .E(n1166), .CK(clk), .Q(data_out_2[59]) );
  EDFFX1 data_out_2_reg_58_ ( .D(N110), .E(n1166), .CK(clk), .Q(data_out_2[58]) );
  EDFFX1 data_out_2_reg_57_ ( .D(N109), .E(n1166), .CK(clk), .Q(data_out_2[57]) );
  EDFFX1 data_out_2_reg_42_ ( .D(N94), .E(n1166), .CK(clk), .Q(data_out_2[42])
         );
  EDFFX1 data_out_2_reg_41_ ( .D(N93), .E(n1166), .CK(clk), .Q(data_out_2[41])
         );
  EDFFX1 data_out_2_reg_40_ ( .D(N92), .E(n1166), .CK(clk), .Q(data_out_2[40])
         );
  EDFFX1 data_out_2_reg_124_ ( .D(N176), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[124]) );
  EDFFX1 data_out_2_reg_123_ ( .D(N175), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[123]) );
  EDFFX1 data_out_2_reg_122_ ( .D(N174), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[122]) );
  EDFFX1 data_out_2_reg_107_ ( .D(N159), .E(n1167), .CK(clk), .Q(
        data_out_2[107]) );
  EDFFX1 data_out_2_reg_106_ ( .D(N158), .E(n1167), .CK(clk), .Q(
        data_out_2[106]) );
  EDFFX1 data_out_2_reg_105_ ( .D(N157), .E(n1167), .CK(clk), .Q(
        data_out_2[105]) );
  EDFFX1 data_out_2_reg_90_ ( .D(N142), .E(n1167), .CK(clk), .Q(data_out_2[90]) );
  EDFFX1 data_out_2_reg_89_ ( .D(N141), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[89]) );
  EDFFX1 data_out_2_reg_88_ ( .D(N140), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[88]) );
  EDFFX1 data_out_2_reg_73_ ( .D(N125), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[73]) );
  EDFFX1 data_out_2_reg_72_ ( .D(N124), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[72]) );
  EDFFX1 data_out_2_reg_71_ ( .D(N123), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[71]) );
  EDFFX1 data_out_2_reg_56_ ( .D(N108), .E(n1166), .CK(clk), .Q(data_out_2[56]) );
  EDFFX1 data_out_2_reg_55_ ( .D(N107), .E(n1166), .CK(clk), .Q(data_out_2[55]) );
  EDFFX1 data_out_2_reg_54_ ( .D(N106), .E(n1166), .CK(clk), .Q(data_out_2[54]) );
  EDFFX1 data_out_2_reg_39_ ( .D(N91), .E(n1166), .CK(clk), .Q(data_out_2[39])
         );
  EDFFX1 data_out_2_reg_38_ ( .D(N90), .E(n1166), .CK(clk), .Q(data_out_2[38])
         );
  EDFFX1 data_out_2_reg_37_ ( .D(N89), .E(n1166), .CK(clk), .Q(data_out_2[37])
         );
  EDFFX1 data_out_2_reg_70_ ( .D(N122), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[70]) );
  EDFFX1 data_out_2_reg_102_ ( .D(N154), .E(n1167), .CK(clk), .Q(
        data_out_2[102]) );
  EDFFX1 data_out_2_reg_68_ ( .D(N120), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[68]) );
  EDFFX1 data_out_2_reg_121_ ( .D(N173), .E(n1167), .CK(clk), .Q(
        data_out_2[121]) );
  EDFFX1 data_out_2_reg_103_ ( .D(N155), .E(n1167), .CK(clk), .Q(
        data_out_2[103]) );
  EDFFX1 data_out_2_reg_87_ ( .D(N139), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[87]) );
  EDFFX1 data_out_2_reg_119_ ( .D(N171), .E(n1167), .CK(clk), .Q(
        data_out_2[119]) );
  EDFFX1 data_out_2_reg_86_ ( .D(N138), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[86]) );
  EDFFX1 data_out_2_reg_120_ ( .D(N172), .E(n1167), .CK(clk), .Q(
        data_out_2[120]) );
  EDFFX1 data_out_2_reg_104_ ( .D(N156), .E(n1167), .CK(clk), .Q(
        data_out_2[104]) );
  EDFFX1 data_out_2_reg_53_ ( .D(N105), .E(n1166), .CK(clk), .Q(data_out_2[53]) );
  EDFFX1 data_out_2_reg_69_ ( .D(N121), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[69]) );
  EDFFX1 data_out_2_reg_36_ ( .D(N88), .E(n1166), .CK(clk), .Q(data_out_2[36])
         );
  EDFFX1 data_out_2_reg_35_ ( .D(N87), .E(n1166), .CK(clk), .Q(data_out_2[35])
         );
  EDFFX1 data_out_2_reg_101_ ( .D(N153), .E(n1167), .CK(clk), .Q(
        data_out_2[101]) );
  EDFFX1 data_out_2_reg_84_ ( .D(N136), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[84]) );
  EDFFX1 data_out_2_reg_34_ ( .D(N86), .E(n1166), .CK(clk), .Q(data_out_2[34])
         );
  EDFFX1 data_out_2_reg_118_ ( .D(N170), .E(n1167), .CK(clk), .Q(
        data_out_2[118]) );
  EDFFX1 data_out_2_reg_135_ ( .D(N187), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[135]) );
  EDFFXL R8_reg_28_ ( .D(data_in_2[28]), .E(n959), .CK(clk), .Q(R8[28]) );
  EDFFXL R8_reg_27_ ( .D(data_in_2[27]), .E(n959), .CK(clk), .Q(R8[27]) );
  EDFFXL R8_reg_11_ ( .D(data_in_2[11]), .E(n960), .CK(clk), .Q(R8[11]) );
  EDFFXL R8_reg_10_ ( .D(data_in_2[10]), .E(n960), .CK(clk), .Q(R8[10]) );
  EDFFXL R12_reg_28_ ( .D(data_in_2[28]), .E(n971), .CK(clk), .Q(R12[28]) );
  EDFFXL R12_reg_27_ ( .D(data_in_2[27]), .E(n1134), .CK(clk), .Q(R12[27]) );
  EDFFXL R12_reg_11_ ( .D(data_in_2[11]), .E(n1134), .CK(clk), .Q(R12[11]) );
  EDFFXL R12_reg_10_ ( .D(data_in_2[10]), .E(n1134), .CK(clk), .Q(R12[10]) );
  EDFFXL R0_reg_28_ ( .D(data_in_2[28]), .E(n1117), .CK(clk), .Q(R0[28]) );
  EDFFXL R0_reg_27_ ( .D(data_in_2[27]), .E(n1117), .CK(clk), .Q(R0[27]) );
  EDFFXL R0_reg_11_ ( .D(data_in_2[11]), .E(n1117), .CK(clk), .Q(R0[11]) );
  EDFFXL R0_reg_10_ ( .D(data_in_2[10]), .E(n1117), .CK(clk), .Q(R0[10]) );
  EDFFXL R4_reg_28_ ( .D(data_in_2[28]), .E(n969), .CK(clk), .Q(R4[28]) );
  EDFFXL R4_reg_27_ ( .D(data_in_2[27]), .E(n969), .CK(clk), .Q(R4[27]) );
  EDFFXL R4_reg_11_ ( .D(data_in_2[11]), .E(n969), .CK(clk), .Q(R4[11]) );
  EDFFXL R4_reg_10_ ( .D(data_in_2[10]), .E(n969), .CK(clk), .Q(R4[10]) );
  EDFFX1 R10_reg_26_ ( .D(data_in_2[94]), .E(n96), .CK(clk), .QN(n727) );
  EDFFX1 R10_reg_25_ ( .D(data_in_2[93]), .E(n960), .CK(clk), .QN(n728) );
  EDFFX1 R10_reg_24_ ( .D(data_in_2[92]), .E(n972), .CK(clk), .QN(n729) );
  EDFFX1 R10_reg_23_ ( .D(data_in_2[91]), .E(n968), .CK(clk), .QN(n730) );
  EDFFX1 R10_reg_11_ ( .D(data_in_2[79]), .E(n968), .CK(clk), .QN(n742) );
  EDFFX1 R10_reg_10_ ( .D(data_in_2[78]), .E(n970), .CK(clk), .QN(n743) );
  EDFFX1 R10_reg_9_ ( .D(data_in_2[77]), .E(n970), .CK(clk), .QN(n744) );
  EDFFX1 R10_reg_8_ ( .D(data_in_2[76]), .E(n970), .CK(clk), .QN(n745) );
  EDFFX1 R10_reg_7_ ( .D(data_in_2[75]), .E(n970), .CK(clk), .QN(n746) );
  EDFFX1 R10_reg_6_ ( .D(data_in_2[74]), .E(n970), .CK(clk), .QN(n747) );
  EDFFX1 R11_reg_28_ ( .D(data_in_2[130]), .E(n963), .CK(clk), .QN(n691) );
  EDFFX1 R11_reg_27_ ( .D(data_in_2[129]), .E(n963), .CK(clk), .QN(n692) );
  EDFFX1 R11_reg_26_ ( .D(data_in_2[128]), .E(n963), .CK(clk), .QN(n693) );
  EDFFX1 R11_reg_25_ ( .D(data_in_2[127]), .E(n963), .CK(clk), .QN(n694) );
  EDFFX1 R11_reg_24_ ( .D(data_in_2[126]), .E(n963), .CK(clk), .QN(n695) );
  EDFFX1 R11_reg_23_ ( .D(data_in_2[125]), .E(n963), .CK(clk), .QN(n696) );
  EDFFX1 R11_reg_11_ ( .D(data_in_2[113]), .E(n967), .CK(clk), .QN(n708) );
  EDFFX1 R11_reg_10_ ( .D(data_in_2[112]), .E(n967), .CK(clk), .QN(n709) );
  EDFFX1 R11_reg_9_ ( .D(data_in_2[111]), .E(n967), .CK(clk), .QN(n710) );
  EDFFX1 R11_reg_8_ ( .D(data_in_2[110]), .E(n967), .CK(clk), .QN(n711) );
  EDFFX1 R11_reg_7_ ( .D(data_in_2[109]), .E(n967), .CK(clk), .QN(n712) );
  EDFFX1 R11_reg_6_ ( .D(data_in_2[108]), .E(n967), .CK(clk), .QN(n713) );
  EDFFX1 data_out_2_reg_85_ ( .D(N137), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[85]) );
  EDFFX1 data_out_2_reg_51_ ( .D(N103), .E(n1166), .CK(clk), .Q(data_out_2[51]) );
  EDFFX1 data_out_2_reg_50_ ( .D(N102), .E(n1166), .CK(clk), .Q(data_out_2[50]) );
  EDFFX1 R5_reg_16_ ( .D(data_in_2[50]), .E(n1136), .CK(clk), .Q(R5[16]) );
  EDFFX1 R1_reg_16_ ( .D(data_in_2[50]), .E(n97), .CK(clk), .Q(R1[16]) );
  EDFFX1 R9_reg_16_ ( .D(data_in_2[50]), .E(n968), .CK(clk), .Q(R9[16]) );
  EDFFX1 R13_reg_16_ ( .D(data_in_2[50]), .E(n1129), .CK(clk), .Q(R13[16]) );
  EDFFXL R12_reg_32_ ( .D(data_in_2[32]), .E(n971), .CK(clk), .Q(R12[32]) );
  EDFFXL R8_reg_32_ ( .D(data_in_2[32]), .E(n96), .CK(clk), .Q(R8[32]) );
  EDFFXL R4_reg_32_ ( .D(data_in_2[32]), .E(n969), .CK(clk), .Q(R4[32]) );
  EDFFXL R0_reg_32_ ( .D(data_in_2[32]), .E(n97), .CK(clk), .Q(R0[32]) );
  EDFFXL data_out_2_reg_52_ ( .D(N104), .E(n1166), .CK(clk), .Q(data_out_2[52]) );
  EDFFXL data_out_2_reg_67_ ( .D(N119), .E(reg_flag_mux), .CK(clk), .Q(
        data_out_2[67]) );
  EDFFXL R12_reg_23_ ( .D(data_in_2[23]), .E(n971), .CK(clk), .Q(R12[23]) );
  EDFFXL R8_reg_23_ ( .D(data_in_2[23]), .E(n96), .CK(clk), .Q(R8[23]) );
  EDFFXL R4_reg_23_ ( .D(data_in_2[23]), .E(n969), .CK(clk), .Q(R4[23]) );
  EDFFXL R0_reg_23_ ( .D(data_in_2[23]), .E(n97), .CK(clk), .Q(R0[23]) );
  EDFFXL R12_reg_6_ ( .D(data_in_2[6]), .E(n971), .CK(clk), .Q(R12[6]) );
  EDFFXL R8_reg_6_ ( .D(data_in_2[6]), .E(n96), .CK(clk), .Q(R8[6]) );
  EDFFXL R4_reg_6_ ( .D(data_in_2[6]), .E(n969), .CK(clk), .Q(R4[6]) );
  EDFFXL R0_reg_6_ ( .D(data_in_2[6]), .E(n97), .CK(clk), .Q(R0[6]) );
  EDFFXL R12_reg_24_ ( .D(data_in_2[24]), .E(n971), .CK(clk), .Q(R12[24]) );
  EDFFXL R8_reg_24_ ( .D(data_in_2[24]), .E(n96), .CK(clk), .Q(R8[24]) );
  EDFFXL R4_reg_24_ ( .D(data_in_2[24]), .E(n969), .CK(clk), .Q(R4[24]) );
  EDFFXL R0_reg_24_ ( .D(data_in_2[24]), .E(n97), .CK(clk), .Q(R0[24]) );
  EDFFXL R12_reg_7_ ( .D(data_in_2[7]), .E(n971), .CK(clk), .Q(R12[7]) );
  EDFFXL R8_reg_7_ ( .D(data_in_2[7]), .E(n96), .CK(clk), .Q(R8[7]) );
  EDFFXL R4_reg_7_ ( .D(data_in_2[7]), .E(n969), .CK(clk), .Q(R4[7]) );
  EDFFXL R0_reg_7_ ( .D(data_in_2[7]), .E(n97), .CK(clk), .Q(R0[7]) );
  EDFFXL R12_reg_8_ ( .D(data_in_2[8]), .E(n971), .CK(clk), .Q(R12[8]) );
  EDFFXL R8_reg_8_ ( .D(data_in_2[8]), .E(n96), .CK(clk), .Q(R8[8]) );
  EDFFXL R4_reg_8_ ( .D(data_in_2[8]), .E(n969), .CK(clk), .Q(R4[8]) );
  EDFFXL R0_reg_8_ ( .D(data_in_2[8]), .E(n97), .CK(clk), .Q(R0[8]) );
  EDFFXL R12_reg_25_ ( .D(data_in_2[25]), .E(n971), .CK(clk), .Q(R12[25]) );
  EDFFXL R8_reg_25_ ( .D(data_in_2[25]), .E(n96), .CK(clk), .Q(R8[25]) );
  EDFFXL R4_reg_25_ ( .D(data_in_2[25]), .E(n969), .CK(clk), .Q(R4[25]) );
  EDFFXL R0_reg_25_ ( .D(data_in_2[25]), .E(n97), .CK(clk), .Q(R0[25]) );
  EDFFXL R12_reg_9_ ( .D(data_in_2[9]), .E(n971), .CK(clk), .Q(R12[9]) );
  EDFFXL R8_reg_9_ ( .D(data_in_2[9]), .E(n96), .CK(clk), .Q(R8[9]) );
  EDFFXL R4_reg_9_ ( .D(data_in_2[9]), .E(n969), .CK(clk), .Q(R4[9]) );
  EDFFXL R0_reg_9_ ( .D(data_in_2[9]), .E(n97), .CK(clk), .Q(R0[9]) );
  EDFFXL R12_reg_26_ ( .D(data_in_2[26]), .E(n971), .CK(clk), .Q(R12[26]) );
  EDFFXL R8_reg_26_ ( .D(data_in_2[26]), .E(n96), .CK(clk), .Q(R8[26]) );
  EDFFXL R4_reg_26_ ( .D(data_in_2[26]), .E(n969), .CK(clk), .Q(R4[26]) );
  EDFFXL R0_reg_26_ ( .D(data_in_2[26]), .E(n97), .CK(clk), .Q(R0[26]) );
  EDFFX1 R7_reg_16_ ( .D(data_in_2[118]), .E(n1138), .CK(clk), .QN(n941) );
  EDFFXL R12_reg_15_ ( .D(data_in_2[15]), .E(n1134), .CK(clk), .Q(R12[15]) );
  EDFFXL R0_reg_15_ ( .D(data_in_2[15]), .E(n1117), .CK(clk), .Q(R0[15]) );
  EDFFXL R8_reg_15_ ( .D(data_in_2[15]), .E(n960), .CK(clk), .Q(R8[15]) );
  EDFFXL R0_reg_16_ ( .D(data_in_2[16]), .E(n1117), .CK(clk), .Q(R0[16]) );
  EDFFXL R12_reg_16_ ( .D(data_in_2[16]), .E(n1134), .CK(clk), .Q(R12[16]) );
  EDFFXL R8_reg_16_ ( .D(data_in_2[16]), .E(n960), .CK(clk), .Q(R8[16]) );
  AND2X2 U3 ( .A(counter2[1]), .B(n1172), .Y(n8) );
  OR2X2 U4 ( .A(counter2[0]), .B(counter2[1]), .Y(n9) );
  OR2X2 U5 ( .A(n1172), .B(counter2[1]), .Y(n10) );
  AND2X2 U6 ( .A(counter2[1]), .B(counter2[0]), .Y(n11) );
  INVX1 U7 ( .A(n1139), .Y(n1137) );
  INVX1 U8 ( .A(n1139), .Y(n1136) );
  INVX1 U9 ( .A(n1139), .Y(n1138) );
  INVX1 U10 ( .A(n10), .Y(n1155) );
  INVX1 U11 ( .A(n10), .Y(n1156) );
  INVX1 U12 ( .A(n10), .Y(n1157) );
  INVX1 U13 ( .A(n10), .Y(n1150) );
  INVX1 U14 ( .A(n10), .Y(n1151) );
  INVX1 U15 ( .A(n10), .Y(n1152) );
  INVX1 U16 ( .A(n10), .Y(n1153) );
  INVX1 U17 ( .A(n10), .Y(n1154) );
  INVX1 U18 ( .A(n9), .Y(n1125) );
  INVX1 U19 ( .A(n9), .Y(n1126) );
  INVX1 U20 ( .A(n9), .Y(n1127) );
  INVX1 U21 ( .A(n9), .Y(n1119) );
  INVX1 U22 ( .A(n9), .Y(n1120) );
  INVX1 U23 ( .A(n9), .Y(n1121) );
  INVX1 U24 ( .A(n9), .Y(n1122) );
  INVX1 U25 ( .A(n9), .Y(n1123) );
  INVX1 U26 ( .A(n9), .Y(n1124) );
  INVX1 U27 ( .A(n8), .Y(n1147) );
  INVX1 U28 ( .A(n8), .Y(n1148) );
  INVX1 U29 ( .A(n8), .Y(n1149) );
  INVX1 U30 ( .A(n8), .Y(n1140) );
  INVX1 U31 ( .A(n8), .Y(n1141) );
  INVX1 U32 ( .A(n8), .Y(n1142) );
  INVX1 U33 ( .A(n8), .Y(n1143) );
  INVX1 U34 ( .A(n8), .Y(n1144) );
  INVX1 U35 ( .A(n8), .Y(n1145) );
  INVX1 U36 ( .A(n8), .Y(n1146) );
  INVX1 U37 ( .A(n1135), .Y(n1128) );
  INVX1 U38 ( .A(n1135), .Y(n1129) );
  INVX1 U39 ( .A(n1135), .Y(n1131) );
  INVX1 U40 ( .A(n1135), .Y(n1132) );
  INVX1 U41 ( .A(n977), .Y(n972) );
  INVX1 U42 ( .A(n977), .Y(n970) );
  INVX1 U43 ( .A(n977), .Y(n968) );
  INVX1 U44 ( .A(n977), .Y(n967) );
  INVX1 U45 ( .A(n977), .Y(n963) );
  INVX1 U46 ( .A(n1135), .Y(n1133) );
  INVX1 U47 ( .A(n1135), .Y(n1130) );
  INVX1 U48 ( .A(n977), .Y(n960) );
  INVX1 U49 ( .A(n977), .Y(n959) );
  INVX1 U50 ( .A(n1135), .Y(n1134) );
  INVX1 U51 ( .A(n969), .Y(n1139) );
  INVX1 U52 ( .A(n11), .Y(n1158) );
  INVX1 U53 ( .A(n11), .Y(n1160) );
  INVX1 U54 ( .A(n11), .Y(n1159) );
  INVX1 U55 ( .A(n11), .Y(n1165) );
  INVX1 U56 ( .A(n11), .Y(n1164) );
  INVX1 U57 ( .A(n11), .Y(n1163) );
  INVX1 U58 ( .A(n11), .Y(n1162) );
  INVX1 U59 ( .A(n11), .Y(n1161) );
  INVX1 U60 ( .A(n966), .Y(n1173) );
  NOR2X1 U61 ( .A(n1171), .B(n1170), .Y(n964) );
  NOR2X1 U62 ( .A(n973), .B(n1171), .Y(n969) );
  INVX1 U63 ( .A(n96), .Y(n977) );
  INVX1 U64 ( .A(n971), .Y(n1135) );
  INVX1 U65 ( .A(n1118), .Y(n1117) );
  INVX1 U66 ( .A(n97), .Y(n1118) );
  INVX1 U67 ( .A(n1168), .Y(n1166) );
  INVX1 U68 ( .A(n1168), .Y(n1167) );
  NOR2X1 U69 ( .A(n961), .B(reg_flag_mux), .Y(n966) );
  OAI2BB2X1 U70 ( .B0(n965), .B1(n961), .A0N(counter2[1]), .A1N(n966), .Y(
        n1113) );
  AOI21X1 U71 ( .A0(n1150), .A1(n1173), .B0(n8), .Y(n965) );
  INVX1 U72 ( .A(n962), .Y(n1169) );
  AOI32X1 U73 ( .A0(reg_flag_mux), .A1(n1158), .A2(rst_n), .B0(n964), .B1(
        rst_n), .Y(n962) );
  OAI32X1 U74 ( .A0(n961), .A1(counter2[0]), .A2(n966), .B0(n1172), .B1(n1173), 
        .Y(n1114) );
  OAI22X1 U75 ( .A0(n1170), .A1(n974), .B0(n961), .B1(n973), .Y(n1116) );
  NAND2BX1 U76 ( .AN(reg_datain_flag), .B(rst_n), .Y(n974) );
  OAI21XL U77 ( .A0(n1171), .A1(n974), .B0(n975), .Y(n1115) );
  OAI21XL U78 ( .A0(n1117), .A1(n969), .B0(rst_n), .Y(n975) );
  OAI221XL U79 ( .A0(n889), .A1(n1160), .B0(n855), .B1(n1149), .C0(n1024), .Y(
        N52) );
  AOI22X1 U80 ( .A0(R1[0]), .A1(n1152), .B0(n1120), .B1(R0[0]), .Y(n1024) );
  OAI221XL U81 ( .A0(n888), .A1(n1159), .B0(n854), .B1(n1144), .C0(n1023), .Y(
        N53) );
  AOI22X1 U82 ( .A0(R1[1]), .A1(n1153), .B0(n1121), .B1(R0[1]), .Y(n1023) );
  OAI221XL U83 ( .A0(n887), .A1(n1163), .B0(n853), .B1(n1145), .C0(n1022), .Y(
        N54) );
  AOI22X1 U84 ( .A0(R1[2]), .A1(n1154), .B0(n1127), .B1(R0[2]), .Y(n1022) );
  OAI221XL U85 ( .A0(n886), .A1(n1158), .B0(n852), .B1(n1147), .C0(n1021), .Y(
        N55) );
  AOI22X1 U86 ( .A0(R1[3]), .A1(n1155), .B0(n1121), .B1(R0[3]), .Y(n1021) );
  OAI221XL U87 ( .A0(n885), .A1(n1161), .B0(n851), .B1(n1146), .C0(n1020), .Y(
        N56) );
  AOI22X1 U88 ( .A0(R1[4]), .A1(n1155), .B0(n1127), .B1(R0[4]), .Y(n1020) );
  OAI221XL U89 ( .A0(n884), .A1(n1164), .B0(n850), .B1(n1148), .C0(n1019), .Y(
        N57) );
  AOI22X1 U90 ( .A0(R1[5]), .A1(n1155), .B0(n1125), .B1(R0[5]), .Y(n1019) );
  OAI221XL U91 ( .A0(n883), .A1(n1160), .B0(n849), .B1(n1140), .C0(n1018), .Y(
        N58) );
  AOI22X1 U92 ( .A0(R1[6]), .A1(n1155), .B0(n1119), .B1(R0[6]), .Y(n1018) );
  OAI221XL U93 ( .A0(n882), .A1(n1159), .B0(n848), .B1(n1149), .C0(n1017), .Y(
        N59) );
  AOI22X1 U94 ( .A0(R1[7]), .A1(n1155), .B0(n1123), .B1(R0[7]), .Y(n1017) );
  OAI221XL U95 ( .A0(n881), .A1(n1163), .B0(n847), .B1(n1147), .C0(n1016), .Y(
        N60) );
  AOI22X1 U96 ( .A0(R1[8]), .A1(n1155), .B0(n1125), .B1(R0[8]), .Y(n1016) );
  OAI221XL U97 ( .A0(n880), .A1(n1165), .B0(n846), .B1(n1147), .C0(n1015), .Y(
        N61) );
  AOI22X1 U98 ( .A0(R1[9]), .A1(n1155), .B0(n1125), .B1(R0[9]), .Y(n1015) );
  OAI221XL U99 ( .A0(n879), .A1(n1160), .B0(n845), .B1(n1147), .C0(n1014), .Y(
        N62) );
  AOI22X1 U100 ( .A0(R1[10]), .A1(n1155), .B0(n1125), .B1(R0[10]), .Y(n1014)
         );
  OAI221XL U101 ( .A0(n878), .A1(n1160), .B0(n844), .B1(n1147), .C0(n1013), 
        .Y(N63) );
  AOI22X1 U102 ( .A0(R1[11]), .A1(n1155), .B0(n1125), .B1(R0[11]), .Y(n1013)
         );
  OAI221XL U103 ( .A0(n877), .A1(n1160), .B0(n843), .B1(n1147), .C0(n1012), 
        .Y(N64) );
  AOI22X1 U104 ( .A0(R1[12]), .A1(n1155), .B0(n1125), .B1(R0[12]), .Y(n1012)
         );
  OAI221XL U105 ( .A0(n876), .A1(n1160), .B0(n842), .B1(n1147), .C0(n1011), 
        .Y(N65) );
  AOI22X1 U106 ( .A0(R1[13]), .A1(n1155), .B0(n1125), .B1(R0[13]), .Y(n1011)
         );
  OAI221XL U107 ( .A0(n875), .A1(n1160), .B0(n841), .B1(n1147), .C0(n1010), 
        .Y(N66) );
  AOI22X1 U108 ( .A0(R1[14]), .A1(n1155), .B0(n1125), .B1(R0[14]), .Y(n1010)
         );
  OAI221XL U109 ( .A0(n874), .A1(n1160), .B0(n840), .B1(n1147), .C0(n1009), 
        .Y(N67) );
  AOI22X1 U110 ( .A0(R1[15]), .A1(n1155), .B0(n1125), .B1(R0[15]), .Y(n1009)
         );
  OAI221XL U111 ( .A0(n873), .A1(n1160), .B0(n839), .B1(n1147), .C0(n1008), 
        .Y(N68) );
  AOI22X1 U112 ( .A0(R1[16]), .A1(n1156), .B0(n1125), .B1(R0[16]), .Y(n1008)
         );
  OAI221XL U113 ( .A0(n872), .A1(n1160), .B0(n838), .B1(n1147), .C0(n1007), 
        .Y(N69) );
  AOI22X1 U114 ( .A0(R1[17]), .A1(n1156), .B0(n1125), .B1(R0[17]), .Y(n1007)
         );
  OAI221XL U115 ( .A0(n871), .A1(n1160), .B0(n837), .B1(n1147), .C0(n1006), 
        .Y(N70) );
  AOI22X1 U116 ( .A0(R1[18]), .A1(n1156), .B0(n1125), .B1(R0[18]), .Y(n1006)
         );
  OAI221XL U117 ( .A0(n870), .A1(n1160), .B0(n836), .B1(n1147), .C0(n1005), 
        .Y(N71) );
  AOI22X1 U118 ( .A0(R1[19]), .A1(n1156), .B0(n1125), .B1(R0[19]), .Y(n1005)
         );
  OAI221XL U119 ( .A0(n869), .A1(n1160), .B0(n835), .B1(n1148), .C0(n1004), 
        .Y(N72) );
  AOI22X1 U120 ( .A0(R1[20]), .A1(n1156), .B0(n1126), .B1(R0[20]), .Y(n1004)
         );
  OAI221XL U121 ( .A0(n868), .A1(n1160), .B0(n834), .B1(n1148), .C0(n1003), 
        .Y(N73) );
  AOI22X1 U122 ( .A0(R1[21]), .A1(n1156), .B0(n1126), .B1(R0[21]), .Y(n1003)
         );
  OAI221XL U123 ( .A0(n867), .A1(n1160), .B0(n833), .B1(n1148), .C0(n1002), 
        .Y(N74) );
  AOI22X1 U124 ( .A0(R1[22]), .A1(n1156), .B0(n1126), .B1(R0[22]), .Y(n1002)
         );
  OAI221XL U125 ( .A0(n866), .A1(n1159), .B0(n832), .B1(n1148), .C0(n1001), 
        .Y(N75) );
  AOI22X1 U126 ( .A0(R1[23]), .A1(n1156), .B0(n1126), .B1(R0[23]), .Y(n1001)
         );
  OAI221XL U127 ( .A0(n865), .A1(n1159), .B0(n831), .B1(n1148), .C0(n1000), 
        .Y(N76) );
  AOI22X1 U128 ( .A0(R1[24]), .A1(n1156), .B0(n1126), .B1(R0[24]), .Y(n1000)
         );
  OAI221XL U129 ( .A0(n864), .A1(n1159), .B0(n830), .B1(n1148), .C0(n999), .Y(
        N77) );
  AOI22X1 U130 ( .A0(R1[25]), .A1(n1156), .B0(n1126), .B1(R0[25]), .Y(n999) );
  OAI221XL U131 ( .A0(n863), .A1(n1159), .B0(n829), .B1(n1148), .C0(n998), .Y(
        N78) );
  AOI22X1 U132 ( .A0(R1[26]), .A1(n1156), .B0(n1126), .B1(R0[26]), .Y(n998) );
  OAI221XL U133 ( .A0(n862), .A1(n1159), .B0(n828), .B1(n1148), .C0(n997), .Y(
        N79) );
  AOI22X1 U134 ( .A0(R1[27]), .A1(n1156), .B0(n1126), .B1(R0[27]), .Y(n997) );
  OAI221XL U135 ( .A0(n861), .A1(n1159), .B0(n827), .B1(n1148), .C0(n996), .Y(
        N80) );
  AOI22X1 U136 ( .A0(R1[28]), .A1(n1156), .B0(n1126), .B1(R0[28]), .Y(n996) );
  OAI221XL U137 ( .A0(n860), .A1(n1159), .B0(n826), .B1(n1148), .C0(n995), .Y(
        N81) );
  AOI22X1 U138 ( .A0(R1[29]), .A1(n1157), .B0(n1126), .B1(R0[29]), .Y(n995) );
  OAI221XL U139 ( .A0(n859), .A1(n1159), .B0(n825), .B1(n1148), .C0(n994), .Y(
        N82) );
  AOI22X1 U140 ( .A0(R1[30]), .A1(n1157), .B0(n1126), .B1(R0[30]), .Y(n994) );
  OAI221XL U141 ( .A0(n858), .A1(n1159), .B0(n824), .B1(n1148), .C0(n993), .Y(
        N83) );
  AOI22X1 U142 ( .A0(R1[31]), .A1(n1157), .B0(n1126), .B1(R0[31]), .Y(n993) );
  OAI221XL U143 ( .A0(n857), .A1(n1159), .B0(n823), .B1(n1149), .C0(n992), .Y(
        N84) );
  AOI22X1 U144 ( .A0(R1[32]), .A1(n1157), .B0(n1127), .B1(R0[32]), .Y(n992) );
  OAI221XL U145 ( .A0(n856), .A1(n1159), .B0(n822), .B1(n1149), .C0(n991), .Y(
        N85) );
  AOI22X1 U146 ( .A0(R1[33]), .A1(n1157), .B0(n1127), .B1(R0[33]), .Y(n991) );
  OAI221XL U147 ( .A0(n957), .A1(n1159), .B0(n923), .B1(n1149), .C0(n990), .Y(
        N86) );
  AOI22X1 U148 ( .A0(R5[0]), .A1(n1157), .B0(n1127), .B1(R4[0]), .Y(n990) );
  OAI221XL U149 ( .A0(n956), .A1(n1159), .B0(n922), .B1(n1149), .C0(n989), .Y(
        N87) );
  AOI22X1 U150 ( .A0(R5[1]), .A1(n1157), .B0(n1127), .B1(R4[1]), .Y(n989) );
  OAI221XL U151 ( .A0(n955), .A1(n1158), .B0(n921), .B1(n1149), .C0(n988), .Y(
        N88) );
  AOI22X1 U152 ( .A0(R5[2]), .A1(n1157), .B0(n1127), .B1(R4[2]), .Y(n988) );
  OAI221XL U153 ( .A0(n954), .A1(n1158), .B0(n920), .B1(n1149), .C0(n987), .Y(
        N89) );
  AOI22X1 U154 ( .A0(R5[3]), .A1(n1157), .B0(n1127), .B1(R4[3]), .Y(n987) );
  OAI221XL U155 ( .A0(n953), .A1(n1158), .B0(n919), .B1(n1149), .C0(n986), .Y(
        N90) );
  AOI22X1 U156 ( .A0(R5[4]), .A1(n1157), .B0(n1127), .B1(R4[4]), .Y(n986) );
  OAI221XL U157 ( .A0(n952), .A1(n1158), .B0(n918), .B1(n1149), .C0(n985), .Y(
        N91) );
  AOI22X1 U158 ( .A0(R5[5]), .A1(n1157), .B0(n1127), .B1(R4[5]), .Y(n985) );
  OAI221XL U159 ( .A0(n951), .A1(n1158), .B0(n917), .B1(n1149), .C0(n984), .Y(
        N92) );
  AOI22X1 U160 ( .A0(R5[6]), .A1(n1157), .B0(n1127), .B1(R4[6]), .Y(n984) );
  OAI221XL U161 ( .A0(n950), .A1(n1158), .B0(n916), .B1(n1149), .C0(n983), .Y(
        N93) );
  AOI22X1 U162 ( .A0(R5[7]), .A1(n1157), .B0(n1127), .B1(R4[7]), .Y(n983) );
  OAI221XL U163 ( .A0(n949), .A1(n1158), .B0(n915), .B1(n1149), .C0(n982), .Y(
        N94) );
  AOI22X1 U164 ( .A0(R5[8]), .A1(n1152), .B0(n1127), .B1(R4[8]), .Y(n982) );
  OAI221XL U165 ( .A0(n948), .A1(n1158), .B0(n914), .B1(n1149), .C0(n981), .Y(
        N95) );
  AOI22X1 U166 ( .A0(R5[9]), .A1(n1153), .B0(n1127), .B1(R4[9]), .Y(n981) );
  OAI221XL U167 ( .A0(n947), .A1(n1158), .B0(n913), .B1(n1141), .C0(n980), .Y(
        N96) );
  AOI22X1 U168 ( .A0(R5[10]), .A1(n1156), .B0(n1126), .B1(R4[10]), .Y(n980) );
  OAI221XL U169 ( .A0(n946), .A1(n1158), .B0(n912), .B1(n1142), .C0(n979), .Y(
        N97) );
  AOI22X1 U170 ( .A0(R5[11]), .A1(n1156), .B0(n1124), .B1(R4[11]), .Y(n979) );
  OAI221XL U171 ( .A0(n945), .A1(n1158), .B0(n911), .B1(n1143), .C0(n978), .Y(
        N98) );
  AOI22X1 U172 ( .A0(R5[12]), .A1(n1154), .B0(n1122), .B1(R4[12]), .Y(n978) );
  OAI221XL U173 ( .A0(n944), .A1(n1158), .B0(n910), .B1(n1141), .C0(n976), .Y(
        N99) );
  AOI22X1 U174 ( .A0(R5[13]), .A1(n1151), .B0(n1126), .B1(R4[13]), .Y(n976) );
  OAI221XL U175 ( .A0(n943), .A1(n1165), .B0(n909), .B1(n1140), .C0(n1112), 
        .Y(N100) );
  AOI22X1 U176 ( .A0(R5[14]), .A1(n1157), .B0(n1119), .B1(R4[14]), .Y(n1112)
         );
  OAI221XL U177 ( .A0(n942), .A1(n1164), .B0(n908), .B1(n1140), .C0(n1111), 
        .Y(N101) );
  AOI22X1 U178 ( .A0(R5[15]), .A1(n1155), .B0(n1119), .B1(R4[15]), .Y(n1111)
         );
  OAI221XL U179 ( .A0(n941), .A1(n1161), .B0(n907), .B1(n1140), .C0(n1110), 
        .Y(N102) );
  AOI22X1 U180 ( .A0(R5[16]), .A1(n1157), .B0(n1119), .B1(R4[16]), .Y(n1110)
         );
  OAI221XL U181 ( .A0(n940), .A1(n1160), .B0(n906), .B1(n1140), .C0(n1109), 
        .Y(N103) );
  AOI22X1 U182 ( .A0(R5[17]), .A1(n1155), .B0(n1119), .B1(R4[17]), .Y(n1109)
         );
  OAI221XL U183 ( .A0(n939), .A1(n1163), .B0(n905), .B1(n1140), .C0(n1108), 
        .Y(N104) );
  AOI22X1 U184 ( .A0(R5[18]), .A1(n1155), .B0(n1119), .B1(R4[18]), .Y(n1108)
         );
  OAI221XL U185 ( .A0(n938), .A1(n1164), .B0(n904), .B1(n1140), .C0(n1107), 
        .Y(N105) );
  AOI22X1 U186 ( .A0(R5[19]), .A1(n1153), .B0(n1119), .B1(R4[19]), .Y(n1107)
         );
  OAI221XL U187 ( .A0(n937), .A1(n1159), .B0(n903), .B1(n1140), .C0(n1106), 
        .Y(N106) );
  AOI22X1 U188 ( .A0(R5[20]), .A1(n1150), .B0(n1119), .B1(R4[20]), .Y(n1106)
         );
  OAI221XL U189 ( .A0(n936), .A1(n1165), .B0(n902), .B1(n1140), .C0(n1105), 
        .Y(N107) );
  AOI22X1 U190 ( .A0(R5[21]), .A1(n1150), .B0(n1119), .B1(R4[21]), .Y(n1105)
         );
  OAI221XL U191 ( .A0(n935), .A1(n1165), .B0(n901), .B1(n1140), .C0(n1104), 
        .Y(N108) );
  AOI22X1 U192 ( .A0(R5[22]), .A1(n1154), .B0(n1119), .B1(R4[22]), .Y(n1104)
         );
  OAI221XL U193 ( .A0(n934), .A1(n1165), .B0(n900), .B1(n1140), .C0(n1103), 
        .Y(N109) );
  AOI22X1 U194 ( .A0(R5[23]), .A1(n1156), .B0(n1119), .B1(R4[23]), .Y(n1103)
         );
  OAI221XL U195 ( .A0(n933), .A1(n1165), .B0(n899), .B1(n1140), .C0(n1102), 
        .Y(N110) );
  AOI22X1 U196 ( .A0(R5[24]), .A1(n1151), .B0(n1119), .B1(R4[24]), .Y(n1102)
         );
  OAI221XL U197 ( .A0(n932), .A1(n1165), .B0(n898), .B1(n1140), .C0(n1101), 
        .Y(N111) );
  AOI22X1 U198 ( .A0(R5[25]), .A1(n1152), .B0(n1119), .B1(R4[25]), .Y(n1101)
         );
  OAI221XL U199 ( .A0(n931), .A1(n1165), .B0(n897), .B1(n1141), .C0(n1100), 
        .Y(N112) );
  AOI22X1 U200 ( .A0(R5[26]), .A1(n1157), .B0(n1120), .B1(R4[26]), .Y(n1100)
         );
  OAI221XL U201 ( .A0(n930), .A1(n1165), .B0(n896), .B1(n1141), .C0(n1099), 
        .Y(N113) );
  AOI22X1 U202 ( .A0(R5[27]), .A1(n1150), .B0(n1120), .B1(R4[27]), .Y(n1099)
         );
  OAI221XL U203 ( .A0(n929), .A1(n1165), .B0(n895), .B1(n1141), .C0(n1098), 
        .Y(N114) );
  AOI22X1 U204 ( .A0(R5[28]), .A1(n1150), .B0(n1120), .B1(R4[28]), .Y(n1098)
         );
  OAI221XL U205 ( .A0(n928), .A1(n1165), .B0(n894), .B1(n1141), .C0(n1097), 
        .Y(N115) );
  AOI22X1 U206 ( .A0(R5[29]), .A1(n1150), .B0(n1120), .B1(R4[29]), .Y(n1097)
         );
  OAI221XL U207 ( .A0(n927), .A1(n1165), .B0(n893), .B1(n1141), .C0(n1096), 
        .Y(N116) );
  AOI22X1 U208 ( .A0(R5[30]), .A1(n1150), .B0(n1120), .B1(R4[30]), .Y(n1096)
         );
  OAI221XL U209 ( .A0(n926), .A1(n1165), .B0(n892), .B1(n1141), .C0(n1095), 
        .Y(N117) );
  AOI22X1 U210 ( .A0(R5[31]), .A1(n1150), .B0(n1120), .B1(R4[31]), .Y(n1095)
         );
  OAI221XL U211 ( .A0(n925), .A1(n1165), .B0(n891), .B1(n1141), .C0(n1094), 
        .Y(N118) );
  AOI22X1 U212 ( .A0(R5[32]), .A1(n1150), .B0(n1120), .B1(R4[32]), .Y(n1094)
         );
  OAI221XL U213 ( .A0(n924), .A1(n1165), .B0(n890), .B1(n1141), .C0(n1093), 
        .Y(N119) );
  AOI22X1 U214 ( .A0(R5[33]), .A1(n1150), .B0(n1120), .B1(R4[33]), .Y(n1093)
         );
  OAI221XL U215 ( .A0(n719), .A1(n1164), .B0(n753), .B1(n1141), .C0(n1092), 
        .Y(N120) );
  AOI22X1 U216 ( .A0(R9[0]), .A1(n1150), .B0(n1120), .B1(R8[0]), .Y(n1092) );
  OAI221XL U217 ( .A0(n718), .A1(n1164), .B0(n752), .B1(n1141), .C0(n1091), 
        .Y(N121) );
  AOI22X1 U218 ( .A0(R9[1]), .A1(n1150), .B0(n1120), .B1(R8[1]), .Y(n1091) );
  OAI221XL U219 ( .A0(n717), .A1(n1164), .B0(n751), .B1(n1141), .C0(n1090), 
        .Y(N122) );
  AOI22X1 U220 ( .A0(R9[2]), .A1(n1150), .B0(n1120), .B1(R8[2]), .Y(n1090) );
  OAI221XL U221 ( .A0(n716), .A1(n1164), .B0(n750), .B1(n1141), .C0(n1089), 
        .Y(N123) );
  AOI22X1 U222 ( .A0(R9[3]), .A1(n1150), .B0(n1120), .B1(R8[3]), .Y(n1089) );
  OAI221XL U223 ( .A0(n715), .A1(n1164), .B0(n749), .B1(n1142), .C0(n1088), 
        .Y(N124) );
  AOI22X1 U224 ( .A0(R9[4]), .A1(n1150), .B0(n1121), .B1(R8[4]), .Y(n1088) );
  OAI221XL U225 ( .A0(n714), .A1(n1164), .B0(n748), .B1(n1142), .C0(n1087), 
        .Y(N125) );
  AOI22X1 U226 ( .A0(R9[5]), .A1(n1150), .B0(n1121), .B1(R8[5]), .Y(n1087) );
  OAI221XL U227 ( .A0(n713), .A1(n1164), .B0(n747), .B1(n1142), .C0(n1086), 
        .Y(N126) );
  AOI22X1 U228 ( .A0(R9[6]), .A1(n1151), .B0(n1121), .B1(R8[6]), .Y(n1086) );
  OAI221XL U229 ( .A0(n712), .A1(n1164), .B0(n746), .B1(n1142), .C0(n1085), 
        .Y(N127) );
  AOI22X1 U230 ( .A0(R9[7]), .A1(n1151), .B0(n1121), .B1(R8[7]), .Y(n1085) );
  OAI221XL U231 ( .A0(n711), .A1(n1164), .B0(n745), .B1(n1142), .C0(n1084), 
        .Y(N128) );
  AOI22X1 U232 ( .A0(R9[8]), .A1(n1151), .B0(n1121), .B1(R8[8]), .Y(n1084) );
  OAI221XL U233 ( .A0(n710), .A1(n1164), .B0(n744), .B1(n1142), .C0(n1083), 
        .Y(N129) );
  AOI22X1 U234 ( .A0(R9[9]), .A1(n1151), .B0(n1121), .B1(R8[9]), .Y(n1083) );
  OAI221XL U235 ( .A0(n709), .A1(n1164), .B0(n743), .B1(n1142), .C0(n1082), 
        .Y(N130) );
  AOI22X1 U236 ( .A0(R9[10]), .A1(n1151), .B0(n1121), .B1(R8[10]), .Y(n1082)
         );
  OAI221XL U237 ( .A0(n708), .A1(n1164), .B0(n742), .B1(n1142), .C0(n1081), 
        .Y(N131) );
  AOI22X1 U238 ( .A0(R9[11]), .A1(n1151), .B0(n1121), .B1(R8[11]), .Y(n1081)
         );
  OAI221XL U239 ( .A0(n707), .A1(n1164), .B0(n741), .B1(n1142), .C0(n1080), 
        .Y(N132) );
  AOI22X1 U240 ( .A0(R9[12]), .A1(n1151), .B0(n1121), .B1(R8[12]), .Y(n1080)
         );
  OAI221XL U241 ( .A0(n706), .A1(n1163), .B0(n740), .B1(n1142), .C0(n1079), 
        .Y(N133) );
  AOI22X1 U242 ( .A0(R9[13]), .A1(n1151), .B0(n1121), .B1(R8[13]), .Y(n1079)
         );
  OAI221XL U243 ( .A0(n705), .A1(n1163), .B0(n739), .B1(n1142), .C0(n1078), 
        .Y(N134) );
  AOI22X1 U244 ( .A0(R9[14]), .A1(n1151), .B0(n1121), .B1(R8[14]), .Y(n1078)
         );
  OAI221XL U245 ( .A0(n704), .A1(n1163), .B0(n738), .B1(n1142), .C0(n1077), 
        .Y(N135) );
  AOI22X1 U246 ( .A0(R9[15]), .A1(n1151), .B0(n1121), .B1(R8[15]), .Y(n1077)
         );
  OAI221XL U247 ( .A0(n703), .A1(n1163), .B0(n737), .B1(n1143), .C0(n1076), 
        .Y(N136) );
  AOI22X1 U248 ( .A0(R9[16]), .A1(n1151), .B0(n1122), .B1(R8[16]), .Y(n1076)
         );
  OAI221XL U249 ( .A0(n702), .A1(n1163), .B0(n736), .B1(n1143), .C0(n1075), 
        .Y(N137) );
  AOI22X1 U250 ( .A0(R9[17]), .A1(n1151), .B0(n1122), .B1(R8[17]), .Y(n1075)
         );
  OAI221XL U251 ( .A0(n701), .A1(n1163), .B0(n735), .B1(n1143), .C0(n1074), 
        .Y(N138) );
  AOI22X1 U252 ( .A0(R9[18]), .A1(n1151), .B0(n1122), .B1(R8[18]), .Y(n1074)
         );
  OAI221XL U253 ( .A0(n700), .A1(n1163), .B0(n734), .B1(n1143), .C0(n1073), 
        .Y(N139) );
  AOI22X1 U254 ( .A0(R9[19]), .A1(n1152), .B0(n1122), .B1(R8[19]), .Y(n1073)
         );
  OAI221XL U255 ( .A0(n699), .A1(n1163), .B0(n733), .B1(n1143), .C0(n1072), 
        .Y(N140) );
  AOI22X1 U256 ( .A0(R9[20]), .A1(n1152), .B0(n1122), .B1(R8[20]), .Y(n1072)
         );
  OAI221XL U257 ( .A0(n698), .A1(n1163), .B0(n732), .B1(n1143), .C0(n1071), 
        .Y(N141) );
  AOI22X1 U258 ( .A0(R9[21]), .A1(n1152), .B0(n1122), .B1(R8[21]), .Y(n1071)
         );
  OAI221XL U259 ( .A0(n697), .A1(n1163), .B0(n731), .B1(n1143), .C0(n1070), 
        .Y(N142) );
  AOI22X1 U260 ( .A0(R9[22]), .A1(n1152), .B0(n1122), .B1(R8[22]), .Y(n1070)
         );
  OAI221XL U261 ( .A0(n696), .A1(n1163), .B0(n730), .B1(n1143), .C0(n1069), 
        .Y(N143) );
  AOI22X1 U262 ( .A0(R9[23]), .A1(n1152), .B0(n1122), .B1(R8[23]), .Y(n1069)
         );
  OAI221XL U263 ( .A0(n695), .A1(n1163), .B0(n729), .B1(n1143), .C0(n1068), 
        .Y(N144) );
  AOI22X1 U264 ( .A0(R9[24]), .A1(n1152), .B0(n1122), .B1(R8[24]), .Y(n1068)
         );
  OAI221XL U265 ( .A0(n694), .A1(n1163), .B0(n728), .B1(n1143), .C0(n1067), 
        .Y(N145) );
  AOI22X1 U266 ( .A0(R9[25]), .A1(n1152), .B0(n1122), .B1(R8[25]), .Y(n1067)
         );
  OAI221XL U267 ( .A0(n693), .A1(n1162), .B0(n727), .B1(n1143), .C0(n1066), 
        .Y(N146) );
  AOI22X1 U268 ( .A0(R9[26]), .A1(n1152), .B0(n1122), .B1(R8[26]), .Y(n1066)
         );
  OAI221XL U269 ( .A0(n692), .A1(n1162), .B0(n726), .B1(n1143), .C0(n1065), 
        .Y(N147) );
  AOI22X1 U270 ( .A0(R9[27]), .A1(n1152), .B0(n1122), .B1(R8[27]), .Y(n1065)
         );
  OAI221XL U271 ( .A0(n691), .A1(n1162), .B0(n725), .B1(n1144), .C0(n1064), 
        .Y(N148) );
  AOI22X1 U272 ( .A0(R9[28]), .A1(n1152), .B0(n1123), .B1(R8[28]), .Y(n1064)
         );
  OAI221XL U273 ( .A0(n690), .A1(n1162), .B0(n724), .B1(n1144), .C0(n1063), 
        .Y(N149) );
  AOI22X1 U274 ( .A0(R9[29]), .A1(n1152), .B0(n1123), .B1(R8[29]), .Y(n1063)
         );
  OAI221XL U275 ( .A0(n689), .A1(n1162), .B0(n723), .B1(n1144), .C0(n1062), 
        .Y(N150) );
  AOI22X1 U276 ( .A0(R9[30]), .A1(n1152), .B0(n1123), .B1(R8[30]), .Y(n1062)
         );
  OAI221XL U277 ( .A0(n688), .A1(n1162), .B0(n722), .B1(n1144), .C0(n1061), 
        .Y(N151) );
  AOI22X1 U278 ( .A0(R9[31]), .A1(n1152), .B0(n1123), .B1(R8[31]), .Y(n1061)
         );
  OAI221XL U279 ( .A0(n687), .A1(n1162), .B0(n721), .B1(n1144), .C0(n1060), 
        .Y(N152) );
  AOI22X1 U280 ( .A0(R9[32]), .A1(n1153), .B0(n1123), .B1(R8[32]), .Y(n1060)
         );
  OAI221XL U281 ( .A0(n686), .A1(n1162), .B0(n720), .B1(n1144), .C0(n1059), 
        .Y(N153) );
  AOI22X1 U282 ( .A0(R9[33]), .A1(n1153), .B0(n1123), .B1(R8[33]), .Y(n1059)
         );
  OAI221XL U283 ( .A0(n821), .A1(n1162), .B0(n787), .B1(n1144), .C0(n1058), 
        .Y(N154) );
  AOI22X1 U284 ( .A0(R13[0]), .A1(n1153), .B0(n1123), .B1(R12[0]), .Y(n1058)
         );
  OAI221XL U285 ( .A0(n820), .A1(n1162), .B0(n786), .B1(n1144), .C0(n1057), 
        .Y(N155) );
  AOI22X1 U286 ( .A0(R13[1]), .A1(n1153), .B0(n1123), .B1(R12[1]), .Y(n1057)
         );
  OAI221XL U287 ( .A0(n819), .A1(n1162), .B0(n785), .B1(n1144), .C0(n1056), 
        .Y(N156) );
  AOI22X1 U288 ( .A0(R13[2]), .A1(n1153), .B0(n1123), .B1(R12[2]), .Y(n1056)
         );
  OAI221XL U289 ( .A0(n818), .A1(n1162), .B0(n784), .B1(n1144), .C0(n1055), 
        .Y(N157) );
  AOI22X1 U290 ( .A0(R13[3]), .A1(n1153), .B0(n1123), .B1(R12[3]), .Y(n1055)
         );
  OAI221XL U291 ( .A0(n817), .A1(n1162), .B0(n783), .B1(n1144), .C0(n1054), 
        .Y(N158) );
  AOI22X1 U292 ( .A0(R13[4]), .A1(n1153), .B0(n1123), .B1(R12[4]), .Y(n1054)
         );
  OAI221XL U293 ( .A0(n816), .A1(n1162), .B0(n782), .B1(n1144), .C0(n1053), 
        .Y(N159) );
  AOI22X1 U294 ( .A0(R13[5]), .A1(n1153), .B0(n1123), .B1(R12[5]), .Y(n1053)
         );
  OAI221XL U295 ( .A0(n815), .A1(n1158), .B0(n781), .B1(n1145), .C0(n1052), 
        .Y(N160) );
  AOI22X1 U296 ( .A0(R13[6]), .A1(n1153), .B0(n1122), .B1(R12[6]), .Y(n1052)
         );
  OAI221XL U297 ( .A0(n814), .A1(n1162), .B0(n780), .B1(n1145), .C0(n1051), 
        .Y(N161) );
  AOI22X1 U298 ( .A0(R13[7]), .A1(n1153), .B0(n1124), .B1(R12[7]), .Y(n1051)
         );
  OAI221XL U299 ( .A0(n813), .A1(n1165), .B0(n779), .B1(n1145), .C0(n1050), 
        .Y(N162) );
  AOI22X1 U300 ( .A0(R13[8]), .A1(n1153), .B0(n1126), .B1(R12[8]), .Y(n1050)
         );
  OAI221XL U301 ( .A0(n812), .A1(n1164), .B0(n778), .B1(n1145), .C0(n1049), 
        .Y(N163) );
  AOI22X1 U303 ( .A0(R13[9]), .A1(n1153), .B0(n1121), .B1(R12[9]), .Y(n1049)
         );
  OAI221XL U304 ( .A0(n811), .A1(n1163), .B0(n777), .B1(n1145), .C0(n1048), 
        .Y(N164) );
  AOI22X1 U305 ( .A0(R13[10]), .A1(n1153), .B0(n1127), .B1(R12[10]), .Y(n1048)
         );
  OAI221XL U306 ( .A0(n810), .A1(n1161), .B0(n776), .B1(n1145), .C0(n1047), 
        .Y(N165) );
  AOI22X1 U307 ( .A0(R13[11]), .A1(n1154), .B0(n1123), .B1(R12[11]), .Y(n1047)
         );
  OAI221XL U308 ( .A0(n809), .A1(n1160), .B0(n775), .B1(n1145), .C0(n1046), 
        .Y(N166) );
  AOI22X1 U309 ( .A0(R13[12]), .A1(n1154), .B0(n1119), .B1(R12[12]), .Y(n1046)
         );
  OAI221XL U310 ( .A0(n808), .A1(n1161), .B0(n774), .B1(n1145), .C0(n1045), 
        .Y(N167) );
  AOI22X1 U311 ( .A0(R13[13]), .A1(n1154), .B0(n1120), .B1(R12[13]), .Y(n1045)
         );
  OAI221XL U312 ( .A0(n807), .A1(n1159), .B0(n773), .B1(n1145), .C0(n1044), 
        .Y(N168) );
  AOI22X1 U313 ( .A0(R13[14]), .A1(n1154), .B0(n1124), .B1(R12[14]), .Y(n1044)
         );
  OAI221XL U314 ( .A0(n806), .A1(n1158), .B0(n772), .B1(n1145), .C0(n1043), 
        .Y(N169) );
  OAI221XL U315 ( .A0(n805), .A1(n1162), .B0(n771), .B1(n1145), .C0(n1042), 
        .Y(N170) );
  AOI22X1 U316 ( .A0(R13[16]), .A1(n1154), .B0(n1122), .B1(R12[16]), .Y(n1042)
         );
  OAI221XL U317 ( .A0(n804), .A1(n1165), .B0(n770), .B1(n1145), .C0(n1041), 
        .Y(N171) );
  AOI22X1 U318 ( .A0(R13[17]), .A1(n1154), .B0(n1124), .B1(R12[17]), .Y(n1041)
         );
  OAI221XL U319 ( .A0(n803), .A1(n1161), .B0(n769), .B1(n1146), .C0(n1040), 
        .Y(N172) );
  AOI22X1 U320 ( .A0(R13[18]), .A1(n1154), .B0(n1124), .B1(R12[18]), .Y(n1040)
         );
  OAI221XL U321 ( .A0(n802), .A1(n1161), .B0(n768), .B1(n1146), .C0(n1039), 
        .Y(N173) );
  AOI22X1 U322 ( .A0(R13[19]), .A1(n1154), .B0(n1124), .B1(R12[19]), .Y(n1039)
         );
  OAI221XL U323 ( .A0(n801), .A1(n1161), .B0(n767), .B1(n1146), .C0(n1038), 
        .Y(N174) );
  AOI22X1 U324 ( .A0(R13[20]), .A1(n1154), .B0(n1124), .B1(R12[20]), .Y(n1038)
         );
  OAI221XL U325 ( .A0(n800), .A1(n1161), .B0(n766), .B1(n1146), .C0(n1037), 
        .Y(N175) );
  AOI22X1 U326 ( .A0(R13[21]), .A1(n1154), .B0(n1124), .B1(R12[21]), .Y(n1037)
         );
  OAI221XL U327 ( .A0(n799), .A1(n1161), .B0(n765), .B1(n1146), .C0(n1036), 
        .Y(N176) );
  AOI22X1 U328 ( .A0(R13[22]), .A1(n1154), .B0(n1124), .B1(R12[22]), .Y(n1036)
         );
  OAI221XL U329 ( .A0(n798), .A1(n1161), .B0(n764), .B1(n1146), .C0(n1035), 
        .Y(N177) );
  AOI22X1 U330 ( .A0(R13[23]), .A1(n1154), .B0(n1124), .B1(R12[23]), .Y(n1035)
         );
  OAI221XL U331 ( .A0(n797), .A1(n1161), .B0(n763), .B1(n1146), .C0(n1034), 
        .Y(N178) );
  AOI22X1 U332 ( .A0(R13[24]), .A1(n1151), .B0(n1124), .B1(R12[24]), .Y(n1034)
         );
  OAI221XL U333 ( .A0(n796), .A1(n1161), .B0(n762), .B1(n1146), .C0(n1033), 
        .Y(N179) );
  AOI22X1 U334 ( .A0(R13[25]), .A1(n1150), .B0(n1124), .B1(R12[25]), .Y(n1033)
         );
  OAI221XL U335 ( .A0(n795), .A1(n1161), .B0(n761), .B1(n1146), .C0(n1032), 
        .Y(N180) );
  AOI22X1 U336 ( .A0(R13[26]), .A1(n1156), .B0(n1124), .B1(R12[26]), .Y(n1032)
         );
  OAI221XL U337 ( .A0(n794), .A1(n1161), .B0(n760), .B1(n1146), .C0(n1031), 
        .Y(N181) );
  AOI22X1 U338 ( .A0(R13[27]), .A1(n1152), .B0(n1124), .B1(R12[27]), .Y(n1031)
         );
  OAI221XL U339 ( .A0(n793), .A1(n1161), .B0(n759), .B1(n1146), .C0(n1030), 
        .Y(N182) );
  AOI22X1 U340 ( .A0(R13[28]), .A1(n1153), .B0(n1124), .B1(R12[28]), .Y(n1030)
         );
  OAI221XL U341 ( .A0(n792), .A1(n1161), .B0(n758), .B1(n1146), .C0(n1029), 
        .Y(N183) );
  AOI22X1 U342 ( .A0(R13[29]), .A1(n1154), .B0(n1124), .B1(R12[29]), .Y(n1029)
         );
  OAI221XL U343 ( .A0(n791), .A1(n1161), .B0(n757), .B1(n1144), .C0(n1028), 
        .Y(N184) );
  AOI22X1 U344 ( .A0(R13[30]), .A1(n1151), .B0(n1125), .B1(R12[30]), .Y(n1028)
         );
  OAI221XL U345 ( .A0(n790), .A1(n1162), .B0(n756), .B1(n1145), .C0(n1027), 
        .Y(N185) );
  AOI22X1 U346 ( .A0(R13[31]), .A1(n1155), .B0(n1119), .B1(R12[31]), .Y(n1027)
         );
  OAI221XL U347 ( .A0(n789), .A1(n1158), .B0(n755), .B1(n1147), .C0(n1026), 
        .Y(N186) );
  AOI22X1 U348 ( .A0(R13[32]), .A1(n1157), .B0(n1123), .B1(R12[32]), .Y(n1026)
         );
  OAI221XL U349 ( .A0(n788), .A1(n1161), .B0(n754), .B1(n1146), .C0(n1025), 
        .Y(N187) );
  AOI22X1 U350 ( .A0(R13[33]), .A1(n1150), .B0(n1120), .B1(R12[33]), .Y(n1025)
         );
  NOR2X1 U351 ( .A(n973), .B(counter1[1]), .Y(n971) );
  NAND2X1 U352 ( .A(reg_datain_flag), .B(n1170), .Y(n973) );
  INVX1 U353 ( .A(counter1[1]), .Y(n1171) );
  INVX1 U354 ( .A(counter1[0]), .Y(n1170) );
  AND2X2 U355 ( .A(reg_datain_flag), .B(n964), .Y(n96) );
  INVX1 U356 ( .A(counter2[0]), .Y(n1172) );
  AND3X2 U357 ( .A(counter1[0]), .B(n1171), .C(reg_datain_flag), .Y(n97) );
  INVX1 U358 ( .A(reg_flag_mux), .Y(n1168) );
  AOI22X1 U359 ( .A0(R13[15]), .A1(n1154), .B0(n1125), .B1(R12[15]), .Y(n1043)
         );
endmodule


module p_s ( clk, rst_n, data_in_3, p_s_flag_in, data_out_3 );
  input [135:0] data_in_3;
  output [33:0] data_out_3;
  input clk, rst_n, p_s_flag_in;
  wire   N26, N50, N52, N119, N120, N121, N122, N123, N124, N125, N126, N127,
         N128, N129, N130, N131, N132, N133, N134, N135, N136, N137, N138,
         N139, N140, N141, N142, N143, N144, N145, N146, N147, N148, N149,
         N150, N151, N152, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n862, n864, n865, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n880, n885, n890, n895, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
         n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
         n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
         n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
         n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
         n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
         n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
         n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
         n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
         n1160, n1161, n1162, n1163, n1164, n1165, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n125, n126, n887, n888,
         n889, n891, n892, n893, n894, n896, n1166, n1167, n1168, n1169, n1170,
         n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
         n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
         n1191, n1192, n1193, n1194, n1195;
  wire   [1:0] counter_1;
  wire   [33:0] R0;
  wire   [33:0] R12;
  wire   [33:0] R1;
  wire   [33:0] R13;
  wire   [33:0] R2;
  wire   [33:0] R14;
  wire   [33:0] R3;
  wire   [33:0] R15;
  wire   [3:0] counter_2;

  EDFFXL R1_reg_33_ ( .D(data_in_3[33]), .E(n1166), .CK(clk), .Q(R1[33]) );
  EDFFXL R0_reg_33_ ( .D(data_in_3[33]), .E(n887), .CK(clk), .Q(R0[33]) );
  EDFFXL R3_reg_33_ ( .D(data_in_3[33]), .E(n865), .CK(clk), .Q(R3[33]) );
  EDFFXL R2_reg_33_ ( .D(data_in_3[33]), .E(n1188), .CK(clk), .Q(R2[33]) );
  EDFFXL R1_reg_14_ ( .D(data_in_3[14]), .E(n1167), .CK(clk), .Q(R1[14]) );
  EDFFXL R0_reg_14_ ( .D(data_in_3[14]), .E(n888), .CK(clk), .Q(R0[14]) );
  EDFFXL R3_reg_14_ ( .D(data_in_3[14]), .E(n1180), .CK(clk), .Q(R3[14]) );
  EDFFXL R2_reg_14_ ( .D(data_in_3[14]), .E(n1188), .CK(clk), .Q(R2[14]) );
  EDFFXL R13_reg_33_ ( .D(data_in_3[135]), .E(n125), .CK(clk), .Q(R13[33]) );
  EDFFXL R12_reg_33_ ( .D(data_in_3[135]), .E(n892), .CK(clk), .Q(R12[33]) );
  EDFFXL R15_reg_33_ ( .D(data_in_3[135]), .E(n1176), .CK(clk), .Q(R15[33]) );
  EDFFXL R14_reg_33_ ( .D(data_in_3[135]), .E(n1187), .CK(clk), .Q(R14[33]) );
  EDFFX1 R7_reg_31_ ( .D(data_in_3[65]), .E(n1179), .CK(clk), .QN(n588) );
  EDFFX1 R7_reg_30_ ( .D(data_in_3[64]), .E(n1181), .CK(clk), .QN(n589) );
  EDFFX1 R7_reg_29_ ( .D(data_in_3[63]), .E(n1179), .CK(clk), .QN(n590) );
  EDFFX1 R7_reg_22_ ( .D(data_in_3[56]), .E(n865), .CK(clk), .QN(n597) );
  EDFFX1 R7_reg_21_ ( .D(data_in_3[55]), .E(n865), .CK(clk), .QN(n598) );
  EDFFX1 R7_reg_20_ ( .D(data_in_3[54]), .E(n1177), .CK(clk), .QN(n599) );
  EDFFX1 R7_reg_19_ ( .D(data_in_3[53]), .E(n1175), .CK(clk), .QN(n600) );
  EDFFX1 R7_reg_18_ ( .D(data_in_3[52]), .E(n1178), .CK(clk), .QN(n601) );
  EDFFX1 R7_reg_17_ ( .D(data_in_3[51]), .E(n1179), .CK(clk), .QN(n602) );
  EDFFX1 R7_reg_16_ ( .D(data_in_3[50]), .E(n1178), .CK(clk), .QN(n603) );
  EDFFX1 R7_reg_15_ ( .D(data_in_3[49]), .E(n1179), .CK(clk), .QN(n604) );
  EDFFX1 R7_reg_14_ ( .D(data_in_3[48]), .E(n1181), .CK(clk), .QN(n605) );
  EDFFX1 R7_reg_13_ ( .D(data_in_3[47]), .E(n1181), .CK(clk), .QN(n606) );
  EDFFX1 R7_reg_12_ ( .D(data_in_3[46]), .E(n1181), .CK(clk), .QN(n607) );
  EDFFX1 R7_reg_5_ ( .D(data_in_3[39]), .E(n1181), .CK(clk), .QN(n614) );
  EDFFX1 R7_reg_4_ ( .D(data_in_3[38]), .E(n1181), .CK(clk), .QN(n615) );
  EDFFX1 R7_reg_3_ ( .D(data_in_3[37]), .E(n1181), .CK(clk), .QN(n616) );
  EDFFX1 R7_reg_2_ ( .D(data_in_3[36]), .E(n1181), .CK(clk), .QN(n617) );
  EDFFX1 R7_reg_1_ ( .D(data_in_3[35]), .E(n1179), .CK(clk), .QN(n618) );
  EDFFX1 R7_reg_0_ ( .D(data_in_3[34]), .E(n1180), .CK(clk), .QN(n619) );
  EDFFX1 R6_reg_31_ ( .D(data_in_3[65]), .E(n864), .CK(clk), .QN(n656) );
  EDFFX1 R6_reg_30_ ( .D(data_in_3[64]), .E(n864), .CK(clk), .QN(n657) );
  EDFFX1 R6_reg_29_ ( .D(data_in_3[63]), .E(n1184), .CK(clk), .QN(n658) );
  EDFFX1 R6_reg_28_ ( .D(data_in_3[62]), .E(n1186), .CK(clk), .QN(n659) );
  EDFFX1 R6_reg_27_ ( .D(data_in_3[61]), .E(n1187), .CK(clk), .QN(n660) );
  EDFFX1 R6_reg_26_ ( .D(data_in_3[60]), .E(n1185), .CK(clk), .QN(n661) );
  EDFFX1 R6_reg_25_ ( .D(data_in_3[59]), .E(n1188), .CK(clk), .QN(n662) );
  EDFFX1 R6_reg_24_ ( .D(data_in_3[58]), .E(n1187), .CK(clk), .QN(n663) );
  EDFFX1 R6_reg_23_ ( .D(data_in_3[57]), .E(n1189), .CK(clk), .QN(n664) );
  EDFFX1 R6_reg_22_ ( .D(data_in_3[56]), .E(n1183), .CK(clk), .QN(n665) );
  EDFFX1 R6_reg_21_ ( .D(data_in_3[55]), .E(n1184), .CK(clk), .QN(n666) );
  EDFFX1 R6_reg_20_ ( .D(data_in_3[54]), .E(n1186), .CK(clk), .QN(n667) );
  EDFFX1 R6_reg_19_ ( .D(data_in_3[53]), .E(n1187), .CK(clk), .QN(n668) );
  EDFFX1 R6_reg_18_ ( .D(data_in_3[52]), .E(n1189), .CK(clk), .QN(n669) );
  EDFFX1 R6_reg_17_ ( .D(data_in_3[51]), .E(n1183), .CK(clk), .QN(n670) );
  EDFFX1 R6_reg_16_ ( .D(data_in_3[50]), .E(n1185), .CK(clk), .QN(n671) );
  EDFFX1 R6_reg_15_ ( .D(data_in_3[49]), .E(n1185), .CK(clk), .QN(n672) );
  EDFFX1 R6_reg_14_ ( .D(data_in_3[48]), .E(n1188), .CK(clk), .QN(n673) );
  EDFFX1 R6_reg_13_ ( .D(data_in_3[47]), .E(n1185), .CK(clk), .QN(n674) );
  EDFFX1 R6_reg_12_ ( .D(data_in_3[46]), .E(n1183), .CK(clk), .QN(n675) );
  EDFFX1 R6_reg_11_ ( .D(data_in_3[45]), .E(n1183), .CK(clk), .QN(n676) );
  EDFFX1 R6_reg_10_ ( .D(data_in_3[44]), .E(n1183), .CK(clk), .QN(n677) );
  EDFFX1 R6_reg_9_ ( .D(data_in_3[43]), .E(n1183), .CK(clk), .QN(n678) );
  EDFFX1 R6_reg_8_ ( .D(data_in_3[42]), .E(n1183), .CK(clk), .QN(n679) );
  EDFFX1 R6_reg_7_ ( .D(data_in_3[41]), .E(n1183), .CK(clk), .QN(n680) );
  EDFFX1 R6_reg_6_ ( .D(data_in_3[40]), .E(n1183), .CK(clk), .QN(n681) );
  EDFFX1 R6_reg_5_ ( .D(data_in_3[39]), .E(n1183), .CK(clk), .QN(n682) );
  EDFFX1 R6_reg_4_ ( .D(data_in_3[38]), .E(n1183), .CK(clk), .QN(n683) );
  EDFFX1 R6_reg_3_ ( .D(data_in_3[37]), .E(n1183), .CK(clk), .QN(n684) );
  EDFFX1 R6_reg_2_ ( .D(data_in_3[36]), .E(n1183), .CK(clk), .QN(n685) );
  EDFFX1 R6_reg_1_ ( .D(data_in_3[35]), .E(n1183), .CK(clk), .QN(n686) );
  EDFFX1 R6_reg_0_ ( .D(data_in_3[34]), .E(n1183), .CK(clk), .QN(n687) );
  EDFFX1 R4_reg_31_ ( .D(data_in_3[65]), .E(n126), .CK(clk), .QN(n724) );
  EDFFX1 R4_reg_30_ ( .D(data_in_3[64]), .E(n126), .CK(clk), .QN(n725) );
  EDFFX1 R4_reg_29_ ( .D(data_in_3[63]), .E(n126), .CK(clk), .QN(n726) );
  EDFFX1 R4_reg_28_ ( .D(data_in_3[62]), .E(n126), .CK(clk), .QN(n727) );
  EDFFX1 R4_reg_27_ ( .D(data_in_3[61]), .E(n126), .CK(clk), .QN(n728) );
  EDFFX1 R4_reg_26_ ( .D(data_in_3[60]), .E(n126), .CK(clk), .QN(n729) );
  EDFFX1 R4_reg_25_ ( .D(data_in_3[59]), .E(n126), .CK(clk), .QN(n730) );
  EDFFX1 R4_reg_24_ ( .D(data_in_3[58]), .E(n126), .CK(clk), .QN(n731) );
  EDFFX1 R4_reg_23_ ( .D(data_in_3[57]), .E(n126), .CK(clk), .QN(n732) );
  EDFFX1 R4_reg_22_ ( .D(data_in_3[56]), .E(n126), .CK(clk), .QN(n733) );
  EDFFX1 R4_reg_21_ ( .D(data_in_3[55]), .E(n893), .CK(clk), .QN(n734) );
  EDFFX1 R4_reg_20_ ( .D(data_in_3[54]), .E(n892), .CK(clk), .QN(n735) );
  EDFFX1 R4_reg_19_ ( .D(data_in_3[53]), .E(n887), .CK(clk), .QN(n736) );
  EDFFX1 R4_reg_18_ ( .D(data_in_3[52]), .E(n891), .CK(clk), .QN(n737) );
  EDFFX1 R4_reg_17_ ( .D(data_in_3[51]), .E(n889), .CK(clk), .QN(n738) );
  EDFFX1 R4_reg_16_ ( .D(data_in_3[50]), .E(n888), .CK(clk), .QN(n739) );
  EDFFX1 R4_reg_15_ ( .D(data_in_3[49]), .E(n889), .CK(clk), .QN(n740) );
  EDFFX1 R4_reg_14_ ( .D(data_in_3[48]), .E(n889), .CK(clk), .QN(n741) );
  EDFFX1 R4_reg_13_ ( .D(data_in_3[47]), .E(n889), .CK(clk), .QN(n742) );
  EDFFX1 R4_reg_12_ ( .D(data_in_3[46]), .E(n889), .CK(clk), .QN(n743) );
  EDFFX1 R4_reg_11_ ( .D(data_in_3[45]), .E(n889), .CK(clk), .QN(n744) );
  EDFFX1 R4_reg_10_ ( .D(data_in_3[44]), .E(n889), .CK(clk), .QN(n745) );
  EDFFX1 R4_reg_9_ ( .D(data_in_3[43]), .E(n889), .CK(clk), .QN(n746) );
  EDFFX1 R4_reg_8_ ( .D(data_in_3[42]), .E(n889), .CK(clk), .QN(n747) );
  EDFFX1 R4_reg_7_ ( .D(data_in_3[41]), .E(n889), .CK(clk), .QN(n748) );
  EDFFX1 R4_reg_6_ ( .D(data_in_3[40]), .E(n889), .CK(clk), .QN(n749) );
  EDFFX1 R4_reg_5_ ( .D(data_in_3[39]), .E(n889), .CK(clk), .QN(n750) );
  EDFFX1 R4_reg_4_ ( .D(data_in_3[38]), .E(n889), .CK(clk), .QN(n751) );
  EDFFX1 R4_reg_3_ ( .D(data_in_3[37]), .E(n889), .CK(clk), .QN(n752) );
  EDFFX1 R4_reg_2_ ( .D(data_in_3[36]), .E(n891), .CK(clk), .QN(n753) );
  EDFFX1 R4_reg_1_ ( .D(data_in_3[35]), .E(n891), .CK(clk), .QN(n754) );
  EDFFX1 R4_reg_0_ ( .D(data_in_3[34]), .E(n891), .CK(clk), .QN(n755) );
  EDFFXL R5_reg_33_ ( .D(data_in_3[67]), .E(n125), .CK(clk), .QN(n790) );
  EDFFXL R5_reg_32_ ( .D(data_in_3[66]), .E(n125), .CK(clk), .QN(n791) );
  EDFFXL R5_reg_31_ ( .D(data_in_3[65]), .E(n125), .CK(clk), .QN(n792) );
  EDFFXL R5_reg_30_ ( .D(data_in_3[64]), .E(n125), .CK(clk), .QN(n793) );
  EDFFXL R5_reg_29_ ( .D(data_in_3[63]), .E(n125), .CK(clk), .QN(n794) );
  EDFFX1 R5_reg_28_ ( .D(data_in_3[62]), .E(n1168), .CK(clk), .QN(n795) );
  EDFFX1 R5_reg_27_ ( .D(data_in_3[61]), .E(n1168), .CK(clk), .QN(n796) );
  EDFFX1 R5_reg_26_ ( .D(data_in_3[60]), .E(n1168), .CK(clk), .QN(n797) );
  EDFFX1 R5_reg_25_ ( .D(data_in_3[59]), .E(n1168), .CK(clk), .QN(n798) );
  EDFFX1 R5_reg_24_ ( .D(data_in_3[58]), .E(n1168), .CK(clk), .QN(n799) );
  EDFFX1 R5_reg_23_ ( .D(data_in_3[57]), .E(n1168), .CK(clk), .QN(n800) );
  EDFFX1 R5_reg_22_ ( .D(data_in_3[56]), .E(n1168), .CK(clk), .QN(n801) );
  EDFFX1 R5_reg_21_ ( .D(data_in_3[55]), .E(n1168), .CK(clk), .QN(n802) );
  EDFFX1 R5_reg_20_ ( .D(data_in_3[54]), .E(n1168), .CK(clk), .QN(n803) );
  EDFFX1 R5_reg_19_ ( .D(data_in_3[53]), .E(n1168), .CK(clk), .QN(n804) );
  EDFFX1 R5_reg_18_ ( .D(data_in_3[52]), .E(n1168), .CK(clk), .QN(n805) );
  EDFFX1 R5_reg_17_ ( .D(data_in_3[51]), .E(n1168), .CK(clk), .QN(n806) );
  EDFFXL R5_reg_15_ ( .D(data_in_3[49]), .E(n1169), .CK(clk), .QN(n808) );
  EDFFXL R5_reg_14_ ( .D(data_in_3[48]), .E(n1169), .CK(clk), .QN(n809) );
  EDFFXL R5_reg_13_ ( .D(data_in_3[47]), .E(n1169), .CK(clk), .QN(n810) );
  EDFFXL R5_reg_12_ ( .D(data_in_3[46]), .E(n1169), .CK(clk), .QN(n811) );
  EDFFX1 R5_reg_11_ ( .D(data_in_3[45]), .E(n1169), .CK(clk), .QN(n812) );
  EDFFX1 R5_reg_10_ ( .D(data_in_3[44]), .E(n1169), .CK(clk), .QN(n813) );
  EDFFX1 R5_reg_9_ ( .D(data_in_3[43]), .E(n1169), .CK(clk), .QN(n814) );
  EDFFX1 R5_reg_8_ ( .D(data_in_3[42]), .E(n1169), .CK(clk), .QN(n815) );
  EDFFX1 R5_reg_7_ ( .D(data_in_3[41]), .E(n1169), .CK(clk), .QN(n816) );
  EDFFX1 R5_reg_6_ ( .D(data_in_3[40]), .E(n1169), .CK(clk), .QN(n817) );
  EDFFX1 R5_reg_5_ ( .D(data_in_3[39]), .E(n1169), .CK(clk), .QN(n818) );
  EDFFX1 R5_reg_4_ ( .D(data_in_3[38]), .E(n1169), .CK(clk), .QN(n819) );
  EDFFX1 R5_reg_3_ ( .D(data_in_3[37]), .E(n1169), .CK(clk), .QN(n820) );
  EDFFX1 R5_reg_2_ ( .D(data_in_3[36]), .E(n1170), .CK(clk), .QN(n821) );
  EDFFX1 R5_reg_1_ ( .D(data_in_3[35]), .E(n1170), .CK(clk), .QN(n822) );
  EDFFX1 R5_reg_0_ ( .D(data_in_3[34]), .E(n1170), .CK(clk), .QN(n823) );
  EDFFXL R10_reg_33_ ( .D(data_in_3[101]), .E(n1189), .CK(clk), .QN(n620) );
  EDFFXL R10_reg_32_ ( .D(data_in_3[100]), .E(n1183), .CK(clk), .QN(n621) );
  EDFFXL R10_reg_31_ ( .D(data_in_3[99]), .E(n1184), .CK(clk), .QN(n622) );
  EDFFXL R10_reg_30_ ( .D(data_in_3[98]), .E(n1185), .CK(clk), .QN(n623) );
  EDFFXL R10_reg_29_ ( .D(data_in_3[97]), .E(n1185), .CK(clk), .QN(n624) );
  EDFFXL R10_reg_28_ ( .D(data_in_3[96]), .E(n1185), .CK(clk), .QN(n625) );
  EDFFXL R10_reg_27_ ( .D(data_in_3[95]), .E(n1185), .CK(clk), .QN(n626) );
  EDFFX1 R10_reg_26_ ( .D(data_in_3[94]), .E(n1185), .CK(clk), .QN(n627) );
  EDFFX1 R10_reg_25_ ( .D(data_in_3[93]), .E(n1185), .CK(clk), .QN(n628) );
  EDFFX1 R10_reg_24_ ( .D(data_in_3[92]), .E(n1185), .CK(clk), .QN(n629) );
  EDFFX1 R10_reg_23_ ( .D(data_in_3[91]), .E(n1185), .CK(clk), .QN(n630) );
  EDFFX1 R10_reg_22_ ( .D(data_in_3[90]), .E(n1185), .CK(clk), .QN(n631) );
  EDFFX1 R10_reg_21_ ( .D(data_in_3[89]), .E(n1185), .CK(clk), .QN(n632) );
  EDFFX1 R10_reg_20_ ( .D(data_in_3[88]), .E(n1185), .CK(clk), .QN(n633) );
  EDFFX1 R10_reg_19_ ( .D(data_in_3[87]), .E(n1185), .CK(clk), .QN(n634) );
  EDFFX1 R10_reg_18_ ( .D(data_in_3[86]), .E(n1185), .CK(clk), .QN(n635) );
  EDFFX1 R10_reg_17_ ( .D(data_in_3[85]), .E(n1184), .CK(clk), .QN(n636) );
  EDFFXL R10_reg_16_ ( .D(data_in_3[84]), .E(n1184), .CK(clk), .QN(n637) );
  EDFFXL R10_reg_15_ ( .D(data_in_3[83]), .E(n1184), .CK(clk), .QN(n638) );
  EDFFXL R10_reg_14_ ( .D(data_in_3[82]), .E(n1184), .CK(clk), .QN(n639) );
  EDFFXL R10_reg_13_ ( .D(data_in_3[81]), .E(n1184), .CK(clk), .QN(n640) );
  EDFFXL R10_reg_12_ ( .D(data_in_3[80]), .E(n1184), .CK(clk), .QN(n641) );
  EDFFX1 R10_reg_11_ ( .D(data_in_3[79]), .E(n1184), .CK(clk), .QN(n642) );
  EDFFX1 R10_reg_10_ ( .D(data_in_3[78]), .E(n1184), .CK(clk), .QN(n643) );
  EDFFX1 R10_reg_9_ ( .D(data_in_3[77]), .E(n1184), .CK(clk), .QN(n644) );
  EDFFX1 R10_reg_8_ ( .D(data_in_3[76]), .E(n1184), .CK(clk), .QN(n645) );
  EDFFX1 R10_reg_7_ ( .D(data_in_3[75]), .E(n1184), .CK(clk), .QN(n646) );
  EDFFX1 R10_reg_6_ ( .D(data_in_3[74]), .E(n1184), .CK(clk), .QN(n647) );
  EDFFX1 R10_reg_5_ ( .D(data_in_3[73]), .E(n1184), .CK(clk), .QN(n648) );
  EDFFX1 R10_reg_4_ ( .D(data_in_3[72]), .E(n1188), .CK(clk), .QN(n649) );
  EDFFX1 R10_reg_3_ ( .D(data_in_3[71]), .E(n1189), .CK(clk), .QN(n650) );
  EDFFX1 R10_reg_2_ ( .D(data_in_3[70]), .E(n1183), .CK(clk), .QN(n651) );
  EDFFX1 R10_reg_1_ ( .D(data_in_3[69]), .E(n1184), .CK(clk), .QN(n652) );
  EDFFX1 R10_reg_0_ ( .D(data_in_3[68]), .E(n1186), .CK(clk), .QN(n653) );
  EDFFXL R11_reg_33_ ( .D(data_in_3[101]), .E(n1179), .CK(clk), .QN(n688) );
  EDFFXL R11_reg_32_ ( .D(data_in_3[100]), .E(n1179), .CK(clk), .QN(n689) );
  EDFFXL R11_reg_31_ ( .D(data_in_3[99]), .E(n1179), .CK(clk), .QN(n690) );
  EDFFXL R11_reg_30_ ( .D(data_in_3[98]), .E(n1178), .CK(clk), .QN(n691) );
  EDFFXL R11_reg_29_ ( .D(data_in_3[97]), .E(n1178), .CK(clk), .QN(n692) );
  EDFFXL R11_reg_28_ ( .D(data_in_3[96]), .E(n1178), .CK(clk), .QN(n693) );
  EDFFXL R11_reg_27_ ( .D(data_in_3[95]), .E(n1178), .CK(clk), .QN(n694) );
  EDFFX1 R11_reg_26_ ( .D(data_in_3[94]), .E(n1178), .CK(clk), .QN(n695) );
  EDFFX1 R11_reg_25_ ( .D(data_in_3[93]), .E(n1178), .CK(clk), .QN(n696) );
  EDFFX1 R11_reg_24_ ( .D(data_in_3[92]), .E(n1178), .CK(clk), .QN(n697) );
  EDFFX1 R11_reg_23_ ( .D(data_in_3[91]), .E(n1178), .CK(clk), .QN(n698) );
  EDFFX1 R11_reg_22_ ( .D(data_in_3[90]), .E(n1178), .CK(clk), .QN(n699) );
  EDFFX1 R11_reg_21_ ( .D(data_in_3[89]), .E(n1178), .CK(clk), .QN(n700) );
  EDFFX1 R11_reg_20_ ( .D(data_in_3[88]), .E(n1178), .CK(clk), .QN(n701) );
  EDFFX1 R11_reg_19_ ( .D(data_in_3[87]), .E(n1178), .CK(clk), .QN(n702) );
  EDFFX1 R11_reg_18_ ( .D(data_in_3[86]), .E(n1178), .CK(clk), .QN(n703) );
  EDFFX1 R11_reg_17_ ( .D(data_in_3[85]), .E(n1177), .CK(clk), .QN(n704) );
  EDFFXL R11_reg_16_ ( .D(data_in_3[84]), .E(n1177), .CK(clk), .QN(n705) );
  EDFFXL R11_reg_15_ ( .D(data_in_3[83]), .E(n1177), .CK(clk), .QN(n706) );
  EDFFXL R11_reg_14_ ( .D(data_in_3[82]), .E(n1177), .CK(clk), .QN(n707) );
  EDFFXL R11_reg_13_ ( .D(data_in_3[81]), .E(n1177), .CK(clk), .QN(n708) );
  EDFFXL R11_reg_12_ ( .D(data_in_3[80]), .E(n1177), .CK(clk), .QN(n709) );
  EDFFX1 R11_reg_11_ ( .D(data_in_3[79]), .E(n1177), .CK(clk), .QN(n710) );
  EDFFX1 R11_reg_10_ ( .D(data_in_3[78]), .E(n1177), .CK(clk), .QN(n711) );
  EDFFX1 R11_reg_9_ ( .D(data_in_3[77]), .E(n1177), .CK(clk), .QN(n712) );
  EDFFX1 R11_reg_8_ ( .D(data_in_3[76]), .E(n1177), .CK(clk), .QN(n713) );
  EDFFX1 R11_reg_7_ ( .D(data_in_3[75]), .E(n1177), .CK(clk), .QN(n714) );
  EDFFX1 R11_reg_6_ ( .D(data_in_3[74]), .E(n1177), .CK(clk), .QN(n715) );
  EDFFX1 R11_reg_5_ ( .D(data_in_3[73]), .E(n1177), .CK(clk), .QN(n716) );
  EDFFX1 R11_reg_4_ ( .D(data_in_3[72]), .E(n1176), .CK(clk), .QN(n717) );
  EDFFX1 R11_reg_3_ ( .D(data_in_3[71]), .E(n1176), .CK(clk), .QN(n718) );
  EDFFX1 R11_reg_2_ ( .D(data_in_3[70]), .E(n1176), .CK(clk), .QN(n719) );
  EDFFX1 R11_reg_1_ ( .D(data_in_3[69]), .E(n1176), .CK(clk), .QN(n720) );
  EDFFX1 R11_reg_0_ ( .D(data_in_3[68]), .E(n1176), .CK(clk), .QN(n721) );
  EDFFXL R8_reg_33_ ( .D(data_in_3[101]), .E(n891), .CK(clk), .QN(n756) );
  EDFFXL R8_reg_32_ ( .D(data_in_3[100]), .E(n891), .CK(clk), .QN(n757) );
  EDFFXL R8_reg_31_ ( .D(data_in_3[99]), .E(n891), .CK(clk), .QN(n758) );
  EDFFXL R8_reg_30_ ( .D(data_in_3[98]), .E(n891), .CK(clk), .QN(n759) );
  EDFFXL R8_reg_29_ ( .D(data_in_3[97]), .E(n891), .CK(clk), .QN(n760) );
  EDFFXL R8_reg_28_ ( .D(data_in_3[96]), .E(n891), .CK(clk), .QN(n761) );
  EDFFXL R8_reg_27_ ( .D(data_in_3[95]), .E(n891), .CK(clk), .QN(n762) );
  EDFFX1 R8_reg_26_ ( .D(data_in_3[94]), .E(n891), .CK(clk), .QN(n763) );
  EDFFX1 R8_reg_25_ ( .D(data_in_3[93]), .E(n891), .CK(clk), .QN(n764) );
  EDFFX1 R8_reg_24_ ( .D(data_in_3[92]), .E(n891), .CK(clk), .QN(n765) );
  EDFFX1 R8_reg_23_ ( .D(data_in_3[91]), .E(n126), .CK(clk), .QN(n766) );
  EDFFX1 R8_reg_22_ ( .D(data_in_3[90]), .E(n126), .CK(clk), .QN(n767) );
  EDFFX1 R8_reg_21_ ( .D(data_in_3[89]), .E(n126), .CK(clk), .QN(n768) );
  EDFFX1 R8_reg_20_ ( .D(data_in_3[88]), .E(n126), .CK(clk), .QN(n769) );
  EDFFX1 R8_reg_19_ ( .D(data_in_3[87]), .E(n126), .CK(clk), .QN(n770) );
  EDFFX1 R8_reg_18_ ( .D(data_in_3[86]), .E(n889), .CK(clk), .QN(n771) );
  EDFFX1 R8_reg_17_ ( .D(data_in_3[85]), .E(n894), .CK(clk), .QN(n772) );
  EDFFXL R8_reg_16_ ( .D(data_in_3[84]), .E(n126), .CK(clk), .QN(n773) );
  EDFFXL R8_reg_15_ ( .D(data_in_3[83]), .E(n126), .CK(clk), .QN(n774) );
  EDFFXL R8_reg_14_ ( .D(data_in_3[82]), .E(n126), .CK(clk), .QN(n775) );
  EDFFXL R8_reg_13_ ( .D(data_in_3[81]), .E(n126), .CK(clk), .QN(n776) );
  EDFFXL R8_reg_12_ ( .D(data_in_3[80]), .E(n126), .CK(clk), .QN(n777) );
  EDFFX1 R8_reg_11_ ( .D(data_in_3[79]), .E(n126), .CK(clk), .QN(n778) );
  EDFFX1 R8_reg_10_ ( .D(data_in_3[78]), .E(n892), .CK(clk), .QN(n779) );
  EDFFX1 R8_reg_9_ ( .D(data_in_3[77]), .E(n892), .CK(clk), .QN(n780) );
  EDFFX1 R8_reg_8_ ( .D(data_in_3[76]), .E(n892), .CK(clk), .QN(n781) );
  EDFFX1 R8_reg_7_ ( .D(data_in_3[75]), .E(n892), .CK(clk), .QN(n782) );
  EDFFX1 R8_reg_6_ ( .D(data_in_3[74]), .E(n892), .CK(clk), .QN(n783) );
  EDFFX1 R8_reg_5_ ( .D(data_in_3[73]), .E(n892), .CK(clk), .QN(n784) );
  EDFFX1 R8_reg_4_ ( .D(data_in_3[72]), .E(n892), .CK(clk), .QN(n785) );
  EDFFX1 R8_reg_3_ ( .D(data_in_3[71]), .E(n892), .CK(clk), .QN(n786) );
  EDFFX1 R8_reg_2_ ( .D(data_in_3[70]), .E(n892), .CK(clk), .QN(n787) );
  EDFFX1 R8_reg_1_ ( .D(data_in_3[69]), .E(n892), .CK(clk), .QN(n788) );
  EDFFX1 R8_reg_0_ ( .D(data_in_3[68]), .E(n892), .CK(clk), .QN(n789) );
  EDFFXL R9_reg_33_ ( .D(data_in_3[101]), .E(n1170), .CK(clk), .QN(n824) );
  EDFFXL R9_reg_32_ ( .D(data_in_3[100]), .E(n1170), .CK(clk), .QN(n825) );
  EDFFXL R9_reg_31_ ( .D(data_in_3[99]), .E(n1170), .CK(clk), .QN(n826) );
  EDFFXL R9_reg_30_ ( .D(data_in_3[98]), .E(n1170), .CK(clk), .QN(n827) );
  EDFFXL R9_reg_29_ ( .D(data_in_3[97]), .E(n1170), .CK(clk), .QN(n828) );
  EDFFXL R9_reg_28_ ( .D(data_in_3[96]), .E(n1170), .CK(clk), .QN(n829) );
  EDFFXL R9_reg_27_ ( .D(data_in_3[95]), .E(n1170), .CK(clk), .QN(n830) );
  EDFFX1 R9_reg_26_ ( .D(data_in_3[94]), .E(n1170), .CK(clk), .QN(n831) );
  EDFFX1 R9_reg_25_ ( .D(data_in_3[93]), .E(n1170), .CK(clk), .QN(n832) );
  EDFFX1 R9_reg_24_ ( .D(data_in_3[92]), .E(n1170), .CK(clk), .QN(n833) );
  EDFFX1 R9_reg_23_ ( .D(data_in_3[91]), .E(n125), .CK(clk), .QN(n834) );
  EDFFX1 R9_reg_22_ ( .D(data_in_3[90]), .E(n125), .CK(clk), .QN(n835) );
  EDFFX1 R9_reg_21_ ( .D(data_in_3[89]), .E(n125), .CK(clk), .QN(n836) );
  EDFFX1 R9_reg_20_ ( .D(data_in_3[88]), .E(n125), .CK(clk), .QN(n837) );
  EDFFX1 R9_reg_19_ ( .D(data_in_3[87]), .E(n1167), .CK(clk), .QN(n838) );
  EDFFX1 R9_reg_18_ ( .D(data_in_3[86]), .E(n1166), .CK(clk), .QN(n839) );
  EDFFX1 R9_reg_17_ ( .D(data_in_3[85]), .E(n1168), .CK(clk), .QN(n840) );
  EDFFXL R9_reg_16_ ( .D(data_in_3[84]), .E(n125), .CK(clk), .QN(n841) );
  EDFFXL R9_reg_15_ ( .D(data_in_3[83]), .E(n125), .CK(clk), .QN(n842) );
  EDFFXL R9_reg_14_ ( .D(data_in_3[82]), .E(n125), .CK(clk), .QN(n843) );
  EDFFXL R9_reg_13_ ( .D(data_in_3[81]), .E(n125), .CK(clk), .QN(n844) );
  EDFFXL R9_reg_12_ ( .D(data_in_3[80]), .E(n125), .CK(clk), .QN(n845) );
  EDFFX1 R9_reg_11_ ( .D(data_in_3[79]), .E(n1170), .CK(clk), .QN(n846) );
  EDFFX1 R9_reg_10_ ( .D(data_in_3[78]), .E(n125), .CK(clk), .QN(n847) );
  EDFFX1 R9_reg_9_ ( .D(data_in_3[77]), .E(n125), .CK(clk), .QN(n848) );
  EDFFX1 R9_reg_8_ ( .D(data_in_3[76]), .E(n125), .CK(clk), .QN(n849) );
  EDFFX1 R9_reg_7_ ( .D(data_in_3[75]), .E(n125), .CK(clk), .QN(n850) );
  EDFFX1 R9_reg_6_ ( .D(data_in_3[74]), .E(n125), .CK(clk), .QN(n851) );
  EDFFX1 R9_reg_5_ ( .D(data_in_3[73]), .E(n1169), .CK(clk), .QN(n852) );
  EDFFX1 R9_reg_4_ ( .D(data_in_3[72]), .E(n1171), .CK(clk), .QN(n853) );
  EDFFX1 R9_reg_3_ ( .D(data_in_3[71]), .E(n1167), .CK(clk), .QN(n854) );
  EDFFX1 R9_reg_2_ ( .D(data_in_3[70]), .E(n1168), .CK(clk), .QN(n855) );
  EDFFX1 R9_reg_1_ ( .D(data_in_3[69]), .E(n1172), .CK(clk), .QN(n856) );
  EDFFX1 R9_reg_0_ ( .D(data_in_3[68]), .E(n1169), .CK(clk), .QN(n857) );
  EDFFXL R14_reg_32_ ( .D(data_in_3[134]), .E(n1187), .CK(clk), .Q(R14[32]) );
  EDFFXL R14_reg_31_ ( .D(data_in_3[133]), .E(n1187), .CK(clk), .Q(R14[31]) );
  EDFFXL R14_reg_30_ ( .D(data_in_3[132]), .E(n1187), .CK(clk), .Q(R14[30]) );
  EDFFXL R14_reg_29_ ( .D(data_in_3[131]), .E(n1187), .CK(clk), .Q(R14[29]) );
  EDFFX1 R14_reg_28_ ( .D(data_in_3[130]), .E(n1187), .CK(clk), .Q(R14[28]) );
  EDFFX1 R14_reg_27_ ( .D(data_in_3[129]), .E(n1187), .CK(clk), .Q(R14[27]) );
  EDFFX1 R14_reg_26_ ( .D(data_in_3[128]), .E(n1187), .CK(clk), .Q(R14[26]) );
  EDFFX1 R14_reg_25_ ( .D(data_in_3[127]), .E(n1187), .CK(clk), .Q(R14[25]) );
  EDFFX1 R14_reg_24_ ( .D(data_in_3[126]), .E(n1187), .CK(clk), .Q(R14[24]) );
  EDFFX1 R14_reg_23_ ( .D(data_in_3[125]), .E(n1187), .CK(clk), .Q(R14[23]) );
  EDFFX1 R14_reg_22_ ( .D(data_in_3[124]), .E(n1186), .CK(clk), .Q(R14[22]) );
  EDFFX1 R14_reg_21_ ( .D(data_in_3[123]), .E(n1186), .CK(clk), .Q(R14[21]) );
  EDFFX1 R14_reg_20_ ( .D(data_in_3[122]), .E(n1186), .CK(clk), .Q(R14[20]) );
  EDFFX1 R14_reg_19_ ( .D(data_in_3[121]), .E(n1186), .CK(clk), .Q(R14[19]) );
  EDFFX1 R14_reg_18_ ( .D(data_in_3[120]), .E(n1186), .CK(clk), .Q(R14[18]) );
  EDFFX1 R14_reg_17_ ( .D(data_in_3[119]), .E(n1186), .CK(clk), .Q(R14[17]) );
  EDFFXL R14_reg_16_ ( .D(data_in_3[118]), .E(n1186), .CK(clk), .Q(R14[16]) );
  EDFFXL R14_reg_15_ ( .D(data_in_3[117]), .E(n1186), .CK(clk), .Q(R14[15]) );
  EDFFXL R14_reg_14_ ( .D(data_in_3[116]), .E(n1186), .CK(clk), .Q(R14[14]) );
  EDFFXL R14_reg_13_ ( .D(data_in_3[115]), .E(n1186), .CK(clk), .Q(R14[13]) );
  EDFFXL R14_reg_12_ ( .D(data_in_3[114]), .E(n1186), .CK(clk), .Q(R14[12]) );
  EDFFX1 R14_reg_11_ ( .D(data_in_3[113]), .E(n1186), .CK(clk), .Q(R14[11]) );
  EDFFX1 R14_reg_10_ ( .D(data_in_3[112]), .E(n1186), .CK(clk), .Q(R14[10]) );
  EDFFX1 R14_reg_9_ ( .D(data_in_3[111]), .E(n1186), .CK(clk), .Q(R14[9]) );
  EDFFX1 R14_reg_8_ ( .D(data_in_3[110]), .E(n1187), .CK(clk), .Q(R14[8]) );
  EDFFX1 R14_reg_7_ ( .D(data_in_3[109]), .E(n1185), .CK(clk), .Q(R14[7]) );
  EDFFX1 R14_reg_6_ ( .D(data_in_3[108]), .E(n1188), .CK(clk), .Q(R14[6]) );
  EDFFX1 R14_reg_5_ ( .D(data_in_3[107]), .E(n1188), .CK(clk), .Q(R14[5]) );
  EDFFX1 R14_reg_4_ ( .D(data_in_3[106]), .E(n1189), .CK(clk), .Q(R14[4]) );
  EDFFX1 R14_reg_3_ ( .D(data_in_3[105]), .E(n1183), .CK(clk), .Q(R14[3]) );
  EDFFX1 R14_reg_2_ ( .D(data_in_3[104]), .E(n1184), .CK(clk), .Q(R14[2]) );
  EDFFX1 R14_reg_1_ ( .D(data_in_3[103]), .E(n1186), .CK(clk), .Q(R14[1]) );
  EDFFX1 R14_reg_0_ ( .D(data_in_3[102]), .E(n1187), .CK(clk), .Q(R14[0]) );
  EDFFXL R15_reg_32_ ( .D(data_in_3[134]), .E(n1176), .CK(clk), .Q(R15[32]) );
  EDFFXL R15_reg_31_ ( .D(data_in_3[133]), .E(n1176), .CK(clk), .Q(R15[31]) );
  EDFFXL R15_reg_30_ ( .D(data_in_3[132]), .E(n1176), .CK(clk), .Q(R15[30]) );
  EDFFXL R15_reg_29_ ( .D(data_in_3[131]), .E(n1176), .CK(clk), .Q(R15[29]) );
  EDFFX1 R15_reg_28_ ( .D(data_in_3[130]), .E(n1176), .CK(clk), .Q(R15[28]) );
  EDFFX1 R15_reg_27_ ( .D(data_in_3[129]), .E(n1176), .CK(clk), .Q(R15[27]) );
  EDFFX1 R15_reg_26_ ( .D(data_in_3[128]), .E(n1176), .CK(clk), .Q(R15[26]) );
  EDFFX1 R15_reg_25_ ( .D(data_in_3[127]), .E(n1175), .CK(clk), .Q(R15[25]) );
  EDFFX1 R15_reg_24_ ( .D(data_in_3[126]), .E(n1175), .CK(clk), .Q(R15[24]) );
  EDFFX1 R15_reg_23_ ( .D(data_in_3[125]), .E(n1175), .CK(clk), .Q(R15[23]) );
  EDFFX1 R15_reg_22_ ( .D(data_in_3[124]), .E(n1175), .CK(clk), .Q(R15[22]) );
  EDFFX1 R15_reg_21_ ( .D(data_in_3[123]), .E(n1175), .CK(clk), .Q(R15[21]) );
  EDFFX1 R15_reg_20_ ( .D(data_in_3[122]), .E(n1175), .CK(clk), .Q(R15[20]) );
  EDFFX1 R15_reg_19_ ( .D(data_in_3[121]), .E(n1175), .CK(clk), .Q(R15[19]) );
  EDFFX1 R15_reg_18_ ( .D(data_in_3[120]), .E(n1175), .CK(clk), .Q(R15[18]) );
  EDFFX1 R15_reg_17_ ( .D(data_in_3[119]), .E(n1175), .CK(clk), .Q(R15[17]) );
  EDFFXL R15_reg_16_ ( .D(data_in_3[118]), .E(n1175), .CK(clk), .Q(R15[16]) );
  EDFFXL R15_reg_15_ ( .D(data_in_3[117]), .E(n1175), .CK(clk), .Q(R15[15]) );
  EDFFXL R15_reg_14_ ( .D(data_in_3[116]), .E(n1175), .CK(clk), .Q(R15[14]) );
  EDFFXL R15_reg_13_ ( .D(data_in_3[115]), .E(n1175), .CK(clk), .Q(R15[13]) );
  EDFFXL R15_reg_12_ ( .D(data_in_3[114]), .E(n1176), .CK(clk), .Q(R15[12]) );
  EDFFX1 R15_reg_11_ ( .D(data_in_3[113]), .E(n1177), .CK(clk), .Q(R15[11]) );
  EDFFX1 R15_reg_10_ ( .D(data_in_3[112]), .E(n1175), .CK(clk), .Q(R15[10]) );
  EDFFX1 R15_reg_9_ ( .D(data_in_3[111]), .E(n1178), .CK(clk), .Q(R15[9]) );
  EDFFX1 R15_reg_8_ ( .D(data_in_3[110]), .E(n1179), .CK(clk), .Q(R15[8]) );
  EDFFX1 R15_reg_7_ ( .D(data_in_3[109]), .E(n1181), .CK(clk), .Q(R15[7]) );
  EDFFX1 R15_reg_6_ ( .D(data_in_3[108]), .E(n1181), .CK(clk), .Q(R15[6]) );
  EDFFX1 R15_reg_5_ ( .D(data_in_3[107]), .E(n1180), .CK(clk), .Q(R15[5]) );
  EDFFX1 R15_reg_4_ ( .D(data_in_3[106]), .E(n1176), .CK(clk), .Q(R15[4]) );
  EDFFX1 R15_reg_3_ ( .D(data_in_3[105]), .E(n1177), .CK(clk), .Q(R15[3]) );
  EDFFX1 R15_reg_2_ ( .D(data_in_3[104]), .E(n1175), .CK(clk), .Q(R15[2]) );
  EDFFX1 R15_reg_1_ ( .D(data_in_3[103]), .E(n1178), .CK(clk), .Q(R15[1]) );
  EDFFX1 R15_reg_0_ ( .D(data_in_3[102]), .E(n1179), .CK(clk), .Q(R15[0]) );
  EDFFXL R12_reg_32_ ( .D(data_in_3[134]), .E(n892), .CK(clk), .Q(R12[32]) );
  EDFFXL R12_reg_31_ ( .D(data_in_3[133]), .E(n893), .CK(clk), .Q(R12[31]) );
  EDFFXL R12_reg_30_ ( .D(data_in_3[132]), .E(n893), .CK(clk), .Q(R12[30]) );
  EDFFXL R12_reg_29_ ( .D(data_in_3[131]), .E(n893), .CK(clk), .Q(R12[29]) );
  EDFFX1 R12_reg_28_ ( .D(data_in_3[130]), .E(n893), .CK(clk), .Q(R12[28]) );
  EDFFX1 R12_reg_27_ ( .D(data_in_3[129]), .E(n893), .CK(clk), .Q(R12[27]) );
  EDFFX1 R12_reg_26_ ( .D(data_in_3[128]), .E(n893), .CK(clk), .Q(R12[26]) );
  EDFFX1 R12_reg_25_ ( .D(data_in_3[127]), .E(n893), .CK(clk), .Q(R12[25]) );
  EDFFX1 R12_reg_24_ ( .D(data_in_3[126]), .E(n893), .CK(clk), .Q(R12[24]) );
  EDFFX1 R12_reg_23_ ( .D(data_in_3[125]), .E(n893), .CK(clk), .Q(R12[23]) );
  EDFFX1 R12_reg_22_ ( .D(data_in_3[124]), .E(n893), .CK(clk), .Q(R12[22]) );
  EDFFX1 R12_reg_21_ ( .D(data_in_3[123]), .E(n893), .CK(clk), .Q(R12[21]) );
  EDFFX1 R12_reg_20_ ( .D(data_in_3[122]), .E(n893), .CK(clk), .Q(R12[20]) );
  EDFFX1 R12_reg_19_ ( .D(data_in_3[121]), .E(n893), .CK(clk), .Q(R12[19]) );
  EDFFX1 R12_reg_18_ ( .D(data_in_3[120]), .E(n894), .CK(clk), .Q(R12[18]) );
  EDFFX1 R12_reg_17_ ( .D(data_in_3[119]), .E(n894), .CK(clk), .Q(R12[17]) );
  EDFFXL R12_reg_16_ ( .D(data_in_3[118]), .E(n894), .CK(clk), .Q(R12[16]) );
  EDFFXL R12_reg_15_ ( .D(data_in_3[117]), .E(n894), .CK(clk), .Q(R12[15]) );
  EDFFXL R12_reg_14_ ( .D(data_in_3[116]), .E(n894), .CK(clk), .Q(R12[14]) );
  EDFFXL R12_reg_13_ ( .D(data_in_3[115]), .E(n894), .CK(clk), .Q(R12[13]) );
  EDFFXL R12_reg_12_ ( .D(data_in_3[114]), .E(n894), .CK(clk), .Q(R12[12]) );
  EDFFX1 R12_reg_11_ ( .D(data_in_3[113]), .E(n894), .CK(clk), .Q(R12[11]) );
  EDFFX1 R12_reg_10_ ( .D(data_in_3[112]), .E(n894), .CK(clk), .Q(R12[10]) );
  EDFFX1 R12_reg_9_ ( .D(data_in_3[111]), .E(n894), .CK(clk), .Q(R12[9]) );
  EDFFX1 R12_reg_8_ ( .D(data_in_3[110]), .E(n894), .CK(clk), .Q(R12[8]) );
  EDFFX1 R12_reg_7_ ( .D(data_in_3[109]), .E(n894), .CK(clk), .Q(R12[7]) );
  EDFFX1 R12_reg_6_ ( .D(data_in_3[108]), .E(n894), .CK(clk), .Q(R12[6]) );
  EDFFX1 R12_reg_5_ ( .D(data_in_3[107]), .E(n888), .CK(clk), .Q(R12[5]) );
  EDFFX1 R12_reg_4_ ( .D(data_in_3[106]), .E(n887), .CK(clk), .Q(R12[4]) );
  EDFFX1 R12_reg_3_ ( .D(data_in_3[105]), .E(n887), .CK(clk), .Q(R12[3]) );
  EDFFX1 R12_reg_2_ ( .D(data_in_3[104]), .E(n888), .CK(clk), .Q(R12[2]) );
  EDFFX1 R12_reg_1_ ( .D(data_in_3[103]), .E(n887), .CK(clk), .Q(R12[1]) );
  EDFFX1 R12_reg_0_ ( .D(data_in_3[102]), .E(n887), .CK(clk), .Q(R12[0]) );
  EDFFXL R13_reg_32_ ( .D(data_in_3[134]), .E(n125), .CK(clk), .Q(R13[32]) );
  EDFFXL R13_reg_31_ ( .D(data_in_3[133]), .E(n1171), .CK(clk), .Q(R13[31]) );
  EDFFXL R13_reg_30_ ( .D(data_in_3[132]), .E(n1171), .CK(clk), .Q(R13[30]) );
  EDFFXL R13_reg_29_ ( .D(data_in_3[131]), .E(n1171), .CK(clk), .Q(R13[29]) );
  EDFFX1 R13_reg_28_ ( .D(data_in_3[130]), .E(n1171), .CK(clk), .Q(R13[28]) );
  EDFFX1 R13_reg_27_ ( .D(data_in_3[129]), .E(n1171), .CK(clk), .Q(R13[27]) );
  EDFFX1 R13_reg_26_ ( .D(data_in_3[128]), .E(n1171), .CK(clk), .Q(R13[26]) );
  EDFFX1 R13_reg_25_ ( .D(data_in_3[127]), .E(n1171), .CK(clk), .Q(R13[25]) );
  EDFFX1 R13_reg_24_ ( .D(data_in_3[126]), .E(n1171), .CK(clk), .Q(R13[24]) );
  EDFFX1 R13_reg_23_ ( .D(data_in_3[125]), .E(n1171), .CK(clk), .Q(R13[23]) );
  EDFFX1 R13_reg_22_ ( .D(data_in_3[124]), .E(n1171), .CK(clk), .Q(R13[22]) );
  EDFFX1 R13_reg_21_ ( .D(data_in_3[123]), .E(n1171), .CK(clk), .Q(R13[21]) );
  EDFFX1 R13_reg_20_ ( .D(data_in_3[122]), .E(n1171), .CK(clk), .Q(R13[20]) );
  EDFFX1 R13_reg_19_ ( .D(data_in_3[121]), .E(n1171), .CK(clk), .Q(R13[19]) );
  EDFFX1 R13_reg_18_ ( .D(data_in_3[120]), .E(n1172), .CK(clk), .Q(R13[18]) );
  EDFFX1 R13_reg_17_ ( .D(data_in_3[119]), .E(n1172), .CK(clk), .Q(R13[17]) );
  EDFFXL R13_reg_15_ ( .D(data_in_3[117]), .E(n1172), .CK(clk), .Q(R13[15]) );
  EDFFXL R13_reg_14_ ( .D(data_in_3[116]), .E(n1172), .CK(clk), .Q(R13[14]) );
  EDFFXL R13_reg_13_ ( .D(data_in_3[115]), .E(n1172), .CK(clk), .Q(R13[13]) );
  EDFFXL R13_reg_12_ ( .D(data_in_3[114]), .E(n1172), .CK(clk), .Q(R13[12]) );
  EDFFX1 R13_reg_11_ ( .D(data_in_3[113]), .E(n1172), .CK(clk), .Q(R13[11]) );
  EDFFX1 R13_reg_10_ ( .D(data_in_3[112]), .E(n1172), .CK(clk), .Q(R13[10]) );
  EDFFX1 R13_reg_9_ ( .D(data_in_3[111]), .E(n1172), .CK(clk), .Q(R13[9]) );
  EDFFX1 R13_reg_8_ ( .D(data_in_3[110]), .E(n1172), .CK(clk), .Q(R13[8]) );
  EDFFX1 R13_reg_7_ ( .D(data_in_3[109]), .E(n1172), .CK(clk), .Q(R13[7]) );
  EDFFX1 R13_reg_6_ ( .D(data_in_3[108]), .E(n1172), .CK(clk), .Q(R13[6]) );
  EDFFX1 R13_reg_5_ ( .D(data_in_3[107]), .E(n1171), .CK(clk), .Q(R13[5]) );
  EDFFX1 R13_reg_4_ ( .D(data_in_3[106]), .E(n1166), .CK(clk), .Q(R13[4]) );
  EDFFX1 R13_reg_3_ ( .D(data_in_3[105]), .E(n1166), .CK(clk), .Q(R13[3]) );
  EDFFX1 R13_reg_2_ ( .D(data_in_3[104]), .E(n1166), .CK(clk), .Q(R13[2]) );
  EDFFX1 R13_reg_1_ ( .D(data_in_3[103]), .E(n1166), .CK(clk), .Q(R13[1]) );
  EDFFX1 R13_reg_0_ ( .D(data_in_3[102]), .E(n1166), .CK(clk), .Q(R13[0]) );
  EDFFXL R2_reg_31_ ( .D(data_in_3[31]), .E(n1189), .CK(clk), .Q(R2[31]) );
  EDFFXL R2_reg_30_ ( .D(data_in_3[30]), .E(n1188), .CK(clk), .Q(R2[30]) );
  EDFFXL R2_reg_29_ ( .D(data_in_3[29]), .E(n1189), .CK(clk), .Q(R2[29]) );
  EDFFX1 R2_reg_22_ ( .D(data_in_3[22]), .E(n1189), .CK(clk), .Q(R2[22]) );
  EDFFX1 R2_reg_21_ ( .D(data_in_3[21]), .E(n1189), .CK(clk), .Q(R2[21]) );
  EDFFX1 R2_reg_20_ ( .D(data_in_3[20]), .E(n1189), .CK(clk), .Q(R2[20]) );
  EDFFX1 R2_reg_19_ ( .D(data_in_3[19]), .E(n1189), .CK(clk), .Q(R2[19]) );
  EDFFX1 R2_reg_18_ ( .D(data_in_3[18]), .E(n1189), .CK(clk), .Q(R2[18]) );
  EDFFX1 R2_reg_17_ ( .D(data_in_3[17]), .E(n1189), .CK(clk), .Q(R2[17]) );
  EDFFXL R2_reg_16_ ( .D(data_in_3[16]), .E(n1189), .CK(clk), .Q(R2[16]) );
  EDFFXL R2_reg_15_ ( .D(data_in_3[15]), .E(n1189), .CK(clk), .Q(R2[15]) );
  EDFFXL R2_reg_13_ ( .D(data_in_3[13]), .E(n1188), .CK(clk), .Q(R2[13]) );
  EDFFXL R2_reg_12_ ( .D(data_in_3[12]), .E(n1188), .CK(clk), .Q(R2[12]) );
  EDFFX1 R2_reg_5_ ( .D(data_in_3[5]), .E(n1188), .CK(clk), .Q(R2[5]) );
  EDFFX1 R2_reg_4_ ( .D(data_in_3[4]), .E(n1188), .CK(clk), .Q(R2[4]) );
  EDFFX1 R2_reg_3_ ( .D(data_in_3[3]), .E(n1188), .CK(clk), .Q(R2[3]) );
  EDFFX1 R2_reg_2_ ( .D(data_in_3[2]), .E(n1188), .CK(clk), .Q(R2[2]) );
  EDFFX1 R2_reg_1_ ( .D(data_in_3[1]), .E(n1187), .CK(clk), .Q(R2[1]) );
  EDFFX1 R2_reg_0_ ( .D(data_in_3[0]), .E(n1187), .CK(clk), .Q(R2[0]) );
  EDFFXL R3_reg_31_ ( .D(data_in_3[31]), .E(n1181), .CK(clk), .Q(R3[31]) );
  EDFFXL R3_reg_30_ ( .D(data_in_3[30]), .E(n1176), .CK(clk), .Q(R3[30]) );
  EDFFXL R3_reg_29_ ( .D(data_in_3[29]), .E(n1177), .CK(clk), .Q(R3[29]) );
  EDFFX1 R3_reg_22_ ( .D(data_in_3[22]), .E(n1180), .CK(clk), .Q(R3[22]) );
  EDFFX1 R3_reg_21_ ( .D(data_in_3[21]), .E(n1180), .CK(clk), .Q(R3[21]) );
  EDFFX1 R3_reg_20_ ( .D(data_in_3[20]), .E(n1180), .CK(clk), .Q(R3[20]) );
  EDFFX1 R3_reg_19_ ( .D(data_in_3[19]), .E(n1180), .CK(clk), .Q(R3[19]) );
  EDFFX1 R3_reg_18_ ( .D(data_in_3[18]), .E(n1180), .CK(clk), .Q(R3[18]) );
  EDFFX1 R3_reg_17_ ( .D(data_in_3[17]), .E(n1180), .CK(clk), .Q(R3[17]) );
  EDFFXL R3_reg_16_ ( .D(data_in_3[16]), .E(n1180), .CK(clk), .Q(R3[16]) );
  EDFFXL R3_reg_15_ ( .D(data_in_3[15]), .E(n1180), .CK(clk), .Q(R3[15]) );
  EDFFXL R3_reg_12_ ( .D(data_in_3[12]), .E(n1180), .CK(clk), .Q(R3[12]) );
  EDFFX1 R3_reg_5_ ( .D(data_in_3[5]), .E(n1179), .CK(clk), .Q(R3[5]) );
  EDFFX1 R3_reg_4_ ( .D(data_in_3[4]), .E(n1179), .CK(clk), .Q(R3[4]) );
  EDFFX1 R3_reg_3_ ( .D(data_in_3[3]), .E(n1179), .CK(clk), .Q(R3[3]) );
  EDFFX1 R3_reg_2_ ( .D(data_in_3[2]), .E(n1179), .CK(clk), .Q(R3[2]) );
  EDFFX1 R3_reg_1_ ( .D(data_in_3[1]), .E(n1179), .CK(clk), .Q(R3[1]) );
  EDFFX1 R3_reg_0_ ( .D(data_in_3[0]), .E(n1179), .CK(clk), .Q(R3[0]) );
  EDFFXL R0_reg_31_ ( .D(data_in_3[31]), .E(n887), .CK(clk), .Q(R0[31]) );
  EDFFXL R0_reg_30_ ( .D(data_in_3[30]), .E(n887), .CK(clk), .Q(R0[30]) );
  EDFFXL R0_reg_29_ ( .D(data_in_3[29]), .E(n887), .CK(clk), .Q(R0[29]) );
  EDFFX1 R0_reg_22_ ( .D(data_in_3[22]), .E(n887), .CK(clk), .Q(R0[22]) );
  EDFFX1 R0_reg_21_ ( .D(data_in_3[21]), .E(n887), .CK(clk), .Q(R0[21]) );
  EDFFX1 R0_reg_20_ ( .D(data_in_3[20]), .E(n888), .CK(clk), .Q(R0[20]) );
  EDFFX1 R0_reg_19_ ( .D(data_in_3[19]), .E(n888), .CK(clk), .Q(R0[19]) );
  EDFFX1 R0_reg_18_ ( .D(data_in_3[18]), .E(n888), .CK(clk), .Q(R0[18]) );
  EDFFX1 R0_reg_17_ ( .D(data_in_3[17]), .E(n888), .CK(clk), .Q(R0[17]) );
  EDFFXL R0_reg_16_ ( .D(data_in_3[16]), .E(n888), .CK(clk), .Q(R0[16]) );
  EDFFXL R0_reg_15_ ( .D(data_in_3[15]), .E(n888), .CK(clk), .Q(R0[15]) );
  EDFFXL R0_reg_13_ ( .D(data_in_3[13]), .E(n888), .CK(clk), .Q(R0[13]) );
  EDFFXL R0_reg_12_ ( .D(data_in_3[12]), .E(n888), .CK(clk), .Q(R0[12]) );
  EDFFX1 R0_reg_5_ ( .D(data_in_3[5]), .E(n126), .CK(clk), .Q(R0[5]) );
  EDFFX1 R0_reg_4_ ( .D(data_in_3[4]), .E(n126), .CK(clk), .Q(R0[4]) );
  EDFFX1 R0_reg_3_ ( .D(data_in_3[3]), .E(n126), .CK(clk), .Q(R0[3]) );
  EDFFX1 R0_reg_2_ ( .D(data_in_3[2]), .E(n126), .CK(clk), .Q(R0[2]) );
  EDFFX1 R0_reg_1_ ( .D(data_in_3[1]), .E(n893), .CK(clk), .Q(R0[1]) );
  EDFFX1 R0_reg_0_ ( .D(data_in_3[0]), .E(n892), .CK(clk), .Q(R0[0]) );
  EDFFXL R1_reg_31_ ( .D(data_in_3[31]), .E(n1166), .CK(clk), .Q(R1[31]) );
  EDFFXL R1_reg_30_ ( .D(data_in_3[30]), .E(n1166), .CK(clk), .Q(R1[30]) );
  EDFFXL R1_reg_29_ ( .D(data_in_3[29]), .E(n1166), .CK(clk), .Q(R1[29]) );
  EDFFX1 R1_reg_22_ ( .D(data_in_3[22]), .E(n1166), .CK(clk), .Q(R1[22]) );
  EDFFX1 R1_reg_21_ ( .D(data_in_3[21]), .E(n1166), .CK(clk), .Q(R1[21]) );
  EDFFX1 R1_reg_20_ ( .D(data_in_3[20]), .E(n1167), .CK(clk), .Q(R1[20]) );
  EDFFX1 R1_reg_19_ ( .D(data_in_3[19]), .E(n1167), .CK(clk), .Q(R1[19]) );
  EDFFX1 R1_reg_18_ ( .D(data_in_3[18]), .E(n1167), .CK(clk), .Q(R1[18]) );
  EDFFX1 R1_reg_17_ ( .D(data_in_3[17]), .E(n1167), .CK(clk), .Q(R1[17]) );
  EDFFXL R1_reg_16_ ( .D(data_in_3[16]), .E(n1167), .CK(clk), .Q(R1[16]) );
  EDFFXL R1_reg_15_ ( .D(data_in_3[15]), .E(n1167), .CK(clk), .Q(R1[15]) );
  EDFFXL R1_reg_13_ ( .D(data_in_3[13]), .E(n1167), .CK(clk), .Q(R1[13]) );
  EDFFXL R1_reg_12_ ( .D(data_in_3[12]), .E(n1167), .CK(clk), .Q(R1[12]) );
  EDFFX1 R1_reg_5_ ( .D(data_in_3[5]), .E(n1170), .CK(clk), .Q(R1[5]) );
  EDFFX1 R1_reg_4_ ( .D(data_in_3[4]), .E(n1167), .CK(clk), .Q(R1[4]) );
  EDFFX1 R1_reg_3_ ( .D(data_in_3[3]), .E(n1166), .CK(clk), .Q(R1[3]) );
  EDFFX1 R1_reg_2_ ( .D(data_in_3[2]), .E(n1168), .CK(clk), .Q(R1[2]) );
  EDFFX1 R1_reg_1_ ( .D(data_in_3[1]), .E(n1172), .CK(clk), .Q(R1[1]) );
  EDFFX1 R1_reg_0_ ( .D(data_in_3[0]), .E(n1167), .CK(clk), .Q(R1[0]) );
  JKFFRXL counter_1_reg_0_ ( .J(1'b1), .K(1'b1), .CK(clk), .RN(rst_n), .Q(
        counter_1[0]), .QN(n585) );
  JKFFRXL counter_2_reg_0_ ( .J(1'b1), .K(1'b1), .CK(clk), .RN(rst_n), .Q(
        counter_2[0]), .QN(n862) );
  DFFRHQX1 counter_2_reg_1_ ( .D(N50), .CK(clk), .RN(rst_n), .Q(counter_2[1])
         );
  DFFRHQX1 counter_2_reg_3_ ( .D(N52), .CK(clk), .RN(rst_n), .Q(counter_2[3])
         );
  DFFRHQX1 counter_2_reg_2_ ( .D(n1192), .CK(clk), .RN(rst_n), .Q(counter_2[2]) );
  DFFRHQX1 counter_1_reg_1_ ( .D(N26), .CK(clk), .RN(rst_n), .Q(counter_1[1])
         );
  EDFFX1 data_out_3_reg_33_ ( .D(N152), .E(n1191), .CK(clk), .Q(data_out_3[33]) );
  EDFFX1 data_out_3_reg_32_ ( .D(N151), .E(n1191), .CK(clk), .Q(data_out_3[32]) );
  EDFFX1 data_out_3_reg_31_ ( .D(N150), .E(n1191), .CK(clk), .Q(data_out_3[31]) );
  EDFFX1 data_out_3_reg_30_ ( .D(N149), .E(n1191), .CK(clk), .Q(data_out_3[30]) );
  EDFFX1 data_out_3_reg_29_ ( .D(N148), .E(n1191), .CK(clk), .Q(data_out_3[29]) );
  EDFFX1 data_out_3_reg_28_ ( .D(N147), .E(n1191), .CK(clk), .Q(data_out_3[28]) );
  EDFFX1 data_out_3_reg_27_ ( .D(N146), .E(n1191), .CK(clk), .Q(data_out_3[27]) );
  EDFFX1 data_out_3_reg_26_ ( .D(N145), .E(n1191), .CK(clk), .Q(data_out_3[26]) );
  EDFFX1 data_out_3_reg_25_ ( .D(N144), .E(n1191), .CK(clk), .Q(data_out_3[25]) );
  EDFFX1 data_out_3_reg_24_ ( .D(N143), .E(n1191), .CK(clk), .Q(data_out_3[24]) );
  EDFFX1 data_out_3_reg_23_ ( .D(N142), .E(n1191), .CK(clk), .Q(data_out_3[23]) );
  EDFFX1 data_out_3_reg_22_ ( .D(N141), .E(n1191), .CK(clk), .Q(data_out_3[22]) );
  EDFFX1 data_out_3_reg_21_ ( .D(N140), .E(n1191), .CK(clk), .Q(data_out_3[21]) );
  EDFFX1 data_out_3_reg_20_ ( .D(N139), .E(n1191), .CK(clk), .Q(data_out_3[20]) );
  EDFFX1 data_out_3_reg_19_ ( .D(N138), .E(n1191), .CK(clk), .Q(data_out_3[19]) );
  EDFFX1 data_out_3_reg_18_ ( .D(N137), .E(n1191), .CK(clk), .Q(data_out_3[18]) );
  EDFFX1 data_out_3_reg_17_ ( .D(N136), .E(n1191), .CK(clk), .Q(data_out_3[17]) );
  EDFFX1 data_out_3_reg_16_ ( .D(N135), .E(n1191), .CK(clk), .Q(data_out_3[16]) );
  EDFFX1 data_out_3_reg_15_ ( .D(N134), .E(n1191), .CK(clk), .Q(data_out_3[15]) );
  EDFFX1 data_out_3_reg_14_ ( .D(N133), .E(n1191), .CK(clk), .Q(data_out_3[14]) );
  EDFFX1 data_out_3_reg_13_ ( .D(N132), .E(n1191), .CK(clk), .Q(data_out_3[13]) );
  EDFFX1 data_out_3_reg_12_ ( .D(N131), .E(n1191), .CK(clk), .Q(data_out_3[12]) );
  EDFFX1 data_out_3_reg_11_ ( .D(N130), .E(n1191), .CK(clk), .Q(data_out_3[11]) );
  EDFFX1 data_out_3_reg_10_ ( .D(N129), .E(n1191), .CK(clk), .Q(data_out_3[10]) );
  EDFFX1 data_out_3_reg_9_ ( .D(N128), .E(n1191), .CK(clk), .Q(data_out_3[9])
         );
  EDFFX1 data_out_3_reg_8_ ( .D(N127), .E(n1191), .CK(clk), .Q(data_out_3[8])
         );
  EDFFX1 data_out_3_reg_7_ ( .D(N126), .E(n1191), .CK(clk), .Q(data_out_3[7])
         );
  EDFFX1 data_out_3_reg_6_ ( .D(N125), .E(n1191), .CK(clk), .Q(data_out_3[6])
         );
  EDFFX1 data_out_3_reg_5_ ( .D(N124), .E(n1191), .CK(clk), .Q(data_out_3[5])
         );
  EDFFX1 data_out_3_reg_4_ ( .D(N123), .E(n1191), .CK(clk), .Q(data_out_3[4])
         );
  EDFFX1 data_out_3_reg_3_ ( .D(N122), .E(n1191), .CK(clk), .Q(data_out_3[3])
         );
  EDFFX1 data_out_3_reg_2_ ( .D(N121), .E(n1191), .CK(clk), .Q(data_out_3[2])
         );
  EDFFX1 data_out_3_reg_1_ ( .D(N120), .E(n1191), .CK(clk), .Q(data_out_3[1])
         );
  EDFFX1 data_out_3_reg_0_ ( .D(N119), .E(n1191), .CK(clk), .Q(data_out_3[0])
         );
  EDFFXL R0_reg_28_ ( .D(data_in_3[28]), .E(n887), .CK(clk), .Q(R0[28]) );
  EDFFXL R0_reg_27_ ( .D(data_in_3[27]), .E(n887), .CK(clk), .Q(R0[27]) );
  EDFFXL R0_reg_26_ ( .D(data_in_3[26]), .E(n887), .CK(clk), .Q(R0[26]) );
  EDFFXL R0_reg_11_ ( .D(data_in_3[11]), .E(n888), .CK(clk), .Q(R0[11]) );
  EDFFXL R0_reg_10_ ( .D(data_in_3[10]), .E(n888), .CK(clk), .Q(R0[10]) );
  EDFFXL R2_reg_28_ ( .D(data_in_3[28]), .E(n1189), .CK(clk), .Q(R2[28]) );
  EDFFXL R2_reg_27_ ( .D(data_in_3[27]), .E(n1189), .CK(clk), .Q(R2[27]) );
  EDFFXL R2_reg_11_ ( .D(data_in_3[11]), .E(n1188), .CK(clk), .Q(R2[11]) );
  EDFFXL R2_reg_10_ ( .D(data_in_3[10]), .E(n1188), .CK(clk), .Q(R2[10]) );
  EDFFXL R3_reg_28_ ( .D(data_in_3[28]), .E(n1175), .CK(clk), .Q(R3[28]) );
  EDFFXL R3_reg_27_ ( .D(data_in_3[27]), .E(n1178), .CK(clk), .Q(R3[27]) );
  EDFFXL R3_reg_11_ ( .D(data_in_3[11]), .E(n1180), .CK(clk), .Q(R3[11]) );
  EDFFXL R3_reg_10_ ( .D(data_in_3[10]), .E(n1180), .CK(clk), .Q(R3[10]) );
  EDFFXL R1_reg_28_ ( .D(data_in_3[28]), .E(n1166), .CK(clk), .Q(R1[28]) );
  EDFFXL R1_reg_27_ ( .D(data_in_3[27]), .E(n1166), .CK(clk), .Q(R1[27]) );
  EDFFXL R1_reg_11_ ( .D(data_in_3[11]), .E(n1167), .CK(clk), .Q(R1[11]) );
  EDFFXL R1_reg_10_ ( .D(data_in_3[10]), .E(n1167), .CK(clk), .Q(R1[10]) );
  EDFFX1 R7_reg_28_ ( .D(data_in_3[62]), .E(n1179), .CK(clk), .QN(n591) );
  EDFFX1 R7_reg_27_ ( .D(data_in_3[61]), .E(n1176), .CK(clk), .QN(n592) );
  EDFFX1 R7_reg_26_ ( .D(data_in_3[60]), .E(n1180), .CK(clk), .QN(n593) );
  EDFFX1 R7_reg_25_ ( .D(data_in_3[59]), .E(n1181), .CK(clk), .QN(n594) );
  EDFFX1 R7_reg_24_ ( .D(data_in_3[58]), .E(n1177), .CK(clk), .QN(n595) );
  EDFFX1 R7_reg_23_ ( .D(data_in_3[57]), .E(n1175), .CK(clk), .QN(n596) );
  EDFFX1 R7_reg_11_ ( .D(data_in_3[45]), .E(n1181), .CK(clk), .QN(n608) );
  EDFFX1 R7_reg_10_ ( .D(data_in_3[44]), .E(n1181), .CK(clk), .QN(n609) );
  EDFFX1 R7_reg_9_ ( .D(data_in_3[43]), .E(n1181), .CK(clk), .QN(n610) );
  EDFFX1 R7_reg_8_ ( .D(data_in_3[42]), .E(n1181), .CK(clk), .QN(n611) );
  EDFFX1 R7_reg_7_ ( .D(data_in_3[41]), .E(n1181), .CK(clk), .QN(n612) );
  EDFFX1 R7_reg_6_ ( .D(data_in_3[40]), .E(n1181), .CK(clk), .QN(n613) );
  EDFFX1 R5_reg_16_ ( .D(data_in_3[50]), .E(n1168), .CK(clk), .QN(n807) );
  EDFFXL R7_reg_33_ ( .D(data_in_3[67]), .E(n1179), .CK(clk), .QN(n586) );
  EDFFXL R6_reg_33_ ( .D(data_in_3[67]), .E(n864), .CK(clk), .QN(n654) );
  EDFFXL R4_reg_33_ ( .D(data_in_3[67]), .E(n126), .CK(clk), .QN(n722) );
  JKFFRXL p_s_flag_out_reg ( .J(n1195), .K(1'b0), .CK(clk), .RN(rst_n), .Q(
        n1191) );
  EDFFXL R2_reg_32_ ( .D(data_in_3[32]), .E(n1188), .CK(clk), .Q(R2[32]) );
  EDFFXL R3_reg_32_ ( .D(data_in_3[32]), .E(n865), .CK(clk), .Q(R3[32]) );
  EDFFXL R1_reg_32_ ( .D(data_in_3[32]), .E(n125), .CK(clk), .Q(R1[32]) );
  EDFFXL R0_reg_32_ ( .D(data_in_3[32]), .E(n126), .CK(clk), .Q(R0[32]) );
  EDFFXL R3_reg_23_ ( .D(data_in_3[23]), .E(n865), .CK(clk), .Q(R3[23]) );
  EDFFXL R2_reg_23_ ( .D(data_in_3[23]), .E(n864), .CK(clk), .Q(R2[23]) );
  EDFFXL R1_reg_23_ ( .D(data_in_3[23]), .E(n125), .CK(clk), .Q(R1[23]) );
  EDFFXL R0_reg_23_ ( .D(data_in_3[23]), .E(n126), .CK(clk), .Q(R0[23]) );
  EDFFXL R3_reg_6_ ( .D(data_in_3[6]), .E(n865), .CK(clk), .Q(R3[6]) );
  EDFFXL R2_reg_6_ ( .D(data_in_3[6]), .E(n864), .CK(clk), .Q(R2[6]) );
  EDFFXL R1_reg_6_ ( .D(data_in_3[6]), .E(n125), .CK(clk), .Q(R1[6]) );
  EDFFXL R0_reg_6_ ( .D(data_in_3[6]), .E(n126), .CK(clk), .Q(R0[6]) );
  EDFFXL R3_reg_24_ ( .D(data_in_3[24]), .E(n865), .CK(clk), .Q(R3[24]) );
  EDFFXL R2_reg_24_ ( .D(data_in_3[24]), .E(n864), .CK(clk), .Q(R2[24]) );
  EDFFXL R1_reg_24_ ( .D(data_in_3[24]), .E(n125), .CK(clk), .Q(R1[24]) );
  EDFFXL R0_reg_24_ ( .D(data_in_3[24]), .E(n126), .CK(clk), .Q(R0[24]) );
  EDFFXL R3_reg_7_ ( .D(data_in_3[7]), .E(n865), .CK(clk), .Q(R3[7]) );
  EDFFXL R2_reg_7_ ( .D(data_in_3[7]), .E(n864), .CK(clk), .Q(R2[7]) );
  EDFFXL R1_reg_7_ ( .D(data_in_3[7]), .E(n125), .CK(clk), .Q(R1[7]) );
  EDFFXL R0_reg_7_ ( .D(data_in_3[7]), .E(n126), .CK(clk), .Q(R0[7]) );
  EDFFXL R3_reg_8_ ( .D(data_in_3[8]), .E(n865), .CK(clk), .Q(R3[8]) );
  EDFFXL R2_reg_8_ ( .D(data_in_3[8]), .E(n864), .CK(clk), .Q(R2[8]) );
  EDFFXL R1_reg_8_ ( .D(data_in_3[8]), .E(n125), .CK(clk), .Q(R1[8]) );
  EDFFXL R0_reg_8_ ( .D(data_in_3[8]), .E(n126), .CK(clk), .Q(R0[8]) );
  EDFFXL R3_reg_25_ ( .D(data_in_3[25]), .E(n865), .CK(clk), .Q(R3[25]) );
  EDFFXL R2_reg_25_ ( .D(data_in_3[25]), .E(n864), .CK(clk), .Q(R2[25]) );
  EDFFXL R1_reg_25_ ( .D(data_in_3[25]), .E(n125), .CK(clk), .Q(R1[25]) );
  EDFFXL R0_reg_25_ ( .D(data_in_3[25]), .E(n126), .CK(clk), .Q(R0[25]) );
  EDFFXL R3_reg_9_ ( .D(data_in_3[9]), .E(n865), .CK(clk), .Q(R3[9]) );
  EDFFXL R2_reg_9_ ( .D(data_in_3[9]), .E(n864), .CK(clk), .Q(R2[9]) );
  EDFFXL R1_reg_9_ ( .D(data_in_3[9]), .E(n125), .CK(clk), .Q(R1[9]) );
  EDFFXL R0_reg_9_ ( .D(data_in_3[9]), .E(n126), .CK(clk), .Q(R0[9]) );
  EDFFXL R3_reg_26_ ( .D(data_in_3[26]), .E(n865), .CK(clk), .Q(R3[26]) );
  EDFFXL R2_reg_26_ ( .D(data_in_3[26]), .E(n864), .CK(clk), .Q(R2[26]) );
  EDFFXL R1_reg_26_ ( .D(data_in_3[26]), .E(n125), .CK(clk), .Q(R1[26]) );
  EDFFX1 R13_reg_16_ ( .D(data_in_3[118]), .E(n1172), .CK(clk), .Q(R13[16]) );
  EDFFX1 R3_reg_13_ ( .D(data_in_3[13]), .E(n1180), .CK(clk), .Q(R3[13]) );
  EDFFXL R4_reg_32_ ( .D(data_in_3[66]), .E(n126), .CK(clk), .QN(n723) );
  EDFFXL R6_reg_32_ ( .D(data_in_3[66]), .E(n864), .CK(clk), .QN(n655) );
  EDFFXL R7_reg_32_ ( .D(data_in_3[66]), .E(n1180), .CK(clk), .QN(n587) );
  AND2X2 U3 ( .A(n1159), .B(n872), .Y(n6) );
  AND2X2 U6 ( .A(n1159), .B(n870), .Y(n7) );
  AND2X2 U7 ( .A(n1163), .B(n872), .Y(n8) );
  AND2X2 U8 ( .A(n1163), .B(n870), .Y(n9) );
  NAND2X1 U9 ( .A(n873), .B(n1159), .Y(n10) );
  NAND2X1 U10 ( .A(n1160), .B(n1159), .Y(n11) );
  NAND2X1 U11 ( .A(n1163), .B(n1160), .Y(n12) );
  NAND2X1 U12 ( .A(n1163), .B(n873), .Y(n13) );
  AND2X2 U13 ( .A(n872), .B(n1164), .Y(n14) );
  AND2X2 U14 ( .A(n1158), .B(n872), .Y(n15) );
  AND2X2 U15 ( .A(n1158), .B(n870), .Y(n16) );
  NAND2X1 U16 ( .A(n1160), .B(n1164), .Y(n17) );
  NAND2X1 U17 ( .A(n873), .B(n1164), .Y(n18) );
  NAND2X1 U18 ( .A(n873), .B(n1158), .Y(n19) );
  NAND2X1 U19 ( .A(n1160), .B(n1158), .Y(n20) );
  INVX1 U21 ( .A(n868), .Y(n1174) );
  INVX1 U22 ( .A(n1173), .Y(n1172) );
  INVX1 U23 ( .A(n1173), .Y(n1171) );
  INVX1 U24 ( .A(n1173), .Y(n1170) );
  INVX1 U25 ( .A(n1173), .Y(n1169) );
  INVX1 U26 ( .A(n1173), .Y(n1168) );
  INVX1 U27 ( .A(n896), .Y(n894) );
  INVX1 U28 ( .A(n896), .Y(n893) );
  INVX1 U29 ( .A(n896), .Y(n891) );
  INVX1 U30 ( .A(n896), .Y(n889) );
  INVX1 U31 ( .A(n1182), .Y(n1175) );
  INVX1 U32 ( .A(n1182), .Y(n1177) );
  INVX1 U33 ( .A(n1182), .Y(n1178) );
  INVX1 U34 ( .A(n1190), .Y(n1183) );
  INVX1 U35 ( .A(n1190), .Y(n1184) );
  INVX1 U36 ( .A(n1190), .Y(n1185) );
  INVX1 U37 ( .A(n1190), .Y(n1186) );
  INVX1 U38 ( .A(n1182), .Y(n1179) );
  INVX1 U39 ( .A(n1182), .Y(n1181) );
  INVX1 U40 ( .A(n1190), .Y(n1189) );
  INVX1 U41 ( .A(n1173), .Y(n1167) );
  INVX1 U42 ( .A(n896), .Y(n892) );
  INVX1 U43 ( .A(n896), .Y(n888) );
  INVX1 U44 ( .A(n1182), .Y(n1176) );
  INVX1 U45 ( .A(n1182), .Y(n1180) );
  INVX1 U46 ( .A(n1190), .Y(n1187) );
  INVX1 U47 ( .A(n1190), .Y(n1188) );
  INVX1 U48 ( .A(n1173), .Y(n1166) );
  INVX1 U49 ( .A(n896), .Y(n887) );
  NOR2X1 U50 ( .A(n1194), .B(n1193), .Y(n870) );
  NAND2X1 U51 ( .A(n1164), .B(n870), .Y(n868) );
  INVX1 U52 ( .A(n865), .Y(n1182) );
  INVX1 U53 ( .A(n125), .Y(n1173) );
  INVX1 U54 ( .A(n126), .Y(n896) );
  INVX1 U55 ( .A(n864), .Y(n1190) );
  NOR3X1 U56 ( .A(counter_1[1]), .B(p_s_flag_in), .C(n585), .Y(n865) );
  NOR3X1 U57 ( .A(counter_1[1]), .B(p_s_flag_in), .C(counter_1[0]), .Y(n864)
         );
  NOR2X1 U58 ( .A(n1194), .B(counter_2[1]), .Y(n873) );
  OAI221XL U59 ( .A0(n711), .A1(n17), .B0(n609), .B1(n12), .C0(n1079), .Y(
        n1074) );
  AOI22X1 U60 ( .A0(n14), .A1(R0[10]), .B0(n8), .B1(R15[10]), .Y(n1079) );
  OAI221XL U61 ( .A0(n710), .A1(n17), .B0(n608), .B1(n12), .C0(n1071), .Y(
        n1066) );
  AOI22X1 U62 ( .A0(n14), .A1(R0[11]), .B0(n8), .B1(R15[11]), .Y(n1071) );
  OAI221XL U63 ( .A0(n709), .A1(n17), .B0(n607), .B1(n12), .C0(n1063), .Y(
        n1058) );
  AOI22X1 U64 ( .A0(n14), .A1(R0[12]), .B0(n8), .B1(R15[12]), .Y(n1063) );
  OAI221XL U65 ( .A0(n708), .A1(n17), .B0(n606), .B1(n12), .C0(n1055), .Y(
        n1050) );
  AOI22X1 U66 ( .A0(n14), .A1(R0[13]), .B0(n8), .B1(R15[13]), .Y(n1055) );
  OAI221XL U67 ( .A0(n706), .A1(n17), .B0(n604), .B1(n12), .C0(n1039), .Y(
        n1034) );
  AOI22X1 U68 ( .A0(n14), .A1(R0[15]), .B0(n8), .B1(R15[15]), .Y(n1039) );
  OAI221XL U69 ( .A0(n705), .A1(n17), .B0(n603), .B1(n12), .C0(n1031), .Y(
        n1026) );
  AOI22X1 U70 ( .A0(n14), .A1(R0[16]), .B0(n8), .B1(R15[16]), .Y(n1031) );
  OAI221XL U71 ( .A0(n704), .A1(n17), .B0(n602), .B1(n12), .C0(n1023), .Y(
        n1018) );
  AOI22X1 U72 ( .A0(n14), .A1(R0[17]), .B0(n8), .B1(R15[17]), .Y(n1023) );
  OAI221XL U73 ( .A0(n703), .A1(n17), .B0(n601), .B1(n12), .C0(n1015), .Y(
        n1010) );
  AOI22X1 U74 ( .A0(n14), .A1(R0[18]), .B0(n8), .B1(R15[18]), .Y(n1015) );
  OAI221XL U75 ( .A0(n702), .A1(n17), .B0(n600), .B1(n12), .C0(n1007), .Y(
        n1002) );
  AOI22X1 U76 ( .A0(n14), .A1(R0[19]), .B0(n8), .B1(R15[19]), .Y(n1007) );
  OAI221XL U77 ( .A0(n701), .A1(n17), .B0(n599), .B1(n12), .C0(n999), .Y(n994)
         );
  AOI22X1 U78 ( .A0(n14), .A1(R0[20]), .B0(n8), .B1(R15[20]), .Y(n999) );
  OAI221XL U79 ( .A0(n700), .A1(n17), .B0(n598), .B1(n12), .C0(n991), .Y(n986)
         );
  AOI22X1 U80 ( .A0(n14), .A1(R0[21]), .B0(n8), .B1(R15[21]), .Y(n991) );
  OAI221XL U81 ( .A0(n699), .A1(n17), .B0(n597), .B1(n12), .C0(n983), .Y(n978)
         );
  AOI22X1 U82 ( .A0(n14), .A1(R0[22]), .B0(n8), .B1(R15[22]), .Y(n983) );
  OAI221XL U83 ( .A0(n698), .A1(n17), .B0(n596), .B1(n12), .C0(n975), .Y(n970)
         );
  AOI22X1 U84 ( .A0(n14), .A1(R0[23]), .B0(n8), .B1(R15[23]), .Y(n975) );
  OAI221XL U85 ( .A0(n697), .A1(n17), .B0(n595), .B1(n12), .C0(n967), .Y(n962)
         );
  AOI22X1 U86 ( .A0(n14), .A1(R0[24]), .B0(n8), .B1(R15[24]), .Y(n967) );
  OAI221XL U87 ( .A0(n696), .A1(n17), .B0(n594), .B1(n12), .C0(n959), .Y(n954)
         );
  AOI22X1 U88 ( .A0(n14), .A1(R0[25]), .B0(n8), .B1(R15[25]), .Y(n959) );
  OAI221XL U89 ( .A0(n695), .A1(n17), .B0(n593), .B1(n12), .C0(n951), .Y(n946)
         );
  AOI22X1 U90 ( .A0(n14), .A1(R0[26]), .B0(n8), .B1(R15[26]), .Y(n951) );
  OAI221XL U91 ( .A0(n694), .A1(n17), .B0(n592), .B1(n12), .C0(n943), .Y(n938)
         );
  AOI22X1 U92 ( .A0(n14), .A1(R0[27]), .B0(n8), .B1(R15[27]), .Y(n943) );
  OAI221XL U93 ( .A0(n693), .A1(n17), .B0(n591), .B1(n12), .C0(n935), .Y(n930)
         );
  AOI22X1 U94 ( .A0(n14), .A1(R0[28]), .B0(n8), .B1(R15[28]), .Y(n935) );
  OAI221XL U95 ( .A0(n692), .A1(n17), .B0(n590), .B1(n12), .C0(n927), .Y(n922)
         );
  AOI22X1 U96 ( .A0(n14), .A1(R0[29]), .B0(n8), .B1(R15[29]), .Y(n927) );
  OAI221XL U97 ( .A0(n691), .A1(n17), .B0(n589), .B1(n12), .C0(n919), .Y(n914)
         );
  AOI22X1 U98 ( .A0(n14), .A1(R0[30]), .B0(n8), .B1(R15[30]), .Y(n919) );
  OAI221XL U99 ( .A0(n690), .A1(n17), .B0(n588), .B1(n12), .C0(n911), .Y(n906)
         );
  AOI22X1 U100 ( .A0(n14), .A1(R0[31]), .B0(n8), .B1(R15[31]), .Y(n911) );
  OAI221XL U101 ( .A0(n689), .A1(n17), .B0(n587), .B1(n12), .C0(n903), .Y(n898) );
  AOI22X1 U102 ( .A0(n14), .A1(R0[32]), .B0(n8), .B1(R15[32]), .Y(n903) );
  OAI221XL U103 ( .A0(n688), .A1(n17), .B0(n586), .B1(n12), .C0(n890), .Y(n875) );
  AOI22X1 U104 ( .A0(n14), .A1(R0[33]), .B0(n8), .B1(R15[33]), .Y(n890) );
  NOR2X1 U105 ( .A(counter_2[2]), .B(counter_2[1]), .Y(n1160) );
  NOR2X1 U106 ( .A(n862), .B(counter_2[3]), .Y(n1164) );
  NOR2X1 U107 ( .A(counter_2[3]), .B(counter_2[0]), .Y(n1163) );
  AOI22X1 U108 ( .A0(n6), .A1(R2[32]), .B0(n15), .B1(R13[32]), .Y(n901) );
  AOI22X1 U109 ( .A0(n7), .A1(R3[32]), .B0(n16), .B1(R14[32]), .Y(n902) );
  AOI22X1 U110 ( .A0(n1174), .A1(R1[32]), .B0(n9), .B1(R12[32]), .Y(n904) );
  AOI22X1 U111 ( .A0(n6), .A1(R2[33]), .B0(n15), .B1(R13[33]), .Y(n880) );
  AOI22X1 U112 ( .A0(n7), .A1(R3[33]), .B0(n16), .B1(R14[33]), .Y(n885) );
  AOI22X1 U113 ( .A0(n1174), .A1(R1[33]), .B0(n9), .B1(R12[33]), .Y(n895) );
  AOI22X1 U114 ( .A0(n6), .A1(R2[14]), .B0(n15), .B1(R13[14]), .Y(n1045) );
  AOI22X1 U115 ( .A0(n7), .A1(R3[14]), .B0(n16), .B1(R14[14]), .Y(n1046) );
  AOI22X1 U116 ( .A0(n1174), .A1(R1[14]), .B0(n9), .B1(R12[14]), .Y(n1048) );
  OAI221XL U117 ( .A0(n707), .A1(n17), .B0(n605), .B1(n12), .C0(n1047), .Y(
        n1042) );
  AOI22X1 U118 ( .A0(n14), .A1(R0[14]), .B0(n8), .B1(R15[14]), .Y(n1047) );
  NOR2X1 U119 ( .A(n1193), .B(counter_2[2]), .Y(n872) );
  AOI22X1 U120 ( .A0(n6), .A1(R2[0]), .B0(n15), .B1(R13[0]), .Y(n1157) );
  AOI22X1 U121 ( .A0(n7), .A1(R3[0]), .B0(n16), .B1(R14[0]), .Y(n1161) );
  AOI22X1 U122 ( .A0(n1174), .A1(R1[0]), .B0(n9), .B1(R12[0]), .Y(n1165) );
  AOI22X1 U123 ( .A0(n6), .A1(R2[1]), .B0(n15), .B1(R13[1]), .Y(n1149) );
  AOI22X1 U124 ( .A0(n7), .A1(R3[1]), .B0(n16), .B1(R14[1]), .Y(n1150) );
  AOI22X1 U125 ( .A0(n1174), .A1(R1[1]), .B0(n9), .B1(R12[1]), .Y(n1152) );
  AOI22X1 U126 ( .A0(n6), .A1(R2[2]), .B0(n15), .B1(R13[2]), .Y(n1141) );
  AOI22X1 U127 ( .A0(n7), .A1(R3[2]), .B0(n16), .B1(R14[2]), .Y(n1142) );
  AOI22X1 U128 ( .A0(n1174), .A1(R1[2]), .B0(n9), .B1(R12[2]), .Y(n1144) );
  AOI22X1 U129 ( .A0(n6), .A1(R2[3]), .B0(n15), .B1(R13[3]), .Y(n1133) );
  AOI22X1 U130 ( .A0(n7), .A1(R3[3]), .B0(n16), .B1(R14[3]), .Y(n1134) );
  AOI22X1 U131 ( .A0(n1174), .A1(R1[3]), .B0(n9), .B1(R12[3]), .Y(n1136) );
  AOI22X1 U132 ( .A0(n6), .A1(R2[4]), .B0(n15), .B1(R13[4]), .Y(n1125) );
  AOI22X1 U133 ( .A0(n7), .A1(R3[4]), .B0(n16), .B1(R14[4]), .Y(n1126) );
  AOI22X1 U134 ( .A0(n1174), .A1(R1[4]), .B0(n9), .B1(R12[4]), .Y(n1128) );
  AOI22X1 U135 ( .A0(n6), .A1(R2[5]), .B0(n15), .B1(R13[5]), .Y(n1117) );
  AOI22X1 U136 ( .A0(n7), .A1(R3[5]), .B0(n16), .B1(R14[5]), .Y(n1118) );
  AOI22X1 U137 ( .A0(n1174), .A1(R1[5]), .B0(n9), .B1(R12[5]), .Y(n1120) );
  AOI22X1 U138 ( .A0(n6), .A1(R2[6]), .B0(n15), .B1(R13[6]), .Y(n1109) );
  AOI22X1 U139 ( .A0(n7), .A1(R3[6]), .B0(n16), .B1(R14[6]), .Y(n1110) );
  AOI22X1 U140 ( .A0(n1174), .A1(R1[6]), .B0(n9), .B1(R12[6]), .Y(n1112) );
  AOI22X1 U141 ( .A0(n6), .A1(R2[7]), .B0(n15), .B1(R13[7]), .Y(n1101) );
  AOI22X1 U142 ( .A0(n7), .A1(R3[7]), .B0(n16), .B1(R14[7]), .Y(n1102) );
  AOI22X1 U143 ( .A0(n1174), .A1(R1[7]), .B0(n9), .B1(R12[7]), .Y(n1104) );
  AOI22X1 U144 ( .A0(n6), .A1(R2[8]), .B0(n15), .B1(R13[8]), .Y(n1093) );
  AOI22X1 U145 ( .A0(n7), .A1(R3[8]), .B0(n16), .B1(R14[8]), .Y(n1094) );
  AOI22X1 U146 ( .A0(n1174), .A1(R1[8]), .B0(n9), .B1(R12[8]), .Y(n1096) );
  AOI22X1 U147 ( .A0(n6), .A1(R2[9]), .B0(n15), .B1(R13[9]), .Y(n1085) );
  AOI22X1 U148 ( .A0(n7), .A1(R3[9]), .B0(n16), .B1(R14[9]), .Y(n1086) );
  AOI22X1 U149 ( .A0(n1174), .A1(R1[9]), .B0(n9), .B1(R12[9]), .Y(n1088) );
  AOI22X1 U150 ( .A0(n6), .A1(R2[10]), .B0(n15), .B1(R13[10]), .Y(n1077) );
  AOI22X1 U151 ( .A0(n7), .A1(R3[10]), .B0(n16), .B1(R14[10]), .Y(n1078) );
  AOI22X1 U152 ( .A0(n1174), .A1(R1[10]), .B0(n9), .B1(R12[10]), .Y(n1080) );
  AOI22X1 U153 ( .A0(n6), .A1(R2[11]), .B0(n15), .B1(R13[11]), .Y(n1069) );
  AOI22X1 U154 ( .A0(n7), .A1(R3[11]), .B0(n16), .B1(R14[11]), .Y(n1070) );
  AOI22X1 U155 ( .A0(n1174), .A1(R1[11]), .B0(n9), .B1(R12[11]), .Y(n1072) );
  AOI22X1 U156 ( .A0(n6), .A1(R2[12]), .B0(n15), .B1(R13[12]), .Y(n1061) );
  AOI22X1 U157 ( .A0(n7), .A1(R3[12]), .B0(n16), .B1(R14[12]), .Y(n1062) );
  AOI22X1 U158 ( .A0(n1174), .A1(R1[12]), .B0(n9), .B1(R12[12]), .Y(n1064) );
  AOI22X1 U159 ( .A0(n6), .A1(R2[13]), .B0(n15), .B1(R13[13]), .Y(n1053) );
  AOI22X1 U160 ( .A0(n7), .A1(R3[13]), .B0(n16), .B1(R14[13]), .Y(n1054) );
  AOI22X1 U161 ( .A0(n1174), .A1(R1[13]), .B0(n9), .B1(R12[13]), .Y(n1056) );
  AOI22X1 U162 ( .A0(n6), .A1(R2[15]), .B0(n15), .B1(R13[15]), .Y(n1037) );
  AOI22X1 U163 ( .A0(n7), .A1(R3[15]), .B0(n16), .B1(R14[15]), .Y(n1038) );
  AOI22X1 U164 ( .A0(n1174), .A1(R1[15]), .B0(n9), .B1(R12[15]), .Y(n1040) );
  AOI22X1 U165 ( .A0(n6), .A1(R2[16]), .B0(n15), .B1(R13[16]), .Y(n1029) );
  AOI22X1 U166 ( .A0(n7), .A1(R3[16]), .B0(n16), .B1(R14[16]), .Y(n1030) );
  AOI22X1 U167 ( .A0(n1174), .A1(R1[16]), .B0(n9), .B1(R12[16]), .Y(n1032) );
  AOI22X1 U168 ( .A0(n6), .A1(R2[17]), .B0(n15), .B1(R13[17]), .Y(n1021) );
  AOI22X1 U169 ( .A0(n7), .A1(R3[17]), .B0(n16), .B1(R14[17]), .Y(n1022) );
  AOI22X1 U170 ( .A0(n1174), .A1(R1[17]), .B0(n9), .B1(R12[17]), .Y(n1024) );
  AOI22X1 U171 ( .A0(n6), .A1(R2[18]), .B0(n15), .B1(R13[18]), .Y(n1013) );
  AOI22X1 U172 ( .A0(n7), .A1(R3[18]), .B0(n16), .B1(R14[18]), .Y(n1014) );
  AOI22X1 U173 ( .A0(n1174), .A1(R1[18]), .B0(n9), .B1(R12[18]), .Y(n1016) );
  AOI22X1 U174 ( .A0(n6), .A1(R2[19]), .B0(n15), .B1(R13[19]), .Y(n1005) );
  AOI22X1 U175 ( .A0(n7), .A1(R3[19]), .B0(n16), .B1(R14[19]), .Y(n1006) );
  AOI22X1 U176 ( .A0(n1174), .A1(R1[19]), .B0(n9), .B1(R12[19]), .Y(n1008) );
  AOI22X1 U177 ( .A0(n6), .A1(R2[20]), .B0(n15), .B1(R13[20]), .Y(n997) );
  AOI22X1 U178 ( .A0(n7), .A1(R3[20]), .B0(n16), .B1(R14[20]), .Y(n998) );
  AOI22X1 U179 ( .A0(n1174), .A1(R1[20]), .B0(n9), .B1(R12[20]), .Y(n1000) );
  AOI22X1 U180 ( .A0(n6), .A1(R2[21]), .B0(n15), .B1(R13[21]), .Y(n989) );
  AOI22X1 U181 ( .A0(n7), .A1(R3[21]), .B0(n16), .B1(R14[21]), .Y(n990) );
  AOI22X1 U182 ( .A0(n1174), .A1(R1[21]), .B0(n9), .B1(R12[21]), .Y(n992) );
  AOI22X1 U183 ( .A0(n6), .A1(R2[22]), .B0(n15), .B1(R13[22]), .Y(n981) );
  AOI22X1 U184 ( .A0(n7), .A1(R3[22]), .B0(n16), .B1(R14[22]), .Y(n982) );
  AOI22X1 U185 ( .A0(n1174), .A1(R1[22]), .B0(n9), .B1(R12[22]), .Y(n984) );
  AOI22X1 U186 ( .A0(n6), .A1(R2[23]), .B0(n15), .B1(R13[23]), .Y(n973) );
  AOI22X1 U187 ( .A0(n7), .A1(R3[23]), .B0(n16), .B1(R14[23]), .Y(n974) );
  AOI22X1 U188 ( .A0(n1174), .A1(R1[23]), .B0(n9), .B1(R12[23]), .Y(n976) );
  AOI22X1 U189 ( .A0(n6), .A1(R2[24]), .B0(n15), .B1(R13[24]), .Y(n965) );
  AOI22X1 U190 ( .A0(n7), .A1(R3[24]), .B0(n16), .B1(R14[24]), .Y(n966) );
  AOI22X1 U191 ( .A0(n1174), .A1(R1[24]), .B0(n9), .B1(R12[24]), .Y(n968) );
  AOI22X1 U192 ( .A0(n6), .A1(R2[25]), .B0(n15), .B1(R13[25]), .Y(n957) );
  AOI22X1 U193 ( .A0(n7), .A1(R3[25]), .B0(n16), .B1(R14[25]), .Y(n958) );
  AOI22X1 U194 ( .A0(n1174), .A1(R1[25]), .B0(n9), .B1(R12[25]), .Y(n960) );
  AOI22X1 U195 ( .A0(n6), .A1(R2[26]), .B0(n15), .B1(R13[26]), .Y(n949) );
  AOI22X1 U196 ( .A0(n7), .A1(R3[26]), .B0(n16), .B1(R14[26]), .Y(n950) );
  AOI22X1 U197 ( .A0(n1174), .A1(R1[26]), .B0(n9), .B1(R12[26]), .Y(n952) );
  AOI22X1 U198 ( .A0(n6), .A1(R2[27]), .B0(n15), .B1(R13[27]), .Y(n941) );
  AOI22X1 U199 ( .A0(n7), .A1(R3[27]), .B0(n16), .B1(R14[27]), .Y(n942) );
  AOI22X1 U200 ( .A0(n1174), .A1(R1[27]), .B0(n9), .B1(R12[27]), .Y(n944) );
  AOI22X1 U201 ( .A0(n6), .A1(R2[28]), .B0(n15), .B1(R13[28]), .Y(n933) );
  AOI22X1 U202 ( .A0(n7), .A1(R3[28]), .B0(n16), .B1(R14[28]), .Y(n934) );
  AOI22X1 U203 ( .A0(n1174), .A1(R1[28]), .B0(n9), .B1(R12[28]), .Y(n936) );
  AOI22X1 U204 ( .A0(n6), .A1(R2[29]), .B0(n15), .B1(R13[29]), .Y(n925) );
  AOI22X1 U205 ( .A0(n7), .A1(R3[29]), .B0(n16), .B1(R14[29]), .Y(n926) );
  AOI22X1 U206 ( .A0(n1174), .A1(R1[29]), .B0(n9), .B1(R12[29]), .Y(n928) );
  AOI22X1 U207 ( .A0(n6), .A1(R2[30]), .B0(n15), .B1(R13[30]), .Y(n917) );
  AOI22X1 U208 ( .A0(n7), .A1(R3[30]), .B0(n16), .B1(R14[30]), .Y(n918) );
  AOI22X1 U209 ( .A0(n1174), .A1(R1[30]), .B0(n9), .B1(R12[30]), .Y(n920) );
  AOI22X1 U210 ( .A0(n6), .A1(R2[31]), .B0(n15), .B1(R13[31]), .Y(n909) );
  AOI22X1 U211 ( .A0(n7), .A1(R3[31]), .B0(n16), .B1(R14[31]), .Y(n910) );
  AOI22X1 U212 ( .A0(n1174), .A1(R1[31]), .B0(n9), .B1(R12[31]), .Y(n912) );
  OAI221XL U213 ( .A0(n721), .A1(n17), .B0(n619), .B1(n12), .C0(n1162), .Y(
        n1154) );
  AOI22X1 U214 ( .A0(n14), .A1(R0[0]), .B0(n8), .B1(R15[0]), .Y(n1162) );
  OAI221XL U215 ( .A0(n720), .A1(n17), .B0(n618), .B1(n12), .C0(n1151), .Y(
        n1146) );
  AOI22X1 U216 ( .A0(n14), .A1(R0[1]), .B0(n8), .B1(R15[1]), .Y(n1151) );
  OAI221XL U217 ( .A0(n719), .A1(n17), .B0(n617), .B1(n12), .C0(n1143), .Y(
        n1138) );
  AOI22X1 U218 ( .A0(n14), .A1(R0[2]), .B0(n8), .B1(R15[2]), .Y(n1143) );
  OAI221XL U219 ( .A0(n718), .A1(n17), .B0(n616), .B1(n12), .C0(n1135), .Y(
        n1130) );
  AOI22X1 U220 ( .A0(n14), .A1(R0[3]), .B0(n8), .B1(R15[3]), .Y(n1135) );
  OAI221XL U221 ( .A0(n717), .A1(n17), .B0(n615), .B1(n12), .C0(n1127), .Y(
        n1122) );
  AOI22X1 U222 ( .A0(n14), .A1(R0[4]), .B0(n8), .B1(R15[4]), .Y(n1127) );
  OAI221XL U223 ( .A0(n716), .A1(n17), .B0(n614), .B1(n12), .C0(n1119), .Y(
        n1114) );
  AOI22X1 U224 ( .A0(n14), .A1(R0[5]), .B0(n8), .B1(R15[5]), .Y(n1119) );
  OAI221XL U225 ( .A0(n715), .A1(n17), .B0(n613), .B1(n12), .C0(n1111), .Y(
        n1106) );
  AOI22X1 U226 ( .A0(n14), .A1(R0[6]), .B0(n8), .B1(R15[6]), .Y(n1111) );
  OAI221XL U227 ( .A0(n714), .A1(n17), .B0(n612), .B1(n12), .C0(n1103), .Y(
        n1098) );
  AOI22X1 U228 ( .A0(n14), .A1(R0[7]), .B0(n8), .B1(R15[7]), .Y(n1103) );
  OAI221XL U229 ( .A0(n713), .A1(n17), .B0(n611), .B1(n12), .C0(n1095), .Y(
        n1090) );
  AOI22X1 U230 ( .A0(n14), .A1(R0[8]), .B0(n8), .B1(R15[8]), .Y(n1095) );
  OAI221XL U231 ( .A0(n712), .A1(n17), .B0(n610), .B1(n12), .C0(n1087), .Y(
        n1082) );
  AOI22X1 U232 ( .A0(n14), .A1(R0[9]), .B0(n8), .B1(R15[9]), .Y(n1087) );
  AND2X2 U233 ( .A(counter_2[3]), .B(counter_2[0]), .Y(n1159) );
  AND2X2 U234 ( .A(counter_2[3]), .B(n862), .Y(n1158) );
  INVX1 U235 ( .A(p_s_flag_in), .Y(n1195) );
  INVX1 U236 ( .A(counter_2[1]), .Y(n1193) );
  INVX1 U237 ( .A(counter_2[2]), .Y(n1194) );
  AND3X2 U238 ( .A(counter_1[0]), .B(n1195), .C(counter_1[1]), .Y(n125) );
  AND3X2 U239 ( .A(n585), .B(n1195), .C(counter_1[1]), .Y(n126) );
  OR4X2 U240 ( .A(n897), .B(n898), .C(n899), .D(n900), .Y(N151) );
  OAI221XL U241 ( .A0(n757), .A1(n18), .B0(n723), .B1(n13), .C0(n904), .Y(n897) );
  OAI221XL U242 ( .A0(n621), .A1(n10), .B0(n655), .B1(n19), .C0(n902), .Y(n899) );
  OAI221XL U243 ( .A0(n825), .A1(n11), .B0(n791), .B1(n20), .C0(n901), .Y(n900) );
  OR4X2 U244 ( .A(n1041), .B(n1042), .C(n1043), .D(n1044), .Y(N133) );
  OAI221XL U245 ( .A0(n775), .A1(n18), .B0(n741), .B1(n13), .C0(n1048), .Y(
        n1041) );
  OAI221XL U246 ( .A0(n639), .A1(n10), .B0(n673), .B1(n19), .C0(n1046), .Y(
        n1043) );
  OAI221XL U247 ( .A0(n843), .A1(n11), .B0(n809), .B1(n20), .C0(n1045), .Y(
        n1044) );
  OR4X2 U248 ( .A(n874), .B(n875), .C(n876), .D(n877), .Y(N152) );
  OAI221XL U249 ( .A0(n756), .A1(n18), .B0(n722), .B1(n13), .C0(n895), .Y(n874) );
  OAI221XL U250 ( .A0(n620), .A1(n10), .B0(n654), .B1(n19), .C0(n885), .Y(n876) );
  OAI221XL U251 ( .A0(n824), .A1(n11), .B0(n790), .B1(n20), .C0(n880), .Y(n877) );
  OR4X2 U252 ( .A(n1153), .B(n1154), .C(n1155), .D(n1156), .Y(N119) );
  OAI221XL U253 ( .A0(n789), .A1(n18), .B0(n755), .B1(n13), .C0(n1165), .Y(
        n1153) );
  OAI221XL U254 ( .A0(n653), .A1(n10), .B0(n687), .B1(n19), .C0(n1161), .Y(
        n1155) );
  OAI221XL U255 ( .A0(n857), .A1(n11), .B0(n823), .B1(n20), .C0(n1157), .Y(
        n1156) );
  OR4X2 U256 ( .A(n1145), .B(n1146), .C(n1147), .D(n1148), .Y(N120) );
  OAI221XL U257 ( .A0(n788), .A1(n18), .B0(n754), .B1(n13), .C0(n1152), .Y(
        n1145) );
  OAI221XL U258 ( .A0(n652), .A1(n10), .B0(n686), .B1(n19), .C0(n1150), .Y(
        n1147) );
  OAI221XL U259 ( .A0(n856), .A1(n11), .B0(n822), .B1(n20), .C0(n1149), .Y(
        n1148) );
  OR4X2 U260 ( .A(n1137), .B(n1138), .C(n1139), .D(n1140), .Y(N121) );
  OAI221XL U261 ( .A0(n787), .A1(n18), .B0(n753), .B1(n13), .C0(n1144), .Y(
        n1137) );
  OAI221XL U262 ( .A0(n651), .A1(n10), .B0(n685), .B1(n19), .C0(n1142), .Y(
        n1139) );
  OAI221XL U263 ( .A0(n855), .A1(n11), .B0(n821), .B1(n20), .C0(n1141), .Y(
        n1140) );
  OR4X2 U264 ( .A(n1129), .B(n1130), .C(n1131), .D(n1132), .Y(N122) );
  OAI221XL U265 ( .A0(n786), .A1(n18), .B0(n752), .B1(n13), .C0(n1136), .Y(
        n1129) );
  OAI221XL U266 ( .A0(n650), .A1(n10), .B0(n684), .B1(n19), .C0(n1134), .Y(
        n1131) );
  OAI221XL U267 ( .A0(n854), .A1(n11), .B0(n820), .B1(n20), .C0(n1133), .Y(
        n1132) );
  OR4X2 U268 ( .A(n1121), .B(n1122), .C(n1123), .D(n1124), .Y(N123) );
  OAI221XL U269 ( .A0(n785), .A1(n18), .B0(n751), .B1(n13), .C0(n1128), .Y(
        n1121) );
  OAI221XL U270 ( .A0(n649), .A1(n10), .B0(n683), .B1(n19), .C0(n1126), .Y(
        n1123) );
  OAI221XL U271 ( .A0(n853), .A1(n11), .B0(n819), .B1(n20), .C0(n1125), .Y(
        n1124) );
  OR4X2 U272 ( .A(n1113), .B(n1114), .C(n1115), .D(n1116), .Y(N124) );
  OAI221XL U273 ( .A0(n784), .A1(n18), .B0(n750), .B1(n13), .C0(n1120), .Y(
        n1113) );
  OAI221XL U274 ( .A0(n648), .A1(n10), .B0(n682), .B1(n19), .C0(n1118), .Y(
        n1115) );
  OAI221XL U275 ( .A0(n852), .A1(n11), .B0(n818), .B1(n20), .C0(n1117), .Y(
        n1116) );
  OR4X2 U276 ( .A(n1105), .B(n1106), .C(n1107), .D(n1108), .Y(N125) );
  OAI221XL U277 ( .A0(n783), .A1(n18), .B0(n749), .B1(n13), .C0(n1112), .Y(
        n1105) );
  OAI221XL U278 ( .A0(n647), .A1(n10), .B0(n681), .B1(n19), .C0(n1110), .Y(
        n1107) );
  OAI221XL U279 ( .A0(n851), .A1(n11), .B0(n817), .B1(n20), .C0(n1109), .Y(
        n1108) );
  OR4X2 U280 ( .A(n1097), .B(n1098), .C(n1099), .D(n1100), .Y(N126) );
  OAI221XL U281 ( .A0(n782), .A1(n18), .B0(n748), .B1(n13), .C0(n1104), .Y(
        n1097) );
  OAI221XL U282 ( .A0(n646), .A1(n10), .B0(n680), .B1(n19), .C0(n1102), .Y(
        n1099) );
  OAI221XL U283 ( .A0(n850), .A1(n11), .B0(n816), .B1(n20), .C0(n1101), .Y(
        n1100) );
  OR4X2 U284 ( .A(n1089), .B(n1090), .C(n1091), .D(n1092), .Y(N127) );
  OAI221XL U285 ( .A0(n781), .A1(n18), .B0(n747), .B1(n13), .C0(n1096), .Y(
        n1089) );
  OAI221XL U286 ( .A0(n645), .A1(n10), .B0(n679), .B1(n19), .C0(n1094), .Y(
        n1091) );
  OAI221XL U287 ( .A0(n849), .A1(n11), .B0(n815), .B1(n20), .C0(n1093), .Y(
        n1092) );
  OR4X2 U288 ( .A(n1081), .B(n1082), .C(n1083), .D(n1084), .Y(N128) );
  OAI221XL U289 ( .A0(n780), .A1(n18), .B0(n746), .B1(n13), .C0(n1088), .Y(
        n1081) );
  OAI221XL U290 ( .A0(n644), .A1(n10), .B0(n678), .B1(n19), .C0(n1086), .Y(
        n1083) );
  OAI221XL U291 ( .A0(n848), .A1(n11), .B0(n814), .B1(n20), .C0(n1085), .Y(
        n1084) );
  OR4X2 U292 ( .A(n1073), .B(n1074), .C(n1075), .D(n1076), .Y(N129) );
  OAI221XL U293 ( .A0(n779), .A1(n18), .B0(n745), .B1(n13), .C0(n1080), .Y(
        n1073) );
  OAI221XL U294 ( .A0(n643), .A1(n10), .B0(n677), .B1(n19), .C0(n1078), .Y(
        n1075) );
  OAI221XL U295 ( .A0(n847), .A1(n11), .B0(n813), .B1(n20), .C0(n1077), .Y(
        n1076) );
  OR4X2 U296 ( .A(n1065), .B(n1066), .C(n1067), .D(n1068), .Y(N130) );
  OAI221XL U297 ( .A0(n778), .A1(n18), .B0(n744), .B1(n13), .C0(n1072), .Y(
        n1065) );
  OAI221XL U298 ( .A0(n642), .A1(n10), .B0(n676), .B1(n19), .C0(n1070), .Y(
        n1067) );
  OAI221XL U299 ( .A0(n846), .A1(n11), .B0(n812), .B1(n20), .C0(n1069), .Y(
        n1068) );
  OR4X2 U300 ( .A(n1057), .B(n1058), .C(n1059), .D(n1060), .Y(N131) );
  OAI221XL U301 ( .A0(n777), .A1(n18), .B0(n743), .B1(n13), .C0(n1064), .Y(
        n1057) );
  OAI221XL U302 ( .A0(n641), .A1(n10), .B0(n675), .B1(n19), .C0(n1062), .Y(
        n1059) );
  OAI221XL U303 ( .A0(n845), .A1(n11), .B0(n811), .B1(n20), .C0(n1061), .Y(
        n1060) );
  OR4X2 U304 ( .A(n1049), .B(n1050), .C(n1051), .D(n1052), .Y(N132) );
  OAI221XL U305 ( .A0(n776), .A1(n18), .B0(n742), .B1(n13), .C0(n1056), .Y(
        n1049) );
  OAI221XL U306 ( .A0(n640), .A1(n10), .B0(n674), .B1(n19), .C0(n1054), .Y(
        n1051) );
  OAI221XL U307 ( .A0(n844), .A1(n11), .B0(n810), .B1(n20), .C0(n1053), .Y(
        n1052) );
  OR4X2 U308 ( .A(n1033), .B(n1034), .C(n1035), .D(n1036), .Y(N134) );
  OAI221XL U309 ( .A0(n774), .A1(n18), .B0(n740), .B1(n13), .C0(n1040), .Y(
        n1033) );
  OAI221XL U310 ( .A0(n638), .A1(n10), .B0(n672), .B1(n19), .C0(n1038), .Y(
        n1035) );
  OAI221XL U311 ( .A0(n842), .A1(n11), .B0(n808), .B1(n20), .C0(n1037), .Y(
        n1036) );
  OR4X2 U312 ( .A(n1025), .B(n1026), .C(n1027), .D(n1028), .Y(N135) );
  OAI221XL U313 ( .A0(n773), .A1(n18), .B0(n739), .B1(n13), .C0(n1032), .Y(
        n1025) );
  OAI221XL U314 ( .A0(n637), .A1(n10), .B0(n671), .B1(n19), .C0(n1030), .Y(
        n1027) );
  OAI221XL U315 ( .A0(n841), .A1(n11), .B0(n807), .B1(n20), .C0(n1029), .Y(
        n1028) );
  OR4X2 U316 ( .A(n1017), .B(n1018), .C(n1019), .D(n1020), .Y(N136) );
  OAI221XL U317 ( .A0(n772), .A1(n18), .B0(n738), .B1(n13), .C0(n1024), .Y(
        n1017) );
  OAI221XL U318 ( .A0(n636), .A1(n10), .B0(n670), .B1(n19), .C0(n1022), .Y(
        n1019) );
  OAI221XL U319 ( .A0(n840), .A1(n11), .B0(n806), .B1(n20), .C0(n1021), .Y(
        n1020) );
  OR4X2 U320 ( .A(n1009), .B(n1010), .C(n1011), .D(n1012), .Y(N137) );
  OAI221XL U321 ( .A0(n771), .A1(n18), .B0(n737), .B1(n13), .C0(n1016), .Y(
        n1009) );
  OAI221XL U322 ( .A0(n635), .A1(n10), .B0(n669), .B1(n19), .C0(n1014), .Y(
        n1011) );
  OAI221XL U323 ( .A0(n839), .A1(n11), .B0(n805), .B1(n20), .C0(n1013), .Y(
        n1012) );
  OR4X2 U324 ( .A(n1001), .B(n1002), .C(n1003), .D(n1004), .Y(N138) );
  OAI221XL U325 ( .A0(n770), .A1(n18), .B0(n736), .B1(n13), .C0(n1008), .Y(
        n1001) );
  OAI221XL U326 ( .A0(n634), .A1(n10), .B0(n668), .B1(n19), .C0(n1006), .Y(
        n1003) );
  OAI221XL U327 ( .A0(n838), .A1(n11), .B0(n804), .B1(n20), .C0(n1005), .Y(
        n1004) );
  OR4X2 U328 ( .A(n993), .B(n994), .C(n995), .D(n996), .Y(N139) );
  OAI221XL U329 ( .A0(n769), .A1(n18), .B0(n735), .B1(n13), .C0(n1000), .Y(
        n993) );
  OAI221XL U330 ( .A0(n633), .A1(n10), .B0(n667), .B1(n19), .C0(n998), .Y(n995) );
  OAI221XL U331 ( .A0(n837), .A1(n11), .B0(n803), .B1(n20), .C0(n997), .Y(n996) );
  OR4X2 U332 ( .A(n985), .B(n986), .C(n987), .D(n988), .Y(N140) );
  OAI221XL U333 ( .A0(n768), .A1(n18), .B0(n734), .B1(n13), .C0(n992), .Y(n985) );
  OAI221XL U334 ( .A0(n632), .A1(n10), .B0(n666), .B1(n19), .C0(n990), .Y(n987) );
  OAI221XL U335 ( .A0(n836), .A1(n11), .B0(n802), .B1(n20), .C0(n989), .Y(n988) );
  OR4X2 U336 ( .A(n977), .B(n978), .C(n979), .D(n980), .Y(N141) );
  OAI221XL U337 ( .A0(n767), .A1(n18), .B0(n733), .B1(n13), .C0(n984), .Y(n977) );
  OAI221XL U338 ( .A0(n631), .A1(n10), .B0(n665), .B1(n19), .C0(n982), .Y(n979) );
  OAI221XL U339 ( .A0(n835), .A1(n11), .B0(n801), .B1(n20), .C0(n981), .Y(n980) );
  OR4X2 U340 ( .A(n969), .B(n970), .C(n971), .D(n972), .Y(N142) );
  OAI221XL U341 ( .A0(n766), .A1(n18), .B0(n732), .B1(n13), .C0(n976), .Y(n969) );
  OAI221XL U342 ( .A0(n630), .A1(n10), .B0(n664), .B1(n19), .C0(n974), .Y(n971) );
  OAI221XL U343 ( .A0(n834), .A1(n11), .B0(n800), .B1(n20), .C0(n973), .Y(n972) );
  OR4X2 U344 ( .A(n961), .B(n962), .C(n963), .D(n964), .Y(N143) );
  OAI221XL U345 ( .A0(n765), .A1(n18), .B0(n731), .B1(n13), .C0(n968), .Y(n961) );
  OAI221XL U346 ( .A0(n629), .A1(n10), .B0(n663), .B1(n19), .C0(n966), .Y(n963) );
  OAI221XL U347 ( .A0(n833), .A1(n11), .B0(n799), .B1(n20), .C0(n965), .Y(n964) );
  OR4X2 U348 ( .A(n953), .B(n954), .C(n955), .D(n956), .Y(N144) );
  OAI221XL U349 ( .A0(n764), .A1(n18), .B0(n730), .B1(n13), .C0(n960), .Y(n953) );
  OAI221XL U350 ( .A0(n628), .A1(n10), .B0(n662), .B1(n19), .C0(n958), .Y(n955) );
  OAI221XL U351 ( .A0(n832), .A1(n11), .B0(n798), .B1(n20), .C0(n957), .Y(n956) );
  OR4X2 U352 ( .A(n945), .B(n946), .C(n947), .D(n948), .Y(N145) );
  OAI221XL U353 ( .A0(n763), .A1(n18), .B0(n729), .B1(n13), .C0(n952), .Y(n945) );
  OAI221XL U354 ( .A0(n627), .A1(n10), .B0(n661), .B1(n19), .C0(n950), .Y(n947) );
  OAI221XL U355 ( .A0(n831), .A1(n11), .B0(n797), .B1(n20), .C0(n949), .Y(n948) );
  OR4X2 U356 ( .A(n937), .B(n938), .C(n939), .D(n940), .Y(N146) );
  OAI221XL U357 ( .A0(n762), .A1(n18), .B0(n728), .B1(n13), .C0(n944), .Y(n937) );
  OAI221XL U358 ( .A0(n626), .A1(n10), .B0(n660), .B1(n19), .C0(n942), .Y(n939) );
  OAI221XL U359 ( .A0(n830), .A1(n11), .B0(n796), .B1(n20), .C0(n941), .Y(n940) );
  OR4X2 U360 ( .A(n929), .B(n930), .C(n931), .D(n932), .Y(N147) );
  OAI221XL U361 ( .A0(n761), .A1(n18), .B0(n727), .B1(n13), .C0(n936), .Y(n929) );
  OAI221XL U362 ( .A0(n625), .A1(n10), .B0(n659), .B1(n19), .C0(n934), .Y(n931) );
  OAI221XL U363 ( .A0(n829), .A1(n11), .B0(n795), .B1(n20), .C0(n933), .Y(n932) );
  OR4X2 U364 ( .A(n921), .B(n922), .C(n923), .D(n924), .Y(N148) );
  OAI221XL U365 ( .A0(n760), .A1(n18), .B0(n726), .B1(n13), .C0(n928), .Y(n921) );
  OAI221XL U366 ( .A0(n624), .A1(n10), .B0(n658), .B1(n19), .C0(n926), .Y(n923) );
  OAI221XL U367 ( .A0(n828), .A1(n11), .B0(n794), .B1(n20), .C0(n925), .Y(n924) );
  OR4X2 U368 ( .A(n913), .B(n914), .C(n915), .D(n916), .Y(N149) );
  OAI221XL U369 ( .A0(n759), .A1(n18), .B0(n725), .B1(n13), .C0(n920), .Y(n913) );
  OAI221XL U370 ( .A0(n623), .A1(n10), .B0(n657), .B1(n19), .C0(n918), .Y(n915) );
  OAI221XL U371 ( .A0(n827), .A1(n11), .B0(n793), .B1(n20), .C0(n917), .Y(n916) );
  OR4X2 U372 ( .A(n905), .B(n906), .C(n907), .D(n908), .Y(N150) );
  OAI221XL U373 ( .A0(n758), .A1(n18), .B0(n724), .B1(n13), .C0(n912), .Y(n905) );
  OAI221XL U374 ( .A0(n622), .A1(n10), .B0(n656), .B1(n19), .C0(n910), .Y(n907) );
  OAI221XL U375 ( .A0(n826), .A1(n11), .B0(n792), .B1(n20), .C0(n909), .Y(n908) );
  NAND2X1 U376 ( .A(n868), .B(n869), .Y(N52) );
  OAI2BB1X1 U377 ( .A0N(n870), .A1N(counter_2[0]), .B0(counter_2[3]), .Y(n869)
         );
  XNOR2X1 U378 ( .A(counter_1[1]), .B(n585), .Y(N26) );
  XNOR2X1 U379 ( .A(n1193), .B(counter_2[0]), .Y(N50) );
  INVX1 U380 ( .A(n871), .Y(n1192) );
  AOI221X1 U381 ( .A0(counter_2[0]), .A1(n872), .B0(n862), .B1(counter_2[2]), 
        .C0(n873), .Y(n871) );
endmodule


module fft ( clk, rst_n, data_in, data_out );
  input [33:0] data_in;
  output [33:0] data_out;
  input clk, rst_n;
  wire   s_p_flag, mux_flag, demux_flag, n1, n2, n3, n4, n5;
  wire   [2:0] rotation;
  wire   [135:0] data_1;
  wire   [135:0] data_2;
  wire   [135:0] data_4;
  wire   [135:0] data_3;

  ctrl ctrl0 ( .clk(clk), .rst_n(rst_n), .s_p_flag_in(s_p_flag), .mux_flag(
        mux_flag), .rotation(rotation), .demux_flag(demux_flag) );
  s_p s_p0 ( .clk(clk), .rst_n(rst_n), .data_in_1(data_in), .data_out_1(data_1), .s_p_flag_out(s_p_flag) );
  mux mux0 ( .mux_flag(n4), .clk(clk), .rst_n(rst_n), .data_in_1(data_2), 
        .data_in_2(data_1), .data_out(data_3), .data_in_3_33_(data_4[33]), 
        .data_in_3_32_(data_4[32]), .data_in_3_31_(n3), .data_in_3_30_(
        data_4[30]), .data_in_3_29_(data_4[29]), .data_in_3_28_(data_4[28]), 
        .data_in_3_27_(data_4[27]), .data_in_3_26_(data_4[26]), 
        .data_in_3_25_(data_4[25]), .data_in_3_24_(data_4[24]), 
        .data_in_3_23_(data_4[23]), .data_in_3_22_(data_4[22]), 
        .data_in_3_21_(data_4[21]), .data_in_3_20_(data_4[20]), 
        .data_in_3_19_(data_4[19]), .data_in_3_18_(data_4[18]), 
        .data_in_3_17_(data_4[17]), .data_in_3_16_(data_4[16]), 
        .data_in_3_15_(data_4[15]), .data_in_3_14_(data_4[14]), 
        .data_in_3_13_(data_4[13]), .data_in_3_12_(data_4[12]), 
        .data_in_3_11_(data_4[11]), .data_in_3_10_(data_4[10]), .data_in_3_9_(
        data_4[9]), .data_in_3_8_(data_4[8]), .data_in_3_7_(data_4[7]), 
        .data_in_3_6_(data_4[6]), .data_in_3_5_(data_4[5]), .data_in_3_4_(
        data_4[4]), .data_in_3_3_(data_4[3]), .data_in_3_2_(data_4[2]), 
        .data_in_3_1_(data_4[1]), .data_in_3_0_(data_4[0]) );
  butterfly butterfly0 ( .calc_in(data_3), .rotation(rotation), .calc_out(
        data_4) );
  reg1 reg10 ( .clk(clk), .rst_n(rst_n), .data_in_2({data_4[135:32], n3, 
        data_4[30:0]}), .reg_datain_flag(demux_flag), .data_out_2(data_2) );
  p_s p_s0 ( .clk(clk), .rst_n(rst_n), .data_in_3({data_4[135:102], n1, 
        data_4[100:32], n3, data_4[30:0]}), .p_s_flag_in(demux_flag), 
        .data_out_3(data_out) );
  INVX8 U1 ( .A(n5), .Y(n4) );
  CLKINVX3 U2 ( .A(data_4[31]), .Y(n2) );
  CLKBUFX3 U3 ( .A(data_4[101]), .Y(n1) );
  INVX4 U4 ( .A(n2), .Y(n3) );
  INVX4 U5 ( .A(mux_flag), .Y(n5) );
endmodule


module fft_chip ( clk, rstn, din, dout );
  input [33:0] din;
  output [33:0] dout;
  input clk, rstn;
  wire   net_clk, net_rstn;
  wire   [33:0] net_din;
  wire   [33:0] net_dout;

  PIW PIW_clk ( .PAD(clk), .C(net_clk) );
  PIW PIW_rstn ( .PAD(rstn), .C(net_rstn) );
  PIW PIW_din0 ( .PAD(din[0]), .C(net_din[0]) );
  PIW PIW_din1 ( .PAD(din[1]), .C(net_din[1]) );
  PIW PIW_din2 ( .PAD(din[2]), .C(net_din[2]) );
  PIW PIW_din3 ( .PAD(din[3]), .C(net_din[3]) );
  PIW PIW_din4 ( .PAD(din[4]), .C(net_din[4]) );
  PIW PIW_din5 ( .PAD(din[5]), .C(net_din[5]) );
  PIW PIW_din6 ( .PAD(din[6]), .C(net_din[6]) );
  PIW PIW_din7 ( .PAD(din[7]), .C(net_din[7]) );
  PIW PIW_din8 ( .PAD(din[8]), .C(net_din[8]) );
  PIW PIW_din9 ( .PAD(din[9]), .C(net_din[9]) );
  PIW PIW_din10 ( .PAD(din[10]), .C(net_din[10]) );
  PIW PIW_din11 ( .PAD(din[11]), .C(net_din[11]) );
  PIW PIW_din12 ( .PAD(din[12]), .C(net_din[12]) );
  PIW PIW_din13 ( .PAD(din[13]), .C(net_din[13]) );
  PIW PIW_din14 ( .PAD(din[14]), .C(net_din[14]) );
  PIW PIW_din15 ( .PAD(din[15]), .C(net_din[15]) );
  PIW PIW_din16 ( .PAD(din[16]), .C(net_din[16]) );
  PIW PIW_din17 ( .PAD(din[17]), .C(net_din[17]) );
  PIW PIW_din18 ( .PAD(din[18]), .C(net_din[18]) );
  PIW PIW_din19 ( .PAD(din[19]), .C(net_din[19]) );
  PIW PIW_din20 ( .PAD(din[20]), .C(net_din[20]) );
  PIW PIW_din21 ( .PAD(din[21]), .C(net_din[21]) );
  PIW PIW_din22 ( .PAD(din[22]), .C(net_din[22]) );
  PIW PIW_din23 ( .PAD(din[23]), .C(net_din[23]) );
  PIW PIW_din24 ( .PAD(din[24]), .C(net_din[24]) );
  PIW PIW_din25 ( .PAD(din[25]), .C(net_din[25]) );
  PIW PIW_din26 ( .PAD(din[26]), .C(net_din[26]) );
  PIW PIW_din27 ( .PAD(din[27]), .C(net_din[27]) );
  PIW PIW_din28 ( .PAD(din[28]), .C(net_din[28]) );
  PIW PIW_din29 ( .PAD(din[29]), .C(net_din[29]) );
  PIW PIW_din30 ( .PAD(din[30]), .C(net_din[30]) );
  PIW PIW_din31 ( .PAD(din[31]), .C(net_din[31]) );
  PIW PIW_din32 ( .PAD(din[32]), .C(net_din[32]) );
  PIW PIW_din33 ( .PAD(din[33]), .C(net_din[33]) );
  PO8W PO8W_dout0 ( .I(net_dout[0]), .PAD(dout[0]) );
  PO8W PO8W_dout1 ( .I(net_dout[1]), .PAD(dout[1]) );
  PO8W PO8W_dout2 ( .I(net_dout[2]), .PAD(dout[2]) );
  PO8W PO8W_dout3 ( .I(net_dout[3]), .PAD(dout[3]) );
  PO8W PO8W_dout4 ( .I(net_dout[4]), .PAD(dout[4]) );
  PO8W PO8W_dout5 ( .I(net_dout[5]), .PAD(dout[5]) );
  PO8W PO8W_dout6 ( .I(net_dout[6]), .PAD(dout[6]) );
  PO8W PO8W_dout7 ( .I(net_dout[7]), .PAD(dout[7]) );
  PO8W PO8W_dout8 ( .I(net_dout[8]), .PAD(dout[8]) );
  PO8W PO8W_dout9 ( .I(net_dout[9]), .PAD(dout[9]) );
  PO8W PO8W_dout10 ( .I(net_dout[10]), .PAD(dout[10]) );
  PO8W PO8W_dout11 ( .I(net_dout[11]), .PAD(dout[11]) );
  PO8W PO8W_dout12 ( .I(net_dout[12]), .PAD(dout[12]) );
  PO8W PO8W_dout13 ( .I(net_dout[13]), .PAD(dout[13]) );
  PO8W PO8W_dout14 ( .I(net_dout[14]), .PAD(dout[14]) );
  PO8W PO8W_dout15 ( .I(net_dout[15]), .PAD(dout[15]) );
  PO8W PO8W_dout16 ( .I(net_dout[16]), .PAD(dout[16]) );
  PO8W PO8W_dout17 ( .I(net_dout[17]), .PAD(dout[17]) );
  PO8W PO8W_dout18 ( .I(net_dout[18]), .PAD(dout[18]) );
  PO8W PO8W_dout19 ( .I(net_dout[19]), .PAD(dout[19]) );
  PO8W PO8W_dout20 ( .I(net_dout[20]), .PAD(dout[20]) );
  PO8W PO8W_dout21 ( .I(net_dout[21]), .PAD(dout[21]) );
  PO8W PO8W_dout22 ( .I(net_dout[22]), .PAD(dout[22]) );
  PO8W PO8W_dout23 ( .I(net_dout[23]), .PAD(dout[23]) );
  PO8W PO8W_dout24 ( .I(net_dout[24]), .PAD(dout[24]) );
  PO8W PO8W_dout25 ( .I(net_dout[25]), .PAD(dout[25]) );
  PO8W PO8W_dout26 ( .I(net_dout[26]), .PAD(dout[26]) );
  PO8W PO8W_dout27 ( .I(net_dout[27]), .PAD(dout[27]) );
  PO8W PO8W_dout28 ( .I(net_dout[28]), .PAD(dout[28]) );
  PO8W PO8W_dout29 ( .I(net_dout[29]), .PAD(dout[29]) );
  PO8W PO8W_dout30 ( .I(net_dout[30]), .PAD(dout[30]) );
  PO8W PO8W_dout31 ( .I(net_dout[31]), .PAD(dout[31]) );
  PO8W PO8W_dout32 ( .I(net_dout[32]), .PAD(dout[32]) );
  PO8W PO8W_dout33 ( .I(net_dout[33]), .PAD(dout[33]) );
  fft inst_fft ( .clk(net_clk), .rst_n(net_rstn), .data_in(net_din), 
        .data_out(net_dout) );
endmodule

