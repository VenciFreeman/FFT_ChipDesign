
module s2p_0 ( clk, rstn, start, mode, din, dout, s2p_ready, mode_out );
  input [1:0] mode;
  input [15:0] din;
  output [255:0] dout;
  output [1:0] mode_out;
  input clk, rstn, start;
  output s2p_ready;
  wire   N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43,
         N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57,
         N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71,
         N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85,
         N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99,
         N100, N101, N102, N103, N104, N105, N106, N107, N108, N109, N110,
         N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121,
         N122, N123, N124, N125, N126, N127, N128, N129, N131, N132, N133,
         N134, N135, N136, N137, N138, N139, N140, N141, N142, N143, N144,
         N145, N146, N147, N148, N149, N150, N151, N152, N153, N154, N155,
         N156, N157, N158, N159, N160, N161, N162, N163, N164, N165, N166,
         N167, N168, N169, N170, N171, N172, N173, N174, N175, N176, N177,
         N178, N179, N180, N181, N182, N183, N184, N185, N186, N187, N188,
         N189, N190, N191, N192, N193, N194, N195, N196, N197, N198, N199,
         N200, N201, N202, N203, N204, N205, N206, N207, N208, N209, N210,
         N211, N212, N213, N214, N215, N216, N217, N218, N219, N220, N221,
         N222, N223, N224, N225, N226, N227, N228, N229, N231, N232, N233,
         N234, N235, N236, N237, N238, N239, N240, N241, N242, N243, N244,
         N245, N246, N247, N248, N249, N250, N251, N252, N253, N254, N255,
         N256, N257, N258, N259, N260, N261, N262, N263, N264, N265, N266,
         N267, N268, N269, N270, N271, N272, N273, N274, N275, N276, N277,
         N278, N279, N280, N281, N282, N283, N284, N285, N286, N287, N288,
         N302, N303, N304, N1114, N1115, N1116, N1117, N1118, N1119, n731,
         n733, n734, n736, n737, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
         n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
         n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
         n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
         n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
         n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
         n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
         n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
         n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
         n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1, n2,
         n3, n4, n5, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n732, n735,
         n738, n739, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
         n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
         n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
         n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
         n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
         n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
         n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
         n1267, n1268, n1269;
  wire   [1:0] mode_reg;
  wire   [63:0] dout4_reg;
  wire   [127:0] dout8_reg;
  wire   [255:0] dout16_reg;
  wire   [4:0] count;
  wire   [4:2] r71_carry;

  OAI2BB2X4 U3 ( .B0(n333), .B1(n335), .A0N(n335), .A1N(mode_out[0]), .Y(
        mode_out[0]) );
  OAI2BB2X4 U4 ( .B0(n335), .B1(n332), .A0N(n335), .A1N(mode_out[1]), .Y(
        mode_out[1]) );
  TLATX1 dout_reg_16_ ( .G(n327), .D(N47), .Q(dout[16]) );
  TLATX1 dout_reg_111_ ( .G(n319), .D(N143), .Q(dout[111]) );
  TLATX1 dout_reg_79_ ( .G(n318), .D(N110), .Q(dout[79]) );
  TLATX1 dout_reg_47_ ( .G(n328), .D(N78), .Q(dout[47]) );
  TLATX1 dout_reg_31_ ( .G(n326), .D(N62), .Q(dout[31]) );
  TLATX1 dout_reg_110_ ( .G(N30), .D(N142), .Q(dout[110]) );
  TLATX1 dout_reg_78_ ( .G(n318), .D(N109), .Q(dout[78]) );
  TLATX1 dout_reg_46_ ( .G(n322), .D(N77), .Q(dout[46]) );
  TLATX1 dout_reg_30_ ( .G(n322), .D(N61), .Q(dout[30]) );
  TLATX1 dout_reg_109_ ( .G(n326), .D(N141), .Q(dout[109]) );
  TLATX1 dout_reg_77_ ( .G(N30), .D(N108), .Q(dout[77]) );
  TLATX1 dout_reg_45_ ( .G(n318), .D(N76), .Q(dout[45]) );
  TLATX1 dout_reg_29_ ( .G(n328), .D(N60), .Q(dout[29]) );
  TLATX1 dout_reg_108_ ( .G(n330), .D(N140), .Q(dout[108]) );
  TLATX1 dout_reg_76_ ( .G(n324), .D(N107), .Q(dout[76]) );
  TLATX1 dout_reg_44_ ( .G(n328), .D(N75), .Q(dout[44]) );
  TLATX1 dout_reg_28_ ( .G(n326), .D(N59), .Q(dout[28]) );
  TLATX1 dout_reg_107_ ( .G(N30), .D(N139), .Q(dout[107]) );
  TLATX1 dout_reg_75_ ( .G(n318), .D(N106), .Q(dout[75]) );
  TLATX1 dout_reg_43_ ( .G(n330), .D(N74), .Q(dout[43]) );
  TLATX1 dout_reg_27_ ( .G(n324), .D(N58), .Q(dout[27]) );
  TLATX1 dout_reg_106_ ( .G(n323), .D(N138), .Q(dout[106]) );
  TLATX1 dout_reg_74_ ( .G(n321), .D(N105), .Q(dout[74]) );
  TLATX1 dout_reg_42_ ( .G(n329), .D(N73), .Q(dout[42]) );
  TLATX1 dout_reg_26_ ( .G(n320), .D(N57), .Q(dout[26]) );
  TLATX1 dout_reg_105_ ( .G(N30), .D(N137), .Q(dout[105]) );
  TLATX1 dout_reg_73_ ( .G(N30), .D(N104), .Q(dout[73]) );
  TLATX1 dout_reg_41_ ( .G(n327), .D(N72), .Q(dout[41]) );
  TLATX1 dout_reg_25_ ( .G(n325), .D(N56), .Q(dout[25]) );
  TLATX1 dout_reg_104_ ( .G(n322), .D(N136), .Q(dout[104]) );
  TLATX1 dout_reg_72_ ( .G(n328), .D(N103), .Q(dout[72]) );
  TLATX1 dout_reg_40_ ( .G(n326), .D(N71), .Q(dout[40]) );
  TLATX1 dout_reg_24_ ( .G(N30), .D(N55), .Q(dout[24]) );
  TLATX1 dout_reg_103_ ( .G(n330), .D(N135), .Q(dout[103]) );
  TLATX1 dout_reg_71_ ( .G(n330), .D(N102), .Q(dout[71]) );
  TLATX1 dout_reg_39_ ( .G(n330), .D(N70), .Q(dout[39]) );
  TLATX1 dout_reg_23_ ( .G(n330), .D(N54), .Q(dout[23]) );
  TLATX1 dout_reg_102_ ( .G(n330), .D(N134), .Q(dout[102]) );
  TLATX1 dout_reg_70_ ( .G(n330), .D(N101), .Q(dout[70]) );
  TLATX1 dout_reg_38_ ( .G(n320), .D(N69), .Q(dout[38]) );
  TLATX1 dout_reg_22_ ( .G(n327), .D(N53), .Q(dout[22]) );
  TLATX1 dout_reg_101_ ( .G(n325), .D(N133), .Q(dout[101]) );
  TLATX1 dout_reg_69_ ( .G(n322), .D(N100), .Q(dout[69]) );
  TLATX1 dout_reg_37_ ( .G(n328), .D(N68), .Q(dout[37]) );
  TLATX1 dout_reg_21_ ( .G(n326), .D(N52), .Q(dout[21]) );
  TLATX1 dout_reg_100_ ( .G(n329), .D(N132), .Q(dout[100]) );
  TLATX1 dout_reg_68_ ( .G(n329), .D(N99), .Q(dout[68]) );
  TLATX1 dout_reg_36_ ( .G(n329), .D(N67), .Q(dout[36]) );
  TLATX1 dout_reg_20_ ( .G(n329), .D(N51), .Q(dout[20]) );
  TLATX1 dout_reg_99_ ( .G(n329), .D(N131), .Q(dout[99]) );
  TLATX1 dout_reg_67_ ( .G(n329), .D(N98), .Q(dout[67]) );
  TLATX1 dout_reg_35_ ( .G(n328), .D(N66), .Q(dout[35]) );
  TLATX1 dout_reg_19_ ( .G(n328), .D(N50), .Q(dout[19]) );
  TLATX1 dout_reg_98_ ( .G(n328), .D(N129), .Q(dout[98]) );
  TLATX1 dout_reg_66_ ( .G(n328), .D(N97), .Q(dout[66]) );
  TLATX1 dout_reg_34_ ( .G(n328), .D(N65), .Q(dout[34]) );
  TLATX1 dout_reg_18_ ( .G(n328), .D(N49), .Q(dout[18]) );
  TLATX1 dout_reg_97_ ( .G(n327), .D(N128), .Q(dout[97]) );
  TLATX1 dout_reg_65_ ( .G(n327), .D(N96), .Q(dout[65]) );
  TLATX1 dout_reg_33_ ( .G(n327), .D(N64), .Q(dout[33]) );
  TLATX1 dout_reg_17_ ( .G(n327), .D(N48), .Q(dout[17]) );
  TLATX1 dout_reg_96_ ( .G(n327), .D(N127), .Q(dout[96]) );
  TLATX1 dout_reg_64_ ( .G(n327), .D(N95), .Q(dout[64]) );
  TLATX1 dout_reg_32_ ( .G(n325), .D(N63), .Q(dout[32]) );
  TLATX1 dout_reg_143_ ( .G(n322), .D(N175), .Q(dout[143]) );
  TLATX1 dout_reg_142_ ( .G(n328), .D(N174), .Q(dout[142]) );
  TLATX1 dout_reg_141_ ( .G(n326), .D(N173), .Q(dout[141]) );
  TLATX1 dout_reg_140_ ( .G(n326), .D(N172), .Q(dout[140]) );
  TLATX1 dout_reg_139_ ( .G(n326), .D(N171), .Q(dout[139]) );
  TLATX1 dout_reg_138_ ( .G(n325), .D(N170), .Q(dout[138]) );
  TLATX1 dout_reg_137_ ( .G(n325), .D(N169), .Q(dout[137]) );
  TLATX1 dout_reg_136_ ( .G(n325), .D(N168), .Q(dout[136]) );
  TLATX1 dout_reg_135_ ( .G(n324), .D(N167), .Q(dout[135]) );
  TLATX1 dout_reg_134_ ( .G(n324), .D(N166), .Q(dout[134]) );
  TLATX1 dout_reg_133_ ( .G(n324), .D(N165), .Q(dout[133]) );
  TLATX1 dout_reg_132_ ( .G(n323), .D(N164), .Q(dout[132]) );
  TLATX1 dout_reg_131_ ( .G(n323), .D(N163), .Q(dout[131]) );
  TLATX1 dout_reg_130_ ( .G(n323), .D(N162), .Q(dout[130]) );
  TLATX1 dout_reg_129_ ( .G(n322), .D(N161), .Q(dout[129]) );
  TLATX1 dout_reg_128_ ( .G(n322), .D(N160), .Q(dout[128]) );
  TLATX1 dout_reg_15_ ( .G(n330), .D(N46), .Q(dout[15]) );
  TLATX1 dout_reg_14_ ( .G(n324), .D(N45), .Q(dout[14]) );
  TLATX1 dout_reg_13_ ( .G(n323), .D(N44), .Q(dout[13]) );
  TLATX1 dout_reg_12_ ( .G(n323), .D(N43), .Q(dout[12]) );
  TLATX1 dout_reg_11_ ( .G(n321), .D(N42), .Q(dout[11]) );
  TLATX1 dout_reg_10_ ( .G(N30), .D(N41), .Q(dout[10]) );
  TLATX1 dout_reg_9_ ( .G(n318), .D(N40), .Q(dout[9]) );
  TLATX1 dout_reg_8_ ( .G(n330), .D(N39), .Q(dout[8]) );
  TLATX1 dout_reg_7_ ( .G(n330), .D(N38), .Q(dout[7]) );
  TLATX1 dout_reg_6_ ( .G(n320), .D(N37), .Q(dout[6]) );
  TLATX1 dout_reg_5_ ( .G(n327), .D(N36), .Q(dout[5]) );
  TLATX1 dout_reg_4_ ( .G(n329), .D(N35), .Q(dout[4]) );
  TLATX1 dout_reg_3_ ( .G(n328), .D(N34), .Q(dout[3]) );
  TLATX1 dout_reg_2_ ( .G(n328), .D(N33), .Q(dout[2]) );
  TLATX1 dout_reg_1_ ( .G(n327), .D(N32), .Q(dout[1]) );
  TLATX1 dout_reg_0_ ( .G(n326), .D(N31), .Q(dout[0]) );
  TLATX1 dout_reg_255_ ( .G(n322), .D(N288), .Q(dout[255]) );
  TLATX1 dout_reg_254_ ( .G(n321), .D(N287), .Q(dout[254]) );
  TLATX1 dout_reg_253_ ( .G(n321), .D(N286), .Q(dout[253]) );
  TLATX1 dout_reg_252_ ( .G(n321), .D(N285), .Q(dout[252]) );
  TLATX1 dout_reg_251_ ( .G(n321), .D(N284), .Q(dout[251]) );
  TLATX1 dout_reg_250_ ( .G(n329), .D(N283), .Q(dout[250]) );
  TLATX1 dout_reg_249_ ( .G(n319), .D(N282), .Q(dout[249]) );
  TLATX1 dout_reg_248_ ( .G(n320), .D(N281), .Q(dout[248]) );
  TLATX1 dout_reg_247_ ( .G(n320), .D(N280), .Q(dout[247]) );
  TLATX1 dout_reg_246_ ( .G(n320), .D(N279), .Q(dout[246]) );
  TLATX1 dout_reg_245_ ( .G(n319), .D(N278), .Q(dout[245]) );
  TLATX1 dout_reg_244_ ( .G(n319), .D(N277), .Q(dout[244]) );
  TLATX1 dout_reg_243_ ( .G(n319), .D(N276), .Q(dout[243]) );
  TLATX1 dout_reg_242_ ( .G(n318), .D(N275), .Q(dout[242]) );
  TLATX1 dout_reg_241_ ( .G(n318), .D(N274), .Q(dout[241]) );
  TLATX1 dout_reg_240_ ( .G(n318), .D(N273), .Q(dout[240]) );
  TLATX1 dout_reg_127_ ( .G(N30), .D(N159), .Q(dout[127]) );
  TLATX1 dout_reg_95_ ( .G(N30), .D(N126), .Q(dout[95]) );
  TLATX1 dout_reg_63_ ( .G(n323), .D(N94), .Q(dout[63]) );
  TLATX1 dout_reg_126_ ( .G(n321), .D(N158), .Q(dout[126]) );
  TLATX1 dout_reg_94_ ( .G(n329), .D(N125), .Q(dout[94]) );
  TLATX1 dout_reg_62_ ( .G(n327), .D(N93), .Q(dout[62]) );
  TLATX1 dout_reg_125_ ( .G(n321), .D(N157), .Q(dout[125]) );
  TLATX1 dout_reg_93_ ( .G(n329), .D(N124), .Q(dout[93]) );
  TLATX1 dout_reg_61_ ( .G(n325), .D(N92), .Q(dout[61]) );
  TLATX1 dout_reg_124_ ( .G(n320), .D(N156), .Q(dout[124]) );
  TLATX1 dout_reg_92_ ( .G(n319), .D(N123), .Q(dout[92]) );
  TLATX1 dout_reg_60_ ( .G(n329), .D(N91), .Q(dout[60]) );
  TLATX1 dout_reg_123_ ( .G(n322), .D(N155), .Q(dout[123]) );
  TLATX1 dout_reg_91_ ( .G(n320), .D(N122), .Q(dout[91]) );
  TLATX1 dout_reg_59_ ( .G(n319), .D(N90), .Q(dout[59]) );
  TLATX1 dout_reg_122_ ( .G(N30), .D(N154), .Q(dout[122]) );
  TLATX1 dout_reg_90_ ( .G(N30), .D(N121), .Q(dout[90]) );
  TLATX1 dout_reg_58_ ( .G(N30), .D(N89), .Q(dout[58]) );
  TLATX1 dout_reg_121_ ( .G(N30), .D(N153), .Q(dout[121]) );
  TLATX1 dout_reg_89_ ( .G(N30), .D(N120), .Q(dout[89]) );
  TLATX1 dout_reg_57_ ( .G(n324), .D(N88), .Q(dout[57]) );
  TLATX1 dout_reg_120_ ( .G(n323), .D(N152), .Q(dout[120]) );
  TLATX1 dout_reg_88_ ( .G(n321), .D(N119), .Q(dout[88]) );
  TLATX1 dout_reg_56_ ( .G(n329), .D(N87), .Q(dout[56]) );
  TLATX1 dout_reg_119_ ( .G(n330), .D(N151), .Q(dout[119]) );
  TLATX1 dout_reg_87_ ( .G(n330), .D(N118), .Q(dout[87]) );
  TLATX1 dout_reg_55_ ( .G(n330), .D(N86), .Q(dout[55]) );
  TLATX1 dout_reg_118_ ( .G(n330), .D(N150), .Q(dout[118]) );
  TLATX1 dout_reg_86_ ( .G(n330), .D(N117), .Q(dout[86]) );
  TLATX1 dout_reg_54_ ( .G(n323), .D(N85), .Q(dout[54]) );
  TLATX1 dout_reg_117_ ( .G(n327), .D(N149), .Q(dout[117]) );
  TLATX1 dout_reg_85_ ( .G(n330), .D(N116), .Q(dout[85]) );
  TLATX1 dout_reg_53_ ( .G(n324), .D(N84), .Q(dout[53]) );
  TLATX1 dout_reg_116_ ( .G(n329), .D(N148), .Q(dout[116]) );
  TLATX1 dout_reg_84_ ( .G(n329), .D(N115), .Q(dout[84]) );
  TLATX1 dout_reg_52_ ( .G(n329), .D(N83), .Q(dout[52]) );
  TLATX1 dout_reg_115_ ( .G(n329), .D(N147), .Q(dout[115]) );
  TLATX1 dout_reg_83_ ( .G(n329), .D(N114), .Q(dout[83]) );
  TLATX1 dout_reg_51_ ( .G(n328), .D(N82), .Q(dout[51]) );
  TLATX1 dout_reg_114_ ( .G(n328), .D(N146), .Q(dout[114]) );
  TLATX1 dout_reg_82_ ( .G(n328), .D(N113), .Q(dout[82]) );
  TLATX1 dout_reg_50_ ( .G(n328), .D(N81), .Q(dout[50]) );
  TLATX1 dout_reg_113_ ( .G(n327), .D(N145), .Q(dout[113]) );
  TLATX1 dout_reg_81_ ( .G(n327), .D(N112), .Q(dout[81]) );
  TLATX1 dout_reg_49_ ( .G(n327), .D(N80), .Q(dout[49]) );
  TLATX1 dout_reg_112_ ( .G(n327), .D(N144), .Q(dout[112]) );
  TLATX1 dout_reg_80_ ( .G(n327), .D(N111), .Q(dout[80]) );
  TLATX1 dout_reg_48_ ( .G(N30), .D(N79), .Q(dout[48]) );
  TLATX1 dout_reg_175_ ( .G(n318), .D(N207), .Q(dout[175]) );
  TLATX1 dout_reg_174_ ( .G(n319), .D(N206), .Q(dout[174]) );
  TLATX1 dout_reg_173_ ( .G(n326), .D(N205), .Q(dout[173]) );
  TLATX1 dout_reg_172_ ( .G(n326), .D(N204), .Q(dout[172]) );
  TLATX1 dout_reg_171_ ( .G(n326), .D(N203), .Q(dout[171]) );
  TLATX1 dout_reg_170_ ( .G(n325), .D(N202), .Q(dout[170]) );
  TLATX1 dout_reg_169_ ( .G(n325), .D(N201), .Q(dout[169]) );
  TLATX1 dout_reg_168_ ( .G(n325), .D(N200), .Q(dout[168]) );
  TLATX1 dout_reg_167_ ( .G(n324), .D(N199), .Q(dout[167]) );
  TLATX1 dout_reg_166_ ( .G(n324), .D(N198), .Q(dout[166]) );
  TLATX1 dout_reg_165_ ( .G(n324), .D(N197), .Q(dout[165]) );
  TLATX1 dout_reg_164_ ( .G(n323), .D(N196), .Q(dout[164]) );
  TLATX1 dout_reg_163_ ( .G(n323), .D(N195), .Q(dout[163]) );
  TLATX1 dout_reg_162_ ( .G(n323), .D(N194), .Q(dout[162]) );
  TLATX1 dout_reg_161_ ( .G(n322), .D(N193), .Q(dout[161]) );
  TLATX1 dout_reg_160_ ( .G(n322), .D(N192), .Q(dout[160]) );
  TLATX1 dout_reg_239_ ( .G(n322), .D(N272), .Q(dout[239]) );
  TLATX1 dout_reg_207_ ( .G(n322), .D(N240), .Q(dout[207]) );
  TLATX1 dout_reg_238_ ( .G(n321), .D(N271), .Q(dout[238]) );
  TLATX1 dout_reg_206_ ( .G(n321), .D(N239), .Q(dout[206]) );
  TLATX1 dout_reg_237_ ( .G(n321), .D(N270), .Q(dout[237]) );
  TLATX1 dout_reg_205_ ( .G(n321), .D(N238), .Q(dout[205]) );
  TLATX1 dout_reg_236_ ( .G(n321), .D(N269), .Q(dout[236]) );
  TLATX1 dout_reg_204_ ( .G(n321), .D(N237), .Q(dout[204]) );
  TLATX1 dout_reg_235_ ( .G(n320), .D(N268), .Q(dout[235]) );
  TLATX1 dout_reg_203_ ( .G(n319), .D(N236), .Q(dout[203]) );
  TLATX1 dout_reg_234_ ( .G(n327), .D(N267), .Q(dout[234]) );
  TLATX1 dout_reg_202_ ( .G(n325), .D(N235), .Q(dout[202]) );
  TLATX1 dout_reg_233_ ( .G(n322), .D(N266), .Q(dout[233]) );
  TLATX1 dout_reg_201_ ( .G(n328), .D(N234), .Q(dout[201]) );
  TLATX1 dout_reg_232_ ( .G(n320), .D(N265), .Q(dout[232]) );
  TLATX1 dout_reg_200_ ( .G(n320), .D(N233), .Q(dout[200]) );
  TLATX1 dout_reg_231_ ( .G(n320), .D(N264), .Q(dout[231]) );
  TLATX1 dout_reg_199_ ( .G(n320), .D(N232), .Q(dout[199]) );
  TLATX1 dout_reg_230_ ( .G(n320), .D(N263), .Q(dout[230]) );
  TLATX1 dout_reg_198_ ( .G(n320), .D(N231), .Q(dout[198]) );
  TLATX1 dout_reg_229_ ( .G(n319), .D(N262), .Q(dout[229]) );
  TLATX1 dout_reg_197_ ( .G(n319), .D(N229), .Q(dout[197]) );
  TLATX1 dout_reg_228_ ( .G(n319), .D(N261), .Q(dout[228]) );
  TLATX1 dout_reg_196_ ( .G(n319), .D(N228), .Q(dout[196]) );
  TLATX1 dout_reg_227_ ( .G(n319), .D(N260), .Q(dout[227]) );
  TLATX1 dout_reg_195_ ( .G(n319), .D(N227), .Q(dout[195]) );
  TLATX1 dout_reg_226_ ( .G(n318), .D(N259), .Q(dout[226]) );
  TLATX1 dout_reg_194_ ( .G(n318), .D(N226), .Q(dout[194]) );
  TLATX1 dout_reg_225_ ( .G(n318), .D(N258), .Q(dout[225]) );
  TLATX1 dout_reg_193_ ( .G(n318), .D(N225), .Q(dout[193]) );
  TLATX1 dout_reg_224_ ( .G(n318), .D(N257), .Q(dout[224]) );
  TLATX1 dout_reg_192_ ( .G(n318), .D(N224), .Q(dout[192]) );
  TLATX1 dout_reg_191_ ( .G(n325), .D(N223), .Q(dout[191]) );
  TLATX1 dout_reg_159_ ( .G(n325), .D(N191), .Q(dout[159]) );
  TLATX1 dout_reg_190_ ( .G(n330), .D(N222), .Q(dout[190]) );
  TLATX1 dout_reg_158_ ( .G(n324), .D(N190), .Q(dout[158]) );
  TLATX1 dout_reg_189_ ( .G(n326), .D(N221), .Q(dout[189]) );
  TLATX1 dout_reg_157_ ( .G(n326), .D(N189), .Q(dout[157]) );
  TLATX1 dout_reg_188_ ( .G(n326), .D(N220), .Q(dout[188]) );
  TLATX1 dout_reg_156_ ( .G(n326), .D(N188), .Q(dout[156]) );
  TLATX1 dout_reg_187_ ( .G(n326), .D(N219), .Q(dout[187]) );
  TLATX1 dout_reg_155_ ( .G(n326), .D(N187), .Q(dout[155]) );
  TLATX1 dout_reg_186_ ( .G(n325), .D(N218), .Q(dout[186]) );
  TLATX1 dout_reg_154_ ( .G(n325), .D(N186), .Q(dout[154]) );
  TLATX1 dout_reg_185_ ( .G(n325), .D(N217), .Q(dout[185]) );
  TLATX1 dout_reg_153_ ( .G(n325), .D(N185), .Q(dout[153]) );
  TLATX1 dout_reg_184_ ( .G(n325), .D(N216), .Q(dout[184]) );
  TLATX1 dout_reg_152_ ( .G(n325), .D(N184), .Q(dout[152]) );
  TLATX1 dout_reg_183_ ( .G(n324), .D(N215), .Q(dout[183]) );
  TLATX1 dout_reg_151_ ( .G(n324), .D(N183), .Q(dout[151]) );
  TLATX1 dout_reg_182_ ( .G(n324), .D(N214), .Q(dout[182]) );
  TLATX1 dout_reg_150_ ( .G(n324), .D(N182), .Q(dout[150]) );
  TLATX1 dout_reg_181_ ( .G(n324), .D(N213), .Q(dout[181]) );
  TLATX1 dout_reg_149_ ( .G(n324), .D(N181), .Q(dout[149]) );
  TLATX1 dout_reg_180_ ( .G(n323), .D(N212), .Q(dout[180]) );
  TLATX1 dout_reg_148_ ( .G(n323), .D(N180), .Q(dout[148]) );
  TLATX1 dout_reg_179_ ( .G(n323), .D(N211), .Q(dout[179]) );
  TLATX1 dout_reg_147_ ( .G(n323), .D(N179), .Q(dout[147]) );
  TLATX1 dout_reg_178_ ( .G(n323), .D(N210), .Q(dout[178]) );
  TLATX1 dout_reg_146_ ( .G(n323), .D(N178), .Q(dout[146]) );
  TLATX1 dout_reg_177_ ( .G(n322), .D(N209), .Q(dout[177]) );
  TLATX1 dout_reg_145_ ( .G(n322), .D(N177), .Q(dout[145]) );
  TLATX1 dout_reg_176_ ( .G(n322), .D(N208), .Q(dout[176]) );
  TLATX1 dout_reg_144_ ( .G(n322), .D(N176), .Q(dout[144]) );
  TLATX1 dout_reg_223_ ( .G(n322), .D(N256), .Q(dout[223]) );
  TLATX1 dout_reg_222_ ( .G(n321), .D(N255), .Q(dout[222]) );
  TLATX1 dout_reg_221_ ( .G(n321), .D(N254), .Q(dout[221]) );
  TLATX1 dout_reg_220_ ( .G(n321), .D(N253), .Q(dout[220]) );
  TLATX1 dout_reg_219_ ( .G(n326), .D(N252), .Q(dout[219]) );
  TLATX1 dout_reg_218_ ( .G(N30), .D(N251), .Q(dout[218]) );
  TLATX1 dout_reg_217_ ( .G(N30), .D(N250), .Q(dout[217]) );
  TLATX1 dout_reg_216_ ( .G(n320), .D(N249), .Q(dout[216]) );
  TLATX1 dout_reg_215_ ( .G(n320), .D(N248), .Q(dout[215]) );
  TLATX1 dout_reg_214_ ( .G(n320), .D(N247), .Q(dout[214]) );
  TLATX1 dout_reg_213_ ( .G(n319), .D(N246), .Q(dout[213]) );
  TLATX1 dout_reg_212_ ( .G(n319), .D(N245), .Q(dout[212]) );
  TLATX1 dout_reg_211_ ( .G(n319), .D(N244), .Q(dout[211]) );
  TLATX1 dout_reg_210_ ( .G(n318), .D(N243), .Q(dout[210]) );
  TLATX1 dout_reg_209_ ( .G(n318), .D(N242), .Q(dout[209]) );
  TLATX1 dout_reg_208_ ( .G(n318), .D(N241), .Q(dout[208]) );
  DFFRHQX1 dout16_reg_reg_207_ ( .D(n991), .CK(clk), .RN(rstn), .Q(
        dout16_reg[207]) );
  DFFRHQX1 dout16_reg_reg_223_ ( .D(n975), .CK(clk), .RN(rstn), .Q(
        dout16_reg[223]) );
  DFFRHQX1 dout16_reg_reg_239_ ( .D(n959), .CK(clk), .RN(rstn), .Q(
        dout16_reg[239]) );
  DFFRHQX1 dout16_reg_reg_255_ ( .D(n943), .CK(clk), .RN(rstn), .Q(
        dout16_reg[255]) );
  DFFRHQX1 dout16_reg_reg_206_ ( .D(n992), .CK(clk), .RN(rstn), .Q(
        dout16_reg[206]) );
  DFFRHQX1 dout16_reg_reg_222_ ( .D(n976), .CK(clk), .RN(rstn), .Q(
        dout16_reg[222]) );
  DFFRHQX1 dout16_reg_reg_238_ ( .D(n960), .CK(clk), .RN(rstn), .Q(
        dout16_reg[238]) );
  DFFRHQX1 dout16_reg_reg_254_ ( .D(n944), .CK(clk), .RN(rstn), .Q(
        dout16_reg[254]) );
  DFFRHQX1 dout16_reg_reg_205_ ( .D(n993), .CK(clk), .RN(rstn), .Q(
        dout16_reg[205]) );
  DFFRHQX1 dout16_reg_reg_221_ ( .D(n977), .CK(clk), .RN(rstn), .Q(
        dout16_reg[221]) );
  DFFRHQX1 dout16_reg_reg_237_ ( .D(n961), .CK(clk), .RN(rstn), .Q(
        dout16_reg[237]) );
  DFFRHQX1 dout16_reg_reg_253_ ( .D(n945), .CK(clk), .RN(rstn), .Q(
        dout16_reg[253]) );
  DFFRHQX1 dout16_reg_reg_204_ ( .D(n994), .CK(clk), .RN(rstn), .Q(
        dout16_reg[204]) );
  DFFRHQX1 dout16_reg_reg_220_ ( .D(n978), .CK(clk), .RN(rstn), .Q(
        dout16_reg[220]) );
  DFFRHQX1 dout16_reg_reg_236_ ( .D(n962), .CK(clk), .RN(rstn), .Q(
        dout16_reg[236]) );
  DFFRHQX1 dout16_reg_reg_252_ ( .D(n946), .CK(clk), .RN(rstn), .Q(
        dout16_reg[252]) );
  DFFRHQX1 dout16_reg_reg_203_ ( .D(n995), .CK(clk), .RN(rstn), .Q(
        dout16_reg[203]) );
  DFFRHQX1 dout16_reg_reg_219_ ( .D(n979), .CK(clk), .RN(rstn), .Q(
        dout16_reg[219]) );
  DFFRHQX1 dout16_reg_reg_235_ ( .D(n963), .CK(clk), .RN(rstn), .Q(
        dout16_reg[235]) );
  DFFRHQX1 dout16_reg_reg_251_ ( .D(n947), .CK(clk), .RN(rstn), .Q(
        dout16_reg[251]) );
  DFFRHQX1 dout16_reg_reg_202_ ( .D(n996), .CK(clk), .RN(rstn), .Q(
        dout16_reg[202]) );
  DFFRHQX1 dout16_reg_reg_218_ ( .D(n980), .CK(clk), .RN(rstn), .Q(
        dout16_reg[218]) );
  DFFRHQX1 dout16_reg_reg_234_ ( .D(n964), .CK(clk), .RN(rstn), .Q(
        dout16_reg[234]) );
  DFFRHQX1 dout16_reg_reg_250_ ( .D(n948), .CK(clk), .RN(rstn), .Q(
        dout16_reg[250]) );
  DFFRHQX1 dout16_reg_reg_201_ ( .D(n997), .CK(clk), .RN(rstn), .Q(
        dout16_reg[201]) );
  DFFRHQX1 dout16_reg_reg_217_ ( .D(n981), .CK(clk), .RN(rstn), .Q(
        dout16_reg[217]) );
  DFFRHQX1 dout16_reg_reg_233_ ( .D(n965), .CK(clk), .RN(rstn), .Q(
        dout16_reg[233]) );
  DFFRHQX1 dout16_reg_reg_249_ ( .D(n949), .CK(clk), .RN(rstn), .Q(
        dout16_reg[249]) );
  DFFRHQX1 dout16_reg_reg_200_ ( .D(n998), .CK(clk), .RN(rstn), .Q(
        dout16_reg[200]) );
  DFFRHQX1 dout16_reg_reg_216_ ( .D(n982), .CK(clk), .RN(rstn), .Q(
        dout16_reg[216]) );
  DFFRHQX1 dout16_reg_reg_232_ ( .D(n966), .CK(clk), .RN(rstn), .Q(
        dout16_reg[232]) );
  DFFRHQX1 dout16_reg_reg_248_ ( .D(n950), .CK(clk), .RN(rstn), .Q(
        dout16_reg[248]) );
  DFFRHQX1 dout16_reg_reg_199_ ( .D(n999), .CK(clk), .RN(rstn), .Q(
        dout16_reg[199]) );
  DFFRHQX1 dout16_reg_reg_215_ ( .D(n983), .CK(clk), .RN(rstn), .Q(
        dout16_reg[215]) );
  DFFRHQX1 dout16_reg_reg_231_ ( .D(n967), .CK(clk), .RN(rstn), .Q(
        dout16_reg[231]) );
  DFFRHQX1 dout16_reg_reg_247_ ( .D(n951), .CK(clk), .RN(rstn), .Q(
        dout16_reg[247]) );
  DFFRHQX1 dout16_reg_reg_198_ ( .D(n1000), .CK(clk), .RN(rstn), .Q(
        dout16_reg[198]) );
  DFFRHQX1 dout16_reg_reg_214_ ( .D(n984), .CK(clk), .RN(rstn), .Q(
        dout16_reg[214]) );
  DFFRHQX1 dout16_reg_reg_230_ ( .D(n968), .CK(clk), .RN(rstn), .Q(
        dout16_reg[230]) );
  DFFRHQX1 dout16_reg_reg_246_ ( .D(n952), .CK(clk), .RN(rstn), .Q(
        dout16_reg[246]) );
  DFFRHQX1 dout16_reg_reg_197_ ( .D(n1001), .CK(clk), .RN(rstn), .Q(
        dout16_reg[197]) );
  DFFRHQX1 dout16_reg_reg_213_ ( .D(n985), .CK(clk), .RN(rstn), .Q(
        dout16_reg[213]) );
  DFFRHQX1 dout16_reg_reg_229_ ( .D(n969), .CK(clk), .RN(rstn), .Q(
        dout16_reg[229]) );
  DFFRHQX1 dout16_reg_reg_245_ ( .D(n953), .CK(clk), .RN(rstn), .Q(
        dout16_reg[245]) );
  DFFRHQX1 dout16_reg_reg_196_ ( .D(n1002), .CK(clk), .RN(rstn), .Q(
        dout16_reg[196]) );
  DFFRHQX1 dout16_reg_reg_212_ ( .D(n986), .CK(clk), .RN(rstn), .Q(
        dout16_reg[212]) );
  DFFRHQX1 dout16_reg_reg_228_ ( .D(n970), .CK(clk), .RN(rstn), .Q(
        dout16_reg[228]) );
  DFFRHQX1 dout16_reg_reg_244_ ( .D(n954), .CK(clk), .RN(rstn), .Q(
        dout16_reg[244]) );
  DFFRHQX1 dout16_reg_reg_195_ ( .D(n1003), .CK(clk), .RN(rstn), .Q(
        dout16_reg[195]) );
  DFFRHQX1 dout16_reg_reg_211_ ( .D(n987), .CK(clk), .RN(rstn), .Q(
        dout16_reg[211]) );
  DFFRHQX1 dout16_reg_reg_227_ ( .D(n971), .CK(clk), .RN(rstn), .Q(
        dout16_reg[227]) );
  DFFRHQX1 dout16_reg_reg_243_ ( .D(n955), .CK(clk), .RN(rstn), .Q(
        dout16_reg[243]) );
  DFFRHQX1 dout16_reg_reg_194_ ( .D(n1004), .CK(clk), .RN(rstn), .Q(
        dout16_reg[194]) );
  DFFRHQX1 dout16_reg_reg_210_ ( .D(n988), .CK(clk), .RN(rstn), .Q(
        dout16_reg[210]) );
  DFFRHQX1 dout16_reg_reg_226_ ( .D(n972), .CK(clk), .RN(rstn), .Q(
        dout16_reg[226]) );
  DFFRHQX1 dout16_reg_reg_242_ ( .D(n956), .CK(clk), .RN(rstn), .Q(
        dout16_reg[242]) );
  DFFRHQX1 dout16_reg_reg_193_ ( .D(n1005), .CK(clk), .RN(rstn), .Q(
        dout16_reg[193]) );
  DFFRHQX1 dout16_reg_reg_209_ ( .D(n989), .CK(clk), .RN(rstn), .Q(
        dout16_reg[209]) );
  DFFRHQX1 dout16_reg_reg_225_ ( .D(n973), .CK(clk), .RN(rstn), .Q(
        dout16_reg[225]) );
  DFFRHQX1 dout16_reg_reg_241_ ( .D(n957), .CK(clk), .RN(rstn), .Q(
        dout16_reg[241]) );
  DFFRHQX1 dout16_reg_reg_192_ ( .D(n1006), .CK(clk), .RN(rstn), .Q(
        dout16_reg[192]) );
  DFFRHQX1 dout16_reg_reg_208_ ( .D(n990), .CK(clk), .RN(rstn), .Q(
        dout16_reg[208]) );
  DFFRHQX1 dout16_reg_reg_224_ ( .D(n974), .CK(clk), .RN(rstn), .Q(
        dout16_reg[224]) );
  DFFRHQX1 dout16_reg_reg_240_ ( .D(n958), .CK(clk), .RN(rstn), .Q(
        dout16_reg[240]) );
  DFFRHQX1 dout8_reg_reg_79_ ( .D(n863), .CK(clk), .RN(rstn), .Q(dout8_reg[79]) );
  DFFRHQX1 dout8_reg_reg_95_ ( .D(n847), .CK(clk), .RN(rstn), .Q(dout8_reg[95]) );
  DFFRHQX1 dout8_reg_reg_111_ ( .D(n831), .CK(clk), .RN(rstn), .Q(
        dout8_reg[111]) );
  DFFRHQX1 dout8_reg_reg_127_ ( .D(n815), .CK(clk), .RN(rstn), .Q(
        dout8_reg[127]) );
  DFFRHQX1 dout8_reg_reg_78_ ( .D(n864), .CK(clk), .RN(rstn), .Q(dout8_reg[78]) );
  DFFRHQX1 dout8_reg_reg_94_ ( .D(n848), .CK(clk), .RN(rstn), .Q(dout8_reg[94]) );
  DFFRHQX1 dout8_reg_reg_110_ ( .D(n832), .CK(clk), .RN(rstn), .Q(
        dout8_reg[110]) );
  DFFRHQX1 dout8_reg_reg_126_ ( .D(n816), .CK(clk), .RN(rstn), .Q(
        dout8_reg[126]) );
  DFFRHQX1 dout8_reg_reg_77_ ( .D(n865), .CK(clk), .RN(rstn), .Q(dout8_reg[77]) );
  DFFRHQX1 dout8_reg_reg_93_ ( .D(n849), .CK(clk), .RN(rstn), .Q(dout8_reg[93]) );
  DFFRHQX1 dout8_reg_reg_109_ ( .D(n833), .CK(clk), .RN(rstn), .Q(
        dout8_reg[109]) );
  DFFRHQX1 dout8_reg_reg_125_ ( .D(n817), .CK(clk), .RN(rstn), .Q(
        dout8_reg[125]) );
  DFFRHQX1 dout8_reg_reg_76_ ( .D(n866), .CK(clk), .RN(rstn), .Q(dout8_reg[76]) );
  DFFRHQX1 dout8_reg_reg_92_ ( .D(n850), .CK(clk), .RN(rstn), .Q(dout8_reg[92]) );
  DFFRHQX1 dout8_reg_reg_108_ ( .D(n834), .CK(clk), .RN(rstn), .Q(
        dout8_reg[108]) );
  DFFRHQX1 dout8_reg_reg_124_ ( .D(n818), .CK(clk), .RN(rstn), .Q(
        dout8_reg[124]) );
  DFFRHQX1 dout8_reg_reg_75_ ( .D(n867), .CK(clk), .RN(rstn), .Q(dout8_reg[75]) );
  DFFRHQX1 dout8_reg_reg_91_ ( .D(n851), .CK(clk), .RN(rstn), .Q(dout8_reg[91]) );
  DFFRHQX1 dout8_reg_reg_107_ ( .D(n835), .CK(clk), .RN(rstn), .Q(
        dout8_reg[107]) );
  DFFRHQX1 dout8_reg_reg_123_ ( .D(n819), .CK(clk), .RN(rstn), .Q(
        dout8_reg[123]) );
  DFFRHQX1 dout8_reg_reg_74_ ( .D(n868), .CK(clk), .RN(rstn), .Q(dout8_reg[74]) );
  DFFRHQX1 dout8_reg_reg_90_ ( .D(n852), .CK(clk), .RN(rstn), .Q(dout8_reg[90]) );
  DFFRHQX1 dout8_reg_reg_106_ ( .D(n836), .CK(clk), .RN(rstn), .Q(
        dout8_reg[106]) );
  DFFRHQX1 dout8_reg_reg_122_ ( .D(n820), .CK(clk), .RN(rstn), .Q(
        dout8_reg[122]) );
  DFFRHQX1 dout8_reg_reg_73_ ( .D(n869), .CK(clk), .RN(rstn), .Q(dout8_reg[73]) );
  DFFRHQX1 dout8_reg_reg_89_ ( .D(n853), .CK(clk), .RN(rstn), .Q(dout8_reg[89]) );
  DFFRHQX1 dout8_reg_reg_105_ ( .D(n837), .CK(clk), .RN(rstn), .Q(
        dout8_reg[105]) );
  DFFRHQX1 dout8_reg_reg_121_ ( .D(n821), .CK(clk), .RN(rstn), .Q(
        dout8_reg[121]) );
  DFFRHQX1 dout8_reg_reg_72_ ( .D(n870), .CK(clk), .RN(rstn), .Q(dout8_reg[72]) );
  DFFRHQX1 dout8_reg_reg_88_ ( .D(n854), .CK(clk), .RN(rstn), .Q(dout8_reg[88]) );
  DFFRHQX1 dout8_reg_reg_104_ ( .D(n838), .CK(clk), .RN(rstn), .Q(
        dout8_reg[104]) );
  DFFRHQX1 dout8_reg_reg_120_ ( .D(n822), .CK(clk), .RN(rstn), .Q(
        dout8_reg[120]) );
  DFFRHQX1 dout8_reg_reg_71_ ( .D(n871), .CK(clk), .RN(rstn), .Q(dout8_reg[71]) );
  DFFRHQX1 dout8_reg_reg_87_ ( .D(n855), .CK(clk), .RN(rstn), .Q(dout8_reg[87]) );
  DFFRHQX1 dout8_reg_reg_103_ ( .D(n839), .CK(clk), .RN(rstn), .Q(
        dout8_reg[103]) );
  DFFRHQX1 dout8_reg_reg_119_ ( .D(n823), .CK(clk), .RN(rstn), .Q(
        dout8_reg[119]) );
  DFFRHQX1 dout8_reg_reg_70_ ( .D(n872), .CK(clk), .RN(rstn), .Q(dout8_reg[70]) );
  DFFRHQX1 dout8_reg_reg_86_ ( .D(n856), .CK(clk), .RN(rstn), .Q(dout8_reg[86]) );
  DFFRHQX1 dout8_reg_reg_102_ ( .D(n840), .CK(clk), .RN(rstn), .Q(
        dout8_reg[102]) );
  DFFRHQX1 dout8_reg_reg_118_ ( .D(n824), .CK(clk), .RN(rstn), .Q(
        dout8_reg[118]) );
  DFFRHQX1 dout8_reg_reg_69_ ( .D(n873), .CK(clk), .RN(rstn), .Q(dout8_reg[69]) );
  DFFRHQX1 dout8_reg_reg_85_ ( .D(n857), .CK(clk), .RN(rstn), .Q(dout8_reg[85]) );
  DFFRHQX1 dout8_reg_reg_101_ ( .D(n841), .CK(clk), .RN(rstn), .Q(
        dout8_reg[101]) );
  DFFRHQX1 dout8_reg_reg_117_ ( .D(n825), .CK(clk), .RN(rstn), .Q(
        dout8_reg[117]) );
  DFFRHQX1 dout8_reg_reg_68_ ( .D(n874), .CK(clk), .RN(rstn), .Q(dout8_reg[68]) );
  DFFRHQX1 dout8_reg_reg_84_ ( .D(n858), .CK(clk), .RN(rstn), .Q(dout8_reg[84]) );
  DFFRHQX1 dout8_reg_reg_100_ ( .D(n842), .CK(clk), .RN(rstn), .Q(
        dout8_reg[100]) );
  DFFRHQX1 dout8_reg_reg_116_ ( .D(n826), .CK(clk), .RN(rstn), .Q(
        dout8_reg[116]) );
  DFFRHQX1 dout8_reg_reg_67_ ( .D(n875), .CK(clk), .RN(rstn), .Q(dout8_reg[67]) );
  DFFRHQX1 dout8_reg_reg_83_ ( .D(n859), .CK(clk), .RN(rstn), .Q(dout8_reg[83]) );
  DFFRHQX1 dout8_reg_reg_99_ ( .D(n843), .CK(clk), .RN(rstn), .Q(dout8_reg[99]) );
  DFFRHQX1 dout8_reg_reg_115_ ( .D(n827), .CK(clk), .RN(rstn), .Q(
        dout8_reg[115]) );
  DFFRHQX1 dout8_reg_reg_66_ ( .D(n876), .CK(clk), .RN(rstn), .Q(dout8_reg[66]) );
  DFFRHQX1 dout8_reg_reg_82_ ( .D(n860), .CK(clk), .RN(rstn), .Q(dout8_reg[82]) );
  DFFRHQX1 dout8_reg_reg_98_ ( .D(n844), .CK(clk), .RN(rstn), .Q(dout8_reg[98]) );
  DFFRHQX1 dout8_reg_reg_114_ ( .D(n828), .CK(clk), .RN(rstn), .Q(
        dout8_reg[114]) );
  DFFRHQX1 dout8_reg_reg_65_ ( .D(n877), .CK(clk), .RN(rstn), .Q(dout8_reg[65]) );
  DFFRHQX1 dout8_reg_reg_81_ ( .D(n861), .CK(clk), .RN(rstn), .Q(dout8_reg[81]) );
  DFFRHQX1 dout8_reg_reg_97_ ( .D(n845), .CK(clk), .RN(rstn), .Q(dout8_reg[97]) );
  DFFRHQX1 dout8_reg_reg_113_ ( .D(n829), .CK(clk), .RN(rstn), .Q(
        dout8_reg[113]) );
  DFFRHQX1 dout8_reg_reg_64_ ( .D(n878), .CK(clk), .RN(rstn), .Q(dout8_reg[64]) );
  DFFRHQX1 dout8_reg_reg_80_ ( .D(n862), .CK(clk), .RN(rstn), .Q(dout8_reg[80]) );
  DFFRHQX1 dout8_reg_reg_96_ ( .D(n846), .CK(clk), .RN(rstn), .Q(dout8_reg[96]) );
  DFFRHQX1 dout8_reg_reg_112_ ( .D(n830), .CK(clk), .RN(rstn), .Q(
        dout8_reg[112]) );
  DFFRHQX1 dout4_reg_reg_15_ ( .D(n799), .CK(clk), .RN(rstn), .Q(dout4_reg[15]) );
  DFFRHQX1 dout4_reg_reg_31_ ( .D(n783), .CK(clk), .RN(rstn), .Q(dout4_reg[31]) );
  DFFRHQX1 dout4_reg_reg_47_ ( .D(n767), .CK(clk), .RN(rstn), .Q(dout4_reg[47]) );
  DFFRHQX1 dout4_reg_reg_63_ ( .D(n751), .CK(clk), .RN(rstn), .Q(dout4_reg[63]) );
  DFFRHQX1 dout4_reg_reg_14_ ( .D(n800), .CK(clk), .RN(rstn), .Q(dout4_reg[14]) );
  DFFRHQX1 dout4_reg_reg_30_ ( .D(n784), .CK(clk), .RN(rstn), .Q(dout4_reg[30]) );
  DFFRHQX1 dout4_reg_reg_46_ ( .D(n768), .CK(clk), .RN(rstn), .Q(dout4_reg[46]) );
  DFFRHQX1 dout4_reg_reg_62_ ( .D(n752), .CK(clk), .RN(rstn), .Q(dout4_reg[62]) );
  DFFRHQX1 dout4_reg_reg_13_ ( .D(n801), .CK(clk), .RN(rstn), .Q(dout4_reg[13]) );
  DFFRHQX1 dout4_reg_reg_29_ ( .D(n785), .CK(clk), .RN(rstn), .Q(dout4_reg[29]) );
  DFFRHQX1 dout4_reg_reg_45_ ( .D(n769), .CK(clk), .RN(rstn), .Q(dout4_reg[45]) );
  DFFRHQX1 dout4_reg_reg_61_ ( .D(n753), .CK(clk), .RN(rstn), .Q(dout4_reg[61]) );
  DFFRHQX1 dout4_reg_reg_12_ ( .D(n802), .CK(clk), .RN(rstn), .Q(dout4_reg[12]) );
  DFFRHQX1 dout4_reg_reg_28_ ( .D(n786), .CK(clk), .RN(rstn), .Q(dout4_reg[28]) );
  DFFRHQX1 dout4_reg_reg_44_ ( .D(n770), .CK(clk), .RN(rstn), .Q(dout4_reg[44]) );
  DFFRHQX1 dout4_reg_reg_60_ ( .D(n754), .CK(clk), .RN(rstn), .Q(dout4_reg[60]) );
  DFFRHQX1 dout4_reg_reg_11_ ( .D(n803), .CK(clk), .RN(rstn), .Q(dout4_reg[11]) );
  DFFRHQX1 dout4_reg_reg_27_ ( .D(n787), .CK(clk), .RN(rstn), .Q(dout4_reg[27]) );
  DFFRHQX1 dout4_reg_reg_43_ ( .D(n771), .CK(clk), .RN(rstn), .Q(dout4_reg[43]) );
  DFFRHQX1 dout4_reg_reg_59_ ( .D(n755), .CK(clk), .RN(rstn), .Q(dout4_reg[59]) );
  DFFRHQX1 dout4_reg_reg_10_ ( .D(n804), .CK(clk), .RN(rstn), .Q(dout4_reg[10]) );
  DFFRHQX1 dout4_reg_reg_26_ ( .D(n788), .CK(clk), .RN(rstn), .Q(dout4_reg[26]) );
  DFFRHQX1 dout4_reg_reg_42_ ( .D(n772), .CK(clk), .RN(rstn), .Q(dout4_reg[42]) );
  DFFRHQX1 dout4_reg_reg_58_ ( .D(n756), .CK(clk), .RN(rstn), .Q(dout4_reg[58]) );
  DFFRHQX1 dout4_reg_reg_9_ ( .D(n805), .CK(clk), .RN(rstn), .Q(dout4_reg[9])
         );
  DFFRHQX1 dout4_reg_reg_25_ ( .D(n789), .CK(clk), .RN(rstn), .Q(dout4_reg[25]) );
  DFFRHQX1 dout4_reg_reg_41_ ( .D(n773), .CK(clk), .RN(rstn), .Q(dout4_reg[41]) );
  DFFRHQX1 dout4_reg_reg_57_ ( .D(n757), .CK(clk), .RN(rstn), .Q(dout4_reg[57]) );
  DFFRHQX1 dout4_reg_reg_8_ ( .D(n806), .CK(clk), .RN(rstn), .Q(dout4_reg[8])
         );
  DFFRHQX1 dout4_reg_reg_24_ ( .D(n790), .CK(clk), .RN(rstn), .Q(dout4_reg[24]) );
  DFFRHQX1 dout4_reg_reg_40_ ( .D(n774), .CK(clk), .RN(rstn), .Q(dout4_reg[40]) );
  DFFRHQX1 dout4_reg_reg_56_ ( .D(n758), .CK(clk), .RN(rstn), .Q(dout4_reg[56]) );
  DFFRHQX1 dout4_reg_reg_7_ ( .D(n807), .CK(clk), .RN(rstn), .Q(dout4_reg[7])
         );
  DFFRHQX1 dout4_reg_reg_23_ ( .D(n791), .CK(clk), .RN(rstn), .Q(dout4_reg[23]) );
  DFFRHQX1 dout4_reg_reg_39_ ( .D(n775), .CK(clk), .RN(rstn), .Q(dout4_reg[39]) );
  DFFRHQX1 dout4_reg_reg_55_ ( .D(n759), .CK(clk), .RN(rstn), .Q(dout4_reg[55]) );
  DFFRHQX1 dout4_reg_reg_6_ ( .D(n808), .CK(clk), .RN(rstn), .Q(dout4_reg[6])
         );
  DFFRHQX1 dout4_reg_reg_22_ ( .D(n792), .CK(clk), .RN(rstn), .Q(dout4_reg[22]) );
  DFFRHQX1 dout4_reg_reg_38_ ( .D(n776), .CK(clk), .RN(rstn), .Q(dout4_reg[38]) );
  DFFRHQX1 dout4_reg_reg_54_ ( .D(n760), .CK(clk), .RN(rstn), .Q(dout4_reg[54]) );
  DFFRHQX1 dout4_reg_reg_5_ ( .D(n809), .CK(clk), .RN(rstn), .Q(dout4_reg[5])
         );
  DFFRHQX1 dout4_reg_reg_21_ ( .D(n793), .CK(clk), .RN(rstn), .Q(dout4_reg[21]) );
  DFFRHQX1 dout4_reg_reg_37_ ( .D(n777), .CK(clk), .RN(rstn), .Q(dout4_reg[37]) );
  DFFRHQX1 dout4_reg_reg_53_ ( .D(n761), .CK(clk), .RN(rstn), .Q(dout4_reg[53]) );
  DFFRHQX1 dout4_reg_reg_4_ ( .D(n810), .CK(clk), .RN(rstn), .Q(dout4_reg[4])
         );
  DFFRHQX1 dout4_reg_reg_20_ ( .D(n794), .CK(clk), .RN(rstn), .Q(dout4_reg[20]) );
  DFFRHQX1 dout4_reg_reg_36_ ( .D(n778), .CK(clk), .RN(rstn), .Q(dout4_reg[36]) );
  DFFRHQX1 dout4_reg_reg_52_ ( .D(n762), .CK(clk), .RN(rstn), .Q(dout4_reg[52]) );
  DFFRHQX1 dout4_reg_reg_3_ ( .D(n811), .CK(clk), .RN(rstn), .Q(dout4_reg[3])
         );
  DFFRHQX1 dout4_reg_reg_19_ ( .D(n795), .CK(clk), .RN(rstn), .Q(dout4_reg[19]) );
  DFFRHQX1 dout4_reg_reg_35_ ( .D(n779), .CK(clk), .RN(rstn), .Q(dout4_reg[35]) );
  DFFRHQX1 dout4_reg_reg_51_ ( .D(n763), .CK(clk), .RN(rstn), .Q(dout4_reg[51]) );
  DFFRHQX1 dout4_reg_reg_2_ ( .D(n812), .CK(clk), .RN(rstn), .Q(dout4_reg[2])
         );
  DFFRHQX1 dout4_reg_reg_18_ ( .D(n796), .CK(clk), .RN(rstn), .Q(dout4_reg[18]) );
  DFFRHQX1 dout4_reg_reg_34_ ( .D(n780), .CK(clk), .RN(rstn), .Q(dout4_reg[34]) );
  DFFRHQX1 dout4_reg_reg_50_ ( .D(n764), .CK(clk), .RN(rstn), .Q(dout4_reg[50]) );
  DFFRHQX1 dout4_reg_reg_1_ ( .D(n813), .CK(clk), .RN(rstn), .Q(dout4_reg[1])
         );
  DFFRHQX1 dout4_reg_reg_17_ ( .D(n797), .CK(clk), .RN(rstn), .Q(dout4_reg[17]) );
  DFFRHQX1 dout4_reg_reg_33_ ( .D(n781), .CK(clk), .RN(rstn), .Q(dout4_reg[33]) );
  DFFRHQX1 dout4_reg_reg_49_ ( .D(n765), .CK(clk), .RN(rstn), .Q(dout4_reg[49]) );
  DFFRHQX1 dout4_reg_reg_0_ ( .D(n814), .CK(clk), .RN(rstn), .Q(dout4_reg[0])
         );
  DFFRHQX1 dout4_reg_reg_16_ ( .D(n798), .CK(clk), .RN(rstn), .Q(dout4_reg[16]) );
  DFFRHQX1 dout4_reg_reg_32_ ( .D(n782), .CK(clk), .RN(rstn), .Q(dout4_reg[32]) );
  DFFRHQX1 dout4_reg_reg_48_ ( .D(n766), .CK(clk), .RN(rstn), .Q(dout4_reg[48]) );
  DFFRHQX1 count_reg_4_ ( .D(N1118), .CK(clk), .RN(rstn), .Q(count[4]) );
  DFFRHQX1 dout16_reg_reg_15_ ( .D(n1183), .CK(clk), .RN(rstn), .Q(
        dout16_reg[15]) );
  DFFRHQX1 dout16_reg_reg_31_ ( .D(n1167), .CK(clk), .RN(rstn), .Q(
        dout16_reg[31]) );
  DFFRHQX1 dout16_reg_reg_47_ ( .D(n1151), .CK(clk), .RN(rstn), .Q(
        dout16_reg[47]) );
  DFFRHQX1 dout16_reg_reg_63_ ( .D(n1135), .CK(clk), .RN(rstn), .Q(
        dout16_reg[63]) );
  DFFRHQX1 dout16_reg_reg_79_ ( .D(n1119), .CK(clk), .RN(rstn), .Q(
        dout16_reg[79]) );
  DFFRHQX1 dout16_reg_reg_95_ ( .D(n1103), .CK(clk), .RN(rstn), .Q(
        dout16_reg[95]) );
  DFFRHQX1 dout16_reg_reg_111_ ( .D(n1087), .CK(clk), .RN(rstn), .Q(
        dout16_reg[111]) );
  DFFRHQX1 dout16_reg_reg_127_ ( .D(n1071), .CK(clk), .RN(rstn), .Q(
        dout16_reg[127]) );
  DFFRHQX1 dout16_reg_reg_143_ ( .D(n1055), .CK(clk), .RN(rstn), .Q(
        dout16_reg[143]) );
  DFFRHQX1 dout16_reg_reg_159_ ( .D(n1039), .CK(clk), .RN(rstn), .Q(
        dout16_reg[159]) );
  DFFRHQX1 dout16_reg_reg_175_ ( .D(n1023), .CK(clk), .RN(rstn), .Q(
        dout16_reg[175]) );
  DFFRHQX1 dout16_reg_reg_191_ ( .D(n1007), .CK(clk), .RN(rstn), .Q(
        dout16_reg[191]) );
  DFFRHQX1 dout16_reg_reg_14_ ( .D(n1184), .CK(clk), .RN(rstn), .Q(
        dout16_reg[14]) );
  DFFRHQX1 dout16_reg_reg_30_ ( .D(n1168), .CK(clk), .RN(rstn), .Q(
        dout16_reg[30]) );
  DFFRHQX1 dout16_reg_reg_46_ ( .D(n1152), .CK(clk), .RN(rstn), .Q(
        dout16_reg[46]) );
  DFFRHQX1 dout16_reg_reg_62_ ( .D(n1136), .CK(clk), .RN(rstn), .Q(
        dout16_reg[62]) );
  DFFRHQX1 dout16_reg_reg_78_ ( .D(n1120), .CK(clk), .RN(rstn), .Q(
        dout16_reg[78]) );
  DFFRHQX1 dout16_reg_reg_94_ ( .D(n1104), .CK(clk), .RN(rstn), .Q(
        dout16_reg[94]) );
  DFFRHQX1 dout16_reg_reg_110_ ( .D(n1088), .CK(clk), .RN(rstn), .Q(
        dout16_reg[110]) );
  DFFRHQX1 dout16_reg_reg_126_ ( .D(n1072), .CK(clk), .RN(rstn), .Q(
        dout16_reg[126]) );
  DFFRHQX1 dout16_reg_reg_142_ ( .D(n1056), .CK(clk), .RN(rstn), .Q(
        dout16_reg[142]) );
  DFFRHQX1 dout16_reg_reg_158_ ( .D(n1040), .CK(clk), .RN(rstn), .Q(
        dout16_reg[158]) );
  DFFRHQX1 dout16_reg_reg_174_ ( .D(n1024), .CK(clk), .RN(rstn), .Q(
        dout16_reg[174]) );
  DFFRHQX1 dout16_reg_reg_190_ ( .D(n1008), .CK(clk), .RN(rstn), .Q(
        dout16_reg[190]) );
  DFFRHQX1 dout16_reg_reg_13_ ( .D(n1185), .CK(clk), .RN(rstn), .Q(
        dout16_reg[13]) );
  DFFRHQX1 dout16_reg_reg_29_ ( .D(n1169), .CK(clk), .RN(rstn), .Q(
        dout16_reg[29]) );
  DFFRHQX1 dout16_reg_reg_45_ ( .D(n1153), .CK(clk), .RN(rstn), .Q(
        dout16_reg[45]) );
  DFFRHQX1 dout16_reg_reg_61_ ( .D(n1137), .CK(clk), .RN(rstn), .Q(
        dout16_reg[61]) );
  DFFRHQX1 dout16_reg_reg_77_ ( .D(n1121), .CK(clk), .RN(rstn), .Q(
        dout16_reg[77]) );
  DFFRHQX1 dout16_reg_reg_93_ ( .D(n1105), .CK(clk), .RN(rstn), .Q(
        dout16_reg[93]) );
  DFFRHQX1 dout16_reg_reg_109_ ( .D(n1089), .CK(clk), .RN(rstn), .Q(
        dout16_reg[109]) );
  DFFRHQX1 dout16_reg_reg_125_ ( .D(n1073), .CK(clk), .RN(rstn), .Q(
        dout16_reg[125]) );
  DFFRHQX1 dout16_reg_reg_141_ ( .D(n1057), .CK(clk), .RN(rstn), .Q(
        dout16_reg[141]) );
  DFFRHQX1 dout16_reg_reg_157_ ( .D(n1041), .CK(clk), .RN(rstn), .Q(
        dout16_reg[157]) );
  DFFRHQX1 dout16_reg_reg_173_ ( .D(n1025), .CK(clk), .RN(rstn), .Q(
        dout16_reg[173]) );
  DFFRHQX1 dout16_reg_reg_189_ ( .D(n1009), .CK(clk), .RN(rstn), .Q(
        dout16_reg[189]) );
  DFFRHQX1 dout16_reg_reg_12_ ( .D(n1186), .CK(clk), .RN(rstn), .Q(
        dout16_reg[12]) );
  DFFRHQX1 dout16_reg_reg_28_ ( .D(n1170), .CK(clk), .RN(rstn), .Q(
        dout16_reg[28]) );
  DFFRHQX1 dout16_reg_reg_44_ ( .D(n1154), .CK(clk), .RN(rstn), .Q(
        dout16_reg[44]) );
  DFFRHQX1 dout16_reg_reg_60_ ( .D(n1138), .CK(clk), .RN(rstn), .Q(
        dout16_reg[60]) );
  DFFRHQX1 dout16_reg_reg_76_ ( .D(n1122), .CK(clk), .RN(rstn), .Q(
        dout16_reg[76]) );
  DFFRHQX1 dout16_reg_reg_92_ ( .D(n1106), .CK(clk), .RN(rstn), .Q(
        dout16_reg[92]) );
  DFFRHQX1 dout16_reg_reg_108_ ( .D(n1090), .CK(clk), .RN(rstn), .Q(
        dout16_reg[108]) );
  DFFRHQX1 dout16_reg_reg_124_ ( .D(n1074), .CK(clk), .RN(rstn), .Q(
        dout16_reg[124]) );
  DFFRHQX1 dout16_reg_reg_140_ ( .D(n1058), .CK(clk), .RN(rstn), .Q(
        dout16_reg[140]) );
  DFFRHQX1 dout16_reg_reg_156_ ( .D(n1042), .CK(clk), .RN(rstn), .Q(
        dout16_reg[156]) );
  DFFRHQX1 dout16_reg_reg_172_ ( .D(n1026), .CK(clk), .RN(rstn), .Q(
        dout16_reg[172]) );
  DFFRHQX1 dout16_reg_reg_188_ ( .D(n1010), .CK(clk), .RN(rstn), .Q(
        dout16_reg[188]) );
  DFFRHQX1 dout16_reg_reg_11_ ( .D(n1187), .CK(clk), .RN(rstn), .Q(
        dout16_reg[11]) );
  DFFRHQX1 dout16_reg_reg_27_ ( .D(n1171), .CK(clk), .RN(rstn), .Q(
        dout16_reg[27]) );
  DFFRHQX1 dout16_reg_reg_43_ ( .D(n1155), .CK(clk), .RN(rstn), .Q(
        dout16_reg[43]) );
  DFFRHQX1 dout16_reg_reg_59_ ( .D(n1139), .CK(clk), .RN(rstn), .Q(
        dout16_reg[59]) );
  DFFRHQX1 dout16_reg_reg_75_ ( .D(n1123), .CK(clk), .RN(rstn), .Q(
        dout16_reg[75]) );
  DFFRHQX1 dout16_reg_reg_91_ ( .D(n1107), .CK(clk), .RN(rstn), .Q(
        dout16_reg[91]) );
  DFFRHQX1 dout16_reg_reg_107_ ( .D(n1091), .CK(clk), .RN(rstn), .Q(
        dout16_reg[107]) );
  DFFRHQX1 dout16_reg_reg_123_ ( .D(n1075), .CK(clk), .RN(rstn), .Q(
        dout16_reg[123]) );
  DFFRHQX1 dout16_reg_reg_139_ ( .D(n1059), .CK(clk), .RN(rstn), .Q(
        dout16_reg[139]) );
  DFFRHQX1 dout16_reg_reg_155_ ( .D(n1043), .CK(clk), .RN(rstn), .Q(
        dout16_reg[155]) );
  DFFRHQX1 dout16_reg_reg_171_ ( .D(n1027), .CK(clk), .RN(rstn), .Q(
        dout16_reg[171]) );
  DFFRHQX1 dout16_reg_reg_187_ ( .D(n1011), .CK(clk), .RN(rstn), .Q(
        dout16_reg[187]) );
  DFFRHQX1 dout16_reg_reg_10_ ( .D(n1188), .CK(clk), .RN(rstn), .Q(
        dout16_reg[10]) );
  DFFRHQX1 dout16_reg_reg_26_ ( .D(n1172), .CK(clk), .RN(rstn), .Q(
        dout16_reg[26]) );
  DFFRHQX1 dout16_reg_reg_42_ ( .D(n1156), .CK(clk), .RN(rstn), .Q(
        dout16_reg[42]) );
  DFFRHQX1 dout16_reg_reg_58_ ( .D(n1140), .CK(clk), .RN(rstn), .Q(
        dout16_reg[58]) );
  DFFRHQX1 dout16_reg_reg_74_ ( .D(n1124), .CK(clk), .RN(rstn), .Q(
        dout16_reg[74]) );
  DFFRHQX1 dout16_reg_reg_90_ ( .D(n1108), .CK(clk), .RN(rstn), .Q(
        dout16_reg[90]) );
  DFFRHQX1 dout16_reg_reg_106_ ( .D(n1092), .CK(clk), .RN(rstn), .Q(
        dout16_reg[106]) );
  DFFRHQX1 dout16_reg_reg_122_ ( .D(n1076), .CK(clk), .RN(rstn), .Q(
        dout16_reg[122]) );
  DFFRHQX1 dout16_reg_reg_138_ ( .D(n1060), .CK(clk), .RN(rstn), .Q(
        dout16_reg[138]) );
  DFFRHQX1 dout16_reg_reg_154_ ( .D(n1044), .CK(clk), .RN(rstn), .Q(
        dout16_reg[154]) );
  DFFRHQX1 dout16_reg_reg_170_ ( .D(n1028), .CK(clk), .RN(rstn), .Q(
        dout16_reg[170]) );
  DFFRHQX1 dout16_reg_reg_186_ ( .D(n1012), .CK(clk), .RN(rstn), .Q(
        dout16_reg[186]) );
  DFFRHQX1 dout16_reg_reg_9_ ( .D(n1189), .CK(clk), .RN(rstn), .Q(
        dout16_reg[9]) );
  DFFRHQX1 dout16_reg_reg_25_ ( .D(n1173), .CK(clk), .RN(rstn), .Q(
        dout16_reg[25]) );
  DFFRHQX1 dout16_reg_reg_41_ ( .D(n1157), .CK(clk), .RN(rstn), .Q(
        dout16_reg[41]) );
  DFFRHQX1 dout16_reg_reg_57_ ( .D(n1141), .CK(clk), .RN(rstn), .Q(
        dout16_reg[57]) );
  DFFRHQX1 dout16_reg_reg_73_ ( .D(n1125), .CK(clk), .RN(rstn), .Q(
        dout16_reg[73]) );
  DFFRHQX1 dout16_reg_reg_89_ ( .D(n1109), .CK(clk), .RN(rstn), .Q(
        dout16_reg[89]) );
  DFFRHQX1 dout16_reg_reg_105_ ( .D(n1093), .CK(clk), .RN(rstn), .Q(
        dout16_reg[105]) );
  DFFRHQX1 dout16_reg_reg_121_ ( .D(n1077), .CK(clk), .RN(rstn), .Q(
        dout16_reg[121]) );
  DFFRHQX1 dout16_reg_reg_137_ ( .D(n1061), .CK(clk), .RN(rstn), .Q(
        dout16_reg[137]) );
  DFFRHQX1 dout16_reg_reg_153_ ( .D(n1045), .CK(clk), .RN(rstn), .Q(
        dout16_reg[153]) );
  DFFRHQX1 dout16_reg_reg_169_ ( .D(n1029), .CK(clk), .RN(rstn), .Q(
        dout16_reg[169]) );
  DFFRHQX1 dout16_reg_reg_185_ ( .D(n1013), .CK(clk), .RN(rstn), .Q(
        dout16_reg[185]) );
  DFFRHQX1 dout16_reg_reg_8_ ( .D(n1190), .CK(clk), .RN(rstn), .Q(
        dout16_reg[8]) );
  DFFRHQX1 dout16_reg_reg_24_ ( .D(n1174), .CK(clk), .RN(rstn), .Q(
        dout16_reg[24]) );
  DFFRHQX1 dout16_reg_reg_40_ ( .D(n1158), .CK(clk), .RN(rstn), .Q(
        dout16_reg[40]) );
  DFFRHQX1 dout16_reg_reg_56_ ( .D(n1142), .CK(clk), .RN(rstn), .Q(
        dout16_reg[56]) );
  DFFRHQX1 dout16_reg_reg_72_ ( .D(n1126), .CK(clk), .RN(rstn), .Q(
        dout16_reg[72]) );
  DFFRHQX1 dout16_reg_reg_88_ ( .D(n1110), .CK(clk), .RN(rstn), .Q(
        dout16_reg[88]) );
  DFFRHQX1 dout16_reg_reg_104_ ( .D(n1094), .CK(clk), .RN(rstn), .Q(
        dout16_reg[104]) );
  DFFRHQX1 dout16_reg_reg_120_ ( .D(n1078), .CK(clk), .RN(rstn), .Q(
        dout16_reg[120]) );
  DFFRHQX1 dout16_reg_reg_136_ ( .D(n1062), .CK(clk), .RN(rstn), .Q(
        dout16_reg[136]) );
  DFFRHQX1 dout16_reg_reg_152_ ( .D(n1046), .CK(clk), .RN(rstn), .Q(
        dout16_reg[152]) );
  DFFRHQX1 dout16_reg_reg_168_ ( .D(n1030), .CK(clk), .RN(rstn), .Q(
        dout16_reg[168]) );
  DFFRHQX1 dout16_reg_reg_184_ ( .D(n1014), .CK(clk), .RN(rstn), .Q(
        dout16_reg[184]) );
  DFFRHQX1 dout16_reg_reg_7_ ( .D(n1191), .CK(clk), .RN(rstn), .Q(
        dout16_reg[7]) );
  DFFRHQX1 dout16_reg_reg_23_ ( .D(n1175), .CK(clk), .RN(rstn), .Q(
        dout16_reg[23]) );
  DFFRHQX1 dout16_reg_reg_39_ ( .D(n1159), .CK(clk), .RN(rstn), .Q(
        dout16_reg[39]) );
  DFFRHQX1 dout16_reg_reg_55_ ( .D(n1143), .CK(clk), .RN(rstn), .Q(
        dout16_reg[55]) );
  DFFRHQX1 dout16_reg_reg_71_ ( .D(n1127), .CK(clk), .RN(rstn), .Q(
        dout16_reg[71]) );
  DFFRHQX1 dout16_reg_reg_87_ ( .D(n1111), .CK(clk), .RN(rstn), .Q(
        dout16_reg[87]) );
  DFFRHQX1 dout16_reg_reg_103_ ( .D(n1095), .CK(clk), .RN(rstn), .Q(
        dout16_reg[103]) );
  DFFRHQX1 dout16_reg_reg_119_ ( .D(n1079), .CK(clk), .RN(rstn), .Q(
        dout16_reg[119]) );
  DFFRHQX1 dout16_reg_reg_135_ ( .D(n1063), .CK(clk), .RN(rstn), .Q(
        dout16_reg[135]) );
  DFFRHQX1 dout16_reg_reg_151_ ( .D(n1047), .CK(clk), .RN(rstn), .Q(
        dout16_reg[151]) );
  DFFRHQX1 dout16_reg_reg_167_ ( .D(n1031), .CK(clk), .RN(rstn), .Q(
        dout16_reg[167]) );
  DFFRHQX1 dout16_reg_reg_183_ ( .D(n1015), .CK(clk), .RN(rstn), .Q(
        dout16_reg[183]) );
  DFFRHQX1 dout16_reg_reg_6_ ( .D(n1192), .CK(clk), .RN(rstn), .Q(
        dout16_reg[6]) );
  DFFRHQX1 dout16_reg_reg_22_ ( .D(n1176), .CK(clk), .RN(rstn), .Q(
        dout16_reg[22]) );
  DFFRHQX1 dout16_reg_reg_38_ ( .D(n1160), .CK(clk), .RN(rstn), .Q(
        dout16_reg[38]) );
  DFFRHQX1 dout16_reg_reg_54_ ( .D(n1144), .CK(clk), .RN(rstn), .Q(
        dout16_reg[54]) );
  DFFRHQX1 dout16_reg_reg_70_ ( .D(n1128), .CK(clk), .RN(rstn), .Q(
        dout16_reg[70]) );
  DFFRHQX1 dout16_reg_reg_86_ ( .D(n1112), .CK(clk), .RN(rstn), .Q(
        dout16_reg[86]) );
  DFFRHQX1 dout16_reg_reg_102_ ( .D(n1096), .CK(clk), .RN(rstn), .Q(
        dout16_reg[102]) );
  DFFRHQX1 dout16_reg_reg_118_ ( .D(n1080), .CK(clk), .RN(rstn), .Q(
        dout16_reg[118]) );
  DFFRHQX1 dout16_reg_reg_134_ ( .D(n1064), .CK(clk), .RN(rstn), .Q(
        dout16_reg[134]) );
  DFFRHQX1 dout16_reg_reg_150_ ( .D(n1048), .CK(clk), .RN(rstn), .Q(
        dout16_reg[150]) );
  DFFRHQX1 dout16_reg_reg_166_ ( .D(n1032), .CK(clk), .RN(rstn), .Q(
        dout16_reg[166]) );
  DFFRHQX1 dout16_reg_reg_182_ ( .D(n1016), .CK(clk), .RN(rstn), .Q(
        dout16_reg[182]) );
  DFFRHQX1 dout16_reg_reg_5_ ( .D(n1193), .CK(clk), .RN(rstn), .Q(
        dout16_reg[5]) );
  DFFRHQX1 dout16_reg_reg_21_ ( .D(n1177), .CK(clk), .RN(rstn), .Q(
        dout16_reg[21]) );
  DFFRHQX1 dout16_reg_reg_37_ ( .D(n1161), .CK(clk), .RN(rstn), .Q(
        dout16_reg[37]) );
  DFFRHQX1 dout16_reg_reg_53_ ( .D(n1145), .CK(clk), .RN(rstn), .Q(
        dout16_reg[53]) );
  DFFRHQX1 dout16_reg_reg_69_ ( .D(n1129), .CK(clk), .RN(rstn), .Q(
        dout16_reg[69]) );
  DFFRHQX1 dout16_reg_reg_85_ ( .D(n1113), .CK(clk), .RN(rstn), .Q(
        dout16_reg[85]) );
  DFFRHQX1 dout16_reg_reg_101_ ( .D(n1097), .CK(clk), .RN(rstn), .Q(
        dout16_reg[101]) );
  DFFRHQX1 dout16_reg_reg_117_ ( .D(n1081), .CK(clk), .RN(rstn), .Q(
        dout16_reg[117]) );
  DFFRHQX1 dout16_reg_reg_133_ ( .D(n1065), .CK(clk), .RN(rstn), .Q(
        dout16_reg[133]) );
  DFFRHQX1 dout16_reg_reg_149_ ( .D(n1049), .CK(clk), .RN(rstn), .Q(
        dout16_reg[149]) );
  DFFRHQX1 dout16_reg_reg_165_ ( .D(n1033), .CK(clk), .RN(rstn), .Q(
        dout16_reg[165]) );
  DFFRHQX1 dout16_reg_reg_181_ ( .D(n1017), .CK(clk), .RN(rstn), .Q(
        dout16_reg[181]) );
  DFFRHQX1 dout16_reg_reg_4_ ( .D(n1194), .CK(clk), .RN(rstn), .Q(
        dout16_reg[4]) );
  DFFRHQX1 dout16_reg_reg_20_ ( .D(n1178), .CK(clk), .RN(rstn), .Q(
        dout16_reg[20]) );
  DFFRHQX1 dout16_reg_reg_36_ ( .D(n1162), .CK(clk), .RN(rstn), .Q(
        dout16_reg[36]) );
  DFFRHQX1 dout16_reg_reg_52_ ( .D(n1146), .CK(clk), .RN(rstn), .Q(
        dout16_reg[52]) );
  DFFRHQX1 dout16_reg_reg_68_ ( .D(n1130), .CK(clk), .RN(rstn), .Q(
        dout16_reg[68]) );
  DFFRHQX1 dout16_reg_reg_84_ ( .D(n1114), .CK(clk), .RN(rstn), .Q(
        dout16_reg[84]) );
  DFFRHQX1 dout16_reg_reg_100_ ( .D(n1098), .CK(clk), .RN(rstn), .Q(
        dout16_reg[100]) );
  DFFRHQX1 dout16_reg_reg_116_ ( .D(n1082), .CK(clk), .RN(rstn), .Q(
        dout16_reg[116]) );
  DFFRHQX1 dout16_reg_reg_132_ ( .D(n1066), .CK(clk), .RN(rstn), .Q(
        dout16_reg[132]) );
  DFFRHQX1 dout16_reg_reg_148_ ( .D(n1050), .CK(clk), .RN(rstn), .Q(
        dout16_reg[148]) );
  DFFRHQX1 dout16_reg_reg_164_ ( .D(n1034), .CK(clk), .RN(rstn), .Q(
        dout16_reg[164]) );
  DFFRHQX1 dout16_reg_reg_180_ ( .D(n1018), .CK(clk), .RN(rstn), .Q(
        dout16_reg[180]) );
  DFFRHQX1 dout16_reg_reg_3_ ( .D(n1195), .CK(clk), .RN(rstn), .Q(
        dout16_reg[3]) );
  DFFRHQX1 dout16_reg_reg_19_ ( .D(n1179), .CK(clk), .RN(rstn), .Q(
        dout16_reg[19]) );
  DFFRHQX1 dout16_reg_reg_35_ ( .D(n1163), .CK(clk), .RN(rstn), .Q(
        dout16_reg[35]) );
  DFFRHQX1 dout16_reg_reg_51_ ( .D(n1147), .CK(clk), .RN(rstn), .Q(
        dout16_reg[51]) );
  DFFRHQX1 dout16_reg_reg_67_ ( .D(n1131), .CK(clk), .RN(rstn), .Q(
        dout16_reg[67]) );
  DFFRHQX1 dout16_reg_reg_83_ ( .D(n1115), .CK(clk), .RN(rstn), .Q(
        dout16_reg[83]) );
  DFFRHQX1 dout16_reg_reg_99_ ( .D(n1099), .CK(clk), .RN(rstn), .Q(
        dout16_reg[99]) );
  DFFRHQX1 dout16_reg_reg_115_ ( .D(n1083), .CK(clk), .RN(rstn), .Q(
        dout16_reg[115]) );
  DFFRHQX1 dout16_reg_reg_131_ ( .D(n1067), .CK(clk), .RN(rstn), .Q(
        dout16_reg[131]) );
  DFFRHQX1 dout16_reg_reg_147_ ( .D(n1051), .CK(clk), .RN(rstn), .Q(
        dout16_reg[147]) );
  DFFRHQX1 dout16_reg_reg_163_ ( .D(n1035), .CK(clk), .RN(rstn), .Q(
        dout16_reg[163]) );
  DFFRHQX1 dout16_reg_reg_179_ ( .D(n1019), .CK(clk), .RN(rstn), .Q(
        dout16_reg[179]) );
  DFFRHQX1 dout16_reg_reg_2_ ( .D(n1196), .CK(clk), .RN(rstn), .Q(
        dout16_reg[2]) );
  DFFRHQX1 dout16_reg_reg_18_ ( .D(n1180), .CK(clk), .RN(rstn), .Q(
        dout16_reg[18]) );
  DFFRHQX1 dout16_reg_reg_34_ ( .D(n1164), .CK(clk), .RN(rstn), .Q(
        dout16_reg[34]) );
  DFFRHQX1 dout16_reg_reg_50_ ( .D(n1148), .CK(clk), .RN(rstn), .Q(
        dout16_reg[50]) );
  DFFRHQX1 dout16_reg_reg_66_ ( .D(n1132), .CK(clk), .RN(rstn), .Q(
        dout16_reg[66]) );
  DFFRHQX1 dout16_reg_reg_82_ ( .D(n1116), .CK(clk), .RN(rstn), .Q(
        dout16_reg[82]) );
  DFFRHQX1 dout16_reg_reg_98_ ( .D(n1100), .CK(clk), .RN(rstn), .Q(
        dout16_reg[98]) );
  DFFRHQX1 dout16_reg_reg_114_ ( .D(n1084), .CK(clk), .RN(rstn), .Q(
        dout16_reg[114]) );
  DFFRHQX1 dout16_reg_reg_130_ ( .D(n1068), .CK(clk), .RN(rstn), .Q(
        dout16_reg[130]) );
  DFFRHQX1 dout16_reg_reg_146_ ( .D(n1052), .CK(clk), .RN(rstn), .Q(
        dout16_reg[146]) );
  DFFRHQX1 dout16_reg_reg_162_ ( .D(n1036), .CK(clk), .RN(rstn), .Q(
        dout16_reg[162]) );
  DFFRHQX1 dout16_reg_reg_178_ ( .D(n1020), .CK(clk), .RN(rstn), .Q(
        dout16_reg[178]) );
  DFFRHQX1 dout16_reg_reg_1_ ( .D(n1197), .CK(clk), .RN(rstn), .Q(
        dout16_reg[1]) );
  DFFRHQX1 dout16_reg_reg_17_ ( .D(n1181), .CK(clk), .RN(rstn), .Q(
        dout16_reg[17]) );
  DFFRHQX1 dout16_reg_reg_33_ ( .D(n1165), .CK(clk), .RN(rstn), .Q(
        dout16_reg[33]) );
  DFFRHQX1 dout16_reg_reg_49_ ( .D(n1149), .CK(clk), .RN(rstn), .Q(
        dout16_reg[49]) );
  DFFRHQX1 dout16_reg_reg_65_ ( .D(n1133), .CK(clk), .RN(rstn), .Q(
        dout16_reg[65]) );
  DFFRHQX1 dout16_reg_reg_81_ ( .D(n1117), .CK(clk), .RN(rstn), .Q(
        dout16_reg[81]) );
  DFFRHQX1 dout16_reg_reg_97_ ( .D(n1101), .CK(clk), .RN(rstn), .Q(
        dout16_reg[97]) );
  DFFRHQX1 dout16_reg_reg_113_ ( .D(n1085), .CK(clk), .RN(rstn), .Q(
        dout16_reg[113]) );
  DFFRHQX1 dout16_reg_reg_129_ ( .D(n1069), .CK(clk), .RN(rstn), .Q(
        dout16_reg[129]) );
  DFFRHQX1 dout16_reg_reg_145_ ( .D(n1053), .CK(clk), .RN(rstn), .Q(
        dout16_reg[145]) );
  DFFRHQX1 dout16_reg_reg_161_ ( .D(n1037), .CK(clk), .RN(rstn), .Q(
        dout16_reg[161]) );
  DFFRHQX1 dout16_reg_reg_177_ ( .D(n1021), .CK(clk), .RN(rstn), .Q(
        dout16_reg[177]) );
  DFFRHQX1 dout16_reg_reg_0_ ( .D(n1198), .CK(clk), .RN(rstn), .Q(
        dout16_reg[0]) );
  DFFRHQX1 dout16_reg_reg_16_ ( .D(n1182), .CK(clk), .RN(rstn), .Q(
        dout16_reg[16]) );
  DFFRHQX1 dout16_reg_reg_32_ ( .D(n1166), .CK(clk), .RN(rstn), .Q(
        dout16_reg[32]) );
  DFFRHQX1 dout16_reg_reg_48_ ( .D(n1150), .CK(clk), .RN(rstn), .Q(
        dout16_reg[48]) );
  DFFRHQX1 dout16_reg_reg_64_ ( .D(n1134), .CK(clk), .RN(rstn), .Q(
        dout16_reg[64]) );
  DFFRHQX1 dout16_reg_reg_80_ ( .D(n1118), .CK(clk), .RN(rstn), .Q(
        dout16_reg[80]) );
  DFFRHQX1 dout16_reg_reg_96_ ( .D(n1102), .CK(clk), .RN(rstn), .Q(
        dout16_reg[96]) );
  DFFRHQX1 dout16_reg_reg_112_ ( .D(n1086), .CK(clk), .RN(rstn), .Q(
        dout16_reg[112]) );
  DFFRHQX1 dout16_reg_reg_128_ ( .D(n1070), .CK(clk), .RN(rstn), .Q(
        dout16_reg[128]) );
  DFFRHQX1 dout16_reg_reg_144_ ( .D(n1054), .CK(clk), .RN(rstn), .Q(
        dout16_reg[144]) );
  DFFRHQX1 dout16_reg_reg_160_ ( .D(n1038), .CK(clk), .RN(rstn), .Q(
        dout16_reg[160]) );
  DFFRHQX1 dout16_reg_reg_176_ ( .D(n1022), .CK(clk), .RN(rstn), .Q(
        dout16_reg[176]) );
  DFFRHQX1 dout8_reg_reg_15_ ( .D(n927), .CK(clk), .RN(rstn), .Q(dout8_reg[15]) );
  DFFRHQX1 dout8_reg_reg_31_ ( .D(n911), .CK(clk), .RN(rstn), .Q(dout8_reg[31]) );
  DFFRHQX1 dout8_reg_reg_47_ ( .D(n895), .CK(clk), .RN(rstn), .Q(dout8_reg[47]) );
  DFFRHQX1 dout8_reg_reg_63_ ( .D(n879), .CK(clk), .RN(rstn), .Q(dout8_reg[63]) );
  DFFRHQX1 dout8_reg_reg_14_ ( .D(n928), .CK(clk), .RN(rstn), .Q(dout8_reg[14]) );
  DFFRHQX1 dout8_reg_reg_30_ ( .D(n912), .CK(clk), .RN(rstn), .Q(dout8_reg[30]) );
  DFFRHQX1 dout8_reg_reg_46_ ( .D(n896), .CK(clk), .RN(rstn), .Q(dout8_reg[46]) );
  DFFRHQX1 dout8_reg_reg_62_ ( .D(n880), .CK(clk), .RN(rstn), .Q(dout8_reg[62]) );
  DFFRHQX1 dout8_reg_reg_13_ ( .D(n929), .CK(clk), .RN(rstn), .Q(dout8_reg[13]) );
  DFFRHQX1 dout8_reg_reg_29_ ( .D(n913), .CK(clk), .RN(rstn), .Q(dout8_reg[29]) );
  DFFRHQX1 dout8_reg_reg_45_ ( .D(n897), .CK(clk), .RN(rstn), .Q(dout8_reg[45]) );
  DFFRHQX1 dout8_reg_reg_61_ ( .D(n881), .CK(clk), .RN(rstn), .Q(dout8_reg[61]) );
  DFFRHQX1 dout8_reg_reg_12_ ( .D(n930), .CK(clk), .RN(rstn), .Q(dout8_reg[12]) );
  DFFRHQX1 dout8_reg_reg_28_ ( .D(n914), .CK(clk), .RN(rstn), .Q(dout8_reg[28]) );
  DFFRHQX1 dout8_reg_reg_44_ ( .D(n898), .CK(clk), .RN(rstn), .Q(dout8_reg[44]) );
  DFFRHQX1 dout8_reg_reg_60_ ( .D(n882), .CK(clk), .RN(rstn), .Q(dout8_reg[60]) );
  DFFRHQX1 dout8_reg_reg_11_ ( .D(n931), .CK(clk), .RN(rstn), .Q(dout8_reg[11]) );
  DFFRHQX1 dout8_reg_reg_27_ ( .D(n915), .CK(clk), .RN(rstn), .Q(dout8_reg[27]) );
  DFFRHQX1 dout8_reg_reg_43_ ( .D(n899), .CK(clk), .RN(rstn), .Q(dout8_reg[43]) );
  DFFRHQX1 dout8_reg_reg_59_ ( .D(n883), .CK(clk), .RN(rstn), .Q(dout8_reg[59]) );
  DFFRHQX1 dout8_reg_reg_10_ ( .D(n932), .CK(clk), .RN(rstn), .Q(dout8_reg[10]) );
  DFFRHQX1 dout8_reg_reg_26_ ( .D(n916), .CK(clk), .RN(rstn), .Q(dout8_reg[26]) );
  DFFRHQX1 dout8_reg_reg_42_ ( .D(n900), .CK(clk), .RN(rstn), .Q(dout8_reg[42]) );
  DFFRHQX1 dout8_reg_reg_58_ ( .D(n884), .CK(clk), .RN(rstn), .Q(dout8_reg[58]) );
  DFFRHQX1 dout8_reg_reg_9_ ( .D(n933), .CK(clk), .RN(rstn), .Q(dout8_reg[9])
         );
  DFFRHQX1 dout8_reg_reg_25_ ( .D(n917), .CK(clk), .RN(rstn), .Q(dout8_reg[25]) );
  DFFRHQX1 dout8_reg_reg_41_ ( .D(n901), .CK(clk), .RN(rstn), .Q(dout8_reg[41]) );
  DFFRHQX1 dout8_reg_reg_57_ ( .D(n885), .CK(clk), .RN(rstn), .Q(dout8_reg[57]) );
  DFFRHQX1 dout8_reg_reg_8_ ( .D(n934), .CK(clk), .RN(rstn), .Q(dout8_reg[8])
         );
  DFFRHQX1 dout8_reg_reg_24_ ( .D(n918), .CK(clk), .RN(rstn), .Q(dout8_reg[24]) );
  DFFRHQX1 dout8_reg_reg_40_ ( .D(n902), .CK(clk), .RN(rstn), .Q(dout8_reg[40]) );
  DFFRHQX1 dout8_reg_reg_56_ ( .D(n886), .CK(clk), .RN(rstn), .Q(dout8_reg[56]) );
  DFFRHQX1 dout8_reg_reg_7_ ( .D(n935), .CK(clk), .RN(rstn), .Q(dout8_reg[7])
         );
  DFFRHQX1 dout8_reg_reg_23_ ( .D(n919), .CK(clk), .RN(rstn), .Q(dout8_reg[23]) );
  DFFRHQX1 dout8_reg_reg_39_ ( .D(n903), .CK(clk), .RN(rstn), .Q(dout8_reg[39]) );
  DFFRHQX1 dout8_reg_reg_55_ ( .D(n887), .CK(clk), .RN(rstn), .Q(dout8_reg[55]) );
  DFFRHQX1 dout8_reg_reg_6_ ( .D(n936), .CK(clk), .RN(rstn), .Q(dout8_reg[6])
         );
  DFFRHQX1 dout8_reg_reg_22_ ( .D(n920), .CK(clk), .RN(rstn), .Q(dout8_reg[22]) );
  DFFRHQX1 dout8_reg_reg_38_ ( .D(n904), .CK(clk), .RN(rstn), .Q(dout8_reg[38]) );
  DFFRHQX1 dout8_reg_reg_54_ ( .D(n888), .CK(clk), .RN(rstn), .Q(dout8_reg[54]) );
  DFFRHQX1 dout8_reg_reg_5_ ( .D(n937), .CK(clk), .RN(rstn), .Q(dout8_reg[5])
         );
  DFFRHQX1 dout8_reg_reg_21_ ( .D(n921), .CK(clk), .RN(rstn), .Q(dout8_reg[21]) );
  DFFRHQX1 dout8_reg_reg_37_ ( .D(n905), .CK(clk), .RN(rstn), .Q(dout8_reg[37]) );
  DFFRHQX1 dout8_reg_reg_53_ ( .D(n889), .CK(clk), .RN(rstn), .Q(dout8_reg[53]) );
  DFFRHQX1 dout8_reg_reg_4_ ( .D(n938), .CK(clk), .RN(rstn), .Q(dout8_reg[4])
         );
  DFFRHQX1 dout8_reg_reg_20_ ( .D(n922), .CK(clk), .RN(rstn), .Q(dout8_reg[20]) );
  DFFRHQX1 dout8_reg_reg_36_ ( .D(n906), .CK(clk), .RN(rstn), .Q(dout8_reg[36]) );
  DFFRHQX1 dout8_reg_reg_52_ ( .D(n890), .CK(clk), .RN(rstn), .Q(dout8_reg[52]) );
  DFFRHQX1 dout8_reg_reg_3_ ( .D(n939), .CK(clk), .RN(rstn), .Q(dout8_reg[3])
         );
  DFFRHQX1 dout8_reg_reg_19_ ( .D(n923), .CK(clk), .RN(rstn), .Q(dout8_reg[19]) );
  DFFRHQX1 dout8_reg_reg_35_ ( .D(n907), .CK(clk), .RN(rstn), .Q(dout8_reg[35]) );
  DFFRHQX1 dout8_reg_reg_51_ ( .D(n891), .CK(clk), .RN(rstn), .Q(dout8_reg[51]) );
  DFFRHQX1 dout8_reg_reg_2_ ( .D(n940), .CK(clk), .RN(rstn), .Q(dout8_reg[2])
         );
  DFFRHQX1 dout8_reg_reg_18_ ( .D(n924), .CK(clk), .RN(rstn), .Q(dout8_reg[18]) );
  DFFRHQX1 dout8_reg_reg_34_ ( .D(n908), .CK(clk), .RN(rstn), .Q(dout8_reg[34]) );
  DFFRHQX1 dout8_reg_reg_50_ ( .D(n892), .CK(clk), .RN(rstn), .Q(dout8_reg[50]) );
  DFFRHQX1 dout8_reg_reg_1_ ( .D(n941), .CK(clk), .RN(rstn), .Q(dout8_reg[1])
         );
  DFFRHQX1 dout8_reg_reg_17_ ( .D(n925), .CK(clk), .RN(rstn), .Q(dout8_reg[17]) );
  DFFRHQX1 dout8_reg_reg_33_ ( .D(n909), .CK(clk), .RN(rstn), .Q(dout8_reg[33]) );
  DFFRHQX1 dout8_reg_reg_49_ ( .D(n893), .CK(clk), .RN(rstn), .Q(dout8_reg[49]) );
  DFFRHQX1 dout8_reg_reg_0_ ( .D(n942), .CK(clk), .RN(rstn), .Q(dout8_reg[0])
         );
  DFFRHQX1 dout8_reg_reg_16_ ( .D(n926), .CK(clk), .RN(rstn), .Q(dout8_reg[16]) );
  DFFRHQX1 dout8_reg_reg_32_ ( .D(n910), .CK(clk), .RN(rstn), .Q(dout8_reg[32]) );
  DFFRHQX1 dout8_reg_reg_48_ ( .D(n894), .CK(clk), .RN(rstn), .Q(dout8_reg[48]) );
  DFFRHQX1 count_reg_0_ ( .D(N1114), .CK(clk), .RN(rstn), .Q(count[0]) );
  DFFRHQX1 count_reg_1_ ( .D(N1115), .CK(clk), .RN(rstn), .Q(count[1]) );
  DFFRHQX1 count_reg_3_ ( .D(N1117), .CK(clk), .RN(rstn), .Q(count[3]) );
  DFFRHQX1 count_reg_2_ ( .D(N1116), .CK(clk), .RN(rstn), .Q(count[2]) );
  DFFRHQX1 mode_reg_reg_1_ ( .D(mode[1]), .CK(clk), .RN(rstn), .Q(mode_reg[1])
         );
  DFFRHQX1 mode_reg_reg_0_ ( .D(mode[0]), .CK(clk), .RN(rstn), .Q(mode_reg[0])
         );
  DFFRHQX1 s2p_ready_reg ( .D(N1119), .CK(clk), .RN(rstn), .Q(s2p_ready) );
  AND2X2 U5 ( .A(n737), .B(n1248), .Y(n1) );
  AND2X2 U6 ( .A(n740), .B(start), .Y(n2) );
  AND2X2 U7 ( .A(n736), .B(start), .Y(n3) );
  AND2X2 U8 ( .A(start), .B(n733), .Y(n4) );
  INVX1 U9 ( .A(n312), .Y(n310) );
  INVX1 U10 ( .A(n312), .Y(n308) );
  INVX1 U11 ( .A(n312), .Y(n309) );
  INVX1 U12 ( .A(n312), .Y(n311) );
  INVX1 U13 ( .A(n1), .Y(n293) );
  INVX1 U14 ( .A(n1), .Y(n301) );
  INVX1 U15 ( .A(n1), .Y(n298) );
  INVX1 U16 ( .A(n1), .Y(n297) );
  INVX1 U17 ( .A(n1), .Y(n296) );
  INVX1 U18 ( .A(n1), .Y(n295) );
  INVX1 U19 ( .A(n1), .Y(n294) );
  INVX1 U20 ( .A(n1), .Y(n292) );
  INVX1 U21 ( .A(n1), .Y(n291) );
  INVX1 U22 ( .A(n1), .Y(n290) );
  INVX1 U23 ( .A(n1), .Y(n303) );
  INVX1 U24 ( .A(n1), .Y(n302) );
  INVX1 U25 ( .A(n1), .Y(n300) );
  INVX1 U26 ( .A(n1), .Y(n299) );
  INVX1 U27 ( .A(n269), .Y(n267) );
  INVX1 U28 ( .A(n269), .Y(n268) );
  INVX1 U29 ( .A(n331), .Y(n319) );
  INVX1 U30 ( .A(n331), .Y(n320) );
  INVX1 U31 ( .A(n331), .Y(n321) );
  INVX1 U32 ( .A(n331), .Y(n322) );
  INVX1 U33 ( .A(n331), .Y(n323) );
  INVX1 U34 ( .A(n331), .Y(n324) );
  INVX1 U35 ( .A(n331), .Y(n325) );
  INVX1 U36 ( .A(n331), .Y(n326) );
  INVX1 U37 ( .A(n331), .Y(n327) );
  INVX1 U38 ( .A(n331), .Y(n328) );
  INVX1 U39 ( .A(n331), .Y(n329) );
  INVX1 U40 ( .A(n331), .Y(n330) );
  INVX1 U41 ( .A(n4), .Y(n313) );
  INVX1 U42 ( .A(n3), .Y(n306) );
  INVX1 U43 ( .A(n3), .Y(n304) );
  INVX1 U44 ( .A(n3), .Y(n305) );
  INVX1 U45 ( .A(n3), .Y(n307) );
  INVX1 U46 ( .A(n2), .Y(n285) );
  INVX1 U47 ( .A(n2), .Y(n281) );
  INVX1 U48 ( .A(n2), .Y(n279) );
  INVX1 U49 ( .A(n2), .Y(n280) );
  INVX1 U50 ( .A(n2), .Y(n282) );
  INVX1 U51 ( .A(n2), .Y(n283) );
  INVX1 U52 ( .A(n2), .Y(n284) );
  INVX1 U53 ( .A(n2), .Y(n286) );
  INVX1 U54 ( .A(n2), .Y(n287) );
  INVX1 U55 ( .A(n2), .Y(n288) );
  INVX1 U56 ( .A(n2), .Y(n289) );
  INVX1 U57 ( .A(n4), .Y(n314) );
  INVX1 U58 ( .A(n317), .Y(n316) );
  INVX1 U59 ( .A(n317), .Y(n315) );
  INVX1 U60 ( .A(n734), .Y(n312) );
  INVX1 U61 ( .A(n278), .Y(n271) );
  INVX1 U62 ( .A(n278), .Y(n270) );
  INVX1 U63 ( .A(n278), .Y(n272) );
  INVX1 U64 ( .A(n278), .Y(n273) );
  INVX1 U65 ( .A(n278), .Y(n274) );
  INVX1 U66 ( .A(n278), .Y(n277) );
  INVX1 U67 ( .A(n278), .Y(n276) );
  INVX1 U68 ( .A(n266), .Y(n265) );
  INVX1 U69 ( .A(n278), .Y(n275) );
  INVX1 U70 ( .A(n266), .Y(n262) );
  INVX1 U71 ( .A(n266), .Y(n264) );
  INVX1 U72 ( .A(n266), .Y(n263) );
  INVX1 U73 ( .A(n331), .Y(n318) );
  INVX1 U74 ( .A(N30), .Y(n331) );
  INVX1 U75 ( .A(n742), .Y(n269) );
  OAI22X1 U76 ( .A0(n311), .A1(n600), .B0(n1255), .B1(n306), .Y(n928) );
  OAI22X1 U77 ( .A0(n310), .A1(n592), .B0(n1254), .B1(n304), .Y(n927) );
  OAI22X1 U78 ( .A0(n295), .A1(n432), .B0(n1260), .B1(n279), .Y(n1189) );
  OAI22X1 U79 ( .A0(n296), .A1(n416), .B0(n1259), .B1(n286), .Y(n1188) );
  OAI22X1 U80 ( .A0(n293), .A1(n400), .B0(n1258), .B1(n287), .Y(n1187) );
  OAI22X1 U81 ( .A0(n294), .A1(n384), .B0(n1257), .B1(n286), .Y(n1186) );
  OAI22X1 U82 ( .A0(n299), .A1(n368), .B0(n1256), .B1(n281), .Y(n1185) );
  OAI22X1 U83 ( .A0(n298), .A1(n352), .B0(n1255), .B1(n286), .Y(n1184) );
  OAI22X1 U84 ( .A0(n297), .A1(n336), .B0(n1254), .B1(n287), .Y(n1183) );
  OAI22X1 U85 ( .A0(n310), .A1(n624), .B0(n1258), .B1(n307), .Y(n931) );
  OAI22X1 U86 ( .A0(n309), .A1(n608), .B0(n1256), .B1(n306), .Y(n929) );
  OAI22X1 U87 ( .A0(n308), .A1(n616), .B0(n1257), .B1(n306), .Y(n930) );
  OAI22X1 U88 ( .A0(n310), .A1(n716), .B0(n305), .B1(n715), .Y(n878) );
  OAI22X1 U89 ( .A0(n309), .A1(n715), .B0(n307), .B1(n714), .Y(n894) );
  OAI22X1 U90 ( .A0(n310), .A1(n714), .B0(n306), .B1(n713), .Y(n910) );
  OAI22X1 U91 ( .A0(n734), .A1(n713), .B0(n306), .B1(n712), .Y(n926) );
  OAI22X1 U92 ( .A0(n308), .A1(n708), .B0(n305), .B1(n707), .Y(n877) );
  OAI22X1 U93 ( .A0(n309), .A1(n707), .B0(n307), .B1(n706), .Y(n893) );
  OAI22X1 U94 ( .A0(n310), .A1(n706), .B0(n305), .B1(n705), .Y(n909) );
  OAI22X1 U95 ( .A0(n734), .A1(n705), .B0(n305), .B1(n704), .Y(n925) );
  OAI22X1 U96 ( .A0(n309), .A1(n700), .B0(n305), .B1(n699), .Y(n876) );
  OAI22X1 U97 ( .A0(n309), .A1(n699), .B0(n306), .B1(n698), .Y(n892) );
  OAI22X1 U98 ( .A0(n310), .A1(n698), .B0(n307), .B1(n697), .Y(n908) );
  OAI22X1 U99 ( .A0(n734), .A1(n697), .B0(n306), .B1(n696), .Y(n924) );
  OAI22X1 U100 ( .A0(n308), .A1(n692), .B0(n305), .B1(n691), .Y(n875) );
  OAI22X1 U101 ( .A0(n309), .A1(n691), .B0(n306), .B1(n690), .Y(n891) );
  OAI22X1 U102 ( .A0(n310), .A1(n690), .B0(n306), .B1(n689), .Y(n907) );
  OAI22X1 U103 ( .A0(n734), .A1(n689), .B0(n304), .B1(n688), .Y(n923) );
  OAI22X1 U104 ( .A0(n308), .A1(n684), .B0(n305), .B1(n683), .Y(n874) );
  OAI22X1 U105 ( .A0(n309), .A1(n683), .B0(n306), .B1(n682), .Y(n890) );
  OAI22X1 U106 ( .A0(n310), .A1(n682), .B0(n304), .B1(n681), .Y(n906) );
  OAI22X1 U107 ( .A0(n311), .A1(n681), .B0(n306), .B1(n680), .Y(n922) );
  OAI22X1 U108 ( .A0(n308), .A1(n676), .B0(n305), .B1(n675), .Y(n873) );
  OAI22X1 U109 ( .A0(n309), .A1(n675), .B0(n306), .B1(n674), .Y(n889) );
  OAI22X1 U110 ( .A0(n310), .A1(n674), .B0(n307), .B1(n673), .Y(n905) );
  OAI22X1 U111 ( .A0(n311), .A1(n673), .B0(n306), .B1(n672), .Y(n921) );
  OAI22X1 U112 ( .A0(n308), .A1(n668), .B0(n305), .B1(n667), .Y(n872) );
  OAI22X1 U113 ( .A0(n309), .A1(n667), .B0(n306), .B1(n666), .Y(n888) );
  OAI22X1 U114 ( .A0(n310), .A1(n666), .B0(n307), .B1(n665), .Y(n904) );
  OAI22X1 U115 ( .A0(n311), .A1(n665), .B0(n304), .B1(n664), .Y(n920) );
  OAI22X1 U116 ( .A0(n308), .A1(n660), .B0(n305), .B1(n659), .Y(n871) );
  OAI22X1 U117 ( .A0(n309), .A1(n659), .B0(n306), .B1(n658), .Y(n887) );
  OAI22X1 U118 ( .A0(n310), .A1(n658), .B0(n307), .B1(n657), .Y(n903) );
  OAI22X1 U119 ( .A0(n311), .A1(n657), .B0(n305), .B1(n656), .Y(n919) );
  OAI22X1 U120 ( .A0(n308), .A1(n652), .B0(n305), .B1(n651), .Y(n870) );
  OAI22X1 U121 ( .A0(n734), .A1(n651), .B0(n306), .B1(n650), .Y(n886) );
  OAI22X1 U122 ( .A0(n310), .A1(n650), .B0(n307), .B1(n649), .Y(n902) );
  OAI22X1 U123 ( .A0(n311), .A1(n649), .B0(n306), .B1(n648), .Y(n918) );
  OAI22X1 U124 ( .A0(n308), .A1(n644), .B0(n305), .B1(n643), .Y(n869) );
  OAI22X1 U125 ( .A0(n734), .A1(n643), .B0(n306), .B1(n642), .Y(n885) );
  OAI22X1 U126 ( .A0(n310), .A1(n642), .B0(n307), .B1(n641), .Y(n901) );
  OAI22X1 U127 ( .A0(n311), .A1(n641), .B0(n305), .B1(n640), .Y(n917) );
  OAI22X1 U128 ( .A0(n308), .A1(n636), .B0(n305), .B1(n635), .Y(n868) );
  OAI22X1 U129 ( .A0(n734), .A1(n635), .B0(n306), .B1(n634), .Y(n884) );
  OAI22X1 U130 ( .A0(n310), .A1(n634), .B0(n307), .B1(n633), .Y(n900) );
  OAI22X1 U131 ( .A0(n311), .A1(n633), .B0(n307), .B1(n632), .Y(n916) );
  OAI22X1 U132 ( .A0(n308), .A1(n628), .B0(n305), .B1(n627), .Y(n867) );
  OAI22X1 U133 ( .A0(n734), .A1(n627), .B0(n306), .B1(n626), .Y(n883) );
  OAI22X1 U134 ( .A0(n310), .A1(n626), .B0(n307), .B1(n625), .Y(n899) );
  OAI22X1 U135 ( .A0(n311), .A1(n625), .B0(n305), .B1(n624), .Y(n915) );
  OAI22X1 U136 ( .A0(n308), .A1(n620), .B0(n304), .B1(n619), .Y(n866) );
  OAI22X1 U137 ( .A0(n734), .A1(n619), .B0(n306), .B1(n618), .Y(n882) );
  OAI22X1 U138 ( .A0(n309), .A1(n618), .B0(n307), .B1(n617), .Y(n898) );
  OAI22X1 U139 ( .A0(n311), .A1(n617), .B0(n304), .B1(n616), .Y(n914) );
  OAI22X1 U140 ( .A0(n308), .A1(n612), .B0(n304), .B1(n611), .Y(n865) );
  OAI22X1 U141 ( .A0(n734), .A1(n611), .B0(n306), .B1(n610), .Y(n881) );
  OAI22X1 U142 ( .A0(n309), .A1(n610), .B0(n307), .B1(n609), .Y(n897) );
  OAI22X1 U143 ( .A0(n311), .A1(n609), .B0(n306), .B1(n608), .Y(n913) );
  OAI22X1 U144 ( .A0(n308), .A1(n604), .B0(n304), .B1(n603), .Y(n864) );
  OAI22X1 U145 ( .A0(n734), .A1(n603), .B0(n306), .B1(n602), .Y(n880) );
  OAI22X1 U146 ( .A0(n309), .A1(n602), .B0(n307), .B1(n601), .Y(n896) );
  OAI22X1 U147 ( .A0(n311), .A1(n601), .B0(n305), .B1(n600), .Y(n912) );
  OAI22X1 U148 ( .A0(n311), .A1(n596), .B0(n304), .B1(n595), .Y(n863) );
  OAI22X1 U149 ( .A0(n311), .A1(n595), .B0(n305), .B1(n594), .Y(n879) );
  OAI22X1 U150 ( .A0(n309), .A1(n594), .B0(n307), .B1(n593), .Y(n895) );
  OAI22X1 U151 ( .A0(n311), .A1(n593), .B0(n307), .B1(n592), .Y(n911) );
  OAI22X1 U152 ( .A0(n294), .A1(n588), .B0(n284), .B1(n587), .Y(n1006) );
  OAI22X1 U153 ( .A0(n293), .A1(n587), .B0(n282), .B1(n586), .Y(n1022) );
  OAI22X1 U154 ( .A0(n291), .A1(n586), .B0(n283), .B1(n585), .Y(n1038) );
  OAI22X1 U155 ( .A0(n290), .A1(n585), .B0(n281), .B1(n584), .Y(n1054) );
  OAI22X1 U156 ( .A0(n300), .A1(n579), .B0(n285), .B1(n578), .Y(n1150) );
  OAI22X1 U157 ( .A0(n299), .A1(n578), .B0(n288), .B1(n577), .Y(n1166) );
  OAI22X1 U158 ( .A0(n302), .A1(n577), .B0(n285), .B1(n576), .Y(n1182) );
  OAI22X1 U159 ( .A0(n294), .A1(n572), .B0(n280), .B1(n571), .Y(n1005) );
  OAI22X1 U160 ( .A0(n293), .A1(n571), .B0(n282), .B1(n570), .Y(n1021) );
  OAI22X1 U161 ( .A0(n291), .A1(n570), .B0(n283), .B1(n569), .Y(n1037) );
  OAI22X1 U162 ( .A0(n290), .A1(n569), .B0(n282), .B1(n568), .Y(n1053) );
  OAI22X1 U163 ( .A0(n298), .A1(n568), .B0(n284), .B1(n567), .Y(n1069) );
  OAI22X1 U164 ( .A0(n301), .A1(n567), .B0(n285), .B1(n566), .Y(n1085) );
  OAI22X1 U165 ( .A0(n303), .A1(n566), .B0(n287), .B1(n565), .Y(n1101) );
  OAI22X1 U166 ( .A0(n302), .A1(n565), .B0(n288), .B1(n564), .Y(n1117) );
  OAI22X1 U167 ( .A0(n301), .A1(n564), .B0(n285), .B1(n563), .Y(n1133) );
  OAI22X1 U168 ( .A0(n300), .A1(n563), .B0(n284), .B1(n562), .Y(n1149) );
  OAI22X1 U169 ( .A0(n299), .A1(n562), .B0(n285), .B1(n561), .Y(n1165) );
  OAI22X1 U170 ( .A0(n290), .A1(n561), .B0(n284), .B1(n560), .Y(n1181) );
  OAI22X1 U171 ( .A0(n294), .A1(n556), .B0(n289), .B1(n555), .Y(n1004) );
  OAI22X1 U172 ( .A0(n293), .A1(n555), .B0(n281), .B1(n554), .Y(n1020) );
  OAI22X1 U173 ( .A0(n291), .A1(n554), .B0(n283), .B1(n553), .Y(n1036) );
  OAI22X1 U174 ( .A0(n290), .A1(n553), .B0(n283), .B1(n552), .Y(n1052) );
  OAI22X1 U175 ( .A0(n300), .A1(n552), .B0(n284), .B1(n551), .Y(n1068) );
  OAI22X1 U176 ( .A0(n302), .A1(n551), .B0(n285), .B1(n550), .Y(n1084) );
  OAI22X1 U177 ( .A0(n303), .A1(n550), .B0(n287), .B1(n549), .Y(n1100) );
  OAI22X1 U178 ( .A0(n302), .A1(n549), .B0(n288), .B1(n548), .Y(n1116) );
  OAI22X1 U179 ( .A0(n301), .A1(n548), .B0(n284), .B1(n547), .Y(n1132) );
  OAI22X1 U180 ( .A0(n300), .A1(n547), .B0(n280), .B1(n546), .Y(n1148) );
  OAI22X1 U181 ( .A0(n299), .A1(n546), .B0(n284), .B1(n545), .Y(n1164) );
  OAI22X1 U182 ( .A0(n298), .A1(n545), .B0(n282), .B1(n544), .Y(n1180) );
  OAI22X1 U183 ( .A0(n294), .A1(n540), .B0(n279), .B1(n539), .Y(n1003) );
  OAI22X1 U184 ( .A0(n293), .A1(n539), .B0(n281), .B1(n538), .Y(n1019) );
  OAI22X1 U185 ( .A0(n291), .A1(n538), .B0(n283), .B1(n537), .Y(n1035) );
  OAI22X1 U186 ( .A0(n290), .A1(n537), .B0(n288), .B1(n536), .Y(n1051) );
  OAI22X1 U187 ( .A0(n296), .A1(n536), .B0(n284), .B1(n535), .Y(n1067) );
  OAI22X1 U188 ( .A0(n301), .A1(n535), .B0(n285), .B1(n534), .Y(n1083) );
  OAI22X1 U189 ( .A0(n303), .A1(n534), .B0(n287), .B1(n533), .Y(n1099) );
  OAI22X1 U190 ( .A0(n302), .A1(n533), .B0(n288), .B1(n532), .Y(n1115) );
  OAI22X1 U191 ( .A0(n301), .A1(n532), .B0(n280), .B1(n531), .Y(n1131) );
  OAI22X1 U192 ( .A0(n300), .A1(n531), .B0(n289), .B1(n530), .Y(n1147) );
  OAI22X1 U193 ( .A0(n299), .A1(n530), .B0(n289), .B1(n529), .Y(n1163) );
  OAI22X1 U194 ( .A0(n298), .A1(n529), .B0(n283), .B1(n528), .Y(n1179) );
  OAI22X1 U195 ( .A0(n294), .A1(n524), .B0(n281), .B1(n523), .Y(n1002) );
  OAI22X1 U196 ( .A0(n293), .A1(n523), .B0(n281), .B1(n522), .Y(n1018) );
  OAI22X1 U197 ( .A0(n292), .A1(n522), .B0(n283), .B1(n521), .Y(n1034) );
  OAI22X1 U198 ( .A0(n290), .A1(n521), .B0(n285), .B1(n520), .Y(n1050) );
  OAI22X1 U199 ( .A0(n293), .A1(n520), .B0(n284), .B1(n519), .Y(n1066) );
  OAI22X1 U200 ( .A0(n303), .A1(n519), .B0(n285), .B1(n518), .Y(n1082) );
  OAI22X1 U201 ( .A0(n303), .A1(n518), .B0(n286), .B1(n517), .Y(n1098) );
  OAI22X1 U202 ( .A0(n302), .A1(n517), .B0(n288), .B1(n516), .Y(n1114) );
  OAI22X1 U203 ( .A0(n301), .A1(n516), .B0(n289), .B1(n515), .Y(n1130) );
  OAI22X1 U204 ( .A0(n300), .A1(n515), .B0(n279), .B1(n514), .Y(n1146) );
  OAI22X1 U205 ( .A0(n299), .A1(n514), .B0(n289), .B1(n513), .Y(n1162) );
  OAI22X1 U206 ( .A0(n298), .A1(n513), .B0(n288), .B1(n512), .Y(n1178) );
  OAI22X1 U207 ( .A0(n294), .A1(n508), .B0(n282), .B1(n507), .Y(n1001) );
  OAI22X1 U208 ( .A0(n293), .A1(n507), .B0(n281), .B1(n506), .Y(n1017) );
  OAI22X1 U209 ( .A0(n292), .A1(n506), .B0(n282), .B1(n505), .Y(n1033) );
  OAI22X1 U210 ( .A0(n290), .A1(n505), .B0(n281), .B1(n504), .Y(n1049) );
  OAI22X1 U211 ( .A0(n294), .A1(n504), .B0(n284), .B1(n503), .Y(n1065) );
  OAI22X1 U212 ( .A0(n290), .A1(n503), .B0(n285), .B1(n502), .Y(n1081) );
  OAI22X1 U213 ( .A0(n303), .A1(n502), .B0(n286), .B1(n501), .Y(n1097) );
  OAI22X1 U214 ( .A0(n302), .A1(n501), .B0(n288), .B1(n500), .Y(n1113) );
  OAI22X1 U215 ( .A0(n301), .A1(n500), .B0(n279), .B1(n499), .Y(n1129) );
  OAI22X1 U216 ( .A0(n300), .A1(n499), .B0(n281), .B1(n498), .Y(n1145) );
  OAI22X1 U217 ( .A0(n299), .A1(n498), .B0(n289), .B1(n497), .Y(n1161) );
  OAI22X1 U218 ( .A0(n298), .A1(n497), .B0(n285), .B1(n496), .Y(n1177) );
  OAI22X1 U219 ( .A0(n294), .A1(n492), .B0(n283), .B1(n491), .Y(n1000) );
  OAI22X1 U220 ( .A0(n293), .A1(n491), .B0(n281), .B1(n490), .Y(n1016) );
  OAI22X1 U221 ( .A0(n292), .A1(n490), .B0(n282), .B1(n489), .Y(n1032) );
  OAI22X1 U222 ( .A0(n290), .A1(n489), .B0(n282), .B1(n488), .Y(n1048) );
  OAI22X1 U223 ( .A0(n299), .A1(n488), .B0(n284), .B1(n487), .Y(n1064) );
  OAI22X1 U224 ( .A0(n295), .A1(n487), .B0(n285), .B1(n486), .Y(n1080) );
  OAI22X1 U225 ( .A0(n293), .A1(n486), .B0(n286), .B1(n485), .Y(n1096) );
  OAI22X1 U226 ( .A0(n302), .A1(n485), .B0(n288), .B1(n484), .Y(n1112) );
  OAI22X1 U227 ( .A0(n301), .A1(n484), .B0(n281), .B1(n483), .Y(n1128) );
  OAI22X1 U228 ( .A0(n294), .A1(n483), .B0(n282), .B1(n482), .Y(n1144) );
  OAI22X1 U229 ( .A0(n299), .A1(n482), .B0(n289), .B1(n481), .Y(n1160) );
  OAI22X1 U230 ( .A0(n298), .A1(n481), .B0(n280), .B1(n480), .Y(n1176) );
  OAI22X1 U231 ( .A0(n295), .A1(n476), .B0(n288), .B1(n475), .Y(n999) );
  OAI22X1 U232 ( .A0(n293), .A1(n475), .B0(n281), .B1(n474), .Y(n1015) );
  OAI22X1 U233 ( .A0(n292), .A1(n474), .B0(n282), .B1(n473), .Y(n1031) );
  OAI22X1 U234 ( .A0(n290), .A1(n473), .B0(n283), .B1(n472), .Y(n1047) );
  OAI22X1 U235 ( .A0(n297), .A1(n456), .B0(n284), .B1(n455), .Y(n1062) );
  OAI22X1 U236 ( .A0(n296), .A1(n455), .B0(n285), .B1(n454), .Y(n1078) );
  OAI22X1 U237 ( .A0(n294), .A1(n454), .B0(n286), .B1(n453), .Y(n1094) );
  OAI22X1 U238 ( .A0(n302), .A1(n453), .B0(n287), .B1(n452), .Y(n1110) );
  OAI22X1 U239 ( .A0(n301), .A1(n452), .B0(n282), .B1(n451), .Y(n1126) );
  OAI22X1 U240 ( .A0(n300), .A1(n451), .B0(n283), .B1(n450), .Y(n1142) );
  OAI22X1 U241 ( .A0(n299), .A1(n450), .B0(n289), .B1(n449), .Y(n1158) );
  OAI22X1 U242 ( .A0(n298), .A1(n449), .B0(n286), .B1(n448), .Y(n1174) );
  OAI22X1 U243 ( .A0(n295), .A1(n444), .B0(n287), .B1(n443), .Y(n997) );
  OAI22X1 U244 ( .A0(n293), .A1(n443), .B0(n281), .B1(n442), .Y(n1013) );
  OAI22X1 U245 ( .A0(n292), .A1(n442), .B0(n282), .B1(n441), .Y(n1029) );
  OAI22X1 U246 ( .A0(n291), .A1(n441), .B0(n283), .B1(n440), .Y(n1045) );
  OAI22X1 U247 ( .A0(n298), .A1(n440), .B0(n284), .B1(n439), .Y(n1061) );
  OAI22X1 U248 ( .A0(n293), .A1(n439), .B0(n285), .B1(n438), .Y(n1077) );
  OAI22X1 U249 ( .A0(n300), .A1(n438), .B0(n286), .B1(n437), .Y(n1093) );
  OAI22X1 U250 ( .A0(n303), .A1(n437), .B0(n287), .B1(n436), .Y(n1109) );
  OAI22X1 U251 ( .A0(n301), .A1(n436), .B0(n283), .B1(n435), .Y(n1125) );
  OAI22X1 U252 ( .A0(n295), .A1(n435), .B0(n287), .B1(n434), .Y(n1141) );
  OAI22X1 U253 ( .A0(n299), .A1(n434), .B0(n289), .B1(n433), .Y(n1157) );
  OAI22X1 U254 ( .A0(n298), .A1(n433), .B0(n287), .B1(n432), .Y(n1173) );
  OAI22X1 U255 ( .A0(n295), .A1(n428), .B0(n284), .B1(n427), .Y(n996) );
  OAI22X1 U256 ( .A0(n293), .A1(n427), .B0(n281), .B1(n426), .Y(n1012) );
  OAI22X1 U257 ( .A0(n292), .A1(n426), .B0(n282), .B1(n425), .Y(n1028) );
  OAI22X1 U258 ( .A0(n291), .A1(n425), .B0(n283), .B1(n424), .Y(n1044) );
  OAI22X1 U259 ( .A0(n301), .A1(n424), .B0(n284), .B1(n423), .Y(n1060) );
  OAI22X1 U260 ( .A0(n294), .A1(n423), .B0(n285), .B1(n422), .Y(n1076) );
  OAI22X1 U261 ( .A0(n295), .A1(n422), .B0(n286), .B1(n421), .Y(n1092) );
  OAI22X1 U262 ( .A0(n303), .A1(n421), .B0(n287), .B1(n420), .Y(n1108) );
  OAI22X1 U263 ( .A0(n301), .A1(n420), .B0(n288), .B1(n419), .Y(n1124) );
  OAI22X1 U264 ( .A0(n298), .A1(n419), .B0(n288), .B1(n418), .Y(n1140) );
  OAI22X1 U265 ( .A0(n300), .A1(n418), .B0(n289), .B1(n417), .Y(n1156) );
  OAI22X1 U266 ( .A0(n298), .A1(n417), .B0(n283), .B1(n416), .Y(n1172) );
  OAI22X1 U267 ( .A0(n295), .A1(n412), .B0(n280), .B1(n411), .Y(n995) );
  OAI22X1 U268 ( .A0(n293), .A1(n411), .B0(n281), .B1(n410), .Y(n1011) );
  OAI22X1 U269 ( .A0(n292), .A1(n410), .B0(n282), .B1(n409), .Y(n1027) );
  OAI22X1 U270 ( .A0(n291), .A1(n409), .B0(n283), .B1(n408), .Y(n1043) );
  OAI22X1 U271 ( .A0(n294), .A1(n395), .B0(n281), .B1(n394), .Y(n1010) );
  OAI22X1 U272 ( .A0(n292), .A1(n394), .B0(n282), .B1(n393), .Y(n1026) );
  OAI22X1 U273 ( .A0(n291), .A1(n393), .B0(n283), .B1(n392), .Y(n1042) );
  OAI22X1 U274 ( .A0(n294), .A1(n584), .B0(n284), .B1(n583), .Y(n1070) );
  OAI22X1 U275 ( .A0(n302), .A1(n583), .B0(n286), .B1(n582), .Y(n1086) );
  OAI22X1 U276 ( .A0(n303), .A1(n582), .B0(n287), .B1(n581), .Y(n1102) );
  OAI22X1 U277 ( .A0(n302), .A1(n581), .B0(n288), .B1(n580), .Y(n1118) );
  OAI22X1 U278 ( .A0(n293), .A1(n580), .B0(n288), .B1(n579), .Y(n1134) );
  OAI22X1 U279 ( .A0(n300), .A1(n472), .B0(n284), .B1(n471), .Y(n1063) );
  OAI22X1 U280 ( .A0(n299), .A1(n471), .B0(n285), .B1(n470), .Y(n1079) );
  OAI22X1 U281 ( .A0(n298), .A1(n470), .B0(n286), .B1(n469), .Y(n1095) );
  OAI22X1 U282 ( .A0(n302), .A1(n469), .B0(n287), .B1(n468), .Y(n1111) );
  OAI22X1 U283 ( .A0(n301), .A1(n468), .B0(n283), .B1(n467), .Y(n1127) );
  OAI22X1 U284 ( .A0(n299), .A1(n467), .B0(n285), .B1(n466), .Y(n1143) );
  OAI22X1 U285 ( .A0(n299), .A1(n466), .B0(n289), .B1(n465), .Y(n1159) );
  OAI22X1 U286 ( .A0(n298), .A1(n465), .B0(n288), .B1(n464), .Y(n1175) );
  OAI22X1 U287 ( .A0(n295), .A1(n460), .B0(n289), .B1(n459), .Y(n998) );
  OAI22X1 U288 ( .A0(n293), .A1(n459), .B0(n281), .B1(n458), .Y(n1014) );
  OAI22X1 U289 ( .A0(n292), .A1(n458), .B0(n282), .B1(n457), .Y(n1030) );
  OAI22X1 U290 ( .A0(n291), .A1(n457), .B0(n283), .B1(n456), .Y(n1046) );
  OAI22X1 U291 ( .A0(n296), .A1(n408), .B0(n288), .B1(n407), .Y(n1059) );
  OAI22X1 U292 ( .A0(n292), .A1(n407), .B0(n285), .B1(n406), .Y(n1075) );
  OAI22X1 U293 ( .A0(n296), .A1(n406), .B0(n286), .B1(n405), .Y(n1091) );
  OAI22X1 U294 ( .A0(n303), .A1(n405), .B0(n287), .B1(n404), .Y(n1107) );
  OAI22X1 U295 ( .A0(n301), .A1(n404), .B0(n288), .B1(n403), .Y(n1123) );
  OAI22X1 U296 ( .A0(n292), .A1(n403), .B0(n284), .B1(n402), .Y(n1139) );
  OAI22X1 U297 ( .A0(n300), .A1(n402), .B0(n289), .B1(n401), .Y(n1155) );
  OAI22X1 U298 ( .A0(n298), .A1(n401), .B0(n285), .B1(n400), .Y(n1171) );
  OAI22X1 U299 ( .A0(n295), .A1(n396), .B0(n280), .B1(n395), .Y(n994) );
  OAI22X1 U300 ( .A0(n290), .A1(n392), .B0(n284), .B1(n391), .Y(n1058) );
  OAI22X1 U301 ( .A0(n290), .A1(n391), .B0(n285), .B1(n390), .Y(n1074) );
  OAI22X1 U302 ( .A0(n299), .A1(n390), .B0(n286), .B1(n389), .Y(n1090) );
  OAI22X1 U303 ( .A0(n303), .A1(n389), .B0(n287), .B1(n388), .Y(n1106) );
  OAI22X1 U304 ( .A0(n301), .A1(n388), .B0(n288), .B1(n387), .Y(n1122) );
  OAI22X1 U305 ( .A0(n290), .A1(n387), .B0(n280), .B1(n386), .Y(n1138) );
  OAI22X1 U306 ( .A0(n300), .A1(n386), .B0(n289), .B1(n385), .Y(n1154) );
  OAI22X1 U307 ( .A0(n298), .A1(n385), .B0(n284), .B1(n384), .Y(n1170) );
  OAI22X1 U308 ( .A0(n295), .A1(n380), .B0(n280), .B1(n379), .Y(n993) );
  OAI22X1 U309 ( .A0(n294), .A1(n379), .B0(n281), .B1(n378), .Y(n1009) );
  OAI22X1 U310 ( .A0(n292), .A1(n378), .B0(n282), .B1(n377), .Y(n1025) );
  OAI22X1 U311 ( .A0(n291), .A1(n377), .B0(n283), .B1(n376), .Y(n1041) );
  OAI22X1 U312 ( .A0(n290), .A1(n376), .B0(n280), .B1(n375), .Y(n1057) );
  OAI22X1 U313 ( .A0(n291), .A1(n375), .B0(n285), .B1(n374), .Y(n1073) );
  OAI22X1 U314 ( .A0(n292), .A1(n374), .B0(n286), .B1(n373), .Y(n1089) );
  OAI22X1 U315 ( .A0(n303), .A1(n373), .B0(n287), .B1(n372), .Y(n1105) );
  OAI22X1 U316 ( .A0(n302), .A1(n372), .B0(n288), .B1(n371), .Y(n1121) );
  OAI22X1 U317 ( .A0(n297), .A1(n371), .B0(n286), .B1(n370), .Y(n1137) );
  OAI22X1 U318 ( .A0(n300), .A1(n370), .B0(n289), .B1(n369), .Y(n1153) );
  OAI22X1 U319 ( .A0(n298), .A1(n369), .B0(n280), .B1(n368), .Y(n1169) );
  OAI22X1 U320 ( .A0(n295), .A1(n364), .B0(n280), .B1(n363), .Y(n992) );
  OAI22X1 U321 ( .A0(n294), .A1(n363), .B0(n281), .B1(n362), .Y(n1008) );
  OAI22X1 U322 ( .A0(n292), .A1(n362), .B0(n282), .B1(n361), .Y(n1024) );
  OAI22X1 U323 ( .A0(n291), .A1(n361), .B0(n283), .B1(n360), .Y(n1040) );
  OAI22X1 U324 ( .A0(n290), .A1(n360), .B0(n289), .B1(n359), .Y(n1056) );
  OAI22X1 U325 ( .A0(n301), .A1(n359), .B0(n284), .B1(n358), .Y(n1072) );
  OAI22X1 U326 ( .A0(n291), .A1(n358), .B0(n286), .B1(n357), .Y(n1088) );
  OAI22X1 U327 ( .A0(n303), .A1(n357), .B0(n287), .B1(n356), .Y(n1104) );
  OAI22X1 U328 ( .A0(n302), .A1(n356), .B0(n288), .B1(n355), .Y(n1120) );
  OAI22X1 U329 ( .A0(n291), .A1(n355), .B0(n287), .B1(n354), .Y(n1136) );
  OAI22X1 U330 ( .A0(n300), .A1(n354), .B0(n289), .B1(n353), .Y(n1152) );
  OAI22X1 U331 ( .A0(n299), .A1(n353), .B0(n289), .B1(n352), .Y(n1168) );
  OAI22X1 U332 ( .A0(n295), .A1(n348), .B0(n280), .B1(n347), .Y(n991) );
  OAI22X1 U333 ( .A0(n294), .A1(n347), .B0(n279), .B1(n346), .Y(n1007) );
  OAI22X1 U334 ( .A0(n292), .A1(n346), .B0(n282), .B1(n345), .Y(n1023) );
  OAI22X1 U335 ( .A0(n291), .A1(n345), .B0(n283), .B1(n344), .Y(n1039) );
  OAI22X1 U336 ( .A0(n290), .A1(n344), .B0(n279), .B1(n343), .Y(n1055) );
  OAI22X1 U337 ( .A0(n303), .A1(n343), .B0(n284), .B1(n342), .Y(n1071) );
  OAI22X1 U338 ( .A0(n302), .A1(n342), .B0(n286), .B1(n341), .Y(n1087) );
  OAI22X1 U339 ( .A0(n303), .A1(n341), .B0(n287), .B1(n340), .Y(n1103) );
  OAI22X1 U340 ( .A0(n302), .A1(n340), .B0(n288), .B1(n339), .Y(n1119) );
  OAI22X1 U341 ( .A0(n294), .A1(n339), .B0(n285), .B1(n338), .Y(n1135) );
  OAI22X1 U342 ( .A0(n300), .A1(n338), .B0(n289), .B1(n337), .Y(n1151) );
  OAI22X1 U343 ( .A0(n299), .A1(n337), .B0(n279), .B1(n336), .Y(n1167) );
  OAI22X1 U344 ( .A0(n734), .A1(n696), .B0(n1267), .B1(n305), .Y(n940) );
  OAI22X1 U345 ( .A0(n734), .A1(n688), .B0(n1266), .B1(n307), .Y(n939) );
  OAI22X1 U346 ( .A0(n734), .A1(n680), .B0(n1265), .B1(n304), .Y(n938) );
  OAI22X1 U347 ( .A0(n734), .A1(n672), .B0(n1264), .B1(n307), .Y(n937) );
  OAI22X1 U348 ( .A0(n734), .A1(n664), .B0(n1263), .B1(n304), .Y(n936) );
  OAI22X1 U349 ( .A0(n311), .A1(n656), .B0(n1262), .B1(n305), .Y(n935) );
  OAI22X1 U350 ( .A0(n734), .A1(n648), .B0(n1261), .B1(n305), .Y(n934) );
  OAI22X1 U351 ( .A0(n308), .A1(n640), .B0(n1260), .B1(n304), .Y(n933) );
  OAI22X1 U352 ( .A0(n734), .A1(n632), .B0(n1259), .B1(n304), .Y(n932) );
  OAI22X1 U353 ( .A0(n731), .A1(n1247), .B0(n314), .B1(n1246), .Y(n766) );
  OAI22X1 U354 ( .A0(n315), .A1(n1246), .B0(n314), .B1(n1245), .Y(n782) );
  OAI22X1 U355 ( .A0(n316), .A1(n1245), .B0(n313), .B1(n1244), .Y(n798) );
  OAI22X1 U356 ( .A0(n316), .A1(n1244), .B0(n313), .B1(n1269), .Y(n814) );
  OAI22X1 U357 ( .A0(n731), .A1(n1243), .B0(n313), .B1(n1242), .Y(n765) );
  OAI22X1 U358 ( .A0(n315), .A1(n1242), .B0(n314), .B1(n1241), .Y(n781) );
  OAI22X1 U359 ( .A0(n731), .A1(n1241), .B0(n314), .B1(n1240), .Y(n797) );
  OAI22X1 U360 ( .A0(n731), .A1(n1240), .B0(n313), .B1(n1268), .Y(n813) );
  OAI22X1 U361 ( .A0(n731), .A1(n1239), .B0(n314), .B1(n1238), .Y(n764) );
  OAI22X1 U362 ( .A0(n315), .A1(n1238), .B0(n313), .B1(n1237), .Y(n780) );
  OAI22X1 U363 ( .A0(n731), .A1(n1237), .B0(n313), .B1(n1236), .Y(n796) );
  OAI22X1 U364 ( .A0(n315), .A1(n1236), .B0(n313), .B1(n1267), .Y(n812) );
  OAI22X1 U365 ( .A0(n731), .A1(n1235), .B0(n313), .B1(n1234), .Y(n763) );
  OAI22X1 U366 ( .A0(n315), .A1(n1234), .B0(n314), .B1(n1233), .Y(n779) );
  OAI22X1 U367 ( .A0(n731), .A1(n1233), .B0(n313), .B1(n1232), .Y(n795) );
  OAI22X1 U368 ( .A0(n316), .A1(n1232), .B0(n313), .B1(n1266), .Y(n811) );
  OAI22X1 U369 ( .A0(n316), .A1(n1231), .B0(n314), .B1(n1230), .Y(n762) );
  OAI22X1 U370 ( .A0(n315), .A1(n1230), .B0(n313), .B1(n1229), .Y(n778) );
  OAI22X1 U371 ( .A0(n731), .A1(n1229), .B0(n313), .B1(n1228), .Y(n794) );
  OAI22X1 U372 ( .A0(n316), .A1(n1228), .B0(n313), .B1(n1265), .Y(n810) );
  OAI22X1 U373 ( .A0(n315), .A1(n1227), .B0(n314), .B1(n1226), .Y(n761) );
  OAI22X1 U374 ( .A0(n315), .A1(n1226), .B0(n313), .B1(n1225), .Y(n777) );
  OAI22X1 U375 ( .A0(n731), .A1(n1225), .B0(n314), .B1(n1224), .Y(n793) );
  OAI22X1 U376 ( .A0(n316), .A1(n1224), .B0(n313), .B1(n1264), .Y(n809) );
  OAI22X1 U377 ( .A0(n316), .A1(n1223), .B0(n314), .B1(n1222), .Y(n760) );
  OAI22X1 U378 ( .A0(n315), .A1(n1222), .B0(n314), .B1(n1221), .Y(n776) );
  OAI22X1 U379 ( .A0(n731), .A1(n1221), .B0(n313), .B1(n1220), .Y(n792) );
  OAI22X1 U380 ( .A0(n316), .A1(n1220), .B0(n313), .B1(n1263), .Y(n808) );
  OAI22X1 U381 ( .A0(n315), .A1(n1219), .B0(n314), .B1(n1218), .Y(n759) );
  OAI22X1 U382 ( .A0(n731), .A1(n1218), .B0(n314), .B1(n1217), .Y(n775) );
  OAI22X1 U383 ( .A0(n731), .A1(n1217), .B0(n314), .B1(n1216), .Y(n791) );
  OAI22X1 U384 ( .A0(n316), .A1(n1216), .B0(n313), .B1(n1262), .Y(n807) );
  OAI22X1 U385 ( .A0(n315), .A1(n1215), .B0(n314), .B1(n1214), .Y(n758) );
  OAI22X1 U386 ( .A0(n731), .A1(n1214), .B0(n313), .B1(n1213), .Y(n774) );
  OAI22X1 U387 ( .A0(n731), .A1(n1213), .B0(n314), .B1(n1212), .Y(n790) );
  OAI22X1 U388 ( .A0(n316), .A1(n1212), .B0(n313), .B1(n1261), .Y(n806) );
  OAI22X1 U389 ( .A0(n315), .A1(n1211), .B0(n314), .B1(n1210), .Y(n757) );
  OAI22X1 U390 ( .A0(n731), .A1(n1210), .B0(n314), .B1(n1209), .Y(n773) );
  OAI22X1 U391 ( .A0(n731), .A1(n1209), .B0(n314), .B1(n1208), .Y(n789) );
  OAI22X1 U392 ( .A0(n316), .A1(n1208), .B0(n313), .B1(n1260), .Y(n805) );
  OAI22X1 U393 ( .A0(n731), .A1(n1207), .B0(n314), .B1(n1206), .Y(n756) );
  OAI22X1 U394 ( .A0(n731), .A1(n1206), .B0(n313), .B1(n1205), .Y(n772) );
  OAI22X1 U395 ( .A0(n731), .A1(n1205), .B0(n314), .B1(n1204), .Y(n788) );
  OAI22X1 U396 ( .A0(n316), .A1(n1204), .B0(n313), .B1(n1259), .Y(n804) );
  OAI22X1 U397 ( .A0(n731), .A1(n1203), .B0(n314), .B1(n1202), .Y(n755) );
  OAI22X1 U398 ( .A0(n731), .A1(n1202), .B0(n314), .B1(n1201), .Y(n771) );
  OAI22X1 U399 ( .A0(n731), .A1(n1201), .B0(n313), .B1(n1200), .Y(n787) );
  OAI22X1 U400 ( .A0(n316), .A1(n1200), .B0(n313), .B1(n1258), .Y(n803) );
  OAI22X1 U401 ( .A0(n731), .A1(n1199), .B0(n314), .B1(n739), .Y(n754) );
  OAI22X1 U402 ( .A0(n731), .A1(n739), .B0(n313), .B1(n738), .Y(n770) );
  OAI22X1 U403 ( .A0(n315), .A1(n738), .B0(n313), .B1(n735), .Y(n786) );
  OAI22X1 U404 ( .A0(n316), .A1(n735), .B0(n313), .B1(n1257), .Y(n802) );
  OAI22X1 U405 ( .A0(n731), .A1(n732), .B0(n314), .B1(n730), .Y(n753) );
  OAI22X1 U406 ( .A0(n731), .A1(n730), .B0(n314), .B1(n729), .Y(n769) );
  OAI22X1 U407 ( .A0(n315), .A1(n729), .B0(n313), .B1(n728), .Y(n785) );
  OAI22X1 U408 ( .A0(n316), .A1(n728), .B0(n314), .B1(n1256), .Y(n801) );
  OAI22X1 U409 ( .A0(n731), .A1(n727), .B0(n314), .B1(n726), .Y(n752) );
  OAI22X1 U410 ( .A0(n731), .A1(n726), .B0(n313), .B1(n725), .Y(n768) );
  OAI22X1 U411 ( .A0(n315), .A1(n725), .B0(n314), .B1(n724), .Y(n784) );
  OAI22X1 U412 ( .A0(n316), .A1(n724), .B0(n313), .B1(n1255), .Y(n800) );
  OAI22X1 U413 ( .A0(n731), .A1(n723), .B0(n314), .B1(n722), .Y(n751) );
  OAI22X1 U414 ( .A0(n311), .A1(n712), .B0(n1269), .B1(n306), .Y(n942) );
  OAI22X1 U415 ( .A0(n734), .A1(n704), .B0(n1268), .B1(n305), .Y(n941) );
  OAI22X1 U416 ( .A0(n722), .A1(n731), .B0(n314), .B1(n721), .Y(n767) );
  OAI22X1 U417 ( .A0(n315), .A1(n721), .B0(n314), .B1(n720), .Y(n783) );
  OAI22X1 U418 ( .A0(n316), .A1(n720), .B0(n313), .B1(n1254), .Y(n799) );
  OAI22X1 U419 ( .A0(n309), .A1(n719), .B0(n305), .B1(n718), .Y(n830) );
  OAI22X1 U420 ( .A0(n311), .A1(n718), .B0(n305), .B1(n717), .Y(n846) );
  OAI22X1 U421 ( .A0(n311), .A1(n717), .B0(n304), .B1(n716), .Y(n862) );
  OAI22X1 U422 ( .A0(n311), .A1(n711), .B0(n305), .B1(n710), .Y(n829) );
  OAI22X1 U423 ( .A0(n309), .A1(n710), .B0(n307), .B1(n709), .Y(n845) );
  OAI22X1 U424 ( .A0(n309), .A1(n709), .B0(n304), .B1(n708), .Y(n861) );
  OAI22X1 U425 ( .A0(n310), .A1(n703), .B0(n307), .B1(n702), .Y(n828) );
  OAI22X1 U426 ( .A0(n310), .A1(n702), .B0(n304), .B1(n701), .Y(n844) );
  OAI22X1 U427 ( .A0(n308), .A1(n701), .B0(n304), .B1(n700), .Y(n860) );
  OAI22X1 U428 ( .A0(n309), .A1(n695), .B0(n304), .B1(n694), .Y(n827) );
  OAI22X1 U429 ( .A0(n734), .A1(n694), .B0(n304), .B1(n693), .Y(n843) );
  OAI22X1 U430 ( .A0(n311), .A1(n693), .B0(n304), .B1(n692), .Y(n859) );
  OAI22X1 U431 ( .A0(n310), .A1(n687), .B0(n306), .B1(n686), .Y(n826) );
  OAI22X1 U432 ( .A0(n309), .A1(n686), .B0(n306), .B1(n685), .Y(n842) );
  OAI22X1 U433 ( .A0(n308), .A1(n685), .B0(n304), .B1(n684), .Y(n858) );
  OAI22X1 U434 ( .A0(n310), .A1(n679), .B0(n305), .B1(n678), .Y(n825) );
  OAI22X1 U435 ( .A0(n308), .A1(n678), .B0(n307), .B1(n677), .Y(n841) );
  OAI22X1 U436 ( .A0(n309), .A1(n677), .B0(n304), .B1(n676), .Y(n857) );
  OAI22X1 U437 ( .A0(n308), .A1(n671), .B0(n307), .B1(n670), .Y(n824) );
  OAI22X1 U438 ( .A0(n310), .A1(n670), .B0(n307), .B1(n669), .Y(n840) );
  OAI22X1 U439 ( .A0(n310), .A1(n669), .B0(n304), .B1(n668), .Y(n856) );
  OAI22X1 U440 ( .A0(n309), .A1(n663), .B0(n304), .B1(n662), .Y(n823) );
  OAI22X1 U441 ( .A0(n308), .A1(n662), .B0(n306), .B1(n661), .Y(n839) );
  OAI22X1 U442 ( .A0(n308), .A1(n661), .B0(n304), .B1(n660), .Y(n855) );
  OAI22X1 U443 ( .A0(n309), .A1(n655), .B0(n306), .B1(n654), .Y(n822) );
  OAI22X1 U444 ( .A0(n311), .A1(n654), .B0(n304), .B1(n653), .Y(n838) );
  OAI22X1 U445 ( .A0(n311), .A1(n653), .B0(n304), .B1(n652), .Y(n854) );
  OAI22X1 U446 ( .A0(n308), .A1(n647), .B0(n305), .B1(n646), .Y(n821) );
  OAI22X1 U447 ( .A0(n309), .A1(n646), .B0(n307), .B1(n645), .Y(n837) );
  OAI22X1 U448 ( .A0(n310), .A1(n645), .B0(n304), .B1(n644), .Y(n853) );
  OAI22X1 U449 ( .A0(n734), .A1(n639), .B0(n307), .B1(n638), .Y(n820) );
  OAI22X1 U450 ( .A0(n310), .A1(n638), .B0(n305), .B1(n637), .Y(n836) );
  OAI22X1 U451 ( .A0(n308), .A1(n637), .B0(n307), .B1(n636), .Y(n852) );
  OAI22X1 U452 ( .A0(n734), .A1(n631), .B0(n304), .B1(n630), .Y(n819) );
  OAI22X1 U453 ( .A0(n311), .A1(n630), .B0(n307), .B1(n629), .Y(n835) );
  OAI22X1 U454 ( .A0(n734), .A1(n629), .B0(n305), .B1(n628), .Y(n851) );
  OAI22X1 U455 ( .A0(n734), .A1(n623), .B0(n306), .B1(n622), .Y(n818) );
  OAI22X1 U456 ( .A0(n308), .A1(n622), .B0(n304), .B1(n621), .Y(n834) );
  OAI22X1 U457 ( .A0(n734), .A1(n621), .B0(n304), .B1(n620), .Y(n850) );
  OAI22X1 U458 ( .A0(n734), .A1(n615), .B0(n305), .B1(n614), .Y(n817) );
  OAI22X1 U459 ( .A0(n309), .A1(n614), .B0(n306), .B1(n613), .Y(n833) );
  OAI22X1 U460 ( .A0(n734), .A1(n613), .B0(n306), .B1(n612), .Y(n849) );
  OAI22X1 U461 ( .A0(n734), .A1(n607), .B0(n307), .B1(n606), .Y(n816) );
  OAI22X1 U462 ( .A0(n310), .A1(n606), .B0(n304), .B1(n605), .Y(n832) );
  OAI22X1 U463 ( .A0(n734), .A1(n605), .B0(n307), .B1(n604), .Y(n848) );
  OAI22X1 U464 ( .A0(n310), .A1(n599), .B0(n307), .B1(n598), .Y(n815) );
  OAI22X1 U465 ( .A0(n598), .A1(n734), .B0(n307), .B1(n597), .Y(n831) );
  OAI22X1 U466 ( .A0(n734), .A1(n597), .B0(n305), .B1(n596), .Y(n847) );
  OAI22X1 U467 ( .A0(n297), .A1(n591), .B0(n285), .B1(n590), .Y(n958) );
  OAI22X1 U468 ( .A0(n299), .A1(n590), .B0(n289), .B1(n589), .Y(n974) );
  OAI22X1 U469 ( .A0(n295), .A1(n589), .B0(n280), .B1(n588), .Y(n990) );
  OAI22X1 U470 ( .A0(n297), .A1(n575), .B0(n284), .B1(n574), .Y(n957) );
  OAI22X1 U471 ( .A0(n292), .A1(n574), .B0(n281), .B1(n573), .Y(n973) );
  OAI22X1 U472 ( .A0(n295), .A1(n573), .B0(n280), .B1(n572), .Y(n989) );
  OAI22X1 U473 ( .A0(n297), .A1(n559), .B0(n280), .B1(n558), .Y(n956) );
  OAI22X1 U474 ( .A0(n296), .A1(n558), .B0(n280), .B1(n557), .Y(n972) );
  OAI22X1 U475 ( .A0(n295), .A1(n557), .B0(n280), .B1(n556), .Y(n988) );
  OAI22X1 U476 ( .A0(n297), .A1(n543), .B0(n279), .B1(n542), .Y(n955) );
  OAI22X1 U477 ( .A0(n300), .A1(n542), .B0(n279), .B1(n541), .Y(n971) );
  OAI22X1 U478 ( .A0(n296), .A1(n541), .B0(n280), .B1(n540), .Y(n987) );
  OAI22X1 U479 ( .A0(n297), .A1(n527), .B0(n279), .B1(n526), .Y(n954) );
  OAI22X1 U480 ( .A0(n293), .A1(n526), .B0(n284), .B1(n525), .Y(n970) );
  OAI22X1 U481 ( .A0(n296), .A1(n525), .B0(n280), .B1(n524), .Y(n986) );
  OAI22X1 U482 ( .A0(n297), .A1(n511), .B0(n279), .B1(n510), .Y(n953) );
  OAI22X1 U483 ( .A0(n303), .A1(n510), .B0(n282), .B1(n509), .Y(n969) );
  OAI22X1 U484 ( .A0(n296), .A1(n509), .B0(n280), .B1(n508), .Y(n985) );
  OAI22X1 U485 ( .A0(n297), .A1(n495), .B0(n279), .B1(n494), .Y(n952) );
  OAI22X1 U486 ( .A0(n291), .A1(n494), .B0(n289), .B1(n493), .Y(n968) );
  OAI22X1 U487 ( .A0(n296), .A1(n493), .B0(n280), .B1(n492), .Y(n984) );
  OAI22X1 U488 ( .A0(n297), .A1(n479), .B0(n279), .B1(n478), .Y(n951) );
  OAI22X1 U489 ( .A0(n290), .A1(n478), .B0(n279), .B1(n477), .Y(n967) );
  OAI22X1 U490 ( .A0(n296), .A1(n477), .B0(n280), .B1(n476), .Y(n983) );
  OAI22X1 U491 ( .A0(n291), .A1(n463), .B0(n279), .B1(n462), .Y(n950) );
  OAI22X1 U492 ( .A0(n295), .A1(n462), .B0(n281), .B1(n461), .Y(n966) );
  OAI22X1 U493 ( .A0(n296), .A1(n461), .B0(n280), .B1(n460), .Y(n982) );
  OAI22X1 U494 ( .A0(n290), .A1(n447), .B0(n279), .B1(n446), .Y(n949) );
  OAI22X1 U495 ( .A0(n298), .A1(n446), .B0(n282), .B1(n445), .Y(n965) );
  OAI22X1 U496 ( .A0(n296), .A1(n445), .B0(n283), .B1(n444), .Y(n981) );
  OAI22X1 U497 ( .A0(n302), .A1(n431), .B0(n279), .B1(n430), .Y(n948) );
  OAI22X1 U498 ( .A0(n301), .A1(n430), .B0(n283), .B1(n429), .Y(n964) );
  OAI22X1 U499 ( .A0(n296), .A1(n429), .B0(n288), .B1(n428), .Y(n980) );
  OAI22X1 U500 ( .A0(n301), .A1(n415), .B0(n279), .B1(n414), .Y(n947) );
  OAI22X1 U501 ( .A0(n297), .A1(n414), .B0(n280), .B1(n413), .Y(n963) );
  OAI22X1 U502 ( .A0(n296), .A1(n413), .B0(n285), .B1(n412), .Y(n979) );
  OAI22X1 U503 ( .A0(n303), .A1(n399), .B0(n279), .B1(n398), .Y(n946) );
  OAI22X1 U504 ( .A0(n297), .A1(n398), .B0(n289), .B1(n397), .Y(n962) );
  OAI22X1 U505 ( .A0(n296), .A1(n397), .B0(n288), .B1(n396), .Y(n978) );
  OAI22X1 U506 ( .A0(n302), .A1(n383), .B0(n279), .B1(n382), .Y(n945) );
  OAI22X1 U507 ( .A0(n297), .A1(n382), .B0(n279), .B1(n381), .Y(n961) );
  OAI22X1 U508 ( .A0(n296), .A1(n381), .B0(n283), .B1(n380), .Y(n977) );
  OAI22X1 U509 ( .A0(n290), .A1(n367), .B0(n279), .B1(n366), .Y(n944) );
  OAI22X1 U510 ( .A0(n297), .A1(n366), .B0(n281), .B1(n365), .Y(n960) );
  OAI22X1 U511 ( .A0(n296), .A1(n365), .B0(n286), .B1(n364), .Y(n976) );
  OAI22X1 U512 ( .A0(n295), .A1(n351), .B0(n279), .B1(n350), .Y(n943) );
  OAI22X1 U513 ( .A0(n350), .A1(n297), .B0(n288), .B1(n349), .Y(n959) );
  OAI22X1 U514 ( .A0(n296), .A1(n349), .B0(n287), .B1(n348), .Y(n975) );
  OAI22X1 U515 ( .A0(n298), .A1(n576), .B0(n1269), .B1(n289), .Y(n1198) );
  OAI22X1 U516 ( .A0(n303), .A1(n560), .B0(n1268), .B1(n287), .Y(n1197) );
  OAI22X1 U517 ( .A0(n292), .A1(n544), .B0(n1267), .B1(n286), .Y(n1196) );
  OAI22X1 U518 ( .A0(n291), .A1(n528), .B0(n1266), .B1(n287), .Y(n1195) );
  OAI22X1 U519 ( .A0(n301), .A1(n512), .B0(n1265), .B1(n286), .Y(n1194) );
  OAI22X1 U520 ( .A0(n292), .A1(n496), .B0(n1264), .B1(n286), .Y(n1193) );
  OAI22X1 U521 ( .A0(n297), .A1(n480), .B0(n1263), .B1(n282), .Y(n1192) );
  OAI22X1 U522 ( .A0(n295), .A1(n464), .B0(n1262), .B1(n286), .Y(n1191) );
  OAI22X1 U523 ( .A0(n300), .A1(n448), .B0(n1261), .B1(n287), .Y(n1190) );
  NAND2X1 U524 ( .A(n737), .B(n1250), .Y(n734) );
  NOR2BX1 U525 ( .AN(N304), .B(n748), .Y(N1117) );
  NOR2BX1 U526 ( .AN(N303), .B(n748), .Y(N1116) );
  NOR2BX1 U527 ( .AN(N302), .B(n748), .Y(N1115) );
  INVX1 U528 ( .A(n736), .Y(n1250) );
  INVX1 U529 ( .A(n740), .Y(n1248) );
  NOR2X1 U530 ( .A(n744), .B(n1253), .Y(N1119) );
  AOI222X1 U531 ( .A0(n745), .A1(n733), .B0(n746), .B1(n740), .C0(n747), .C1(
        n736), .Y(n744) );
  INVX1 U532 ( .A(n733), .Y(n1251) );
  INVX1 U533 ( .A(n731), .Y(n317) );
  OAI222XL U534 ( .A0(n588), .A1(n275), .B0(n1244), .B1(n267), .C0(n716), .C1(
        n263), .Y(N224) );
  OAI222XL U535 ( .A0(n589), .A1(n277), .B0(n1245), .B1(n742), .C0(n717), .C1(
        n265), .Y(N241) );
  OAI222XL U536 ( .A0(n590), .A1(n277), .B0(n1246), .B1(n267), .C0(n718), .C1(
        n265), .Y(N257) );
  OAI222XL U537 ( .A0(n591), .A1(n276), .B0(n1247), .B1(n268), .C0(n719), .C1(
        n265), .Y(N273) );
  OAI222XL U538 ( .A0(n572), .A1(n275), .B0(n1240), .B1(n267), .C0(n708), .C1(
        n743), .Y(N225) );
  OAI222XL U539 ( .A0(n573), .A1(n277), .B0(n1241), .B1(n268), .C0(n709), .C1(
        n265), .Y(N242) );
  OAI222XL U540 ( .A0(n574), .A1(n277), .B0(n1242), .B1(n267), .C0(n710), .C1(
        n265), .Y(N258) );
  OAI222XL U541 ( .A0(n575), .A1(n276), .B0(n1243), .B1(n268), .C0(n711), .C1(
        n264), .Y(N274) );
  OAI222XL U542 ( .A0(n556), .A1(n275), .B0(n1236), .B1(n267), .C0(n700), .C1(
        n265), .Y(N226) );
  OAI222XL U543 ( .A0(n557), .A1(n277), .B0(n1237), .B1(n267), .C0(n701), .C1(
        n265), .Y(N243) );
  OAI222XL U544 ( .A0(n558), .A1(n276), .B0(n1238), .B1(n742), .C0(n702), .C1(
        n265), .Y(N259) );
  OAI222XL U545 ( .A0(n559), .A1(n276), .B0(n1239), .B1(n268), .C0(n703), .C1(
        n262), .Y(N275) );
  OAI222XL U546 ( .A0(n540), .A1(n275), .B0(n1232), .B1(n267), .C0(n692), .C1(
        n264), .Y(N227) );
  OAI222XL U547 ( .A0(n541), .A1(n277), .B0(n1233), .B1(n742), .C0(n693), .C1(
        n265), .Y(N244) );
  OAI222XL U548 ( .A0(n542), .A1(n276), .B0(n1234), .B1(n268), .C0(n694), .C1(
        n263), .Y(N260) );
  OAI222XL U549 ( .A0(n543), .A1(n276), .B0(n1235), .B1(n268), .C0(n695), .C1(
        n265), .Y(N276) );
  OAI222XL U550 ( .A0(n524), .A1(n275), .B0(n1228), .B1(n267), .C0(n684), .C1(
        n262), .Y(N228) );
  OAI222XL U551 ( .A0(n525), .A1(n277), .B0(n1229), .B1(n268), .C0(n685), .C1(
        n265), .Y(N245) );
  OAI222XL U552 ( .A0(n526), .A1(n276), .B0(n1230), .B1(n742), .C0(n686), .C1(
        n265), .Y(N261) );
  OAI222XL U553 ( .A0(n527), .A1(n276), .B0(n1231), .B1(n268), .C0(n687), .C1(
        n264), .Y(N277) );
  OAI222XL U554 ( .A0(n508), .A1(n275), .B0(n1224), .B1(n267), .C0(n676), .C1(
        n263), .Y(N229) );
  OAI222XL U555 ( .A0(n509), .A1(n277), .B0(n1225), .B1(n267), .C0(n677), .C1(
        n265), .Y(N246) );
  OAI222XL U556 ( .A0(n510), .A1(n276), .B0(n1226), .B1(n742), .C0(n678), .C1(
        n262), .Y(N262) );
  OAI222XL U557 ( .A0(n511), .A1(n276), .B0(n1227), .B1(n268), .C0(n679), .C1(
        n263), .Y(N278) );
  OAI222XL U558 ( .A0(n492), .A1(n275), .B0(n1220), .B1(n267), .C0(n668), .C1(
        n743), .Y(N231) );
  OAI222XL U559 ( .A0(n493), .A1(n277), .B0(n1221), .B1(n742), .C0(n669), .C1(
        n265), .Y(N247) );
  OAI222XL U560 ( .A0(n494), .A1(n276), .B0(n1222), .B1(n742), .C0(n670), .C1(
        n743), .Y(N263) );
  OAI222XL U561 ( .A0(n495), .A1(n276), .B0(n1223), .B1(n268), .C0(n671), .C1(
        n264), .Y(N279) );
  OAI222XL U562 ( .A0(n476), .A1(n275), .B0(n1216), .B1(n267), .C0(n660), .C1(
        n265), .Y(N232) );
  OAI222XL U563 ( .A0(n477), .A1(n277), .B0(n1217), .B1(n268), .C0(n661), .C1(
        n265), .Y(N248) );
  OAI222XL U564 ( .A0(n478), .A1(n276), .B0(n1218), .B1(n742), .C0(n662), .C1(
        n265), .Y(N264) );
  OAI222XL U565 ( .A0(n479), .A1(n276), .B0(n1219), .B1(n268), .C0(n663), .C1(
        n264), .Y(N280) );
  OAI222XL U566 ( .A0(n460), .A1(n275), .B0(n1212), .B1(n267), .C0(n652), .C1(
        n264), .Y(N233) );
  OAI222XL U567 ( .A0(n461), .A1(n277), .B0(n1213), .B1(n267), .C0(n653), .C1(
        n265), .Y(N249) );
  OAI222XL U568 ( .A0(n462), .A1(n275), .B0(n1214), .B1(n742), .C0(n654), .C1(
        n262), .Y(N265) );
  OAI222XL U569 ( .A0(n463), .A1(n276), .B0(n1215), .B1(n268), .C0(n655), .C1(
        n743), .Y(N281) );
  OAI222XL U570 ( .A0(n444), .A1(n275), .B0(n1208), .B1(n267), .C0(n644), .C1(
        n262), .Y(N234) );
  OAI222XL U571 ( .A0(n445), .A1(n277), .B0(n1209), .B1(n742), .C0(n645), .C1(
        n265), .Y(N250) );
  OAI222XL U572 ( .A0(n446), .A1(n276), .B0(n1210), .B1(n742), .C0(n646), .C1(
        n263), .Y(N266) );
  OAI222XL U573 ( .A0(n447), .A1(n275), .B0(n1211), .B1(n268), .C0(n647), .C1(
        n743), .Y(N282) );
  OAI222XL U574 ( .A0(n428), .A1(n275), .B0(n1204), .B1(n267), .C0(n636), .C1(
        n263), .Y(N235) );
  OAI222XL U575 ( .A0(n429), .A1(n277), .B0(n1205), .B1(n742), .C0(n637), .C1(
        n265), .Y(N251) );
  OAI222XL U576 ( .A0(n430), .A1(n276), .B0(n1206), .B1(n742), .C0(n638), .C1(
        n743), .Y(N267) );
  OAI222XL U577 ( .A0(n431), .A1(n275), .B0(n1207), .B1(n268), .C0(n639), .C1(
        n743), .Y(N283) );
  OAI222XL U578 ( .A0(n412), .A1(n275), .B0(n1200), .B1(n267), .C0(n628), .C1(
        n743), .Y(N236) );
  OAI222XL U579 ( .A0(n413), .A1(n277), .B0(n1201), .B1(n268), .C0(n629), .C1(
        n265), .Y(N252) );
  OAI222XL U580 ( .A0(n414), .A1(n276), .B0(n1202), .B1(n268), .C0(n630), .C1(
        n262), .Y(N268) );
  OAI222XL U581 ( .A0(n415), .A1(n275), .B0(n1203), .B1(n268), .C0(n631), .C1(
        n743), .Y(N284) );
  OAI222XL U582 ( .A0(n396), .A1(n277), .B0(n735), .B1(n267), .C0(n620), .C1(
        n265), .Y(N237) );
  OAI222XL U583 ( .A0(n397), .A1(n277), .B0(n738), .B1(n267), .C0(n621), .C1(
        n265), .Y(N253) );
  OAI222XL U584 ( .A0(n398), .A1(n276), .B0(n739), .B1(n267), .C0(n622), .C1(
        n265), .Y(N269) );
  OAI222XL U585 ( .A0(n399), .A1(n275), .B0(n1199), .B1(n742), .C0(n623), .C1(
        n743), .Y(N285) );
  OAI222XL U586 ( .A0(n380), .A1(n277), .B0(n728), .B1(n742), .C0(n612), .C1(
        n264), .Y(N238) );
  OAI222XL U587 ( .A0(n381), .A1(n277), .B0(n729), .B1(n268), .C0(n613), .C1(
        n265), .Y(N254) );
  OAI222XL U588 ( .A0(n382), .A1(n276), .B0(n730), .B1(n267), .C0(n614), .C1(
        n264), .Y(N270) );
  OAI222XL U589 ( .A0(n383), .A1(n275), .B0(n732), .B1(n742), .C0(n615), .C1(
        n743), .Y(N286) );
  OAI222XL U590 ( .A0(n364), .A1(n277), .B0(n724), .B1(n268), .C0(n604), .C1(
        n265), .Y(N239) );
  OAI222XL U591 ( .A0(n365), .A1(n277), .B0(n725), .B1(n742), .C0(n605), .C1(
        n265), .Y(N255) );
  OAI222XL U592 ( .A0(n366), .A1(n276), .B0(n726), .B1(n268), .C0(n606), .C1(
        n262), .Y(N271) );
  OAI222XL U593 ( .A0(n367), .A1(n275), .B0(n727), .B1(n742), .C0(n607), .C1(
        n743), .Y(N287) );
  OAI222XL U594 ( .A0(n348), .A1(n277), .B0(n720), .B1(n267), .C0(n596), .C1(
        n265), .Y(N240) );
  OAI222XL U595 ( .A0(n349), .A1(n277), .B0(n721), .B1(n268), .C0(n597), .C1(
        n265), .Y(N256) );
  OAI222XL U596 ( .A0(n350), .A1(n276), .B0(n722), .B1(n742), .C0(n598), .C1(
        n263), .Y(N272) );
  OAI222XL U597 ( .A0(n351), .A1(n275), .B0(n723), .B1(n742), .C0(n599), .C1(
        n743), .Y(N288) );
  OAI21XL U598 ( .A0(n333), .A1(n332), .B0(n335), .Y(N30) );
  OAI22X1 U599 ( .A0(n712), .A1(n262), .B0(n584), .B1(n271), .Y(N160) );
  OAI22X1 U600 ( .A0(n713), .A1(n263), .B0(n585), .B1(n274), .Y(N176) );
  OAI22X1 U601 ( .A0(n714), .A1(n263), .B0(n586), .B1(n741), .Y(N192) );
  OAI22X1 U602 ( .A0(n715), .A1(n264), .B0(n587), .B1(n271), .Y(N208) );
  OAI22X1 U603 ( .A0(n704), .A1(n262), .B0(n568), .B1(n277), .Y(N161) );
  OAI22X1 U604 ( .A0(n705), .A1(n263), .B0(n569), .B1(n270), .Y(N177) );
  OAI22X1 U605 ( .A0(n706), .A1(n743), .B0(n570), .B1(n274), .Y(N193) );
  OAI22X1 U606 ( .A0(n707), .A1(n264), .B0(n571), .B1(n271), .Y(N209) );
  OAI22X1 U607 ( .A0(n696), .A1(n262), .B0(n552), .B1(n275), .Y(N162) );
  OAI22X1 U608 ( .A0(n697), .A1(n263), .B0(n553), .B1(n275), .Y(N178) );
  OAI22X1 U609 ( .A0(n698), .A1(n264), .B0(n554), .B1(n273), .Y(N194) );
  OAI22X1 U610 ( .A0(n699), .A1(n264), .B0(n555), .B1(n271), .Y(N210) );
  OAI22X1 U611 ( .A0(n688), .A1(n262), .B0(n536), .B1(n741), .Y(N163) );
  OAI22X1 U612 ( .A0(n689), .A1(n263), .B0(n537), .B1(n741), .Y(N179) );
  OAI22X1 U613 ( .A0(n690), .A1(n262), .B0(n538), .B1(n274), .Y(N195) );
  OAI22X1 U614 ( .A0(n691), .A1(n264), .B0(n539), .B1(n270), .Y(N211) );
  OAI22X1 U615 ( .A0(n680), .A1(n262), .B0(n520), .B1(n276), .Y(N164) );
  OAI22X1 U616 ( .A0(n681), .A1(n263), .B0(n521), .B1(n273), .Y(N180) );
  OAI22X1 U617 ( .A0(n682), .A1(n743), .B0(n522), .B1(n272), .Y(N196) );
  OAI22X1 U618 ( .A0(n683), .A1(n264), .B0(n523), .B1(n270), .Y(N212) );
  OAI22X1 U619 ( .A0(n672), .A1(n262), .B0(n504), .B1(n272), .Y(N165) );
  OAI22X1 U620 ( .A0(n673), .A1(n263), .B0(n505), .B1(n272), .Y(N181) );
  OAI22X1 U621 ( .A0(n674), .A1(n743), .B0(n506), .B1(n277), .Y(N197) );
  OAI22X1 U622 ( .A0(n675), .A1(n264), .B0(n507), .B1(n270), .Y(N213) );
  OAI22X1 U623 ( .A0(n664), .A1(n262), .B0(n488), .B1(n272), .Y(N166) );
  OAI22X1 U624 ( .A0(n665), .A1(n263), .B0(n489), .B1(n271), .Y(N182) );
  OAI22X1 U625 ( .A0(n666), .A1(n743), .B0(n490), .B1(n271), .Y(N198) );
  OAI22X1 U626 ( .A0(n667), .A1(n264), .B0(n491), .B1(n270), .Y(N214) );
  OAI22X1 U627 ( .A0(n656), .A1(n262), .B0(n472), .B1(n277), .Y(N167) );
  OAI22X1 U628 ( .A0(n657), .A1(n263), .B0(n473), .B1(n277), .Y(N183) );
  OAI22X1 U629 ( .A0(n658), .A1(n743), .B0(n474), .B1(n271), .Y(N199) );
  OAI22X1 U630 ( .A0(n659), .A1(n264), .B0(n475), .B1(n270), .Y(N215) );
  OAI22X1 U631 ( .A0(n648), .A1(n262), .B0(n456), .B1(n276), .Y(N168) );
  OAI22X1 U632 ( .A0(n649), .A1(n263), .B0(n457), .B1(n276), .Y(N184) );
  OAI22X1 U633 ( .A0(n650), .A1(n743), .B0(n458), .B1(n271), .Y(N200) );
  OAI22X1 U634 ( .A0(n651), .A1(n264), .B0(n459), .B1(n270), .Y(N216) );
  OAI22X1 U635 ( .A0(n640), .A1(n262), .B0(n440), .B1(n274), .Y(N169) );
  OAI22X1 U636 ( .A0(n641), .A1(n743), .B0(n441), .B1(n270), .Y(N185) );
  OAI22X1 U637 ( .A0(n642), .A1(n743), .B0(n442), .B1(n271), .Y(N201) );
  OAI22X1 U638 ( .A0(n643), .A1(n264), .B0(n443), .B1(n270), .Y(N217) );
  OAI22X1 U639 ( .A0(n632), .A1(n262), .B0(n424), .B1(n273), .Y(N170) );
  OAI22X1 U640 ( .A0(n633), .A1(n743), .B0(n425), .B1(n270), .Y(N186) );
  OAI22X1 U641 ( .A0(n634), .A1(n264), .B0(n426), .B1(n271), .Y(N202) );
  OAI22X1 U642 ( .A0(n635), .A1(n264), .B0(n427), .B1(n270), .Y(N218) );
  OAI22X1 U643 ( .A0(n624), .A1(n262), .B0(n408), .B1(n270), .Y(N171) );
  OAI22X1 U644 ( .A0(n625), .A1(n264), .B0(n409), .B1(n271), .Y(N187) );
  OAI22X1 U645 ( .A0(n626), .A1(n262), .B0(n410), .B1(n271), .Y(N203) );
  OAI22X1 U646 ( .A0(n627), .A1(n264), .B0(n411), .B1(n270), .Y(N219) );
  OAI22X1 U647 ( .A0(n616), .A1(n263), .B0(n392), .B1(n274), .Y(N172) );
  OAI22X1 U648 ( .A0(n617), .A1(n262), .B0(n393), .B1(n276), .Y(N188) );
  OAI22X1 U649 ( .A0(n618), .A1(n263), .B0(n394), .B1(n271), .Y(N204) );
  OAI22X1 U650 ( .A0(n619), .A1(n264), .B0(n395), .B1(n270), .Y(N220) );
  OAI22X1 U651 ( .A0(n608), .A1(n263), .B0(n376), .B1(n270), .Y(N173) );
  OAI22X1 U652 ( .A0(n609), .A1(n263), .B0(n377), .B1(n741), .Y(N189) );
  OAI22X1 U653 ( .A0(n610), .A1(n262), .B0(n378), .B1(n271), .Y(N205) );
  OAI22X1 U654 ( .A0(n611), .A1(n262), .B0(n379), .B1(n270), .Y(N221) );
  OAI22X1 U655 ( .A0(n600), .A1(n263), .B0(n360), .B1(n275), .Y(N174) );
  OAI22X1 U656 ( .A0(n601), .A1(n265), .B0(n361), .B1(n274), .Y(N190) );
  OAI22X1 U657 ( .A0(n602), .A1(n743), .B0(n362), .B1(n271), .Y(N206) );
  OAI22X1 U658 ( .A0(n603), .A1(n263), .B0(n363), .B1(n270), .Y(N222) );
  OAI22X1 U659 ( .A0(n592), .A1(n263), .B0(n344), .B1(n741), .Y(N175) );
  OAI22X1 U660 ( .A0(n593), .A1(n743), .B0(n345), .B1(n273), .Y(N191) );
  OAI22X1 U661 ( .A0(n594), .A1(n264), .B0(n346), .B1(n271), .Y(N207) );
  OAI22X1 U662 ( .A0(n595), .A1(n743), .B0(n347), .B1(n270), .Y(N223) );
  NOR2X1 U663 ( .A(n576), .B(n272), .Y(N31) );
  NOR2X1 U664 ( .A(n577), .B(n272), .Y(N47) );
  NOR2X1 U665 ( .A(n578), .B(n273), .Y(N63) );
  NOR2X1 U666 ( .A(n579), .B(n270), .Y(N79) );
  NOR2X1 U667 ( .A(n580), .B(n270), .Y(N95) );
  NOR2X1 U668 ( .A(n581), .B(n277), .Y(N111) );
  NOR2X1 U669 ( .A(n582), .B(n274), .Y(N127) );
  NOR2X1 U670 ( .A(n583), .B(n741), .Y(N144) );
  NOR2X1 U671 ( .A(n560), .B(n741), .Y(N32) );
  NOR2X1 U672 ( .A(n561), .B(n272), .Y(N48) );
  NOR2X1 U673 ( .A(n562), .B(n273), .Y(N64) );
  NOR2X1 U674 ( .A(n563), .B(n275), .Y(N80) );
  NOR2X1 U675 ( .A(n564), .B(n271), .Y(N96) );
  NOR2X1 U676 ( .A(n565), .B(n272), .Y(N112) );
  NOR2X1 U677 ( .A(n566), .B(n274), .Y(N128) );
  NOR2X1 U678 ( .A(n567), .B(n741), .Y(N145) );
  NOR2X1 U679 ( .A(n544), .B(n273), .Y(N33) );
  NOR2X1 U680 ( .A(n545), .B(n272), .Y(N49) );
  NOR2X1 U681 ( .A(n546), .B(n273), .Y(N65) );
  NOR2X1 U682 ( .A(n547), .B(n741), .Y(N81) );
  NOR2X1 U683 ( .A(n548), .B(n272), .Y(N97) );
  NOR2X1 U684 ( .A(n549), .B(n271), .Y(N113) );
  NOR2X1 U685 ( .A(n550), .B(n274), .Y(N129) );
  NOR2X1 U686 ( .A(n551), .B(n741), .Y(N146) );
  NOR2X1 U687 ( .A(n528), .B(n272), .Y(N34) );
  NOR2X1 U688 ( .A(n529), .B(n272), .Y(N50) );
  NOR2X1 U689 ( .A(n530), .B(n273), .Y(N66) );
  NOR2X1 U690 ( .A(n531), .B(n273), .Y(N82) );
  NOR2X1 U691 ( .A(n532), .B(n277), .Y(N98) );
  NOR2X1 U692 ( .A(n533), .B(n271), .Y(N114) );
  NOR2X1 U693 ( .A(n534), .B(n274), .Y(N131) );
  NOR2X1 U694 ( .A(n535), .B(n741), .Y(N147) );
  NOR2X1 U695 ( .A(n512), .B(n276), .Y(N35) );
  NOR2X1 U696 ( .A(n513), .B(n272), .Y(N51) );
  NOR2X1 U697 ( .A(n514), .B(n273), .Y(N67) );
  NOR2X1 U698 ( .A(n515), .B(n274), .Y(N83) );
  NOR2X1 U699 ( .A(n516), .B(n274), .Y(N99) );
  NOR2X1 U700 ( .A(n517), .B(n274), .Y(N115) );
  NOR2X1 U701 ( .A(n518), .B(n273), .Y(N132) );
  NOR2X1 U702 ( .A(n519), .B(n741), .Y(N148) );
  NOR2X1 U703 ( .A(n496), .B(n270), .Y(N36) );
  NOR2X1 U704 ( .A(n497), .B(n272), .Y(N52) );
  NOR2X1 U705 ( .A(n498), .B(n273), .Y(N68) );
  NOR2X1 U706 ( .A(n499), .B(n271), .Y(N84) );
  NOR2X1 U707 ( .A(n500), .B(n275), .Y(N100) );
  NOR2X1 U708 ( .A(n501), .B(n274), .Y(N116) );
  NOR2X1 U709 ( .A(n502), .B(n273), .Y(N133) );
  NOR2X1 U710 ( .A(n503), .B(n275), .Y(N149) );
  NOR2X1 U711 ( .A(n480), .B(n741), .Y(N37) );
  NOR2X1 U712 ( .A(n481), .B(n272), .Y(N53) );
  NOR2X1 U713 ( .A(n482), .B(n276), .Y(N69) );
  NOR2X1 U714 ( .A(n483), .B(n741), .Y(N85) );
  NOR2X1 U715 ( .A(n484), .B(n272), .Y(N101) );
  NOR2X1 U716 ( .A(n485), .B(n274), .Y(N117) );
  NOR2X1 U717 ( .A(n486), .B(n271), .Y(N134) );
  NOR2X1 U718 ( .A(n487), .B(n741), .Y(N150) );
  NOR2X1 U719 ( .A(n464), .B(n273), .Y(N38) );
  NOR2X1 U720 ( .A(n465), .B(n272), .Y(N54) );
  NOR2X1 U721 ( .A(n466), .B(n274), .Y(N70) );
  NOR2X1 U722 ( .A(n467), .B(n274), .Y(N86) );
  NOR2X1 U723 ( .A(n468), .B(n275), .Y(N102) );
  NOR2X1 U724 ( .A(n469), .B(n274), .Y(N118) );
  NOR2X1 U725 ( .A(n470), .B(n271), .Y(N135) );
  NOR2X1 U726 ( .A(n471), .B(n741), .Y(N151) );
  NOR2X1 U727 ( .A(n448), .B(n272), .Y(N39) );
  NOR2X1 U728 ( .A(n449), .B(n273), .Y(N55) );
  NOR2X1 U729 ( .A(n450), .B(n273), .Y(N71) );
  NOR2X1 U730 ( .A(n451), .B(n273), .Y(N87) );
  NOR2X1 U731 ( .A(n452), .B(n270), .Y(N103) );
  NOR2X1 U732 ( .A(n453), .B(n274), .Y(N119) );
  NOR2X1 U733 ( .A(n454), .B(n741), .Y(N136) );
  NOR2X1 U734 ( .A(n455), .B(n741), .Y(N152) );
  NOR2X1 U735 ( .A(n432), .B(n271), .Y(N40) );
  NOR2X1 U736 ( .A(n433), .B(n273), .Y(N56) );
  NOR2X1 U737 ( .A(n434), .B(n272), .Y(N72) );
  NOR2X1 U738 ( .A(n435), .B(n273), .Y(N88) );
  NOR2X1 U739 ( .A(n436), .B(n271), .Y(N104) );
  NOR2X1 U740 ( .A(n437), .B(n274), .Y(N120) );
  NOR2X1 U741 ( .A(n438), .B(n274), .Y(N137) );
  NOR2X1 U742 ( .A(n439), .B(n741), .Y(N153) );
  NOR2X1 U743 ( .A(n416), .B(n272), .Y(N41) );
  NOR2X1 U744 ( .A(n417), .B(n273), .Y(N57) );
  NOR2X1 U745 ( .A(n418), .B(n271), .Y(N73) );
  NOR2X1 U746 ( .A(n419), .B(n272), .Y(N89) );
  NOR2X1 U747 ( .A(n420), .B(n275), .Y(N105) );
  NOR2X1 U748 ( .A(n421), .B(n274), .Y(N121) );
  NOR2X1 U749 ( .A(n422), .B(n270), .Y(N138) );
  NOR2X1 U750 ( .A(n423), .B(n741), .Y(N154) );
  NOR2X1 U751 ( .A(n400), .B(n272), .Y(N42) );
  NOR2X1 U752 ( .A(n401), .B(n273), .Y(N58) );
  NOR2X1 U753 ( .A(n402), .B(n277), .Y(N74) );
  NOR2X1 U754 ( .A(n403), .B(n273), .Y(N90) );
  NOR2X1 U755 ( .A(n404), .B(n272), .Y(N106) );
  NOR2X1 U756 ( .A(n405), .B(n274), .Y(N122) );
  NOR2X1 U757 ( .A(n406), .B(n271), .Y(N139) );
  NOR2X1 U758 ( .A(n407), .B(n741), .Y(N155) );
  NOR2X1 U759 ( .A(n384), .B(n272), .Y(N43) );
  NOR2X1 U760 ( .A(n385), .B(n273), .Y(N59) );
  NOR2X1 U761 ( .A(n386), .B(n277), .Y(N75) );
  NOR2X1 U762 ( .A(n387), .B(n276), .Y(N91) );
  NOR2X1 U763 ( .A(n388), .B(n741), .Y(N107) );
  NOR2X1 U764 ( .A(n389), .B(n274), .Y(N123) );
  NOR2X1 U765 ( .A(n390), .B(n741), .Y(N140) );
  NOR2X1 U766 ( .A(n391), .B(n741), .Y(N156) );
  NOR2X1 U767 ( .A(n368), .B(n272), .Y(N44) );
  NOR2X1 U768 ( .A(n369), .B(n273), .Y(N60) );
  NOR2X1 U769 ( .A(n370), .B(n270), .Y(N76) );
  NOR2X1 U770 ( .A(n371), .B(n270), .Y(N92) );
  NOR2X1 U771 ( .A(n372), .B(n274), .Y(N108) );
  NOR2X1 U772 ( .A(n373), .B(n274), .Y(N124) );
  NOR2X1 U773 ( .A(n374), .B(n276), .Y(N141) );
  NOR2X1 U774 ( .A(n375), .B(n741), .Y(N157) );
  NOR2X1 U775 ( .A(n352), .B(n272), .Y(N45) );
  NOR2X1 U776 ( .A(n353), .B(n273), .Y(N61) );
  NOR2X1 U777 ( .A(n354), .B(n275), .Y(N77) );
  NOR2X1 U778 ( .A(n355), .B(n271), .Y(N93) );
  NOR2X1 U779 ( .A(n356), .B(n273), .Y(N109) );
  NOR2X1 U780 ( .A(n357), .B(n270), .Y(N125) );
  NOR2X1 U781 ( .A(n358), .B(n741), .Y(N142) );
  NOR2X1 U782 ( .A(n359), .B(n275), .Y(N158) );
  NOR2X1 U783 ( .A(n336), .B(n272), .Y(N46) );
  NOR2X1 U784 ( .A(n337), .B(n273), .Y(N62) );
  NOR2X1 U785 ( .A(n338), .B(n741), .Y(N78) );
  NOR2X1 U786 ( .A(n339), .B(n270), .Y(N94) );
  NOR2X1 U787 ( .A(n340), .B(n272), .Y(N110) );
  NOR2X1 U788 ( .A(n341), .B(n274), .Y(N126) );
  NOR2X1 U789 ( .A(n342), .B(n274), .Y(N143) );
  NOR2X1 U790 ( .A(n343), .B(n741), .Y(N159) );
  NAND2X1 U791 ( .A(n333), .B(n332), .Y(n742) );
  INVX1 U792 ( .A(n741), .Y(n278) );
  INVX1 U793 ( .A(n743), .Y(n266) );
  OAI211X1 U794 ( .A0(n1252), .A1(n1249), .B0(n1251), .C0(start), .Y(n731) );
  NAND2X1 U795 ( .A(start), .B(n749), .Y(n748) );
  OAI222XL U796 ( .A0(n747), .A1(n1250), .B0(n746), .B1(n1248), .C0(n745), 
        .C1(n1251), .Y(n749) );
  NOR2X1 U797 ( .A(mode[0]), .B(mode[1]), .Y(n733) );
  NOR2X1 U798 ( .A(n1252), .B(mode[1]), .Y(n736) );
  NOR2X1 U799 ( .A(n1249), .B(mode[0]), .Y(n740) );
  AOI21X1 U800 ( .A0(mode[0]), .A1(mode[1]), .B0(n1253), .Y(n737) );
  NOR2X1 U801 ( .A(n5), .B(n748), .Y(N1118) );
  XNOR2X1 U802 ( .A(r71_carry[4]), .B(count[4]), .Y(n5) );
  NOR2X1 U803 ( .A(count[0]), .B(n748), .Y(N1114) );
  INVX1 U804 ( .A(start), .Y(n1253) );
  INVX1 U805 ( .A(mode[0]), .Y(n1252) );
  INVX1 U806 ( .A(mode[1]), .Y(n1249) );
  INVX1 U807 ( .A(s2p_ready), .Y(n335) );
  INVX1 U808 ( .A(din[0]), .Y(n1269) );
  INVX1 U809 ( .A(din[1]), .Y(n1268) );
  INVX1 U810 ( .A(din[2]), .Y(n1267) );
  INVX1 U811 ( .A(din[3]), .Y(n1266) );
  INVX1 U812 ( .A(din[4]), .Y(n1265) );
  INVX1 U813 ( .A(din[5]), .Y(n1264) );
  INVX1 U814 ( .A(din[6]), .Y(n1263) );
  INVX1 U815 ( .A(din[7]), .Y(n1262) );
  INVX1 U816 ( .A(din[8]), .Y(n1261) );
  INVX1 U817 ( .A(din[9]), .Y(n1260) );
  INVX1 U818 ( .A(din[10]), .Y(n1259) );
  INVX1 U819 ( .A(din[11]), .Y(n1258) );
  INVX1 U820 ( .A(din[12]), .Y(n1257) );
  INVX1 U821 ( .A(din[13]), .Y(n1256) );
  INVX1 U822 ( .A(din[14]), .Y(n1255) );
  INVX1 U823 ( .A(din[15]), .Y(n1254) );
  INVX1 U824 ( .A(mode_reg[0]), .Y(n333) );
  INVX1 U825 ( .A(mode_reg[1]), .Y(n332) );
  NAND3BX1 U826 ( .AN(count[4]), .B(count[0]), .C(count[1]), .Y(n750) );
  NOR3X1 U827 ( .A(count[2]), .B(count[3]), .C(n750), .Y(n745) );
  NOR3X1 U828 ( .A(n750), .B(count[3]), .C(n334), .Y(n747) );
  NOR3BX1 U829 ( .AN(count[3]), .B(n334), .C(n750), .Y(n746) );
  INVX1 U830 ( .A(dout16_reg[176]), .Y(n587) );
  INVX1 U831 ( .A(dout16_reg[160]), .Y(n586) );
  INVX1 U832 ( .A(dout16_reg[144]), .Y(n585) );
  INVX1 U833 ( .A(dout16_reg[128]), .Y(n584) );
  INVX1 U834 ( .A(dout16_reg[177]), .Y(n571) );
  INVX1 U835 ( .A(dout16_reg[161]), .Y(n570) );
  INVX1 U836 ( .A(dout16_reg[145]), .Y(n569) );
  INVX1 U837 ( .A(dout16_reg[129]), .Y(n568) );
  INVX1 U838 ( .A(dout16_reg[178]), .Y(n555) );
  INVX1 U839 ( .A(dout16_reg[162]), .Y(n554) );
  INVX1 U840 ( .A(dout16_reg[146]), .Y(n553) );
  INVX1 U841 ( .A(dout16_reg[130]), .Y(n552) );
  INVX1 U842 ( .A(dout16_reg[179]), .Y(n539) );
  INVX1 U843 ( .A(dout16_reg[163]), .Y(n538) );
  INVX1 U844 ( .A(dout16_reg[147]), .Y(n537) );
  INVX1 U845 ( .A(dout16_reg[131]), .Y(n536) );
  INVX1 U846 ( .A(dout16_reg[180]), .Y(n523) );
  INVX1 U847 ( .A(dout16_reg[164]), .Y(n522) );
  INVX1 U848 ( .A(dout16_reg[148]), .Y(n521) );
  INVX1 U849 ( .A(dout16_reg[132]), .Y(n520) );
  INVX1 U850 ( .A(dout16_reg[181]), .Y(n507) );
  INVX1 U851 ( .A(dout16_reg[165]), .Y(n506) );
  INVX1 U852 ( .A(dout16_reg[149]), .Y(n505) );
  INVX1 U853 ( .A(dout16_reg[133]), .Y(n504) );
  INVX1 U854 ( .A(dout16_reg[182]), .Y(n491) );
  INVX1 U855 ( .A(dout16_reg[166]), .Y(n490) );
  INVX1 U856 ( .A(dout16_reg[150]), .Y(n489) );
  INVX1 U857 ( .A(dout16_reg[134]), .Y(n488) );
  INVX1 U858 ( .A(dout16_reg[183]), .Y(n475) );
  INVX1 U859 ( .A(dout16_reg[167]), .Y(n474) );
  INVX1 U860 ( .A(dout16_reg[151]), .Y(n473) );
  INVX1 U861 ( .A(dout16_reg[135]), .Y(n472) );
  INVX1 U862 ( .A(dout16_reg[184]), .Y(n459) );
  INVX1 U863 ( .A(dout16_reg[168]), .Y(n458) );
  INVX1 U864 ( .A(dout16_reg[152]), .Y(n457) );
  INVX1 U865 ( .A(dout16_reg[136]), .Y(n456) );
  INVX1 U866 ( .A(dout16_reg[185]), .Y(n443) );
  INVX1 U867 ( .A(dout16_reg[169]), .Y(n442) );
  INVX1 U868 ( .A(dout16_reg[153]), .Y(n441) );
  INVX1 U869 ( .A(dout16_reg[137]), .Y(n440) );
  INVX1 U870 ( .A(dout16_reg[186]), .Y(n427) );
  INVX1 U871 ( .A(dout16_reg[170]), .Y(n426) );
  INVX1 U872 ( .A(dout16_reg[154]), .Y(n425) );
  INVX1 U873 ( .A(dout16_reg[138]), .Y(n424) );
  INVX1 U874 ( .A(dout16_reg[187]), .Y(n411) );
  INVX1 U875 ( .A(dout16_reg[171]), .Y(n410) );
  INVX1 U876 ( .A(dout16_reg[155]), .Y(n409) );
  INVX1 U877 ( .A(dout16_reg[139]), .Y(n408) );
  INVX1 U878 ( .A(dout16_reg[188]), .Y(n395) );
  INVX1 U879 ( .A(dout16_reg[172]), .Y(n394) );
  INVX1 U880 ( .A(dout16_reg[156]), .Y(n393) );
  INVX1 U881 ( .A(dout16_reg[140]), .Y(n392) );
  INVX1 U882 ( .A(dout16_reg[189]), .Y(n379) );
  INVX1 U883 ( .A(dout16_reg[173]), .Y(n378) );
  INVX1 U884 ( .A(dout16_reg[157]), .Y(n377) );
  INVX1 U885 ( .A(dout16_reg[141]), .Y(n376) );
  INVX1 U886 ( .A(dout16_reg[190]), .Y(n363) );
  INVX1 U887 ( .A(dout16_reg[174]), .Y(n362) );
  INVX1 U888 ( .A(dout16_reg[158]), .Y(n361) );
  INVX1 U889 ( .A(dout16_reg[142]), .Y(n360) );
  INVX1 U890 ( .A(dout16_reg[191]), .Y(n347) );
  INVX1 U891 ( .A(dout16_reg[175]), .Y(n346) );
  INVX1 U892 ( .A(dout16_reg[159]), .Y(n345) );
  INVX1 U893 ( .A(dout16_reg[143]), .Y(n344) );
  INVX1 U894 ( .A(dout8_reg[48]), .Y(n715) );
  INVX1 U895 ( .A(dout8_reg[32]), .Y(n714) );
  INVX1 U896 ( .A(dout8_reg[16]), .Y(n713) );
  INVX1 U897 ( .A(dout8_reg[0]), .Y(n712) );
  INVX1 U898 ( .A(dout8_reg[49]), .Y(n707) );
  INVX1 U899 ( .A(dout8_reg[33]), .Y(n706) );
  INVX1 U900 ( .A(dout8_reg[17]), .Y(n705) );
  INVX1 U901 ( .A(dout8_reg[1]), .Y(n704) );
  INVX1 U902 ( .A(dout8_reg[50]), .Y(n699) );
  INVX1 U903 ( .A(dout8_reg[34]), .Y(n698) );
  INVX1 U904 ( .A(dout8_reg[18]), .Y(n697) );
  INVX1 U905 ( .A(dout8_reg[2]), .Y(n696) );
  INVX1 U906 ( .A(dout8_reg[51]), .Y(n691) );
  INVX1 U907 ( .A(dout8_reg[35]), .Y(n690) );
  INVX1 U908 ( .A(dout8_reg[19]), .Y(n689) );
  INVX1 U909 ( .A(dout8_reg[3]), .Y(n688) );
  INVX1 U910 ( .A(dout8_reg[52]), .Y(n683) );
  INVX1 U911 ( .A(dout8_reg[36]), .Y(n682) );
  INVX1 U912 ( .A(dout8_reg[20]), .Y(n681) );
  INVX1 U913 ( .A(dout8_reg[4]), .Y(n680) );
  INVX1 U914 ( .A(dout8_reg[53]), .Y(n675) );
  INVX1 U915 ( .A(dout8_reg[37]), .Y(n674) );
  INVX1 U916 ( .A(dout8_reg[21]), .Y(n673) );
  INVX1 U917 ( .A(dout8_reg[5]), .Y(n672) );
  INVX1 U918 ( .A(dout8_reg[54]), .Y(n667) );
  INVX1 U919 ( .A(dout8_reg[38]), .Y(n666) );
  INVX1 U920 ( .A(dout8_reg[22]), .Y(n665) );
  INVX1 U921 ( .A(dout8_reg[6]), .Y(n664) );
  INVX1 U922 ( .A(dout8_reg[55]), .Y(n659) );
  INVX1 U923 ( .A(dout8_reg[39]), .Y(n658) );
  INVX1 U924 ( .A(dout8_reg[23]), .Y(n657) );
  INVX1 U925 ( .A(dout8_reg[7]), .Y(n656) );
  INVX1 U926 ( .A(dout8_reg[56]), .Y(n651) );
  INVX1 U927 ( .A(dout8_reg[40]), .Y(n650) );
  INVX1 U928 ( .A(dout8_reg[24]), .Y(n649) );
  INVX1 U929 ( .A(dout8_reg[8]), .Y(n648) );
  INVX1 U930 ( .A(dout8_reg[57]), .Y(n643) );
  INVX1 U931 ( .A(dout8_reg[41]), .Y(n642) );
  INVX1 U932 ( .A(dout8_reg[25]), .Y(n641) );
  INVX1 U933 ( .A(dout8_reg[9]), .Y(n640) );
  INVX1 U934 ( .A(dout8_reg[58]), .Y(n635) );
  INVX1 U935 ( .A(dout8_reg[42]), .Y(n634) );
  INVX1 U936 ( .A(dout8_reg[26]), .Y(n633) );
  INVX1 U937 ( .A(dout8_reg[10]), .Y(n632) );
  INVX1 U938 ( .A(dout8_reg[59]), .Y(n627) );
  INVX1 U939 ( .A(dout8_reg[43]), .Y(n626) );
  INVX1 U940 ( .A(dout8_reg[27]), .Y(n625) );
  INVX1 U941 ( .A(dout8_reg[11]), .Y(n624) );
  INVX1 U942 ( .A(dout8_reg[60]), .Y(n619) );
  INVX1 U943 ( .A(dout8_reg[44]), .Y(n618) );
  INVX1 U944 ( .A(dout8_reg[28]), .Y(n617) );
  INVX1 U945 ( .A(dout8_reg[12]), .Y(n616) );
  INVX1 U946 ( .A(dout8_reg[61]), .Y(n611) );
  INVX1 U947 ( .A(dout8_reg[45]), .Y(n610) );
  INVX1 U948 ( .A(dout8_reg[29]), .Y(n609) );
  INVX1 U949 ( .A(dout8_reg[13]), .Y(n608) );
  INVX1 U950 ( .A(dout8_reg[62]), .Y(n603) );
  INVX1 U951 ( .A(dout8_reg[46]), .Y(n602) );
  INVX1 U952 ( .A(dout8_reg[30]), .Y(n601) );
  INVX1 U953 ( .A(dout8_reg[14]), .Y(n600) );
  INVX1 U954 ( .A(dout8_reg[63]), .Y(n595) );
  INVX1 U955 ( .A(dout8_reg[47]), .Y(n594) );
  INVX1 U956 ( .A(dout8_reg[31]), .Y(n593) );
  INVX1 U957 ( .A(dout8_reg[15]), .Y(n592) );
  INVX1 U958 ( .A(dout16_reg[112]), .Y(n583) );
  INVX1 U959 ( .A(dout16_reg[96]), .Y(n582) );
  INVX1 U960 ( .A(dout16_reg[80]), .Y(n581) );
  INVX1 U961 ( .A(dout16_reg[64]), .Y(n580) );
  INVX1 U962 ( .A(dout16_reg[48]), .Y(n579) );
  INVX1 U963 ( .A(dout16_reg[32]), .Y(n578) );
  INVX1 U964 ( .A(dout16_reg[16]), .Y(n577) );
  INVX1 U965 ( .A(dout16_reg[0]), .Y(n576) );
  INVX1 U966 ( .A(dout16_reg[113]), .Y(n567) );
  INVX1 U967 ( .A(dout16_reg[97]), .Y(n566) );
  INVX1 U968 ( .A(dout16_reg[81]), .Y(n565) );
  INVX1 U969 ( .A(dout16_reg[65]), .Y(n564) );
  INVX1 U970 ( .A(dout16_reg[49]), .Y(n563) );
  INVX1 U971 ( .A(dout16_reg[33]), .Y(n562) );
  INVX1 U972 ( .A(dout16_reg[17]), .Y(n561) );
  INVX1 U973 ( .A(dout16_reg[1]), .Y(n560) );
  INVX1 U974 ( .A(dout16_reg[114]), .Y(n551) );
  INVX1 U975 ( .A(dout16_reg[98]), .Y(n550) );
  INVX1 U976 ( .A(dout16_reg[82]), .Y(n549) );
  INVX1 U977 ( .A(dout16_reg[66]), .Y(n548) );
  INVX1 U978 ( .A(dout16_reg[50]), .Y(n547) );
  INVX1 U979 ( .A(dout16_reg[34]), .Y(n546) );
  INVX1 U980 ( .A(dout16_reg[18]), .Y(n545) );
  INVX1 U981 ( .A(dout16_reg[2]), .Y(n544) );
  INVX1 U982 ( .A(dout16_reg[115]), .Y(n535) );
  INVX1 U983 ( .A(dout16_reg[99]), .Y(n534) );
  INVX1 U984 ( .A(dout16_reg[83]), .Y(n533) );
  INVX1 U985 ( .A(dout16_reg[67]), .Y(n532) );
  INVX1 U986 ( .A(dout16_reg[51]), .Y(n531) );
  INVX1 U987 ( .A(dout16_reg[35]), .Y(n530) );
  INVX1 U988 ( .A(dout16_reg[19]), .Y(n529) );
  INVX1 U989 ( .A(dout16_reg[3]), .Y(n528) );
  INVX1 U990 ( .A(dout16_reg[116]), .Y(n519) );
  INVX1 U991 ( .A(dout16_reg[100]), .Y(n518) );
  INVX1 U992 ( .A(dout16_reg[84]), .Y(n517) );
  INVX1 U993 ( .A(dout16_reg[68]), .Y(n516) );
  INVX1 U994 ( .A(dout16_reg[52]), .Y(n515) );
  INVX1 U995 ( .A(dout16_reg[36]), .Y(n514) );
  INVX1 U996 ( .A(dout16_reg[20]), .Y(n513) );
  INVX1 U997 ( .A(dout16_reg[4]), .Y(n512) );
  INVX1 U998 ( .A(dout16_reg[117]), .Y(n503) );
  INVX1 U999 ( .A(dout16_reg[101]), .Y(n502) );
  INVX1 U1000 ( .A(dout16_reg[85]), .Y(n501) );
  INVX1 U1001 ( .A(dout16_reg[69]), .Y(n500) );
  INVX1 U1002 ( .A(dout16_reg[53]), .Y(n499) );
  INVX1 U1003 ( .A(dout16_reg[37]), .Y(n498) );
  INVX1 U1004 ( .A(dout16_reg[21]), .Y(n497) );
  INVX1 U1005 ( .A(dout16_reg[5]), .Y(n496) );
  INVX1 U1006 ( .A(dout16_reg[118]), .Y(n487) );
  INVX1 U1007 ( .A(dout16_reg[102]), .Y(n486) );
  INVX1 U1008 ( .A(dout16_reg[86]), .Y(n485) );
  INVX1 U1009 ( .A(dout16_reg[70]), .Y(n484) );
  INVX1 U1010 ( .A(dout16_reg[54]), .Y(n483) );
  INVX1 U1011 ( .A(dout16_reg[38]), .Y(n482) );
  INVX1 U1012 ( .A(dout16_reg[22]), .Y(n481) );
  INVX1 U1013 ( .A(dout16_reg[6]), .Y(n480) );
  INVX1 U1014 ( .A(dout16_reg[119]), .Y(n471) );
  INVX1 U1015 ( .A(dout16_reg[103]), .Y(n470) );
  INVX1 U1016 ( .A(dout16_reg[87]), .Y(n469) );
  INVX1 U1017 ( .A(dout16_reg[71]), .Y(n468) );
  INVX1 U1018 ( .A(dout16_reg[55]), .Y(n467) );
  INVX1 U1019 ( .A(dout16_reg[39]), .Y(n466) );
  INVX1 U1020 ( .A(dout16_reg[23]), .Y(n465) );
  INVX1 U1021 ( .A(dout16_reg[7]), .Y(n464) );
  INVX1 U1022 ( .A(dout16_reg[120]), .Y(n455) );
  INVX1 U1023 ( .A(dout16_reg[104]), .Y(n454) );
  INVX1 U1024 ( .A(dout16_reg[88]), .Y(n453) );
  INVX1 U1025 ( .A(dout16_reg[72]), .Y(n452) );
  INVX1 U1026 ( .A(dout16_reg[56]), .Y(n451) );
  INVX1 U1027 ( .A(dout16_reg[40]), .Y(n450) );
  INVX1 U1028 ( .A(dout16_reg[24]), .Y(n449) );
  INVX1 U1029 ( .A(dout16_reg[8]), .Y(n448) );
  INVX1 U1030 ( .A(dout16_reg[121]), .Y(n439) );
  INVX1 U1031 ( .A(dout16_reg[105]), .Y(n438) );
  INVX1 U1032 ( .A(dout16_reg[89]), .Y(n437) );
  INVX1 U1033 ( .A(dout16_reg[73]), .Y(n436) );
  INVX1 U1034 ( .A(dout16_reg[57]), .Y(n435) );
  INVX1 U1035 ( .A(dout16_reg[41]), .Y(n434) );
  INVX1 U1036 ( .A(dout16_reg[25]), .Y(n433) );
  INVX1 U1037 ( .A(dout16_reg[9]), .Y(n432) );
  INVX1 U1038 ( .A(dout16_reg[122]), .Y(n423) );
  INVX1 U1039 ( .A(dout16_reg[106]), .Y(n422) );
  INVX1 U1040 ( .A(dout16_reg[90]), .Y(n421) );
  INVX1 U1041 ( .A(dout16_reg[74]), .Y(n420) );
  INVX1 U1042 ( .A(dout16_reg[58]), .Y(n419) );
  INVX1 U1043 ( .A(dout16_reg[42]), .Y(n418) );
  INVX1 U1044 ( .A(dout16_reg[26]), .Y(n417) );
  INVX1 U1045 ( .A(dout16_reg[10]), .Y(n416) );
  INVX1 U1046 ( .A(dout16_reg[123]), .Y(n407) );
  INVX1 U1047 ( .A(dout16_reg[107]), .Y(n406) );
  INVX1 U1048 ( .A(dout16_reg[91]), .Y(n405) );
  INVX1 U1049 ( .A(dout16_reg[75]), .Y(n404) );
  INVX1 U1050 ( .A(dout16_reg[59]), .Y(n403) );
  INVX1 U1051 ( .A(dout16_reg[43]), .Y(n402) );
  INVX1 U1052 ( .A(dout16_reg[27]), .Y(n401) );
  INVX1 U1053 ( .A(dout16_reg[11]), .Y(n400) );
  INVX1 U1054 ( .A(dout16_reg[124]), .Y(n391) );
  INVX1 U1055 ( .A(dout16_reg[108]), .Y(n390) );
  INVX1 U1056 ( .A(dout16_reg[92]), .Y(n389) );
  INVX1 U1057 ( .A(dout16_reg[76]), .Y(n388) );
  INVX1 U1058 ( .A(dout16_reg[60]), .Y(n387) );
  INVX1 U1059 ( .A(dout16_reg[44]), .Y(n386) );
  INVX1 U1060 ( .A(dout16_reg[28]), .Y(n385) );
  INVX1 U1061 ( .A(dout16_reg[12]), .Y(n384) );
  INVX1 U1062 ( .A(dout16_reg[125]), .Y(n375) );
  INVX1 U1063 ( .A(dout16_reg[109]), .Y(n374) );
  INVX1 U1064 ( .A(dout16_reg[93]), .Y(n373) );
  INVX1 U1065 ( .A(dout16_reg[77]), .Y(n372) );
  INVX1 U1066 ( .A(dout16_reg[61]), .Y(n371) );
  INVX1 U1067 ( .A(dout16_reg[45]), .Y(n370) );
  INVX1 U1068 ( .A(dout16_reg[29]), .Y(n369) );
  INVX1 U1069 ( .A(dout16_reg[13]), .Y(n368) );
  INVX1 U1070 ( .A(dout16_reg[126]), .Y(n359) );
  INVX1 U1071 ( .A(dout16_reg[110]), .Y(n358) );
  INVX1 U1072 ( .A(dout16_reg[94]), .Y(n357) );
  INVX1 U1073 ( .A(dout16_reg[78]), .Y(n356) );
  INVX1 U1074 ( .A(dout16_reg[62]), .Y(n355) );
  INVX1 U1075 ( .A(dout16_reg[46]), .Y(n354) );
  INVX1 U1076 ( .A(dout16_reg[30]), .Y(n353) );
  INVX1 U1077 ( .A(dout16_reg[14]), .Y(n352) );
  INVX1 U1078 ( .A(dout16_reg[127]), .Y(n343) );
  INVX1 U1079 ( .A(dout16_reg[111]), .Y(n342) );
  INVX1 U1080 ( .A(dout16_reg[95]), .Y(n341) );
  INVX1 U1081 ( .A(dout16_reg[79]), .Y(n340) );
  INVX1 U1082 ( .A(dout16_reg[63]), .Y(n339) );
  INVX1 U1083 ( .A(dout16_reg[47]), .Y(n338) );
  INVX1 U1084 ( .A(dout16_reg[31]), .Y(n337) );
  INVX1 U1085 ( .A(dout16_reg[15]), .Y(n336) );
  INVX1 U1086 ( .A(count[2]), .Y(n334) );
  ADDHXL U1087 ( .A(count[2]), .B(r71_carry[2]), .CO(r71_carry[3]), .S(N303)
         );
  ADDHXL U1088 ( .A(count[1]), .B(count[0]), .CO(r71_carry[2]), .S(N302) );
  ADDHXL U1089 ( .A(count[3]), .B(r71_carry[3]), .CO(r71_carry[4]), .S(N304)
         );
  INVX1 U1090 ( .A(dout16_reg[239]), .Y(n350) );
  INVX1 U1091 ( .A(dout8_reg[111]), .Y(n598) );
  INVX1 U1092 ( .A(dout4_reg[47]), .Y(n722) );
  INVX1 U1093 ( .A(dout16_reg[224]), .Y(n590) );
  INVX1 U1094 ( .A(dout16_reg[208]), .Y(n589) );
  INVX1 U1095 ( .A(dout16_reg[192]), .Y(n588) );
  INVX1 U1096 ( .A(dout16_reg[225]), .Y(n574) );
  INVX1 U1097 ( .A(dout16_reg[209]), .Y(n573) );
  INVX1 U1098 ( .A(dout16_reg[193]), .Y(n572) );
  INVX1 U1099 ( .A(dout16_reg[226]), .Y(n558) );
  INVX1 U1100 ( .A(dout16_reg[210]), .Y(n557) );
  INVX1 U1101 ( .A(dout16_reg[194]), .Y(n556) );
  INVX1 U1102 ( .A(dout16_reg[227]), .Y(n542) );
  INVX1 U1103 ( .A(dout16_reg[211]), .Y(n541) );
  INVX1 U1104 ( .A(dout16_reg[195]), .Y(n540) );
  INVX1 U1105 ( .A(dout16_reg[228]), .Y(n526) );
  INVX1 U1106 ( .A(dout16_reg[212]), .Y(n525) );
  INVX1 U1107 ( .A(dout16_reg[196]), .Y(n524) );
  INVX1 U1108 ( .A(dout16_reg[229]), .Y(n510) );
  INVX1 U1109 ( .A(dout16_reg[213]), .Y(n509) );
  INVX1 U1110 ( .A(dout16_reg[197]), .Y(n508) );
  INVX1 U1111 ( .A(dout16_reg[230]), .Y(n494) );
  INVX1 U1112 ( .A(dout16_reg[214]), .Y(n493) );
  INVX1 U1113 ( .A(dout16_reg[198]), .Y(n492) );
  INVX1 U1114 ( .A(dout16_reg[231]), .Y(n478) );
  INVX1 U1115 ( .A(dout16_reg[215]), .Y(n477) );
  INVX1 U1116 ( .A(dout16_reg[199]), .Y(n476) );
  INVX1 U1117 ( .A(dout16_reg[232]), .Y(n462) );
  INVX1 U1118 ( .A(dout16_reg[216]), .Y(n461) );
  INVX1 U1119 ( .A(dout16_reg[200]), .Y(n460) );
  INVX1 U1120 ( .A(dout16_reg[233]), .Y(n446) );
  INVX1 U1121 ( .A(dout16_reg[217]), .Y(n445) );
  INVX1 U1122 ( .A(dout16_reg[201]), .Y(n444) );
  INVX1 U1123 ( .A(dout16_reg[234]), .Y(n430) );
  INVX1 U1124 ( .A(dout16_reg[218]), .Y(n429) );
  INVX1 U1125 ( .A(dout16_reg[202]), .Y(n428) );
  INVX1 U1126 ( .A(dout16_reg[235]), .Y(n414) );
  INVX1 U1127 ( .A(dout16_reg[219]), .Y(n413) );
  INVX1 U1128 ( .A(dout16_reg[203]), .Y(n412) );
  INVX1 U1129 ( .A(dout16_reg[236]), .Y(n398) );
  INVX1 U1130 ( .A(dout16_reg[220]), .Y(n397) );
  INVX1 U1131 ( .A(dout16_reg[204]), .Y(n396) );
  INVX1 U1132 ( .A(dout16_reg[237]), .Y(n382) );
  INVX1 U1133 ( .A(dout16_reg[221]), .Y(n381) );
  INVX1 U1134 ( .A(dout16_reg[205]), .Y(n380) );
  INVX1 U1135 ( .A(dout16_reg[238]), .Y(n366) );
  INVX1 U1136 ( .A(dout16_reg[222]), .Y(n365) );
  INVX1 U1137 ( .A(dout16_reg[206]), .Y(n364) );
  INVX1 U1138 ( .A(dout16_reg[223]), .Y(n349) );
  INVX1 U1139 ( .A(dout16_reg[207]), .Y(n348) );
  INVX1 U1140 ( .A(dout8_reg[96]), .Y(n718) );
  INVX1 U1141 ( .A(dout8_reg[80]), .Y(n717) );
  INVX1 U1142 ( .A(dout8_reg[64]), .Y(n716) );
  INVX1 U1143 ( .A(dout8_reg[97]), .Y(n710) );
  INVX1 U1144 ( .A(dout8_reg[81]), .Y(n709) );
  INVX1 U1145 ( .A(dout8_reg[65]), .Y(n708) );
  INVX1 U1146 ( .A(dout8_reg[98]), .Y(n702) );
  INVX1 U1147 ( .A(dout8_reg[82]), .Y(n701) );
  INVX1 U1148 ( .A(dout8_reg[66]), .Y(n700) );
  INVX1 U1149 ( .A(dout8_reg[99]), .Y(n694) );
  INVX1 U1150 ( .A(dout8_reg[83]), .Y(n693) );
  INVX1 U1151 ( .A(dout8_reg[67]), .Y(n692) );
  INVX1 U1152 ( .A(dout8_reg[100]), .Y(n686) );
  INVX1 U1153 ( .A(dout8_reg[84]), .Y(n685) );
  INVX1 U1154 ( .A(dout8_reg[68]), .Y(n684) );
  INVX1 U1155 ( .A(dout8_reg[101]), .Y(n678) );
  INVX1 U1156 ( .A(dout8_reg[85]), .Y(n677) );
  INVX1 U1157 ( .A(dout8_reg[69]), .Y(n676) );
  INVX1 U1158 ( .A(dout8_reg[102]), .Y(n670) );
  INVX1 U1159 ( .A(dout8_reg[86]), .Y(n669) );
  INVX1 U1160 ( .A(dout8_reg[70]), .Y(n668) );
  INVX1 U1161 ( .A(dout8_reg[103]), .Y(n662) );
  INVX1 U1162 ( .A(dout8_reg[87]), .Y(n661) );
  INVX1 U1163 ( .A(dout8_reg[71]), .Y(n660) );
  INVX1 U1164 ( .A(dout8_reg[104]), .Y(n654) );
  INVX1 U1165 ( .A(dout8_reg[88]), .Y(n653) );
  INVX1 U1166 ( .A(dout8_reg[72]), .Y(n652) );
  INVX1 U1167 ( .A(dout8_reg[105]), .Y(n646) );
  INVX1 U1168 ( .A(dout8_reg[89]), .Y(n645) );
  INVX1 U1169 ( .A(dout8_reg[73]), .Y(n644) );
  INVX1 U1170 ( .A(dout8_reg[106]), .Y(n638) );
  INVX1 U1171 ( .A(dout8_reg[90]), .Y(n637) );
  INVX1 U1172 ( .A(dout8_reg[74]), .Y(n636) );
  INVX1 U1173 ( .A(dout8_reg[107]), .Y(n630) );
  INVX1 U1174 ( .A(dout8_reg[91]), .Y(n629) );
  INVX1 U1175 ( .A(dout8_reg[75]), .Y(n628) );
  INVX1 U1176 ( .A(dout8_reg[108]), .Y(n622) );
  INVX1 U1177 ( .A(dout8_reg[92]), .Y(n621) );
  INVX1 U1178 ( .A(dout8_reg[76]), .Y(n620) );
  INVX1 U1179 ( .A(dout8_reg[109]), .Y(n614) );
  INVX1 U1180 ( .A(dout8_reg[93]), .Y(n613) );
  INVX1 U1181 ( .A(dout8_reg[77]), .Y(n612) );
  INVX1 U1182 ( .A(dout8_reg[110]), .Y(n606) );
  INVX1 U1183 ( .A(dout8_reg[94]), .Y(n605) );
  INVX1 U1184 ( .A(dout8_reg[78]), .Y(n604) );
  INVX1 U1185 ( .A(dout8_reg[95]), .Y(n597) );
  INVX1 U1186 ( .A(dout8_reg[79]), .Y(n596) );
  INVX1 U1187 ( .A(dout4_reg[32]), .Y(n1246) );
  INVX1 U1188 ( .A(dout4_reg[16]), .Y(n1245) );
  INVX1 U1189 ( .A(dout4_reg[0]), .Y(n1244) );
  INVX1 U1190 ( .A(dout4_reg[33]), .Y(n1242) );
  INVX1 U1191 ( .A(dout4_reg[17]), .Y(n1241) );
  INVX1 U1192 ( .A(dout4_reg[1]), .Y(n1240) );
  INVX1 U1193 ( .A(dout4_reg[34]), .Y(n1238) );
  INVX1 U1194 ( .A(dout4_reg[18]), .Y(n1237) );
  INVX1 U1195 ( .A(dout4_reg[2]), .Y(n1236) );
  INVX1 U1196 ( .A(dout4_reg[35]), .Y(n1234) );
  INVX1 U1197 ( .A(dout4_reg[19]), .Y(n1233) );
  INVX1 U1198 ( .A(dout4_reg[3]), .Y(n1232) );
  INVX1 U1199 ( .A(dout4_reg[36]), .Y(n1230) );
  INVX1 U1200 ( .A(dout4_reg[20]), .Y(n1229) );
  INVX1 U1201 ( .A(dout4_reg[4]), .Y(n1228) );
  INVX1 U1202 ( .A(dout4_reg[37]), .Y(n1226) );
  INVX1 U1203 ( .A(dout4_reg[21]), .Y(n1225) );
  INVX1 U1204 ( .A(dout4_reg[5]), .Y(n1224) );
  INVX1 U1205 ( .A(dout4_reg[38]), .Y(n1222) );
  INVX1 U1206 ( .A(dout4_reg[22]), .Y(n1221) );
  INVX1 U1207 ( .A(dout4_reg[6]), .Y(n1220) );
  INVX1 U1208 ( .A(dout4_reg[39]), .Y(n1218) );
  INVX1 U1209 ( .A(dout4_reg[23]), .Y(n1217) );
  INVX1 U1210 ( .A(dout4_reg[7]), .Y(n1216) );
  INVX1 U1211 ( .A(dout4_reg[40]), .Y(n1214) );
  INVX1 U1212 ( .A(dout4_reg[24]), .Y(n1213) );
  INVX1 U1213 ( .A(dout4_reg[8]), .Y(n1212) );
  INVX1 U1214 ( .A(dout4_reg[41]), .Y(n1210) );
  INVX1 U1215 ( .A(dout4_reg[25]), .Y(n1209) );
  INVX1 U1216 ( .A(dout4_reg[9]), .Y(n1208) );
  INVX1 U1217 ( .A(dout4_reg[42]), .Y(n1206) );
  INVX1 U1218 ( .A(dout4_reg[26]), .Y(n1205) );
  INVX1 U1219 ( .A(dout4_reg[10]), .Y(n1204) );
  INVX1 U1220 ( .A(dout4_reg[43]), .Y(n1202) );
  INVX1 U1221 ( .A(dout4_reg[27]), .Y(n1201) );
  INVX1 U1222 ( .A(dout4_reg[11]), .Y(n1200) );
  INVX1 U1223 ( .A(dout4_reg[44]), .Y(n739) );
  INVX1 U1224 ( .A(dout4_reg[28]), .Y(n738) );
  INVX1 U1225 ( .A(dout4_reg[12]), .Y(n735) );
  INVX1 U1226 ( .A(dout4_reg[45]), .Y(n730) );
  INVX1 U1227 ( .A(dout4_reg[29]), .Y(n729) );
  INVX1 U1228 ( .A(dout4_reg[13]), .Y(n728) );
  INVX1 U1229 ( .A(dout4_reg[46]), .Y(n726) );
  INVX1 U1230 ( .A(dout4_reg[30]), .Y(n725) );
  INVX1 U1231 ( .A(dout4_reg[14]), .Y(n724) );
  INVX1 U1232 ( .A(dout4_reg[31]), .Y(n721) );
  INVX1 U1233 ( .A(dout4_reg[15]), .Y(n720) );
  INVX1 U1234 ( .A(dout16_reg[240]), .Y(n591) );
  INVX1 U1235 ( .A(dout16_reg[241]), .Y(n575) );
  INVX1 U1236 ( .A(dout16_reg[242]), .Y(n559) );
  INVX1 U1237 ( .A(dout16_reg[243]), .Y(n543) );
  INVX1 U1238 ( .A(dout16_reg[244]), .Y(n527) );
  INVX1 U1239 ( .A(dout16_reg[245]), .Y(n511) );
  INVX1 U1240 ( .A(dout16_reg[246]), .Y(n495) );
  INVX1 U1241 ( .A(dout16_reg[247]), .Y(n479) );
  INVX1 U1242 ( .A(dout16_reg[248]), .Y(n463) );
  INVX1 U1243 ( .A(dout16_reg[249]), .Y(n447) );
  INVX1 U1244 ( .A(dout16_reg[250]), .Y(n431) );
  INVX1 U1245 ( .A(dout16_reg[251]), .Y(n415) );
  INVX1 U1246 ( .A(dout16_reg[252]), .Y(n399) );
  INVX1 U1247 ( .A(dout16_reg[253]), .Y(n383) );
  INVX1 U1248 ( .A(dout16_reg[254]), .Y(n367) );
  INVX1 U1249 ( .A(dout16_reg[255]), .Y(n351) );
  INVX1 U1250 ( .A(dout8_reg[112]), .Y(n719) );
  INVX1 U1251 ( .A(dout8_reg[113]), .Y(n711) );
  INVX1 U1252 ( .A(dout8_reg[114]), .Y(n703) );
  INVX1 U1253 ( .A(dout8_reg[115]), .Y(n695) );
  INVX1 U1254 ( .A(dout8_reg[116]), .Y(n687) );
  INVX1 U1255 ( .A(dout8_reg[117]), .Y(n679) );
  INVX1 U1256 ( .A(dout8_reg[118]), .Y(n671) );
  INVX1 U1257 ( .A(dout8_reg[119]), .Y(n663) );
  INVX1 U1258 ( .A(dout8_reg[120]), .Y(n655) );
  INVX1 U1259 ( .A(dout8_reg[121]), .Y(n647) );
  INVX1 U1260 ( .A(dout8_reg[122]), .Y(n639) );
  INVX1 U1261 ( .A(dout8_reg[123]), .Y(n631) );
  INVX1 U1262 ( .A(dout8_reg[124]), .Y(n623) );
  INVX1 U1263 ( .A(dout8_reg[125]), .Y(n615) );
  INVX1 U1264 ( .A(dout8_reg[126]), .Y(n607) );
  INVX1 U1265 ( .A(dout8_reg[127]), .Y(n599) );
  INVX1 U1266 ( .A(dout4_reg[48]), .Y(n1247) );
  INVX1 U1267 ( .A(dout4_reg[49]), .Y(n1243) );
  INVX1 U1268 ( .A(dout4_reg[50]), .Y(n1239) );
  INVX1 U1269 ( .A(dout4_reg[51]), .Y(n1235) );
  INVX1 U1270 ( .A(dout4_reg[52]), .Y(n1231) );
  INVX1 U1271 ( .A(dout4_reg[53]), .Y(n1227) );
  INVX1 U1272 ( .A(dout4_reg[54]), .Y(n1223) );
  INVX1 U1273 ( .A(dout4_reg[55]), .Y(n1219) );
  INVX1 U1274 ( .A(dout4_reg[56]), .Y(n1215) );
  INVX1 U1275 ( .A(dout4_reg[57]), .Y(n1211) );
  INVX1 U1276 ( .A(dout4_reg[58]), .Y(n1207) );
  INVX1 U1277 ( .A(dout4_reg[59]), .Y(n1203) );
  INVX1 U1278 ( .A(dout4_reg[60]), .Y(n1199) );
  INVX1 U1279 ( .A(dout4_reg[61]), .Y(n732) );
  INVX1 U1280 ( .A(dout4_reg[62]), .Y(n727) );
  INVX1 U1281 ( .A(dout4_reg[63]), .Y(n723) );
  NAND2X1 U1282 ( .A(mode_reg[1]), .B(n333), .Y(n741) );
  NAND2X1 U1283 ( .A(mode_reg[0]), .B(n332), .Y(n743) );
endmodule


module even_odd_0 ( clk, rstn, mode, start, din, dout, even_odd_ready, 
        mode_out );
  input [1:0] mode;
  input [255:0] din;
  output [255:0] dout;
  output [1:0] mode_out;
  input clk, rstn, start;
  output even_odd_ready;
  wire   N275, n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n153, n156, n159, n162, n165, n168, n171,
         n174, n177, n180, n183, n186, n189, n192, n195, n198, n200, n202,
         n204, n206, n208, n210, n212, n214, n216, n218, n220, n222, n224,
         n226, n228, n230, n233, n236, n239, n242, n245, n248, n251, n254,
         n257, n260, n263, n266, n269, n272, n275, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n296, n298, n300, n302, n304, n306, n308, n310, n312,
         n314, n316, n318, n320, n322, n324, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n2, n19, n20, n149, n150, n151,
         n152, n154, n155, n157, n158, n160, n161, n163, n164, n166, n167,
         n169, n170, n172, n173, n175, n176, n178, n179, n181, n182, n184,
         n185, n187, n188, n190, n191, n193, n194, n196, n197, n199, n201,
         n203, n205, n207, n209, n211, n213, n215, n217, n219, n221, n223,
         n225, n227, n229, n231, n232, n234, n235, n237, n238, n240, n241,
         n243, n244, n246, n247, n249, n250, n252, n253, n255, n256, n258,
         n259, n261, n262, n264, n265, n267, n268, n270, n271, n273, n274,
         n276, n277, n295, n297, n299, n301, n303, n305, n307, n309, n311,
         n313, n315, n317, n319, n321, n323, n325, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649;

  DFFRHQX1 dout_reg_15_ ( .D(n380), .CK(clk), .RN(rstn), .Q(dout[15]) );
  DFFRHQX1 dout_reg_14_ ( .D(n379), .CK(clk), .RN(rstn), .Q(dout[14]) );
  DFFRHQX1 dout_reg_13_ ( .D(n378), .CK(clk), .RN(rstn), .Q(dout[13]) );
  DFFRHQX1 dout_reg_12_ ( .D(n377), .CK(clk), .RN(rstn), .Q(dout[12]) );
  DFFRHQX1 dout_reg_11_ ( .D(n376), .CK(clk), .RN(rstn), .Q(dout[11]) );
  DFFRHQX1 dout_reg_10_ ( .D(n375), .CK(clk), .RN(rstn), .Q(dout[10]) );
  DFFRHQX1 dout_reg_9_ ( .D(n374), .CK(clk), .RN(rstn), .Q(dout[9]) );
  DFFRHQX1 dout_reg_8_ ( .D(n373), .CK(clk), .RN(rstn), .Q(dout[8]) );
  DFFRHQX1 dout_reg_7_ ( .D(n372), .CK(clk), .RN(rstn), .Q(dout[7]) );
  DFFRHQX1 dout_reg_6_ ( .D(n371), .CK(clk), .RN(rstn), .Q(dout[6]) );
  DFFRHQX1 dout_reg_5_ ( .D(n370), .CK(clk), .RN(rstn), .Q(dout[5]) );
  DFFRHQX1 dout_reg_4_ ( .D(n369), .CK(clk), .RN(rstn), .Q(dout[4]) );
  DFFRHQX1 dout_reg_3_ ( .D(n368), .CK(clk), .RN(rstn), .Q(dout[3]) );
  DFFRHQX1 dout_reg_2_ ( .D(n367), .CK(clk), .RN(rstn), .Q(dout[2]) );
  DFFRHQX1 dout_reg_1_ ( .D(n366), .CK(clk), .RN(rstn), .Q(dout[1]) );
  DFFRHQX1 dout_reg_0_ ( .D(n365), .CK(clk), .RN(rstn), .Q(dout[0]) );
  DFFRHQX1 mode_out_reg_1_ ( .D(n622), .CK(clk), .RN(rstn), .Q(mode_out[1]) );
  DFFRHQX1 mode_out_reg_0_ ( .D(n621), .CK(clk), .RN(rstn), .Q(mode_out[0]) );
  DFFRHQX1 dout_reg_255_ ( .D(n620), .CK(clk), .RN(rstn), .Q(dout[255]) );
  DFFRHQX1 dout_reg_254_ ( .D(n619), .CK(clk), .RN(rstn), .Q(dout[254]) );
  DFFRHQX1 dout_reg_253_ ( .D(n618), .CK(clk), .RN(rstn), .Q(dout[253]) );
  DFFRHQX1 dout_reg_252_ ( .D(n617), .CK(clk), .RN(rstn), .Q(dout[252]) );
  DFFRHQX1 dout_reg_251_ ( .D(n616), .CK(clk), .RN(rstn), .Q(dout[251]) );
  DFFRHQX1 dout_reg_250_ ( .D(n615), .CK(clk), .RN(rstn), .Q(dout[250]) );
  DFFRHQX1 dout_reg_249_ ( .D(n614), .CK(clk), .RN(rstn), .Q(dout[249]) );
  DFFRHQX1 dout_reg_248_ ( .D(n613), .CK(clk), .RN(rstn), .Q(dout[248]) );
  DFFRHQX1 dout_reg_247_ ( .D(n612), .CK(clk), .RN(rstn), .Q(dout[247]) );
  DFFRHQX1 dout_reg_246_ ( .D(n611), .CK(clk), .RN(rstn), .Q(dout[246]) );
  DFFRHQX1 dout_reg_245_ ( .D(n610), .CK(clk), .RN(rstn), .Q(dout[245]) );
  DFFRHQX1 dout_reg_244_ ( .D(n609), .CK(clk), .RN(rstn), .Q(dout[244]) );
  DFFRHQX1 dout_reg_243_ ( .D(n608), .CK(clk), .RN(rstn), .Q(dout[243]) );
  DFFRHQX1 dout_reg_242_ ( .D(n607), .CK(clk), .RN(rstn), .Q(dout[242]) );
  DFFRHQX1 dout_reg_241_ ( .D(n606), .CK(clk), .RN(rstn), .Q(dout[241]) );
  DFFRHQX1 dout_reg_240_ ( .D(n605), .CK(clk), .RN(rstn), .Q(dout[240]) );
  DFFRHQX1 dout_reg_127_ ( .D(n492), .CK(clk), .RN(rstn), .Q(dout[127]) );
  DFFRHQX1 dout_reg_126_ ( .D(n491), .CK(clk), .RN(rstn), .Q(dout[126]) );
  DFFRHQX1 dout_reg_125_ ( .D(n490), .CK(clk), .RN(rstn), .Q(dout[125]) );
  DFFRHQX1 dout_reg_124_ ( .D(n489), .CK(clk), .RN(rstn), .Q(dout[124]) );
  DFFRHQX1 dout_reg_123_ ( .D(n488), .CK(clk), .RN(rstn), .Q(dout[123]) );
  DFFRHQX1 dout_reg_122_ ( .D(n487), .CK(clk), .RN(rstn), .Q(dout[122]) );
  DFFRHQX1 dout_reg_121_ ( .D(n486), .CK(clk), .RN(rstn), .Q(dout[121]) );
  DFFRHQX1 dout_reg_120_ ( .D(n485), .CK(clk), .RN(rstn), .Q(dout[120]) );
  DFFRHQX1 dout_reg_119_ ( .D(n484), .CK(clk), .RN(rstn), .Q(dout[119]) );
  DFFRHQX1 dout_reg_118_ ( .D(n483), .CK(clk), .RN(rstn), .Q(dout[118]) );
  DFFRHQX1 dout_reg_117_ ( .D(n482), .CK(clk), .RN(rstn), .Q(dout[117]) );
  DFFRHQX1 dout_reg_116_ ( .D(n481), .CK(clk), .RN(rstn), .Q(dout[116]) );
  DFFRHQX1 dout_reg_115_ ( .D(n480), .CK(clk), .RN(rstn), .Q(dout[115]) );
  DFFRHQX1 dout_reg_114_ ( .D(n479), .CK(clk), .RN(rstn), .Q(dout[114]) );
  DFFRHQX1 dout_reg_113_ ( .D(n478), .CK(clk), .RN(rstn), .Q(dout[113]) );
  DFFRHQX1 dout_reg_112_ ( .D(n477), .CK(clk), .RN(rstn), .Q(dout[112]) );
  DFFRHQX1 dout_reg_111_ ( .D(n476), .CK(clk), .RN(rstn), .Q(dout[111]) );
  DFFRHQX1 dout_reg_110_ ( .D(n475), .CK(clk), .RN(rstn), .Q(dout[110]) );
  DFFRHQX1 dout_reg_109_ ( .D(n474), .CK(clk), .RN(rstn), .Q(dout[109]) );
  DFFRHQX1 dout_reg_108_ ( .D(n473), .CK(clk), .RN(rstn), .Q(dout[108]) );
  DFFRHQX1 dout_reg_107_ ( .D(n472), .CK(clk), .RN(rstn), .Q(dout[107]) );
  DFFRHQX1 dout_reg_106_ ( .D(n471), .CK(clk), .RN(rstn), .Q(dout[106]) );
  DFFRHQX1 dout_reg_105_ ( .D(n470), .CK(clk), .RN(rstn), .Q(dout[105]) );
  DFFRHQX1 dout_reg_104_ ( .D(n469), .CK(clk), .RN(rstn), .Q(dout[104]) );
  DFFRHQX1 dout_reg_103_ ( .D(n468), .CK(clk), .RN(rstn), .Q(dout[103]) );
  DFFRHQX1 dout_reg_102_ ( .D(n467), .CK(clk), .RN(rstn), .Q(dout[102]) );
  DFFRHQX1 dout_reg_101_ ( .D(n466), .CK(clk), .RN(rstn), .Q(dout[101]) );
  DFFRHQX1 dout_reg_100_ ( .D(n465), .CK(clk), .RN(rstn), .Q(dout[100]) );
  DFFRHQX1 dout_reg_99_ ( .D(n464), .CK(clk), .RN(rstn), .Q(dout[99]) );
  DFFRHQX1 dout_reg_98_ ( .D(n463), .CK(clk), .RN(rstn), .Q(dout[98]) );
  DFFRHQX1 dout_reg_97_ ( .D(n462), .CK(clk), .RN(rstn), .Q(dout[97]) );
  DFFRHQX1 dout_reg_96_ ( .D(n461), .CK(clk), .RN(rstn), .Q(dout[96]) );
  DFFRHQX1 dout_reg_95_ ( .D(n460), .CK(clk), .RN(rstn), .Q(dout[95]) );
  DFFRHQX1 dout_reg_94_ ( .D(n459), .CK(clk), .RN(rstn), .Q(dout[94]) );
  DFFRHQX1 dout_reg_93_ ( .D(n458), .CK(clk), .RN(rstn), .Q(dout[93]) );
  DFFRHQX1 dout_reg_92_ ( .D(n457), .CK(clk), .RN(rstn), .Q(dout[92]) );
  DFFRHQX1 dout_reg_91_ ( .D(n456), .CK(clk), .RN(rstn), .Q(dout[91]) );
  DFFRHQX1 dout_reg_90_ ( .D(n455), .CK(clk), .RN(rstn), .Q(dout[90]) );
  DFFRHQX1 dout_reg_89_ ( .D(n454), .CK(clk), .RN(rstn), .Q(dout[89]) );
  DFFRHQX1 dout_reg_88_ ( .D(n453), .CK(clk), .RN(rstn), .Q(dout[88]) );
  DFFRHQX1 dout_reg_87_ ( .D(n452), .CK(clk), .RN(rstn), .Q(dout[87]) );
  DFFRHQX1 dout_reg_86_ ( .D(n451), .CK(clk), .RN(rstn), .Q(dout[86]) );
  DFFRHQX1 dout_reg_85_ ( .D(n450), .CK(clk), .RN(rstn), .Q(dout[85]) );
  DFFRHQX1 dout_reg_84_ ( .D(n449), .CK(clk), .RN(rstn), .Q(dout[84]) );
  DFFRHQX1 dout_reg_83_ ( .D(n448), .CK(clk), .RN(rstn), .Q(dout[83]) );
  DFFRHQX1 dout_reg_82_ ( .D(n447), .CK(clk), .RN(rstn), .Q(dout[82]) );
  DFFRHQX1 dout_reg_81_ ( .D(n446), .CK(clk), .RN(rstn), .Q(dout[81]) );
  DFFRHQX1 dout_reg_80_ ( .D(n445), .CK(clk), .RN(rstn), .Q(dout[80]) );
  DFFRHQX1 dout_reg_79_ ( .D(n444), .CK(clk), .RN(rstn), .Q(dout[79]) );
  DFFRHQX1 dout_reg_78_ ( .D(n443), .CK(clk), .RN(rstn), .Q(dout[78]) );
  DFFRHQX1 dout_reg_77_ ( .D(n442), .CK(clk), .RN(rstn), .Q(dout[77]) );
  DFFRHQX1 dout_reg_76_ ( .D(n441), .CK(clk), .RN(rstn), .Q(dout[76]) );
  DFFRHQX1 dout_reg_75_ ( .D(n440), .CK(clk), .RN(rstn), .Q(dout[75]) );
  DFFRHQX1 dout_reg_74_ ( .D(n439), .CK(clk), .RN(rstn), .Q(dout[74]) );
  DFFRHQX1 dout_reg_73_ ( .D(n438), .CK(clk), .RN(rstn), .Q(dout[73]) );
  DFFRHQX1 dout_reg_72_ ( .D(n437), .CK(clk), .RN(rstn), .Q(dout[72]) );
  DFFRHQX1 dout_reg_71_ ( .D(n436), .CK(clk), .RN(rstn), .Q(dout[71]) );
  DFFRHQX1 dout_reg_70_ ( .D(n435), .CK(clk), .RN(rstn), .Q(dout[70]) );
  DFFRHQX1 dout_reg_69_ ( .D(n434), .CK(clk), .RN(rstn), .Q(dout[69]) );
  DFFRHQX1 dout_reg_68_ ( .D(n433), .CK(clk), .RN(rstn), .Q(dout[68]) );
  DFFRHQX1 dout_reg_67_ ( .D(n432), .CK(clk), .RN(rstn), .Q(dout[67]) );
  DFFRHQX1 dout_reg_66_ ( .D(n431), .CK(clk), .RN(rstn), .Q(dout[66]) );
  DFFRHQX1 dout_reg_65_ ( .D(n430), .CK(clk), .RN(rstn), .Q(dout[65]) );
  DFFRHQX1 dout_reg_64_ ( .D(n429), .CK(clk), .RN(rstn), .Q(dout[64]) );
  DFFRHQX1 dout_reg_63_ ( .D(n428), .CK(clk), .RN(rstn), .Q(dout[63]) );
  DFFRHQX1 dout_reg_62_ ( .D(n427), .CK(clk), .RN(rstn), .Q(dout[62]) );
  DFFRHQX1 dout_reg_61_ ( .D(n426), .CK(clk), .RN(rstn), .Q(dout[61]) );
  DFFRHQX1 dout_reg_60_ ( .D(n425), .CK(clk), .RN(rstn), .Q(dout[60]) );
  DFFRHQX1 dout_reg_59_ ( .D(n424), .CK(clk), .RN(rstn), .Q(dout[59]) );
  DFFRHQX1 dout_reg_58_ ( .D(n423), .CK(clk), .RN(rstn), .Q(dout[58]) );
  DFFRHQX1 dout_reg_57_ ( .D(n422), .CK(clk), .RN(rstn), .Q(dout[57]) );
  DFFRHQX1 dout_reg_56_ ( .D(n421), .CK(clk), .RN(rstn), .Q(dout[56]) );
  DFFRHQX1 dout_reg_55_ ( .D(n420), .CK(clk), .RN(rstn), .Q(dout[55]) );
  DFFRHQX1 dout_reg_54_ ( .D(n419), .CK(clk), .RN(rstn), .Q(dout[54]) );
  DFFRHQX1 dout_reg_53_ ( .D(n418), .CK(clk), .RN(rstn), .Q(dout[53]) );
  DFFRHQX1 dout_reg_52_ ( .D(n417), .CK(clk), .RN(rstn), .Q(dout[52]) );
  DFFRHQX1 dout_reg_51_ ( .D(n416), .CK(clk), .RN(rstn), .Q(dout[51]) );
  DFFRHQX1 dout_reg_50_ ( .D(n415), .CK(clk), .RN(rstn), .Q(dout[50]) );
  DFFRHQX1 dout_reg_49_ ( .D(n414), .CK(clk), .RN(rstn), .Q(dout[49]) );
  DFFRHQX1 dout_reg_48_ ( .D(n413), .CK(clk), .RN(rstn), .Q(dout[48]) );
  DFFRHQX1 dout_reg_47_ ( .D(n412), .CK(clk), .RN(rstn), .Q(dout[47]) );
  DFFRHQX1 dout_reg_46_ ( .D(n411), .CK(clk), .RN(rstn), .Q(dout[46]) );
  DFFRHQX1 dout_reg_45_ ( .D(n410), .CK(clk), .RN(rstn), .Q(dout[45]) );
  DFFRHQX1 dout_reg_44_ ( .D(n409), .CK(clk), .RN(rstn), .Q(dout[44]) );
  DFFRHQX1 dout_reg_43_ ( .D(n408), .CK(clk), .RN(rstn), .Q(dout[43]) );
  DFFRHQX1 dout_reg_42_ ( .D(n407), .CK(clk), .RN(rstn), .Q(dout[42]) );
  DFFRHQX1 dout_reg_41_ ( .D(n406), .CK(clk), .RN(rstn), .Q(dout[41]) );
  DFFRHQX1 dout_reg_40_ ( .D(n405), .CK(clk), .RN(rstn), .Q(dout[40]) );
  DFFRHQX1 dout_reg_39_ ( .D(n404), .CK(clk), .RN(rstn), .Q(dout[39]) );
  DFFRHQX1 dout_reg_38_ ( .D(n403), .CK(clk), .RN(rstn), .Q(dout[38]) );
  DFFRHQX1 dout_reg_37_ ( .D(n402), .CK(clk), .RN(rstn), .Q(dout[37]) );
  DFFRHQX1 dout_reg_36_ ( .D(n401), .CK(clk), .RN(rstn), .Q(dout[36]) );
  DFFRHQX1 dout_reg_35_ ( .D(n400), .CK(clk), .RN(rstn), .Q(dout[35]) );
  DFFRHQX1 dout_reg_34_ ( .D(n399), .CK(clk), .RN(rstn), .Q(dout[34]) );
  DFFRHQX1 dout_reg_33_ ( .D(n398), .CK(clk), .RN(rstn), .Q(dout[33]) );
  DFFRHQX1 dout_reg_32_ ( .D(n397), .CK(clk), .RN(rstn), .Q(dout[32]) );
  DFFRHQX1 dout_reg_31_ ( .D(n396), .CK(clk), .RN(rstn), .Q(dout[31]) );
  DFFRHQX1 dout_reg_30_ ( .D(n395), .CK(clk), .RN(rstn), .Q(dout[30]) );
  DFFRHQX1 dout_reg_29_ ( .D(n394), .CK(clk), .RN(rstn), .Q(dout[29]) );
  DFFRHQX1 dout_reg_28_ ( .D(n393), .CK(clk), .RN(rstn), .Q(dout[28]) );
  DFFRHQX1 dout_reg_27_ ( .D(n392), .CK(clk), .RN(rstn), .Q(dout[27]) );
  DFFRHQX1 dout_reg_26_ ( .D(n391), .CK(clk), .RN(rstn), .Q(dout[26]) );
  DFFRHQX1 dout_reg_25_ ( .D(n390), .CK(clk), .RN(rstn), .Q(dout[25]) );
  DFFRHQX1 dout_reg_24_ ( .D(n389), .CK(clk), .RN(rstn), .Q(dout[24]) );
  DFFRHQX1 dout_reg_23_ ( .D(n388), .CK(clk), .RN(rstn), .Q(dout[23]) );
  DFFRHQX1 dout_reg_22_ ( .D(n387), .CK(clk), .RN(rstn), .Q(dout[22]) );
  DFFRHQX1 dout_reg_21_ ( .D(n386), .CK(clk), .RN(rstn), .Q(dout[21]) );
  DFFRHQX1 dout_reg_20_ ( .D(n385), .CK(clk), .RN(rstn), .Q(dout[20]) );
  DFFRHQX1 dout_reg_19_ ( .D(n384), .CK(clk), .RN(rstn), .Q(dout[19]) );
  DFFRHQX1 dout_reg_18_ ( .D(n383), .CK(clk), .RN(rstn), .Q(dout[18]) );
  DFFRHQX1 dout_reg_17_ ( .D(n382), .CK(clk), .RN(rstn), .Q(dout[17]) );
  DFFRHQX1 dout_reg_16_ ( .D(n381), .CK(clk), .RN(rstn), .Q(dout[16]) );
  DFFRHQX1 dout_reg_223_ ( .D(n588), .CK(clk), .RN(rstn), .Q(dout[223]) );
  DFFRHQX1 dout_reg_222_ ( .D(n587), .CK(clk), .RN(rstn), .Q(dout[222]) );
  DFFRHQX1 dout_reg_221_ ( .D(n586), .CK(clk), .RN(rstn), .Q(dout[221]) );
  DFFRHQX1 dout_reg_220_ ( .D(n585), .CK(clk), .RN(rstn), .Q(dout[220]) );
  DFFRHQX1 dout_reg_219_ ( .D(n584), .CK(clk), .RN(rstn), .Q(dout[219]) );
  DFFRHQX1 dout_reg_218_ ( .D(n583), .CK(clk), .RN(rstn), .Q(dout[218]) );
  DFFRHQX1 dout_reg_217_ ( .D(n582), .CK(clk), .RN(rstn), .Q(dout[217]) );
  DFFRHQX1 dout_reg_216_ ( .D(n581), .CK(clk), .RN(rstn), .Q(dout[216]) );
  DFFRHQX1 dout_reg_215_ ( .D(n580), .CK(clk), .RN(rstn), .Q(dout[215]) );
  DFFRHQX1 dout_reg_214_ ( .D(n579), .CK(clk), .RN(rstn), .Q(dout[214]) );
  DFFRHQX1 dout_reg_213_ ( .D(n578), .CK(clk), .RN(rstn), .Q(dout[213]) );
  DFFRHQX1 dout_reg_212_ ( .D(n577), .CK(clk), .RN(rstn), .Q(dout[212]) );
  DFFRHQX1 dout_reg_211_ ( .D(n576), .CK(clk), .RN(rstn), .Q(dout[211]) );
  DFFRHQX1 dout_reg_210_ ( .D(n575), .CK(clk), .RN(rstn), .Q(dout[210]) );
  DFFRHQX1 dout_reg_209_ ( .D(n574), .CK(clk), .RN(rstn), .Q(dout[209]) );
  DFFRHQX1 dout_reg_208_ ( .D(n573), .CK(clk), .RN(rstn), .Q(dout[208]) );
  DFFRHQX1 dout_reg_143_ ( .D(n508), .CK(clk), .RN(rstn), .Q(dout[143]) );
  DFFRHQX1 dout_reg_191_ ( .D(n556), .CK(clk), .RN(rstn), .Q(dout[191]) );
  DFFRHQX1 dout_reg_175_ ( .D(n540), .CK(clk), .RN(rstn), .Q(dout[175]) );
  DFFRHQX1 dout_reg_159_ ( .D(n524), .CK(clk), .RN(rstn), .Q(dout[159]) );
  DFFRHQX1 dout_reg_142_ ( .D(n507), .CK(clk), .RN(rstn), .Q(dout[142]) );
  DFFRHQX1 dout_reg_141_ ( .D(n506), .CK(clk), .RN(rstn), .Q(dout[141]) );
  DFFRHQX1 dout_reg_239_ ( .D(n604), .CK(clk), .RN(rstn), .Q(dout[239]) );
  DFFRHQX1 dout_reg_207_ ( .D(n572), .CK(clk), .RN(rstn), .Q(dout[207]) );
  DFFRHQX1 dout_reg_190_ ( .D(n555), .CK(clk), .RN(rstn), .Q(dout[190]) );
  DFFRHQX1 dout_reg_189_ ( .D(n554), .CK(clk), .RN(rstn), .Q(dout[189]) );
  DFFRHQX1 dout_reg_174_ ( .D(n539), .CK(clk), .RN(rstn), .Q(dout[174]) );
  DFFRHQX1 dout_reg_173_ ( .D(n538), .CK(clk), .RN(rstn), .Q(dout[173]) );
  DFFRHQX1 dout_reg_158_ ( .D(n523), .CK(clk), .RN(rstn), .Q(dout[158]) );
  DFFRHQX1 dout_reg_157_ ( .D(n522), .CK(clk), .RN(rstn), .Q(dout[157]) );
  DFFRHQX1 dout_reg_238_ ( .D(n603), .CK(clk), .RN(rstn), .Q(dout[238]) );
  DFFRHQX1 dout_reg_237_ ( .D(n602), .CK(clk), .RN(rstn), .Q(dout[237]) );
  DFFRHQX1 dout_reg_206_ ( .D(n571), .CK(clk), .RN(rstn), .Q(dout[206]) );
  DFFRHQX1 dout_reg_205_ ( .D(n570), .CK(clk), .RN(rstn), .Q(dout[205]) );
  DFFRHQX1 dout_reg_140_ ( .D(n505), .CK(clk), .RN(rstn), .Q(dout[140]) );
  DFFRHQX1 dout_reg_139_ ( .D(n504), .CK(clk), .RN(rstn), .Q(dout[139]) );
  DFFRHQX1 dout_reg_138_ ( .D(n503), .CK(clk), .RN(rstn), .Q(dout[138]) );
  DFFRHQX1 dout_reg_137_ ( .D(n502), .CK(clk), .RN(rstn), .Q(dout[137]) );
  DFFRHQX1 dout_reg_188_ ( .D(n553), .CK(clk), .RN(rstn), .Q(dout[188]) );
  DFFRHQX1 dout_reg_187_ ( .D(n552), .CK(clk), .RN(rstn), .Q(dout[187]) );
  DFFRHQX1 dout_reg_186_ ( .D(n551), .CK(clk), .RN(rstn), .Q(dout[186]) );
  DFFRHQX1 dout_reg_185_ ( .D(n550), .CK(clk), .RN(rstn), .Q(dout[185]) );
  DFFRHQX1 dout_reg_172_ ( .D(n537), .CK(clk), .RN(rstn), .Q(dout[172]) );
  DFFRHQX1 dout_reg_171_ ( .D(n536), .CK(clk), .RN(rstn), .Q(dout[171]) );
  DFFRHQX1 dout_reg_170_ ( .D(n535), .CK(clk), .RN(rstn), .Q(dout[170]) );
  DFFRHQX1 dout_reg_169_ ( .D(n534), .CK(clk), .RN(rstn), .Q(dout[169]) );
  DFFRHQX1 dout_reg_156_ ( .D(n521), .CK(clk), .RN(rstn), .Q(dout[156]) );
  DFFRHQX1 dout_reg_155_ ( .D(n520), .CK(clk), .RN(rstn), .Q(dout[155]) );
  DFFRHQX1 dout_reg_154_ ( .D(n519), .CK(clk), .RN(rstn), .Q(dout[154]) );
  DFFRHQX1 dout_reg_153_ ( .D(n518), .CK(clk), .RN(rstn), .Q(dout[153]) );
  DFFRHQX1 dout_reg_236_ ( .D(n601), .CK(clk), .RN(rstn), .Q(dout[236]) );
  DFFRHQX1 dout_reg_235_ ( .D(n600), .CK(clk), .RN(rstn), .Q(dout[235]) );
  DFFRHQX1 dout_reg_234_ ( .D(n599), .CK(clk), .RN(rstn), .Q(dout[234]) );
  DFFRHQX1 dout_reg_233_ ( .D(n598), .CK(clk), .RN(rstn), .Q(dout[233]) );
  DFFRHQX1 dout_reg_204_ ( .D(n569), .CK(clk), .RN(rstn), .Q(dout[204]) );
  DFFRHQX1 dout_reg_203_ ( .D(n568), .CK(clk), .RN(rstn), .Q(dout[203]) );
  DFFRHQX1 dout_reg_202_ ( .D(n567), .CK(clk), .RN(rstn), .Q(dout[202]) );
  DFFRHQX1 dout_reg_201_ ( .D(n566), .CK(clk), .RN(rstn), .Q(dout[201]) );
  DFFRHQX1 dout_reg_136_ ( .D(n501), .CK(clk), .RN(rstn), .Q(dout[136]) );
  DFFRHQX1 dout_reg_135_ ( .D(n500), .CK(clk), .RN(rstn), .Q(dout[135]) );
  DFFRHQX1 dout_reg_134_ ( .D(n499), .CK(clk), .RN(rstn), .Q(dout[134]) );
  DFFRHQX1 dout_reg_133_ ( .D(n498), .CK(clk), .RN(rstn), .Q(dout[133]) );
  DFFRHQX1 dout_reg_132_ ( .D(n497), .CK(clk), .RN(rstn), .Q(dout[132]) );
  DFFRHQX1 dout_reg_131_ ( .D(n496), .CK(clk), .RN(rstn), .Q(dout[131]) );
  DFFRHQX1 dout_reg_130_ ( .D(n495), .CK(clk), .RN(rstn), .Q(dout[130]) );
  DFFRHQX1 dout_reg_184_ ( .D(n549), .CK(clk), .RN(rstn), .Q(dout[184]) );
  DFFRHQX1 dout_reg_183_ ( .D(n548), .CK(clk), .RN(rstn), .Q(dout[183]) );
  DFFRHQX1 dout_reg_182_ ( .D(n547), .CK(clk), .RN(rstn), .Q(dout[182]) );
  DFFRHQX1 dout_reg_181_ ( .D(n546), .CK(clk), .RN(rstn), .Q(dout[181]) );
  DFFRHQX1 dout_reg_180_ ( .D(n545), .CK(clk), .RN(rstn), .Q(dout[180]) );
  DFFRHQX1 dout_reg_179_ ( .D(n544), .CK(clk), .RN(rstn), .Q(dout[179]) );
  DFFRHQX1 dout_reg_178_ ( .D(n543), .CK(clk), .RN(rstn), .Q(dout[178]) );
  DFFRHQX1 dout_reg_168_ ( .D(n533), .CK(clk), .RN(rstn), .Q(dout[168]) );
  DFFRHQX1 dout_reg_167_ ( .D(n532), .CK(clk), .RN(rstn), .Q(dout[167]) );
  DFFRHQX1 dout_reg_166_ ( .D(n531), .CK(clk), .RN(rstn), .Q(dout[166]) );
  DFFRHQX1 dout_reg_165_ ( .D(n530), .CK(clk), .RN(rstn), .Q(dout[165]) );
  DFFRHQX1 dout_reg_164_ ( .D(n529), .CK(clk), .RN(rstn), .Q(dout[164]) );
  DFFRHQX1 dout_reg_163_ ( .D(n528), .CK(clk), .RN(rstn), .Q(dout[163]) );
  DFFRHQX1 dout_reg_162_ ( .D(n527), .CK(clk), .RN(rstn), .Q(dout[162]) );
  DFFRHQX1 dout_reg_152_ ( .D(n517), .CK(clk), .RN(rstn), .Q(dout[152]) );
  DFFRHQX1 dout_reg_151_ ( .D(n516), .CK(clk), .RN(rstn), .Q(dout[151]) );
  DFFRHQX1 dout_reg_150_ ( .D(n515), .CK(clk), .RN(rstn), .Q(dout[150]) );
  DFFRHQX1 dout_reg_149_ ( .D(n514), .CK(clk), .RN(rstn), .Q(dout[149]) );
  DFFRHQX1 dout_reg_148_ ( .D(n513), .CK(clk), .RN(rstn), .Q(dout[148]) );
  DFFRHQX1 dout_reg_147_ ( .D(n512), .CK(clk), .RN(rstn), .Q(dout[147]) );
  DFFRHQX1 dout_reg_146_ ( .D(n511), .CK(clk), .RN(rstn), .Q(dout[146]) );
  DFFRHQX1 dout_reg_224_ ( .D(n589), .CK(clk), .RN(rstn), .Q(dout[224]) );
  DFFRHQX1 dout_reg_192_ ( .D(n557), .CK(clk), .RN(rstn), .Q(dout[192]) );
  DFFRHQX1 dout_reg_226_ ( .D(n591), .CK(clk), .RN(rstn), .Q(dout[226]) );
  DFFRHQX1 dout_reg_225_ ( .D(n590), .CK(clk), .RN(rstn), .Q(dout[225]) );
  DFFRHQX1 dout_reg_194_ ( .D(n559), .CK(clk), .RN(rstn), .Q(dout[194]) );
  DFFRHQX1 dout_reg_193_ ( .D(n558), .CK(clk), .RN(rstn), .Q(dout[193]) );
  DFFRHQX1 dout_reg_227_ ( .D(n592), .CK(clk), .RN(rstn), .Q(dout[227]) );
  DFFRHQX1 dout_reg_195_ ( .D(n560), .CK(clk), .RN(rstn), .Q(dout[195]) );
  DFFRHQX1 dout_reg_128_ ( .D(n493), .CK(clk), .RN(rstn), .Q(dout[128]) );
  DFFRHQX1 dout_reg_176_ ( .D(n541), .CK(clk), .RN(rstn), .Q(dout[176]) );
  DFFRHQX1 dout_reg_160_ ( .D(n525), .CK(clk), .RN(rstn), .Q(dout[160]) );
  DFFRHQX1 dout_reg_144_ ( .D(n509), .CK(clk), .RN(rstn), .Q(dout[144]) );
  DFFRHQX1 dout_reg_129_ ( .D(n494), .CK(clk), .RN(rstn), .Q(dout[129]) );
  DFFRHQX1 dout_reg_177_ ( .D(n542), .CK(clk), .RN(rstn), .Q(dout[177]) );
  DFFRHQX1 dout_reg_161_ ( .D(n526), .CK(clk), .RN(rstn), .Q(dout[161]) );
  DFFRHQX1 dout_reg_145_ ( .D(n510), .CK(clk), .RN(rstn), .Q(dout[145]) );
  DFFRHQX1 dout_reg_229_ ( .D(n594), .CK(clk), .RN(rstn), .Q(dout[229]) );
  DFFRHQX1 dout_reg_228_ ( .D(n593), .CK(clk), .RN(rstn), .Q(dout[228]) );
  DFFRHQX1 dout_reg_197_ ( .D(n562), .CK(clk), .RN(rstn), .Q(dout[197]) );
  DFFRHQX1 dout_reg_196_ ( .D(n561), .CK(clk), .RN(rstn), .Q(dout[196]) );
  DFFRHQX1 dout_reg_230_ ( .D(n595), .CK(clk), .RN(rstn), .Q(dout[230]) );
  DFFRHQX1 dout_reg_198_ ( .D(n563), .CK(clk), .RN(rstn), .Q(dout[198]) );
  DFFRHQX1 dout_reg_232_ ( .D(n597), .CK(clk), .RN(rstn), .Q(dout[232]) );
  DFFRHQX1 dout_reg_231_ ( .D(n596), .CK(clk), .RN(rstn), .Q(dout[231]) );
  DFFRHQX1 dout_reg_200_ ( .D(n565), .CK(clk), .RN(rstn), .Q(dout[200]) );
  DFFRHQX1 dout_reg_199_ ( .D(n564), .CK(clk), .RN(rstn), .Q(dout[199]) );
  DFFRHQX1 even_odd_ready_reg ( .D(N275), .CK(clk), .RN(rstn), .Q(
        even_odd_ready) );
  NAND2X1 U3 ( .A(n343), .B(start), .Y(n2) );
  NAND2X1 U4 ( .A(n148), .B(start), .Y(n19) );
  AND2X2 U5 ( .A(n345), .B(start), .Y(n20) );
  AND2X2 U6 ( .A(n344), .B(start), .Y(n149) );
  INVX1 U7 ( .A(n19), .Y(n170) );
  INVX1 U8 ( .A(n19), .Y(n172) );
  INVX1 U9 ( .A(n19), .Y(n173) );
  INVX1 U10 ( .A(n19), .Y(n175) );
  INVX1 U11 ( .A(n188), .Y(n187) );
  INVX1 U12 ( .A(n2), .Y(n176) );
  INVX1 U13 ( .A(n2), .Y(n178) );
  INVX1 U14 ( .A(n2), .Y(n179) );
  INVX1 U15 ( .A(n2), .Y(n181) );
  INVX1 U16 ( .A(start), .Y(n154) );
  INVX1 U17 ( .A(start), .Y(n150) );
  INVX1 U18 ( .A(start), .Y(n151) );
  INVX1 U19 ( .A(start), .Y(n152) );
  INVX1 U20 ( .A(n20), .Y(n166) );
  INVX1 U21 ( .A(n20), .Y(n167) );
  INVX1 U22 ( .A(n20), .Y(n169) );
  INVX1 U23 ( .A(n149), .Y(n164) );
  INVX1 U24 ( .A(n149), .Y(n163) );
  INVX1 U25 ( .A(n149), .Y(n161) );
  INVX1 U26 ( .A(n2), .Y(n182) );
  INVX1 U27 ( .A(n2), .Y(n184) );
  INVX1 U28 ( .A(n2), .Y(n185) );
  INVX1 U29 ( .A(start), .Y(n155) );
  INVX1 U30 ( .A(start), .Y(n157) );
  INVX1 U31 ( .A(start), .Y(n158) );
  INVX1 U32 ( .A(start), .Y(n160) );
  OR2X2 U33 ( .A(n345), .B(n344), .Y(n148) );
  INVX1 U34 ( .A(N275), .Y(n188) );
  AOI2BB1X1 U35 ( .A0N(n343), .A1N(n148), .B0(n154), .Y(N275) );
  NOR2X1 U36 ( .A(mode[0]), .B(mode[1]), .Y(n345) );
  NOR2X1 U37 ( .A(n362), .B(mode[1]), .Y(n344) );
  INVX1 U38 ( .A(mode[0]), .Y(n362) );
  INVX1 U39 ( .A(n18), .Y(n381) );
  AOI222X1 U40 ( .A0(n178), .A1(din[32]), .B0(n170), .B1(din[16]), .C0(n154), 
        .C1(dout[16]), .Y(n18) );
  INVX1 U41 ( .A(n21), .Y(n382) );
  AOI222X1 U42 ( .A0(n181), .A1(din[33]), .B0(n170), .B1(din[17]), .C0(n157), 
        .C1(dout[17]), .Y(n21) );
  INVX1 U43 ( .A(n22), .Y(n383) );
  AOI222X1 U44 ( .A0(n184), .A1(din[34]), .B0(n170), .B1(din[18]), .C0(n154), 
        .C1(dout[18]), .Y(n22) );
  INVX1 U45 ( .A(n23), .Y(n384) );
  AOI222X1 U46 ( .A0(n179), .A1(din[35]), .B0(n170), .B1(din[19]), .C0(n154), 
        .C1(dout[19]), .Y(n23) );
  INVX1 U47 ( .A(n24), .Y(n385) );
  AOI222X1 U48 ( .A0(n176), .A1(din[36]), .B0(n170), .B1(din[20]), .C0(n154), 
        .C1(dout[20]), .Y(n24) );
  INVX1 U49 ( .A(n25), .Y(n386) );
  AOI222X1 U50 ( .A0(n178), .A1(din[37]), .B0(n170), .B1(din[21]), .C0(n154), 
        .C1(dout[21]), .Y(n25) );
  INVX1 U51 ( .A(n26), .Y(n387) );
  AOI222X1 U52 ( .A0(n181), .A1(din[38]), .B0(n170), .B1(din[22]), .C0(n154), 
        .C1(dout[22]), .Y(n26) );
  INVX1 U53 ( .A(n27), .Y(n388) );
  AOI222X1 U54 ( .A0(n179), .A1(din[39]), .B0(n170), .B1(din[23]), .C0(n154), 
        .C1(dout[23]), .Y(n27) );
  INVX1 U55 ( .A(n28), .Y(n389) );
  AOI222X1 U56 ( .A0(n176), .A1(din[40]), .B0(n170), .B1(din[24]), .C0(n154), 
        .C1(dout[24]), .Y(n28) );
  INVX1 U57 ( .A(n29), .Y(n390) );
  AOI222X1 U58 ( .A0(n178), .A1(din[41]), .B0(n170), .B1(din[25]), .C0(n154), 
        .C1(dout[25]), .Y(n29) );
  INVX1 U59 ( .A(n30), .Y(n391) );
  AOI222X1 U60 ( .A0(n181), .A1(din[42]), .B0(n170), .B1(din[26]), .C0(n155), 
        .C1(dout[26]), .Y(n30) );
  INVX1 U61 ( .A(n31), .Y(n392) );
  AOI222X1 U62 ( .A0(n179), .A1(din[43]), .B0(n170), .B1(din[27]), .C0(n155), 
        .C1(dout[27]), .Y(n31) );
  INVX1 U63 ( .A(n32), .Y(n393) );
  AOI222X1 U64 ( .A0(n182), .A1(din[44]), .B0(n172), .B1(din[28]), .C0(n155), 
        .C1(dout[28]), .Y(n32) );
  INVX1 U65 ( .A(n33), .Y(n394) );
  AOI222X1 U66 ( .A0(n182), .A1(din[45]), .B0(n172), .B1(din[29]), .C0(n155), 
        .C1(dout[29]), .Y(n33) );
  INVX1 U67 ( .A(n34), .Y(n395) );
  AOI222X1 U68 ( .A0(n182), .A1(din[46]), .B0(n172), .B1(din[30]), .C0(n155), 
        .C1(dout[30]), .Y(n34) );
  INVX1 U69 ( .A(n35), .Y(n396) );
  AOI222X1 U70 ( .A0(n182), .A1(din[47]), .B0(n172), .B1(din[31]), .C0(n155), 
        .C1(dout[31]), .Y(n35) );
  INVX1 U71 ( .A(n36), .Y(n397) );
  AOI222X1 U72 ( .A0(n182), .A1(din[64]), .B0(n172), .B1(din[32]), .C0(n155), 
        .C1(dout[32]), .Y(n36) );
  INVX1 U73 ( .A(n37), .Y(n398) );
  AOI222X1 U74 ( .A0(n182), .A1(din[65]), .B0(n172), .B1(din[33]), .C0(n155), 
        .C1(dout[33]), .Y(n37) );
  INVX1 U75 ( .A(n38), .Y(n399) );
  AOI222X1 U76 ( .A0(n182), .A1(din[66]), .B0(n172), .B1(din[34]), .C0(n155), 
        .C1(dout[34]), .Y(n38) );
  INVX1 U77 ( .A(n39), .Y(n400) );
  AOI222X1 U78 ( .A0(n182), .A1(din[67]), .B0(n172), .B1(din[35]), .C0(n155), 
        .C1(dout[35]), .Y(n39) );
  INVX1 U79 ( .A(n40), .Y(n401) );
  AOI222X1 U80 ( .A0(n182), .A1(din[68]), .B0(n172), .B1(din[36]), .C0(n155), 
        .C1(dout[36]), .Y(n40) );
  INVX1 U81 ( .A(n41), .Y(n402) );
  AOI222X1 U82 ( .A0(n182), .A1(din[69]), .B0(n172), .B1(din[37]), .C0(n155), 
        .C1(dout[37]), .Y(n41) );
  INVX1 U83 ( .A(n42), .Y(n403) );
  AOI222X1 U84 ( .A0(n182), .A1(din[70]), .B0(n172), .B1(din[38]), .C0(n155), 
        .C1(dout[38]), .Y(n42) );
  INVX1 U85 ( .A(n43), .Y(n404) );
  AOI222X1 U86 ( .A0(n182), .A1(din[71]), .B0(n172), .B1(din[39]), .C0(n155), 
        .C1(dout[39]), .Y(n43) );
  INVX1 U87 ( .A(n140), .Y(n501) );
  AOI222X1 U88 ( .A0(n176), .A1(din[24]), .B0(n172), .B1(din[136]), .C0(n160), 
        .C1(dout[136]), .Y(n140) );
  INVX1 U89 ( .A(n141), .Y(n502) );
  AOI222X1 U90 ( .A0(n178), .A1(din[25]), .B0(n172), .B1(din[137]), .C0(n154), 
        .C1(dout[137]), .Y(n141) );
  INVX1 U91 ( .A(n142), .Y(n503) );
  AOI222X1 U92 ( .A0(n181), .A1(din[26]), .B0(n172), .B1(din[138]), .C0(n154), 
        .C1(dout[138]), .Y(n142) );
  INVX1 U93 ( .A(n143), .Y(n504) );
  AOI222X1 U94 ( .A0(n179), .A1(din[27]), .B0(n170), .B1(din[139]), .C0(n154), 
        .C1(dout[139]), .Y(n143) );
  INVX1 U95 ( .A(n144), .Y(n505) );
  AOI222X1 U96 ( .A0(n176), .A1(din[28]), .B0(n170), .B1(din[140]), .C0(n154), 
        .C1(dout[140]), .Y(n144) );
  INVX1 U97 ( .A(n145), .Y(n506) );
  AOI222X1 U98 ( .A0(n178), .A1(din[29]), .B0(n173), .B1(din[141]), .C0(n154), 
        .C1(dout[141]), .Y(n145) );
  INVX1 U99 ( .A(n146), .Y(n507) );
  AOI222X1 U100 ( .A0(n181), .A1(din[30]), .B0(n175), .B1(din[142]), .C0(n154), 
        .C1(dout[142]), .Y(n146) );
  INVX1 U101 ( .A(n147), .Y(n508) );
  AOI222X1 U102 ( .A0(n179), .A1(din[31]), .B0(n170), .B1(din[143]), .C0(n154), 
        .C1(dout[143]), .Y(n147) );
  INVX1 U103 ( .A(n44), .Y(n405) );
  AOI222X1 U104 ( .A0(n182), .A1(din[72]), .B0(n173), .B1(din[40]), .C0(n155), 
        .C1(dout[40]), .Y(n44) );
  INVX1 U105 ( .A(n45), .Y(n406) );
  AOI222X1 U106 ( .A0(n182), .A1(din[73]), .B0(n173), .B1(din[41]), .C0(n155), 
        .C1(dout[41]), .Y(n45) );
  INVX1 U107 ( .A(n46), .Y(n407) );
  AOI222X1 U108 ( .A0(n182), .A1(din[74]), .B0(n173), .B1(din[42]), .C0(n155), 
        .C1(dout[42]), .Y(n46) );
  INVX1 U109 ( .A(n47), .Y(n408) );
  AOI222X1 U110 ( .A0(n182), .A1(din[75]), .B0(n173), .B1(din[43]), .C0(n155), 
        .C1(dout[43]), .Y(n47) );
  INVX1 U111 ( .A(n48), .Y(n409) );
  AOI222X1 U112 ( .A0(n182), .A1(din[76]), .B0(n173), .B1(din[44]), .C0(n155), 
        .C1(dout[44]), .Y(n48) );
  INVX1 U113 ( .A(n49), .Y(n410) );
  AOI222X1 U114 ( .A0(n182), .A1(din[77]), .B0(n173), .B1(din[45]), .C0(n155), 
        .C1(dout[45]), .Y(n49) );
  INVX1 U115 ( .A(n50), .Y(n411) );
  AOI222X1 U116 ( .A0(n182), .A1(din[78]), .B0(n173), .B1(din[46]), .C0(n155), 
        .C1(dout[46]), .Y(n50) );
  INVX1 U117 ( .A(n51), .Y(n412) );
  AOI222X1 U118 ( .A0(n182), .A1(din[79]), .B0(n173), .B1(din[47]), .C0(n155), 
        .C1(dout[47]), .Y(n51) );
  INVX1 U119 ( .A(n68), .Y(n429) );
  AOI222X1 U120 ( .A0(n184), .A1(din[128]), .B0(n175), .B1(din[64]), .C0(n154), 
        .C1(dout[64]), .Y(n68) );
  INVX1 U121 ( .A(n69), .Y(n430) );
  AOI222X1 U122 ( .A0(n184), .A1(din[129]), .B0(n175), .B1(din[65]), .C0(n157), 
        .C1(dout[65]), .Y(n69) );
  INVX1 U123 ( .A(n70), .Y(n431) );
  AOI222X1 U124 ( .A0(n184), .A1(din[130]), .B0(n175), .B1(din[66]), .C0(n157), 
        .C1(dout[66]), .Y(n70) );
  INVX1 U125 ( .A(n71), .Y(n432) );
  AOI222X1 U126 ( .A0(n184), .A1(din[131]), .B0(n175), .B1(din[67]), .C0(n157), 
        .C1(dout[67]), .Y(n71) );
  INVX1 U127 ( .A(n72), .Y(n433) );
  AOI222X1 U128 ( .A0(n184), .A1(din[132]), .B0(n175), .B1(din[68]), .C0(n157), 
        .C1(dout[68]), .Y(n72) );
  INVX1 U129 ( .A(n73), .Y(n434) );
  AOI222X1 U130 ( .A0(n184), .A1(din[133]), .B0(n175), .B1(din[69]), .C0(n157), 
        .C1(dout[69]), .Y(n73) );
  INVX1 U131 ( .A(n74), .Y(n435) );
  AOI222X1 U132 ( .A0(n184), .A1(din[134]), .B0(n175), .B1(din[70]), .C0(n157), 
        .C1(dout[70]), .Y(n74) );
  INVX1 U133 ( .A(n75), .Y(n436) );
  AOI222X1 U134 ( .A0(n184), .A1(din[135]), .B0(n175), .B1(din[71]), .C0(n157), 
        .C1(dout[71]), .Y(n75) );
  INVX1 U135 ( .A(n76), .Y(n437) );
  AOI222X1 U136 ( .A0(n184), .A1(din[136]), .B0(n175), .B1(din[72]), .C0(n157), 
        .C1(dout[72]), .Y(n76) );
  INVX1 U137 ( .A(n77), .Y(n438) );
  AOI222X1 U138 ( .A0(n184), .A1(din[137]), .B0(n175), .B1(din[73]), .C0(n157), 
        .C1(dout[73]), .Y(n77) );
  INVX1 U139 ( .A(n78), .Y(n439) );
  AOI222X1 U140 ( .A0(n184), .A1(din[138]), .B0(n175), .B1(din[74]), .C0(n157), 
        .C1(dout[74]), .Y(n78) );
  INVX1 U141 ( .A(n79), .Y(n440) );
  AOI222X1 U142 ( .A0(n184), .A1(din[139]), .B0(n175), .B1(din[75]), .C0(n157), 
        .C1(dout[75]), .Y(n79) );
  INVX1 U143 ( .A(n80), .Y(n441) );
  AOI222X1 U144 ( .A0(n184), .A1(din[140]), .B0(n173), .B1(din[76]), .C0(n157), 
        .C1(dout[76]), .Y(n80) );
  INVX1 U145 ( .A(n81), .Y(n442) );
  AOI222X1 U146 ( .A0(n184), .A1(din[141]), .B0(n170), .B1(din[77]), .C0(n157), 
        .C1(dout[77]), .Y(n81) );
  INVX1 U147 ( .A(n82), .Y(n443) );
  AOI222X1 U148 ( .A0(n184), .A1(din[142]), .B0(n170), .B1(din[78]), .C0(n157), 
        .C1(dout[78]), .Y(n82) );
  INVX1 U149 ( .A(n83), .Y(n444) );
  AOI222X1 U150 ( .A0(n184), .A1(din[143]), .B0(n175), .B1(din[79]), .C0(n157), 
        .C1(dout[79]), .Y(n83) );
  INVX1 U151 ( .A(n100), .Y(n461) );
  AOI222X1 U152 ( .A0(n185), .A1(din[192]), .B0(n170), .B1(din[96]), .C0(n158), 
        .C1(dout[96]), .Y(n100) );
  INVX1 U153 ( .A(n101), .Y(n462) );
  AOI222X1 U154 ( .A0(n185), .A1(din[193]), .B0(n173), .B1(din[97]), .C0(n158), 
        .C1(dout[97]), .Y(n101) );
  INVX1 U155 ( .A(n102), .Y(n463) );
  AOI222X1 U156 ( .A0(n185), .A1(din[194]), .B0(n172), .B1(din[98]), .C0(n158), 
        .C1(dout[98]), .Y(n102) );
  INVX1 U157 ( .A(n103), .Y(n464) );
  AOI222X1 U158 ( .A0(n185), .A1(din[195]), .B0(n173), .B1(din[99]), .C0(n158), 
        .C1(dout[99]), .Y(n103) );
  INVX1 U159 ( .A(n104), .Y(n465) );
  AOI222X1 U160 ( .A0(n185), .A1(din[196]), .B0(n173), .B1(din[100]), .C0(n158), .C1(dout[100]), .Y(n104) );
  INVX1 U161 ( .A(n105), .Y(n466) );
  AOI222X1 U162 ( .A0(n185), .A1(din[197]), .B0(n173), .B1(din[101]), .C0(n158), .C1(dout[101]), .Y(n105) );
  INVX1 U163 ( .A(n106), .Y(n467) );
  AOI222X1 U164 ( .A0(n185), .A1(din[198]), .B0(n172), .B1(din[102]), .C0(n158), .C1(dout[102]), .Y(n106) );
  INVX1 U165 ( .A(n107), .Y(n468) );
  AOI222X1 U166 ( .A0(n185), .A1(din[199]), .B0(n170), .B1(din[103]), .C0(n158), .C1(dout[103]), .Y(n107) );
  INVX1 U167 ( .A(n108), .Y(n469) );
  AOI222X1 U168 ( .A0(n185), .A1(din[200]), .B0(n175), .B1(din[104]), .C0(n158), .C1(dout[104]), .Y(n108) );
  INVX1 U169 ( .A(n109), .Y(n470) );
  AOI222X1 U170 ( .A0(n185), .A1(din[201]), .B0(n173), .B1(din[105]), .C0(n158), .C1(dout[105]), .Y(n109) );
  INVX1 U171 ( .A(n110), .Y(n471) );
  AOI222X1 U172 ( .A0(n185), .A1(din[202]), .B0(n173), .B1(din[106]), .C0(n158), .C1(dout[106]), .Y(n110) );
  INVX1 U173 ( .A(n111), .Y(n472) );
  AOI222X1 U174 ( .A0(n185), .A1(din[203]), .B0(n172), .B1(din[107]), .C0(n158), .C1(dout[107]), .Y(n111) );
  INVX1 U175 ( .A(n112), .Y(n473) );
  AOI222X1 U176 ( .A0(n185), .A1(din[204]), .B0(n170), .B1(din[108]), .C0(n158), .C1(dout[108]), .Y(n112) );
  INVX1 U177 ( .A(n113), .Y(n474) );
  AOI222X1 U178 ( .A0(n185), .A1(din[205]), .B0(n175), .B1(din[109]), .C0(n158), .C1(dout[109]), .Y(n113) );
  INVX1 U179 ( .A(n114), .Y(n475) );
  AOI222X1 U180 ( .A0(n185), .A1(din[206]), .B0(n173), .B1(din[110]), .C0(n158), .C1(dout[110]), .Y(n114) );
  INVX1 U181 ( .A(n115), .Y(n476) );
  AOI222X1 U182 ( .A0(n185), .A1(din[207]), .B0(n172), .B1(din[111]), .C0(n158), .C1(dout[111]), .Y(n115) );
  INVX1 U183 ( .A(n132), .Y(n493) );
  AOI222X1 U184 ( .A0(din[16]), .A1(n176), .B0(n175), .B1(din[128]), .C0(n160), 
        .C1(dout[128]), .Y(n132) );
  INVX1 U185 ( .A(n133), .Y(n494) );
  AOI222X1 U186 ( .A0(n179), .A1(din[17]), .B0(n175), .B1(din[129]), .C0(n160), 
        .C1(dout[129]), .Y(n133) );
  INVX1 U187 ( .A(n134), .Y(n495) );
  AOI222X1 U188 ( .A0(n176), .A1(din[18]), .B0(n172), .B1(din[130]), .C0(n160), 
        .C1(dout[130]), .Y(n134) );
  INVX1 U189 ( .A(n135), .Y(n496) );
  AOI222X1 U190 ( .A0(n178), .A1(din[19]), .B0(n173), .B1(din[131]), .C0(n160), 
        .C1(dout[131]), .Y(n135) );
  INVX1 U191 ( .A(n136), .Y(n497) );
  AOI222X1 U192 ( .A0(n181), .A1(din[20]), .B0(n172), .B1(din[132]), .C0(n160), 
        .C1(dout[132]), .Y(n136) );
  INVX1 U193 ( .A(n137), .Y(n498) );
  AOI222X1 U194 ( .A0(n179), .A1(din[21]), .B0(n175), .B1(din[133]), .C0(n160), 
        .C1(dout[133]), .Y(n137) );
  INVX1 U195 ( .A(n138), .Y(n499) );
  AOI222X1 U196 ( .A0(n176), .A1(din[22]), .B0(n170), .B1(din[134]), .C0(n160), 
        .C1(dout[134]), .Y(n138) );
  INVX1 U197 ( .A(n139), .Y(n500) );
  AOI222X1 U198 ( .A0(n178), .A1(din[23]), .B0(n173), .B1(din[135]), .C0(n160), 
        .C1(dout[135]), .Y(n139) );
  INVX1 U199 ( .A(n52), .Y(n413) );
  AOI222X1 U200 ( .A0(n182), .A1(din[96]), .B0(n173), .B1(din[48]), .C0(n155), 
        .C1(dout[48]), .Y(n52) );
  INVX1 U201 ( .A(n53), .Y(n414) );
  AOI222X1 U202 ( .A0(n182), .A1(din[97]), .B0(n173), .B1(din[49]), .C0(n155), 
        .C1(dout[49]), .Y(n53) );
  INVX1 U203 ( .A(n54), .Y(n415) );
  AOI222X1 U204 ( .A0(n182), .A1(din[98]), .B0(n173), .B1(din[50]), .C0(n155), 
        .C1(dout[50]), .Y(n54) );
  INVX1 U205 ( .A(n55), .Y(n416) );
  AOI222X1 U206 ( .A0(n182), .A1(din[99]), .B0(n173), .B1(din[51]), .C0(n155), 
        .C1(dout[51]), .Y(n55) );
  INVX1 U207 ( .A(n56), .Y(n417) );
  AOI222X1 U208 ( .A0(n182), .A1(din[100]), .B0(n172), .B1(din[52]), .C0(n155), 
        .C1(dout[52]), .Y(n56) );
  INVX1 U209 ( .A(n57), .Y(n418) );
  AOI222X1 U210 ( .A0(n182), .A1(din[101]), .B0(n175), .B1(din[53]), .C0(n155), 
        .C1(dout[53]), .Y(n57) );
  INVX1 U211 ( .A(n58), .Y(n419) );
  AOI222X1 U212 ( .A0(n182), .A1(din[102]), .B0(n170), .B1(din[54]), .C0(n155), 
        .C1(dout[54]), .Y(n58) );
  INVX1 U213 ( .A(n59), .Y(n420) );
  AOI222X1 U214 ( .A0(n182), .A1(din[103]), .B0(n173), .B1(din[55]), .C0(n155), 
        .C1(dout[55]), .Y(n59) );
  INVX1 U215 ( .A(n60), .Y(n421) );
  AOI222X1 U216 ( .A0(n182), .A1(din[104]), .B0(n172), .B1(din[56]), .C0(n155), 
        .C1(dout[56]), .Y(n60) );
  INVX1 U217 ( .A(n61), .Y(n422) );
  AOI222X1 U218 ( .A0(n182), .A1(din[105]), .B0(n175), .B1(din[57]), .C0(n155), 
        .C1(dout[57]), .Y(n61) );
  INVX1 U219 ( .A(n62), .Y(n423) );
  AOI222X1 U220 ( .A0(n182), .A1(din[106]), .B0(n170), .B1(din[58]), .C0(n157), 
        .C1(dout[58]), .Y(n62) );
  INVX1 U221 ( .A(n63), .Y(n424) );
  AOI222X1 U222 ( .A0(n182), .A1(din[107]), .B0(n173), .B1(din[59]), .C0(n157), 
        .C1(dout[59]), .Y(n63) );
  INVX1 U223 ( .A(n64), .Y(n425) );
  AOI222X1 U224 ( .A0(n184), .A1(din[108]), .B0(n172), .B1(din[60]), .C0(n157), 
        .C1(dout[60]), .Y(n64) );
  INVX1 U225 ( .A(n65), .Y(n426) );
  AOI222X1 U226 ( .A0(n184), .A1(din[109]), .B0(n175), .B1(din[61]), .C0(n157), 
        .C1(dout[61]), .Y(n65) );
  INVX1 U227 ( .A(n66), .Y(n427) );
  AOI222X1 U228 ( .A0(n184), .A1(din[110]), .B0(n170), .B1(din[62]), .C0(n157), 
        .C1(dout[62]), .Y(n66) );
  INVX1 U229 ( .A(n67), .Y(n428) );
  AOI222X1 U230 ( .A0(n184), .A1(din[111]), .B0(n173), .B1(din[63]), .C0(n157), 
        .C1(dout[63]), .Y(n67) );
  INVX1 U231 ( .A(n84), .Y(n445) );
  AOI222X1 U232 ( .A0(n184), .A1(din[160]), .B0(n172), .B1(din[80]), .C0(n157), 
        .C1(dout[80]), .Y(n84) );
  INVX1 U233 ( .A(n85), .Y(n446) );
  AOI222X1 U234 ( .A0(n184), .A1(din[161]), .B0(n172), .B1(din[81]), .C0(n157), 
        .C1(dout[81]), .Y(n85) );
  INVX1 U235 ( .A(n86), .Y(n447) );
  AOI222X1 U236 ( .A0(n184), .A1(din[162]), .B0(n173), .B1(din[82]), .C0(n157), 
        .C1(dout[82]), .Y(n86) );
  INVX1 U237 ( .A(n87), .Y(n448) );
  AOI222X1 U238 ( .A0(n184), .A1(din[163]), .B0(n173), .B1(din[83]), .C0(n157), 
        .C1(dout[83]), .Y(n87) );
  INVX1 U239 ( .A(n88), .Y(n449) );
  AOI222X1 U240 ( .A0(n184), .A1(din[164]), .B0(n170), .B1(din[84]), .C0(n157), 
        .C1(dout[84]), .Y(n88) );
  INVX1 U241 ( .A(n89), .Y(n450) );
  AOI222X1 U242 ( .A0(n184), .A1(din[165]), .B0(n175), .B1(din[85]), .C0(n157), 
        .C1(dout[85]), .Y(n89) );
  INVX1 U243 ( .A(n90), .Y(n451) );
  AOI222X1 U244 ( .A0(n184), .A1(din[166]), .B0(n172), .B1(din[86]), .C0(n157), 
        .C1(dout[86]), .Y(n90) );
  INVX1 U245 ( .A(n91), .Y(n452) );
  AOI222X1 U246 ( .A0(n184), .A1(din[167]), .B0(n170), .B1(din[87]), .C0(n157), 
        .C1(dout[87]), .Y(n91) );
  INVX1 U247 ( .A(n92), .Y(n453) );
  AOI222X1 U248 ( .A0(n184), .A1(din[168]), .B0(n175), .B1(din[88]), .C0(n157), 
        .C1(dout[88]), .Y(n92) );
  INVX1 U249 ( .A(n93), .Y(n454) );
  AOI222X1 U250 ( .A0(n184), .A1(din[169]), .B0(n172), .B1(din[89]), .C0(n157), 
        .C1(dout[89]), .Y(n93) );
  INVX1 U251 ( .A(n94), .Y(n455) );
  AOI222X1 U252 ( .A0(n184), .A1(din[170]), .B0(n172), .B1(din[90]), .C0(n158), 
        .C1(dout[90]), .Y(n94) );
  INVX1 U253 ( .A(n95), .Y(n456) );
  AOI222X1 U254 ( .A0(n185), .A1(din[171]), .B0(n170), .B1(din[91]), .C0(n158), 
        .C1(dout[91]), .Y(n95) );
  INVX1 U255 ( .A(n96), .Y(n457) );
  AOI222X1 U256 ( .A0(n185), .A1(din[172]), .B0(n173), .B1(din[92]), .C0(n158), 
        .C1(dout[92]), .Y(n96) );
  INVX1 U257 ( .A(n97), .Y(n458) );
  AOI222X1 U258 ( .A0(n185), .A1(din[173]), .B0(n175), .B1(din[93]), .C0(n158), 
        .C1(dout[93]), .Y(n97) );
  INVX1 U259 ( .A(n98), .Y(n459) );
  AOI222X1 U260 ( .A0(n185), .A1(din[174]), .B0(n175), .B1(din[94]), .C0(n158), 
        .C1(dout[94]), .Y(n98) );
  INVX1 U261 ( .A(n99), .Y(n460) );
  AOI222X1 U262 ( .A0(n185), .A1(din[175]), .B0(n175), .B1(din[95]), .C0(n158), 
        .C1(dout[95]), .Y(n99) );
  INVX1 U263 ( .A(n116), .Y(n477) );
  AOI222X1 U264 ( .A0(n185), .A1(din[224]), .B0(n172), .B1(din[112]), .C0(n158), .C1(dout[112]), .Y(n116) );
  INVX1 U265 ( .A(n117), .Y(n478) );
  AOI222X1 U266 ( .A0(n185), .A1(din[225]), .B0(n170), .B1(din[113]), .C0(n158), .C1(dout[113]), .Y(n117) );
  INVX1 U267 ( .A(n118), .Y(n479) );
  AOI222X1 U268 ( .A0(n185), .A1(din[226]), .B0(n170), .B1(din[114]), .C0(n158), .C1(dout[114]), .Y(n118) );
  INVX1 U269 ( .A(n119), .Y(n480) );
  AOI222X1 U270 ( .A0(n185), .A1(din[227]), .B0(n173), .B1(din[115]), .C0(n158), .C1(dout[115]), .Y(n119) );
  INVX1 U271 ( .A(n120), .Y(n481) );
  AOI222X1 U272 ( .A0(n185), .A1(din[228]), .B0(n170), .B1(din[116]), .C0(n158), .C1(dout[116]), .Y(n120) );
  INVX1 U273 ( .A(n121), .Y(n482) );
  AOI222X1 U274 ( .A0(n185), .A1(din[229]), .B0(n175), .B1(din[117]), .C0(n158), .C1(dout[117]), .Y(n121) );
  INVX1 U275 ( .A(n122), .Y(n483) );
  AOI222X1 U276 ( .A0(n185), .A1(din[230]), .B0(n175), .B1(din[118]), .C0(n158), .C1(dout[118]), .Y(n122) );
  INVX1 U277 ( .A(n123), .Y(n484) );
  AOI222X1 U278 ( .A0(n185), .A1(din[231]), .B0(n170), .B1(din[119]), .C0(n158), .C1(dout[119]), .Y(n123) );
  INVX1 U279 ( .A(n124), .Y(n485) );
  AOI222X1 U280 ( .A0(n185), .A1(din[232]), .B0(n173), .B1(din[120]), .C0(n158), .C1(dout[120]), .Y(n124) );
  INVX1 U281 ( .A(n125), .Y(n486) );
  AOI222X1 U282 ( .A0(n185), .A1(din[233]), .B0(n173), .B1(din[121]), .C0(n158), .C1(dout[121]), .Y(n125) );
  INVX1 U283 ( .A(n126), .Y(n487) );
  AOI222X1 U284 ( .A0(n185), .A1(din[234]), .B0(n175), .B1(din[122]), .C0(n160), .C1(dout[122]), .Y(n126) );
  INVX1 U285 ( .A(n127), .Y(n488) );
  AOI222X1 U286 ( .A0(n176), .A1(din[235]), .B0(n175), .B1(din[123]), .C0(n160), .C1(dout[123]), .Y(n127) );
  INVX1 U287 ( .A(n128), .Y(n489) );
  AOI222X1 U288 ( .A0(n179), .A1(din[236]), .B0(n170), .B1(din[124]), .C0(n160), .C1(dout[124]), .Y(n128) );
  INVX1 U289 ( .A(n129), .Y(n490) );
  AOI222X1 U290 ( .A0(n181), .A1(din[237]), .B0(n172), .B1(din[125]), .C0(n160), .C1(dout[125]), .Y(n129) );
  INVX1 U291 ( .A(n130), .Y(n491) );
  AOI222X1 U292 ( .A0(n178), .A1(din[238]), .B0(n175), .B1(din[126]), .C0(n160), .C1(dout[126]), .Y(n130) );
  INVX1 U293 ( .A(n131), .Y(n492) );
  AOI222X1 U294 ( .A0(n178), .A1(din[239]), .B0(n172), .B1(din[127]), .C0(n160), .C1(dout[127]), .Y(n131) );
  OAI221XL U295 ( .A0(n646), .A1(n167), .B0(n161), .B1(n265), .C0(n280), .Y(
        n558) );
  AOI22X1 U296 ( .A0(din[49]), .A1(n179), .B0(dout[193]), .B1(n151), .Y(n280)
         );
  OAI221XL U297 ( .A0(n643), .A1(n169), .B0(n161), .B1(n261), .C0(n281), .Y(
        n559) );
  AOI22X1 U298 ( .A0(din[50]), .A1(n181), .B0(dout[194]), .B1(n150), .Y(n281)
         );
  OAI221XL U299 ( .A0(n640), .A1(n169), .B0(n164), .B1(n256), .C0(n282), .Y(
        n560) );
  AOI22X1 U300 ( .A0(din[51]), .A1(n178), .B0(dout[195]), .B1(n160), .Y(n282)
         );
  OAI221XL U301 ( .A0(n637), .A1(n166), .B0(n163), .B1(n252), .C0(n283), .Y(
        n561) );
  AOI22X1 U302 ( .A0(din[52]), .A1(n178), .B0(dout[196]), .B1(n151), .Y(n283)
         );
  OAI221XL U303 ( .A0(n634), .A1(n169), .B0(n164), .B1(n247), .C0(n284), .Y(
        n562) );
  AOI22X1 U304 ( .A0(din[53]), .A1(n178), .B0(dout[197]), .B1(n152), .Y(n284)
         );
  OAI221XL U305 ( .A0(n631), .A1(n169), .B0(n161), .B1(n243), .C0(n285), .Y(
        n563) );
  AOI22X1 U306 ( .A0(din[54]), .A1(n178), .B0(dout[198]), .B1(n151), .Y(n285)
         );
  OAI221XL U307 ( .A0(n628), .A1(n169), .B0(n164), .B1(n238), .C0(n286), .Y(
        n564) );
  AOI22X1 U308 ( .A0(din[55]), .A1(n178), .B0(dout[199]), .B1(n150), .Y(n286)
         );
  OAI221XL U309 ( .A0(n625), .A1(n167), .B0(n163), .B1(n234), .C0(n287), .Y(
        n565) );
  AOI22X1 U310 ( .A0(din[56]), .A1(n178), .B0(dout[200]), .B1(n160), .Y(n287)
         );
  OAI221XL U311 ( .A0(n325), .A1(n169), .B0(n164), .B1(n229), .C0(n288), .Y(
        n566) );
  AOI22X1 U312 ( .A0(din[57]), .A1(n178), .B0(dout[201]), .B1(n160), .Y(n288)
         );
  OAI221XL U313 ( .A0(n319), .A1(n166), .B0(n164), .B1(n223), .C0(n289), .Y(
        n567) );
  AOI22X1 U314 ( .A0(din[58]), .A1(n178), .B0(dout[202]), .B1(n160), .Y(n289)
         );
  OAI221XL U315 ( .A0(n313), .A1(n167), .B0(n164), .B1(n217), .C0(n290), .Y(
        n568) );
  AOI22X1 U316 ( .A0(din[59]), .A1(n178), .B0(dout[203]), .B1(n152), .Y(n290)
         );
  OAI221XL U317 ( .A0(n307), .A1(n169), .B0(n164), .B1(n211), .C0(n291), .Y(
        n569) );
  AOI22X1 U318 ( .A0(din[60]), .A1(n178), .B0(dout[204]), .B1(n151), .Y(n291)
         );
  OAI221XL U319 ( .A0(n301), .A1(n169), .B0(n164), .B1(n205), .C0(n292), .Y(
        n570) );
  AOI22X1 U320 ( .A0(din[61]), .A1(n178), .B0(dout[205]), .B1(n151), .Y(n292)
         );
  OAI221XL U321 ( .A0(n295), .A1(n169), .B0(n164), .B1(n199), .C0(n293), .Y(
        n571) );
  AOI22X1 U322 ( .A0(din[62]), .A1(n178), .B0(dout[206]), .B1(n151), .Y(n293)
         );
  OAI221XL U323 ( .A0(n274), .A1(n169), .B0(n164), .B1(n194), .C0(n294), .Y(
        n572) );
  AOI22X1 U324 ( .A0(din[63]), .A1(n178), .B0(dout[207]), .B1(n151), .Y(n294)
         );
  OAI221XL U325 ( .A0(n167), .A1(n648), .B0(n164), .B1(n267), .C0(n296), .Y(
        n573) );
  AOI22X1 U326 ( .A0(din[112]), .A1(n179), .B0(dout[208]), .B1(n151), .Y(n296)
         );
  OAI221XL U327 ( .A0(n169), .A1(n645), .B0(n164), .B1(n262), .C0(n298), .Y(
        n574) );
  AOI22X1 U328 ( .A0(din[113]), .A1(n179), .B0(dout[209]), .B1(n151), .Y(n298)
         );
  OAI221XL U329 ( .A0(n166), .A1(n642), .B0(n164), .B1(n258), .C0(n300), .Y(
        n575) );
  AOI22X1 U330 ( .A0(din[114]), .A1(n179), .B0(dout[210]), .B1(n151), .Y(n300)
         );
  OAI221XL U331 ( .A0(n167), .A1(n639), .B0(n164), .B1(n253), .C0(n302), .Y(
        n576) );
  AOI22X1 U332 ( .A0(din[115]), .A1(n179), .B0(dout[211]), .B1(n151), .Y(n302)
         );
  OAI221XL U333 ( .A0(n166), .A1(n636), .B0(n164), .B1(n249), .C0(n304), .Y(
        n577) );
  AOI22X1 U334 ( .A0(din[116]), .A1(n179), .B0(dout[212]), .B1(n151), .Y(n304)
         );
  OAI221XL U335 ( .A0(n167), .A1(n633), .B0(n164), .B1(n244), .C0(n306), .Y(
        n578) );
  AOI22X1 U336 ( .A0(din[117]), .A1(n179), .B0(dout[213]), .B1(n151), .Y(n306)
         );
  OAI221XL U337 ( .A0(n169), .A1(n630), .B0(n163), .B1(n240), .C0(n308), .Y(
        n579) );
  AOI22X1 U338 ( .A0(din[118]), .A1(n179), .B0(dout[214]), .B1(n152), .Y(n308)
         );
  OAI221XL U339 ( .A0(n169), .A1(n627), .B0(n163), .B1(n235), .C0(n310), .Y(
        n580) );
  AOI22X1 U340 ( .A0(din[119]), .A1(n179), .B0(dout[215]), .B1(n152), .Y(n310)
         );
  OAI221XL U341 ( .A0(n167), .A1(n624), .B0(n163), .B1(n231), .C0(n312), .Y(
        n581) );
  AOI22X1 U342 ( .A0(din[120]), .A1(n179), .B0(dout[216]), .B1(n152), .Y(n312)
         );
  OAI221XL U343 ( .A0(n166), .A1(n323), .B0(n163), .B1(n225), .C0(n314), .Y(
        n582) );
  AOI22X1 U344 ( .A0(din[121]), .A1(n179), .B0(dout[217]), .B1(n152), .Y(n314)
         );
  OAI221XL U345 ( .A0(n167), .A1(n317), .B0(n163), .B1(n219), .C0(n316), .Y(
        n583) );
  AOI22X1 U346 ( .A0(din[122]), .A1(n179), .B0(dout[218]), .B1(n152), .Y(n316)
         );
  OAI221XL U347 ( .A0(n169), .A1(n311), .B0(n163), .B1(n213), .C0(n318), .Y(
        n584) );
  AOI22X1 U348 ( .A0(din[123]), .A1(n179), .B0(dout[219]), .B1(n152), .Y(n318)
         );
  OAI221XL U349 ( .A0(n169), .A1(n305), .B0(n163), .B1(n207), .C0(n320), .Y(
        n585) );
  AOI22X1 U350 ( .A0(din[124]), .A1(n179), .B0(dout[220]), .B1(n152), .Y(n320)
         );
  OAI221XL U351 ( .A0(n166), .A1(n299), .B0(n163), .B1(n201), .C0(n322), .Y(
        n586) );
  AOI22X1 U352 ( .A0(din[125]), .A1(n181), .B0(dout[221]), .B1(n152), .Y(n322)
         );
  OAI221XL U353 ( .A0(n166), .A1(n277), .B0(n163), .B1(n196), .C0(n324), .Y(
        n587) );
  AOI22X1 U354 ( .A0(din[126]), .A1(n181), .B0(dout[222]), .B1(n151), .Y(n324)
         );
  OAI221XL U355 ( .A0(n167), .A1(n273), .B0(n163), .B1(n191), .C0(n326), .Y(
        n588) );
  AOI22X1 U356 ( .A0(din[127]), .A1(n181), .B0(dout[223]), .B1(n152), .Y(n326)
         );
  OAI221XL U357 ( .A0(n647), .A1(n169), .B0(n163), .B1(n648), .C0(n327), .Y(
        n589) );
  AOI22X1 U358 ( .A0(din[176]), .A1(n181), .B0(dout[224]), .B1(n152), .Y(n327)
         );
  OAI221XL U359 ( .A0(n644), .A1(n167), .B0(n163), .B1(n645), .C0(n328), .Y(
        n590) );
  AOI22X1 U360 ( .A0(din[177]), .A1(n181), .B0(dout[225]), .B1(n152), .Y(n328)
         );
  OAI221XL U361 ( .A0(n641), .A1(n167), .B0(n163), .B1(n642), .C0(n329), .Y(
        n591) );
  AOI22X1 U362 ( .A0(din[178]), .A1(n181), .B0(dout[226]), .B1(n151), .Y(n329)
         );
  OAI221XL U363 ( .A0(n638), .A1(n166), .B0(n161), .B1(n639), .C0(n330), .Y(
        n592) );
  AOI22X1 U364 ( .A0(din[179]), .A1(n181), .B0(dout[227]), .B1(n151), .Y(n330)
         );
  OAI221XL U365 ( .A0(n635), .A1(n169), .B0(n161), .B1(n636), .C0(n331), .Y(
        n593) );
  AOI22X1 U366 ( .A0(din[180]), .A1(n181), .B0(dout[228]), .B1(n151), .Y(n331)
         );
  OAI221XL U367 ( .A0(n632), .A1(n166), .B0(n161), .B1(n633), .C0(n332), .Y(
        n594) );
  AOI22X1 U368 ( .A0(din[181]), .A1(n181), .B0(dout[229]), .B1(n152), .Y(n332)
         );
  OAI221XL U369 ( .A0(n629), .A1(n167), .B0(n161), .B1(n630), .C0(n333), .Y(
        n595) );
  AOI22X1 U370 ( .A0(din[182]), .A1(n181), .B0(dout[230]), .B1(n150), .Y(n333)
         );
  OAI221XL U371 ( .A0(n626), .A1(n166), .B0(n161), .B1(n627), .C0(n334), .Y(
        n596) );
  AOI22X1 U372 ( .A0(din[183]), .A1(n181), .B0(dout[231]), .B1(n150), .Y(n334)
         );
  OAI221XL U373 ( .A0(n623), .A1(n169), .B0(n161), .B1(n624), .C0(n335), .Y(
        n597) );
  AOI22X1 U374 ( .A0(din[184]), .A1(n181), .B0(dout[232]), .B1(n151), .Y(n335)
         );
  OAI221XL U375 ( .A0(n321), .A1(n169), .B0(n161), .B1(n323), .C0(n336), .Y(
        n598) );
  AOI22X1 U376 ( .A0(din[185]), .A1(n181), .B0(dout[233]), .B1(n151), .Y(n336)
         );
  OAI221XL U377 ( .A0(n315), .A1(n167), .B0(n161), .B1(n317), .C0(n337), .Y(
        n599) );
  AOI22X1 U378 ( .A0(din[186]), .A1(n176), .B0(dout[234]), .B1(n150), .Y(n337)
         );
  OAI221XL U379 ( .A0(n309), .A1(n169), .B0(n161), .B1(n311), .C0(n338), .Y(
        n600) );
  AOI22X1 U380 ( .A0(din[187]), .A1(n181), .B0(dout[235]), .B1(n152), .Y(n338)
         );
  OAI221XL U381 ( .A0(n303), .A1(n169), .B0(n161), .B1(n305), .C0(n339), .Y(
        n601) );
  AOI22X1 U382 ( .A0(din[188]), .A1(n178), .B0(dout[236]), .B1(n152), .Y(n339)
         );
  OAI221XL U383 ( .A0(n297), .A1(n167), .B0(n161), .B1(n299), .C0(n340), .Y(
        n602) );
  AOI22X1 U384 ( .A0(din[189]), .A1(n179), .B0(dout[237]), .B1(n150), .Y(n340)
         );
  OAI221XL U385 ( .A0(n276), .A1(n169), .B0(n161), .B1(n277), .C0(n341), .Y(
        n603) );
  AOI22X1 U386 ( .A0(din[190]), .A1(n181), .B0(dout[238]), .B1(n152), .Y(n341)
         );
  OAI221XL U387 ( .A0(n271), .A1(n169), .B0(n161), .B1(n273), .C0(n342), .Y(
        n604) );
  AOI22X1 U388 ( .A0(din[191]), .A1(n179), .B0(dout[239]), .B1(n152), .Y(n342)
         );
  OAI221XL U389 ( .A0(n169), .A1(n270), .B0(n268), .B1(n164), .C0(n153), .Y(
        n509) );
  AOI22X1 U390 ( .A0(din[80]), .A1(n176), .B0(dout[144]), .B1(n150), .Y(n153)
         );
  OAI221XL U391 ( .A0(n166), .A1(n265), .B0(n264), .B1(n161), .C0(n156), .Y(
        n510) );
  AOI22X1 U392 ( .A0(din[81]), .A1(n176), .B0(dout[145]), .B1(n150), .Y(n156)
         );
  OAI221XL U393 ( .A0(n167), .A1(n261), .B0(n259), .B1(n163), .C0(n159), .Y(
        n511) );
  AOI22X1 U394 ( .A0(din[82]), .A1(n176), .B0(dout[146]), .B1(n150), .Y(n159)
         );
  OAI221XL U395 ( .A0(n167), .A1(n256), .B0(n255), .B1(n164), .C0(n162), .Y(
        n512) );
  AOI22X1 U396 ( .A0(din[83]), .A1(n176), .B0(dout[147]), .B1(n160), .Y(n162)
         );
  OAI221XL U397 ( .A0(n167), .A1(n252), .B0(n250), .B1(n161), .C0(n165), .Y(
        n513) );
  AOI22X1 U398 ( .A0(din[84]), .A1(n176), .B0(dout[148]), .B1(n151), .Y(n165)
         );
  OAI221XL U399 ( .A0(n167), .A1(n247), .B0(n246), .B1(n163), .C0(n168), .Y(
        n514) );
  AOI22X1 U400 ( .A0(din[85]), .A1(n176), .B0(dout[149]), .B1(n154), .Y(n168)
         );
  OAI221XL U401 ( .A0(n166), .A1(n243), .B0(n241), .B1(n163), .C0(n171), .Y(
        n515) );
  AOI22X1 U402 ( .A0(din[86]), .A1(n176), .B0(dout[150]), .B1(n152), .Y(n171)
         );
  OAI221XL U403 ( .A0(n167), .A1(n238), .B0(n237), .B1(n161), .C0(n174), .Y(
        n516) );
  AOI22X1 U404 ( .A0(din[87]), .A1(n176), .B0(dout[151]), .B1(n151), .Y(n174)
         );
  OAI221XL U405 ( .A0(n167), .A1(n234), .B0(n232), .B1(n164), .C0(n177), .Y(
        n517) );
  AOI22X1 U406 ( .A0(din[88]), .A1(n176), .B0(dout[152]), .B1(n152), .Y(n177)
         );
  OAI221XL U407 ( .A0(n167), .A1(n229), .B0(n227), .B1(n163), .C0(n180), .Y(
        n518) );
  AOI22X1 U408 ( .A0(din[89]), .A1(n176), .B0(dout[153]), .B1(n150), .Y(n180)
         );
  OAI221XL U409 ( .A0(n166), .A1(n223), .B0(n221), .B1(n161), .C0(n183), .Y(
        n519) );
  AOI22X1 U410 ( .A0(din[90]), .A1(n176), .B0(dout[154]), .B1(n151), .Y(n183)
         );
  OAI221XL U411 ( .A0(n166), .A1(n217), .B0(n215), .B1(n164), .C0(n186), .Y(
        n520) );
  AOI22X1 U412 ( .A0(din[91]), .A1(n176), .B0(dout[155]), .B1(n150), .Y(n186)
         );
  OAI221XL U413 ( .A0(n166), .A1(n211), .B0(n209), .B1(n163), .C0(n189), .Y(
        n521) );
  AOI22X1 U414 ( .A0(din[92]), .A1(n176), .B0(dout[156]), .B1(n150), .Y(n189)
         );
  OAI221XL U415 ( .A0(n167), .A1(n205), .B0(n203), .B1(n161), .C0(n192), .Y(
        n522) );
  AOI22X1 U416 ( .A0(din[93]), .A1(n178), .B0(dout[157]), .B1(n150), .Y(n192)
         );
  OAI221XL U417 ( .A0(n166), .A1(n199), .B0(n197), .B1(n161), .C0(n195), .Y(
        n523) );
  AOI22X1 U418 ( .A0(din[94]), .A1(n181), .B0(dout[158]), .B1(n150), .Y(n195)
         );
  OAI221XL U419 ( .A0(n167), .A1(n194), .B0(n193), .B1(n164), .C0(n198), .Y(
        n524) );
  AOI22X1 U420 ( .A0(din[95]), .A1(n176), .B0(dout[159]), .B1(n150), .Y(n198)
         );
  OAI221XL U421 ( .A0(n268), .A1(n166), .B0(n649), .B1(n163), .C0(n200), .Y(
        n525) );
  AOI22X1 U422 ( .A0(din[144]), .A1(n181), .B0(dout[160]), .B1(n150), .Y(n200)
         );
  OAI221XL U423 ( .A0(n264), .A1(n169), .B0(n646), .B1(n164), .C0(n202), .Y(
        n526) );
  AOI22X1 U424 ( .A0(din[145]), .A1(n181), .B0(dout[161]), .B1(n150), .Y(n202)
         );
  OAI221XL U425 ( .A0(n259), .A1(n169), .B0(n643), .B1(n163), .C0(n204), .Y(
        n527) );
  AOI22X1 U426 ( .A0(din[146]), .A1(n178), .B0(dout[162]), .B1(n150), .Y(n204)
         );
  OAI221XL U427 ( .A0(n255), .A1(n167), .B0(n640), .B1(n161), .C0(n206), .Y(
        n528) );
  AOI22X1 U428 ( .A0(din[147]), .A1(n179), .B0(dout[163]), .B1(n150), .Y(n206)
         );
  OAI221XL U429 ( .A0(n250), .A1(n169), .B0(n637), .B1(n164), .C0(n208), .Y(
        n529) );
  AOI22X1 U430 ( .A0(din[148]), .A1(n181), .B0(dout[164]), .B1(n150), .Y(n208)
         );
  OAI221XL U431 ( .A0(n246), .A1(n169), .B0(n634), .B1(n163), .C0(n210), .Y(
        n530) );
  AOI22X1 U432 ( .A0(din[149]), .A1(n176), .B0(dout[165]), .B1(n150), .Y(n210)
         );
  OAI221XL U433 ( .A0(n241), .A1(n166), .B0(n631), .B1(n161), .C0(n212), .Y(
        n531) );
  AOI22X1 U434 ( .A0(din[150]), .A1(n181), .B0(dout[166]), .B1(n150), .Y(n212)
         );
  OAI221XL U435 ( .A0(n237), .A1(n167), .B0(n628), .B1(n164), .C0(n214), .Y(
        n532) );
  AOI22X1 U436 ( .A0(din[151]), .A1(n179), .B0(dout[167]), .B1(n152), .Y(n214)
         );
  OAI221XL U437 ( .A0(n232), .A1(n169), .B0(n625), .B1(n161), .C0(n216), .Y(
        n533) );
  AOI22X1 U438 ( .A0(din[152]), .A1(n178), .B0(dout[168]), .B1(n152), .Y(n216)
         );
  OAI221XL U439 ( .A0(n227), .A1(n167), .B0(n325), .B1(n163), .C0(n218), .Y(
        n534) );
  AOI22X1 U440 ( .A0(din[153]), .A1(n179), .B0(dout[169]), .B1(n150), .Y(n218)
         );
  OAI221XL U441 ( .A0(n221), .A1(n169), .B0(n319), .B1(n161), .C0(n220), .Y(
        n535) );
  AOI22X1 U442 ( .A0(din[154]), .A1(n179), .B0(dout[170]), .B1(n150), .Y(n220)
         );
  OAI221XL U443 ( .A0(n215), .A1(n167), .B0(n313), .B1(n164), .C0(n222), .Y(
        n536) );
  AOI22X1 U444 ( .A0(din[155]), .A1(n181), .B0(dout[171]), .B1(n151), .Y(n222)
         );
  OAI221XL U445 ( .A0(n209), .A1(n167), .B0(n307), .B1(n164), .C0(n224), .Y(
        n537) );
  AOI22X1 U446 ( .A0(din[156]), .A1(n176), .B0(dout[172]), .B1(n160), .Y(n224)
         );
  OAI221XL U447 ( .A0(n203), .A1(n167), .B0(n301), .B1(n161), .C0(n226), .Y(
        n538) );
  AOI22X1 U448 ( .A0(din[157]), .A1(n178), .B0(dout[173]), .B1(n160), .Y(n226)
         );
  OAI221XL U449 ( .A0(n197), .A1(n166), .B0(n295), .B1(n163), .C0(n228), .Y(
        n539) );
  AOI22X1 U450 ( .A0(din[158]), .A1(n178), .B0(dout[174]), .B1(n152), .Y(n228)
         );
  OAI221XL U451 ( .A0(n193), .A1(n167), .B0(n274), .B1(n161), .C0(n230), .Y(
        n540) );
  AOI22X1 U452 ( .A0(din[159]), .A1(n176), .B0(dout[175]), .B1(n160), .Y(n230)
         );
  OAI221XL U453 ( .A0(n166), .A1(n267), .B0(n647), .B1(n164), .C0(n233), .Y(
        n541) );
  AOI22X1 U454 ( .A0(din[208]), .A1(n179), .B0(dout[176]), .B1(n154), .Y(n233)
         );
  OAI221XL U455 ( .A0(n166), .A1(n262), .B0(n644), .B1(n163), .C0(n236), .Y(
        n542) );
  AOI22X1 U456 ( .A0(din[209]), .A1(n176), .B0(dout[177]), .B1(n160), .Y(n236)
         );
  OAI221XL U457 ( .A0(n166), .A1(n258), .B0(n641), .B1(n161), .C0(n239), .Y(
        n543) );
  AOI22X1 U458 ( .A0(din[210]), .A1(n179), .B0(dout[178]), .B1(n151), .Y(n239)
         );
  OAI221XL U459 ( .A0(n166), .A1(n253), .B0(n638), .B1(n164), .C0(n242), .Y(
        n544) );
  AOI22X1 U460 ( .A0(din[211]), .A1(n176), .B0(dout[179]), .B1(n152), .Y(n242)
         );
  OAI221XL U461 ( .A0(n166), .A1(n249), .B0(n635), .B1(n161), .C0(n245), .Y(
        n545) );
  AOI22X1 U462 ( .A0(din[212]), .A1(n178), .B0(dout[180]), .B1(n151), .Y(n245)
         );
  OAI221XL U463 ( .A0(n166), .A1(n244), .B0(n632), .B1(n164), .C0(n248), .Y(
        n546) );
  AOI22X1 U464 ( .A0(din[213]), .A1(n181), .B0(dout[181]), .B1(n160), .Y(n248)
         );
  OAI221XL U465 ( .A0(n166), .A1(n240), .B0(n629), .B1(n163), .C0(n251), .Y(
        n547) );
  AOI22X1 U466 ( .A0(din[214]), .A1(n176), .B0(dout[182]), .B1(n152), .Y(n251)
         );
  OAI221XL U467 ( .A0(n166), .A1(n235), .B0(n626), .B1(n164), .C0(n254), .Y(
        n548) );
  AOI22X1 U468 ( .A0(din[215]), .A1(n178), .B0(dout[183]), .B1(n160), .Y(n254)
         );
  OAI221XL U469 ( .A0(n166), .A1(n231), .B0(n623), .B1(n163), .C0(n257), .Y(
        n549) );
  AOI22X1 U470 ( .A0(din[216]), .A1(n181), .B0(dout[184]), .B1(n150), .Y(n257)
         );
  OAI221XL U471 ( .A0(n167), .A1(n225), .B0(n321), .B1(n164), .C0(n260), .Y(
        n550) );
  AOI22X1 U472 ( .A0(din[217]), .A1(n181), .B0(dout[185]), .B1(n190), .Y(n260)
         );
  OAI221XL U473 ( .A0(n166), .A1(n219), .B0(n315), .B1(n163), .C0(n263), .Y(
        n551) );
  AOI22X1 U474 ( .A0(din[218]), .A1(n179), .B0(dout[186]), .B1(n160), .Y(n263)
         );
  OAI221XL U475 ( .A0(n169), .A1(n213), .B0(n309), .B1(n163), .C0(n266), .Y(
        n552) );
  AOI22X1 U476 ( .A0(din[219]), .A1(n179), .B0(dout[187]), .B1(n150), .Y(n266)
         );
  OAI221XL U477 ( .A0(n166), .A1(n207), .B0(n303), .B1(n163), .C0(n269), .Y(
        n553) );
  AOI22X1 U478 ( .A0(din[220]), .A1(n176), .B0(dout[188]), .B1(n151), .Y(n269)
         );
  OAI221XL U479 ( .A0(n167), .A1(n201), .B0(n297), .B1(n161), .C0(n272), .Y(
        n554) );
  AOI22X1 U480 ( .A0(din[221]), .A1(n178), .B0(dout[189]), .B1(n152), .Y(n272)
         );
  OAI221XL U481 ( .A0(n169), .A1(n196), .B0(n276), .B1(n164), .C0(n275), .Y(
        n555) );
  AOI22X1 U482 ( .A0(din[222]), .A1(n176), .B0(dout[190]), .B1(n160), .Y(n275)
         );
  OAI221XL U483 ( .A0(n166), .A1(n191), .B0(n271), .B1(n163), .C0(n278), .Y(
        n556) );
  AOI22X1 U484 ( .A0(din[223]), .A1(n178), .B0(dout[191]), .B1(n160), .Y(n278)
         );
  OAI221XL U485 ( .A0(n649), .A1(n166), .B0(n270), .B1(n161), .C0(n279), .Y(
        n557) );
  AOI22X1 U486 ( .A0(din[48]), .A1(n176), .B0(dout[192]), .B1(n152), .Y(n279)
         );
  INVX1 U487 ( .A(start), .Y(n190) );
  INVX1 U488 ( .A(mode[1]), .Y(n364) );
  NOR2X1 U489 ( .A(n364), .B(mode[0]), .Y(n343) );
  INVX1 U490 ( .A(n1), .Y(n365) );
  AOI22X1 U491 ( .A0(din[0]), .A1(n187), .B0(dout[0]), .B1(n150), .Y(n1) );
  INVX1 U492 ( .A(n3), .Y(n366) );
  AOI22X1 U493 ( .A0(din[1]), .A1(n187), .B0(dout[1]), .B1(n150), .Y(n3) );
  INVX1 U494 ( .A(n4), .Y(n367) );
  AOI22X1 U495 ( .A0(din[2]), .A1(n187), .B0(dout[2]), .B1(n154), .Y(n4) );
  INVX1 U496 ( .A(n5), .Y(n368) );
  AOI22X1 U497 ( .A0(din[3]), .A1(n187), .B0(dout[3]), .B1(n154), .Y(n5) );
  INVX1 U498 ( .A(n6), .Y(n369) );
  AOI22X1 U499 ( .A0(din[4]), .A1(n187), .B0(dout[4]), .B1(n154), .Y(n6) );
  INVX1 U500 ( .A(n7), .Y(n370) );
  AOI22X1 U501 ( .A0(din[5]), .A1(n187), .B0(dout[5]), .B1(n154), .Y(n7) );
  INVX1 U502 ( .A(n8), .Y(n371) );
  AOI22X1 U503 ( .A0(din[6]), .A1(n187), .B0(dout[6]), .B1(n154), .Y(n8) );
  INVX1 U504 ( .A(n9), .Y(n372) );
  AOI22X1 U505 ( .A0(din[7]), .A1(n187), .B0(dout[7]), .B1(n154), .Y(n9) );
  INVX1 U506 ( .A(n10), .Y(n373) );
  AOI22X1 U507 ( .A0(din[8]), .A1(n187), .B0(dout[8]), .B1(n154), .Y(n10) );
  INVX1 U508 ( .A(n11), .Y(n374) );
  AOI22X1 U509 ( .A0(din[9]), .A1(n187), .B0(dout[9]), .B1(n150), .Y(n11) );
  INVX1 U510 ( .A(n12), .Y(n375) );
  AOI22X1 U511 ( .A0(din[10]), .A1(n187), .B0(dout[10]), .B1(n154), .Y(n12) );
  INVX1 U512 ( .A(n13), .Y(n376) );
  AOI22X1 U513 ( .A0(din[11]), .A1(n187), .B0(dout[11]), .B1(n160), .Y(n13) );
  INVX1 U514 ( .A(n14), .Y(n377) );
  AOI22X1 U515 ( .A0(din[12]), .A1(n187), .B0(dout[12]), .B1(n151), .Y(n14) );
  INVX1 U516 ( .A(n15), .Y(n378) );
  AOI22X1 U517 ( .A0(din[13]), .A1(N275), .B0(dout[13]), .B1(n150), .Y(n15) );
  INVX1 U518 ( .A(n16), .Y(n379) );
  AOI22X1 U519 ( .A0(din[14]), .A1(N275), .B0(dout[14]), .B1(n152), .Y(n16) );
  INVX1 U520 ( .A(n17), .Y(n380) );
  AOI22X1 U521 ( .A0(din[15]), .A1(N275), .B0(dout[15]), .B1(n152), .Y(n17) );
  INVX1 U522 ( .A(n346), .Y(n605) );
  AOI22X1 U523 ( .A0(din[240]), .A1(N275), .B0(dout[240]), .B1(n151), .Y(n346)
         );
  INVX1 U524 ( .A(n347), .Y(n606) );
  AOI22X1 U525 ( .A0(din[241]), .A1(N275), .B0(dout[241]), .B1(n151), .Y(n347)
         );
  INVX1 U526 ( .A(n348), .Y(n607) );
  AOI22X1 U527 ( .A0(din[242]), .A1(N275), .B0(dout[242]), .B1(n152), .Y(n348)
         );
  INVX1 U528 ( .A(n349), .Y(n608) );
  AOI22X1 U529 ( .A0(din[243]), .A1(N275), .B0(dout[243]), .B1(n190), .Y(n349)
         );
  INVX1 U530 ( .A(n350), .Y(n609) );
  AOI22X1 U531 ( .A0(din[244]), .A1(N275), .B0(dout[244]), .B1(n151), .Y(n350)
         );
  INVX1 U532 ( .A(n351), .Y(n610) );
  AOI22X1 U533 ( .A0(din[245]), .A1(N275), .B0(dout[245]), .B1(n190), .Y(n351)
         );
  INVX1 U534 ( .A(n352), .Y(n611) );
  AOI22X1 U535 ( .A0(din[246]), .A1(N275), .B0(dout[246]), .B1(n150), .Y(n352)
         );
  INVX1 U536 ( .A(n353), .Y(n612) );
  AOI22X1 U537 ( .A0(din[247]), .A1(N275), .B0(dout[247]), .B1(n152), .Y(n353)
         );
  INVX1 U538 ( .A(n354), .Y(n613) );
  AOI22X1 U539 ( .A0(din[248]), .A1(N275), .B0(dout[248]), .B1(n151), .Y(n354)
         );
  INVX1 U540 ( .A(n355), .Y(n614) );
  AOI22X1 U541 ( .A0(din[249]), .A1(N275), .B0(dout[249]), .B1(n152), .Y(n355)
         );
  INVX1 U542 ( .A(n356), .Y(n615) );
  AOI22X1 U543 ( .A0(din[250]), .A1(n187), .B0(dout[250]), .B1(n190), .Y(n356)
         );
  INVX1 U544 ( .A(n357), .Y(n616) );
  AOI22X1 U545 ( .A0(din[251]), .A1(n187), .B0(dout[251]), .B1(n150), .Y(n357)
         );
  INVX1 U546 ( .A(n358), .Y(n617) );
  AOI22X1 U547 ( .A0(din[252]), .A1(N275), .B0(dout[252]), .B1(n160), .Y(n358)
         );
  INVX1 U548 ( .A(n359), .Y(n618) );
  AOI22X1 U549 ( .A0(din[253]), .A1(N275), .B0(dout[253]), .B1(n160), .Y(n359)
         );
  INVX1 U550 ( .A(n360), .Y(n619) );
  AOI22X1 U551 ( .A0(din[254]), .A1(N275), .B0(dout[254]), .B1(n190), .Y(n360)
         );
  INVX1 U552 ( .A(n361), .Y(n620) );
  AOI22X1 U553 ( .A0(din[255]), .A1(N275), .B0(dout[255]), .B1(n151), .Y(n361)
         );
  OAI21XL U554 ( .A0(n362), .A1(n364), .B0(start), .Y(n363) );
  OAI2BB2X1 U555 ( .B0(n362), .B1(n363), .A0N(mode_out[0]), .A1N(n363), .Y(
        n621) );
  OAI2BB2X1 U556 ( .B0(n364), .B1(n363), .A0N(mode_out[1]), .A1N(n363), .Y(
        n622) );
  INVX1 U557 ( .A(din[144]), .Y(n270) );
  INVX1 U558 ( .A(din[145]), .Y(n265) );
  INVX1 U559 ( .A(din[146]), .Y(n261) );
  INVX1 U560 ( .A(din[147]), .Y(n256) );
  INVX1 U561 ( .A(din[148]), .Y(n252) );
  INVX1 U562 ( .A(din[149]), .Y(n247) );
  INVX1 U563 ( .A(din[150]), .Y(n243) );
  INVX1 U564 ( .A(din[151]), .Y(n238) );
  INVX1 U565 ( .A(din[152]), .Y(n234) );
  INVX1 U566 ( .A(din[153]), .Y(n229) );
  INVX1 U567 ( .A(din[154]), .Y(n223) );
  INVX1 U568 ( .A(din[155]), .Y(n217) );
  INVX1 U569 ( .A(din[156]), .Y(n211) );
  INVX1 U570 ( .A(din[157]), .Y(n205) );
  INVX1 U571 ( .A(din[158]), .Y(n199) );
  INVX1 U572 ( .A(din[159]), .Y(n194) );
  INVX1 U573 ( .A(din[176]), .Y(n267) );
  INVX1 U574 ( .A(din[177]), .Y(n262) );
  INVX1 U575 ( .A(din[178]), .Y(n258) );
  INVX1 U576 ( .A(din[179]), .Y(n253) );
  INVX1 U577 ( .A(din[180]), .Y(n249) );
  INVX1 U578 ( .A(din[181]), .Y(n244) );
  INVX1 U579 ( .A(din[182]), .Y(n240) );
  INVX1 U580 ( .A(din[183]), .Y(n235) );
  INVX1 U581 ( .A(din[184]), .Y(n231) );
  INVX1 U582 ( .A(din[185]), .Y(n225) );
  INVX1 U583 ( .A(din[186]), .Y(n219) );
  INVX1 U584 ( .A(din[187]), .Y(n213) );
  INVX1 U585 ( .A(din[188]), .Y(n207) );
  INVX1 U586 ( .A(din[189]), .Y(n201) );
  INVX1 U587 ( .A(din[190]), .Y(n196) );
  INVX1 U588 ( .A(din[191]), .Y(n191) );
  INVX1 U589 ( .A(din[208]), .Y(n648) );
  INVX1 U590 ( .A(din[209]), .Y(n645) );
  INVX1 U591 ( .A(din[210]), .Y(n642) );
  INVX1 U592 ( .A(din[211]), .Y(n639) );
  INVX1 U593 ( .A(din[212]), .Y(n636) );
  INVX1 U594 ( .A(din[213]), .Y(n633) );
  INVX1 U595 ( .A(din[214]), .Y(n630) );
  INVX1 U596 ( .A(din[215]), .Y(n627) );
  INVX1 U597 ( .A(din[216]), .Y(n624) );
  INVX1 U598 ( .A(din[217]), .Y(n323) );
  INVX1 U599 ( .A(din[218]), .Y(n317) );
  INVX1 U600 ( .A(din[219]), .Y(n311) );
  INVX1 U601 ( .A(din[220]), .Y(n305) );
  INVX1 U602 ( .A(din[221]), .Y(n299) );
  INVX1 U603 ( .A(din[222]), .Y(n277) );
  INVX1 U604 ( .A(din[223]), .Y(n273) );
  INVX1 U605 ( .A(din[160]), .Y(n268) );
  INVX1 U606 ( .A(din[161]), .Y(n264) );
  INVX1 U607 ( .A(din[162]), .Y(n259) );
  INVX1 U608 ( .A(din[163]), .Y(n255) );
  INVX1 U609 ( .A(din[164]), .Y(n250) );
  INVX1 U610 ( .A(din[165]), .Y(n246) );
  INVX1 U611 ( .A(din[166]), .Y(n241) );
  INVX1 U612 ( .A(din[167]), .Y(n237) );
  INVX1 U613 ( .A(din[168]), .Y(n232) );
  INVX1 U614 ( .A(din[169]), .Y(n227) );
  INVX1 U615 ( .A(din[170]), .Y(n221) );
  INVX1 U616 ( .A(din[171]), .Y(n215) );
  INVX1 U617 ( .A(din[172]), .Y(n209) );
  INVX1 U618 ( .A(din[173]), .Y(n203) );
  INVX1 U619 ( .A(din[174]), .Y(n197) );
  INVX1 U620 ( .A(din[175]), .Y(n193) );
  INVX1 U621 ( .A(din[192]), .Y(n649) );
  INVX1 U622 ( .A(din[193]), .Y(n646) );
  INVX1 U623 ( .A(din[194]), .Y(n643) );
  INVX1 U624 ( .A(din[195]), .Y(n640) );
  INVX1 U625 ( .A(din[196]), .Y(n637) );
  INVX1 U626 ( .A(din[197]), .Y(n634) );
  INVX1 U627 ( .A(din[198]), .Y(n631) );
  INVX1 U628 ( .A(din[199]), .Y(n628) );
  INVX1 U629 ( .A(din[200]), .Y(n625) );
  INVX1 U630 ( .A(din[201]), .Y(n325) );
  INVX1 U631 ( .A(din[202]), .Y(n319) );
  INVX1 U632 ( .A(din[203]), .Y(n313) );
  INVX1 U633 ( .A(din[204]), .Y(n307) );
  INVX1 U634 ( .A(din[205]), .Y(n301) );
  INVX1 U635 ( .A(din[206]), .Y(n295) );
  INVX1 U636 ( .A(din[207]), .Y(n274) );
  INVX1 U637 ( .A(din[224]), .Y(n647) );
  INVX1 U638 ( .A(din[225]), .Y(n644) );
  INVX1 U639 ( .A(din[226]), .Y(n641) );
  INVX1 U640 ( .A(din[227]), .Y(n638) );
  INVX1 U641 ( .A(din[228]), .Y(n635) );
  INVX1 U642 ( .A(din[229]), .Y(n632) );
  INVX1 U643 ( .A(din[230]), .Y(n629) );
  INVX1 U644 ( .A(din[231]), .Y(n626) );
  INVX1 U645 ( .A(din[232]), .Y(n623) );
  INVX1 U646 ( .A(din[233]), .Y(n321) );
  INVX1 U647 ( .A(din[234]), .Y(n315) );
  INVX1 U648 ( .A(din[235]), .Y(n309) );
  INVX1 U649 ( .A(din[236]), .Y(n303) );
  INVX1 U650 ( .A(din[237]), .Y(n297) );
  INVX1 U651 ( .A(din[238]), .Y(n276) );
  INVX1 U652 ( .A(din[239]), .Y(n271) );
endmodule


module idct4_shift7_add64_DW01_add_4 ( A, B, SUM );
  input [24:0] A;
  input [24:0] B;
  output [24:0] SUM;
  wire   n2;
  wire   [24:1] carry;

  XOR3X2 U1_24 ( .A(A[24]), .B(B[24]), .C(carry[24]), .Y(SUM[24]) );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_5 ( .A(1'b0), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(1'b0), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(1'b0), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(1'b0), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_1 ( .A(1'b0), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  CLKINVX8 U1 ( .A(n2), .Y(carry[1]) );
  CLKINVX8 U2 ( .A(B[0]), .Y(SUM[0]) );
  INVX1 U4 ( .A(B[0]), .Y(n2) );
endmodule


module idct4_shift7_add64_DW01_add_5 ( A, B, SUM );
  input [24:0] A;
  input [24:0] B;
  output [24:0] SUM;
  wire   n2;
  wire   [24:1] carry;

  XOR3X2 U1_24 ( .A(A[24]), .B(B[24]), .C(carry[24]), .Y(SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(1'b0), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(1'b0), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(1'b0), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(1'b0), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_1 ( .A(1'b0), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  CLKINVX8 U1 ( .A(n2), .Y(carry[1]) );
  CLKINVX8 U2 ( .A(B[0]), .Y(SUM[0]) );
  INVX1 U4 ( .A(B[0]), .Y(n2) );
endmodule


module idct4_shift7_add64_DW01_add_6 ( A, B, SUM );
  input [24:0] A;
  input [24:0] B;
  output [24:0] SUM;

  wire   [24:1] carry;

  XOR3X2 U1_24 ( .A(A[24]), .B(B[24]), .C(carry[24]), .Y(SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_1 ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(SUM[1]) );
  ADDFX2 U1_5 ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(SUM[5]) );
  ADDFX2 U1_4 ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(SUM[4]) );
  ADDFX2 U1_3 ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(SUM[3]) );
  ADDFX2 U1_2 ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(SUM[2]) );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(1'b0), .CO(carry[7]), .S(SUM[6]) );
  XOR2X1 U1 ( .A(B[0]), .B(1'b0), .Y(SUM[0]) );
endmodule


module idct4_shift7_add64_DW01_add_7 ( A, B, SUM );
  input [24:0] A;
  input [24:0] B;
  output [24:0] SUM;

  wire   [24:1] carry;

  XOR3X2 U1_24 ( .A(A[24]), .B(B[24]), .C(carry[24]), .Y(SUM[24]) );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_1 ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(SUM[1]) );
  ADDFX2 U1_5 ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(SUM[5]) );
  ADDFX2 U1_4 ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(SUM[4]) );
  ADDFX2 U1_3 ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(SUM[3]) );
  ADDFX2 U1_2 ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(SUM[2]) );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(1'b0), .CO(carry[7]), .S(SUM[6]) );
  XOR2X1 U1 ( .A(B[0]), .B(1'b0), .Y(SUM[0]) );
endmodule


module idct4_shift7_add64_DW01_add_8 ( A, B, SUM );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;

  wire   [23:1] carry;

  XOR3X2 U1_23 ( .A(A[23]), .B(B[23]), .C(carry[23]), .Y(SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_1 ( .A(A[1]), .B(1'b0), .CI(1'b0), .S(SUM[1]) );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(1'b0), .CO(carry[3]), .S(SUM[2]) );
  XOR2X1 U1 ( .A(1'b0), .B(A[0]), .Y(SUM[0]) );
endmodule


module idct4_shift7_add64_DW01_add_9 ( A, B, SUM );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  wire   n2;
  wire   [23:1] carry;

  XOR3X2 U1_23 ( .A(A[23]), .B(B[23]), .C(carry[23]), .Y(SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_1 ( .A(1'b0), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  CLKINVX8 U1 ( .A(n2), .Y(carry[1]) );
  CLKINVX8 U2 ( .A(B[0]), .Y(SUM[0]) );
  INVX1 U4 ( .A(B[0]), .Y(n2) );
endmodule


module idct4_shift7_add64_DW01_add_12 ( A, B, SUM );
  input [22:0] A;
  input [22:0] B;
  output [22:0] SUM;

  wire   [22:1] carry;

  XOR3X2 U1_22 ( .A(A[22]), .B(B[22]), .C(carry[22]), .Y(SUM[22]) );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(1'b0), .CO(carry[2]), .S(SUM[1]) );
  XOR2X1 U1 ( .A(1'b0), .B(A[0]), .Y(SUM[0]) );
endmodule


module idct4_shift7_add64_DW01_add_13 ( A, B, SUM );
  input [22:0] A;
  input [22:0] B;
  output [22:0] SUM;

  wire   [22:1] carry;

  XOR3X2 U1_22 ( .A(A[22]), .B(B[22]), .C(carry[22]), .Y(SUM[22]) );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(1'b0), .CO(carry[2]), .S(SUM[1]) );
  XOR2X1 U1 ( .A(1'b0), .B(A[0]), .Y(SUM[0]) );
endmodule


module idct4_shift7_add64 ( clk, rstn, mode, start, x0, x1, x2, x3, y0, y1, y2, 
        y3, idct4_ready );
  input [1:0] mode;
  input [15:0] x0;
  input [15:0] x1;
  input [15:0] x2;
  input [15:0] x3;
  output [24:0] y0;
  output [24:0] y1;
  output [24:0] y2;
  output [24:0] y3;
  input clk, rstn, start;
  output idct4_ready;
  wire   idct4_ready_delay1, idct4_ready_delay2, idct4_ready_delay3, N14, N15,
         N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29,
         N30, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48,
         N49, N50, N51, N52, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68,
         N69, N70, N71, N72, N73, N74, N80, N81, N82, N83, N84, N85, N86, N87,
         N88, N89, N90, N91, N92, N93, N94, N95, N103, N104, N105, N106, N107,
         N108, N109, N110, N111, N112, N113, N114, N115, N116, N117, N118,
         N124, N125, N126, N127, N128, N129, N130, N131, N132, N133, N134,
         N135, N136, N137, N138, N139, N141, N142, N143, N144, N145, N146,
         N147, N148, N149, N150, N151, N152, N153, N154, N155, N156, N157,
         N158, N159, N160, N161, N162, N163, N164, N165, N166, N167, N168,
         N169, N170, N171, N172, N173, N174, N175, N176, N177, N178, N179,
         N180, N181, N182, N183, N184, N185, N186, N193, N194, N195, N196,
         N197, N198, N199, N200, N201, N202, N203, N204, N205, N206, N207,
         N208, N209, N261, N262, N263, N264, N265, N266, N267, N268, N269,
         N270, N271, N272, N273, N274, N275, N276, N277, N325, N326, N327,
         N328, N329, N330, N331, N332, N333, N334, N335, N336, N337, N338,
         N339, N340, N341, N342, N343, N344, N345, N346, N347, N348, N349,
         N350, N351, N352, N353, N354, N355, N356, N357, N358, N359, N360,
         N361, N362, N363, N364, N365, N366, N367, N368, N369, N370, N371,
         N372, N373, N374, N375, N376, N377, N378, N379, N380, N381, N382,
         N383, N384, N385, N386, N387, N388, N389, N390, N391, N392, N393,
         N394, N395, N396, N397, N398, N399, N400, N401, N402, N403, N404,
         N405, N406, N407, N408, N409, N410, N411, N412, N413, N414, N415,
         N416, N417, N418, N419, N420, N421, N422, N472, N473, N474, N475,
         N476, N477, N478, N479, N480, N481, N482, N483, N484, N485, N486,
         N487, N488, N489, N490, N491, N492, N493, N494, N495, N496, N546,
         N547, N548, N549, N550, N551, N552, N553, N554, N555, N556, N557,
         N558, N559, N560, N561, N562, N563, N564, N565, N566, N567, N568,
         N569, N570, N571, N572, N573, N574, N575, N576, N577, N578, N579,
         N580, N581, N582, N583, N584, N585, N586, N587, N588, N589, N590,
         N591, N592, N593, N594, N595, N596, N597, N598, N599, N600, N601,
         N602, N603, N604, N605, N606, N607, N608, N609, N610, N611, N612,
         N613, N614, N615, N616, N617, N618, N619, N620, N621, N622, N623,
         N624, N625, N626, N627, N628, N629, N630, N631, N632, N633, N634,
         N635, N636, N637, N638, N639, N640, N641, N642, N643, N644, N645,
         N646, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, add_125_carry_8_, add_125_carry_9_, add_125_carry_10_,
         add_125_carry_11_, add_125_carry_12_, add_125_carry_13_,
         add_125_carry_14_, add_125_carry_15_, add_125_carry_16_,
         add_125_carry_17_, add_125_carry_18_, add_125_carry_19_,
         add_125_carry_20_, add_125_carry_21_, add_125_carry_22_,
         add_125_carry_23_, add_125_carry_24_, add_125_carry_25_,
         add_124_carry_8_, add_124_carry_9_, add_124_carry_10_,
         add_124_carry_11_, add_124_carry_12_, add_124_carry_13_,
         add_124_carry_14_, add_124_carry_15_, add_124_carry_16_,
         add_124_carry_17_, add_124_carry_18_, add_124_carry_19_,
         add_124_carry_20_, add_124_carry_21_, add_124_carry_22_,
         add_124_carry_23_, add_124_carry_24_, add_124_carry_25_,
         add_123_carry_8_, add_123_carry_9_, add_123_carry_10_,
         add_123_carry_11_, add_123_carry_12_, add_123_carry_13_,
         add_123_carry_14_, add_123_carry_15_, add_123_carry_16_,
         add_123_carry_17_, add_123_carry_18_, add_123_carry_19_,
         add_123_carry_20_, add_123_carry_21_, add_123_carry_22_,
         add_123_carry_23_, add_123_carry_24_, add_123_carry_25_,
         add_122_carry_8_, add_122_carry_9_, add_122_carry_10_,
         add_122_carry_11_, add_122_carry_12_, add_122_carry_13_,
         add_122_carry_14_, add_122_carry_15_, add_122_carry_16_,
         add_122_carry_17_, add_122_carry_18_, add_122_carry_19_,
         add_122_carry_20_, add_122_carry_21_, add_122_carry_22_,
         add_122_carry_23_, add_122_carry_24_, add_122_carry_25_,
         add_1_root_add_112_2_B_6_, add_1_root_add_112_2_B_7_,
         add_1_root_add_112_2_B_8_, add_1_root_add_112_2_B_9_,
         add_1_root_add_112_2_B_10_, add_1_root_add_112_2_B_11_,
         add_1_root_add_112_2_B_12_, add_1_root_add_112_2_B_13_,
         add_1_root_add_112_2_B_14_, add_1_root_add_112_2_B_15_,
         add_1_root_add_112_2_B_16_, add_1_root_add_112_2_B_17_,
         add_1_root_add_112_2_B_18_, add_1_root_add_112_2_B_19_,
         add_1_root_add_112_2_B_20_, add_1_root_add_112_2_B_21_,
         add_88_carry_10_, add_88_carry_11_, add_88_carry_12_,
         add_88_carry_13_, add_88_carry_14_, add_88_carry_15_,
         add_88_carry_16_, add_88_carry_17_, add_88_carry_18_, add_88_carry_5_,
         add_88_carry_6_, add_88_carry_7_, add_88_carry_8_, add_88_carry_9_,
         add_87_carry_10_, add_87_carry_11_, add_87_carry_12_,
         add_87_carry_13_, add_87_carry_14_, add_87_carry_15_,
         add_87_carry_16_, add_87_carry_17_, add_87_carry_18_,
         add_87_carry_19_, add_87_carry_20_, add_87_carry_7_, add_87_carry_8_,
         add_87_carry_9_, add_86_carry_10_, add_86_carry_11_, add_86_carry_12_,
         add_86_carry_13_, add_86_carry_14_, add_86_carry_15_,
         add_86_carry_16_, add_86_carry_17_, add_86_carry_18_, add_86_carry_5_,
         add_86_carry_6_, add_86_carry_7_, add_86_carry_8_, add_86_carry_9_,
         add_85_carry_10_, add_85_carry_11_, add_85_carry_12_,
         add_85_carry_13_, add_85_carry_14_, add_85_carry_15_,
         add_85_carry_16_, add_85_carry_17_, add_85_carry_18_,
         add_85_carry_19_, add_85_carry_20_, add_85_carry_7_, add_85_carry_8_,
         add_85_carry_9_, add_81_carry_10_, add_81_carry_11_, add_81_carry_12_,
         add_81_carry_13_, add_81_carry_14_, add_81_carry_15_,
         add_81_carry_16_, add_81_carry_17_, add_81_carry_18_,
         add_81_carry_19_, add_81_carry_6_, add_81_carry_7_, add_81_carry_8_,
         add_81_carry_9_, add_80_carry_10_, add_80_carry_11_, add_80_carry_12_,
         add_80_carry_13_, add_80_carry_14_, add_80_carry_15_,
         add_80_carry_16_, add_80_carry_17_, add_80_carry_18_,
         add_80_carry_19_, add_80_carry_6_, add_80_carry_7_, add_80_carry_8_,
         add_80_carry_9_, n1, n2, n3, n4, n8, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120;
  wire   [1:0] mode_delay2;
  wire   [1:0] mode_delay1;
  wire   [20:0] x1_o0_tmp2;
  wire   [20:0] x3_o1_tmp2;
  wire   [21:6] x0_e;
  wire   [21:6] x2_e;
  wire   [21:0] x1_o1;
  wire   [21:0] x3_o0;
  wire   [22:0] x1_o0;
  wire   [22:0] x3_o1;
  wire   [21:2] x3_o0_tmp;
  wire   [21:2] x1_o1_tmp;
  wire   [21:6] x2_e_tmp;
  wire   [21:6] x0_e_tmp;
  wire   [22:0] x3_o1_tmp1;
  wire   [22:0] x1_o0_tmp1;
  wire   [22:0] e0;
  wire   [23:0] o0;
  wire   [22:0] e1;
  wire   [23:0] o1;
  wire   [24:0] y0_tmp;
  wire   [24:0] y1_tmp;
  wire   [24:0] y2_tmp;
  wire   [24:0] y3_tmp;
  wire   [22:7] add_1_root_add_112_2_carry;
  wire   [22:7] add_111_carry;

  idct4_shift7_add64_DW01_add_4 add_1_root_add_119_2 ( .A({e0[22], e0[22], 
        e0[22:6], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({n97, n97, n98, n99, 
        n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, 
        n112, n113, n114, n115, n116, n117, n118, n119, n120}), .SUM({N570, 
        N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, 
        N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546}) );
  idct4_shift7_add64_DW01_add_5 add_1_root_add_118_2 ( .A({e1[22], e1[22], 
        e1[22:6], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({n73, n73, n74, n75, 
        n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, 
        n90, n91, n92, n93, n94, n95, n96}), .SUM({N496, N495, N494, N493, 
        N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, 
        N480, N479, N478, N477, N476, N475, N474, N473, N472}) );
  idct4_shift7_add64_DW01_add_6 add_117 ( .A({e1[22], e1[22], e1[22:6], 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({o1[23], o1}), .SUM({N422, N421, 
        N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, 
        N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398}) );
  idct4_shift7_add64_DW01_add_7 add_116 ( .A({e0[22], e0[22], e0[22:6], 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({o0[23], o0}), .SUM({N397, N396, 
        N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, 
        N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373}) );
  idct4_shift7_add64_DW01_add_8 add_114 ( .A({x1_o0[22], x1_o0}), .B({
        x3_o0[21], x3_o0[21], x3_o0[21:2], 1'b0, 1'b0}), .SUM({N372, N371, 
        N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, 
        N358, N357, N356, N355, N354, N353, N352, N351, N350, N349}) );
  idct4_shift7_add64_DW01_add_9 add_1_root_add_113_2 ( .A({x1_o1[21], 
        x1_o1[21], x1_o1[21:2], 1'b0, 1'b0}), .B({n50, n50, n51, n52, n53, n54, 
        n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, 
        n69, n70, n71, n72}), .SUM({N348, N347, N346, N345, N344, N343, N342, 
        N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, 
        N329, N328, N327, N326, N325}) );
  idct4_shift7_add64_DW01_add_12 add_90 ( .A(x3_o1_tmp1), .B({x3_o1_tmp2[20], 
        x3_o1_tmp2[20], x3_o1_tmp2[20:1], 1'b0}), .SUM({N186, N185, N184, N183, 
        N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, 
        N170, N169, N168, N167, N166, N165, N164}) );
  idct4_shift7_add64_DW01_add_13 add_89 ( .A(x1_o0_tmp1), .B({x1_o0_tmp2[20], 
        x1_o0_tmp2[20], x1_o0_tmp2[20:1], 1'b0}), .SUM({N163, N162, N161, N160, 
        N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, 
        N147, N146, N145, N144, N143, N142, N141}) );
  DFFRHQX1 x3_o1_tmp1_reg_22_ ( .D(N52), .CK(clk), .RN(rstn), .Q(
        x3_o1_tmp1[22]) );
  DFFRHQX1 x3_o1_tmp1_reg_21_ ( .D(N118), .CK(clk), .RN(rstn), .Q(
        x3_o1_tmp1[21]) );
  DFFRHQX1 x3_o1_tmp1_reg_20_ ( .D(N117), .CK(clk), .RN(rstn), .Q(
        x3_o1_tmp1[20]) );
  DFFRHQX1 x3_o1_tmp1_reg_19_ ( .D(N116), .CK(clk), .RN(rstn), .Q(
        x3_o1_tmp1[19]) );
  DFFRHQX1 x1_o0_tmp1_reg_22_ ( .D(N30), .CK(clk), .RN(rstn), .Q(
        x1_o0_tmp1[22]) );
  DFFRHQX1 x1_o0_tmp1_reg_21_ ( .D(N74), .CK(clk), .RN(rstn), .Q(
        x1_o0_tmp1[21]) );
  DFFRHQX1 x1_o0_tmp1_reg_20_ ( .D(N73), .CK(clk), .RN(rstn), .Q(
        x1_o0_tmp1[20]) );
  DFFRHQX1 x1_o0_tmp1_reg_19_ ( .D(N72), .CK(clk), .RN(rstn), .Q(
        x1_o0_tmp1[19]) );
  DFFRHQX1 x1_o0_reg_20_ ( .D(N161), .CK(clk), .RN(rstn), .Q(x1_o0[20]) );
  DFFRHQX1 x1_o0_reg_21_ ( .D(N162), .CK(clk), .RN(rstn), .Q(x1_o0[21]) );
  DFFRHQX1 x1_o1_reg_20_ ( .D(x1_o1_tmp[20]), .CK(clk), .RN(rstn), .Q(
        x1_o1[20]) );
  DFFRHQX1 x3_o1_reg_22_ ( .D(N186), .CK(clk), .RN(rstn), .Q(x3_o1[22]) );
  DFFRHQX1 x3_o1_reg_21_ ( .D(N185), .CK(clk), .RN(rstn), .Q(x3_o1[21]) );
  DFFRHQX1 x3_o1_reg_20_ ( .D(N184), .CK(clk), .RN(rstn), .Q(x3_o1[20]) );
  DFFRHQX1 x1_o0_reg_22_ ( .D(N163), .CK(clk), .RN(rstn), .Q(x1_o0[22]) );
  DFFRHQX1 x0_e_reg_20_ ( .D(x0_e_tmp[20]), .CK(clk), .RN(rstn), .Q(x0_e[20])
         );
  DFFRHQX1 x0_e_reg_19_ ( .D(x0_e_tmp[19]), .CK(clk), .RN(rstn), .Q(x0_e[19])
         );
  DFFRHQX1 e1_reg_21_ ( .D(N276), .CK(clk), .RN(rstn), .Q(e1[21]) );
  DFFRHQX1 e0_reg_21_ ( .D(N208), .CK(clk), .RN(rstn), .Q(e0[21]) );
  DFFRHQX1 x3_o1_tmp2_reg_19_ ( .D(N139), .CK(clk), .RN(rstn), .Q(
        x3_o1_tmp2[19]) );
  DFFRHQX1 x1_o0_tmp2_reg_19_ ( .D(N95), .CK(clk), .RN(rstn), .Q(
        x1_o0_tmp2[19]) );
  DFFRHQX1 x3_o0_reg_20_ ( .D(x3_o0_tmp[20]), .CK(clk), .RN(rstn), .Q(
        x3_o0[20]) );
  DFFRHQX1 x3_o1_tmp1_reg_0_ ( .D(x3[0]), .CK(clk), .RN(rstn), .Q(
        x3_o1_tmp1[0]) );
  DFFRHQX1 x1_o0_tmp1_reg_0_ ( .D(x1[0]), .CK(clk), .RN(rstn), .Q(
        x1_o0_tmp1[0]) );
  DFFRHQX1 x1_o0_reg_0_ ( .D(N141), .CK(clk), .RN(rstn), .Q(x1_o0[0]) );
  DFFRHQX1 x1_o1_reg_21_ ( .D(x1_o1_tmp[21]), .CK(clk), .RN(rstn), .Q(
        x1_o1[21]) );
  DFFRHQX1 x0_e_reg_21_ ( .D(x0_e_tmp[21]), .CK(clk), .RN(rstn), .Q(x0_e[21])
         );
  DFFRHQX1 x2_e_reg_20_ ( .D(x2_e_tmp[20]), .CK(clk), .RN(rstn), .Q(x2_e[20])
         );
  DFFRHQX1 o1_reg_22_ ( .D(N347), .CK(clk), .RN(rstn), .Q(o1[22]) );
  DFFRHQX1 o0_reg_22_ ( .D(N371), .CK(clk), .RN(rstn), .Q(o0[22]) );
  DFFRHQX1 e1_reg_22_ ( .D(N277), .CK(clk), .RN(rstn), .Q(e1[22]) );
  DFFRHQX1 e0_reg_22_ ( .D(N209), .CK(clk), .RN(rstn), .Q(e0[22]) );
  DFFRHQX1 x2_e_reg_21_ ( .D(x2_e_tmp[21]), .CK(clk), .RN(rstn), .Q(x2_e[21])
         );
  DFFRHQX1 o1_reg_23_ ( .D(N348), .CK(clk), .RN(rstn), .Q(o1[23]) );
  DFFRHQX1 o0_reg_23_ ( .D(N372), .CK(clk), .RN(rstn), .Q(o0[23]) );
  DFFRHQX1 x3_o1_tmp2_reg_20_ ( .D(N52), .CK(clk), .RN(rstn), .Q(
        x3_o1_tmp2[20]) );
  DFFRHQX1 x1_o0_tmp2_reg_20_ ( .D(N30), .CK(clk), .RN(rstn), .Q(
        x1_o0_tmp2[20]) );
  DFFRHQX1 x3_o0_reg_21_ ( .D(x3_o0_tmp[21]), .CK(clk), .RN(rstn), .Q(
        x3_o0[21]) );
  DFFRHQX1 x3_o1_tmp1_reg_18_ ( .D(N115), .CK(clk), .RN(rstn), .Q(
        x3_o1_tmp1[18]) );
  DFFRHQX1 x3_o1_tmp1_reg_17_ ( .D(N114), .CK(clk), .RN(rstn), .Q(
        x3_o1_tmp1[17]) );
  DFFRHQX1 x3_o1_tmp1_reg_16_ ( .D(N113), .CK(clk), .RN(rstn), .Q(
        x3_o1_tmp1[16]) );
  DFFRHQX1 x3_o1_tmp1_reg_15_ ( .D(N112), .CK(clk), .RN(rstn), .Q(
        x3_o1_tmp1[15]) );
  DFFRHQX1 x1_o0_tmp1_reg_18_ ( .D(N71), .CK(clk), .RN(rstn), .Q(
        x1_o0_tmp1[18]) );
  DFFRHQX1 x1_o0_tmp1_reg_17_ ( .D(N70), .CK(clk), .RN(rstn), .Q(
        x1_o0_tmp1[17]) );
  DFFRHQX1 x1_o0_tmp1_reg_16_ ( .D(N69), .CK(clk), .RN(rstn), .Q(
        x1_o0_tmp1[16]) );
  DFFRHQX1 x1_o0_tmp1_reg_15_ ( .D(N68), .CK(clk), .RN(rstn), .Q(
        x1_o0_tmp1[15]) );
  DFFRHQX1 x1_o0_reg_16_ ( .D(N157), .CK(clk), .RN(rstn), .Q(x1_o0[16]) );
  DFFRHQX1 x1_o0_reg_17_ ( .D(N158), .CK(clk), .RN(rstn), .Q(x1_o0[17]) );
  DFFRHQX1 x1_o0_reg_18_ ( .D(N159), .CK(clk), .RN(rstn), .Q(x1_o0[18]) );
  DFFRHQX1 x1_o0_reg_19_ ( .D(N160), .CK(clk), .RN(rstn), .Q(x1_o0[19]) );
  DFFRHQX1 x1_o1_reg_19_ ( .D(x1_o1_tmp[19]), .CK(clk), .RN(rstn), .Q(
        x1_o1[19]) );
  DFFRHQX1 x1_o1_reg_18_ ( .D(x1_o1_tmp[18]), .CK(clk), .RN(rstn), .Q(
        x1_o1[18]) );
  DFFRHQX1 x1_o1_reg_17_ ( .D(x1_o1_tmp[17]), .CK(clk), .RN(rstn), .Q(
        x1_o1[17]) );
  DFFRHQX1 x1_o1_reg_16_ ( .D(x1_o1_tmp[16]), .CK(clk), .RN(rstn), .Q(
        x1_o1[16]) );
  DFFRHQX1 x3_o1_reg_19_ ( .D(N183), .CK(clk), .RN(rstn), .Q(x3_o1[19]) );
  DFFRHQX1 x3_o1_reg_18_ ( .D(N182), .CK(clk), .RN(rstn), .Q(x3_o1[18]) );
  DFFRHQX1 x3_o1_reg_17_ ( .D(N181), .CK(clk), .RN(rstn), .Q(x3_o1[17]) );
  DFFRHQX1 x3_o1_reg_16_ ( .D(N180), .CK(clk), .RN(rstn), .Q(x3_o1[16]) );
  DFFRHQX1 x0_e_reg_18_ ( .D(x0_e_tmp[18]), .CK(clk), .RN(rstn), .Q(x0_e[18])
         );
  DFFRHQX1 x0_e_reg_17_ ( .D(x0_e_tmp[17]), .CK(clk), .RN(rstn), .Q(x0_e[17])
         );
  DFFRHQX1 x0_e_reg_16_ ( .D(x0_e_tmp[16]), .CK(clk), .RN(rstn), .Q(x0_e[16])
         );
  DFFRHQX1 x0_e_reg_15_ ( .D(x0_e_tmp[15]), .CK(clk), .RN(rstn), .Q(x0_e[15])
         );
  DFFRHQX1 e1_reg_20_ ( .D(N275), .CK(clk), .RN(rstn), .Q(e1[20]) );
  DFFRHQX1 e1_reg_19_ ( .D(N274), .CK(clk), .RN(rstn), .Q(e1[19]) );
  DFFRHQX1 e1_reg_18_ ( .D(N273), .CK(clk), .RN(rstn), .Q(e1[18]) );
  DFFRHQX1 e1_reg_17_ ( .D(N272), .CK(clk), .RN(rstn), .Q(e1[17]) );
  DFFRHQX1 e0_reg_20_ ( .D(N207), .CK(clk), .RN(rstn), .Q(e0[20]) );
  DFFRHQX1 e0_reg_19_ ( .D(N206), .CK(clk), .RN(rstn), .Q(e0[19]) );
  DFFRHQX1 e0_reg_18_ ( .D(N205), .CK(clk), .RN(rstn), .Q(e0[18]) );
  DFFRHQX1 e0_reg_17_ ( .D(N204), .CK(clk), .RN(rstn), .Q(e0[17]) );
  DFFRHQX1 x3_o1_tmp2_reg_18_ ( .D(N138), .CK(clk), .RN(rstn), .Q(
        x3_o1_tmp2[18]) );
  DFFRHQX1 x3_o1_tmp2_reg_17_ ( .D(N137), .CK(clk), .RN(rstn), .Q(
        x3_o1_tmp2[17]) );
  DFFRHQX1 x3_o1_tmp2_reg_16_ ( .D(N136), .CK(clk), .RN(rstn), .Q(
        x3_o1_tmp2[16]) );
  DFFRHQX1 x3_o1_tmp2_reg_15_ ( .D(N135), .CK(clk), .RN(rstn), .Q(
        x3_o1_tmp2[15]) );
  DFFRHQX1 x3_o1_tmp2_reg_14_ ( .D(N134), .CK(clk), .RN(rstn), .Q(
        x3_o1_tmp2[14]) );
  DFFRHQX1 x1_o0_tmp2_reg_18_ ( .D(N94), .CK(clk), .RN(rstn), .Q(
        x1_o0_tmp2[18]) );
  DFFRHQX1 x1_o0_tmp2_reg_17_ ( .D(N93), .CK(clk), .RN(rstn), .Q(
        x1_o0_tmp2[17]) );
  DFFRHQX1 x1_o0_tmp2_reg_16_ ( .D(N92), .CK(clk), .RN(rstn), .Q(
        x1_o0_tmp2[16]) );
  DFFRHQX1 x1_o0_tmp2_reg_15_ ( .D(N91), .CK(clk), .RN(rstn), .Q(
        x1_o0_tmp2[15]) );
  DFFRHQX1 x1_o0_tmp2_reg_14_ ( .D(N90), .CK(clk), .RN(rstn), .Q(
        x1_o0_tmp2[14]) );
  DFFRHQX1 x3_o0_reg_19_ ( .D(x3_o0_tmp[19]), .CK(clk), .RN(rstn), .Q(
        x3_o0[19]) );
  DFFRHQX1 x3_o0_reg_18_ ( .D(x3_o0_tmp[18]), .CK(clk), .RN(rstn), .Q(
        x3_o0[18]) );
  DFFRHQX1 x3_o0_reg_17_ ( .D(x3_o0_tmp[17]), .CK(clk), .RN(rstn), .Q(
        x3_o0[17]) );
  DFFRHQX1 x3_o0_reg_16_ ( .D(x3_o0_tmp[16]), .CK(clk), .RN(rstn), .Q(
        x3_o0[16]) );
  DFFRHQX1 x3_o0_reg_15_ ( .D(x3_o0_tmp[15]), .CK(clk), .RN(rstn), .Q(
        x3_o0[15]) );
  DFFRHQX1 x2_e_reg_19_ ( .D(x2_e_tmp[19]), .CK(clk), .RN(rstn), .Q(x2_e[19])
         );
  DFFRHQX1 x2_e_reg_18_ ( .D(x2_e_tmp[18]), .CK(clk), .RN(rstn), .Q(x2_e[18])
         );
  DFFRHQX1 x2_e_reg_17_ ( .D(x2_e_tmp[17]), .CK(clk), .RN(rstn), .Q(x2_e[17])
         );
  DFFRHQX1 x2_e_reg_16_ ( .D(x2_e_tmp[16]), .CK(clk), .RN(rstn), .Q(x2_e[16])
         );
  DFFRHQX1 x2_e_reg_15_ ( .D(x2_e_tmp[15]), .CK(clk), .RN(rstn), .Q(x2_e[15])
         );
  DFFRHQX1 o1_reg_21_ ( .D(N346), .CK(clk), .RN(rstn), .Q(o1[21]) );
  DFFRHQX1 o1_reg_20_ ( .D(N345), .CK(clk), .RN(rstn), .Q(o1[20]) );
  DFFRHQX1 o1_reg_19_ ( .D(N344), .CK(clk), .RN(rstn), .Q(o1[19]) );
  DFFRHQX1 o1_reg_18_ ( .D(N343), .CK(clk), .RN(rstn), .Q(o1[18]) );
  DFFRHQX1 o1_reg_17_ ( .D(N342), .CK(clk), .RN(rstn), .Q(o1[17]) );
  DFFRHQX1 o0_reg_21_ ( .D(N370), .CK(clk), .RN(rstn), .Q(o0[21]) );
  DFFRHQX1 o0_reg_20_ ( .D(N369), .CK(clk), .RN(rstn), .Q(o0[20]) );
  DFFRHQX1 o0_reg_19_ ( .D(N368), .CK(clk), .RN(rstn), .Q(o0[19]) );
  DFFRHQX1 o0_reg_18_ ( .D(N367), .CK(clk), .RN(rstn), .Q(o0[18]) );
  DFFRHQX1 o0_reg_17_ ( .D(N366), .CK(clk), .RN(rstn), .Q(o0[17]) );
  DFFRHQX1 x3_o1_tmp1_reg_14_ ( .D(N111), .CK(clk), .RN(rstn), .Q(
        x3_o1_tmp1[14]) );
  DFFRHQX1 x3_o1_tmp1_reg_13_ ( .D(N110), .CK(clk), .RN(rstn), .Q(
        x3_o1_tmp1[13]) );
  DFFRHQX1 x3_o1_tmp1_reg_12_ ( .D(N109), .CK(clk), .RN(rstn), .Q(
        x3_o1_tmp1[12]) );
  DFFRHQX1 x3_o1_tmp1_reg_11_ ( .D(N108), .CK(clk), .RN(rstn), .Q(
        x3_o1_tmp1[11]) );
  DFFRHQX1 x3_o1_tmp1_reg_10_ ( .D(N107), .CK(clk), .RN(rstn), .Q(
        x3_o1_tmp1[10]) );
  DFFRHQX1 x1_o0_tmp1_reg_14_ ( .D(N67), .CK(clk), .RN(rstn), .Q(
        x1_o0_tmp1[14]) );
  DFFRHQX1 x1_o0_tmp1_reg_13_ ( .D(N66), .CK(clk), .RN(rstn), .Q(
        x1_o0_tmp1[13]) );
  DFFRHQX1 x1_o0_tmp1_reg_12_ ( .D(N65), .CK(clk), .RN(rstn), .Q(
        x1_o0_tmp1[12]) );
  DFFRHQX1 x1_o0_tmp1_reg_11_ ( .D(N64), .CK(clk), .RN(rstn), .Q(
        x1_o0_tmp1[11]) );
  DFFRHQX1 x1_o0_tmp1_reg_10_ ( .D(N63), .CK(clk), .RN(rstn), .Q(
        x1_o0_tmp1[10]) );
  DFFRHQX1 x1_o0_reg_11_ ( .D(N152), .CK(clk), .RN(rstn), .Q(x1_o0[11]) );
  DFFRHQX1 x1_o0_reg_12_ ( .D(N153), .CK(clk), .RN(rstn), .Q(x1_o0[12]) );
  DFFRHQX1 x1_o0_reg_13_ ( .D(N154), .CK(clk), .RN(rstn), .Q(x1_o0[13]) );
  DFFRHQX1 x1_o0_reg_14_ ( .D(N155), .CK(clk), .RN(rstn), .Q(x1_o0[14]) );
  DFFRHQX1 x1_o0_reg_15_ ( .D(N156), .CK(clk), .RN(rstn), .Q(x1_o0[15]) );
  DFFRHQX1 x1_o1_reg_15_ ( .D(x1_o1_tmp[15]), .CK(clk), .RN(rstn), .Q(
        x1_o1[15]) );
  DFFRHQX1 x1_o1_reg_14_ ( .D(x1_o1_tmp[14]), .CK(clk), .RN(rstn), .Q(
        x1_o1[14]) );
  DFFRHQX1 x1_o1_reg_13_ ( .D(x1_o1_tmp[13]), .CK(clk), .RN(rstn), .Q(
        x1_o1[13]) );
  DFFRHQX1 x1_o1_reg_12_ ( .D(x1_o1_tmp[12]), .CK(clk), .RN(rstn), .Q(
        x1_o1[12]) );
  DFFRHQX1 x1_o1_reg_11_ ( .D(x1_o1_tmp[11]), .CK(clk), .RN(rstn), .Q(
        x1_o1[11]) );
  DFFRHQX1 y1_tmp_reg_23_ ( .D(N421), .CK(clk), .RN(rstn), .Q(y1_tmp[23]) );
  DFFRHQX1 y2_tmp_reg_23_ ( .D(N495), .CK(clk), .RN(rstn), .Q(y2_tmp[23]) );
  DFFRHQX1 y0_tmp_reg_23_ ( .D(N396), .CK(clk), .RN(rstn), .Q(y0_tmp[23]) );
  DFFRHQX1 y3_tmp_reg_23_ ( .D(N569), .CK(clk), .RN(rstn), .Q(y3_tmp[23]) );
  DFFRHQX1 y1_tmp_reg_24_ ( .D(N422), .CK(clk), .RN(rstn), .Q(y1_tmp[24]) );
  DFFRHQX1 y2_tmp_reg_24_ ( .D(N496), .CK(clk), .RN(rstn), .Q(y2_tmp[24]) );
  DFFRHQX1 y0_tmp_reg_24_ ( .D(N397), .CK(clk), .RN(rstn), .Q(y0_tmp[24]) );
  DFFRHQX1 y3_tmp_reg_24_ ( .D(N570), .CK(clk), .RN(rstn), .Q(y3_tmp[24]) );
  DFFRHQX1 x3_o1_reg_15_ ( .D(N179), .CK(clk), .RN(rstn), .Q(x3_o1[15]) );
  DFFRHQX1 x3_o1_reg_14_ ( .D(N178), .CK(clk), .RN(rstn), .Q(x3_o1[14]) );
  DFFRHQX1 x3_o1_reg_13_ ( .D(N177), .CK(clk), .RN(rstn), .Q(x3_o1[13]) );
  DFFRHQX1 x3_o1_reg_12_ ( .D(N176), .CK(clk), .RN(rstn), .Q(x3_o1[12]) );
  DFFRHQX1 x0_e_reg_14_ ( .D(x0_e_tmp[14]), .CK(clk), .RN(rstn), .Q(x0_e[14])
         );
  DFFRHQX1 x0_e_reg_13_ ( .D(x0_e_tmp[13]), .CK(clk), .RN(rstn), .Q(x0_e[13])
         );
  DFFRHQX1 x0_e_reg_12_ ( .D(x0_e_tmp[12]), .CK(clk), .RN(rstn), .Q(x0_e[12])
         );
  DFFRHQX1 x0_e_reg_11_ ( .D(x0_e_tmp[11]), .CK(clk), .RN(rstn), .Q(x0_e[11])
         );
  DFFRHQX1 e1_reg_16_ ( .D(N271), .CK(clk), .RN(rstn), .Q(e1[16]) );
  DFFRHQX1 e1_reg_15_ ( .D(N270), .CK(clk), .RN(rstn), .Q(e1[15]) );
  DFFRHQX1 e1_reg_14_ ( .D(N269), .CK(clk), .RN(rstn), .Q(e1[14]) );
  DFFRHQX1 e1_reg_13_ ( .D(N268), .CK(clk), .RN(rstn), .Q(e1[13]) );
  DFFRHQX1 e0_reg_16_ ( .D(N203), .CK(clk), .RN(rstn), .Q(e0[16]) );
  DFFRHQX1 e0_reg_15_ ( .D(N202), .CK(clk), .RN(rstn), .Q(e0[15]) );
  DFFRHQX1 e0_reg_14_ ( .D(N201), .CK(clk), .RN(rstn), .Q(e0[14]) );
  DFFRHQX1 e0_reg_13_ ( .D(N200), .CK(clk), .RN(rstn), .Q(e0[13]) );
  DFFRHQX1 x3_o1_tmp2_reg_13_ ( .D(N133), .CK(clk), .RN(rstn), .Q(
        x3_o1_tmp2[13]) );
  DFFRHQX1 x3_o1_tmp2_reg_12_ ( .D(N132), .CK(clk), .RN(rstn), .Q(
        x3_o1_tmp2[12]) );
  DFFRHQX1 x3_o1_tmp2_reg_11_ ( .D(N131), .CK(clk), .RN(rstn), .Q(
        x3_o1_tmp2[11]) );
  DFFRHQX1 x3_o1_tmp2_reg_10_ ( .D(N130), .CK(clk), .RN(rstn), .Q(
        x3_o1_tmp2[10]) );
  DFFRHQX1 x1_o0_tmp2_reg_13_ ( .D(N89), .CK(clk), .RN(rstn), .Q(
        x1_o0_tmp2[13]) );
  DFFRHQX1 x1_o0_tmp2_reg_12_ ( .D(N88), .CK(clk), .RN(rstn), .Q(
        x1_o0_tmp2[12]) );
  DFFRHQX1 x1_o0_tmp2_reg_11_ ( .D(N87), .CK(clk), .RN(rstn), .Q(
        x1_o0_tmp2[11]) );
  DFFRHQX1 x1_o0_tmp2_reg_10_ ( .D(N86), .CK(clk), .RN(rstn), .Q(
        x1_o0_tmp2[10]) );
  DFFRHQX1 x3_o0_reg_14_ ( .D(x3_o0_tmp[14]), .CK(clk), .RN(rstn), .Q(
        x3_o0[14]) );
  DFFRHQX1 x3_o0_reg_13_ ( .D(x3_o0_tmp[13]), .CK(clk), .RN(rstn), .Q(
        x3_o0[13]) );
  DFFRHQX1 x3_o0_reg_12_ ( .D(x3_o0_tmp[12]), .CK(clk), .RN(rstn), .Q(
        x3_o0[12]) );
  DFFRHQX1 x3_o0_reg_11_ ( .D(x3_o0_tmp[11]), .CK(clk), .RN(rstn), .Q(
        x3_o0[11]) );
  DFFRHQX1 x2_e_reg_14_ ( .D(x2_e_tmp[14]), .CK(clk), .RN(rstn), .Q(x2_e[14])
         );
  DFFRHQX1 x2_e_reg_13_ ( .D(x2_e_tmp[13]), .CK(clk), .RN(rstn), .Q(x2_e[13])
         );
  DFFRHQX1 x2_e_reg_12_ ( .D(x2_e_tmp[12]), .CK(clk), .RN(rstn), .Q(x2_e[12])
         );
  DFFRHQX1 x2_e_reg_11_ ( .D(x2_e_tmp[11]), .CK(clk), .RN(rstn), .Q(x2_e[11])
         );
  DFFRHQX1 o1_reg_16_ ( .D(N341), .CK(clk), .RN(rstn), .Q(o1[16]) );
  DFFRHQX1 o1_reg_15_ ( .D(N340), .CK(clk), .RN(rstn), .Q(o1[15]) );
  DFFRHQX1 o1_reg_14_ ( .D(N339), .CK(clk), .RN(rstn), .Q(o1[14]) );
  DFFRHQX1 o1_reg_13_ ( .D(N338), .CK(clk), .RN(rstn), .Q(o1[13]) );
  DFFRHQX1 o0_reg_16_ ( .D(N365), .CK(clk), .RN(rstn), .Q(o0[16]) );
  DFFRHQX1 o0_reg_15_ ( .D(N364), .CK(clk), .RN(rstn), .Q(o0[15]) );
  DFFRHQX1 o0_reg_14_ ( .D(N363), .CK(clk), .RN(rstn), .Q(o0[14]) );
  DFFRHQX1 o0_reg_13_ ( .D(N362), .CK(clk), .RN(rstn), .Q(o0[13]) );
  DFFRHQX1 x3_o1_tmp1_reg_9_ ( .D(N106), .CK(clk), .RN(rstn), .Q(x3_o1_tmp1[9]) );
  DFFRHQX1 x3_o1_tmp1_reg_8_ ( .D(N105), .CK(clk), .RN(rstn), .Q(x3_o1_tmp1[8]) );
  DFFRHQX1 x3_o1_tmp1_reg_7_ ( .D(N104), .CK(clk), .RN(rstn), .Q(x3_o1_tmp1[7]) );
  DFFRHQX1 x3_o1_tmp1_reg_6_ ( .D(N103), .CK(clk), .RN(rstn), .Q(x3_o1_tmp1[6]) );
  DFFRHQX1 x1_o0_tmp1_reg_9_ ( .D(N62), .CK(clk), .RN(rstn), .Q(x1_o0_tmp1[9])
         );
  DFFRHQX1 x1_o0_tmp1_reg_8_ ( .D(N61), .CK(clk), .RN(rstn), .Q(x1_o0_tmp1[8])
         );
  DFFRHQX1 x1_o0_tmp1_reg_7_ ( .D(N60), .CK(clk), .RN(rstn), .Q(x1_o0_tmp1[7])
         );
  DFFRHQX1 x1_o0_tmp1_reg_6_ ( .D(N59), .CK(clk), .RN(rstn), .Q(x1_o0_tmp1[6])
         );
  DFFRHQX1 x1_o0_reg_7_ ( .D(N148), .CK(clk), .RN(rstn), .Q(x1_o0[7]) );
  DFFRHQX1 x1_o0_reg_8_ ( .D(N149), .CK(clk), .RN(rstn), .Q(x1_o0[8]) );
  DFFRHQX1 x1_o0_reg_9_ ( .D(N150), .CK(clk), .RN(rstn), .Q(x1_o0[9]) );
  DFFRHQX1 x1_o0_reg_10_ ( .D(N151), .CK(clk), .RN(rstn), .Q(x1_o0[10]) );
  DFFRHQX1 x1_o1_reg_10_ ( .D(x1_o1_tmp[10]), .CK(clk), .RN(rstn), .Q(
        x1_o1[10]) );
  DFFRHQX1 x1_o1_reg_9_ ( .D(x1_o1_tmp[9]), .CK(clk), .RN(rstn), .Q(x1_o1[9])
         );
  DFFRHQX1 x1_o1_reg_8_ ( .D(x1_o1_tmp[8]), .CK(clk), .RN(rstn), .Q(x1_o1[8])
         );
  DFFRHQX1 x1_o1_reg_7_ ( .D(x1_o1_tmp[7]), .CK(clk), .RN(rstn), .Q(x1_o1[7])
         );
  DFFRHQX1 y1_tmp_reg_22_ ( .D(N420), .CK(clk), .RN(rstn), .Q(y1_tmp[22]) );
  DFFRHQX1 y1_tmp_reg_21_ ( .D(N419), .CK(clk), .RN(rstn), .Q(y1_tmp[21]) );
  DFFRHQX1 y1_tmp_reg_20_ ( .D(N418), .CK(clk), .RN(rstn), .Q(y1_tmp[20]) );
  DFFRHQX1 y1_tmp_reg_19_ ( .D(N417), .CK(clk), .RN(rstn), .Q(y1_tmp[19]) );
  DFFRHQX1 y2_tmp_reg_22_ ( .D(N494), .CK(clk), .RN(rstn), .Q(y2_tmp[22]) );
  DFFRHQX1 y2_tmp_reg_21_ ( .D(N493), .CK(clk), .RN(rstn), .Q(y2_tmp[21]) );
  DFFRHQX1 y2_tmp_reg_20_ ( .D(N492), .CK(clk), .RN(rstn), .Q(y2_tmp[20]) );
  DFFRHQX1 y2_tmp_reg_19_ ( .D(N491), .CK(clk), .RN(rstn), .Q(y2_tmp[19]) );
  DFFRHQX1 y0_tmp_reg_19_ ( .D(N392), .CK(clk), .RN(rstn), .Q(y0_tmp[19]) );
  DFFRHQX1 y0_tmp_reg_20_ ( .D(N393), .CK(clk), .RN(rstn), .Q(y0_tmp[20]) );
  DFFRHQX1 y0_tmp_reg_21_ ( .D(N394), .CK(clk), .RN(rstn), .Q(y0_tmp[21]) );
  DFFRHQX1 y0_tmp_reg_22_ ( .D(N395), .CK(clk), .RN(rstn), .Q(y0_tmp[22]) );
  DFFRHQX1 y3_tmp_reg_19_ ( .D(N565), .CK(clk), .RN(rstn), .Q(y3_tmp[19]) );
  DFFRHQX1 y3_tmp_reg_20_ ( .D(N566), .CK(clk), .RN(rstn), .Q(y3_tmp[20]) );
  DFFRHQX1 y3_tmp_reg_21_ ( .D(N567), .CK(clk), .RN(rstn), .Q(y3_tmp[21]) );
  DFFRHQX1 y3_tmp_reg_22_ ( .D(N568), .CK(clk), .RN(rstn), .Q(y3_tmp[22]) );
  DFFRHQX1 x0_e_reg_6_ ( .D(x0_e_tmp[6]), .CK(clk), .RN(rstn), .Q(x0_e[6]) );
  DFFRHQX1 idct4_ready_reg ( .D(idct4_ready_delay3), .CK(clk), .RN(rstn), .Q(
        idct4_ready) );
  DFFRHQX1 x3_o1_reg_11_ ( .D(N175), .CK(clk), .RN(rstn), .Q(x3_o1[11]) );
  DFFRHQX1 x3_o1_reg_10_ ( .D(N174), .CK(clk), .RN(rstn), .Q(x3_o1[10]) );
  DFFRHQX1 x3_o1_reg_9_ ( .D(N173), .CK(clk), .RN(rstn), .Q(x3_o1[9]) );
  DFFRHQX1 x3_o1_reg_8_ ( .D(N172), .CK(clk), .RN(rstn), .Q(x3_o1[8]) );
  DFFRHQX1 x3_o1_reg_7_ ( .D(N171), .CK(clk), .RN(rstn), .Q(x3_o1[7]) );
  DFFRHQX1 x0_e_reg_10_ ( .D(x0_e_tmp[10]), .CK(clk), .RN(rstn), .Q(x0_e[10])
         );
  DFFRHQX1 x0_e_reg_9_ ( .D(x0_e_tmp[9]), .CK(clk), .RN(rstn), .Q(x0_e[9]) );
  DFFRHQX1 x0_e_reg_8_ ( .D(x0_e_tmp[8]), .CK(clk), .RN(rstn), .Q(x0_e[8]) );
  DFFRHQX1 x0_e_reg_7_ ( .D(x0_e_tmp[7]), .CK(clk), .RN(rstn), .Q(x0_e[7]) );
  DFFRHQX1 e1_reg_12_ ( .D(N267), .CK(clk), .RN(rstn), .Q(e1[12]) );
  DFFRHQX1 e1_reg_11_ ( .D(N266), .CK(clk), .RN(rstn), .Q(e1[11]) );
  DFFRHQX1 e1_reg_10_ ( .D(N265), .CK(clk), .RN(rstn), .Q(e1[10]) );
  DFFRHQX1 e1_reg_9_ ( .D(N264), .CK(clk), .RN(rstn), .Q(e1[9]) );
  DFFRHQX1 e1_reg_8_ ( .D(N263), .CK(clk), .RN(rstn), .Q(e1[8]) );
  DFFRHQX1 e0_reg_12_ ( .D(N199), .CK(clk), .RN(rstn), .Q(e0[12]) );
  DFFRHQX1 e0_reg_11_ ( .D(N198), .CK(clk), .RN(rstn), .Q(e0[11]) );
  DFFRHQX1 e0_reg_10_ ( .D(N197), .CK(clk), .RN(rstn), .Q(e0[10]) );
  DFFRHQX1 e0_reg_9_ ( .D(N196), .CK(clk), .RN(rstn), .Q(e0[9]) );
  DFFRHQX1 e0_reg_8_ ( .D(N195), .CK(clk), .RN(rstn), .Q(e0[8]) );
  DFFRHQX1 x3_o1_tmp2_reg_9_ ( .D(N129), .CK(clk), .RN(rstn), .Q(x3_o1_tmp2[9]) );
  DFFRHQX1 x3_o1_tmp2_reg_8_ ( .D(N128), .CK(clk), .RN(rstn), .Q(x3_o1_tmp2[8]) );
  DFFRHQX1 x3_o1_tmp2_reg_7_ ( .D(N127), .CK(clk), .RN(rstn), .Q(x3_o1_tmp2[7]) );
  DFFRHQX1 x3_o1_tmp2_reg_6_ ( .D(N126), .CK(clk), .RN(rstn), .Q(x3_o1_tmp2[6]) );
  DFFRHQX1 x1_o0_tmp2_reg_9_ ( .D(N85), .CK(clk), .RN(rstn), .Q(x1_o0_tmp2[9])
         );
  DFFRHQX1 x1_o0_tmp2_reg_8_ ( .D(N84), .CK(clk), .RN(rstn), .Q(x1_o0_tmp2[8])
         );
  DFFRHQX1 x1_o0_tmp2_reg_7_ ( .D(N83), .CK(clk), .RN(rstn), .Q(x1_o0_tmp2[7])
         );
  DFFRHQX1 x1_o0_tmp2_reg_6_ ( .D(N82), .CK(clk), .RN(rstn), .Q(x1_o0_tmp2[6])
         );
  DFFRHQX1 x3_o0_reg_10_ ( .D(x3_o0_tmp[10]), .CK(clk), .RN(rstn), .Q(
        x3_o0[10]) );
  DFFRHQX1 x3_o0_reg_9_ ( .D(x3_o0_tmp[9]), .CK(clk), .RN(rstn), .Q(x3_o0[9])
         );
  DFFRHQX1 x3_o0_reg_8_ ( .D(x3_o0_tmp[8]), .CK(clk), .RN(rstn), .Q(x3_o0[8])
         );
  DFFRHQX1 x3_o0_reg_7_ ( .D(x3_o0_tmp[7]), .CK(clk), .RN(rstn), .Q(x3_o0[7])
         );
  DFFRHQX1 x2_e_reg_6_ ( .D(x2_e_tmp[6]), .CK(clk), .RN(rstn), .Q(x2_e[6]) );
  DFFRHQX1 x2_e_reg_10_ ( .D(x2_e_tmp[10]), .CK(clk), .RN(rstn), .Q(x2_e[10])
         );
  DFFRHQX1 x2_e_reg_9_ ( .D(x2_e_tmp[9]), .CK(clk), .RN(rstn), .Q(x2_e[9]) );
  DFFRHQX1 x2_e_reg_8_ ( .D(x2_e_tmp[8]), .CK(clk), .RN(rstn), .Q(x2_e[8]) );
  DFFRHQX1 x2_e_reg_7_ ( .D(x2_e_tmp[7]), .CK(clk), .RN(rstn), .Q(x2_e[7]) );
  DFFRHQX1 o1_reg_12_ ( .D(N337), .CK(clk), .RN(rstn), .Q(o1[12]) );
  DFFRHQX1 o1_reg_11_ ( .D(N336), .CK(clk), .RN(rstn), .Q(o1[11]) );
  DFFRHQX1 o1_reg_10_ ( .D(N335), .CK(clk), .RN(rstn), .Q(o1[10]) );
  DFFRHQX1 o1_reg_9_ ( .D(N334), .CK(clk), .RN(rstn), .Q(o1[9]) );
  DFFRHQX1 o0_reg_12_ ( .D(N361), .CK(clk), .RN(rstn), .Q(o0[12]) );
  DFFRHQX1 o0_reg_11_ ( .D(N360), .CK(clk), .RN(rstn), .Q(o0[11]) );
  DFFRHQX1 o0_reg_10_ ( .D(N359), .CK(clk), .RN(rstn), .Q(o0[10]) );
  DFFRHQX1 o0_reg_9_ ( .D(N358), .CK(clk), .RN(rstn), .Q(o0[9]) );
  DFFRHQX1 x3_o1_tmp1_reg_5_ ( .D(x3[5]), .CK(clk), .RN(rstn), .Q(
        x3_o1_tmp1[5]) );
  DFFRHQX1 x3_o1_tmp1_reg_4_ ( .D(x3[4]), .CK(clk), .RN(rstn), .Q(
        x3_o1_tmp1[4]) );
  DFFRHQX1 x3_o1_tmp1_reg_3_ ( .D(x3[3]), .CK(clk), .RN(rstn), .Q(
        x3_o1_tmp1[3]) );
  DFFRHQX1 x3_o1_tmp1_reg_2_ ( .D(x3[2]), .CK(clk), .RN(rstn), .Q(
        x3_o1_tmp1[2]) );
  DFFRHQX1 x1_o0_tmp1_reg_5_ ( .D(x1[5]), .CK(clk), .RN(rstn), .Q(
        x1_o0_tmp1[5]) );
  DFFRHQX1 x1_o0_tmp1_reg_4_ ( .D(x1[4]), .CK(clk), .RN(rstn), .Q(
        x1_o0_tmp1[4]) );
  DFFRHQX1 x1_o0_tmp1_reg_3_ ( .D(x1[3]), .CK(clk), .RN(rstn), .Q(
        x1_o0_tmp1[3]) );
  DFFRHQX1 x1_o0_tmp1_reg_2_ ( .D(x1[2]), .CK(clk), .RN(rstn), .Q(
        x1_o0_tmp1[2]) );
  DFFRHQX1 x1_o0_reg_3_ ( .D(N144), .CK(clk), .RN(rstn), .Q(x1_o0[3]) );
  DFFRHQX1 x1_o0_reg_4_ ( .D(N145), .CK(clk), .RN(rstn), .Q(x1_o0[4]) );
  DFFRHQX1 x1_o0_reg_5_ ( .D(N146), .CK(clk), .RN(rstn), .Q(x1_o0[5]) );
  DFFRHQX1 x1_o0_reg_6_ ( .D(N147), .CK(clk), .RN(rstn), .Q(x1_o0[6]) );
  DFFRHQX1 x1_o1_reg_6_ ( .D(x1_o1_tmp[6]), .CK(clk), .RN(rstn), .Q(x1_o1[6])
         );
  DFFRHQX1 x1_o1_reg_5_ ( .D(x1_o1_tmp[5]), .CK(clk), .RN(rstn), .Q(x1_o1[5])
         );
  DFFRHQX1 x1_o1_reg_4_ ( .D(x1_o1_tmp[4]), .CK(clk), .RN(rstn), .Q(x1_o1[4])
         );
  DFFRHQX1 x1_o1_reg_3_ ( .D(x1_o1_tmp[3]), .CK(clk), .RN(rstn), .Q(x1_o1[3])
         );
  DFFRHQX1 y1_tmp_reg_18_ ( .D(N416), .CK(clk), .RN(rstn), .Q(y1_tmp[18]) );
  DFFRHQX1 y2_tmp_reg_18_ ( .D(N490), .CK(clk), .RN(rstn), .Q(y2_tmp[18]) );
  DFFRHQX1 y0_tmp_reg_18_ ( .D(N391), .CK(clk), .RN(rstn), .Q(y0_tmp[18]) );
  DFFRHQX1 y3_tmp_reg_18_ ( .D(N564), .CK(clk), .RN(rstn), .Q(y3_tmp[18]) );
  DFFRHQX1 x3_o1_reg_6_ ( .D(N170), .CK(clk), .RN(rstn), .Q(x3_o1[6]) );
  DFFRHQX1 x3_o1_reg_5_ ( .D(N169), .CK(clk), .RN(rstn), .Q(x3_o1[5]) );
  DFFRHQX1 x3_o1_reg_4_ ( .D(N168), .CK(clk), .RN(rstn), .Q(x3_o1[4]) );
  DFFRHQX1 x3_o1_reg_3_ ( .D(N167), .CK(clk), .RN(rstn), .Q(x3_o1[3]) );
  DFFRHQX1 e1_reg_7_ ( .D(N262), .CK(clk), .RN(rstn), .Q(e1[7]) );
  DFFRHQX1 e1_reg_6_ ( .D(N261), .CK(clk), .RN(rstn), .Q(e1[6]) );
  DFFRHQX1 e0_reg_7_ ( .D(N194), .CK(clk), .RN(rstn), .Q(e0[7]) );
  DFFRHQX1 e0_reg_6_ ( .D(N193), .CK(clk), .RN(rstn), .Q(e0[6]) );
  DFFRHQX1 y1_tmp_reg_17_ ( .D(N415), .CK(clk), .RN(rstn), .Q(y1_tmp[17]) );
  DFFRHQX1 y1_tmp_reg_16_ ( .D(N414), .CK(clk), .RN(rstn), .Q(y1_tmp[16]) );
  DFFRHQX1 y1_tmp_reg_15_ ( .D(N413), .CK(clk), .RN(rstn), .Q(y1_tmp[15]) );
  DFFRHQX1 y2_tmp_reg_17_ ( .D(N489), .CK(clk), .RN(rstn), .Q(y2_tmp[17]) );
  DFFRHQX1 y2_tmp_reg_16_ ( .D(N488), .CK(clk), .RN(rstn), .Q(y2_tmp[16]) );
  DFFRHQX1 y2_tmp_reg_15_ ( .D(N487), .CK(clk), .RN(rstn), .Q(y2_tmp[15]) );
  DFFRHQX1 y0_tmp_reg_15_ ( .D(N388), .CK(clk), .RN(rstn), .Q(y0_tmp[15]) );
  DFFRHQX1 y0_tmp_reg_16_ ( .D(N389), .CK(clk), .RN(rstn), .Q(y0_tmp[16]) );
  DFFRHQX1 y0_tmp_reg_17_ ( .D(N390), .CK(clk), .RN(rstn), .Q(y0_tmp[17]) );
  DFFRHQX1 y3_tmp_reg_15_ ( .D(N561), .CK(clk), .RN(rstn), .Q(y3_tmp[15]) );
  DFFRHQX1 y3_tmp_reg_16_ ( .D(N562), .CK(clk), .RN(rstn), .Q(y3_tmp[16]) );
  DFFRHQX1 y3_tmp_reg_17_ ( .D(N563), .CK(clk), .RN(rstn), .Q(y3_tmp[17]) );
  DFFRHQX1 x3_o1_tmp2_reg_5_ ( .D(N125), .CK(clk), .RN(rstn), .Q(x3_o1_tmp2[5]) );
  DFFRHQX1 x3_o1_tmp2_reg_4_ ( .D(N124), .CK(clk), .RN(rstn), .Q(x3_o1_tmp2[4]) );
  DFFRHQX1 x3_o1_tmp2_reg_3_ ( .D(x3[2]), .CK(clk), .RN(rstn), .Q(
        x3_o1_tmp2[3]) );
  DFFRHQX1 x3_o1_tmp2_reg_2_ ( .D(x3[1]), .CK(clk), .RN(rstn), .Q(
        x3_o1_tmp2[2]) );
  DFFRHQX1 x3_o1_tmp2_reg_1_ ( .D(x3[0]), .CK(clk), .RN(rstn), .Q(
        x3_o1_tmp2[1]) );
  DFFRHQX1 x1_o0_tmp2_reg_5_ ( .D(N81), .CK(clk), .RN(rstn), .Q(x1_o0_tmp2[5])
         );
  DFFRHQX1 x1_o0_tmp2_reg_4_ ( .D(N80), .CK(clk), .RN(rstn), .Q(x1_o0_tmp2[4])
         );
  DFFRHQX1 x1_o0_tmp2_reg_3_ ( .D(x1[2]), .CK(clk), .RN(rstn), .Q(
        x1_o0_tmp2[3]) );
  DFFRHQX1 x1_o0_tmp2_reg_2_ ( .D(x1[1]), .CK(clk), .RN(rstn), .Q(
        x1_o0_tmp2[2]) );
  DFFRHQX1 x1_o0_tmp2_reg_1_ ( .D(x1[0]), .CK(clk), .RN(rstn), .Q(
        x1_o0_tmp2[1]) );
  DFFRHQX1 x3_o0_reg_6_ ( .D(x3_o0_tmp[6]), .CK(clk), .RN(rstn), .Q(x3_o0[6])
         );
  DFFRHQX1 x3_o0_reg_5_ ( .D(x3_o0_tmp[5]), .CK(clk), .RN(rstn), .Q(x3_o0[5])
         );
  DFFRHQX1 x3_o0_reg_4_ ( .D(x3_o0_tmp[4]), .CK(clk), .RN(rstn), .Q(x3_o0[4])
         );
  DFFRHQX1 x3_o0_reg_3_ ( .D(x3_o0_tmp[3]), .CK(clk), .RN(rstn), .Q(x3_o0[3])
         );
  DFFRHQX1 x3_o0_reg_2_ ( .D(x3_o0_tmp[2]), .CK(clk), .RN(rstn), .Q(x3_o0[2])
         );
  DFFRHQX1 o1_reg_8_ ( .D(N333), .CK(clk), .RN(rstn), .Q(o1[8]) );
  DFFRHQX1 o1_reg_7_ ( .D(N332), .CK(clk), .RN(rstn), .Q(o1[7]) );
  DFFRHQX1 o1_reg_6_ ( .D(N331), .CK(clk), .RN(rstn), .Q(o1[6]) );
  DFFRHQX1 o1_reg_5_ ( .D(N330), .CK(clk), .RN(rstn), .Q(o1[5]) );
  DFFRHQX1 o1_reg_4_ ( .D(N329), .CK(clk), .RN(rstn), .Q(o1[4]) );
  DFFRHQX1 o0_reg_8_ ( .D(N357), .CK(clk), .RN(rstn), .Q(o0[8]) );
  DFFRHQX1 o0_reg_7_ ( .D(N356), .CK(clk), .RN(rstn), .Q(o0[7]) );
  DFFRHQX1 o0_reg_6_ ( .D(N355), .CK(clk), .RN(rstn), .Q(o0[6]) );
  DFFRHQX1 o0_reg_5_ ( .D(N354), .CK(clk), .RN(rstn), .Q(o0[5]) );
  DFFRHQX1 o0_reg_4_ ( .D(N353), .CK(clk), .RN(rstn), .Q(o0[4]) );
  DFFRHQX1 x3_o1_tmp1_reg_1_ ( .D(x3[1]), .CK(clk), .RN(rstn), .Q(
        x3_o1_tmp1[1]) );
  DFFRHQX1 x1_o0_tmp1_reg_1_ ( .D(x1[1]), .CK(clk), .RN(rstn), .Q(
        x1_o0_tmp1[1]) );
  DFFRHQX1 x1_o0_reg_1_ ( .D(N142), .CK(clk), .RN(rstn), .Q(x1_o0[1]) );
  DFFRHQX1 x1_o0_reg_2_ ( .D(N143), .CK(clk), .RN(rstn), .Q(x1_o0[2]) );
  DFFRHQX1 x1_o1_reg_2_ ( .D(x1_o1_tmp[2]), .CK(clk), .RN(rstn), .Q(x1_o1[2])
         );
  DFFRHQX1 y1_tmp_reg_5_ ( .D(N403), .CK(clk), .RN(rstn), .Q(y1_tmp[5]) );
  DFFRHQX1 y1_tmp_reg_4_ ( .D(N402), .CK(clk), .RN(rstn), .Q(y1_tmp[4]) );
  DFFRHQX1 y1_tmp_reg_3_ ( .D(N401), .CK(clk), .RN(rstn), .Q(y1_tmp[3]) );
  DFFRHQX1 y1_tmp_reg_2_ ( .D(N400), .CK(clk), .RN(rstn), .Q(y1_tmp[2]) );
  DFFRHQX1 y2_tmp_reg_5_ ( .D(N477), .CK(clk), .RN(rstn), .Q(y2_tmp[5]) );
  DFFRHQX1 y2_tmp_reg_4_ ( .D(N476), .CK(clk), .RN(rstn), .Q(y2_tmp[4]) );
  DFFRHQX1 y2_tmp_reg_3_ ( .D(N475), .CK(clk), .RN(rstn), .Q(y2_tmp[3]) );
  DFFRHQX1 y2_tmp_reg_2_ ( .D(N474), .CK(clk), .RN(rstn), .Q(y2_tmp[2]) );
  DFFRHQX1 y0_tmp_reg_2_ ( .D(N375), .CK(clk), .RN(rstn), .Q(y0_tmp[2]) );
  DFFRHQX1 y0_tmp_reg_3_ ( .D(N376), .CK(clk), .RN(rstn), .Q(y0_tmp[3]) );
  DFFRHQX1 y0_tmp_reg_4_ ( .D(N377), .CK(clk), .RN(rstn), .Q(y0_tmp[4]) );
  DFFRHQX1 y0_tmp_reg_5_ ( .D(N378), .CK(clk), .RN(rstn), .Q(y0_tmp[5]) );
  DFFRHQX1 y3_tmp_reg_2_ ( .D(N548), .CK(clk), .RN(rstn), .Q(y3_tmp[2]) );
  DFFRHQX1 y3_tmp_reg_3_ ( .D(N549), .CK(clk), .RN(rstn), .Q(y3_tmp[3]) );
  DFFRHQX1 y3_tmp_reg_4_ ( .D(N550), .CK(clk), .RN(rstn), .Q(y3_tmp[4]) );
  DFFRHQX1 y3_tmp_reg_5_ ( .D(N551), .CK(clk), .RN(rstn), .Q(y3_tmp[5]) );
  DFFRHQX1 x3_o1_reg_2_ ( .D(N166), .CK(clk), .RN(rstn), .Q(x3_o1[2]) );
  DFFRHQX1 x3_o1_reg_1_ ( .D(N165), .CK(clk), .RN(rstn), .Q(x3_o1[1]) );
  DFFRHQX1 x3_o1_reg_0_ ( .D(N164), .CK(clk), .RN(rstn), .Q(x3_o1[0]) );
  DFFRHQX1 y1_tmp_reg_14_ ( .D(N412), .CK(clk), .RN(rstn), .Q(y1_tmp[14]) );
  DFFRHQX1 y1_tmp_reg_13_ ( .D(N411), .CK(clk), .RN(rstn), .Q(y1_tmp[13]) );
  DFFRHQX1 y1_tmp_reg_12_ ( .D(N410), .CK(clk), .RN(rstn), .Q(y1_tmp[12]) );
  DFFRHQX1 y1_tmp_reg_11_ ( .D(N409), .CK(clk), .RN(rstn), .Q(y1_tmp[11]) );
  DFFRHQX1 y2_tmp_reg_14_ ( .D(N486), .CK(clk), .RN(rstn), .Q(y2_tmp[14]) );
  DFFRHQX1 y2_tmp_reg_13_ ( .D(N485), .CK(clk), .RN(rstn), .Q(y2_tmp[13]) );
  DFFRHQX1 y2_tmp_reg_12_ ( .D(N484), .CK(clk), .RN(rstn), .Q(y2_tmp[12]) );
  DFFRHQX1 y2_tmp_reg_11_ ( .D(N483), .CK(clk), .RN(rstn), .Q(y2_tmp[11]) );
  DFFRHQX1 y0_tmp_reg_11_ ( .D(N384), .CK(clk), .RN(rstn), .Q(y0_tmp[11]) );
  DFFRHQX1 y0_tmp_reg_12_ ( .D(N385), .CK(clk), .RN(rstn), .Q(y0_tmp[12]) );
  DFFRHQX1 y0_tmp_reg_13_ ( .D(N386), .CK(clk), .RN(rstn), .Q(y0_tmp[13]) );
  DFFRHQX1 y0_tmp_reg_14_ ( .D(N387), .CK(clk), .RN(rstn), .Q(y0_tmp[14]) );
  DFFRHQX1 y3_tmp_reg_11_ ( .D(N557), .CK(clk), .RN(rstn), .Q(y3_tmp[11]) );
  DFFRHQX1 y3_tmp_reg_12_ ( .D(N558), .CK(clk), .RN(rstn), .Q(y3_tmp[12]) );
  DFFRHQX1 y3_tmp_reg_13_ ( .D(N559), .CK(clk), .RN(rstn), .Q(y3_tmp[13]) );
  DFFRHQX1 y3_tmp_reg_14_ ( .D(N560), .CK(clk), .RN(rstn), .Q(y3_tmp[14]) );
  DFFRHQX1 o1_reg_0_ ( .D(N325), .CK(clk), .RN(rstn), .Q(o1[0]) );
  DFFRHQX1 o0_reg_0_ ( .D(N349), .CK(clk), .RN(rstn), .Q(o0[0]) );
  DFFRHQX1 o1_reg_3_ ( .D(N328), .CK(clk), .RN(rstn), .Q(o1[3]) );
  DFFRHQX1 o1_reg_2_ ( .D(N327), .CK(clk), .RN(rstn), .Q(o1[2]) );
  DFFRHQX1 o1_reg_1_ ( .D(N326), .CK(clk), .RN(rstn), .Q(o1[1]) );
  DFFRHQX1 o0_reg_3_ ( .D(N352), .CK(clk), .RN(rstn), .Q(o0[3]) );
  DFFRHQX1 o0_reg_2_ ( .D(N351), .CK(clk), .RN(rstn), .Q(o0[2]) );
  DFFRHQX1 o0_reg_1_ ( .D(N350), .CK(clk), .RN(rstn), .Q(o0[1]) );
  DFFRHQX1 y1_tmp_reg_1_ ( .D(N399), .CK(clk), .RN(rstn), .Q(y1_tmp[1]) );
  DFFRHQX1 y1_tmp_reg_0_ ( .D(N398), .CK(clk), .RN(rstn), .Q(y1_tmp[0]) );
  DFFRHQX1 y2_tmp_reg_1_ ( .D(N473), .CK(clk), .RN(rstn), .Q(y2_tmp[1]) );
  DFFRHQX1 y2_tmp_reg_0_ ( .D(N472), .CK(clk), .RN(rstn), .Q(y2_tmp[0]) );
  DFFRHQX1 y0_tmp_reg_0_ ( .D(N373), .CK(clk), .RN(rstn), .Q(y0_tmp[0]) );
  DFFRHQX1 y0_tmp_reg_1_ ( .D(N374), .CK(clk), .RN(rstn), .Q(y0_tmp[1]) );
  DFFRHQX1 y3_tmp_reg_0_ ( .D(N546), .CK(clk), .RN(rstn), .Q(y3_tmp[0]) );
  DFFRHQX1 y3_tmp_reg_1_ ( .D(N547), .CK(clk), .RN(rstn), .Q(y3_tmp[1]) );
  DFFRHQX1 y1_tmp_reg_10_ ( .D(N408), .CK(clk), .RN(rstn), .Q(y1_tmp[10]) );
  DFFRHQX1 y1_tmp_reg_9_ ( .D(N407), .CK(clk), .RN(rstn), .Q(y1_tmp[9]) );
  DFFRHQX1 y1_tmp_reg_8_ ( .D(N406), .CK(clk), .RN(rstn), .Q(y1_tmp[8]) );
  DFFRHQX1 y1_tmp_reg_7_ ( .D(N405), .CK(clk), .RN(rstn), .Q(y1_tmp[7]) );
  DFFRHQX1 y2_tmp_reg_10_ ( .D(N482), .CK(clk), .RN(rstn), .Q(y2_tmp[10]) );
  DFFRHQX1 y2_tmp_reg_9_ ( .D(N481), .CK(clk), .RN(rstn), .Q(y2_tmp[9]) );
  DFFRHQX1 y2_tmp_reg_8_ ( .D(N480), .CK(clk), .RN(rstn), .Q(y2_tmp[8]) );
  DFFRHQX1 y2_tmp_reg_7_ ( .D(N479), .CK(clk), .RN(rstn), .Q(y2_tmp[7]) );
  DFFRHQX1 y0_tmp_reg_7_ ( .D(N380), .CK(clk), .RN(rstn), .Q(y0_tmp[7]) );
  DFFRHQX1 y0_tmp_reg_8_ ( .D(N381), .CK(clk), .RN(rstn), .Q(y0_tmp[8]) );
  DFFRHQX1 y0_tmp_reg_9_ ( .D(N382), .CK(clk), .RN(rstn), .Q(y0_tmp[9]) );
  DFFRHQX1 y0_tmp_reg_10_ ( .D(N383), .CK(clk), .RN(rstn), .Q(y0_tmp[10]) );
  DFFRHQX1 y3_tmp_reg_7_ ( .D(N553), .CK(clk), .RN(rstn), .Q(y3_tmp[7]) );
  DFFRHQX1 y3_tmp_reg_8_ ( .D(N554), .CK(clk), .RN(rstn), .Q(y3_tmp[8]) );
  DFFRHQX1 y3_tmp_reg_9_ ( .D(N555), .CK(clk), .RN(rstn), .Q(y3_tmp[9]) );
  DFFRHQX1 y3_tmp_reg_10_ ( .D(N556), .CK(clk), .RN(rstn), .Q(y3_tmp[10]) );
  DFFRHQX1 y1_tmp_reg_6_ ( .D(N404), .CK(clk), .RN(rstn), .Q(y1_tmp[6]) );
  DFFRHQX1 y2_tmp_reg_6_ ( .D(N478), .CK(clk), .RN(rstn), .Q(y2_tmp[6]) );
  DFFRHQX1 y0_tmp_reg_6_ ( .D(N379), .CK(clk), .RN(rstn), .Q(y0_tmp[6]) );
  DFFRHQX1 y3_tmp_reg_6_ ( .D(N552), .CK(clk), .RN(rstn), .Q(y3_tmp[6]) );
  DFFRHQX1 mode_delay2_reg_1_ ( .D(mode_delay1[1]), .CK(clk), .RN(rstn), .Q(
        mode_delay2[1]) );
  DFFRHQX1 mode_delay2_reg_0_ ( .D(mode_delay1[0]), .CK(clk), .RN(rstn), .Q(
        mode_delay2[0]) );
  DFFRHQX1 x1_o1_tmp_reg_21_ ( .D(N30), .CK(clk), .RN(rstn), .Q(x1_o1_tmp[21])
         );
  DFFRHQX1 x1_o1_tmp_reg_20_ ( .D(N29), .CK(clk), .RN(rstn), .Q(x1_o1_tmp[20])
         );
  DFFRHQX1 x1_o1_tmp_reg_19_ ( .D(N28), .CK(clk), .RN(rstn), .Q(x1_o1_tmp[19])
         );
  DFFRHQX1 x1_o1_tmp_reg_18_ ( .D(N27), .CK(clk), .RN(rstn), .Q(x1_o1_tmp[18])
         );
  DFFRHQX1 x1_o1_tmp_reg_17_ ( .D(N26), .CK(clk), .RN(rstn), .Q(x1_o1_tmp[17])
         );
  DFFRHQX1 x1_o1_tmp_reg_16_ ( .D(N25), .CK(clk), .RN(rstn), .Q(x1_o1_tmp[16])
         );
  DFFRHQX1 x1_o1_tmp_reg_15_ ( .D(N24), .CK(clk), .RN(rstn), .Q(x1_o1_tmp[15])
         );
  DFFRHQX1 x1_o1_tmp_reg_14_ ( .D(N23), .CK(clk), .RN(rstn), .Q(x1_o1_tmp[14])
         );
  DFFRHQX1 x1_o1_tmp_reg_13_ ( .D(N22), .CK(clk), .RN(rstn), .Q(x1_o1_tmp[13])
         );
  DFFRHQX1 x1_o1_tmp_reg_12_ ( .D(N21), .CK(clk), .RN(rstn), .Q(x1_o1_tmp[12])
         );
  DFFRHQX1 x1_o1_tmp_reg_11_ ( .D(N20), .CK(clk), .RN(rstn), .Q(x1_o1_tmp[11])
         );
  DFFRHQX1 x1_o1_tmp_reg_10_ ( .D(N19), .CK(clk), .RN(rstn), .Q(x1_o1_tmp[10])
         );
  DFFRHQX1 x1_o1_tmp_reg_9_ ( .D(N18), .CK(clk), .RN(rstn), .Q(x1_o1_tmp[9])
         );
  DFFRHQX1 x1_o1_tmp_reg_8_ ( .D(N17), .CK(clk), .RN(rstn), .Q(x1_o1_tmp[8])
         );
  DFFRHQX1 x1_o1_tmp_reg_7_ ( .D(N16), .CK(clk), .RN(rstn), .Q(x1_o1_tmp[7])
         );
  DFFRHQX1 x1_o1_tmp_reg_6_ ( .D(N15), .CK(clk), .RN(rstn), .Q(x1_o1_tmp[6])
         );
  DFFRHQX1 x1_o1_tmp_reg_5_ ( .D(N14), .CK(clk), .RN(rstn), .Q(x1_o1_tmp[5])
         );
  DFFRHQX1 x3_o0_tmp_reg_21_ ( .D(N52), .CK(clk), .RN(rstn), .Q(x3_o0_tmp[21])
         );
  DFFRHQX1 x3_o0_tmp_reg_20_ ( .D(N51), .CK(clk), .RN(rstn), .Q(x3_o0_tmp[20])
         );
  DFFRHQX1 x3_o0_tmp_reg_19_ ( .D(N50), .CK(clk), .RN(rstn), .Q(x3_o0_tmp[19])
         );
  DFFRHQX1 x3_o0_tmp_reg_18_ ( .D(N49), .CK(clk), .RN(rstn), .Q(x3_o0_tmp[18])
         );
  DFFRHQX1 x3_o0_tmp_reg_17_ ( .D(N48), .CK(clk), .RN(rstn), .Q(x3_o0_tmp[17])
         );
  DFFRHQX1 x3_o0_tmp_reg_16_ ( .D(N47), .CK(clk), .RN(rstn), .Q(x3_o0_tmp[16])
         );
  DFFRHQX1 x3_o0_tmp_reg_15_ ( .D(N46), .CK(clk), .RN(rstn), .Q(x3_o0_tmp[15])
         );
  DFFRHQX1 x3_o0_tmp_reg_14_ ( .D(N45), .CK(clk), .RN(rstn), .Q(x3_o0_tmp[14])
         );
  DFFRHQX1 x3_o0_tmp_reg_13_ ( .D(N44), .CK(clk), .RN(rstn), .Q(x3_o0_tmp[13])
         );
  DFFRHQX1 x3_o0_tmp_reg_12_ ( .D(N43), .CK(clk), .RN(rstn), .Q(x3_o0_tmp[12])
         );
  DFFRHQX1 x3_o0_tmp_reg_11_ ( .D(N42), .CK(clk), .RN(rstn), .Q(x3_o0_tmp[11])
         );
  DFFRHQX1 x3_o0_tmp_reg_10_ ( .D(N41), .CK(clk), .RN(rstn), .Q(x3_o0_tmp[10])
         );
  DFFRHQX1 x3_o0_tmp_reg_9_ ( .D(N40), .CK(clk), .RN(rstn), .Q(x3_o0_tmp[9])
         );
  DFFRHQX1 x3_o0_tmp_reg_8_ ( .D(N39), .CK(clk), .RN(rstn), .Q(x3_o0_tmp[8])
         );
  DFFRHQX1 x3_o0_tmp_reg_7_ ( .D(N38), .CK(clk), .RN(rstn), .Q(x3_o0_tmp[7])
         );
  DFFRHQX1 x3_o0_tmp_reg_6_ ( .D(N37), .CK(clk), .RN(rstn), .Q(x3_o0_tmp[6])
         );
  DFFRHQX1 x3_o0_tmp_reg_5_ ( .D(N36), .CK(clk), .RN(rstn), .Q(x3_o0_tmp[5])
         );
  DFFRHQX1 mode_delay1_reg_1_ ( .D(mode[1]), .CK(clk), .RN(rstn), .Q(
        mode_delay1[1]) );
  DFFRHQX1 mode_delay1_reg_0_ ( .D(mode[0]), .CK(clk), .RN(rstn), .Q(
        mode_delay1[0]) );
  DFFRHQX1 idct4_ready_delay3_reg ( .D(idct4_ready_delay2), .CK(clk), .RN(rstn), .Q(idct4_ready_delay3) );
  DFFRHQX1 x1_o1_tmp_reg_4_ ( .D(x1[2]), .CK(clk), .RN(rstn), .Q(x1_o1_tmp[4])
         );
  DFFRHQX1 x1_o1_tmp_reg_3_ ( .D(x1[1]), .CK(clk), .RN(rstn), .Q(x1_o1_tmp[3])
         );
  DFFRHQX1 x1_o1_tmp_reg_2_ ( .D(x1[0]), .CK(clk), .RN(rstn), .Q(x1_o1_tmp[2])
         );
  DFFRHQX1 x2_e_tmp_reg_21_ ( .D(x2[15]), .CK(clk), .RN(rstn), .Q(x2_e_tmp[21]) );
  DFFRHQX1 x2_e_tmp_reg_20_ ( .D(x2[14]), .CK(clk), .RN(rstn), .Q(x2_e_tmp[20]) );
  DFFRHQX1 x2_e_tmp_reg_19_ ( .D(x2[13]), .CK(clk), .RN(rstn), .Q(x2_e_tmp[19]) );
  DFFRHQX1 x2_e_tmp_reg_18_ ( .D(x2[12]), .CK(clk), .RN(rstn), .Q(x2_e_tmp[18]) );
  DFFRHQX1 x2_e_tmp_reg_17_ ( .D(x2[11]), .CK(clk), .RN(rstn), .Q(x2_e_tmp[17]) );
  DFFRHQX1 x2_e_tmp_reg_16_ ( .D(x2[10]), .CK(clk), .RN(rstn), .Q(x2_e_tmp[16]) );
  DFFRHQX1 x2_e_tmp_reg_15_ ( .D(x2[9]), .CK(clk), .RN(rstn), .Q(x2_e_tmp[15])
         );
  DFFRHQX1 x2_e_tmp_reg_14_ ( .D(x2[8]), .CK(clk), .RN(rstn), .Q(x2_e_tmp[14])
         );
  DFFRHQX1 x2_e_tmp_reg_13_ ( .D(x2[7]), .CK(clk), .RN(rstn), .Q(x2_e_tmp[13])
         );
  DFFRHQX1 x2_e_tmp_reg_12_ ( .D(x2[6]), .CK(clk), .RN(rstn), .Q(x2_e_tmp[12])
         );
  DFFRHQX1 x2_e_tmp_reg_11_ ( .D(x2[5]), .CK(clk), .RN(rstn), .Q(x2_e_tmp[11])
         );
  DFFRHQX1 x2_e_tmp_reg_10_ ( .D(x2[4]), .CK(clk), .RN(rstn), .Q(x2_e_tmp[10])
         );
  DFFRHQX1 x2_e_tmp_reg_9_ ( .D(x2[3]), .CK(clk), .RN(rstn), .Q(x2_e_tmp[9])
         );
  DFFRHQX1 x2_e_tmp_reg_8_ ( .D(x2[2]), .CK(clk), .RN(rstn), .Q(x2_e_tmp[8])
         );
  DFFRHQX1 x2_e_tmp_reg_7_ ( .D(x2[1]), .CK(clk), .RN(rstn), .Q(x2_e_tmp[7])
         );
  DFFRHQX1 x2_e_tmp_reg_6_ ( .D(x2[0]), .CK(clk), .RN(rstn), .Q(x2_e_tmp[6])
         );
  DFFRHQX1 x0_e_tmp_reg_21_ ( .D(x0[15]), .CK(clk), .RN(rstn), .Q(x0_e_tmp[21]) );
  DFFRHQX1 x0_e_tmp_reg_20_ ( .D(x0[14]), .CK(clk), .RN(rstn), .Q(x0_e_tmp[20]) );
  DFFRHQX1 x0_e_tmp_reg_19_ ( .D(x0[13]), .CK(clk), .RN(rstn), .Q(x0_e_tmp[19]) );
  DFFRHQX1 x0_e_tmp_reg_18_ ( .D(x0[12]), .CK(clk), .RN(rstn), .Q(x0_e_tmp[18]) );
  DFFRHQX1 x0_e_tmp_reg_17_ ( .D(x0[11]), .CK(clk), .RN(rstn), .Q(x0_e_tmp[17]) );
  DFFRHQX1 x0_e_tmp_reg_16_ ( .D(x0[10]), .CK(clk), .RN(rstn), .Q(x0_e_tmp[16]) );
  DFFRHQX1 x0_e_tmp_reg_15_ ( .D(x0[9]), .CK(clk), .RN(rstn), .Q(x0_e_tmp[15])
         );
  DFFRHQX1 x0_e_tmp_reg_14_ ( .D(x0[8]), .CK(clk), .RN(rstn), .Q(x0_e_tmp[14])
         );
  DFFRHQX1 x0_e_tmp_reg_13_ ( .D(x0[7]), .CK(clk), .RN(rstn), .Q(x0_e_tmp[13])
         );
  DFFRHQX1 x0_e_tmp_reg_12_ ( .D(x0[6]), .CK(clk), .RN(rstn), .Q(x0_e_tmp[12])
         );
  DFFRHQX1 x0_e_tmp_reg_11_ ( .D(x0[5]), .CK(clk), .RN(rstn), .Q(x0_e_tmp[11])
         );
  DFFRHQX1 x0_e_tmp_reg_10_ ( .D(x0[4]), .CK(clk), .RN(rstn), .Q(x0_e_tmp[10])
         );
  DFFRHQX1 x0_e_tmp_reg_9_ ( .D(x0[3]), .CK(clk), .RN(rstn), .Q(x0_e_tmp[9])
         );
  DFFRHQX1 x0_e_tmp_reg_8_ ( .D(x0[2]), .CK(clk), .RN(rstn), .Q(x0_e_tmp[8])
         );
  DFFRHQX1 x0_e_tmp_reg_7_ ( .D(x0[1]), .CK(clk), .RN(rstn), .Q(x0_e_tmp[7])
         );
  DFFRHQX1 x0_e_tmp_reg_6_ ( .D(x0[0]), .CK(clk), .RN(rstn), .Q(x0_e_tmp[6])
         );
  DFFRHQX1 x3_o0_tmp_reg_4_ ( .D(x3[2]), .CK(clk), .RN(rstn), .Q(x3_o0_tmp[4])
         );
  DFFRHQX1 x3_o0_tmp_reg_3_ ( .D(x3[1]), .CK(clk), .RN(rstn), .Q(x3_o0_tmp[3])
         );
  DFFRHQX1 x3_o0_tmp_reg_2_ ( .D(x3[0]), .CK(clk), .RN(rstn), .Q(x3_o0_tmp[2])
         );
  DFFRHQX1 idct4_ready_delay1_reg ( .D(start), .CK(clk), .RN(rstn), .Q(
        idct4_ready_delay1) );
  DFFRHQX1 idct4_ready_delay2_reg ( .D(idct4_ready_delay1), .CK(clk), .RN(rstn), .Q(idct4_ready_delay2) );
  INVX1 U3 ( .A(n36), .Y(n3) );
  INVX1 U4 ( .A(n37), .Y(n4) );
  INVX1 U5 ( .A(n35), .Y(n2) );
  INVX1 U6 ( .A(n37), .Y(n12) );
  INVX1 U7 ( .A(n37), .Y(n11) );
  INVX1 U8 ( .A(n37), .Y(n8) );
  INVX1 U9 ( .A(n38), .Y(n37) );
  INVX1 U10 ( .A(n38), .Y(n36) );
  INVX1 U11 ( .A(n39), .Y(n35) );
  INVX1 U15 ( .A(n49), .Y(n15) );
  INVX1 U18 ( .A(n49), .Y(n14) );
  INVX1 U19 ( .A(n47), .Y(n21) );
  INVX1 U20 ( .A(n47), .Y(n20) );
  INVX1 U21 ( .A(n48), .Y(n17) );
  INVX1 U22 ( .A(n44), .Y(n26) );
  INVX1 U23 ( .A(n44), .Y(n25) );
  INVX1 U24 ( .A(n45), .Y(n22) );
  INVX1 U25 ( .A(n41), .Y(n32) );
  INVX1 U26 ( .A(n41), .Y(n31) );
  INVX1 U27 ( .A(n39), .Y(n34) );
  INVX1 U28 ( .A(n40), .Y(n33) );
  INVX1 U29 ( .A(n42), .Y(n28) );
  INVX1 U30 ( .A(n43), .Y(n27) );
  INVX1 U31 ( .A(n49), .Y(n13) );
  INVX1 U32 ( .A(n47), .Y(n19) );
  INVX1 U33 ( .A(n48), .Y(n18) );
  INVX1 U34 ( .A(n44), .Y(n24) );
  INVX1 U35 ( .A(n45), .Y(n23) );
  INVX1 U36 ( .A(n41), .Y(n30) );
  INVX1 U37 ( .A(n42), .Y(n29) );
  INVX1 U38 ( .A(n46), .Y(n16) );
  INVX1 U39 ( .A(n176), .Y(n38) );
  INVX1 U40 ( .A(n176), .Y(n39) );
  INVX1 U41 ( .A(n176), .Y(n49) );
  INVX1 U42 ( .A(n176), .Y(n47) );
  INVX1 U43 ( .A(n176), .Y(n48) );
  INVX1 U44 ( .A(n176), .Y(n44) );
  INVX1 U45 ( .A(n176), .Y(n45) );
  INVX1 U46 ( .A(n176), .Y(n41) );
  INVX1 U47 ( .A(n176), .Y(n40) );
  INVX1 U48 ( .A(n176), .Y(n42) );
  INVX1 U49 ( .A(n176), .Y(n43) );
  INVX1 U50 ( .A(n176), .Y(n46) );
  INVX1 U51 ( .A(n213), .Y(y2[0]) );
  AOI22X1 U52 ( .A0(N609), .A1(n22), .B0(y2_tmp[0]), .B1(n4), .Y(n213) );
  INVX1 U53 ( .A(n194), .Y(y3[0]) );
  AOI22X1 U54 ( .A0(N628), .A1(n17), .B0(y3_tmp[0]), .B1(n3), .Y(n194) );
  INVX1 U55 ( .A(n251), .Y(y0[0]) );
  AOI22X1 U56 ( .A0(N571), .A1(n34), .B0(y0_tmp[0]), .B1(n2), .Y(n251) );
  INVX1 U57 ( .A(n232), .Y(y1[0]) );
  AOI22X1 U58 ( .A0(N590), .A1(n28), .B0(y1_tmp[0]), .B1(n12), .Y(n232) );
  INVX1 U59 ( .A(n185), .Y(y3[1]) );
  AOI22X1 U60 ( .A0(N629), .A1(n15), .B0(y3_tmp[1]), .B1(n2), .Y(n185) );
  INVX1 U61 ( .A(n204), .Y(y2[1]) );
  AOI22X1 U62 ( .A0(N610), .A1(n21), .B0(y2_tmp[1]), .B1(n4), .Y(n204) );
  INVX1 U63 ( .A(n223), .Y(y1[1]) );
  AOI22X1 U64 ( .A0(N591), .A1(n27), .B0(y1_tmp[1]), .B1(n11), .Y(n223) );
  INVX1 U65 ( .A(n242), .Y(y0[1]) );
  AOI22X1 U66 ( .A0(N572), .A1(n33), .B0(y0_tmp[1]), .B1(n12), .Y(n242) );
  OR2X2 U67 ( .A(mode_delay2[0]), .B(mode_delay2[1]), .Y(n1) );
  INVX1 U68 ( .A(n1), .Y(n176) );
  NAND2X1 U69 ( .A(N646), .B(n36), .Y(n184) );
  NAND2X1 U70 ( .A(N627), .B(n35), .Y(n203) );
  NAND2X1 U71 ( .A(N589), .B(n36), .Y(n241) );
  NAND2X1 U72 ( .A(N608), .B(n35), .Y(n222) );
  INVX1 U73 ( .A(n192), .Y(y3[11]) );
  AOI22X1 U74 ( .A0(N639), .A1(n16), .B0(y3_tmp[11]), .B1(n3), .Y(n192) );
  INVX1 U75 ( .A(n191), .Y(y3[12]) );
  AOI22X1 U76 ( .A0(N640), .A1(n16), .B0(y3_tmp[12]), .B1(n3), .Y(n191) );
  INVX1 U77 ( .A(n186), .Y(y3[17]) );
  AOI22X1 U78 ( .A0(N645), .A1(n16), .B0(y3_tmp[17]), .B1(n2), .Y(n186) );
  INVX1 U79 ( .A(n211), .Y(y2[11]) );
  AOI22X1 U80 ( .A0(N620), .A1(n16), .B0(y2_tmp[11]), .B1(n4), .Y(n211) );
  INVX1 U81 ( .A(n210), .Y(y2[12]) );
  AOI22X1 U82 ( .A0(N621), .A1(n16), .B0(y2_tmp[12]), .B1(n4), .Y(n210) );
  INVX1 U83 ( .A(n205), .Y(y2[17]) );
  AOI22X1 U84 ( .A0(N626), .A1(n16), .B0(y2_tmp[17]), .B1(n4), .Y(n205) );
  INVX1 U85 ( .A(n230), .Y(y1[11]) );
  AOI22X1 U86 ( .A0(N601), .A1(n16), .B0(y1_tmp[11]), .B1(n11), .Y(n230) );
  INVX1 U87 ( .A(n229), .Y(y1[12]) );
  AOI22X1 U88 ( .A0(N602), .A1(n16), .B0(y1_tmp[12]), .B1(n11), .Y(n229) );
  INVX1 U89 ( .A(n249), .Y(y0[11]) );
  AOI22X1 U90 ( .A0(N582), .A1(n16), .B0(y0_tmp[11]), .B1(n12), .Y(n249) );
  INVX1 U91 ( .A(n248), .Y(y0[12]) );
  AOI22X1 U92 ( .A0(N583), .A1(n16), .B0(y0_tmp[12]), .B1(n12), .Y(n248) );
  INVX1 U93 ( .A(n243), .Y(y0[17]) );
  AOI22X1 U94 ( .A0(N588), .A1(n33), .B0(y0_tmp[17]), .B1(n12), .Y(n243) );
  INVX1 U95 ( .A(n224), .Y(y1[17]) );
  AOI22X1 U96 ( .A0(N607), .A1(n27), .B0(y1_tmp[17]), .B1(n8), .Y(n224) );
  OAI2BB1X1 U97 ( .A0N(y3_tmp[18]), .A1N(n46), .B0(n184), .Y(y3[18]) );
  OAI2BB1X1 U98 ( .A0N(y3_tmp[19]), .A1N(n46), .B0(n184), .Y(y3[19]) );
  OAI2BB1X1 U99 ( .A0N(y3_tmp[20]), .A1N(n46), .B0(n184), .Y(y3[20]) );
  OAI2BB1X1 U100 ( .A0N(y2_tmp[18]), .A1N(n46), .B0(n203), .Y(y2[18]) );
  OAI2BB1X1 U101 ( .A0N(y2_tmp[19]), .A1N(n46), .B0(n203), .Y(y2[19]) );
  OAI2BB1X1 U102 ( .A0N(y2_tmp[20]), .A1N(n46), .B0(n203), .Y(y2[20]) );
  OAI2BB1X1 U103 ( .A0N(y0_tmp[18]), .A1N(n46), .B0(n241), .Y(y0[18]) );
  OAI2BB1X1 U104 ( .A0N(y0_tmp[19]), .A1N(n46), .B0(n241), .Y(y0[19]) );
  OAI2BB1X1 U105 ( .A0N(y0_tmp[20]), .A1N(n46), .B0(n241), .Y(y0[20]) );
  OAI2BB1X1 U106 ( .A0N(y1_tmp[18]), .A1N(n46), .B0(n222), .Y(y1[18]) );
  OAI2BB1X1 U107 ( .A0N(y1_tmp[19]), .A1N(n46), .B0(n222), .Y(y1[19]) );
  OAI2BB1X1 U108 ( .A0N(y1_tmp[20]), .A1N(n46), .B0(n222), .Y(y1[20]) );
  INVX1 U109 ( .A(n183), .Y(y3[2]) );
  AOI22X1 U110 ( .A0(N630), .A1(n15), .B0(y3_tmp[2]), .B1(n2), .Y(n183) );
  INVX1 U111 ( .A(n182), .Y(y3[3]) );
  AOI22X1 U112 ( .A0(N631), .A1(n14), .B0(y3_tmp[3]), .B1(n2), .Y(n182) );
  INVX1 U113 ( .A(n181), .Y(y3[4]) );
  AOI22X1 U114 ( .A0(N632), .A1(n14), .B0(y3_tmp[4]), .B1(n2), .Y(n181) );
  INVX1 U115 ( .A(n180), .Y(y3[5]) );
  AOI22X1 U116 ( .A0(N633), .A1(n13), .B0(y3_tmp[5]), .B1(n2), .Y(n180) );
  INVX1 U117 ( .A(n179), .Y(y3[6]) );
  AOI22X1 U118 ( .A0(N634), .A1(n13), .B0(y3_tmp[6]), .B1(n2), .Y(n179) );
  INVX1 U119 ( .A(n178), .Y(y3[7]) );
  AOI22X1 U120 ( .A0(N635), .A1(n18), .B0(y3_tmp[7]), .B1(n2), .Y(n178) );
  INVX1 U121 ( .A(n177), .Y(y3[8]) );
  AOI22X1 U122 ( .A0(N636), .A1(n29), .B0(y3_tmp[8]), .B1(n2), .Y(n177) );
  INVX1 U123 ( .A(n175), .Y(y3[9]) );
  AOI22X1 U124 ( .A0(N637), .A1(n25), .B0(y3_tmp[9]), .B1(n8), .Y(n175) );
  INVX1 U125 ( .A(n193), .Y(y3[10]) );
  AOI22X1 U126 ( .A0(N638), .A1(n29), .B0(y3_tmp[10]), .B1(n3), .Y(n193) );
  INVX1 U127 ( .A(n190), .Y(y3[13]) );
  AOI22X1 U128 ( .A0(N641), .A1(n16), .B0(y3_tmp[13]), .B1(n3), .Y(n190) );
  INVX1 U129 ( .A(n189), .Y(y3[14]) );
  AOI22X1 U130 ( .A0(N642), .A1(n16), .B0(y3_tmp[14]), .B1(n3), .Y(n189) );
  INVX1 U131 ( .A(n188), .Y(y3[15]) );
  AOI22X1 U132 ( .A0(N643), .A1(n16), .B0(y3_tmp[15]), .B1(n2), .Y(n188) );
  INVX1 U133 ( .A(n202), .Y(y2[2]) );
  AOI22X1 U134 ( .A0(N611), .A1(n21), .B0(y2_tmp[2]), .B1(n4), .Y(n202) );
  INVX1 U135 ( .A(n201), .Y(y2[3]) );
  AOI22X1 U136 ( .A0(N612), .A1(n20), .B0(y2_tmp[3]), .B1(n4), .Y(n201) );
  INVX1 U137 ( .A(n200), .Y(y2[4]) );
  AOI22X1 U138 ( .A0(N613), .A1(n20), .B0(y2_tmp[4]), .B1(n3), .Y(n200) );
  INVX1 U139 ( .A(n199), .Y(y2[5]) );
  AOI22X1 U140 ( .A0(N614), .A1(n19), .B0(y2_tmp[5]), .B1(n3), .Y(n199) );
  INVX1 U141 ( .A(n198), .Y(y2[6]) );
  AOI22X1 U142 ( .A0(N615), .A1(n19), .B0(y2_tmp[6]), .B1(n3), .Y(n198) );
  INVX1 U143 ( .A(n197), .Y(y2[7]) );
  AOI22X1 U144 ( .A0(N616), .A1(n18), .B0(y2_tmp[7]), .B1(n3), .Y(n197) );
  INVX1 U145 ( .A(n196), .Y(y2[8]) );
  AOI22X1 U146 ( .A0(N617), .A1(n18), .B0(y2_tmp[8]), .B1(n3), .Y(n196) );
  INVX1 U147 ( .A(n195), .Y(y2[9]) );
  AOI22X1 U148 ( .A0(N618), .A1(n17), .B0(y2_tmp[9]), .B1(n3), .Y(n195) );
  INVX1 U149 ( .A(n212), .Y(y2[10]) );
  AOI22X1 U150 ( .A0(N619), .A1(n29), .B0(y2_tmp[10]), .B1(n4), .Y(n212) );
  INVX1 U151 ( .A(n209), .Y(y2[13]) );
  AOI22X1 U152 ( .A0(N622), .A1(n16), .B0(y2_tmp[13]), .B1(n4), .Y(n209) );
  INVX1 U153 ( .A(n208), .Y(y2[14]) );
  AOI22X1 U154 ( .A0(N623), .A1(n16), .B0(y2_tmp[14]), .B1(n4), .Y(n208) );
  INVX1 U155 ( .A(n207), .Y(y2[15]) );
  AOI22X1 U156 ( .A0(N624), .A1(n16), .B0(y2_tmp[15]), .B1(n4), .Y(n207) );
  INVX1 U157 ( .A(n221), .Y(y1[2]) );
  AOI22X1 U158 ( .A0(N592), .A1(n26), .B0(y1_tmp[2]), .B1(n8), .Y(n221) );
  INVX1 U159 ( .A(n220), .Y(y1[3]) );
  AOI22X1 U160 ( .A0(N593), .A1(n26), .B0(y1_tmp[3]), .B1(n8), .Y(n220) );
  INVX1 U161 ( .A(n219), .Y(y1[4]) );
  AOI22X1 U162 ( .A0(N594), .A1(n25), .B0(y1_tmp[4]), .B1(n8), .Y(n219) );
  INVX1 U163 ( .A(n218), .Y(y1[5]) );
  AOI22X1 U164 ( .A0(N595), .A1(n24), .B0(y1_tmp[5]), .B1(n8), .Y(n218) );
  INVX1 U165 ( .A(n217), .Y(y1[6]) );
  AOI22X1 U166 ( .A0(N596), .A1(n24), .B0(y1_tmp[6]), .B1(n8), .Y(n217) );
  INVX1 U167 ( .A(n216), .Y(y1[7]) );
  AOI22X1 U168 ( .A0(N597), .A1(n23), .B0(y1_tmp[7]), .B1(n8), .Y(n216) );
  INVX1 U169 ( .A(n215), .Y(y1[8]) );
  AOI22X1 U170 ( .A0(N598), .A1(n23), .B0(y1_tmp[8]), .B1(n8), .Y(n215) );
  INVX1 U171 ( .A(n214), .Y(y1[9]) );
  AOI22X1 U172 ( .A0(N599), .A1(n22), .B0(y1_tmp[9]), .B1(n8), .Y(n214) );
  INVX1 U173 ( .A(n231), .Y(y1[10]) );
  AOI22X1 U174 ( .A0(N600), .A1(n28), .B0(y1_tmp[10]), .B1(n11), .Y(n231) );
  INVX1 U175 ( .A(n228), .Y(y1[13]) );
  AOI22X1 U176 ( .A0(N603), .A1(n16), .B0(y1_tmp[13]), .B1(n11), .Y(n228) );
  INVX1 U177 ( .A(n227), .Y(y1[14]) );
  AOI22X1 U178 ( .A0(N604), .A1(n16), .B0(y1_tmp[14]), .B1(n11), .Y(n227) );
  INVX1 U179 ( .A(n226), .Y(y1[15]) );
  AOI22X1 U180 ( .A0(N605), .A1(n16), .B0(y1_tmp[15]), .B1(n8), .Y(n226) );
  INVX1 U181 ( .A(n240), .Y(y0[2]) );
  AOI22X1 U182 ( .A0(N573), .A1(n32), .B0(y0_tmp[2]), .B1(n12), .Y(n240) );
  INVX1 U183 ( .A(n239), .Y(y0[3]) );
  AOI22X1 U184 ( .A0(N574), .A1(n32), .B0(y0_tmp[3]), .B1(n12), .Y(n239) );
  INVX1 U185 ( .A(n238), .Y(y0[4]) );
  AOI22X1 U186 ( .A0(N575), .A1(n31), .B0(y0_tmp[4]), .B1(n8), .Y(n238) );
  INVX1 U187 ( .A(n237), .Y(y0[5]) );
  AOI22X1 U188 ( .A0(N576), .A1(n31), .B0(y0_tmp[5]), .B1(n11), .Y(n237) );
  INVX1 U189 ( .A(n236), .Y(y0[6]) );
  AOI22X1 U190 ( .A0(N577), .A1(n30), .B0(y0_tmp[6]), .B1(n12), .Y(n236) );
  INVX1 U191 ( .A(n235), .Y(y0[7]) );
  AOI22X1 U192 ( .A0(N578), .A1(n30), .B0(y0_tmp[7]), .B1(n11), .Y(n235) );
  INVX1 U193 ( .A(n234), .Y(y0[8]) );
  AOI22X1 U194 ( .A0(N579), .A1(n29), .B0(y0_tmp[8]), .B1(n12), .Y(n234) );
  INVX1 U195 ( .A(n233), .Y(y0[9]) );
  AOI22X1 U196 ( .A0(N580), .A1(n29), .B0(y0_tmp[9]), .B1(n11), .Y(n233) );
  INVX1 U197 ( .A(n250), .Y(y0[10]) );
  AOI22X1 U198 ( .A0(N581), .A1(n34), .B0(y0_tmp[10]), .B1(n11), .Y(n250) );
  INVX1 U199 ( .A(n247), .Y(y0[13]) );
  AOI22X1 U200 ( .A0(N584), .A1(n16), .B0(y0_tmp[13]), .B1(n12), .Y(n247) );
  INVX1 U201 ( .A(n246), .Y(y0[14]) );
  AOI22X1 U202 ( .A0(N585), .A1(n16), .B0(y0_tmp[14]), .B1(n12), .Y(n246) );
  INVX1 U203 ( .A(n245), .Y(y0[15]) );
  AOI22X1 U204 ( .A0(N586), .A1(n16), .B0(y0_tmp[15]), .B1(n11), .Y(n245) );
  INVX1 U205 ( .A(n187), .Y(y3[16]) );
  AOI22X1 U206 ( .A0(N644), .A1(n16), .B0(y3_tmp[16]), .B1(n2), .Y(n187) );
  INVX1 U207 ( .A(n206), .Y(y2[16]) );
  AOI22X1 U208 ( .A0(N625), .A1(n16), .B0(y2_tmp[16]), .B1(n4), .Y(n206) );
  INVX1 U209 ( .A(n244), .Y(y0[16]) );
  AOI22X1 U210 ( .A0(N587), .A1(n16), .B0(y0_tmp[16]), .B1(n12), .Y(n244) );
  INVX1 U211 ( .A(n225), .Y(y1[16]) );
  AOI22X1 U212 ( .A0(N606), .A1(n16), .B0(y1_tmp[16]), .B1(n11), .Y(n225) );
  OAI2BB1X1 U213 ( .A0N(y3_tmp[24]), .A1N(n46), .B0(n184), .Y(y3[24]) );
  OAI2BB1X1 U214 ( .A0N(y2_tmp[24]), .A1N(n46), .B0(n203), .Y(y2[24]) );
  OAI2BB1X1 U215 ( .A0N(y0_tmp[24]), .A1N(n46), .B0(n241), .Y(y0[24]) );
  OAI2BB1X1 U216 ( .A0N(y1_tmp[24]), .A1N(n46), .B0(n222), .Y(y1[24]) );
  OAI2BB1X1 U217 ( .A0N(y3_tmp[21]), .A1N(n46), .B0(n184), .Y(y3[21]) );
  OAI2BB1X1 U218 ( .A0N(y3_tmp[22]), .A1N(n46), .B0(n184), .Y(y3[22]) );
  OAI2BB1X1 U219 ( .A0N(y3_tmp[23]), .A1N(n46), .B0(n184), .Y(y3[23]) );
  OAI2BB1X1 U220 ( .A0N(y2_tmp[21]), .A1N(n46), .B0(n203), .Y(y2[21]) );
  OAI2BB1X1 U221 ( .A0N(y2_tmp[22]), .A1N(n46), .B0(n203), .Y(y2[22]) );
  OAI2BB1X1 U222 ( .A0N(y2_tmp[23]), .A1N(n46), .B0(n203), .Y(y2[23]) );
  OAI2BB1X1 U223 ( .A0N(y0_tmp[21]), .A1N(n46), .B0(n241), .Y(y0[21]) );
  OAI2BB1X1 U224 ( .A0N(y0_tmp[22]), .A1N(n46), .B0(n241), .Y(y0[22]) );
  OAI2BB1X1 U225 ( .A0N(y0_tmp[23]), .A1N(n46), .B0(n241), .Y(y0[23]) );
  OAI2BB1X1 U226 ( .A0N(y1_tmp[21]), .A1N(n46), .B0(n222), .Y(y1[21]) );
  OAI2BB1X1 U227 ( .A0N(y1_tmp[22]), .A1N(n46), .B0(n222), .Y(y1[22]) );
  OAI2BB1X1 U228 ( .A0N(y1_tmp[23]), .A1N(n46), .B0(n222), .Y(y1[23]) );
  INVX1 U229 ( .A(o0[0]), .Y(n120) );
  INVX1 U230 ( .A(o1[0]), .Y(n96) );
  INVX1 U231 ( .A(x3_o1[0]), .Y(n72) );
  INVX1 U232 ( .A(o0[1]), .Y(n119) );
  INVX1 U233 ( .A(o1[1]), .Y(n95) );
  INVX1 U234 ( .A(o0[22]), .Y(n98) );
  INVX1 U235 ( .A(o0[21]), .Y(n99) );
  INVX1 U236 ( .A(o0[20]), .Y(n100) );
  INVX1 U237 ( .A(o0[19]), .Y(n101) );
  INVX1 U238 ( .A(o0[18]), .Y(n102) );
  INVX1 U239 ( .A(o0[17]), .Y(n103) );
  INVX1 U240 ( .A(o0[16]), .Y(n104) );
  INVX1 U241 ( .A(o0[15]), .Y(n105) );
  INVX1 U242 ( .A(o0[14]), .Y(n106) );
  INVX1 U243 ( .A(o0[13]), .Y(n107) );
  INVX1 U244 ( .A(o0[12]), .Y(n108) );
  INVX1 U245 ( .A(o0[11]), .Y(n109) );
  INVX1 U246 ( .A(o0[10]), .Y(n110) );
  INVX1 U247 ( .A(o0[9]), .Y(n111) );
  INVX1 U248 ( .A(o0[8]), .Y(n112) );
  INVX1 U249 ( .A(o0[7]), .Y(n113) );
  INVX1 U250 ( .A(o0[6]), .Y(n114) );
  INVX1 U251 ( .A(o0[5]), .Y(n115) );
  INVX1 U252 ( .A(o0[4]), .Y(n116) );
  INVX1 U253 ( .A(o0[3]), .Y(n117) );
  INVX1 U254 ( .A(o0[2]), .Y(n118) );
  INVX1 U255 ( .A(o1[2]), .Y(n94) );
  INVX1 U256 ( .A(o1[3]), .Y(n93) );
  INVX1 U257 ( .A(o1[4]), .Y(n92) );
  INVX1 U258 ( .A(o1[5]), .Y(n91) );
  INVX1 U259 ( .A(o1[6]), .Y(n90) );
  INVX1 U260 ( .A(o1[7]), .Y(n89) );
  INVX1 U261 ( .A(o1[8]), .Y(n88) );
  INVX1 U262 ( .A(o1[9]), .Y(n87) );
  INVX1 U263 ( .A(o1[10]), .Y(n86) );
  INVX1 U264 ( .A(o1[11]), .Y(n85) );
  INVX1 U265 ( .A(o1[12]), .Y(n84) );
  INVX1 U266 ( .A(o1[13]), .Y(n83) );
  INVX1 U267 ( .A(o1[14]), .Y(n82) );
  INVX1 U268 ( .A(o1[15]), .Y(n81) );
  INVX1 U269 ( .A(o1[16]), .Y(n80) );
  INVX1 U270 ( .A(o1[17]), .Y(n79) );
  INVX1 U271 ( .A(o1[18]), .Y(n78) );
  INVX1 U272 ( .A(o1[19]), .Y(n77) );
  INVX1 U273 ( .A(o1[20]), .Y(n76) );
  INVX1 U274 ( .A(o1[21]), .Y(n75) );
  INVX1 U275 ( .A(o1[22]), .Y(n74) );
  INVX1 U276 ( .A(x3_o1[2]), .Y(n70) );
  INVX1 U277 ( .A(x3_o1[3]), .Y(n69) );
  INVX1 U278 ( .A(x3_o1[4]), .Y(n68) );
  INVX1 U279 ( .A(x3_o1[5]), .Y(n67) );
  INVX1 U280 ( .A(x3_o1[6]), .Y(n66) );
  INVX1 U281 ( .A(x3_o1[7]), .Y(n65) );
  INVX1 U282 ( .A(x3_o1[8]), .Y(n64) );
  INVX1 U283 ( .A(x3_o1[9]), .Y(n63) );
  INVX1 U284 ( .A(x3_o1[10]), .Y(n62) );
  INVX1 U285 ( .A(x3_o1[11]), .Y(n61) );
  INVX1 U286 ( .A(x3_o1[12]), .Y(n60) );
  INVX1 U287 ( .A(x3_o1[13]), .Y(n59) );
  INVX1 U288 ( .A(x3_o1[14]), .Y(n58) );
  INVX1 U289 ( .A(x3_o1[15]), .Y(n57) );
  INVX1 U290 ( .A(x3_o1[16]), .Y(n56) );
  INVX1 U291 ( .A(x3_o1[17]), .Y(n55) );
  INVX1 U292 ( .A(x3_o1[18]), .Y(n54) );
  INVX1 U293 ( .A(x3_o1[19]), .Y(n53) );
  INVX1 U294 ( .A(x3_o1[20]), .Y(n52) );
  INVX1 U295 ( .A(x3_o1[21]), .Y(n51) );
  INVX1 U296 ( .A(x3_o1[1]), .Y(n71) );
  ADDFX2 U297 ( .A(x1[1]), .B(x1[7]), .CI(add_85_carry_7_), .CO(
        add_85_carry_8_), .S(N60) );
  ADDFX2 U298 ( .A(x3[1]), .B(x3[7]), .CI(add_87_carry_7_), .CO(
        add_87_carry_8_), .S(N104) );
  ADDFX2 U299 ( .A(x3[1]), .B(x3[4]), .CI(add_81_carry_6_), .CO(
        add_81_carry_7_), .S(N37) );
  ADDFX2 U300 ( .A(x1[1]), .B(x1[4]), .CI(add_80_carry_6_), .CO(
        add_80_carry_7_), .S(N15) );
  ADDFX2 U301 ( .A(x1[1]), .B(x1[4]), .CI(add_86_carry_5_), .CO(
        add_86_carry_6_), .S(N81) );
  ADDFX2 U302 ( .A(x3[1]), .B(x3[4]), .CI(add_88_carry_5_), .CO(
        add_88_carry_6_), .S(N125) );
  ADDFX2 U303 ( .A(x0_e[7]), .B(add_1_root_add_112_2_B_7_), .CI(
        add_1_root_add_112_2_carry[7]), .CO(add_1_root_add_112_2_carry[8]), 
        .S(N262) );
  INVX1 U304 ( .A(x2_e[7]), .Y(add_1_root_add_112_2_B_7_) );
  ADDFX2 U305 ( .A(x0_e[7]), .B(x2_e[7]), .CI(add_111_carry[7]), .CO(
        add_111_carry[8]), .S(N194) );
  ADDFX2 U306 ( .A(x0_e[8]), .B(x2_e[8]), .CI(add_111_carry[8]), .CO(
        add_111_carry[9]), .S(N195) );
  ADDFX2 U307 ( .A(x0_e[9]), .B(x2_e[9]), .CI(add_111_carry[9]), .CO(
        add_111_carry[10]), .S(N196) );
  ADDFX2 U308 ( .A(x0_e[10]), .B(x2_e[10]), .CI(add_111_carry[10]), .CO(
        add_111_carry[11]), .S(N197) );
  ADDFX2 U309 ( .A(x0_e[11]), .B(x2_e[11]), .CI(add_111_carry[11]), .CO(
        add_111_carry[12]), .S(N198) );
  ADDFX2 U310 ( .A(x0_e[12]), .B(x2_e[12]), .CI(add_111_carry[12]), .CO(
        add_111_carry[13]), .S(N199) );
  ADDFX2 U311 ( .A(x0_e[13]), .B(x2_e[13]), .CI(add_111_carry[13]), .CO(
        add_111_carry[14]), .S(N200) );
  ADDFX2 U312 ( .A(x0_e[14]), .B(x2_e[14]), .CI(add_111_carry[14]), .CO(
        add_111_carry[15]), .S(N201) );
  ADDFX2 U313 ( .A(x0_e[15]), .B(x2_e[15]), .CI(add_111_carry[15]), .CO(
        add_111_carry[16]), .S(N202) );
  ADDFX2 U314 ( .A(x0_e[16]), .B(x2_e[16]), .CI(add_111_carry[16]), .CO(
        add_111_carry[17]), .S(N203) );
  ADDFX2 U315 ( .A(x0_e[17]), .B(x2_e[17]), .CI(add_111_carry[17]), .CO(
        add_111_carry[18]), .S(N204) );
  ADDFX2 U316 ( .A(x0_e[18]), .B(x2_e[18]), .CI(add_111_carry[18]), .CO(
        add_111_carry[19]), .S(N205) );
  ADDFX2 U317 ( .A(x0_e[19]), .B(x2_e[19]), .CI(add_111_carry[19]), .CO(
        add_111_carry[20]), .S(N206) );
  ADDFX2 U318 ( .A(x0_e[20]), .B(x2_e[20]), .CI(add_111_carry[20]), .CO(
        add_111_carry[21]), .S(N207) );
  ADDFX2 U319 ( .A(x0_e[21]), .B(x2_e[21]), .CI(add_111_carry[21]), .CO(
        add_111_carry[22]), .S(N208) );
  ADDFX2 U320 ( .A(x0_e[8]), .B(add_1_root_add_112_2_B_8_), .CI(
        add_1_root_add_112_2_carry[8]), .CO(add_1_root_add_112_2_carry[9]), 
        .S(N263) );
  INVX1 U321 ( .A(x2_e[8]), .Y(add_1_root_add_112_2_B_8_) );
  ADDFX2 U322 ( .A(x0_e[9]), .B(add_1_root_add_112_2_B_9_), .CI(
        add_1_root_add_112_2_carry[9]), .CO(add_1_root_add_112_2_carry[10]), 
        .S(N264) );
  INVX1 U323 ( .A(x2_e[9]), .Y(add_1_root_add_112_2_B_9_) );
  ADDFX2 U324 ( .A(x0_e[10]), .B(add_1_root_add_112_2_B_10_), .CI(
        add_1_root_add_112_2_carry[10]), .CO(add_1_root_add_112_2_carry[11]), 
        .S(N265) );
  INVX1 U325 ( .A(x2_e[10]), .Y(add_1_root_add_112_2_B_10_) );
  ADDFX2 U326 ( .A(x0_e[11]), .B(add_1_root_add_112_2_B_11_), .CI(
        add_1_root_add_112_2_carry[11]), .CO(add_1_root_add_112_2_carry[12]), 
        .S(N266) );
  INVX1 U327 ( .A(x2_e[11]), .Y(add_1_root_add_112_2_B_11_) );
  ADDFX2 U328 ( .A(x0_e[12]), .B(add_1_root_add_112_2_B_12_), .CI(
        add_1_root_add_112_2_carry[12]), .CO(add_1_root_add_112_2_carry[13]), 
        .S(N267) );
  INVX1 U329 ( .A(x2_e[12]), .Y(add_1_root_add_112_2_B_12_) );
  ADDFX2 U330 ( .A(x0_e[13]), .B(add_1_root_add_112_2_B_13_), .CI(
        add_1_root_add_112_2_carry[13]), .CO(add_1_root_add_112_2_carry[14]), 
        .S(N268) );
  INVX1 U331 ( .A(x2_e[13]), .Y(add_1_root_add_112_2_B_13_) );
  ADDFX2 U332 ( .A(x0_e[14]), .B(add_1_root_add_112_2_B_14_), .CI(
        add_1_root_add_112_2_carry[14]), .CO(add_1_root_add_112_2_carry[15]), 
        .S(N269) );
  INVX1 U333 ( .A(x2_e[14]), .Y(add_1_root_add_112_2_B_14_) );
  ADDFX2 U334 ( .A(x0_e[15]), .B(add_1_root_add_112_2_B_15_), .CI(
        add_1_root_add_112_2_carry[15]), .CO(add_1_root_add_112_2_carry[16]), 
        .S(N270) );
  INVX1 U335 ( .A(x2_e[15]), .Y(add_1_root_add_112_2_B_15_) );
  ADDFX2 U336 ( .A(x0_e[16]), .B(add_1_root_add_112_2_B_16_), .CI(
        add_1_root_add_112_2_carry[16]), .CO(add_1_root_add_112_2_carry[17]), 
        .S(N271) );
  INVX1 U337 ( .A(x2_e[16]), .Y(add_1_root_add_112_2_B_16_) );
  ADDFX2 U338 ( .A(x0_e[17]), .B(add_1_root_add_112_2_B_17_), .CI(
        add_1_root_add_112_2_carry[17]), .CO(add_1_root_add_112_2_carry[18]), 
        .S(N272) );
  INVX1 U339 ( .A(x2_e[17]), .Y(add_1_root_add_112_2_B_17_) );
  ADDFX2 U340 ( .A(x0_e[18]), .B(add_1_root_add_112_2_B_18_), .CI(
        add_1_root_add_112_2_carry[18]), .CO(add_1_root_add_112_2_carry[19]), 
        .S(N273) );
  INVX1 U341 ( .A(x2_e[18]), .Y(add_1_root_add_112_2_B_18_) );
  ADDFX2 U342 ( .A(x0_e[19]), .B(add_1_root_add_112_2_B_19_), .CI(
        add_1_root_add_112_2_carry[19]), .CO(add_1_root_add_112_2_carry[20]), 
        .S(N274) );
  INVX1 U343 ( .A(x2_e[19]), .Y(add_1_root_add_112_2_B_19_) );
  ADDFX2 U344 ( .A(x0_e[20]), .B(add_1_root_add_112_2_B_20_), .CI(
        add_1_root_add_112_2_carry[20]), .CO(add_1_root_add_112_2_carry[21]), 
        .S(N275) );
  INVX1 U345 ( .A(x2_e[20]), .Y(add_1_root_add_112_2_B_20_) );
  ADDFX2 U346 ( .A(x0_e[21]), .B(add_1_root_add_112_2_B_21_), .CI(
        add_1_root_add_112_2_carry[21]), .CO(add_1_root_add_112_2_carry[22]), 
        .S(N276) );
  ADDFX2 U347 ( .A(x1[2]), .B(x1[8]), .CI(add_85_carry_8_), .CO(
        add_85_carry_9_), .S(N61) );
  ADDFX2 U348 ( .A(x1[3]), .B(x1[9]), .CI(add_85_carry_9_), .CO(
        add_85_carry_10_), .S(N62) );
  ADDFX2 U349 ( .A(x1[4]), .B(x1[10]), .CI(add_85_carry_10_), .CO(
        add_85_carry_11_), .S(N63) );
  ADDFX2 U350 ( .A(x1[5]), .B(x1[11]), .CI(add_85_carry_11_), .CO(
        add_85_carry_12_), .S(N64) );
  ADDFX2 U351 ( .A(x1[6]), .B(x1[12]), .CI(add_85_carry_12_), .CO(
        add_85_carry_13_), .S(N65) );
  ADDFX2 U352 ( .A(x1[7]), .B(x1[13]), .CI(add_85_carry_13_), .CO(
        add_85_carry_14_), .S(N66) );
  ADDFX2 U353 ( .A(x1[8]), .B(x1[14]), .CI(add_85_carry_14_), .CO(
        add_85_carry_15_), .S(N67) );
  ADDFX2 U354 ( .A(x1[9]), .B(N30), .CI(add_85_carry_15_), .CO(
        add_85_carry_16_), .S(N68) );
  ADDFX2 U355 ( .A(x1[10]), .B(N30), .CI(add_85_carry_16_), .CO(
        add_85_carry_17_), .S(N69) );
  ADDFX2 U356 ( .A(x1[11]), .B(N30), .CI(add_85_carry_17_), .CO(
        add_85_carry_18_), .S(N70) );
  ADDFX2 U357 ( .A(x1[12]), .B(N30), .CI(add_85_carry_18_), .CO(
        add_85_carry_19_), .S(N71) );
  ADDFX2 U358 ( .A(x1[13]), .B(N30), .CI(add_85_carry_19_), .CO(
        add_85_carry_20_), .S(N72) );
  ADDFX2 U359 ( .A(x3[2]), .B(x3[5]), .CI(add_81_carry_7_), .CO(
        add_81_carry_8_), .S(N38) );
  ADDFX2 U360 ( .A(x3[3]), .B(x3[6]), .CI(add_81_carry_8_), .CO(
        add_81_carry_9_), .S(N39) );
  ADDFX2 U361 ( .A(x3[4]), .B(x3[7]), .CI(add_81_carry_9_), .CO(
        add_81_carry_10_), .S(N40) );
  ADDFX2 U362 ( .A(x3[5]), .B(x3[8]), .CI(add_81_carry_10_), .CO(
        add_81_carry_11_), .S(N41) );
  ADDFX2 U363 ( .A(x3[6]), .B(x3[9]), .CI(add_81_carry_11_), .CO(
        add_81_carry_12_), .S(N42) );
  ADDFX2 U364 ( .A(x3[7]), .B(x3[10]), .CI(add_81_carry_12_), .CO(
        add_81_carry_13_), .S(N43) );
  ADDFX2 U365 ( .A(x3[8]), .B(x3[11]), .CI(add_81_carry_13_), .CO(
        add_81_carry_14_), .S(N44) );
  ADDFX2 U366 ( .A(x3[9]), .B(x3[12]), .CI(add_81_carry_14_), .CO(
        add_81_carry_15_), .S(N45) );
  ADDFX2 U367 ( .A(x3[10]), .B(x3[13]), .CI(add_81_carry_15_), .CO(
        add_81_carry_16_), .S(N46) );
  ADDFX2 U368 ( .A(x3[11]), .B(x3[14]), .CI(add_81_carry_16_), .CO(
        add_81_carry_17_), .S(N47) );
  ADDFX2 U369 ( .A(x3[12]), .B(N52), .CI(add_81_carry_17_), .CO(
        add_81_carry_18_), .S(N48) );
  ADDFX2 U370 ( .A(x3[13]), .B(N52), .CI(add_81_carry_18_), .CO(
        add_81_carry_19_), .S(N49) );
  ADDFX2 U371 ( .A(x1[2]), .B(x1[5]), .CI(add_80_carry_7_), .CO(
        add_80_carry_8_), .S(N16) );
  ADDFX2 U372 ( .A(x1[3]), .B(x1[6]), .CI(add_80_carry_8_), .CO(
        add_80_carry_9_), .S(N17) );
  ADDFX2 U373 ( .A(x1[4]), .B(x1[7]), .CI(add_80_carry_9_), .CO(
        add_80_carry_10_), .S(N18) );
  ADDFX2 U374 ( .A(x1[5]), .B(x1[8]), .CI(add_80_carry_10_), .CO(
        add_80_carry_11_), .S(N19) );
  ADDFX2 U375 ( .A(x1[6]), .B(x1[9]), .CI(add_80_carry_11_), .CO(
        add_80_carry_12_), .S(N20) );
  ADDFX2 U376 ( .A(x1[7]), .B(x1[10]), .CI(add_80_carry_12_), .CO(
        add_80_carry_13_), .S(N21) );
  ADDFX2 U377 ( .A(x1[8]), .B(x1[11]), .CI(add_80_carry_13_), .CO(
        add_80_carry_14_), .S(N22) );
  ADDFX2 U378 ( .A(x1[9]), .B(x1[12]), .CI(add_80_carry_14_), .CO(
        add_80_carry_15_), .S(N23) );
  ADDFX2 U379 ( .A(x1[10]), .B(x1[13]), .CI(add_80_carry_15_), .CO(
        add_80_carry_16_), .S(N24) );
  ADDFX2 U380 ( .A(x1[11]), .B(x1[14]), .CI(add_80_carry_16_), .CO(
        add_80_carry_17_), .S(N25) );
  ADDFX2 U381 ( .A(x1[12]), .B(N30), .CI(add_80_carry_17_), .CO(
        add_80_carry_18_), .S(N26) );
  ADDFX2 U382 ( .A(x1[13]), .B(N30), .CI(add_80_carry_18_), .CO(
        add_80_carry_19_), .S(N27) );
  ADDFX2 U383 ( .A(x1[2]), .B(x1[5]), .CI(add_86_carry_6_), .CO(
        add_86_carry_7_), .S(N82) );
  ADDFX2 U384 ( .A(x1[3]), .B(x1[6]), .CI(add_86_carry_7_), .CO(
        add_86_carry_8_), .S(N83) );
  ADDFX2 U385 ( .A(x1[4]), .B(x1[7]), .CI(add_86_carry_8_), .CO(
        add_86_carry_9_), .S(N84) );
  ADDFX2 U386 ( .A(x1[5]), .B(x1[8]), .CI(add_86_carry_9_), .CO(
        add_86_carry_10_), .S(N85) );
  ADDFX2 U387 ( .A(x1[6]), .B(x1[9]), .CI(add_86_carry_10_), .CO(
        add_86_carry_11_), .S(N86) );
  ADDFX2 U388 ( .A(x1[7]), .B(x1[10]), .CI(add_86_carry_11_), .CO(
        add_86_carry_12_), .S(N87) );
  ADDFX2 U389 ( .A(x1[8]), .B(x1[11]), .CI(add_86_carry_12_), .CO(
        add_86_carry_13_), .S(N88) );
  ADDFX2 U390 ( .A(x1[9]), .B(x1[12]), .CI(add_86_carry_13_), .CO(
        add_86_carry_14_), .S(N89) );
  ADDFX2 U391 ( .A(x1[10]), .B(x1[13]), .CI(add_86_carry_14_), .CO(
        add_86_carry_15_), .S(N90) );
  ADDFX2 U392 ( .A(x1[11]), .B(x1[14]), .CI(add_86_carry_15_), .CO(
        add_86_carry_16_), .S(N91) );
  ADDFX2 U393 ( .A(x1[12]), .B(N30), .CI(add_86_carry_16_), .CO(
        add_86_carry_17_), .S(N92) );
  ADDFX2 U394 ( .A(x1[13]), .B(N30), .CI(add_86_carry_17_), .CO(
        add_86_carry_18_), .S(N93) );
  ADDFX2 U395 ( .A(x3[2]), .B(x3[8]), .CI(add_87_carry_8_), .CO(
        add_87_carry_9_), .S(N105) );
  ADDFX2 U396 ( .A(x3[3]), .B(x3[9]), .CI(add_87_carry_9_), .CO(
        add_87_carry_10_), .S(N106) );
  ADDFX2 U397 ( .A(x3[4]), .B(x3[10]), .CI(add_87_carry_10_), .CO(
        add_87_carry_11_), .S(N107) );
  ADDFX2 U398 ( .A(x3[5]), .B(x3[11]), .CI(add_87_carry_11_), .CO(
        add_87_carry_12_), .S(N108) );
  ADDFX2 U399 ( .A(x3[6]), .B(x3[12]), .CI(add_87_carry_12_), .CO(
        add_87_carry_13_), .S(N109) );
  ADDFX2 U400 ( .A(x3[7]), .B(x3[13]), .CI(add_87_carry_13_), .CO(
        add_87_carry_14_), .S(N110) );
  ADDFX2 U401 ( .A(x3[8]), .B(x3[14]), .CI(add_87_carry_14_), .CO(
        add_87_carry_15_), .S(N111) );
  ADDFX2 U402 ( .A(x3[9]), .B(N52), .CI(add_87_carry_15_), .CO(
        add_87_carry_16_), .S(N112) );
  ADDFX2 U403 ( .A(x3[10]), .B(N52), .CI(add_87_carry_16_), .CO(
        add_87_carry_17_), .S(N113) );
  ADDFX2 U404 ( .A(x3[11]), .B(N52), .CI(add_87_carry_17_), .CO(
        add_87_carry_18_), .S(N114) );
  ADDFX2 U405 ( .A(x3[12]), .B(N52), .CI(add_87_carry_18_), .CO(
        add_87_carry_19_), .S(N115) );
  ADDFX2 U406 ( .A(x3[13]), .B(N52), .CI(add_87_carry_19_), .CO(
        add_87_carry_20_), .S(N116) );
  ADDFX2 U407 ( .A(x3[2]), .B(x3[5]), .CI(add_88_carry_6_), .CO(
        add_88_carry_7_), .S(N126) );
  ADDFX2 U408 ( .A(x3[3]), .B(x3[6]), .CI(add_88_carry_7_), .CO(
        add_88_carry_8_), .S(N127) );
  ADDFX2 U409 ( .A(x3[4]), .B(x3[7]), .CI(add_88_carry_8_), .CO(
        add_88_carry_9_), .S(N128) );
  ADDFX2 U410 ( .A(x3[5]), .B(x3[8]), .CI(add_88_carry_9_), .CO(
        add_88_carry_10_), .S(N129) );
  ADDFX2 U411 ( .A(x3[6]), .B(x3[9]), .CI(add_88_carry_10_), .CO(
        add_88_carry_11_), .S(N130) );
  ADDFX2 U412 ( .A(x3[7]), .B(x3[10]), .CI(add_88_carry_11_), .CO(
        add_88_carry_12_), .S(N131) );
  ADDFX2 U413 ( .A(x3[8]), .B(x3[11]), .CI(add_88_carry_12_), .CO(
        add_88_carry_13_), .S(N132) );
  ADDFX2 U414 ( .A(x3[9]), .B(x3[12]), .CI(add_88_carry_13_), .CO(
        add_88_carry_14_), .S(N133) );
  ADDFX2 U415 ( .A(x3[10]), .B(x3[13]), .CI(add_88_carry_14_), .CO(
        add_88_carry_15_), .S(N134) );
  ADDFX2 U416 ( .A(x3[11]), .B(x3[14]), .CI(add_88_carry_15_), .CO(
        add_88_carry_16_), .S(N135) );
  ADDFX2 U417 ( .A(x3[12]), .B(N52), .CI(add_88_carry_16_), .CO(
        add_88_carry_17_), .S(N136) );
  ADDFX2 U418 ( .A(x3[13]), .B(N52), .CI(add_88_carry_17_), .CO(
        add_88_carry_18_), .S(N137) );
  XOR3X2 U419 ( .A(x0_e[21]), .B(x2_e[21]), .C(add_111_carry[22]), .Y(N209) );
  XOR3X2 U420 ( .A(x0_e[21]), .B(add_1_root_add_112_2_B_21_), .C(
        add_1_root_add_112_2_carry[22]), .Y(N277) );
  ADDFX2 U421 ( .A(x1[14]), .B(N30), .CI(add_85_carry_20_), .CO(N74), .S(N73)
         );
  ADDFX2 U422 ( .A(x3[14]), .B(N52), .CI(add_81_carry_19_), .CO(N51), .S(N50)
         );
  ADDFX2 U423 ( .A(x1[14]), .B(N30), .CI(add_80_carry_19_), .CO(N29), .S(N28)
         );
  ADDFX2 U424 ( .A(x1[14]), .B(N30), .CI(add_86_carry_18_), .CO(N95), .S(N94)
         );
  ADDFX2 U425 ( .A(x3[14]), .B(N52), .CI(add_87_carry_20_), .CO(N118), .S(N117) );
  ADDFX2 U426 ( .A(x3[14]), .B(N52), .CI(add_88_carry_18_), .CO(N139), .S(N138) );
  INVX1 U427 ( .A(x2_e[6]), .Y(add_1_root_add_112_2_B_6_) );
  BUFX3 U428 ( .A(x1[15]), .Y(N30) );
  BUFX3 U429 ( .A(x3[15]), .Y(N52) );
  INVX1 U430 ( .A(o0[23]), .Y(n97) );
  INVX1 U431 ( .A(o1[23]), .Y(n73) );
  INVX1 U432 ( .A(x2_e[21]), .Y(add_1_root_add_112_2_B_21_) );
  INVX1 U433 ( .A(x3_o1[22]), .Y(n50) );
  XOR2X1 U452 ( .A(y3_tmp[24]), .B(add_125_carry_25_), .Y(N646) );
  AND2X1 U453 ( .A(add_125_carry_24_), .B(y3_tmp[24]), .Y(add_125_carry_25_)
         );
  XOR2X1 U454 ( .A(y3_tmp[24]), .B(add_125_carry_24_), .Y(N645) );
  AND2X1 U455 ( .A(add_125_carry_23_), .B(y3_tmp[23]), .Y(add_125_carry_24_)
         );
  XOR2X1 U456 ( .A(y3_tmp[23]), .B(add_125_carry_23_), .Y(N644) );
  XOR2X1 U457 ( .A(y2_tmp[24]), .B(add_124_carry_25_), .Y(N627) );
  AND2X1 U458 ( .A(add_124_carry_24_), .B(y2_tmp[24]), .Y(add_124_carry_25_)
         );
  XOR2X1 U459 ( .A(y2_tmp[24]), .B(add_124_carry_24_), .Y(N626) );
  AND2X1 U460 ( .A(add_124_carry_23_), .B(y2_tmp[23]), .Y(add_124_carry_24_)
         );
  XOR2X1 U461 ( .A(y2_tmp[23]), .B(add_124_carry_23_), .Y(N625) );
  XOR2X1 U462 ( .A(y0_tmp[24]), .B(add_122_carry_25_), .Y(N589) );
  AND2X1 U463 ( .A(add_122_carry_24_), .B(y0_tmp[24]), .Y(add_122_carry_25_)
         );
  XOR2X1 U464 ( .A(y0_tmp[24]), .B(add_122_carry_24_), .Y(N588) );
  AND2X1 U465 ( .A(add_122_carry_23_), .B(y0_tmp[23]), .Y(add_122_carry_24_)
         );
  XOR2X1 U466 ( .A(y0_tmp[23]), .B(add_122_carry_23_), .Y(N587) );
  XOR2X1 U467 ( .A(y1_tmp[24]), .B(add_123_carry_25_), .Y(N608) );
  AND2X1 U468 ( .A(add_123_carry_24_), .B(y1_tmp[24]), .Y(add_123_carry_25_)
         );
  XOR2X1 U469 ( .A(y1_tmp[24]), .B(add_123_carry_24_), .Y(N607) );
  AND2X1 U470 ( .A(add_123_carry_23_), .B(y1_tmp[23]), .Y(add_123_carry_24_)
         );
  XOR2X1 U471 ( .A(y1_tmp[23]), .B(add_123_carry_23_), .Y(N606) );
  AND2X1 U472 ( .A(x0_e[6]), .B(x2_e[6]), .Y(add_111_carry[7]) );
  XOR2X1 U473 ( .A(x2_e[6]), .B(x0_e[6]), .Y(N193) );
  OR2X1 U474 ( .A(add_1_root_add_112_2_B_6_), .B(x0_e[6]), .Y(
        add_1_root_add_112_2_carry[7]) );
  XNOR2X1 U475 ( .A(x0_e[6]), .B(add_1_root_add_112_2_B_6_), .Y(N261) );
  AND2X1 U476 ( .A(x1[0]), .B(x1[6]), .Y(add_85_carry_7_) );
  XOR2X1 U477 ( .A(x1[6]), .B(x1[0]), .Y(N59) );
  AND2X1 U478 ( .A(x3[0]), .B(x3[3]), .Y(add_81_carry_6_) );
  XOR2X1 U479 ( .A(x3[3]), .B(x3[0]), .Y(N36) );
  AND2X1 U480 ( .A(x1[0]), .B(x1[3]), .Y(add_80_carry_6_) );
  XOR2X1 U481 ( .A(x1[3]), .B(x1[0]), .Y(N14) );
  AND2X1 U482 ( .A(x1[0]), .B(x1[3]), .Y(add_86_carry_5_) );
  XOR2X1 U483 ( .A(x1[3]), .B(x1[0]), .Y(N80) );
  AND2X1 U484 ( .A(x3[0]), .B(x3[6]), .Y(add_87_carry_7_) );
  XOR2X1 U485 ( .A(x3[6]), .B(x3[0]), .Y(N103) );
  AND2X1 U486 ( .A(x3[0]), .B(x3[3]), .Y(add_88_carry_5_) );
  XOR2X1 U487 ( .A(x3[3]), .B(x3[0]), .Y(N124) );
  AND2X1 U488 ( .A(add_122_carry_22_), .B(y0_tmp[22]), .Y(add_122_carry_23_)
         );
  XOR2X1 U489 ( .A(y0_tmp[22]), .B(add_122_carry_22_), .Y(N586) );
  AND2X1 U490 ( .A(add_122_carry_21_), .B(y0_tmp[21]), .Y(add_122_carry_22_)
         );
  XOR2X1 U491 ( .A(y0_tmp[21]), .B(add_122_carry_21_), .Y(N585) );
  AND2X1 U492 ( .A(add_122_carry_20_), .B(y0_tmp[20]), .Y(add_122_carry_21_)
         );
  XOR2X1 U493 ( .A(y0_tmp[20]), .B(add_122_carry_20_), .Y(N584) );
  AND2X1 U494 ( .A(add_122_carry_19_), .B(y0_tmp[19]), .Y(add_122_carry_20_)
         );
  XOR2X1 U495 ( .A(y0_tmp[19]), .B(add_122_carry_19_), .Y(N583) );
  AND2X1 U496 ( .A(add_122_carry_18_), .B(y0_tmp[18]), .Y(add_122_carry_19_)
         );
  XOR2X1 U497 ( .A(y0_tmp[18]), .B(add_122_carry_18_), .Y(N582) );
  AND2X1 U498 ( .A(add_122_carry_17_), .B(y0_tmp[17]), .Y(add_122_carry_18_)
         );
  XOR2X1 U499 ( .A(y0_tmp[17]), .B(add_122_carry_17_), .Y(N581) );
  AND2X1 U500 ( .A(add_122_carry_16_), .B(y0_tmp[16]), .Y(add_122_carry_17_)
         );
  XOR2X1 U501 ( .A(y0_tmp[16]), .B(add_122_carry_16_), .Y(N580) );
  AND2X1 U502 ( .A(add_122_carry_15_), .B(y0_tmp[15]), .Y(add_122_carry_16_)
         );
  XOR2X1 U503 ( .A(y0_tmp[15]), .B(add_122_carry_15_), .Y(N579) );
  AND2X1 U504 ( .A(add_122_carry_14_), .B(y0_tmp[14]), .Y(add_122_carry_15_)
         );
  XOR2X1 U505 ( .A(y0_tmp[14]), .B(add_122_carry_14_), .Y(N578) );
  AND2X1 U506 ( .A(add_122_carry_13_), .B(y0_tmp[13]), .Y(add_122_carry_14_)
         );
  XOR2X1 U507 ( .A(y0_tmp[13]), .B(add_122_carry_13_), .Y(N577) );
  AND2X1 U508 ( .A(add_122_carry_12_), .B(y0_tmp[12]), .Y(add_122_carry_13_)
         );
  XOR2X1 U509 ( .A(y0_tmp[12]), .B(add_122_carry_12_), .Y(N576) );
  AND2X1 U510 ( .A(add_122_carry_11_), .B(y0_tmp[11]), .Y(add_122_carry_12_)
         );
  XOR2X1 U511 ( .A(y0_tmp[11]), .B(add_122_carry_11_), .Y(N575) );
  AND2X1 U512 ( .A(add_122_carry_10_), .B(y0_tmp[10]), .Y(add_122_carry_11_)
         );
  XOR2X1 U513 ( .A(y0_tmp[10]), .B(add_122_carry_10_), .Y(N574) );
  AND2X1 U514 ( .A(add_122_carry_9_), .B(y0_tmp[9]), .Y(add_122_carry_10_) );
  XOR2X1 U515 ( .A(y0_tmp[9]), .B(add_122_carry_9_), .Y(N573) );
  AND2X1 U516 ( .A(add_122_carry_8_), .B(y0_tmp[8]), .Y(add_122_carry_9_) );
  XOR2X1 U517 ( .A(y0_tmp[8]), .B(add_122_carry_8_), .Y(N572) );
  AND2X1 U518 ( .A(y0_tmp[6]), .B(y0_tmp[7]), .Y(add_122_carry_8_) );
  XOR2X1 U519 ( .A(y0_tmp[7]), .B(y0_tmp[6]), .Y(N571) );
  AND2X1 U520 ( .A(add_123_carry_22_), .B(y1_tmp[22]), .Y(add_123_carry_23_)
         );
  XOR2X1 U521 ( .A(y1_tmp[22]), .B(add_123_carry_22_), .Y(N605) );
  AND2X1 U522 ( .A(add_123_carry_21_), .B(y1_tmp[21]), .Y(add_123_carry_22_)
         );
  XOR2X1 U523 ( .A(y1_tmp[21]), .B(add_123_carry_21_), .Y(N604) );
  AND2X1 U524 ( .A(add_123_carry_20_), .B(y1_tmp[20]), .Y(add_123_carry_21_)
         );
  XOR2X1 U525 ( .A(y1_tmp[20]), .B(add_123_carry_20_), .Y(N603) );
  AND2X1 U526 ( .A(add_123_carry_19_), .B(y1_tmp[19]), .Y(add_123_carry_20_)
         );
  XOR2X1 U527 ( .A(y1_tmp[19]), .B(add_123_carry_19_), .Y(N602) );
  AND2X1 U528 ( .A(add_123_carry_18_), .B(y1_tmp[18]), .Y(add_123_carry_19_)
         );
  XOR2X1 U529 ( .A(y1_tmp[18]), .B(add_123_carry_18_), .Y(N601) );
  AND2X1 U530 ( .A(add_123_carry_17_), .B(y1_tmp[17]), .Y(add_123_carry_18_)
         );
  XOR2X1 U531 ( .A(y1_tmp[17]), .B(add_123_carry_17_), .Y(N600) );
  AND2X1 U532 ( .A(add_123_carry_16_), .B(y1_tmp[16]), .Y(add_123_carry_17_)
         );
  XOR2X1 U533 ( .A(y1_tmp[16]), .B(add_123_carry_16_), .Y(N599) );
  AND2X1 U534 ( .A(add_123_carry_15_), .B(y1_tmp[15]), .Y(add_123_carry_16_)
         );
  XOR2X1 U535 ( .A(y1_tmp[15]), .B(add_123_carry_15_), .Y(N598) );
  AND2X1 U536 ( .A(add_123_carry_14_), .B(y1_tmp[14]), .Y(add_123_carry_15_)
         );
  XOR2X1 U537 ( .A(y1_tmp[14]), .B(add_123_carry_14_), .Y(N597) );
  AND2X1 U538 ( .A(add_123_carry_13_), .B(y1_tmp[13]), .Y(add_123_carry_14_)
         );
  XOR2X1 U539 ( .A(y1_tmp[13]), .B(add_123_carry_13_), .Y(N596) );
  AND2X1 U540 ( .A(add_123_carry_12_), .B(y1_tmp[12]), .Y(add_123_carry_13_)
         );
  XOR2X1 U541 ( .A(y1_tmp[12]), .B(add_123_carry_12_), .Y(N595) );
  AND2X1 U542 ( .A(add_123_carry_11_), .B(y1_tmp[11]), .Y(add_123_carry_12_)
         );
  XOR2X1 U543 ( .A(y1_tmp[11]), .B(add_123_carry_11_), .Y(N594) );
  AND2X1 U544 ( .A(add_123_carry_10_), .B(y1_tmp[10]), .Y(add_123_carry_11_)
         );
  XOR2X1 U545 ( .A(y1_tmp[10]), .B(add_123_carry_10_), .Y(N593) );
  AND2X1 U546 ( .A(add_123_carry_9_), .B(y1_tmp[9]), .Y(add_123_carry_10_) );
  XOR2X1 U547 ( .A(y1_tmp[9]), .B(add_123_carry_9_), .Y(N592) );
  AND2X1 U548 ( .A(add_123_carry_8_), .B(y1_tmp[8]), .Y(add_123_carry_9_) );
  XOR2X1 U549 ( .A(y1_tmp[8]), .B(add_123_carry_8_), .Y(N591) );
  AND2X1 U550 ( .A(y1_tmp[6]), .B(y1_tmp[7]), .Y(add_123_carry_8_) );
  XOR2X1 U551 ( .A(y1_tmp[7]), .B(y1_tmp[6]), .Y(N590) );
  AND2X1 U552 ( .A(add_124_carry_22_), .B(y2_tmp[22]), .Y(add_124_carry_23_)
         );
  XOR2X1 U553 ( .A(y2_tmp[22]), .B(add_124_carry_22_), .Y(N624) );
  AND2X1 U554 ( .A(add_124_carry_21_), .B(y2_tmp[21]), .Y(add_124_carry_22_)
         );
  XOR2X1 U555 ( .A(y2_tmp[21]), .B(add_124_carry_21_), .Y(N623) );
  AND2X1 U556 ( .A(add_124_carry_20_), .B(y2_tmp[20]), .Y(add_124_carry_21_)
         );
  XOR2X1 U557 ( .A(y2_tmp[20]), .B(add_124_carry_20_), .Y(N622) );
  AND2X1 U558 ( .A(add_124_carry_19_), .B(y2_tmp[19]), .Y(add_124_carry_20_)
         );
  XOR2X1 U559 ( .A(y2_tmp[19]), .B(add_124_carry_19_), .Y(N621) );
  AND2X1 U560 ( .A(add_124_carry_18_), .B(y2_tmp[18]), .Y(add_124_carry_19_)
         );
  XOR2X1 U561 ( .A(y2_tmp[18]), .B(add_124_carry_18_), .Y(N620) );
  AND2X1 U562 ( .A(add_124_carry_17_), .B(y2_tmp[17]), .Y(add_124_carry_18_)
         );
  XOR2X1 U563 ( .A(y2_tmp[17]), .B(add_124_carry_17_), .Y(N619) );
  AND2X1 U564 ( .A(add_124_carry_16_), .B(y2_tmp[16]), .Y(add_124_carry_17_)
         );
  XOR2X1 U565 ( .A(y2_tmp[16]), .B(add_124_carry_16_), .Y(N618) );
  AND2X1 U566 ( .A(add_124_carry_15_), .B(y2_tmp[15]), .Y(add_124_carry_16_)
         );
  XOR2X1 U567 ( .A(y2_tmp[15]), .B(add_124_carry_15_), .Y(N617) );
  AND2X1 U568 ( .A(add_124_carry_14_), .B(y2_tmp[14]), .Y(add_124_carry_15_)
         );
  XOR2X1 U569 ( .A(y2_tmp[14]), .B(add_124_carry_14_), .Y(N616) );
  AND2X1 U570 ( .A(add_124_carry_13_), .B(y2_tmp[13]), .Y(add_124_carry_14_)
         );
  XOR2X1 U571 ( .A(y2_tmp[13]), .B(add_124_carry_13_), .Y(N615) );
  AND2X1 U572 ( .A(add_124_carry_12_), .B(y2_tmp[12]), .Y(add_124_carry_13_)
         );
  XOR2X1 U573 ( .A(y2_tmp[12]), .B(add_124_carry_12_), .Y(N614) );
  AND2X1 U574 ( .A(add_124_carry_11_), .B(y2_tmp[11]), .Y(add_124_carry_12_)
         );
  XOR2X1 U575 ( .A(y2_tmp[11]), .B(add_124_carry_11_), .Y(N613) );
  AND2X1 U576 ( .A(add_124_carry_10_), .B(y2_tmp[10]), .Y(add_124_carry_11_)
         );
  XOR2X1 U577 ( .A(y2_tmp[10]), .B(add_124_carry_10_), .Y(N612) );
  AND2X1 U578 ( .A(add_124_carry_9_), .B(y2_tmp[9]), .Y(add_124_carry_10_) );
  XOR2X1 U579 ( .A(y2_tmp[9]), .B(add_124_carry_9_), .Y(N611) );
  AND2X1 U580 ( .A(add_124_carry_8_), .B(y2_tmp[8]), .Y(add_124_carry_9_) );
  XOR2X1 U581 ( .A(y2_tmp[8]), .B(add_124_carry_8_), .Y(N610) );
  AND2X1 U582 ( .A(y2_tmp[6]), .B(y2_tmp[7]), .Y(add_124_carry_8_) );
  XOR2X1 U583 ( .A(y2_tmp[7]), .B(y2_tmp[6]), .Y(N609) );
  AND2X1 U584 ( .A(add_125_carry_22_), .B(y3_tmp[22]), .Y(add_125_carry_23_)
         );
  XOR2X1 U585 ( .A(y3_tmp[22]), .B(add_125_carry_22_), .Y(N643) );
  AND2X1 U586 ( .A(add_125_carry_21_), .B(y3_tmp[21]), .Y(add_125_carry_22_)
         );
  XOR2X1 U587 ( .A(y3_tmp[21]), .B(add_125_carry_21_), .Y(N642) );
  AND2X1 U588 ( .A(add_125_carry_20_), .B(y3_tmp[20]), .Y(add_125_carry_21_)
         );
  XOR2X1 U589 ( .A(y3_tmp[20]), .B(add_125_carry_20_), .Y(N641) );
  AND2X1 U590 ( .A(add_125_carry_19_), .B(y3_tmp[19]), .Y(add_125_carry_20_)
         );
  XOR2X1 U591 ( .A(y3_tmp[19]), .B(add_125_carry_19_), .Y(N640) );
  AND2X1 U592 ( .A(add_125_carry_18_), .B(y3_tmp[18]), .Y(add_125_carry_19_)
         );
  XOR2X1 U593 ( .A(y3_tmp[18]), .B(add_125_carry_18_), .Y(N639) );
  AND2X1 U594 ( .A(add_125_carry_17_), .B(y3_tmp[17]), .Y(add_125_carry_18_)
         );
  XOR2X1 U595 ( .A(y3_tmp[17]), .B(add_125_carry_17_), .Y(N638) );
  AND2X1 U596 ( .A(add_125_carry_16_), .B(y3_tmp[16]), .Y(add_125_carry_17_)
         );
  XOR2X1 U597 ( .A(y3_tmp[16]), .B(add_125_carry_16_), .Y(N637) );
  AND2X1 U598 ( .A(add_125_carry_15_), .B(y3_tmp[15]), .Y(add_125_carry_16_)
         );
  XOR2X1 U599 ( .A(y3_tmp[15]), .B(add_125_carry_15_), .Y(N636) );
  AND2X1 U600 ( .A(add_125_carry_14_), .B(y3_tmp[14]), .Y(add_125_carry_15_)
         );
  XOR2X1 U601 ( .A(y3_tmp[14]), .B(add_125_carry_14_), .Y(N635) );
  AND2X1 U602 ( .A(add_125_carry_13_), .B(y3_tmp[13]), .Y(add_125_carry_14_)
         );
  XOR2X1 U603 ( .A(y3_tmp[13]), .B(add_125_carry_13_), .Y(N634) );
  AND2X1 U604 ( .A(add_125_carry_12_), .B(y3_tmp[12]), .Y(add_125_carry_13_)
         );
  XOR2X1 U605 ( .A(y3_tmp[12]), .B(add_125_carry_12_), .Y(N633) );
  AND2X1 U606 ( .A(add_125_carry_11_), .B(y3_tmp[11]), .Y(add_125_carry_12_)
         );
  XOR2X1 U607 ( .A(y3_tmp[11]), .B(add_125_carry_11_), .Y(N632) );
  AND2X1 U608 ( .A(add_125_carry_10_), .B(y3_tmp[10]), .Y(add_125_carry_11_)
         );
  XOR2X1 U609 ( .A(y3_tmp[10]), .B(add_125_carry_10_), .Y(N631) );
  AND2X1 U610 ( .A(add_125_carry_9_), .B(y3_tmp[9]), .Y(add_125_carry_10_) );
  XOR2X1 U611 ( .A(y3_tmp[9]), .B(add_125_carry_9_), .Y(N630) );
  AND2X1 U612 ( .A(add_125_carry_8_), .B(y3_tmp[8]), .Y(add_125_carry_9_) );
  XOR2X1 U613 ( .A(y3_tmp[8]), .B(add_125_carry_8_), .Y(N629) );
  AND2X1 U614 ( .A(y3_tmp[6]), .B(y3_tmp[7]), .Y(add_125_carry_8_) );
  XOR2X1 U615 ( .A(y3_tmp[7]), .B(y3_tmp[6]), .Y(N628) );
endmodule


module idct8_shift7_add64_DW01_add_0 ( A, SUM );
  input [28:0] A;
  output [28:0] SUM;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  AND2X2 U1 ( .A(A[27]), .B(n18), .Y(SUM[28]) );
  XOR2X1 U2 ( .A(A[20]), .B(n14), .Y(SUM[20]) );
  XOR2X1 U3 ( .A(A[21]), .B(n15), .Y(SUM[21]) );
  XOR2X1 U4 ( .A(A[22]), .B(n16), .Y(SUM[22]) );
  AND2X2 U5 ( .A(A[9]), .B(n4), .Y(n2) );
  AND2X2 U6 ( .A(A[7]), .B(A[6]), .Y(n3) );
  AND2X2 U7 ( .A(A[8]), .B(n3), .Y(n4) );
  AND2X2 U8 ( .A(A[10]), .B(n2), .Y(n5) );
  AND2X2 U9 ( .A(A[11]), .B(n5), .Y(n6) );
  AND2X2 U10 ( .A(A[12]), .B(n6), .Y(n7) );
  AND2X2 U11 ( .A(A[13]), .B(n7), .Y(n8) );
  AND2X2 U12 ( .A(A[14]), .B(n8), .Y(n9) );
  AND2X2 U13 ( .A(A[15]), .B(n9), .Y(n10) );
  AND2X2 U14 ( .A(A[16]), .B(n10), .Y(n11) );
  AND2X2 U15 ( .A(A[17]), .B(n11), .Y(n12) );
  AND2X2 U16 ( .A(A[18]), .B(n12), .Y(n13) );
  AND2X2 U17 ( .A(A[19]), .B(n13), .Y(n14) );
  AND2X2 U18 ( .A(A[20]), .B(n14), .Y(n15) );
  AND2X2 U19 ( .A(A[21]), .B(n15), .Y(n16) );
  XOR2X1 U20 ( .A(A[15]), .B(n9), .Y(SUM[15]) );
  XOR2X1 U21 ( .A(A[16]), .B(n10), .Y(SUM[16]) );
  XOR2X1 U22 ( .A(A[17]), .B(n11), .Y(SUM[17]) );
  XOR2X1 U23 ( .A(A[18]), .B(n12), .Y(SUM[18]) );
  XOR2X1 U24 ( .A(A[19]), .B(n13), .Y(SUM[19]) );
  XOR2X1 U25 ( .A(A[7]), .B(A[6]), .Y(SUM[7]) );
  XOR2X1 U26 ( .A(A[8]), .B(n3), .Y(SUM[8]) );
  XOR2X1 U27 ( .A(A[9]), .B(n4), .Y(SUM[9]) );
  XOR2X1 U28 ( .A(A[10]), .B(n2), .Y(SUM[10]) );
  XOR2X1 U29 ( .A(A[11]), .B(n5), .Y(SUM[11]) );
  XOR2X1 U30 ( .A(A[12]), .B(n6), .Y(SUM[12]) );
  XOR2X1 U31 ( .A(A[13]), .B(n7), .Y(SUM[13]) );
  XOR2X1 U32 ( .A(A[14]), .B(n8), .Y(SUM[14]) );
  XOR2X1 U33 ( .A(A[23]), .B(n19), .Y(SUM[23]) );
  XOR2X1 U34 ( .A(A[24]), .B(n20), .Y(SUM[24]) );
  XOR2X1 U35 ( .A(A[25]), .B(n21), .Y(SUM[25]) );
  XOR2X1 U36 ( .A(A[26]), .B(n17), .Y(SUM[26]) );
  XOR2X1 U37 ( .A(A[27]), .B(n18), .Y(SUM[27]) );
  AND2X2 U38 ( .A(A[25]), .B(n21), .Y(n17) );
  AND2X2 U39 ( .A(A[26]), .B(n17), .Y(n18) );
  AND2X2 U40 ( .A(A[22]), .B(n16), .Y(n19) );
  AND2X2 U41 ( .A(A[23]), .B(n19), .Y(n20) );
  AND2X2 U42 ( .A(A[24]), .B(n20), .Y(n21) );
endmodule


module idct8_shift7_add64_DW01_add_1 ( A, SUM );
  input [28:0] A;
  output [28:0] SUM;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  AND2X2 U1 ( .A(A[27]), .B(n18), .Y(SUM[28]) );
  XOR2X1 U2 ( .A(A[20]), .B(n14), .Y(SUM[20]) );
  XOR2X1 U3 ( .A(A[21]), .B(n15), .Y(SUM[21]) );
  XOR2X1 U4 ( .A(A[22]), .B(n16), .Y(SUM[22]) );
  AND2X2 U5 ( .A(A[9]), .B(n4), .Y(n2) );
  AND2X2 U6 ( .A(A[7]), .B(A[6]), .Y(n3) );
  AND2X2 U7 ( .A(A[8]), .B(n3), .Y(n4) );
  AND2X2 U8 ( .A(A[10]), .B(n2), .Y(n5) );
  AND2X2 U9 ( .A(A[11]), .B(n5), .Y(n6) );
  AND2X2 U10 ( .A(A[12]), .B(n6), .Y(n7) );
  AND2X2 U11 ( .A(A[13]), .B(n7), .Y(n8) );
  AND2X2 U12 ( .A(A[14]), .B(n8), .Y(n9) );
  AND2X2 U13 ( .A(A[15]), .B(n9), .Y(n10) );
  AND2X2 U14 ( .A(A[16]), .B(n10), .Y(n11) );
  AND2X2 U15 ( .A(A[17]), .B(n11), .Y(n12) );
  AND2X2 U16 ( .A(A[18]), .B(n12), .Y(n13) );
  AND2X2 U17 ( .A(A[19]), .B(n13), .Y(n14) );
  AND2X2 U18 ( .A(A[20]), .B(n14), .Y(n15) );
  AND2X2 U19 ( .A(A[21]), .B(n15), .Y(n16) );
  XOR2X1 U20 ( .A(A[15]), .B(n9), .Y(SUM[15]) );
  XOR2X1 U21 ( .A(A[16]), .B(n10), .Y(SUM[16]) );
  XOR2X1 U22 ( .A(A[17]), .B(n11), .Y(SUM[17]) );
  XOR2X1 U23 ( .A(A[18]), .B(n12), .Y(SUM[18]) );
  XOR2X1 U24 ( .A(A[19]), .B(n13), .Y(SUM[19]) );
  XOR2X1 U25 ( .A(A[7]), .B(A[6]), .Y(SUM[7]) );
  XOR2X1 U26 ( .A(A[8]), .B(n3), .Y(SUM[8]) );
  XOR2X1 U27 ( .A(A[9]), .B(n4), .Y(SUM[9]) );
  XOR2X1 U28 ( .A(A[10]), .B(n2), .Y(SUM[10]) );
  XOR2X1 U29 ( .A(A[11]), .B(n5), .Y(SUM[11]) );
  XOR2X1 U30 ( .A(A[12]), .B(n6), .Y(SUM[12]) );
  XOR2X1 U31 ( .A(A[13]), .B(n7), .Y(SUM[13]) );
  XOR2X1 U32 ( .A(A[14]), .B(n8), .Y(SUM[14]) );
  XOR2X1 U33 ( .A(A[23]), .B(n19), .Y(SUM[23]) );
  XOR2X1 U34 ( .A(A[24]), .B(n20), .Y(SUM[24]) );
  XOR2X1 U35 ( .A(A[25]), .B(n21), .Y(SUM[25]) );
  XOR2X1 U36 ( .A(A[26]), .B(n17), .Y(SUM[26]) );
  XOR2X1 U37 ( .A(A[27]), .B(n18), .Y(SUM[27]) );
  AND2X2 U38 ( .A(A[25]), .B(n21), .Y(n17) );
  AND2X2 U39 ( .A(A[26]), .B(n17), .Y(n18) );
  AND2X2 U40 ( .A(A[22]), .B(n16), .Y(n19) );
  AND2X2 U41 ( .A(A[23]), .B(n19), .Y(n20) );
  AND2X2 U42 ( .A(A[24]), .B(n20), .Y(n21) );
endmodule


module idct8_shift7_add64_DW01_add_2 ( A, SUM );
  input [28:0] A;
  output [28:0] SUM;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  AND2X2 U1 ( .A(A[27]), .B(n18), .Y(SUM[28]) );
  XOR2X1 U2 ( .A(A[20]), .B(n14), .Y(SUM[20]) );
  XOR2X1 U3 ( .A(A[21]), .B(n15), .Y(SUM[21]) );
  XOR2X1 U4 ( .A(A[22]), .B(n16), .Y(SUM[22]) );
  AND2X2 U5 ( .A(A[9]), .B(n4), .Y(n2) );
  AND2X2 U6 ( .A(A[7]), .B(A[6]), .Y(n3) );
  AND2X2 U7 ( .A(A[8]), .B(n3), .Y(n4) );
  AND2X2 U8 ( .A(A[10]), .B(n2), .Y(n5) );
  AND2X2 U9 ( .A(A[11]), .B(n5), .Y(n6) );
  AND2X2 U10 ( .A(A[12]), .B(n6), .Y(n7) );
  AND2X2 U11 ( .A(A[13]), .B(n7), .Y(n8) );
  AND2X2 U12 ( .A(A[14]), .B(n8), .Y(n9) );
  AND2X2 U13 ( .A(A[15]), .B(n9), .Y(n10) );
  AND2X2 U14 ( .A(A[16]), .B(n10), .Y(n11) );
  AND2X2 U15 ( .A(A[17]), .B(n11), .Y(n12) );
  AND2X2 U16 ( .A(A[18]), .B(n12), .Y(n13) );
  AND2X2 U17 ( .A(A[19]), .B(n13), .Y(n14) );
  AND2X2 U18 ( .A(A[20]), .B(n14), .Y(n15) );
  AND2X2 U19 ( .A(A[21]), .B(n15), .Y(n16) );
  XOR2X1 U20 ( .A(A[15]), .B(n9), .Y(SUM[15]) );
  XOR2X1 U21 ( .A(A[16]), .B(n10), .Y(SUM[16]) );
  XOR2X1 U22 ( .A(A[17]), .B(n11), .Y(SUM[17]) );
  XOR2X1 U23 ( .A(A[18]), .B(n12), .Y(SUM[18]) );
  XOR2X1 U24 ( .A(A[19]), .B(n13), .Y(SUM[19]) );
  XOR2X1 U25 ( .A(A[7]), .B(A[6]), .Y(SUM[7]) );
  XOR2X1 U26 ( .A(A[8]), .B(n3), .Y(SUM[8]) );
  XOR2X1 U27 ( .A(A[9]), .B(n4), .Y(SUM[9]) );
  XOR2X1 U28 ( .A(A[10]), .B(n2), .Y(SUM[10]) );
  XOR2X1 U29 ( .A(A[11]), .B(n5), .Y(SUM[11]) );
  XOR2X1 U30 ( .A(A[12]), .B(n6), .Y(SUM[12]) );
  XOR2X1 U31 ( .A(A[13]), .B(n7), .Y(SUM[13]) );
  XOR2X1 U32 ( .A(A[14]), .B(n8), .Y(SUM[14]) );
  XOR2X1 U33 ( .A(A[23]), .B(n19), .Y(SUM[23]) );
  XOR2X1 U34 ( .A(A[24]), .B(n20), .Y(SUM[24]) );
  XOR2X1 U35 ( .A(A[25]), .B(n21), .Y(SUM[25]) );
  XOR2X1 U36 ( .A(A[26]), .B(n17), .Y(SUM[26]) );
  XOR2X1 U37 ( .A(A[27]), .B(n18), .Y(SUM[27]) );
  AND2X2 U38 ( .A(A[25]), .B(n21), .Y(n17) );
  AND2X2 U39 ( .A(A[26]), .B(n17), .Y(n18) );
  AND2X2 U40 ( .A(A[22]), .B(n16), .Y(n19) );
  AND2X2 U41 ( .A(A[23]), .B(n19), .Y(n20) );
  AND2X2 U42 ( .A(A[24]), .B(n20), .Y(n21) );
endmodule


module idct8_shift7_add64_DW01_add_3 ( A, SUM );
  input [28:0] A;
  output [28:0] SUM;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  AND2X2 U1 ( .A(A[27]), .B(n18), .Y(SUM[28]) );
  XOR2X1 U2 ( .A(A[20]), .B(n14), .Y(SUM[20]) );
  XOR2X1 U3 ( .A(A[21]), .B(n15), .Y(SUM[21]) );
  XOR2X1 U4 ( .A(A[22]), .B(n16), .Y(SUM[22]) );
  AND2X2 U5 ( .A(A[9]), .B(n4), .Y(n2) );
  AND2X2 U6 ( .A(A[7]), .B(A[6]), .Y(n3) );
  AND2X2 U7 ( .A(A[8]), .B(n3), .Y(n4) );
  AND2X2 U8 ( .A(A[10]), .B(n2), .Y(n5) );
  AND2X2 U9 ( .A(A[11]), .B(n5), .Y(n6) );
  AND2X2 U10 ( .A(A[12]), .B(n6), .Y(n7) );
  AND2X2 U11 ( .A(A[13]), .B(n7), .Y(n8) );
  AND2X2 U12 ( .A(A[14]), .B(n8), .Y(n9) );
  AND2X2 U13 ( .A(A[15]), .B(n9), .Y(n10) );
  AND2X2 U14 ( .A(A[16]), .B(n10), .Y(n11) );
  AND2X2 U15 ( .A(A[17]), .B(n11), .Y(n12) );
  AND2X2 U16 ( .A(A[18]), .B(n12), .Y(n13) );
  AND2X2 U17 ( .A(A[19]), .B(n13), .Y(n14) );
  AND2X2 U18 ( .A(A[20]), .B(n14), .Y(n15) );
  AND2X2 U19 ( .A(A[21]), .B(n15), .Y(n16) );
  XOR2X1 U20 ( .A(A[15]), .B(n9), .Y(SUM[15]) );
  XOR2X1 U21 ( .A(A[16]), .B(n10), .Y(SUM[16]) );
  XOR2X1 U22 ( .A(A[17]), .B(n11), .Y(SUM[17]) );
  XOR2X1 U23 ( .A(A[18]), .B(n12), .Y(SUM[18]) );
  XOR2X1 U24 ( .A(A[19]), .B(n13), .Y(SUM[19]) );
  XOR2X1 U25 ( .A(A[7]), .B(A[6]), .Y(SUM[7]) );
  XOR2X1 U26 ( .A(A[8]), .B(n3), .Y(SUM[8]) );
  XOR2X1 U27 ( .A(A[9]), .B(n4), .Y(SUM[9]) );
  XOR2X1 U28 ( .A(A[10]), .B(n2), .Y(SUM[10]) );
  XOR2X1 U29 ( .A(A[11]), .B(n5), .Y(SUM[11]) );
  XOR2X1 U30 ( .A(A[12]), .B(n6), .Y(SUM[12]) );
  XOR2X1 U31 ( .A(A[13]), .B(n7), .Y(SUM[13]) );
  XOR2X1 U32 ( .A(A[14]), .B(n8), .Y(SUM[14]) );
  XOR2X1 U33 ( .A(A[23]), .B(n19), .Y(SUM[23]) );
  XOR2X1 U34 ( .A(A[24]), .B(n20), .Y(SUM[24]) );
  XOR2X1 U35 ( .A(A[25]), .B(n21), .Y(SUM[25]) );
  XOR2X1 U36 ( .A(A[26]), .B(n17), .Y(SUM[26]) );
  XOR2X1 U37 ( .A(A[27]), .B(n18), .Y(SUM[27]) );
  AND2X2 U38 ( .A(A[25]), .B(n21), .Y(n17) );
  AND2X2 U39 ( .A(A[26]), .B(n17), .Y(n18) );
  AND2X2 U40 ( .A(A[22]), .B(n16), .Y(n19) );
  AND2X2 U41 ( .A(A[23]), .B(n19), .Y(n20) );
  AND2X2 U42 ( .A(A[24]), .B(n20), .Y(n21) );
endmodule


module idct8_shift7_add64_DW01_add_4 ( A, SUM );
  input [28:0] A;
  output [28:0] SUM;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  AND2X2 U1 ( .A(A[27]), .B(n18), .Y(SUM[28]) );
  AND2X2 U2 ( .A(A[7]), .B(A[6]), .Y(n2) );
  AND2X2 U3 ( .A(A[8]), .B(n2), .Y(n3) );
  AND2X2 U4 ( .A(A[9]), .B(n3), .Y(n4) );
  AND2X2 U5 ( .A(A[10]), .B(n4), .Y(n5) );
  AND2X2 U6 ( .A(A[11]), .B(n5), .Y(n6) );
  AND2X2 U7 ( .A(A[12]), .B(n6), .Y(n7) );
  AND2X2 U8 ( .A(A[13]), .B(n7), .Y(n8) );
  AND2X2 U9 ( .A(A[14]), .B(n8), .Y(n9) );
  AND2X2 U10 ( .A(A[15]), .B(n9), .Y(n10) );
  AND2X2 U11 ( .A(A[16]), .B(n10), .Y(n11) );
  AND2X2 U12 ( .A(A[17]), .B(n11), .Y(n12) );
  AND2X2 U13 ( .A(A[18]), .B(n12), .Y(n13) );
  AND2X2 U14 ( .A(A[19]), .B(n13), .Y(n14) );
  AND2X2 U15 ( .A(A[20]), .B(n14), .Y(n15) );
  AND2X2 U16 ( .A(A[21]), .B(n15), .Y(n16) );
  XOR2X1 U17 ( .A(A[18]), .B(n12), .Y(SUM[18]) );
  XOR2X1 U18 ( .A(A[19]), .B(n13), .Y(SUM[19]) );
  XOR2X1 U19 ( .A(A[20]), .B(n14), .Y(SUM[20]) );
  XOR2X1 U20 ( .A(A[21]), .B(n15), .Y(SUM[21]) );
  XOR2X1 U21 ( .A(A[22]), .B(n16), .Y(SUM[22]) );
  XOR2X1 U22 ( .A(A[13]), .B(n7), .Y(SUM[13]) );
  XOR2X1 U23 ( .A(A[14]), .B(n8), .Y(SUM[14]) );
  XOR2X1 U24 ( .A(A[15]), .B(n9), .Y(SUM[15]) );
  XOR2X1 U25 ( .A(A[16]), .B(n10), .Y(SUM[16]) );
  XOR2X1 U26 ( .A(A[17]), .B(n11), .Y(SUM[17]) );
  XOR2X1 U27 ( .A(A[7]), .B(A[6]), .Y(SUM[7]) );
  XOR2X1 U28 ( .A(A[8]), .B(n2), .Y(SUM[8]) );
  XOR2X1 U29 ( .A(A[9]), .B(n3), .Y(SUM[9]) );
  XOR2X1 U30 ( .A(A[10]), .B(n4), .Y(SUM[10]) );
  XOR2X1 U31 ( .A(A[11]), .B(n5), .Y(SUM[11]) );
  XOR2X1 U32 ( .A(A[12]), .B(n6), .Y(SUM[12]) );
  XOR2X1 U33 ( .A(A[23]), .B(n19), .Y(SUM[23]) );
  XOR2X1 U34 ( .A(A[24]), .B(n20), .Y(SUM[24]) );
  XOR2X1 U35 ( .A(A[25]), .B(n21), .Y(SUM[25]) );
  XOR2X1 U36 ( .A(A[26]), .B(n17), .Y(SUM[26]) );
  XOR2X1 U37 ( .A(A[27]), .B(n18), .Y(SUM[27]) );
  AND2X2 U38 ( .A(A[25]), .B(n21), .Y(n17) );
  AND2X2 U39 ( .A(A[26]), .B(n17), .Y(n18) );
  AND2X2 U40 ( .A(A[22]), .B(n16), .Y(n19) );
  AND2X2 U41 ( .A(A[23]), .B(n19), .Y(n20) );
  AND2X2 U42 ( .A(A[24]), .B(n20), .Y(n21) );
endmodule


module idct8_shift7_add64_DW01_add_5 ( A, SUM );
  input [28:0] A;
  output [28:0] SUM;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  AND2X2 U1 ( .A(A[27]), .B(n18), .Y(SUM[28]) );
  AND2X2 U2 ( .A(A[7]), .B(A[6]), .Y(n2) );
  AND2X2 U3 ( .A(A[8]), .B(n2), .Y(n3) );
  AND2X2 U4 ( .A(A[9]), .B(n3), .Y(n4) );
  AND2X2 U5 ( .A(A[10]), .B(n4), .Y(n5) );
  AND2X2 U6 ( .A(A[11]), .B(n5), .Y(n6) );
  AND2X2 U7 ( .A(A[12]), .B(n6), .Y(n7) );
  AND2X2 U8 ( .A(A[13]), .B(n7), .Y(n8) );
  AND2X2 U9 ( .A(A[14]), .B(n8), .Y(n9) );
  AND2X2 U10 ( .A(A[15]), .B(n9), .Y(n10) );
  AND2X2 U11 ( .A(A[16]), .B(n10), .Y(n11) );
  AND2X2 U12 ( .A(A[17]), .B(n11), .Y(n12) );
  AND2X2 U13 ( .A(A[18]), .B(n12), .Y(n13) );
  AND2X2 U14 ( .A(A[19]), .B(n13), .Y(n14) );
  AND2X2 U15 ( .A(A[20]), .B(n14), .Y(n15) );
  AND2X2 U16 ( .A(A[21]), .B(n15), .Y(n16) );
  XOR2X1 U17 ( .A(A[18]), .B(n12), .Y(SUM[18]) );
  XOR2X1 U18 ( .A(A[19]), .B(n13), .Y(SUM[19]) );
  XOR2X1 U19 ( .A(A[20]), .B(n14), .Y(SUM[20]) );
  XOR2X1 U20 ( .A(A[21]), .B(n15), .Y(SUM[21]) );
  XOR2X1 U21 ( .A(A[22]), .B(n16), .Y(SUM[22]) );
  XOR2X1 U22 ( .A(A[13]), .B(n7), .Y(SUM[13]) );
  XOR2X1 U23 ( .A(A[14]), .B(n8), .Y(SUM[14]) );
  XOR2X1 U24 ( .A(A[15]), .B(n9), .Y(SUM[15]) );
  XOR2X1 U25 ( .A(A[16]), .B(n10), .Y(SUM[16]) );
  XOR2X1 U26 ( .A(A[17]), .B(n11), .Y(SUM[17]) );
  XOR2X1 U27 ( .A(A[7]), .B(A[6]), .Y(SUM[7]) );
  XOR2X1 U28 ( .A(A[8]), .B(n2), .Y(SUM[8]) );
  XOR2X1 U29 ( .A(A[9]), .B(n3), .Y(SUM[9]) );
  XOR2X1 U30 ( .A(A[10]), .B(n4), .Y(SUM[10]) );
  XOR2X1 U31 ( .A(A[11]), .B(n5), .Y(SUM[11]) );
  XOR2X1 U32 ( .A(A[12]), .B(n6), .Y(SUM[12]) );
  XOR2X1 U33 ( .A(A[23]), .B(n19), .Y(SUM[23]) );
  XOR2X1 U34 ( .A(A[24]), .B(n20), .Y(SUM[24]) );
  XOR2X1 U35 ( .A(A[25]), .B(n21), .Y(SUM[25]) );
  XOR2X1 U36 ( .A(A[26]), .B(n17), .Y(SUM[26]) );
  XOR2X1 U37 ( .A(A[27]), .B(n18), .Y(SUM[27]) );
  AND2X2 U38 ( .A(A[25]), .B(n21), .Y(n17) );
  AND2X2 U39 ( .A(A[26]), .B(n17), .Y(n18) );
  AND2X2 U40 ( .A(A[22]), .B(n16), .Y(n19) );
  AND2X2 U41 ( .A(A[23]), .B(n19), .Y(n20) );
  AND2X2 U42 ( .A(A[24]), .B(n20), .Y(n21) );
endmodule


module idct8_shift7_add64_DW01_add_6 ( A, SUM );
  input [28:0] A;
  output [28:0] SUM;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  AND2X2 U1 ( .A(A[27]), .B(n18), .Y(SUM[28]) );
  AND2X2 U2 ( .A(A[7]), .B(A[6]), .Y(n2) );
  AND2X2 U3 ( .A(A[8]), .B(n2), .Y(n3) );
  AND2X2 U4 ( .A(A[9]), .B(n3), .Y(n4) );
  AND2X2 U5 ( .A(A[10]), .B(n4), .Y(n5) );
  AND2X2 U6 ( .A(A[11]), .B(n5), .Y(n6) );
  AND2X2 U7 ( .A(A[12]), .B(n6), .Y(n7) );
  AND2X2 U8 ( .A(A[13]), .B(n7), .Y(n8) );
  AND2X2 U9 ( .A(A[14]), .B(n8), .Y(n9) );
  AND2X2 U10 ( .A(A[15]), .B(n9), .Y(n10) );
  AND2X2 U11 ( .A(A[16]), .B(n10), .Y(n11) );
  AND2X2 U12 ( .A(A[17]), .B(n11), .Y(n12) );
  AND2X2 U13 ( .A(A[18]), .B(n12), .Y(n13) );
  AND2X2 U14 ( .A(A[19]), .B(n13), .Y(n14) );
  AND2X2 U15 ( .A(A[20]), .B(n14), .Y(n15) );
  AND2X2 U16 ( .A(A[21]), .B(n15), .Y(n16) );
  XOR2X1 U17 ( .A(A[18]), .B(n12), .Y(SUM[18]) );
  XOR2X1 U18 ( .A(A[19]), .B(n13), .Y(SUM[19]) );
  XOR2X1 U19 ( .A(A[20]), .B(n14), .Y(SUM[20]) );
  XOR2X1 U20 ( .A(A[21]), .B(n15), .Y(SUM[21]) );
  XOR2X1 U21 ( .A(A[22]), .B(n16), .Y(SUM[22]) );
  XOR2X1 U22 ( .A(A[13]), .B(n7), .Y(SUM[13]) );
  XOR2X1 U23 ( .A(A[14]), .B(n8), .Y(SUM[14]) );
  XOR2X1 U24 ( .A(A[15]), .B(n9), .Y(SUM[15]) );
  XOR2X1 U25 ( .A(A[16]), .B(n10), .Y(SUM[16]) );
  XOR2X1 U26 ( .A(A[17]), .B(n11), .Y(SUM[17]) );
  XOR2X1 U27 ( .A(A[7]), .B(A[6]), .Y(SUM[7]) );
  XOR2X1 U28 ( .A(A[8]), .B(n2), .Y(SUM[8]) );
  XOR2X1 U29 ( .A(A[9]), .B(n3), .Y(SUM[9]) );
  XOR2X1 U30 ( .A(A[10]), .B(n4), .Y(SUM[10]) );
  XOR2X1 U31 ( .A(A[11]), .B(n5), .Y(SUM[11]) );
  XOR2X1 U32 ( .A(A[12]), .B(n6), .Y(SUM[12]) );
  XOR2X1 U33 ( .A(A[23]), .B(n19), .Y(SUM[23]) );
  XOR2X1 U34 ( .A(A[24]), .B(n20), .Y(SUM[24]) );
  XOR2X1 U35 ( .A(A[25]), .B(n21), .Y(SUM[25]) );
  XOR2X1 U36 ( .A(A[26]), .B(n17), .Y(SUM[26]) );
  XOR2X1 U37 ( .A(A[27]), .B(n18), .Y(SUM[27]) );
  AND2X2 U38 ( .A(A[25]), .B(n21), .Y(n17) );
  AND2X2 U39 ( .A(A[26]), .B(n17), .Y(n18) );
  AND2X2 U40 ( .A(A[22]), .B(n16), .Y(n19) );
  AND2X2 U41 ( .A(A[23]), .B(n19), .Y(n20) );
  AND2X2 U42 ( .A(A[24]), .B(n20), .Y(n21) );
endmodule


module idct8_shift7_add64_DW01_add_7 ( A, SUM );
  input [28:0] A;
  output [28:0] SUM;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  AND2X2 U1 ( .A(A[27]), .B(n18), .Y(SUM[28]) );
  AND2X2 U2 ( .A(A[7]), .B(A[6]), .Y(n2) );
  AND2X2 U3 ( .A(A[8]), .B(n2), .Y(n3) );
  AND2X2 U4 ( .A(A[9]), .B(n3), .Y(n4) );
  AND2X2 U5 ( .A(A[10]), .B(n4), .Y(n5) );
  AND2X2 U6 ( .A(A[11]), .B(n5), .Y(n6) );
  AND2X2 U7 ( .A(A[12]), .B(n6), .Y(n7) );
  AND2X2 U8 ( .A(A[13]), .B(n7), .Y(n8) );
  AND2X2 U9 ( .A(A[14]), .B(n8), .Y(n9) );
  AND2X2 U10 ( .A(A[15]), .B(n9), .Y(n10) );
  AND2X2 U11 ( .A(A[16]), .B(n10), .Y(n11) );
  AND2X2 U12 ( .A(A[17]), .B(n11), .Y(n12) );
  AND2X2 U13 ( .A(A[18]), .B(n12), .Y(n13) );
  AND2X2 U14 ( .A(A[19]), .B(n13), .Y(n14) );
  AND2X2 U15 ( .A(A[20]), .B(n14), .Y(n15) );
  AND2X2 U16 ( .A(A[21]), .B(n15), .Y(n16) );
  XOR2X1 U17 ( .A(A[18]), .B(n12), .Y(SUM[18]) );
  XOR2X1 U18 ( .A(A[19]), .B(n13), .Y(SUM[19]) );
  XOR2X1 U19 ( .A(A[20]), .B(n14), .Y(SUM[20]) );
  XOR2X1 U20 ( .A(A[21]), .B(n15), .Y(SUM[21]) );
  XOR2X1 U21 ( .A(A[22]), .B(n16), .Y(SUM[22]) );
  XOR2X1 U22 ( .A(A[13]), .B(n7), .Y(SUM[13]) );
  XOR2X1 U23 ( .A(A[14]), .B(n8), .Y(SUM[14]) );
  XOR2X1 U24 ( .A(A[15]), .B(n9), .Y(SUM[15]) );
  XOR2X1 U25 ( .A(A[16]), .B(n10), .Y(SUM[16]) );
  XOR2X1 U26 ( .A(A[17]), .B(n11), .Y(SUM[17]) );
  XOR2X1 U27 ( .A(A[7]), .B(A[6]), .Y(SUM[7]) );
  XOR2X1 U28 ( .A(A[8]), .B(n2), .Y(SUM[8]) );
  XOR2X1 U29 ( .A(A[9]), .B(n3), .Y(SUM[9]) );
  XOR2X1 U30 ( .A(A[10]), .B(n4), .Y(SUM[10]) );
  XOR2X1 U31 ( .A(A[11]), .B(n5), .Y(SUM[11]) );
  XOR2X1 U32 ( .A(A[12]), .B(n6), .Y(SUM[12]) );
  XOR2X1 U33 ( .A(A[23]), .B(n19), .Y(SUM[23]) );
  XOR2X1 U34 ( .A(A[24]), .B(n20), .Y(SUM[24]) );
  XOR2X1 U35 ( .A(A[25]), .B(n21), .Y(SUM[25]) );
  XOR2X1 U36 ( .A(A[26]), .B(n17), .Y(SUM[26]) );
  XOR2X1 U37 ( .A(A[27]), .B(n18), .Y(SUM[27]) );
  AND2X2 U38 ( .A(A[25]), .B(n21), .Y(n17) );
  AND2X2 U39 ( .A(A[26]), .B(n17), .Y(n18) );
  AND2X2 U40 ( .A(A[22]), .B(n16), .Y(n19) );
  AND2X2 U41 ( .A(A[23]), .B(n19), .Y(n20) );
  AND2X2 U42 ( .A(A[24]), .B(n20), .Y(n21) );
endmodule


module idct8_shift7_add64_DW01_add_8 ( A, B, SUM );
  input [25:0] A;
  input [25:0] B;
  output [25:0] SUM;
  wire   n1, n2;
  wire   [25:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  XOR3X2 U1_25 ( .A(A[25]), .B(B[25]), .C(carry[25]), .Y(SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  INVX1 U1 ( .A(A[0]), .Y(n2) );
  XNOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  NAND2X1 U3 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U4 ( .A(B[0]), .Y(n1) );
endmodule


module idct8_shift7_add64_DW01_add_9 ( A, B, SUM );
  input [25:0] A;
  input [25:0] B;
  output [25:0] SUM;
  wire   n1, n2;
  wire   [25:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  XOR3X2 U1_25 ( .A(A[25]), .B(B[25]), .C(carry[25]), .Y(SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  INVX1 U1 ( .A(A[0]), .Y(n2) );
  XNOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  NAND2X1 U3 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U4 ( .A(B[0]), .Y(n1) );
endmodule


module idct8_shift7_add64_DW01_add_10 ( A, B, SUM );
  input [25:0] A;
  input [25:0] B;
  output [25:0] SUM;
  wire   n1, n2;
  wire   [25:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  XOR3X2 U1_25 ( .A(A[25]), .B(B[25]), .C(carry[25]), .Y(SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  INVX1 U1 ( .A(A[0]), .Y(n2) );
  XNOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  NAND2X1 U3 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U4 ( .A(B[0]), .Y(n1) );
endmodule


module idct8_shift7_add64_DW01_add_11 ( A, B, SUM );
  input [25:0] A;
  input [25:0] B;
  output [25:0] SUM;
  wire   n1, n2;
  wire   [25:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  XOR3X2 U1_25 ( .A(A[25]), .B(B[25]), .C(carry[25]), .Y(SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  INVX1 U1 ( .A(A[0]), .Y(n2) );
  XNOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  NAND2X1 U3 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U4 ( .A(B[0]), .Y(n1) );
endmodule


module idct8_shift7_add64_DW01_add_12 ( A, B, SUM );
  input [25:0] A;
  input [25:0] B;
  output [25:0] SUM;
  wire   n1;
  wire   [25:2] carry;

  XOR3X2 U1_25 ( .A(A[25]), .B(B[25]), .C(carry[25]), .Y(SUM[25]) );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module idct8_shift7_add64_DW01_add_13 ( A, B, SUM );
  input [25:0] A;
  input [25:0] B;
  output [25:0] SUM;
  wire   n1;
  wire   [25:2] carry;

  XOR3X2 U1_25 ( .A(A[25]), .B(B[25]), .C(carry[25]), .Y(SUM[25]) );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module idct8_shift7_add64_DW01_add_14 ( A, B, SUM );
  input [25:0] A;
  input [25:0] B;
  output [25:0] SUM;
  wire   n1;
  wire   [25:2] carry;

  XOR3X2 U1_25 ( .A(A[25]), .B(B[25]), .C(carry[25]), .Y(SUM[25]) );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module idct8_shift7_add64_DW01_add_15 ( A, B, SUM );
  input [25:0] A;
  input [25:0] B;
  output [25:0] SUM;
  wire   n1;
  wire   [25:2] carry;

  XOR3X2 U1_25 ( .A(A[25]), .B(B[25]), .C(carry[25]), .Y(SUM[25]) );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module idct8_shift7_add64_DW01_add_16 ( A, B, SUM );
  input [24:0] A;
  input [24:0] B;
  output [24:0] SUM;
  wire   n1;
  wire   [24:2] carry;

  XOR3X2 U1_24 ( .A(A[24]), .B(B[24]), .C(carry[24]), .Y(SUM[24]) );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module idct8_shift7_add64_DW01_add_17 ( A, B, SUM );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  wire   n1;
  wire   [23:2] carry;

  XOR3X2 U1_23 ( .A(A[23]), .B(B[23]), .C(carry[23]), .Y(SUM[23]) );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module idct8_shift7_add64_DW01_add_18 ( A, B, SUM );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;

  wire   [23:1] carry;

  XOR3X2 U1_23 ( .A(A[23]), .B(B[23]), .C(carry[23]), .Y(SUM[23]) );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(1'b0), .CO(carry[2]), .S(SUM[1]) );
  XOR2X1 U1 ( .A(1'b0), .B(A[0]), .Y(SUM[0]) );
endmodule


module idct8_shift7_add64_DW01_add_19 ( A, B, SUM );
  input [24:0] A;
  input [24:0] B;
  output [24:0] SUM;
  wire   n1;
  wire   [24:2] carry;

  XOR3X2 U1_24 ( .A(A[24]), .B(B[24]), .C(carry[24]), .Y(SUM[24]) );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module idct8_shift7_add64_DW01_add_20 ( A, B, SUM );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  wire   n1, n2;
  wire   [23:1] carry;

  XOR3X2 U1_23 ( .A(A[23]), .B(B[23]), .C(carry[23]), .Y(SUM[23]) );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  INVX1 U1 ( .A(B[0]), .Y(n1) );
  NAND2X1 U2 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U3 ( .A(A[0]), .Y(n2) );
  XNOR2X1 U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module idct8_shift7_add64_DW01_add_21 ( A, B, SUM );
  input [24:0] A;
  input [24:0] B;
  output [24:0] SUM;
  wire   n1;
  wire   [24:2] carry;

  XOR3X2 U1_24 ( .A(A[24]), .B(B[24]), .C(carry[24]), .Y(SUM[24]) );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module idct8_shift7_add64_DW01_add_22 ( A, B, SUM );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  wire   n1;
  wire   [23:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  XOR3X2 U1_23 ( .A(A[23]), .B(B[23]), .C(carry[23]), .Y(SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  CLKINVX8 U1 ( .A(n1), .Y(carry[1]) );
  CLKINVX8 U2 ( .A(B[0]), .Y(SUM[0]) );
  INVX1 U3 ( .A(B[0]), .Y(n1) );
endmodule


module idct8_shift7_add64_DW01_add_23 ( A, B, SUM );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  wire   n1;
  wire   [23:2] carry;

  XOR3X2 U1_23 ( .A(A[23]), .B(B[23]), .C(carry[23]), .Y(SUM[23]) );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module idct8_shift7_add64_DW01_add_24 ( A, B, SUM );
  input [24:0] A;
  input [24:0] B;
  output [24:0] SUM;
  wire   n1;
  wire   [24:2] carry;

  XOR3X2 U1_24 ( .A(A[24]), .B(B[24]), .C(carry[24]), .Y(SUM[24]) );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module idct8_shift7_add64_DW01_add_25 ( A, B, SUM );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  wire   n1, n2;
  wire   [23:1] carry;

  XOR3X2 U1_23 ( .A(A[23]), .B(B[23]), .C(carry[23]), .Y(SUM[23]) );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  INVX1 U1 ( .A(B[0]), .Y(n1) );
  NAND2X1 U2 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U3 ( .A(A[0]), .Y(n2) );
  XNOR2X1 U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module idct8_shift7_add64_DW01_add_26 ( A, B, SUM );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  wire   n1;
  wire   [23:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  XOR3X2 U1_23 ( .A(A[23]), .B(B[23]), .C(carry[23]), .Y(SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  CLKINVX8 U1 ( .A(n1), .Y(carry[1]) );
  CLKINVX8 U2 ( .A(B[0]), .Y(SUM[0]) );
  INVX1 U3 ( .A(B[0]), .Y(n1) );
endmodule


module idct8_shift7_add64_DW01_add_27 ( A, B, SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n1;
  wire   [20:6] carry;

  XOR3X2 U1_20 ( .A(A[20]), .B(B[20]), .C(carry[20]), .Y(SUM[20]) );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(n1), .CO(carry[6]), .S(SUM[5]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  AND2X2 U1 ( .A(B[4]), .B(A[4]), .Y(n1) );
  XOR2X1 U2 ( .A(B[4]), .B(A[4]), .Y(SUM[4]) );
  BUFX3 U3 ( .A(B[1]), .Y(SUM[1]) );
  BUFX3 U4 ( .A(B[2]), .Y(SUM[2]) );
  BUFX3 U5 ( .A(B[3]), .Y(SUM[3]) );
endmodule


module idct8_shift7_add64_DW01_add_28 ( A, B, SUM );
  input [21:0] A;
  input [21:0] B;
  output [21:0] SUM;
  wire   n1;
  wire   [21:7] carry;

  XOR3X2 U1_21 ( .A(A[21]), .B(B[21]), .C(carry[21]), .Y(SUM[21]) );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(n1), .CO(carry[7]), .S(SUM[6]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  AND2X2 U1 ( .A(B[5]), .B(A[5]), .Y(n1) );
  XOR2X1 U2 ( .A(B[5]), .B(A[5]), .Y(SUM[5]) );
  BUFX3 U3 ( .A(B[1]), .Y(SUM[1]) );
  BUFX3 U4 ( .A(B[2]), .Y(SUM[2]) );
  BUFX3 U5 ( .A(B[3]), .Y(SUM[3]) );
  BUFX3 U6 ( .A(B[4]), .Y(SUM[4]) );
endmodule


module idct8_shift7_add64_DW01_add_29 ( A, B, SUM );
  input [22:0] A;
  input [22:0] B;
  output [22:0] SUM;

  wire   [22:1] carry;

  XOR3X2 U1_22 ( .A(A[22]), .B(B[22]), .C(carry[22]), .Y(SUM[22]) );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(1'b0), .CO(carry[2]), .S(SUM[1]) );
  XOR2X1 U1 ( .A(1'b0), .B(A[0]), .Y(SUM[0]) );
endmodule


module idct8_shift7_add64_DW01_add_30 ( A, B, SUM );
  input [22:0] A;
  input [22:0] B;
  output [22:0] SUM;

  wire   [22:1] carry;

  XOR3X2 U1_22 ( .A(A[22]), .B(B[22]), .C(carry[22]), .Y(SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_1 ( .A(A[1]), .B(1'b0), .CI(1'b0), .S(SUM[1]) );
  ADDFX2 U1_2 ( .A(A[2]), .B(1'b0), .CI(1'b0), .S(SUM[2]) );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(1'b0), .CO(carry[4]), .S(SUM[3]) );
  XOR2X1 U1 ( .A(1'b0), .B(A[0]), .Y(SUM[0]) );
endmodule


module idct8_shift7_add64_DW01_add_31 ( A, B, SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n1;
  wire   [20:6] carry;

  XOR3X2 U1_20 ( .A(A[20]), .B(B[20]), .C(carry[20]), .Y(SUM[20]) );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(n1), .CO(carry[6]), .S(SUM[5]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  AND2X2 U1 ( .A(B[4]), .B(A[4]), .Y(n1) );
  XOR2X1 U2 ( .A(B[4]), .B(A[4]), .Y(SUM[4]) );
  BUFX3 U3 ( .A(B[1]), .Y(SUM[1]) );
  BUFX3 U4 ( .A(B[2]), .Y(SUM[2]) );
  BUFX3 U5 ( .A(B[3]), .Y(SUM[3]) );
endmodule


module idct8_shift7_add64_DW01_add_32 ( A, B, SUM );
  input [21:0] A;
  input [21:0] B;
  output [21:0] SUM;
  wire   n1;
  wire   [21:7] carry;

  XOR3X2 U1_21 ( .A(A[21]), .B(B[21]), .C(carry[21]), .Y(SUM[21]) );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(n1), .CO(carry[7]), .S(SUM[6]) );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  AND2X2 U1 ( .A(B[5]), .B(A[5]), .Y(n1) );
  XOR2X1 U2 ( .A(B[5]), .B(A[5]), .Y(SUM[5]) );
  BUFX3 U3 ( .A(B[4]), .Y(SUM[4]) );
  BUFX3 U4 ( .A(B[3]), .Y(SUM[3]) );
  BUFX3 U5 ( .A(B[2]), .Y(SUM[2]) );
  BUFX3 U6 ( .A(B[1]), .Y(SUM[1]) );
endmodule


module idct8_shift7_add64_DW01_add_33 ( A, B, SUM );
  input [22:0] A;
  input [22:0] B;
  output [22:0] SUM;

  wire   [22:1] carry;

  XOR3X2 U1_22 ( .A(A[22]), .B(B[22]), .C(carry[22]), .Y(SUM[22]) );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(1'b0), .CO(carry[2]), .S(SUM[1]) );
  XOR2X1 U1 ( .A(1'b0), .B(A[0]), .Y(SUM[0]) );
endmodule


module idct8_shift7_add64_DW01_add_34 ( A, B, SUM );
  input [22:0] A;
  input [22:0] B;
  output [22:0] SUM;

  wire   [22:1] carry;

  XOR3X2 U1_22 ( .A(A[22]), .B(B[22]), .C(carry[22]), .Y(SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_1 ( .A(A[1]), .B(1'b0), .CI(1'b0), .S(SUM[1]) );
  ADDFX2 U1_2 ( .A(A[2]), .B(1'b0), .CI(1'b0), .S(SUM[2]) );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(1'b0), .CO(carry[4]), .S(SUM[3]) );
  XOR2X1 U1 ( .A(1'b0), .B(A[0]), .Y(SUM[0]) );
endmodule


module idct8_shift7_add64_DW01_add_35 ( A, B, SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n1;
  wire   [20:6] carry;

  XOR3X2 U1_20 ( .A(A[20]), .B(B[20]), .C(carry[20]), .Y(SUM[20]) );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(n1), .CO(carry[6]), .S(SUM[5]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  AND2X2 U1 ( .A(B[4]), .B(A[4]), .Y(n1) );
  XOR2X1 U2 ( .A(B[4]), .B(A[4]), .Y(SUM[4]) );
  BUFX3 U3 ( .A(B[1]), .Y(SUM[1]) );
  BUFX3 U4 ( .A(B[2]), .Y(SUM[2]) );
  BUFX3 U5 ( .A(B[3]), .Y(SUM[3]) );
endmodule


module idct8_shift7_add64_DW01_add_36 ( A, B, SUM );
  input [21:0] A;
  input [21:0] B;
  output [21:0] SUM;
  wire   n1;
  wire   [21:7] carry;

  XOR3X2 U1_21 ( .A(A[21]), .B(B[21]), .C(carry[21]), .Y(SUM[21]) );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(n1), .CO(carry[7]), .S(SUM[6]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  AND2X2 U1 ( .A(B[5]), .B(A[5]), .Y(n1) );
  XOR2X1 U2 ( .A(B[5]), .B(A[5]), .Y(SUM[5]) );
  BUFX3 U3 ( .A(B[1]), .Y(SUM[1]) );
  BUFX3 U4 ( .A(B[2]), .Y(SUM[2]) );
  BUFX3 U5 ( .A(B[3]), .Y(SUM[3]) );
  BUFX3 U6 ( .A(B[4]), .Y(SUM[4]) );
endmodule


module idct8_shift7_add64_DW01_add_37 ( A, B, SUM );
  input [22:0] A;
  input [22:0] B;
  output [22:0] SUM;

  wire   [22:1] carry;

  XOR3X2 U1_22 ( .A(A[22]), .B(B[22]), .C(carry[22]), .Y(SUM[22]) );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(1'b0), .CO(carry[2]), .S(SUM[1]) );
  XOR2X1 U1 ( .A(1'b0), .B(A[0]), .Y(SUM[0]) );
endmodule


module idct8_shift7_add64_DW01_add_38 ( A, B, SUM );
  input [22:0] A;
  input [22:0] B;
  output [22:0] SUM;

  wire   [22:1] carry;

  XOR3X2 U1_22 ( .A(A[22]), .B(B[22]), .C(carry[22]), .Y(SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_1 ( .A(A[1]), .B(1'b0), .CI(1'b0), .S(SUM[1]) );
  ADDFX2 U1_2 ( .A(A[2]), .B(1'b0), .CI(1'b0), .S(SUM[2]) );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(1'b0), .CO(carry[4]), .S(SUM[3]) );
  XOR2X1 U1 ( .A(1'b0), .B(A[0]), .Y(SUM[0]) );
endmodule


module idct8_shift7_add64_DW01_add_39 ( A, B, SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n1;
  wire   [20:6] carry;

  XOR3X2 U1_20 ( .A(A[20]), .B(B[20]), .C(carry[20]), .Y(SUM[20]) );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(n1), .CO(carry[6]), .S(SUM[5]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  AND2X2 U1 ( .A(B[4]), .B(A[4]), .Y(n1) );
  XOR2X1 U2 ( .A(B[4]), .B(A[4]), .Y(SUM[4]) );
  BUFX3 U3 ( .A(B[1]), .Y(SUM[1]) );
  BUFX3 U4 ( .A(B[2]), .Y(SUM[2]) );
  BUFX3 U5 ( .A(B[3]), .Y(SUM[3]) );
endmodule


module idct8_shift7_add64_DW01_add_40 ( A, B, SUM );
  input [21:0] A;
  input [21:0] B;
  output [21:0] SUM;
  wire   n1;
  wire   [21:7] carry;

  XOR3X2 U1_21 ( .A(A[21]), .B(B[21]), .C(carry[21]), .Y(SUM[21]) );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(n1), .CO(carry[7]), .S(SUM[6]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  AND2X2 U1 ( .A(B[5]), .B(A[5]), .Y(n1) );
  XOR2X1 U2 ( .A(B[5]), .B(A[5]), .Y(SUM[5]) );
  BUFX3 U3 ( .A(B[1]), .Y(SUM[1]) );
  BUFX3 U4 ( .A(B[2]), .Y(SUM[2]) );
  BUFX3 U5 ( .A(B[3]), .Y(SUM[3]) );
  BUFX3 U6 ( .A(B[4]), .Y(SUM[4]) );
endmodule


module idct8_shift7_add64_DW01_add_41 ( A, B, SUM );
  input [22:0] A;
  input [22:0] B;
  output [22:0] SUM;

  wire   [22:1] carry;

  XOR3X2 U1_22 ( .A(A[22]), .B(B[22]), .C(carry[22]), .Y(SUM[22]) );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(1'b0), .CO(carry[2]), .S(SUM[1]) );
  XOR2X1 U1 ( .A(1'b0), .B(A[0]), .Y(SUM[0]) );
endmodule


module idct8_shift7_add64_DW01_add_42 ( A, B, SUM );
  input [22:0] A;
  input [22:0] B;
  output [22:0] SUM;

  wire   [22:1] carry;

  XOR3X2 U1_22 ( .A(A[22]), .B(B[22]), .C(carry[22]), .Y(SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_1 ( .A(A[1]), .B(1'b0), .CI(1'b0), .S(SUM[1]) );
  ADDFX2 U1_2 ( .A(A[2]), .B(1'b0), .CI(1'b0), .S(SUM[2]) );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(1'b0), .CO(carry[4]), .S(SUM[3]) );
  XOR2X1 U1 ( .A(1'b0), .B(A[0]), .Y(SUM[0]) );
endmodule


module idct8_shift7_add64_DW01_add_59 ( A, B, SUM );
  input [24:0] A;
  input [24:0] B;
  output [24:0] SUM;

  wire   [23:1] carry;

  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  XOR3X2 U1_23 ( .A(A[23]), .B(B[23]), .C(carry[23]), .Y(SUM[23]) );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(1'b0), .CO(carry[2]), .S(SUM[1]) );
  XOR2X1 U1 ( .A(B[0]), .B(1'b0), .Y(SUM[0]) );
endmodule


module idct8_shift7_add64_DW01_sub_0 ( B, DIFF );
  input [23:0] B;
  output [23:0] DIFF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46;

  AND2X2 U1 ( .A(n35), .B(n21), .Y(n1) );
  AND2X2 U2 ( .A(n34), .B(n1), .Y(n2) );
  AND2X2 U3 ( .A(n33), .B(n2), .Y(n3) );
  AND2X2 U4 ( .A(n32), .B(n3), .Y(n4) );
  AND2X2 U5 ( .A(n31), .B(n4), .Y(n5) );
  AND2X2 U6 ( .A(n30), .B(n5), .Y(n6) );
  AND2X2 U7 ( .A(n29), .B(n6), .Y(n7) );
  AND2X2 U8 ( .A(n28), .B(n7), .Y(n8) );
  AND2X2 U9 ( .A(n27), .B(n8), .Y(n9) );
  AND2X2 U10 ( .A(n26), .B(n9), .Y(n10) );
  AND2X2 U11 ( .A(n25), .B(n10), .Y(n11) );
  XOR2X1 U12 ( .A(n25), .B(n10), .Y(DIFF[21]) );
  XOR2X1 U13 ( .A(n24), .B(n11), .Y(DIFF[22]) );
  AND2X2 U14 ( .A(n45), .B(n46), .Y(n12) );
  AND2X2 U15 ( .A(n44), .B(n12), .Y(n13) );
  AND2X2 U16 ( .A(n43), .B(n13), .Y(n14) );
  AND2X2 U17 ( .A(n42), .B(n14), .Y(n15) );
  AND2X2 U18 ( .A(n41), .B(n15), .Y(n16) );
  AND2X2 U19 ( .A(n40), .B(n16), .Y(n17) );
  AND2X2 U20 ( .A(n39), .B(n17), .Y(n18) );
  AND2X2 U21 ( .A(n38), .B(n18), .Y(n19) );
  AND2X2 U22 ( .A(n37), .B(n19), .Y(n20) );
  AND2X2 U23 ( .A(n36), .B(n20), .Y(n21) );
  XOR2X1 U24 ( .A(n29), .B(n6), .Y(DIFF[17]) );
  XOR2X1 U25 ( .A(n28), .B(n7), .Y(DIFF[18]) );
  XOR2X1 U26 ( .A(n27), .B(n8), .Y(DIFF[19]) );
  XOR2X1 U27 ( .A(n26), .B(n9), .Y(DIFF[20]) );
  XOR2X1 U28 ( .A(n34), .B(n1), .Y(DIFF[12]) );
  XOR2X1 U29 ( .A(n33), .B(n2), .Y(DIFF[13]) );
  XOR2X1 U30 ( .A(n32), .B(n3), .Y(DIFF[14]) );
  XOR2X1 U31 ( .A(n31), .B(n4), .Y(DIFF[15]) );
  XOR2X1 U32 ( .A(n30), .B(n5), .Y(DIFF[16]) );
  XOR2X1 U33 ( .A(n38), .B(n18), .Y(DIFF[8]) );
  XOR2X1 U34 ( .A(n37), .B(n19), .Y(DIFF[9]) );
  XOR2X1 U35 ( .A(n36), .B(n20), .Y(DIFF[10]) );
  XOR2X1 U36 ( .A(n35), .B(n21), .Y(DIFF[11]) );
  XOR2X1 U37 ( .A(n43), .B(n13), .Y(DIFF[3]) );
  XOR2X1 U38 ( .A(n42), .B(n14), .Y(DIFF[4]) );
  XOR2X1 U39 ( .A(n41), .B(n15), .Y(DIFF[5]) );
  XOR2X1 U40 ( .A(n40), .B(n16), .Y(DIFF[6]) );
  XOR2X1 U41 ( .A(n39), .B(n17), .Y(DIFF[7]) );
  XOR2X1 U42 ( .A(n44), .B(n12), .Y(DIFF[2]) );
  XOR2X1 U43 ( .A(n45), .B(n46), .Y(DIFF[1]) );
  INVX1 U44 ( .A(B[11]), .Y(n35) );
  INVX1 U45 ( .A(B[12]), .Y(n34) );
  INVX1 U46 ( .A(B[13]), .Y(n33) );
  INVX1 U47 ( .A(B[14]), .Y(n32) );
  INVX1 U48 ( .A(B[15]), .Y(n31) );
  INVX1 U49 ( .A(B[16]), .Y(n30) );
  INVX1 U50 ( .A(B[17]), .Y(n29) );
  INVX1 U51 ( .A(B[18]), .Y(n28) );
  INVX1 U52 ( .A(B[19]), .Y(n27) );
  INVX1 U53 ( .A(B[20]), .Y(n26) );
  INVX1 U54 ( .A(B[21]), .Y(n25) );
  INVX1 U55 ( .A(B[22]), .Y(n24) );
  XOR2X1 U56 ( .A(B[23]), .B(n23), .Y(DIFF[23]) );
  NAND2X1 U57 ( .A(n24), .B(n11), .Y(n23) );
  INVX1 U58 ( .A(B[0]), .Y(n46) );
  INVX1 U59 ( .A(B[1]), .Y(n45) );
  INVX1 U60 ( .A(B[2]), .Y(n44) );
  INVX1 U61 ( .A(B[3]), .Y(n43) );
  INVX1 U62 ( .A(B[4]), .Y(n42) );
  INVX1 U63 ( .A(B[5]), .Y(n41) );
  INVX1 U64 ( .A(B[6]), .Y(n40) );
  INVX1 U65 ( .A(B[7]), .Y(n39) );
  INVX1 U66 ( .A(B[8]), .Y(n38) );
  INVX1 U67 ( .A(B[9]), .Y(n37) );
  INVX1 U68 ( .A(B[10]), .Y(n36) );
  BUFX3 U69 ( .A(B[0]), .Y(DIFF[0]) );
endmodule


module idct8_shift7_add64 ( clk, rstn, mode, start, x0, x1, x2, x3, x4, x5, x6, 
        x7, y0, y1, y2, y3, y4, y5, y6, y7, idct8_ready );
  input [1:0] mode;
  input [24:0] x0;
  input [24:0] x1;
  input [24:0] x2;
  input [24:0] x3;
  input [15:0] x4;
  input [15:0] x5;
  input [15:0] x6;
  input [15:0] x7;
  output [25:0] y0;
  output [25:0] y1;
  output [25:0] y2;
  output [25:0] y3;
  output [25:0] y4;
  output [25:0] y5;
  output [25:0] y6;
  output [25:0] y7;
  input clk, rstn, start;
  output idct8_ready;
  wire   N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36,
         N37, N38, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55,
         N56, N57, N58, N59, N60, N64, N65, N66, N67, N68, N69, N70, N71, N72,
         N73, N74, N75, N76, N77, N78, N79, N80, N85, N86, N87, N88, N89, N90,
         N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N108, N109,
         N110, N111, N112, N113, N114, N115, N116, N117, N118, N119, N120,
         N121, N122, N123, N129, N130, N131, N132, N133, N134, N135, N136,
         N137, N138, N139, N140, N141, N142, N143, N144, N145, N149, N150,
         N151, N152, N153, N154, N155, N156, N157, N158, N159, N160, N161,
         N162, N163, N164, N165, N170, N171, N172, N173, N174, N175, N176,
         N177, N178, N179, N180, N181, N182, N183, N184, N185, N186, N193,
         N194, N195, N196, N197, N198, N199, N200, N201, N202, N203, N204,
         N205, N206, N207, N208, N214, N215, N216, N217, N218, N219, N220,
         N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N234,
         N235, N236, N237, N238, N239, N240, N241, N242, N243, N244, N245,
         N246, N247, N248, N249, N250, N255, N256, N257, N258, N259, N260,
         N261, N262, N263, N264, N265, N266, N267, N268, N269, N270, N271,
         N278, N279, N280, N281, N282, N283, N284, N285, N286, N287, N288,
         N289, N290, N291, N292, N293, N299, N300, N301, N302, N303, N304,
         N305, N306, N307, N308, N309, N310, N311, N312, N313, N314, N315,
         N319, N320, N321, N322, N323, N324, N325, N326, N327, N328, N329,
         N330, N331, N332, N333, N334, N335, N340, N341, N342, N343, N344,
         N345, N346, N347, N348, N349, N350, N351, N352, N353, N354, N355,
         N356, N357, N358, N359, N360, N361, N362, N363, N364, N365, N366,
         N367, N368, N369, N370, N371, N372, N373, N374, N375, N376, N377,
         N378, N379, N380, N381, N382, N383, N384, N385, N386, N387, N388,
         N389, N390, N391, N392, N393, N394, N395, N396, N397, N398, N399,
         N400, N401, N402, N404, N405, N406, N407, N408, N409, N410, N411,
         N412, N413, N414, N415, N416, N417, N418, N419, N420, N421, N422,
         N423, N424, N426, N427, N428, N429, N430, N431, N432, N433, N434,
         N435, N436, N437, N438, N439, N440, N441, N442, N443, N444, N445,
         N446, N447, N448, N449, N450, N451, N452, N453, N454, N455, N456,
         N457, N458, N459, N460, N461, N462, N463, N464, N465, N466, N467,
         N468, N469, N470, N471, N472, N473, N474, N475, N476, N477, N478,
         N479, N480, N481, N482, N483, N484, N485, N486, N487, N488, N489,
         N490, N491, N493, N494, N495, N496, N497, N498, N499, N500, N501,
         N502, N503, N504, N505, N506, N507, N508, N509, N510, N511, N512,
         N513, N515, N516, N517, N518, N519, N520, N521, N522, N523, N524,
         N525, N526, N527, N528, N529, N530, N531, N532, N533, N534, N535,
         N536, N537, N538, N539, N540, N541, N542, N543, N544, N545, N546,
         N547, N548, N549, N550, N551, N552, N553, N554, N555, N556, N557,
         N558, N559, N560, N561, N562, N563, N564, N565, N566, N567, N568,
         N569, N570, N571, N572, N573, N574, N575, N576, N577, N578, N579,
         N580, N582, N583, N584, N585, N586, N587, N588, N589, N590, N591,
         N592, N593, N594, N595, N596, N597, N598, N599, N600, N601, N602,
         N604, N605, N606, N607, N608, N609, N610, N611, N612, N613, N614,
         N615, N616, N617, N618, N619, N620, N621, N622, N623, N624, N625,
         N626, N627, N628, N629, N630, N631, N632, N633, N634, N635, N636,
         N637, N638, N639, N640, N641, N642, N643, N644, N645, N646, N647,
         N648, N649, N650, N651, N652, N653, N654, N655, N656, N657, N658,
         N659, N660, N661, N662, N663, N664, N665, N666, N667, N668, N669,
         N671, N672, N673, N674, N675, N676, N677, N678, N679, N680, N681,
         N682, N683, N684, N685, N686, N687, N688, N689, N690, N691, N693,
         N694, N695, N696, N697, N698, N699, N700, N701, N702, N703, N704,
         N705, N706, N707, N708, N709, N710, N711, N712, N760, N761, N762,
         N763, N764, N765, N766, N767, N768, N769, N770, N771, N772, N773,
         N774, N775, N776, N777, N778, N779, N780, N781, N782, N783, N830,
         N831, N832, N833, N834, N835, N836, N837, N838, N839, N840, N841,
         N842, N843, N844, N845, N846, N847, N848, N849, N850, N851, N852,
         N853, N854, N855, N856, N857, N858, N859, N860, N861, N862, N863,
         N864, N865, N866, N867, N868, N869, N870, N871, N872, N873, N874,
         N875, N876, N877, N878, N879, N880, N881, N882, N883, N884, N885,
         N886, N887, N888, N889, N890, N891, N892, N893, N894, N895, N896,
         N897, N898, N899, N900, N901, N902, N950, N951, N952, N953, N954,
         N955, N956, N957, N958, N959, N960, N961, N962, N963, N964, N965,
         N966, N967, N968, N969, N970, N971, N972, N973, N974, N975, N976,
         N977, N978, N979, N980, N981, N982, N983, N984, N985, N986, N987,
         N988, N989, N990, N991, N992, N993, N994, N995, N996, N997, N998,
         N1045, N1046, N1047, N1048, N1049, N1050, N1051, N1052, N1053, N1054,
         N1055, N1056, N1057, N1058, N1059, N1060, N1061, N1062, N1063, N1064,
         N1065, N1066, N1067, N1068, N1093, N1094, N1095, N1096, N1097, N1098,
         N1099, N1100, N1101, N1102, N1103, N1104, N1105, N1106, N1107, N1108,
         N1109, N1110, N1111, N1112, N1113, N1114, N1115, N1116, N1117, N1118,
         N1119, N1120, N1121, N1122, N1123, N1124, N1125, N1126, N1127, N1128,
         N1129, N1130, N1131, N1132, N1133, N1134, N1135, N1136, N1137, N1138,
         N1139, N1140, N1141, N1142, N1143, N1144, N1145, N1146, N1147, N1148,
         N1149, N1150, N1151, N1152, N1153, N1154, N1155, N1156, N1157, N1158,
         N1159, N1160, N1161, N1162, N1163, N1164, N1165, N1166, N1167, N1168,
         N1169, N1170, N1171, N1172, N1173, N1174, N1175, N1176, N1177, N1178,
         N1179, N1180, N1181, N1182, N1183, N1184, N1185, N1186, N1187, N1188,
         N1189, N1190, N1191, N1192, N1193, N1194, N1195, N1196, N1197, N1198,
         N1199, N1200, N1201, N1202, N1203, N1204, N1205, N1206, N1207, N1208,
         N1209, N1210, N1211, N1212, N1213, N1214, N1215, N1216, N1217, N1218,
         N1219, N1220, N1221, N1222, N1223, N1224, N1225, N1226, N1227, N1228,
         N1229, N1230, N1231, N1232, N1233, N1234, N1235, N1236, N1237, N1238,
         N1239, N1240, N1241, N1242, N1243, N1244, N1245, N1246, N1247, N1248,
         N1249, N1250, N1251, N1252, N1253, N1254, N1255, N1256, N1257, N1258,
         N1259, N1260, N1261, N1262, N1263, N1264, N1265, N1266, N1267, N1268,
         N1269, N1270, N1271, N1272, N1273, N1274, N1275, N1276, N1277, N1278,
         N1279, N1280, N1281, N1282, N1283, N1284, N1285, N1286, N1287, N1288,
         N1289, N1290, N1291, N1292, N1293, N1294, N1295, N1296, N1297, N1298,
         N1299, N1300, N1301, N1302, N1303, N1304, N1305, N1306, N1307, N1308,
         N1309, N1310, N1311, N1312, N1313, N1314, N1315, N1316, N1317, N1318,
         N1370, N1371, N1372, N1373, N1374, N1375, N1376, N1377, N1378, N1379,
         N1380, N1381, N1382, N1383, N1384, N1385, N1386, N1387, N1388, N1389,
         N1390, N1391, N1392, N1393, N1394, N1395, N1447, N1448, N1449, N1450,
         N1451, N1452, N1453, N1454, N1455, N1456, N1457, N1458, N1459, N1460,
         N1461, N1462, N1463, N1464, N1465, N1466, N1467, N1468, N1469, N1470,
         N1471, N1472, N1524, N1525, N1526, N1527, N1528, N1529, N1530, N1531,
         N1532, N1533, N1534, N1535, N1536, N1537, N1538, N1539, N1540, N1541,
         N1542, N1543, N1544, N1545, N1546, N1547, N1548, N1549, N1601, N1602,
         N1603, N1604, N1605, N1606, N1607, N1608, N1609, N1610, N1611, N1612,
         N1613, N1614, N1615, N1616, N1617, N1618, N1619, N1620, N1621, N1622,
         N1623, N1624, N1625, N1626, N1627, N1628, N1629, N1630, N1631, N1632,
         N1633, N1634, N1635, N1636, N1637, N1638, N1639, N1640, N1641, N1642,
         N1643, N1644, N1645, N1646, N1647, N1648, N1649, N1650, N1651, N1652,
         N1653, N1654, N1655, N1656, N1657, N1658, N1659, N1660, N1661, N1662,
         N1663, N1664, N1665, N1666, N1667, N1668, N1669, N1670, N1671, N1672,
         N1673, N1674, N1675, N1676, N1677, N1678, N1679, N1680, N1681, N1682,
         N1683, N1684, N1685, N1686, N1687, N1688, N1689, N1690, N1691, N1692,
         N1693, N1694, N1695, N1696, N1697, N1698, N1699, N1700, N1701, N1702,
         N1703, N1704, N1705, N1706, N1707, N1708, N1709, N1710, N1711, N1712,
         N1713, N1714, N1715, N1716, N1717, N1718, N1719, N1720, N1721, N1722,
         N1723, N1724, N1725, N1726, N1727, N1728, N1729, N1730, N1731, N1732,
         N1733, N1734, N1735, N1736, N1737, N1738, N1739, N1740, N1741, N1742,
         N1743, N1744, N1745, N1746, N1747, N1748, N1749, N1750, N1751, N1752,
         N1753, N1754, N1755, N1756, N1757, N1758, N1759, N1760, N1761, N1762,
         N1763, N1764, N1765, N1766, N1767, N1768, N1769, N1770, N1771, N1772,
         N1773, N1774, N1775, N1776, N1777, N1778, N1779, N1780, N1781, N1782,
         N1783, N1784, N1785, N1786, N1787, N1788, N1789, N1790, N1791, N1792,
         N1793, N1794, N1795, N1796, N1797, N1798, N1799, N1800, N1801, N1802,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, N1092, N1091, N1090, N1089, N1088, N1087, N1086, N1085, N1084,
         N1083, N1082, N1081, N1080, N1079, N1078, N1077, N1076, N1075, N1074,
         N1073, N1072, N1071, N1070, N1069, add_104_carry_10_,
         add_104_carry_11_, add_104_carry_12_, add_104_carry_13_,
         add_104_carry_14_, add_104_carry_15_, add_104_carry_16_,
         add_104_carry_17_, add_104_carry_18_, add_104_carry_5_,
         add_104_carry_6_, add_104_carry_7_, add_104_carry_8_,
         add_104_carry_9_, add_102_carry_10_, add_102_carry_11_,
         add_102_carry_12_, add_102_carry_13_, add_102_carry_14_,
         add_102_carry_15_, add_102_carry_16_, add_102_carry_17_,
         add_102_carry_4_, add_102_carry_5_, add_102_carry_6_,
         add_102_carry_7_, add_102_carry_8_, add_102_carry_9_,
         add_100_carry_10_, add_100_carry_11_, add_100_carry_12_,
         add_100_carry_13_, add_100_carry_14_, add_100_carry_15_,
         add_100_carry_16_, add_100_carry_17_, add_100_carry_18_,
         add_100_carry_5_, add_100_carry_6_, add_100_carry_7_,
         add_100_carry_8_, add_100_carry_9_, add_99_carry_10_,
         add_99_carry_11_, add_99_carry_12_, add_99_carry_13_,
         add_99_carry_14_, add_99_carry_15_, add_99_carry_16_,
         add_99_carry_17_, add_99_carry_18_, add_99_carry_19_,
         add_99_carry_20_, add_99_carry_7_, add_99_carry_8_, add_99_carry_9_,
         add_95_carry_10_, add_95_carry_11_, add_95_carry_12_,
         add_95_carry_13_, add_95_carry_14_, add_95_carry_15_,
         add_95_carry_16_, add_95_carry_17_, add_95_carry_18_, add_95_carry_5_,
         add_95_carry_6_, add_95_carry_7_, add_95_carry_8_, add_95_carry_9_,
         add_93_carry_10_, add_93_carry_11_, add_93_carry_12_,
         add_93_carry_13_, add_93_carry_14_, add_93_carry_15_,
         add_93_carry_16_, add_93_carry_17_, add_93_carry_4_, add_93_carry_5_,
         add_93_carry_6_, add_93_carry_7_, add_93_carry_8_, add_93_carry_9_,
         add_91_carry_10_, add_91_carry_11_, add_91_carry_12_,
         add_91_carry_13_, add_91_carry_14_, add_91_carry_15_,
         add_91_carry_16_, add_91_carry_17_, add_91_carry_18_, add_91_carry_5_,
         add_91_carry_6_, add_91_carry_7_, add_91_carry_8_, add_91_carry_9_,
         add_90_carry_10_, add_90_carry_11_, add_90_carry_12_,
         add_90_carry_13_, add_90_carry_14_, add_90_carry_15_,
         add_90_carry_16_, add_90_carry_17_, add_90_carry_18_,
         add_90_carry_19_, add_90_carry_20_, add_90_carry_7_, add_90_carry_8_,
         add_90_carry_9_, add_86_carry_10_, add_86_carry_11_, add_86_carry_12_,
         add_86_carry_13_, add_86_carry_14_, add_86_carry_15_,
         add_86_carry_16_, add_86_carry_17_, add_86_carry_18_, add_86_carry_5_,
         add_86_carry_6_, add_86_carry_7_, add_86_carry_8_, add_86_carry_9_,
         add_84_carry_10_, add_84_carry_11_, add_84_carry_12_,
         add_84_carry_13_, add_84_carry_14_, add_84_carry_15_,
         add_84_carry_16_, add_84_carry_17_, add_84_carry_4_, add_84_carry_5_,
         add_84_carry_6_, add_84_carry_7_, add_84_carry_8_, add_84_carry_9_,
         add_82_carry_10_, add_82_carry_11_, add_82_carry_12_,
         add_82_carry_13_, add_82_carry_14_, add_82_carry_15_,
         add_82_carry_16_, add_82_carry_17_, add_82_carry_18_, add_82_carry_5_,
         add_82_carry_6_, add_82_carry_7_, add_82_carry_8_, add_82_carry_9_,
         add_81_carry_10_, add_81_carry_11_, add_81_carry_12_,
         add_81_carry_13_, add_81_carry_14_, add_81_carry_15_,
         add_81_carry_16_, add_81_carry_17_, add_81_carry_18_,
         add_81_carry_19_, add_81_carry_20_, add_81_carry_7_, add_81_carry_8_,
         add_81_carry_9_, add_77_carry_10_, add_77_carry_11_, add_77_carry_12_,
         add_77_carry_13_, add_77_carry_14_, add_77_carry_15_,
         add_77_carry_16_, add_77_carry_17_, add_77_carry_18_, add_77_carry_5_,
         add_77_carry_6_, add_77_carry_7_, add_77_carry_8_, add_77_carry_9_,
         add_75_carry_10_, add_75_carry_11_, add_75_carry_12_,
         add_75_carry_13_, add_75_carry_14_, add_75_carry_15_,
         add_75_carry_16_, add_75_carry_17_, add_75_carry_4_, add_75_carry_5_,
         add_75_carry_6_, add_75_carry_7_, add_75_carry_8_, add_75_carry_9_,
         add_73_carry_10_, add_73_carry_11_, add_73_carry_12_,
         add_73_carry_13_, add_73_carry_14_, add_73_carry_15_,
         add_73_carry_16_, add_73_carry_17_, add_73_carry_18_, add_73_carry_5_,
         add_73_carry_6_, add_73_carry_7_, add_73_carry_8_, add_73_carry_9_,
         add_72_carry_10_, add_72_carry_11_, add_72_carry_12_,
         add_72_carry_13_, add_72_carry_14_, add_72_carry_15_,
         add_72_carry_16_, add_72_carry_17_, add_72_carry_18_,
         add_72_carry_19_, add_72_carry_20_, add_72_carry_7_, add_72_carry_8_,
         add_72_carry_9_, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n590, n591, n592;
  wire   [1:0] mode_delay2;
  wire   [1:0] mode_delay1;
  wire   [20:0] x4_89_tmp2;
  wire   [19:0] x4_75_tmp2;
  wire   [20:0] x4_50_tmp1;
  wire   [20:0] x4_50_tmp2;
  wire   [19:0] x4_18_tmp1;
  wire   [16:0] x4_18_tmp2;
  wire   [20:0] x5_89_tmp2;
  wire   [19:0] x5_75_tmp2;
  wire   [20:0] x5_50_tmp1;
  wire   [20:0] x5_50_tmp2;
  wire   [19:0] x5_18_tmp1;
  wire   [16:0] x5_18_tmp2;
  wire   [20:0] x6_89_tmp2;
  wire   [19:0] x6_75_tmp2;
  wire   [20:0] x6_50_tmp1;
  wire   [20:0] x6_50_tmp2;
  wire   [19:0] x6_18_tmp1;
  wire   [16:0] x6_18_tmp2;
  wire   [20:0] x7_89_tmp2;
  wire   [19:0] x7_75_tmp2;
  wire   [20:0] x7_50_tmp1;
  wire   [20:0] x7_50_tmp2;
  wire   [19:0] x7_18_tmp1;
  wire   [16:0] x7_18_tmp2;
  wire   [22:0] x4_89;
  wire   [22:0] x5_89;
  wire   [22:0] x6_89;
  wire   [22:0] x7_89;
  wire   [22:0] x4_75;
  wire   [22:0] x5_75;
  wire   [22:0] x6_75;
  wire   [22:0] x7_75;
  wire   [21:0] x4_50;
  wire   [21:0] x5_50;
  wire   [21:0] x6_50;
  wire   [21:0] x7_50;
  wire   [20:0] x4_18;
  wire   [20:0] x5_18;
  wire   [20:0] x6_18;
  wire   [20:0] x7_18;
  wire   [22:0] x7_75_tmp1;
  wire   [22:0] x6_75_tmp1;
  wire   [22:0] x5_75_tmp1;
  wire   [22:0] x4_75_tmp1;
  wire   [22:0] x7_89_tmp1;
  wire   [22:0] x6_89_tmp1;
  wire   [22:0] x5_89_tmp1;
  wire   [22:0] x4_89_tmp1;
  wire   [23:0] x4_tmp1;
  wire   [23:0] x4_tmp2;
  wire   [23:0] x5_tmp1;
  wire   [23:0] x5_tmp2;
  wire   [23:0] x6_tmp1;
  wire   [23:0] x6_tmp2;
  wire   [23:0] x7_tmp1;
  wire   [23:0] x7_tmp2;
  wire   [24:0] x4_tmp;
  wire   [24:0] x5_tmp;
  wire   [24:0] x6_tmp;
  wire   [24:0] x7_tmp;
  wire   [25:0] y0_tmp;
  wire   [25:0] y1_tmp;
  wire   [25:0] y2_tmp;
  wire   [25:0] y3_tmp;
  wire   [25:0] y4_tmp;
  wire   [25:0] y5_tmp;
  wire   [25:0] y6_tmp;
  wire   [25:0] y7_tmp;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64;

  idct8_shift7_add64_DW01_add_0 add_187 ( .A({1'b0, y7_tmp[25], y7_tmp[25], 
        y7_tmp}), .SUM({N1802, N1801, N1800, N1799, N1798, N1797, N1796, N1795, 
        N1794, N1793, N1792, N1791, N1790, N1789, N1788, N1787, N1786, N1785, 
        N1784, N1783, N1782, N1781, SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6}) );
  idct8_shift7_add64_DW01_add_1 add_186 ( .A({1'b0, y6_tmp[25], y6_tmp[25], 
        y6_tmp}), .SUM({N1780, N1779, N1778, N1777, N1776, N1775, N1774, N1773, 
        N1772, N1771, N1770, N1769, N1768, N1767, N1766, N1765, N1764, N1763, 
        N1762, N1761, N1760, N1759, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13}) );
  idct8_shift7_add64_DW01_add_2 add_185 ( .A({1'b0, y5_tmp[25], y5_tmp[25], 
        y5_tmp}), .SUM({N1758, N1757, N1756, N1755, N1754, N1753, N1752, N1751, 
        N1750, N1749, N1748, N1747, N1746, N1745, N1744, N1743, N1742, N1741, 
        N1740, N1739, N1738, N1737, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, SYNOPSYS_UNCONNECTED__16, 
        SYNOPSYS_UNCONNECTED__17, SYNOPSYS_UNCONNECTED__18, 
        SYNOPSYS_UNCONNECTED__19, SYNOPSYS_UNCONNECTED__20}) );
  idct8_shift7_add64_DW01_add_3 add_184 ( .A({1'b0, y4_tmp[25], y4_tmp[25], 
        y4_tmp}), .SUM({N1736, N1735, N1734, N1733, N1732, N1731, N1730, N1729, 
        N1728, N1727, N1726, N1725, N1724, N1723, N1722, N1721, N1720, N1719, 
        N1718, N1717, N1716, N1715, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27}) );
  idct8_shift7_add64_DW01_add_4 add_183 ( .A({1'b0, y3_tmp[25], y3_tmp[25], 
        y3_tmp}), .SUM({N1714, N1713, N1712, N1711, N1710, N1709, N1708, N1707, 
        N1706, N1705, N1704, N1703, N1702, N1701, N1700, N1699, N1698, N1697, 
        N1696, N1695, N1694, N1693, SYNOPSYS_UNCONNECTED__28, 
        SYNOPSYS_UNCONNECTED__29, SYNOPSYS_UNCONNECTED__30, 
        SYNOPSYS_UNCONNECTED__31, SYNOPSYS_UNCONNECTED__32, 
        SYNOPSYS_UNCONNECTED__33, SYNOPSYS_UNCONNECTED__34}) );
  idct8_shift7_add64_DW01_add_5 add_182 ( .A({1'b0, y2_tmp[25], y2_tmp[25], 
        y2_tmp}), .SUM({N1692, N1691, N1690, N1689, N1688, N1687, N1686, N1685, 
        N1684, N1683, N1682, N1681, N1680, N1679, N1678, N1677, N1676, N1675, 
        N1674, N1673, N1672, N1671, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41}) );
  idct8_shift7_add64_DW01_add_6 add_181 ( .A({1'b0, y1_tmp[25], y1_tmp[25], 
        y1_tmp}), .SUM({N1670, N1669, N1668, N1667, N1666, N1665, N1664, N1663, 
        N1662, N1661, N1660, N1659, N1658, N1657, N1656, N1655, N1654, N1653, 
        N1652, N1651, N1650, N1649, SYNOPSYS_UNCONNECTED__42, 
        SYNOPSYS_UNCONNECTED__43, SYNOPSYS_UNCONNECTED__44, 
        SYNOPSYS_UNCONNECTED__45, SYNOPSYS_UNCONNECTED__46, 
        SYNOPSYS_UNCONNECTED__47, SYNOPSYS_UNCONNECTED__48}) );
  idct8_shift7_add64_DW01_add_7 add_180 ( .A({1'b0, y0_tmp[25], y0_tmp[25], 
        y0_tmp}), .SUM({N1648, N1647, N1646, N1645, N1644, N1643, N1642, N1641, 
        N1640, N1639, N1638, N1637, N1636, N1635, N1634, N1633, N1632, N1631, 
        N1630, N1629, N1628, N1627, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55}) );
  idct8_shift7_add64_DW01_add_8 add_1_root_add_177_2 ( .A({x0[24], x0}), .B({
        n340, n340, n339, n338, n337, n336, n335, n334, n333, n332, n331, n330, 
        n329, n328, n327, n326, n325, n324, n323, n322, n321, n320, n319, n318, 
        n317, n316}), .SUM({N1626, N1625, N1624, N1623, N1622, N1621, N1620, 
        N1619, N1618, N1617, N1616, N1615, N1614, N1613, N1612, N1611, N1610, 
        N1609, N1608, N1607, N1606, N1605, N1604, N1603, N1602, N1601}) );
  idct8_shift7_add64_DW01_add_9 add_1_root_add_176_2 ( .A({x1[24], x1}), .B({
        n366, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, 
        n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, 
        n389, n390}), .SUM({N1549, N1548, N1547, N1546, N1545, N1544, N1543, 
        N1542, N1541, N1540, N1539, N1538, N1537, N1536, N1535, N1534, N1533, 
        N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524}) );
  idct8_shift7_add64_DW01_add_10 add_1_root_add_175_2 ( .A({x2[24], x2}), .B({
        n341, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, 
        n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, 
        n364, n365}), .SUM({N1472, N1471, N1470, N1469, N1468, N1467, N1466, 
        N1465, N1464, N1463, N1462, N1461, N1460, N1459, N1458, N1457, N1456, 
        N1455, N1454, N1453, N1452, N1451, N1450, N1449, N1448, N1447}) );
  idct8_shift7_add64_DW01_add_11 add_1_root_add_174_2 ( .A({x3[24], x3}), .B({
        n592, n592, n591, n590, n412, n411, n410, n409, n408, n407, n406, n405, 
        n404, n403, n402, n401, n400, n399, n398, n397, n396, n395, n394, n393, 
        n392, n391}), .SUM({N1395, N1394, N1393, N1392, N1391, N1390, N1389, 
        N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, 
        N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370}) );
  idct8_shift7_add64_DW01_add_12 add_173 ( .A({x3[24], x3}), .B({x4_tmp[24], 
        x4_tmp}), .SUM({N1318, N1317, N1316, N1315, N1314, N1313, N1312, N1311, 
        N1310, N1309, N1308, N1307, N1306, N1305, N1304, N1303, N1302, N1301, 
        N1300, N1299, N1298, N1297, N1296, N1295, N1294, N1293}) );
  idct8_shift7_add64_DW01_add_13 add_172 ( .A({x2[24], x2}), .B({x5_tmp[24], 
        x5_tmp}), .SUM({N1292, N1291, N1290, N1289, N1288, N1287, N1286, N1285, 
        N1284, N1283, N1282, N1281, N1280, N1279, N1278, N1277, N1276, N1275, 
        N1274, N1273, N1272, N1271, N1270, N1269, N1268, N1267}) );
  idct8_shift7_add64_DW01_add_14 add_171 ( .A({x1[24], x1}), .B({x6_tmp[24], 
        x6_tmp}), .SUM({N1266, N1265, N1264, N1263, N1262, N1261, N1260, N1259, 
        N1258, N1257, N1256, N1255, N1254, N1253, N1252, N1251, N1250, N1249, 
        N1248, N1247, N1246, N1245, N1244, N1243, N1242, N1241}) );
  idct8_shift7_add64_DW01_add_15 add_170 ( .A({x0[24], x0}), .B({x7_tmp[24], 
        x7_tmp}), .SUM({N1240, N1239, N1238, N1237, N1236, N1235, N1234, N1233, 
        N1232, N1231, N1230, N1229, N1228, N1227, N1226, N1225, N1224, N1223, 
        N1222, N1221, N1220, N1219, N1218, N1217, N1216, N1215}) );
  idct8_shift7_add64_DW01_add_16 add_157 ( .A({x7_tmp1[23], x7_tmp1}), .B({
        x7_tmp2[23], x7_tmp2}), .SUM({N1214, N1213, N1212, N1211, N1210, N1209, 
        N1208, N1207, N1206, N1205, N1204, N1203, N1202, N1201, N1200, N1199, 
        N1198, N1197, N1196, N1195, N1194, N1193, N1192, N1191, N1190}) );
  idct8_shift7_add64_DW01_add_17 add_156 ( .A({x5_75[22], x5_75}), .B({
        x6_50[21], x6_50[21], x6_50}), .SUM({N1189, N1188, N1187, N1186, N1185, 
        N1184, N1183, N1182, N1181, N1180, N1179, N1178, N1177, N1176, N1175, 
        N1174, N1173, N1172, N1171, N1170, N1169, N1168, N1167, N1166}) );
  idct8_shift7_add64_DW01_add_18 add_155 ( .A({x4_89[22], x4_89}), .B({
        x7_18[20], x7_18[20], x7_18[20], x7_18[20:1], 1'b0}), .SUM({N1165, 
        N1164, N1163, N1162, N1161, N1160, N1159, N1158, N1157, N1156, N1155, 
        N1154, N1153, N1152, N1151, N1150, N1149, N1148, N1147, N1146, N1145, 
        N1144, N1143, N1142}) );
  idct8_shift7_add64_DW01_add_19 add_153 ( .A({x6_tmp1[23], x6_tmp1}), .B({
        x6_tmp2[23], x6_tmp2}), .SUM({N1141, N1140, N1139, N1138, N1137, N1136, 
        N1135, N1134, N1133, N1132, N1131, N1130, N1129, N1128, N1127, N1126, 
        N1125, N1124, N1123, N1122, N1121, N1120, N1119, N1118, N1117}) );
  idct8_shift7_add64_DW01_add_20 add_1_root_add_151_2 ( .A({x4_75[22], x4_75}), 
        .B({n226, n226, n226, n227, n228, n229, n230, n231, n232, n233, n234, 
        n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, 
        n247}), .SUM({N1068, N1067, N1066, N1065, N1064, N1063, N1062, N1061, 
        N1060, N1059, N1058, N1057, N1056, N1055, N1054, N1053, N1052, N1051, 
        N1050, N1049, N1048, N1047, N1046, N1045}) );
  idct8_shift7_add64_DW01_add_21 add_149 ( .A({x5_tmp1[23], x5_tmp1}), .B({
        x5_tmp2[23], x5_tmp2}), .SUM({N998, N997, N996, N995, N994, N993, N992, 
        N991, N990, N989, N988, N987, N986, N985, N984, N983, N982, N981, N980, 
        N979, N978, N977, N976, N975, N974}) );
  idct8_shift7_add64_DW01_add_22 add_1_root_add_148_2 ( .A({x6_18[20], 
        x6_18[20], x6_18[20], x6_18[20:1], 1'b0}), .B({n248, n248, n249, n250, 
        n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, 
        n263, n264, n265, n266, n267, n268, n269, n270}), .SUM({N973, N972, 
        N971, N970, N969, N968, N967, N966, N965, N964, N963, N962, N961, N960, 
        N959, N958, N957, N956, N955, N954, N953, N952, N951, N950}) );
  idct8_shift7_add64_DW01_add_23 add_147 ( .A({x4_50[21], x4_50[21], x4_50}), 
        .B({x7_75[22], x7_75}), .SUM({N902, N901, N900, N899, N898, N897, N896, 
        N895, N894, N893, N892, N891, N890, N889, N888, N887, N886, N885, N884, 
        N883, N882, N881, N880, N879}) );
  idct8_shift7_add64_DW01_add_24 add_145 ( .A({x4_tmp1[23], x4_tmp1}), .B({
        x4_tmp2[23], x4_tmp2}), .SUM({N878, N877, N876, N875, N874, N873, N872, 
        N871, N870, N869, N868, N867, N866, N865, N864, N863, N862, N861, N860, 
        N859, N858, N857, N856, N855, N854}) );
  idct8_shift7_add64_DW01_add_25 add_1_root_add_144_2 ( .A({x6_75[22], x6_75}), 
        .B({n294, n294, n294, n295, n296, n297, n298, n299, n300, n301, n302, 
        n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, 
        n315}), .SUM({N853, N852, N851, N850, N849, N848, N847, N846, N845, 
        N844, N843, N842, N841, N840, N839, N838, N837, N836, N835, N834, N833, 
        N832, N831, N830}) );
  idct8_shift7_add64_DW01_add_26 add_1_root_add_143_2 ( .A({x4_18[20], 
        x4_18[20], x4_18[20], x4_18[20:1], 1'b0}), .B({n271, n271, n272, n273, 
        n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, 
        n286, n287, n288, n289, n290, n291, n292, n293}), .SUM({N783, N782, 
        N781, N780, N779, N778, N777, N776, N775, N774, N773, N772, N771, N770, 
        N769, N768, N767, N766, N765, N764, N763, N762, N761, N760}) );
  idct8_shift7_add64_DW01_add_27 add_127 ( .A({x7_18_tmp1[19], 
        x7_18_tmp1[19:4], 1'b0, 1'b0, 1'b0, 1'b0}), .B({x7_18_tmp2[16], 
        x7_18_tmp2[16], x7_18_tmp2[16], x7_18_tmp2[16], x7_18_tmp2[16:1], 1'b0}), .SUM({N712, N711, N710, N709, N708, N707, N706, N705, N704, N703, N702, 
        N701, N700, N699, N698, N697, N696, N695, N694, N693, 
        SYNOPSYS_UNCONNECTED__56}) );
  idct8_shift7_add64_DW01_add_28 add_126 ( .A({x7_50_tmp1[20], 
        x7_50_tmp1[20:5], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({x7_50_tmp2[20], 
        x7_50_tmp2[20:1], 1'b0}), .SUM({N691, N690, N689, N688, N687, N686, 
        N685, N684, N683, N682, N681, N680, N679, N678, N677, N676, N675, N674, 
        N673, N672, N671, SYNOPSYS_UNCONNECTED__57}) );
  idct8_shift7_add64_DW01_add_29 add_125 ( .A(x7_75_tmp1), .B({x7_75_tmp2[19], 
        x7_75_tmp2[19], x7_75_tmp2[19], x7_75_tmp2[19:1], 1'b0}), .SUM({N669, 
        N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, 
        N656, N655, N654, N653, N652, N651, N650, N649, N648, N647}) );
  idct8_shift7_add64_DW01_add_30 add_124 ( .A(x7_89_tmp1), .B({x7_89_tmp2[20], 
        x7_89_tmp2[20], x7_89_tmp2[20:3], 1'b0, 1'b0, 1'b0}), .SUM({N646, N645, 
        N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, 
        N632, N631, N630, N629, N628, N627, N626, N625, N624}) );
  idct8_shift7_add64_DW01_add_31 add_122 ( .A({x6_18_tmp1[19], 
        x6_18_tmp1[19:4], 1'b0, 1'b0, 1'b0, 1'b0}), .B({x6_18_tmp2[16], 
        x6_18_tmp2[16], x6_18_tmp2[16], x6_18_tmp2[16], x6_18_tmp2[16:1], 1'b0}), .SUM({N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, 
        N612, N611, N610, N609, N608, N607, N606, N605, N604, 
        SYNOPSYS_UNCONNECTED__58}) );
  idct8_shift7_add64_DW01_add_32 add_121 ( .A({x6_50_tmp1[20], 
        x6_50_tmp1[20:5], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({x6_50_tmp2[20], 
        x6_50_tmp2[20:1], 1'b0}), .SUM({N602, N601, N600, N599, N598, N597, 
        N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, 
        N584, N583, N582, SYNOPSYS_UNCONNECTED__59}) );
  idct8_shift7_add64_DW01_add_33 add_120 ( .A(x6_75_tmp1), .B({x6_75_tmp2[19], 
        x6_75_tmp2[19], x6_75_tmp2[19], x6_75_tmp2[19:1], 1'b0}), .SUM({N580, 
        N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, 
        N567, N566, N565, N564, N563, N562, N561, N560, N559, N558}) );
  idct8_shift7_add64_DW01_add_34 add_119 ( .A(x6_89_tmp1), .B({x6_89_tmp2[20], 
        x6_89_tmp2[20], x6_89_tmp2[20:3], 1'b0, 1'b0, 1'b0}), .SUM({N557, N556, 
        N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, 
        N543, N542, N541, N540, N539, N538, N537, N536, N535}) );
  idct8_shift7_add64_DW01_add_35 add_117 ( .A({x5_18_tmp1[19], 
        x5_18_tmp1[19:4], 1'b0, 1'b0, 1'b0, 1'b0}), .B({x5_18_tmp2[16], 
        x5_18_tmp2[16], x5_18_tmp2[16], x5_18_tmp2[16], x5_18_tmp2[16:1], 1'b0}), .SUM({N534, N533, N532, N531, N530, N529, N528, N527, N526, N525, N524, 
        N523, N522, N521, N520, N519, N518, N517, N516, N515, 
        SYNOPSYS_UNCONNECTED__60}) );
  idct8_shift7_add64_DW01_add_36 add_116 ( .A({x5_50_tmp1[20], 
        x5_50_tmp1[20:5], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({x5_50_tmp2[20], 
        x5_50_tmp2[20:1], 1'b0}), .SUM({N513, N512, N511, N510, N509, N508, 
        N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, 
        N495, N494, N493, SYNOPSYS_UNCONNECTED__61}) );
  idct8_shift7_add64_DW01_add_37 add_115 ( .A(x5_75_tmp1), .B({x5_75_tmp2[19], 
        x5_75_tmp2[19], x5_75_tmp2[19], x5_75_tmp2[19:1], 1'b0}), .SUM({N491, 
        N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, 
        N478, N477, N476, N475, N474, N473, N472, N471, N470, N469}) );
  idct8_shift7_add64_DW01_add_38 add_114 ( .A(x5_89_tmp1), .B({x5_89_tmp2[20], 
        x5_89_tmp2[20], x5_89_tmp2[20:3], 1'b0, 1'b0, 1'b0}), .SUM({N468, N467, 
        N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, 
        N454, N453, N452, N451, N450, N449, N448, N447, N446}) );
  idct8_shift7_add64_DW01_add_39 add_112 ( .A({x4_18_tmp1[19], 
        x4_18_tmp1[19:4], 1'b0, 1'b0, 1'b0, 1'b0}), .B({x4_18_tmp2[16], 
        x4_18_tmp2[16], x4_18_tmp2[16], x4_18_tmp2[16], x4_18_tmp2[16:1], 1'b0}), .SUM({N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, 
        N434, N433, N432, N431, N430, N429, N428, N427, N426, 
        SYNOPSYS_UNCONNECTED__62}) );
  idct8_shift7_add64_DW01_add_40 add_111 ( .A({x4_50_tmp1[20], 
        x4_50_tmp1[20:5], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({x4_50_tmp2[20], 
        x4_50_tmp2[20:1], 1'b0}), .SUM({N424, N423, N422, N421, N420, N419, 
        N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, 
        N406, N405, N404, SYNOPSYS_UNCONNECTED__63}) );
  idct8_shift7_add64_DW01_add_41 add_110 ( .A(x4_75_tmp1), .B({x4_75_tmp2[19], 
        x4_75_tmp2[19], x4_75_tmp2[19], x4_75_tmp2[19:1], 1'b0}), .SUM({N402, 
        N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, 
        N389, N388, N387, N386, N385, N384, N383, N382, N381, N380}) );
  idct8_shift7_add64_DW01_add_42 add_109 ( .A(x4_89_tmp1), .B({x4_89_tmp2[20], 
        x4_89_tmp2[20], x4_89_tmp2[20:3], 1'b0, 1'b0, 1'b0}), .SUM({N379, N378, 
        N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, 
        N365, N364, N363, N362, N361, N360, N359, N358, N357}) );
  idct8_shift7_add64_DW01_add_59 add_152 ( .A({1'b0, x5_18[20], x5_18[20], 
        x5_18[20], x5_18[20:1], 1'b0}), .B({1'b0, x6_89[22], x6_89}), .SUM({
        SYNOPSYS_UNCONNECTED__64, N1092, N1091, N1090, N1089, N1088, N1087, 
        N1086, N1085, N1084, N1083, N1082, N1081, N1080, N1079, N1078, N1077, 
        N1076, N1075, N1074, N1073, N1072, N1071, N1070, N1069}) );
  idct8_shift7_add64_DW01_sub_0 sub_add_152_2_b0 ( .B({N1092, N1091, N1090, 
        N1089, N1088, N1087, N1086, N1085, N1084, N1083, N1082, N1081, N1080, 
        N1079, N1078, N1077, N1076, N1075, N1074, N1073, N1072, N1071, N1070, 
        N1069}), .DIFF({N1116, N1115, N1114, N1113, N1112, N1111, N1110, N1109, 
        N1108, N1107, N1106, N1105, N1104, N1103, N1102, N1101, N1100, N1099, 
        N1098, N1097, N1096, N1095, N1094, N1093}) );
  DFFRHQX1 y6_tmp_reg_24_ ( .D(N1548), .CK(clk), .RN(rstn), .Q(y6_tmp[24]) );
  DFFRHQX1 y6_tmp_reg_23_ ( .D(N1547), .CK(clk), .RN(rstn), .Q(y6_tmp[23]) );
  DFFRHQX1 y7_tmp_reg_24_ ( .D(N1625), .CK(clk), .RN(rstn), .Q(y7_tmp[24]) );
  DFFRHQX1 y7_tmp_reg_23_ ( .D(N1624), .CK(clk), .RN(rstn), .Q(y7_tmp[23]) );
  DFFRHQX1 y0_tmp_reg_24_ ( .D(N1239), .CK(clk), .RN(rstn), .Q(y0_tmp[24]) );
  DFFRHQX1 y0_tmp_reg_23_ ( .D(N1238), .CK(clk), .RN(rstn), .Q(y0_tmp[23]) );
  DFFRHQX1 y1_tmp_reg_24_ ( .D(N1265), .CK(clk), .RN(rstn), .Q(y1_tmp[24]) );
  DFFRHQX1 y1_tmp_reg_23_ ( .D(N1264), .CK(clk), .RN(rstn), .Q(y1_tmp[23]) );
  DFFRHQX1 y2_tmp_reg_24_ ( .D(N1291), .CK(clk), .RN(rstn), .Q(y2_tmp[24]) );
  DFFRHQX1 y2_tmp_reg_23_ ( .D(N1290), .CK(clk), .RN(rstn), .Q(y2_tmp[23]) );
  DFFRHQX1 y3_tmp_reg_24_ ( .D(N1317), .CK(clk), .RN(rstn), .Q(y3_tmp[24]) );
  DFFRHQX1 y3_tmp_reg_23_ ( .D(N1316), .CK(clk), .RN(rstn), .Q(y3_tmp[23]) );
  DFFRHQX1 y4_tmp_reg_24_ ( .D(N1394), .CK(clk), .RN(rstn), .Q(y4_tmp[24]) );
  DFFRHQX1 y4_tmp_reg_23_ ( .D(N1393), .CK(clk), .RN(rstn), .Q(y4_tmp[23]) );
  DFFRHQX1 y5_tmp_reg_24_ ( .D(N1471), .CK(clk), .RN(rstn), .Q(y5_tmp[24]) );
  DFFRHQX1 y5_tmp_reg_23_ ( .D(N1470), .CK(clk), .RN(rstn), .Q(y5_tmp[23]) );
  DFFRHQX1 y6_tmp_reg_25_ ( .D(N1549), .CK(clk), .RN(rstn), .Q(y6_tmp[25]) );
  DFFRHQX1 y7_tmp_reg_25_ ( .D(N1626), .CK(clk), .RN(rstn), .Q(y7_tmp[25]) );
  DFFRHQX1 y0_tmp_reg_25_ ( .D(N1240), .CK(clk), .RN(rstn), .Q(y0_tmp[25]) );
  DFFRHQX1 y1_tmp_reg_25_ ( .D(N1266), .CK(clk), .RN(rstn), .Q(y1_tmp[25]) );
  DFFRHQX1 y2_tmp_reg_25_ ( .D(N1292), .CK(clk), .RN(rstn), .Q(y2_tmp[25]) );
  DFFRHQX1 y3_tmp_reg_25_ ( .D(N1318), .CK(clk), .RN(rstn), .Q(y3_tmp[25]) );
  DFFRHQX1 y4_tmp_reg_25_ ( .D(N1395), .CK(clk), .RN(rstn), .Q(y4_tmp[25]) );
  DFFRHQX1 y5_tmp_reg_25_ ( .D(N1472), .CK(clk), .RN(rstn), .Q(y5_tmp[25]) );
  DFFRHQX1 x4_50_tmp2_reg_4_ ( .D(N85), .CK(clk), .RN(rstn), .Q(x4_50_tmp2[4])
         );
  DFFRHQX1 x4_50_tmp2_reg_3_ ( .D(n76), .CK(clk), .RN(rstn), .Q(x4_50_tmp2[3])
         );
  DFFRHQX1 x4_50_tmp2_reg_2_ ( .D(x4[1]), .CK(clk), .RN(rstn), .Q(
        x4_50_tmp2[2]) );
  DFFRHQX1 x4_50_tmp2_reg_1_ ( .D(x4[0]), .CK(clk), .RN(rstn), .Q(
        x4_50_tmp2[1]) );
  DFFRHQX1 x6_50_tmp2_reg_4_ ( .D(N255), .CK(clk), .RN(rstn), .Q(x6_50_tmp2[4]) );
  DFFRHQX1 x6_50_tmp2_reg_3_ ( .D(n50), .CK(clk), .RN(rstn), .Q(x6_50_tmp2[3])
         );
  DFFRHQX1 x6_50_tmp2_reg_2_ ( .D(x6[1]), .CK(clk), .RN(rstn), .Q(
        x6_50_tmp2[2]) );
  DFFRHQX1 x6_50_tmp2_reg_1_ ( .D(x6[0]), .CK(clk), .RN(rstn), .Q(
        x6_50_tmp2[1]) );
  DFFRHQX1 x5_50_tmp2_reg_4_ ( .D(N170), .CK(clk), .RN(rstn), .Q(x5_50_tmp2[4]) );
  DFFRHQX1 x5_50_tmp2_reg_3_ ( .D(n63), .CK(clk), .RN(rstn), .Q(x5_50_tmp2[3])
         );
  DFFRHQX1 x5_50_tmp2_reg_2_ ( .D(x5[1]), .CK(clk), .RN(rstn), .Q(
        x5_50_tmp2[2]) );
  DFFRHQX1 x5_50_tmp2_reg_1_ ( .D(x5[0]), .CK(clk), .RN(rstn), .Q(
        x5_50_tmp2[1]) );
  DFFRHQX1 x7_50_tmp2_reg_4_ ( .D(N340), .CK(clk), .RN(rstn), .Q(x7_50_tmp2[4]) );
  DFFRHQX1 x7_50_tmp2_reg_3_ ( .D(n37), .CK(clk), .RN(rstn), .Q(x7_50_tmp2[3])
         );
  DFFRHQX1 x7_50_tmp2_reg_2_ ( .D(x7[1]), .CK(clk), .RN(rstn), .Q(
        x7_50_tmp2[2]) );
  DFFRHQX1 x7_50_tmp2_reg_1_ ( .D(x7[0]), .CK(clk), .RN(rstn), .Q(
        x7_50_tmp2[1]) );
  DFFRHQX1 x4_18_tmp2_reg_3_ ( .D(n76), .CK(clk), .RN(rstn), .Q(x4_18_tmp2[3])
         );
  DFFRHQX1 x4_18_tmp2_reg_2_ ( .D(x4[1]), .CK(clk), .RN(rstn), .Q(
        x4_18_tmp2[2]) );
  DFFRHQX1 x4_18_tmp2_reg_1_ ( .D(x4[0]), .CK(clk), .RN(rstn), .Q(
        x4_18_tmp2[1]) );
  DFFRHQX1 x6_18_tmp2_reg_3_ ( .D(n50), .CK(clk), .RN(rstn), .Q(x6_18_tmp2[3])
         );
  DFFRHQX1 x6_18_tmp2_reg_2_ ( .D(x6[1]), .CK(clk), .RN(rstn), .Q(
        x6_18_tmp2[2]) );
  DFFRHQX1 x6_18_tmp2_reg_1_ ( .D(x6[0]), .CK(clk), .RN(rstn), .Q(
        x6_18_tmp2[1]) );
  DFFRHQX1 x5_18_tmp2_reg_3_ ( .D(n63), .CK(clk), .RN(rstn), .Q(x5_18_tmp2[3])
         );
  DFFRHQX1 x5_18_tmp2_reg_2_ ( .D(x5[1]), .CK(clk), .RN(rstn), .Q(
        x5_18_tmp2[2]) );
  DFFRHQX1 x5_18_tmp2_reg_1_ ( .D(x5[0]), .CK(clk), .RN(rstn), .Q(
        x5_18_tmp2[1]) );
  DFFRHQX1 x7_18_tmp2_reg_3_ ( .D(n37), .CK(clk), .RN(rstn), .Q(x7_18_tmp2[3])
         );
  DFFRHQX1 x7_18_tmp2_reg_2_ ( .D(x7[1]), .CK(clk), .RN(rstn), .Q(
        x7_18_tmp2[2]) );
  DFFRHQX1 x7_18_tmp2_reg_1_ ( .D(x7[0]), .CK(clk), .RN(rstn), .Q(
        x7_18_tmp2[1]) );
  DFFRHQX1 x7_89_tmp1_reg_22_ ( .D(x7[15]), .CK(clk), .RN(rstn), .Q(
        x7_89_tmp1[22]) );
  DFFRHQX1 x7_89_tmp1_reg_21_ ( .D(N293), .CK(clk), .RN(rstn), .Q(
        x7_89_tmp1[21]) );
  DFFRHQX1 x7_89_tmp1_reg_20_ ( .D(N292), .CK(clk), .RN(rstn), .Q(
        x7_89_tmp1[20]) );
  DFFRHQX1 x7_89_tmp1_reg_19_ ( .D(N291), .CK(clk), .RN(rstn), .Q(
        x7_89_tmp1[19]) );
  DFFRHQX1 x6_89_tmp1_reg_22_ ( .D(x6[15]), .CK(clk), .RN(rstn), .Q(
        x6_89_tmp1[22]) );
  DFFRHQX1 x6_89_tmp1_reg_21_ ( .D(N208), .CK(clk), .RN(rstn), .Q(
        x6_89_tmp1[21]) );
  DFFRHQX1 x6_89_tmp1_reg_20_ ( .D(N207), .CK(clk), .RN(rstn), .Q(
        x6_89_tmp1[20]) );
  DFFRHQX1 x6_89_tmp1_reg_19_ ( .D(N206), .CK(clk), .RN(rstn), .Q(
        x6_89_tmp1[19]) );
  DFFRHQX1 x5_89_tmp1_reg_22_ ( .D(x5[15]), .CK(clk), .RN(rstn), .Q(
        x5_89_tmp1[22]) );
  DFFRHQX1 x5_89_tmp1_reg_21_ ( .D(N123), .CK(clk), .RN(rstn), .Q(
        x5_89_tmp1[21]) );
  DFFRHQX1 x5_89_tmp1_reg_20_ ( .D(N122), .CK(clk), .RN(rstn), .Q(
        x5_89_tmp1[20]) );
  DFFRHQX1 x5_89_tmp1_reg_19_ ( .D(N121), .CK(clk), .RN(rstn), .Q(
        x5_89_tmp1[19]) );
  DFFRHQX1 x5_75_tmp1_reg_22_ ( .D(x5[15]), .CK(clk), .RN(rstn), .Q(
        x5_75_tmp1[22]) );
  DFFRHQX1 x5_75_tmp1_reg_21_ ( .D(N123), .CK(clk), .RN(rstn), .Q(
        x5_75_tmp1[21]) );
  DFFRHQX1 x5_75_tmp1_reg_20_ ( .D(N122), .CK(clk), .RN(rstn), .Q(
        x5_75_tmp1[20]) );
  DFFRHQX1 x5_75_tmp1_reg_19_ ( .D(N121), .CK(clk), .RN(rstn), .Q(
        x5_75_tmp1[19]) );
  DFFRHQX1 x4_75_tmp1_reg_22_ ( .D(x4[15]), .CK(clk), .RN(rstn), .Q(
        x4_75_tmp1[22]) );
  DFFRHQX1 x4_75_tmp1_reg_21_ ( .D(N38), .CK(clk), .RN(rstn), .Q(
        x4_75_tmp1[21]) );
  DFFRHQX1 x4_75_tmp1_reg_20_ ( .D(N37), .CK(clk), .RN(rstn), .Q(
        x4_75_tmp1[20]) );
  DFFRHQX1 x4_75_tmp1_reg_19_ ( .D(N36), .CK(clk), .RN(rstn), .Q(
        x4_75_tmp1[19]) );
  DFFRHQX1 x7_75_tmp1_reg_22_ ( .D(x7[15]), .CK(clk), .RN(rstn), .Q(
        x7_75_tmp1[22]) );
  DFFRHQX1 x7_75_tmp1_reg_21_ ( .D(N293), .CK(clk), .RN(rstn), .Q(
        x7_75_tmp1[21]) );
  DFFRHQX1 x7_75_tmp1_reg_20_ ( .D(N292), .CK(clk), .RN(rstn), .Q(
        x7_75_tmp1[20]) );
  DFFRHQX1 x7_75_tmp1_reg_19_ ( .D(N291), .CK(clk), .RN(rstn), .Q(
        x7_75_tmp1[19]) );
  DFFRHQX1 x6_75_tmp1_reg_22_ ( .D(x6[15]), .CK(clk), .RN(rstn), .Q(
        x6_75_tmp1[22]) );
  DFFRHQX1 x6_75_tmp1_reg_21_ ( .D(N208), .CK(clk), .RN(rstn), .Q(
        x6_75_tmp1[21]) );
  DFFRHQX1 x6_75_tmp1_reg_20_ ( .D(N207), .CK(clk), .RN(rstn), .Q(
        x6_75_tmp1[20]) );
  DFFRHQX1 x6_75_tmp1_reg_19_ ( .D(N206), .CK(clk), .RN(rstn), .Q(
        x6_75_tmp1[19]) );
  DFFRHQX1 x4_50_tmp1_reg_19_ ( .D(n88), .CK(clk), .RN(rstn), .Q(
        x4_50_tmp1[19]) );
  DFFRHQX1 x4_50_tmp1_reg_18_ ( .D(n87), .CK(clk), .RN(rstn), .Q(
        x4_50_tmp1[18]) );
  DFFRHQX1 x6_50_tmp1_reg_19_ ( .D(n62), .CK(clk), .RN(rstn), .Q(
        x6_50_tmp1[19]) );
  DFFRHQX1 x6_50_tmp1_reg_18_ ( .D(n61), .CK(clk), .RN(rstn), .Q(
        x6_50_tmp1[18]) );
  DFFRHQX1 x5_50_tmp1_reg_19_ ( .D(n75), .CK(clk), .RN(rstn), .Q(
        x5_50_tmp1[19]) );
  DFFRHQX1 x5_50_tmp1_reg_18_ ( .D(n74), .CK(clk), .RN(rstn), .Q(
        x5_50_tmp1[18]) );
  DFFRHQX1 x7_50_tmp1_reg_19_ ( .D(n49), .CK(clk), .RN(rstn), .Q(
        x7_50_tmp1[19]) );
  DFFRHQX1 x7_50_tmp1_reg_18_ ( .D(n48), .CK(clk), .RN(rstn), .Q(
        x7_50_tmp1[18]) );
  DFFRHQX1 x4_18_tmp1_reg_18_ ( .D(n88), .CK(clk), .RN(rstn), .Q(
        x4_18_tmp1[18]) );
  DFFRHQX1 x4_18_tmp1_reg_17_ ( .D(n87), .CK(clk), .RN(rstn), .Q(
        x4_18_tmp1[17]) );
  DFFRHQX1 x5_18_tmp1_reg_18_ ( .D(n75), .CK(clk), .RN(rstn), .Q(
        x5_18_tmp1[18]) );
  DFFRHQX1 x5_18_tmp1_reg_17_ ( .D(n74), .CK(clk), .RN(rstn), .Q(
        x5_18_tmp1[17]) );
  DFFRHQX1 x6_18_tmp1_reg_18_ ( .D(n62), .CK(clk), .RN(rstn), .Q(
        x6_18_tmp1[18]) );
  DFFRHQX1 x6_18_tmp1_reg_17_ ( .D(n61), .CK(clk), .RN(rstn), .Q(
        x6_18_tmp1[17]) );
  DFFRHQX1 x7_18_tmp1_reg_18_ ( .D(n49), .CK(clk), .RN(rstn), .Q(
        x7_18_tmp1[18]) );
  DFFRHQX1 x7_18_tmp1_reg_17_ ( .D(n48), .CK(clk), .RN(rstn), .Q(
        x7_18_tmp1[17]) );
  DFFRHQX1 x4_89_tmp1_reg_22_ ( .D(x4[15]), .CK(clk), .RN(rstn), .Q(
        x4_89_tmp1[22]) );
  DFFRHQX1 x4_89_tmp1_reg_21_ ( .D(N38), .CK(clk), .RN(rstn), .Q(
        x4_89_tmp1[21]) );
  DFFRHQX1 x4_89_tmp1_reg_20_ ( .D(N37), .CK(clk), .RN(rstn), .Q(
        x4_89_tmp1[20]) );
  DFFRHQX1 x4_89_tmp1_reg_19_ ( .D(N36), .CK(clk), .RN(rstn), .Q(
        x4_89_tmp1[19]) );
  DFFRHQX1 x4_89_reg_21_ ( .D(N378), .CK(clk), .RN(rstn), .Q(x4_89[21]) );
  DFFRHQX1 x4_89_reg_20_ ( .D(N377), .CK(clk), .RN(rstn), .Q(x4_89[20]) );
  DFFRHQX1 x4_75_reg_21_ ( .D(N401), .CK(clk), .RN(rstn), .Q(x4_75[21]) );
  DFFRHQX1 x4_75_reg_20_ ( .D(N400), .CK(clk), .RN(rstn), .Q(x4_75[20]) );
  DFFRHQX1 x5_75_reg_21_ ( .D(N490), .CK(clk), .RN(rstn), .Q(x5_75[21]) );
  DFFRHQX1 x5_75_reg_20_ ( .D(N489), .CK(clk), .RN(rstn), .Q(x5_75[20]) );
  DFFRHQX1 x6_75_reg_21_ ( .D(N579), .CK(clk), .RN(rstn), .Q(x6_75[21]) );
  DFFRHQX1 x6_75_reg_20_ ( .D(N578), .CK(clk), .RN(rstn), .Q(x6_75[20]) );
  DFFRHQX1 x4_50_reg_20_ ( .D(N423), .CK(clk), .RN(rstn), .Q(x4_50[20]) );
  DFFRHQX1 x5_tmp1_reg_22_ ( .D(N901), .CK(clk), .RN(rstn), .Q(x5_tmp1[22]) );
  DFFRHQX1 x5_tmp1_reg_21_ ( .D(N900), .CK(clk), .RN(rstn), .Q(x5_tmp1[21]) );
  DFFRHQX1 x6_tmp1_reg_22_ ( .D(N1067), .CK(clk), .RN(rstn), .Q(x6_tmp1[22])
         );
  DFFRHQX1 x6_tmp1_reg_21_ ( .D(N1066), .CK(clk), .RN(rstn), .Q(x6_tmp1[21])
         );
  DFFRHQX1 x7_tmp1_reg_22_ ( .D(N1164), .CK(clk), .RN(rstn), .Q(x7_tmp1[22])
         );
  DFFRHQX1 x7_tmp1_reg_21_ ( .D(N1163), .CK(clk), .RN(rstn), .Q(x7_tmp1[21])
         );
  DFFRHQX1 x4_tmp1_reg_22_ ( .D(N782), .CK(clk), .RN(rstn), .Q(x4_tmp1[22]) );
  DFFRHQX1 x4_tmp1_reg_21_ ( .D(N781), .CK(clk), .RN(rstn), .Q(x4_tmp1[21]) );
  DFFRHQX1 y6_tmp_reg_5_ ( .D(N1529), .CK(clk), .RN(rstn), .Q(y6_tmp[5]) );
  DFFRHQX1 y6_tmp_reg_4_ ( .D(N1528), .CK(clk), .RN(rstn), .Q(y6_tmp[4]) );
  DFFRHQX1 y6_tmp_reg_3_ ( .D(N1527), .CK(clk), .RN(rstn), .Q(y6_tmp[3]) );
  DFFRHQX1 y6_tmp_reg_2_ ( .D(N1526), .CK(clk), .RN(rstn), .Q(y6_tmp[2]) );
  DFFRHQX1 y6_tmp_reg_1_ ( .D(N1525), .CK(clk), .RN(rstn), .Q(y6_tmp[1]) );
  DFFRHQX1 y6_tmp_reg_0_ ( .D(N1524), .CK(clk), .RN(rstn), .Q(y6_tmp[0]) );
  DFFRHQX1 y7_tmp_reg_5_ ( .D(N1606), .CK(clk), .RN(rstn), .Q(y7_tmp[5]) );
  DFFRHQX1 y7_tmp_reg_4_ ( .D(N1605), .CK(clk), .RN(rstn), .Q(y7_tmp[4]) );
  DFFRHQX1 y7_tmp_reg_3_ ( .D(N1604), .CK(clk), .RN(rstn), .Q(y7_tmp[3]) );
  DFFRHQX1 y7_tmp_reg_2_ ( .D(N1603), .CK(clk), .RN(rstn), .Q(y7_tmp[2]) );
  DFFRHQX1 y7_tmp_reg_1_ ( .D(N1602), .CK(clk), .RN(rstn), .Q(y7_tmp[1]) );
  DFFRHQX1 y7_tmp_reg_0_ ( .D(N1601), .CK(clk), .RN(rstn), .Q(y7_tmp[0]) );
  DFFRHQX1 y0_tmp_reg_5_ ( .D(N1220), .CK(clk), .RN(rstn), .Q(y0_tmp[5]) );
  DFFRHQX1 y0_tmp_reg_4_ ( .D(N1219), .CK(clk), .RN(rstn), .Q(y0_tmp[4]) );
  DFFRHQX1 y0_tmp_reg_3_ ( .D(N1218), .CK(clk), .RN(rstn), .Q(y0_tmp[3]) );
  DFFRHQX1 y0_tmp_reg_2_ ( .D(N1217), .CK(clk), .RN(rstn), .Q(y0_tmp[2]) );
  DFFRHQX1 y0_tmp_reg_1_ ( .D(N1216), .CK(clk), .RN(rstn), .Q(y0_tmp[1]) );
  DFFRHQX1 y0_tmp_reg_0_ ( .D(N1215), .CK(clk), .RN(rstn), .Q(y0_tmp[0]) );
  DFFRHQX1 y1_tmp_reg_5_ ( .D(N1246), .CK(clk), .RN(rstn), .Q(y1_tmp[5]) );
  DFFRHQX1 y1_tmp_reg_4_ ( .D(N1245), .CK(clk), .RN(rstn), .Q(y1_tmp[4]) );
  DFFRHQX1 y1_tmp_reg_3_ ( .D(N1244), .CK(clk), .RN(rstn), .Q(y1_tmp[3]) );
  DFFRHQX1 y1_tmp_reg_2_ ( .D(N1243), .CK(clk), .RN(rstn), .Q(y1_tmp[2]) );
  DFFRHQX1 y1_tmp_reg_1_ ( .D(N1242), .CK(clk), .RN(rstn), .Q(y1_tmp[1]) );
  DFFRHQX1 y1_tmp_reg_0_ ( .D(N1241), .CK(clk), .RN(rstn), .Q(y1_tmp[0]) );
  DFFRHQX1 y2_tmp_reg_5_ ( .D(N1272), .CK(clk), .RN(rstn), .Q(y2_tmp[5]) );
  DFFRHQX1 y2_tmp_reg_4_ ( .D(N1271), .CK(clk), .RN(rstn), .Q(y2_tmp[4]) );
  DFFRHQX1 y2_tmp_reg_3_ ( .D(N1270), .CK(clk), .RN(rstn), .Q(y2_tmp[3]) );
  DFFRHQX1 y2_tmp_reg_2_ ( .D(N1269), .CK(clk), .RN(rstn), .Q(y2_tmp[2]) );
  DFFRHQX1 y2_tmp_reg_1_ ( .D(N1268), .CK(clk), .RN(rstn), .Q(y2_tmp[1]) );
  DFFRHQX1 y2_tmp_reg_0_ ( .D(N1267), .CK(clk), .RN(rstn), .Q(y2_tmp[0]) );
  DFFRHQX1 y3_tmp_reg_5_ ( .D(N1298), .CK(clk), .RN(rstn), .Q(y3_tmp[5]) );
  DFFRHQX1 y3_tmp_reg_4_ ( .D(N1297), .CK(clk), .RN(rstn), .Q(y3_tmp[4]) );
  DFFRHQX1 y3_tmp_reg_3_ ( .D(N1296), .CK(clk), .RN(rstn), .Q(y3_tmp[3]) );
  DFFRHQX1 y3_tmp_reg_2_ ( .D(N1295), .CK(clk), .RN(rstn), .Q(y3_tmp[2]) );
  DFFRHQX1 y3_tmp_reg_1_ ( .D(N1294), .CK(clk), .RN(rstn), .Q(y3_tmp[1]) );
  DFFRHQX1 y3_tmp_reg_0_ ( .D(N1293), .CK(clk), .RN(rstn), .Q(y3_tmp[0]) );
  DFFRHQX1 y4_tmp_reg_5_ ( .D(N1375), .CK(clk), .RN(rstn), .Q(y4_tmp[5]) );
  DFFRHQX1 y4_tmp_reg_4_ ( .D(N1374), .CK(clk), .RN(rstn), .Q(y4_tmp[4]) );
  DFFRHQX1 y4_tmp_reg_3_ ( .D(N1373), .CK(clk), .RN(rstn), .Q(y4_tmp[3]) );
  DFFRHQX1 y4_tmp_reg_2_ ( .D(N1372), .CK(clk), .RN(rstn), .Q(y4_tmp[2]) );
  DFFRHQX1 y4_tmp_reg_1_ ( .D(N1371), .CK(clk), .RN(rstn), .Q(y4_tmp[1]) );
  DFFRHQX1 y4_tmp_reg_0_ ( .D(N1370), .CK(clk), .RN(rstn), .Q(y4_tmp[0]) );
  DFFRHQX1 y5_tmp_reg_5_ ( .D(N1452), .CK(clk), .RN(rstn), .Q(y5_tmp[5]) );
  DFFRHQX1 y5_tmp_reg_4_ ( .D(N1451), .CK(clk), .RN(rstn), .Q(y5_tmp[4]) );
  DFFRHQX1 y5_tmp_reg_3_ ( .D(N1450), .CK(clk), .RN(rstn), .Q(y5_tmp[3]) );
  DFFRHQX1 y5_tmp_reg_2_ ( .D(N1449), .CK(clk), .RN(rstn), .Q(y5_tmp[2]) );
  DFFRHQX1 y5_tmp_reg_1_ ( .D(N1448), .CK(clk), .RN(rstn), .Q(y5_tmp[1]) );
  DFFRHQX1 y5_tmp_reg_0_ ( .D(N1447), .CK(clk), .RN(rstn), .Q(y5_tmp[0]) );
  DFFRHQX1 x7_50_reg_21_ ( .D(N691), .CK(clk), .RN(rstn), .Q(x7_50[21]) );
  DFFRHQX1 x7_50_reg_20_ ( .D(N690), .CK(clk), .RN(rstn), .Q(x7_50[20]) );
  DFFRHQX1 x5_89_reg_22_ ( .D(N468), .CK(clk), .RN(rstn), .Q(x5_89[22]) );
  DFFRHQX1 x5_89_reg_21_ ( .D(N467), .CK(clk), .RN(rstn), .Q(x5_89[21]) );
  DFFRHQX1 x5_89_reg_20_ ( .D(N466), .CK(clk), .RN(rstn), .Q(x5_89[20]) );
  DFFRHQX1 x7_89_reg_22_ ( .D(N646), .CK(clk), .RN(rstn), .Q(x7_89[22]) );
  DFFRHQX1 x7_89_reg_21_ ( .D(N645), .CK(clk), .RN(rstn), .Q(x7_89[21]) );
  DFFRHQX1 x7_89_reg_20_ ( .D(N644), .CK(clk), .RN(rstn), .Q(x7_89[20]) );
  DFFRHQX1 x5_50_reg_21_ ( .D(N513), .CK(clk), .RN(rstn), .Q(x5_50[21]) );
  DFFRHQX1 x5_50_reg_20_ ( .D(N512), .CK(clk), .RN(rstn), .Q(x5_50[20]) );
  DFFRHQX1 x4_50_tmp1_reg_20_ ( .D(x4[15]), .CK(clk), .RN(rstn), .Q(
        x4_50_tmp1[20]) );
  DFFRHQX1 x6_50_tmp1_reg_20_ ( .D(x6[15]), .CK(clk), .RN(rstn), .Q(
        x6_50_tmp1[20]) );
  DFFRHQX1 x5_50_tmp1_reg_20_ ( .D(x5[15]), .CK(clk), .RN(rstn), .Q(
        x5_50_tmp1[20]) );
  DFFRHQX1 x7_50_tmp1_reg_20_ ( .D(x7[15]), .CK(clk), .RN(rstn), .Q(
        x7_50_tmp1[20]) );
  DFFRHQX1 x4_18_tmp1_reg_19_ ( .D(x4[15]), .CK(clk), .RN(rstn), .Q(
        x4_18_tmp1[19]) );
  DFFRHQX1 x5_18_tmp1_reg_19_ ( .D(x5[15]), .CK(clk), .RN(rstn), .Q(
        x5_18_tmp1[19]) );
  DFFRHQX1 x6_18_tmp1_reg_19_ ( .D(x6[15]), .CK(clk), .RN(rstn), .Q(
        x6_18_tmp1[19]) );
  DFFRHQX1 x7_18_tmp1_reg_19_ ( .D(x7[15]), .CK(clk), .RN(rstn), .Q(
        x7_18_tmp1[19]) );
  DFFRHQX1 x4_89_reg_22_ ( .D(N379), .CK(clk), .RN(rstn), .Q(x4_89[22]) );
  DFFRHQX1 x4_75_reg_22_ ( .D(N402), .CK(clk), .RN(rstn), .Q(x4_75[22]) );
  DFFRHQX1 x5_75_reg_22_ ( .D(N491), .CK(clk), .RN(rstn), .Q(x5_75[22]) );
  DFFRHQX1 x6_75_reg_22_ ( .D(N580), .CK(clk), .RN(rstn), .Q(x6_75[22]) );
  DFFRHQX1 x5_tmp1_reg_23_ ( .D(N902), .CK(clk), .RN(rstn), .Q(x5_tmp1[23]) );
  DFFRHQX1 x6_tmp1_reg_23_ ( .D(N1068), .CK(clk), .RN(rstn), .Q(x6_tmp1[23])
         );
  DFFRHQX1 x7_tmp1_reg_23_ ( .D(N1165), .CK(clk), .RN(rstn), .Q(x7_tmp1[23])
         );
  DFFRHQX1 x4_tmp1_reg_23_ ( .D(N783), .CK(clk), .RN(rstn), .Q(x4_tmp1[23]) );
  DFFRHQX1 x6_89_tmp2_reg_19_ ( .D(N229), .CK(clk), .RN(rstn), .Q(
        x6_89_tmp2[19]) );
  DFFRHQX1 x5_89_tmp2_reg_19_ ( .D(N144), .CK(clk), .RN(rstn), .Q(
        x5_89_tmp2[19]) );
  DFFRHQX1 x4_89_tmp2_reg_19_ ( .D(N59), .CK(clk), .RN(rstn), .Q(
        x4_89_tmp2[19]) );
  DFFRHQX1 x7_89_tmp2_reg_19_ ( .D(N314), .CK(clk), .RN(rstn), .Q(
        x7_89_tmp2[19]) );
  DFFRHQX1 x4_50_tmp2_reg_19_ ( .D(N100), .CK(clk), .RN(rstn), .Q(
        x4_50_tmp2[19]) );
  DFFRHQX1 x4_50_tmp2_reg_18_ ( .D(N99), .CK(clk), .RN(rstn), .Q(
        x4_50_tmp2[18]) );
  DFFRHQX1 x6_50_tmp2_reg_19_ ( .D(N270), .CK(clk), .RN(rstn), .Q(
        x6_50_tmp2[19]) );
  DFFRHQX1 x6_50_tmp2_reg_18_ ( .D(N269), .CK(clk), .RN(rstn), .Q(
        x6_50_tmp2[18]) );
  DFFRHQX1 x6_50_reg_20_ ( .D(N601), .CK(clk), .RN(rstn), .Q(x6_50[20]) );
  DFFRHQX1 x5_50_tmp2_reg_19_ ( .D(N185), .CK(clk), .RN(rstn), .Q(
        x5_50_tmp2[19]) );
  DFFRHQX1 x5_50_tmp2_reg_18_ ( .D(N184), .CK(clk), .RN(rstn), .Q(
        x5_50_tmp2[18]) );
  DFFRHQX1 x7_50_tmp2_reg_19_ ( .D(N355), .CK(clk), .RN(rstn), .Q(
        x7_50_tmp2[19]) );
  DFFRHQX1 x7_50_tmp2_reg_18_ ( .D(N354), .CK(clk), .RN(rstn), .Q(
        x7_50_tmp2[18]) );
  DFFRHQX1 x6_89_reg_21_ ( .D(N556), .CK(clk), .RN(rstn), .Q(x6_89[21]) );
  DFFRHQX1 x7_75_reg_21_ ( .D(N668), .CK(clk), .RN(rstn), .Q(x7_75[21]) );
  DFFRHQX1 x7_75_reg_20_ ( .D(N667), .CK(clk), .RN(rstn), .Q(x7_75[20]) );
  DFFRHQX1 x4_tmp2_reg_22_ ( .D(N852), .CK(clk), .RN(rstn), .Q(x4_tmp2[22]) );
  DFFRHQX1 x4_tmp2_reg_21_ ( .D(N851), .CK(clk), .RN(rstn), .Q(x4_tmp2[21]) );
  DFFRHQX1 x5_tmp2_reg_22_ ( .D(N972), .CK(clk), .RN(rstn), .Q(x5_tmp2[22]) );
  DFFRHQX1 x5_tmp2_reg_21_ ( .D(N971), .CK(clk), .RN(rstn), .Q(x5_tmp2[21]) );
  DFFRHQX1 x6_tmp2_reg_22_ ( .D(N1115), .CK(clk), .RN(rstn), .Q(x6_tmp2[22])
         );
  DFFRHQX1 x6_tmp2_reg_21_ ( .D(N1114), .CK(clk), .RN(rstn), .Q(x6_tmp2[21])
         );
  DFFRHQX1 x7_tmp2_reg_22_ ( .D(N1188), .CK(clk), .RN(rstn), .Q(x7_tmp2[22])
         );
  DFFRHQX1 x7_tmp2_reg_21_ ( .D(N1187), .CK(clk), .RN(rstn), .Q(x7_tmp2[21])
         );
  DFFRHQX1 x7_89_tmp1_reg_0_ ( .D(x7[0]), .CK(clk), .RN(rstn), .Q(
        x7_89_tmp1[0]) );
  DFFRHQX1 x6_89_tmp1_reg_0_ ( .D(x6[0]), .CK(clk), .RN(rstn), .Q(
        x6_89_tmp1[0]) );
  DFFRHQX1 x5_89_tmp1_reg_0_ ( .D(x5[0]), .CK(clk), .RN(rstn), .Q(
        x5_89_tmp1[0]) );
  DFFRHQX1 x5_75_tmp1_reg_0_ ( .D(x5[0]), .CK(clk), .RN(rstn), .Q(
        x5_75_tmp1[0]) );
  DFFRHQX1 x4_75_tmp1_reg_0_ ( .D(x4[0]), .CK(clk), .RN(rstn), .Q(
        x4_75_tmp1[0]) );
  DFFRHQX1 x7_75_tmp1_reg_0_ ( .D(x7[0]), .CK(clk), .RN(rstn), .Q(
        x7_75_tmp1[0]) );
  DFFRHQX1 x6_75_tmp1_reg_0_ ( .D(x6[0]), .CK(clk), .RN(rstn), .Q(
        x6_75_tmp1[0]) );
  DFFRHQX1 x4_89_tmp1_reg_0_ ( .D(x4[0]), .CK(clk), .RN(rstn), .Q(
        x4_89_tmp1[0]) );
  DFFRHQX1 x4_89_reg_0_ ( .D(N357), .CK(clk), .RN(rstn), .Q(x4_89[0]) );
  DFFRHQX1 x4_50_reg_21_ ( .D(N424), .CK(clk), .RN(rstn), .Q(x4_50[21]) );
  DFFRHQX1 y6_tmp_reg_22_ ( .D(N1546), .CK(clk), .RN(rstn), .Q(y6_tmp[22]) );
  DFFRHQX1 y7_tmp_reg_22_ ( .D(N1623), .CK(clk), .RN(rstn), .Q(y7_tmp[22]) );
  DFFRHQX1 y4_tmp_reg_22_ ( .D(N1392), .CK(clk), .RN(rstn), .Q(y4_tmp[22]) );
  DFFRHQX1 y5_tmp_reg_22_ ( .D(N1469), .CK(clk), .RN(rstn), .Q(y5_tmp[22]) );
  DFFRHQX1 x7_tmp_reg_23_ ( .D(N1213), .CK(clk), .RN(rstn), .Q(x7_tmp[23]) );
  DFFRHQX1 x5_tmp_reg_23_ ( .D(N997), .CK(clk), .RN(rstn), .Q(x5_tmp[23]) );
  DFFRHQX1 x6_tmp_reg_23_ ( .D(N1140), .CK(clk), .RN(rstn), .Q(x6_tmp[23]) );
  DFFRHQX1 x4_tmp_reg_23_ ( .D(N877), .CK(clk), .RN(rstn), .Q(x4_tmp[23]) );
  DFFRHQX1 y6_tmp_reg_21_ ( .D(N1545), .CK(clk), .RN(rstn), .Q(y6_tmp[21]) );
  DFFRHQX1 y7_tmp_reg_21_ ( .D(N1622), .CK(clk), .RN(rstn), .Q(y7_tmp[21]) );
  DFFRHQX1 y4_tmp_reg_21_ ( .D(N1391), .CK(clk), .RN(rstn), .Q(y4_tmp[21]) );
  DFFRHQX1 y5_tmp_reg_21_ ( .D(N1468), .CK(clk), .RN(rstn), .Q(y5_tmp[21]) );
  DFFRHQX1 x4_50_tmp2_reg_20_ ( .D(N101), .CK(clk), .RN(rstn), .Q(
        x4_50_tmp2[20]) );
  DFFRHQX1 x6_50_tmp2_reg_20_ ( .D(N271), .CK(clk), .RN(rstn), .Q(
        x6_50_tmp2[20]) );
  DFFRHQX1 x5_50_tmp2_reg_20_ ( .D(N186), .CK(clk), .RN(rstn), .Q(
        x5_50_tmp2[20]) );
  DFFRHQX1 x7_50_tmp2_reg_20_ ( .D(N356), .CK(clk), .RN(rstn), .Q(
        x7_50_tmp2[20]) );
  DFFRHQX1 x6_89_reg_22_ ( .D(N557), .CK(clk), .RN(rstn), .Q(x6_89[22]) );
  DFFRHQX1 x7_75_reg_22_ ( .D(N669), .CK(clk), .RN(rstn), .Q(x7_75[22]) );
  DFFRHQX1 x4_tmp2_reg_23_ ( .D(N853), .CK(clk), .RN(rstn), .Q(x4_tmp2[23]) );
  DFFRHQX1 x5_tmp2_reg_23_ ( .D(N973), .CK(clk), .RN(rstn), .Q(x5_tmp2[23]) );
  DFFRHQX1 x6_tmp2_reg_23_ ( .D(N1116), .CK(clk), .RN(rstn), .Q(x6_tmp2[23])
         );
  DFFRHQX1 x7_tmp2_reg_23_ ( .D(N1189), .CK(clk), .RN(rstn), .Q(x7_tmp2[23])
         );
  DFFRHQX1 x7_tmp_reg_24_ ( .D(N1214), .CK(clk), .RN(rstn), .Q(x7_tmp[24]) );
  DFFRHQX1 x5_tmp_reg_24_ ( .D(N998), .CK(clk), .RN(rstn), .Q(x5_tmp[24]) );
  DFFRHQX1 x6_tmp_reg_24_ ( .D(N1141), .CK(clk), .RN(rstn), .Q(x6_tmp[24]) );
  DFFRHQX1 x4_tmp_reg_24_ ( .D(N878), .CK(clk), .RN(rstn), .Q(x4_tmp[24]) );
  DFFRHQX1 x6_89_tmp2_reg_20_ ( .D(N230), .CK(clk), .RN(rstn), .Q(
        x6_89_tmp2[20]) );
  DFFRHQX1 x5_89_tmp2_reg_20_ ( .D(N145), .CK(clk), .RN(rstn), .Q(
        x5_89_tmp2[20]) );
  DFFRHQX1 x4_89_tmp2_reg_20_ ( .D(N60), .CK(clk), .RN(rstn), .Q(
        x4_89_tmp2[20]) );
  DFFRHQX1 x7_89_tmp2_reg_20_ ( .D(N315), .CK(clk), .RN(rstn), .Q(
        x7_89_tmp2[20]) );
  DFFRHQX1 x6_50_reg_21_ ( .D(N602), .CK(clk), .RN(rstn), .Q(x6_50[21]) );
  DFFRHQX1 x7_89_tmp1_reg_18_ ( .D(N290), .CK(clk), .RN(rstn), .Q(
        x7_89_tmp1[18]) );
  DFFRHQX1 x7_89_tmp1_reg_17_ ( .D(N289), .CK(clk), .RN(rstn), .Q(
        x7_89_tmp1[17]) );
  DFFRHQX1 x7_89_tmp1_reg_16_ ( .D(N288), .CK(clk), .RN(rstn), .Q(
        x7_89_tmp1[16]) );
  DFFRHQX1 x7_89_tmp1_reg_15_ ( .D(N287), .CK(clk), .RN(rstn), .Q(
        x7_89_tmp1[15]) );
  DFFRHQX1 x6_89_tmp1_reg_18_ ( .D(N205), .CK(clk), .RN(rstn), .Q(
        x6_89_tmp1[18]) );
  DFFRHQX1 x6_89_tmp1_reg_17_ ( .D(N204), .CK(clk), .RN(rstn), .Q(
        x6_89_tmp1[17]) );
  DFFRHQX1 x6_89_tmp1_reg_16_ ( .D(N203), .CK(clk), .RN(rstn), .Q(
        x6_89_tmp1[16]) );
  DFFRHQX1 x6_89_tmp1_reg_15_ ( .D(N202), .CK(clk), .RN(rstn), .Q(
        x6_89_tmp1[15]) );
  DFFRHQX1 x5_89_tmp1_reg_18_ ( .D(N120), .CK(clk), .RN(rstn), .Q(
        x5_89_tmp1[18]) );
  DFFRHQX1 x5_89_tmp1_reg_17_ ( .D(N119), .CK(clk), .RN(rstn), .Q(
        x5_89_tmp1[17]) );
  DFFRHQX1 x5_89_tmp1_reg_16_ ( .D(N118), .CK(clk), .RN(rstn), .Q(
        x5_89_tmp1[16]) );
  DFFRHQX1 x5_89_tmp1_reg_15_ ( .D(N117), .CK(clk), .RN(rstn), .Q(
        x5_89_tmp1[15]) );
  DFFRHQX1 x5_75_tmp1_reg_18_ ( .D(N120), .CK(clk), .RN(rstn), .Q(
        x5_75_tmp1[18]) );
  DFFRHQX1 x5_75_tmp1_reg_17_ ( .D(N119), .CK(clk), .RN(rstn), .Q(
        x5_75_tmp1[17]) );
  DFFRHQX1 x5_75_tmp1_reg_16_ ( .D(N118), .CK(clk), .RN(rstn), .Q(
        x5_75_tmp1[16]) );
  DFFRHQX1 x5_75_tmp1_reg_15_ ( .D(N117), .CK(clk), .RN(rstn), .Q(
        x5_75_tmp1[15]) );
  DFFRHQX1 x4_75_tmp1_reg_18_ ( .D(N35), .CK(clk), .RN(rstn), .Q(
        x4_75_tmp1[18]) );
  DFFRHQX1 x4_75_tmp1_reg_17_ ( .D(N34), .CK(clk), .RN(rstn), .Q(
        x4_75_tmp1[17]) );
  DFFRHQX1 x4_75_tmp1_reg_16_ ( .D(N33), .CK(clk), .RN(rstn), .Q(
        x4_75_tmp1[16]) );
  DFFRHQX1 x4_75_tmp1_reg_15_ ( .D(N32), .CK(clk), .RN(rstn), .Q(
        x4_75_tmp1[15]) );
  DFFRHQX1 x7_75_tmp1_reg_18_ ( .D(N290), .CK(clk), .RN(rstn), .Q(
        x7_75_tmp1[18]) );
  DFFRHQX1 x7_75_tmp1_reg_17_ ( .D(N289), .CK(clk), .RN(rstn), .Q(
        x7_75_tmp1[17]) );
  DFFRHQX1 x7_75_tmp1_reg_16_ ( .D(N288), .CK(clk), .RN(rstn), .Q(
        x7_75_tmp1[16]) );
  DFFRHQX1 x7_75_tmp1_reg_15_ ( .D(N287), .CK(clk), .RN(rstn), .Q(
        x7_75_tmp1[15]) );
  DFFRHQX1 x6_75_tmp1_reg_18_ ( .D(N205), .CK(clk), .RN(rstn), .Q(
        x6_75_tmp1[18]) );
  DFFRHQX1 x6_75_tmp1_reg_17_ ( .D(N204), .CK(clk), .RN(rstn), .Q(
        x6_75_tmp1[17]) );
  DFFRHQX1 x6_75_tmp1_reg_16_ ( .D(N203), .CK(clk), .RN(rstn), .Q(
        x6_75_tmp1[16]) );
  DFFRHQX1 x6_75_tmp1_reg_15_ ( .D(N202), .CK(clk), .RN(rstn), .Q(
        x6_75_tmp1[15]) );
  DFFRHQX1 x4_50_tmp1_reg_17_ ( .D(n86), .CK(clk), .RN(rstn), .Q(
        x4_50_tmp1[17]) );
  DFFRHQX1 x4_50_tmp1_reg_16_ ( .D(n85), .CK(clk), .RN(rstn), .Q(
        x4_50_tmp1[16]) );
  DFFRHQX1 x4_50_tmp1_reg_15_ ( .D(n84), .CK(clk), .RN(rstn), .Q(
        x4_50_tmp1[15]) );
  DFFRHQX1 x4_50_tmp1_reg_14_ ( .D(n83), .CK(clk), .RN(rstn), .Q(
        x4_50_tmp1[14]) );
  DFFRHQX1 x6_50_tmp1_reg_17_ ( .D(n60), .CK(clk), .RN(rstn), .Q(
        x6_50_tmp1[17]) );
  DFFRHQX1 x6_50_tmp1_reg_16_ ( .D(n59), .CK(clk), .RN(rstn), .Q(
        x6_50_tmp1[16]) );
  DFFRHQX1 x6_50_tmp1_reg_15_ ( .D(n58), .CK(clk), .RN(rstn), .Q(
        x6_50_tmp1[15]) );
  DFFRHQX1 x6_50_tmp1_reg_14_ ( .D(n57), .CK(clk), .RN(rstn), .Q(
        x6_50_tmp1[14]) );
  DFFRHQX1 x5_50_tmp1_reg_17_ ( .D(n73), .CK(clk), .RN(rstn), .Q(
        x5_50_tmp1[17]) );
  DFFRHQX1 x5_50_tmp1_reg_16_ ( .D(n72), .CK(clk), .RN(rstn), .Q(
        x5_50_tmp1[16]) );
  DFFRHQX1 x5_50_tmp1_reg_15_ ( .D(n71), .CK(clk), .RN(rstn), .Q(
        x5_50_tmp1[15]) );
  DFFRHQX1 x5_50_tmp1_reg_14_ ( .D(n70), .CK(clk), .RN(rstn), .Q(
        x5_50_tmp1[14]) );
  DFFRHQX1 x7_50_tmp1_reg_17_ ( .D(n47), .CK(clk), .RN(rstn), .Q(
        x7_50_tmp1[17]) );
  DFFRHQX1 x7_50_tmp1_reg_16_ ( .D(n46), .CK(clk), .RN(rstn), .Q(
        x7_50_tmp1[16]) );
  DFFRHQX1 x7_50_tmp1_reg_15_ ( .D(n45), .CK(clk), .RN(rstn), .Q(
        x7_50_tmp1[15]) );
  DFFRHQX1 x7_50_tmp1_reg_14_ ( .D(n44), .CK(clk), .RN(rstn), .Q(
        x7_50_tmp1[14]) );
  DFFRHQX1 x4_18_tmp1_reg_16_ ( .D(n86), .CK(clk), .RN(rstn), .Q(
        x4_18_tmp1[16]) );
  DFFRHQX1 x4_18_tmp1_reg_15_ ( .D(n85), .CK(clk), .RN(rstn), .Q(
        x4_18_tmp1[15]) );
  DFFRHQX1 x4_18_tmp1_reg_14_ ( .D(n84), .CK(clk), .RN(rstn), .Q(
        x4_18_tmp1[14]) );
  DFFRHQX1 x4_18_tmp1_reg_13_ ( .D(n83), .CK(clk), .RN(rstn), .Q(
        x4_18_tmp1[13]) );
  DFFRHQX1 x5_18_tmp1_reg_16_ ( .D(n73), .CK(clk), .RN(rstn), .Q(
        x5_18_tmp1[16]) );
  DFFRHQX1 x5_18_tmp1_reg_15_ ( .D(n72), .CK(clk), .RN(rstn), .Q(
        x5_18_tmp1[15]) );
  DFFRHQX1 x5_18_tmp1_reg_14_ ( .D(n71), .CK(clk), .RN(rstn), .Q(
        x5_18_tmp1[14]) );
  DFFRHQX1 x5_18_tmp1_reg_13_ ( .D(n70), .CK(clk), .RN(rstn), .Q(
        x5_18_tmp1[13]) );
  DFFRHQX1 x6_18_tmp1_reg_16_ ( .D(n60), .CK(clk), .RN(rstn), .Q(
        x6_18_tmp1[16]) );
  DFFRHQX1 x6_18_tmp1_reg_15_ ( .D(n59), .CK(clk), .RN(rstn), .Q(
        x6_18_tmp1[15]) );
  DFFRHQX1 x6_18_tmp1_reg_14_ ( .D(n58), .CK(clk), .RN(rstn), .Q(
        x6_18_tmp1[14]) );
  DFFRHQX1 x6_18_tmp1_reg_13_ ( .D(n57), .CK(clk), .RN(rstn), .Q(
        x6_18_tmp1[13]) );
  DFFRHQX1 x7_18_tmp1_reg_16_ ( .D(n47), .CK(clk), .RN(rstn), .Q(
        x7_18_tmp1[16]) );
  DFFRHQX1 x7_18_tmp1_reg_15_ ( .D(n46), .CK(clk), .RN(rstn), .Q(
        x7_18_tmp1[15]) );
  DFFRHQX1 x7_18_tmp1_reg_14_ ( .D(n45), .CK(clk), .RN(rstn), .Q(
        x7_18_tmp1[14]) );
  DFFRHQX1 x7_18_tmp1_reg_13_ ( .D(n44), .CK(clk), .RN(rstn), .Q(
        x7_18_tmp1[13]) );
  DFFRHQX1 x5_18_reg_19_ ( .D(N533), .CK(clk), .RN(rstn), .Q(x5_18[19]) );
  DFFRHQX1 x5_18_reg_18_ ( .D(N532), .CK(clk), .RN(rstn), .Q(x5_18[18]) );
  DFFRHQX1 x5_18_reg_17_ ( .D(N531), .CK(clk), .RN(rstn), .Q(x5_18[17]) );
  DFFRHQX1 x6_18_reg_19_ ( .D(N622), .CK(clk), .RN(rstn), .Q(x6_18[19]) );
  DFFRHQX1 x6_18_reg_18_ ( .D(N621), .CK(clk), .RN(rstn), .Q(x6_18[18]) );
  DFFRHQX1 x6_18_reg_17_ ( .D(N620), .CK(clk), .RN(rstn), .Q(x6_18[17]) );
  DFFRHQX1 x6_18_reg_16_ ( .D(N619), .CK(clk), .RN(rstn), .Q(x6_18[16]) );
  DFFRHQX1 x4_18_reg_19_ ( .D(N444), .CK(clk), .RN(rstn), .Q(x4_18[19]) );
  DFFRHQX1 x4_18_reg_18_ ( .D(N443), .CK(clk), .RN(rstn), .Q(x4_18[18]) );
  DFFRHQX1 x4_18_reg_17_ ( .D(N442), .CK(clk), .RN(rstn), .Q(x4_18[17]) );
  DFFRHQX1 x4_18_reg_16_ ( .D(N441), .CK(clk), .RN(rstn), .Q(x4_18[16]) );
  DFFRHQX1 x4_89_tmp1_reg_18_ ( .D(N35), .CK(clk), .RN(rstn), .Q(
        x4_89_tmp1[18]) );
  DFFRHQX1 x4_89_tmp1_reg_17_ ( .D(N34), .CK(clk), .RN(rstn), .Q(
        x4_89_tmp1[17]) );
  DFFRHQX1 x4_89_tmp1_reg_16_ ( .D(N33), .CK(clk), .RN(rstn), .Q(
        x4_89_tmp1[16]) );
  DFFRHQX1 x4_89_tmp1_reg_15_ ( .D(N32), .CK(clk), .RN(rstn), .Q(
        x4_89_tmp1[15]) );
  DFFRHQX1 x4_89_reg_19_ ( .D(N376), .CK(clk), .RN(rstn), .Q(x4_89[19]) );
  DFFRHQX1 x4_89_reg_18_ ( .D(N375), .CK(clk), .RN(rstn), .Q(x4_89[18]) );
  DFFRHQX1 x4_89_reg_17_ ( .D(N374), .CK(clk), .RN(rstn), .Q(x4_89[17]) );
  DFFRHQX1 x4_89_reg_16_ ( .D(N373), .CK(clk), .RN(rstn), .Q(x4_89[16]) );
  DFFRHQX1 x4_75_reg_19_ ( .D(N399), .CK(clk), .RN(rstn), .Q(x4_75[19]) );
  DFFRHQX1 x4_75_reg_18_ ( .D(N398), .CK(clk), .RN(rstn), .Q(x4_75[18]) );
  DFFRHQX1 x4_75_reg_17_ ( .D(N397), .CK(clk), .RN(rstn), .Q(x4_75[17]) );
  DFFRHQX1 x4_75_reg_16_ ( .D(N396), .CK(clk), .RN(rstn), .Q(x4_75[16]) );
  DFFRHQX1 x5_75_reg_19_ ( .D(N488), .CK(clk), .RN(rstn), .Q(x5_75[19]) );
  DFFRHQX1 x5_75_reg_18_ ( .D(N487), .CK(clk), .RN(rstn), .Q(x5_75[18]) );
  DFFRHQX1 x5_75_reg_17_ ( .D(N486), .CK(clk), .RN(rstn), .Q(x5_75[17]) );
  DFFRHQX1 x5_75_reg_16_ ( .D(N485), .CK(clk), .RN(rstn), .Q(x5_75[16]) );
  DFFRHQX1 x6_75_reg_19_ ( .D(N577), .CK(clk), .RN(rstn), .Q(x6_75[19]) );
  DFFRHQX1 x6_75_reg_18_ ( .D(N576), .CK(clk), .RN(rstn), .Q(x6_75[18]) );
  DFFRHQX1 x6_75_reg_17_ ( .D(N575), .CK(clk), .RN(rstn), .Q(x6_75[17]) );
  DFFRHQX1 x6_75_reg_16_ ( .D(N574), .CK(clk), .RN(rstn), .Q(x6_75[16]) );
  DFFRHQX1 x4_50_reg_19_ ( .D(N422), .CK(clk), .RN(rstn), .Q(x4_50[19]) );
  DFFRHQX1 x4_50_reg_18_ ( .D(N421), .CK(clk), .RN(rstn), .Q(x4_50[18]) );
  DFFRHQX1 x4_50_reg_17_ ( .D(N420), .CK(clk), .RN(rstn), .Q(x4_50[17]) );
  DFFRHQX1 x4_50_reg_16_ ( .D(N419), .CK(clk), .RN(rstn), .Q(x4_50[16]) );
  DFFRHQX1 x5_tmp1_reg_20_ ( .D(N899), .CK(clk), .RN(rstn), .Q(x5_tmp1[20]) );
  DFFRHQX1 x5_tmp1_reg_19_ ( .D(N898), .CK(clk), .RN(rstn), .Q(x5_tmp1[19]) );
  DFFRHQX1 x5_tmp1_reg_18_ ( .D(N897), .CK(clk), .RN(rstn), .Q(x5_tmp1[18]) );
  DFFRHQX1 x5_tmp1_reg_17_ ( .D(N896), .CK(clk), .RN(rstn), .Q(x5_tmp1[17]) );
  DFFRHQX1 x6_tmp1_reg_20_ ( .D(N1065), .CK(clk), .RN(rstn), .Q(x6_tmp1[20])
         );
  DFFRHQX1 x6_tmp1_reg_19_ ( .D(N1064), .CK(clk), .RN(rstn), .Q(x6_tmp1[19])
         );
  DFFRHQX1 x6_tmp1_reg_18_ ( .D(N1063), .CK(clk), .RN(rstn), .Q(x6_tmp1[18])
         );
  DFFRHQX1 x6_tmp1_reg_17_ ( .D(N1062), .CK(clk), .RN(rstn), .Q(x6_tmp1[17])
         );
  DFFRHQX1 x7_tmp1_reg_20_ ( .D(N1162), .CK(clk), .RN(rstn), .Q(x7_tmp1[20])
         );
  DFFRHQX1 x7_tmp1_reg_19_ ( .D(N1161), .CK(clk), .RN(rstn), .Q(x7_tmp1[19])
         );
  DFFRHQX1 x7_tmp1_reg_18_ ( .D(N1160), .CK(clk), .RN(rstn), .Q(x7_tmp1[18])
         );
  DFFRHQX1 x7_tmp1_reg_17_ ( .D(N1159), .CK(clk), .RN(rstn), .Q(x7_tmp1[17])
         );
  DFFRHQX1 x4_tmp1_reg_20_ ( .D(N780), .CK(clk), .RN(rstn), .Q(x4_tmp1[20]) );
  DFFRHQX1 x4_tmp1_reg_19_ ( .D(N779), .CK(clk), .RN(rstn), .Q(x4_tmp1[19]) );
  DFFRHQX1 x4_tmp1_reg_18_ ( .D(N778), .CK(clk), .RN(rstn), .Q(x4_tmp1[18]) );
  DFFRHQX1 x4_tmp1_reg_17_ ( .D(N777), .CK(clk), .RN(rstn), .Q(x4_tmp1[17]) );
  DFFRHQX1 x7_50_reg_19_ ( .D(N689), .CK(clk), .RN(rstn), .Q(x7_50[19]) );
  DFFRHQX1 x7_50_reg_18_ ( .D(N688), .CK(clk), .RN(rstn), .Q(x7_50[18]) );
  DFFRHQX1 x7_50_reg_17_ ( .D(N687), .CK(clk), .RN(rstn), .Q(x7_50[17]) );
  DFFRHQX1 x7_50_reg_16_ ( .D(N686), .CK(clk), .RN(rstn), .Q(x7_50[16]) );
  DFFRHQX1 x5_89_reg_19_ ( .D(N465), .CK(clk), .RN(rstn), .Q(x5_89[19]) );
  DFFRHQX1 x5_89_reg_18_ ( .D(N464), .CK(clk), .RN(rstn), .Q(x5_89[18]) );
  DFFRHQX1 x5_89_reg_17_ ( .D(N463), .CK(clk), .RN(rstn), .Q(x5_89[17]) );
  DFFRHQX1 x5_89_reg_16_ ( .D(N462), .CK(clk), .RN(rstn), .Q(x5_89[16]) );
  DFFRHQX1 x7_89_reg_19_ ( .D(N643), .CK(clk), .RN(rstn), .Q(x7_89[19]) );
  DFFRHQX1 x7_89_reg_18_ ( .D(N642), .CK(clk), .RN(rstn), .Q(x7_89[18]) );
  DFFRHQX1 x7_89_reg_17_ ( .D(N641), .CK(clk), .RN(rstn), .Q(x7_89[17]) );
  DFFRHQX1 x7_89_reg_16_ ( .D(N640), .CK(clk), .RN(rstn), .Q(x7_89[16]) );
  DFFRHQX1 x5_50_reg_19_ ( .D(N511), .CK(clk), .RN(rstn), .Q(x5_50[19]) );
  DFFRHQX1 x5_50_reg_18_ ( .D(N510), .CK(clk), .RN(rstn), .Q(x5_50[18]) );
  DFFRHQX1 x5_50_reg_17_ ( .D(N509), .CK(clk), .RN(rstn), .Q(x5_50[17]) );
  DFFRHQX1 x5_50_reg_16_ ( .D(N508), .CK(clk), .RN(rstn), .Q(x5_50[16]) );
  DFFRHQX1 x6_89_tmp2_reg_18_ ( .D(N228), .CK(clk), .RN(rstn), .Q(
        x6_89_tmp2[18]) );
  DFFRHQX1 x6_89_tmp2_reg_17_ ( .D(N227), .CK(clk), .RN(rstn), .Q(
        x6_89_tmp2[17]) );
  DFFRHQX1 x6_89_tmp2_reg_16_ ( .D(N226), .CK(clk), .RN(rstn), .Q(
        x6_89_tmp2[16]) );
  DFFRHQX1 x6_89_tmp2_reg_15_ ( .D(N225), .CK(clk), .RN(rstn), .Q(
        x6_89_tmp2[15]) );
  DFFRHQX1 x6_89_tmp2_reg_14_ ( .D(N224), .CK(clk), .RN(rstn), .Q(
        x6_89_tmp2[14]) );
  DFFRHQX1 x5_89_tmp2_reg_18_ ( .D(N143), .CK(clk), .RN(rstn), .Q(
        x5_89_tmp2[18]) );
  DFFRHQX1 x5_89_tmp2_reg_17_ ( .D(N142), .CK(clk), .RN(rstn), .Q(
        x5_89_tmp2[17]) );
  DFFRHQX1 x5_89_tmp2_reg_16_ ( .D(N141), .CK(clk), .RN(rstn), .Q(
        x5_89_tmp2[16]) );
  DFFRHQX1 x5_89_tmp2_reg_15_ ( .D(N140), .CK(clk), .RN(rstn), .Q(
        x5_89_tmp2[15]) );
  DFFRHQX1 x5_89_tmp2_reg_14_ ( .D(N139), .CK(clk), .RN(rstn), .Q(
        x5_89_tmp2[14]) );
  DFFRHQX1 x4_89_tmp2_reg_18_ ( .D(N58), .CK(clk), .RN(rstn), .Q(
        x4_89_tmp2[18]) );
  DFFRHQX1 x4_89_tmp2_reg_17_ ( .D(N57), .CK(clk), .RN(rstn), .Q(
        x4_89_tmp2[17]) );
  DFFRHQX1 x4_89_tmp2_reg_16_ ( .D(N56), .CK(clk), .RN(rstn), .Q(
        x4_89_tmp2[16]) );
  DFFRHQX1 x4_89_tmp2_reg_15_ ( .D(N55), .CK(clk), .RN(rstn), .Q(
        x4_89_tmp2[15]) );
  DFFRHQX1 x4_89_tmp2_reg_14_ ( .D(N54), .CK(clk), .RN(rstn), .Q(
        x4_89_tmp2[14]) );
  DFFRHQX1 x7_89_tmp2_reg_18_ ( .D(N313), .CK(clk), .RN(rstn), .Q(
        x7_89_tmp2[18]) );
  DFFRHQX1 x7_89_tmp2_reg_17_ ( .D(N312), .CK(clk), .RN(rstn), .Q(
        x7_89_tmp2[17]) );
  DFFRHQX1 x7_89_tmp2_reg_16_ ( .D(N311), .CK(clk), .RN(rstn), .Q(
        x7_89_tmp2[16]) );
  DFFRHQX1 x7_89_tmp2_reg_15_ ( .D(N310), .CK(clk), .RN(rstn), .Q(
        x7_89_tmp2[15]) );
  DFFRHQX1 x7_89_tmp2_reg_14_ ( .D(N309), .CK(clk), .RN(rstn), .Q(
        x7_89_tmp2[14]) );
  DFFRHQX1 x4_75_tmp2_reg_18_ ( .D(N79), .CK(clk), .RN(rstn), .Q(
        x4_75_tmp2[18]) );
  DFFRHQX1 x4_75_tmp2_reg_17_ ( .D(N78), .CK(clk), .RN(rstn), .Q(
        x4_75_tmp2[17]) );
  DFFRHQX1 x4_75_tmp2_reg_16_ ( .D(N77), .CK(clk), .RN(rstn), .Q(
        x4_75_tmp2[16]) );
  DFFRHQX1 x4_75_tmp2_reg_15_ ( .D(N76), .CK(clk), .RN(rstn), .Q(
        x4_75_tmp2[15]) );
  DFFRHQX1 x4_75_tmp2_reg_14_ ( .D(N75), .CK(clk), .RN(rstn), .Q(
        x4_75_tmp2[14]) );
  DFFRHQX1 x5_75_tmp2_reg_18_ ( .D(N164), .CK(clk), .RN(rstn), .Q(
        x5_75_tmp2[18]) );
  DFFRHQX1 x5_75_tmp2_reg_17_ ( .D(N163), .CK(clk), .RN(rstn), .Q(
        x5_75_tmp2[17]) );
  DFFRHQX1 x5_75_tmp2_reg_16_ ( .D(N162), .CK(clk), .RN(rstn), .Q(
        x5_75_tmp2[16]) );
  DFFRHQX1 x5_75_tmp2_reg_15_ ( .D(N161), .CK(clk), .RN(rstn), .Q(
        x5_75_tmp2[15]) );
  DFFRHQX1 x5_75_tmp2_reg_14_ ( .D(N160), .CK(clk), .RN(rstn), .Q(
        x5_75_tmp2[14]) );
  DFFRHQX1 x6_75_tmp2_reg_18_ ( .D(N249), .CK(clk), .RN(rstn), .Q(
        x6_75_tmp2[18]) );
  DFFRHQX1 x6_75_tmp2_reg_17_ ( .D(N248), .CK(clk), .RN(rstn), .Q(
        x6_75_tmp2[17]) );
  DFFRHQX1 x6_75_tmp2_reg_16_ ( .D(N247), .CK(clk), .RN(rstn), .Q(
        x6_75_tmp2[16]) );
  DFFRHQX1 x6_75_tmp2_reg_15_ ( .D(N246), .CK(clk), .RN(rstn), .Q(
        x6_75_tmp2[15]) );
  DFFRHQX1 x6_75_tmp2_reg_14_ ( .D(N245), .CK(clk), .RN(rstn), .Q(
        x6_75_tmp2[14]) );
  DFFRHQX1 x7_75_tmp2_reg_18_ ( .D(N334), .CK(clk), .RN(rstn), .Q(
        x7_75_tmp2[18]) );
  DFFRHQX1 x7_75_tmp2_reg_17_ ( .D(N333), .CK(clk), .RN(rstn), .Q(
        x7_75_tmp2[17]) );
  DFFRHQX1 x7_75_tmp2_reg_16_ ( .D(N332), .CK(clk), .RN(rstn), .Q(
        x7_75_tmp2[16]) );
  DFFRHQX1 x7_75_tmp2_reg_15_ ( .D(N331), .CK(clk), .RN(rstn), .Q(
        x7_75_tmp2[15]) );
  DFFRHQX1 x7_75_tmp2_reg_14_ ( .D(N330), .CK(clk), .RN(rstn), .Q(
        x7_75_tmp2[14]) );
  DFFRHQX1 x4_50_tmp2_reg_17_ ( .D(N98), .CK(clk), .RN(rstn), .Q(
        x4_50_tmp2[17]) );
  DFFRHQX1 x4_50_tmp2_reg_16_ ( .D(N97), .CK(clk), .RN(rstn), .Q(
        x4_50_tmp2[16]) );
  DFFRHQX1 x4_50_tmp2_reg_15_ ( .D(N96), .CK(clk), .RN(rstn), .Q(
        x4_50_tmp2[15]) );
  DFFRHQX1 x4_50_tmp2_reg_14_ ( .D(N95), .CK(clk), .RN(rstn), .Q(
        x4_50_tmp2[14]) );
  DFFRHQX1 x4_50_tmp2_reg_13_ ( .D(N94), .CK(clk), .RN(rstn), .Q(
        x4_50_tmp2[13]) );
  DFFRHQX1 x6_50_tmp2_reg_17_ ( .D(N268), .CK(clk), .RN(rstn), .Q(
        x6_50_tmp2[17]) );
  DFFRHQX1 x6_50_tmp2_reg_16_ ( .D(N267), .CK(clk), .RN(rstn), .Q(
        x6_50_tmp2[16]) );
  DFFRHQX1 x6_50_tmp2_reg_15_ ( .D(N266), .CK(clk), .RN(rstn), .Q(
        x6_50_tmp2[15]) );
  DFFRHQX1 x6_50_tmp2_reg_14_ ( .D(N265), .CK(clk), .RN(rstn), .Q(
        x6_50_tmp2[14]) );
  DFFRHQX1 x6_50_tmp2_reg_13_ ( .D(N264), .CK(clk), .RN(rstn), .Q(
        x6_50_tmp2[13]) );
  DFFRHQX1 x6_50_reg_15_ ( .D(N596), .CK(clk), .RN(rstn), .Q(x6_50[15]) );
  DFFRHQX1 x6_50_reg_16_ ( .D(N597), .CK(clk), .RN(rstn), .Q(x6_50[16]) );
  DFFRHQX1 x6_50_reg_17_ ( .D(N598), .CK(clk), .RN(rstn), .Q(x6_50[17]) );
  DFFRHQX1 x6_50_reg_18_ ( .D(N599), .CK(clk), .RN(rstn), .Q(x6_50[18]) );
  DFFRHQX1 x6_50_reg_19_ ( .D(N600), .CK(clk), .RN(rstn), .Q(x6_50[19]) );
  DFFRHQX1 x5_50_tmp2_reg_17_ ( .D(N183), .CK(clk), .RN(rstn), .Q(
        x5_50_tmp2[17]) );
  DFFRHQX1 x5_50_tmp2_reg_16_ ( .D(N182), .CK(clk), .RN(rstn), .Q(
        x5_50_tmp2[16]) );
  DFFRHQX1 x5_50_tmp2_reg_15_ ( .D(N181), .CK(clk), .RN(rstn), .Q(
        x5_50_tmp2[15]) );
  DFFRHQX1 x5_50_tmp2_reg_14_ ( .D(N180), .CK(clk), .RN(rstn), .Q(
        x5_50_tmp2[14]) );
  DFFRHQX1 x5_50_tmp2_reg_13_ ( .D(N179), .CK(clk), .RN(rstn), .Q(
        x5_50_tmp2[13]) );
  DFFRHQX1 x7_50_tmp2_reg_17_ ( .D(N353), .CK(clk), .RN(rstn), .Q(
        x7_50_tmp2[17]) );
  DFFRHQX1 x7_50_tmp2_reg_16_ ( .D(N352), .CK(clk), .RN(rstn), .Q(
        x7_50_tmp2[16]) );
  DFFRHQX1 x7_50_tmp2_reg_15_ ( .D(N351), .CK(clk), .RN(rstn), .Q(
        x7_50_tmp2[15]) );
  DFFRHQX1 x7_50_tmp2_reg_14_ ( .D(N350), .CK(clk), .RN(rstn), .Q(
        x7_50_tmp2[14]) );
  DFFRHQX1 x7_50_tmp2_reg_13_ ( .D(N349), .CK(clk), .RN(rstn), .Q(
        x7_50_tmp2[13]) );
  DFFRHQX1 x4_18_tmp2_reg_15_ ( .D(n88), .CK(clk), .RN(rstn), .Q(
        x4_18_tmp2[15]) );
  DFFRHQX1 x4_18_tmp2_reg_14_ ( .D(n87), .CK(clk), .RN(rstn), .Q(
        x4_18_tmp2[14]) );
  DFFRHQX1 x4_18_tmp2_reg_13_ ( .D(n86), .CK(clk), .RN(rstn), .Q(
        x4_18_tmp2[13]) );
  DFFRHQX1 x4_18_tmp2_reg_12_ ( .D(n85), .CK(clk), .RN(rstn), .Q(
        x4_18_tmp2[12]) );
  DFFRHQX1 x6_18_tmp2_reg_15_ ( .D(n62), .CK(clk), .RN(rstn), .Q(
        x6_18_tmp2[15]) );
  DFFRHQX1 x6_18_tmp2_reg_14_ ( .D(n61), .CK(clk), .RN(rstn), .Q(
        x6_18_tmp2[14]) );
  DFFRHQX1 x6_18_tmp2_reg_13_ ( .D(n60), .CK(clk), .RN(rstn), .Q(
        x6_18_tmp2[13]) );
  DFFRHQX1 x6_18_tmp2_reg_12_ ( .D(n59), .CK(clk), .RN(rstn), .Q(
        x6_18_tmp2[12]) );
  DFFRHQX1 x5_18_tmp2_reg_15_ ( .D(n75), .CK(clk), .RN(rstn), .Q(
        x5_18_tmp2[15]) );
  DFFRHQX1 x5_18_tmp2_reg_14_ ( .D(n74), .CK(clk), .RN(rstn), .Q(
        x5_18_tmp2[14]) );
  DFFRHQX1 x5_18_tmp2_reg_13_ ( .D(n73), .CK(clk), .RN(rstn), .Q(
        x5_18_tmp2[13]) );
  DFFRHQX1 x5_18_tmp2_reg_12_ ( .D(n72), .CK(clk), .RN(rstn), .Q(
        x5_18_tmp2[12]) );
  DFFRHQX1 x7_18_tmp2_reg_15_ ( .D(n49), .CK(clk), .RN(rstn), .Q(
        x7_18_tmp2[15]) );
  DFFRHQX1 x7_18_tmp2_reg_14_ ( .D(n48), .CK(clk), .RN(rstn), .Q(
        x7_18_tmp2[14]) );
  DFFRHQX1 x7_18_tmp2_reg_13_ ( .D(n47), .CK(clk), .RN(rstn), .Q(
        x7_18_tmp2[13]) );
  DFFRHQX1 x7_18_tmp2_reg_12_ ( .D(n46), .CK(clk), .RN(rstn), .Q(
        x7_18_tmp2[12]) );
  DFFRHQX1 x7_18_reg_19_ ( .D(N711), .CK(clk), .RN(rstn), .Q(x7_18[19]) );
  DFFRHQX1 x7_18_reg_18_ ( .D(N710), .CK(clk), .RN(rstn), .Q(x7_18[18]) );
  DFFRHQX1 x7_18_reg_17_ ( .D(N709), .CK(clk), .RN(rstn), .Q(x7_18[17]) );
  DFFRHQX1 x7_18_reg_16_ ( .D(N708), .CK(clk), .RN(rstn), .Q(x7_18[16]) );
  DFFRHQX1 x7_18_reg_15_ ( .D(N707), .CK(clk), .RN(rstn), .Q(x7_18[15]) );
  DFFRHQX1 x6_89_reg_20_ ( .D(N555), .CK(clk), .RN(rstn), .Q(x6_89[20]) );
  DFFRHQX1 x6_89_reg_19_ ( .D(N554), .CK(clk), .RN(rstn), .Q(x6_89[19]) );
  DFFRHQX1 x6_89_reg_18_ ( .D(N553), .CK(clk), .RN(rstn), .Q(x6_89[18]) );
  DFFRHQX1 x6_89_reg_17_ ( .D(N552), .CK(clk), .RN(rstn), .Q(x6_89[17]) );
  DFFRHQX1 x7_75_reg_19_ ( .D(N666), .CK(clk), .RN(rstn), .Q(x7_75[19]) );
  DFFRHQX1 x7_75_reg_18_ ( .D(N665), .CK(clk), .RN(rstn), .Q(x7_75[18]) );
  DFFRHQX1 x7_75_reg_17_ ( .D(N664), .CK(clk), .RN(rstn), .Q(x7_75[17]) );
  DFFRHQX1 x7_75_reg_16_ ( .D(N663), .CK(clk), .RN(rstn), .Q(x7_75[16]) );
  DFFRHQX1 x7_75_reg_15_ ( .D(N662), .CK(clk), .RN(rstn), .Q(x7_75[15]) );
  DFFRHQX1 x4_tmp2_reg_20_ ( .D(N850), .CK(clk), .RN(rstn), .Q(x4_tmp2[20]) );
  DFFRHQX1 x4_tmp2_reg_19_ ( .D(N849), .CK(clk), .RN(rstn), .Q(x4_tmp2[19]) );
  DFFRHQX1 x4_tmp2_reg_18_ ( .D(N848), .CK(clk), .RN(rstn), .Q(x4_tmp2[18]) );
  DFFRHQX1 x4_tmp2_reg_17_ ( .D(N847), .CK(clk), .RN(rstn), .Q(x4_tmp2[17]) );
  DFFRHQX1 x4_tmp2_reg_16_ ( .D(N846), .CK(clk), .RN(rstn), .Q(x4_tmp2[16]) );
  DFFRHQX1 x5_tmp2_reg_20_ ( .D(N970), .CK(clk), .RN(rstn), .Q(x5_tmp2[20]) );
  DFFRHQX1 x5_tmp2_reg_19_ ( .D(N969), .CK(clk), .RN(rstn), .Q(x5_tmp2[19]) );
  DFFRHQX1 x5_tmp2_reg_18_ ( .D(N968), .CK(clk), .RN(rstn), .Q(x5_tmp2[18]) );
  DFFRHQX1 x5_tmp2_reg_17_ ( .D(N967), .CK(clk), .RN(rstn), .Q(x5_tmp2[17]) );
  DFFRHQX1 x5_tmp2_reg_16_ ( .D(N966), .CK(clk), .RN(rstn), .Q(x5_tmp2[16]) );
  DFFRHQX1 x6_tmp2_reg_20_ ( .D(N1113), .CK(clk), .RN(rstn), .Q(x6_tmp2[20])
         );
  DFFRHQX1 x6_tmp2_reg_19_ ( .D(N1112), .CK(clk), .RN(rstn), .Q(x6_tmp2[19])
         );
  DFFRHQX1 x6_tmp2_reg_18_ ( .D(N1111), .CK(clk), .RN(rstn), .Q(x6_tmp2[18])
         );
  DFFRHQX1 x6_tmp2_reg_17_ ( .D(N1110), .CK(clk), .RN(rstn), .Q(x6_tmp2[17])
         );
  DFFRHQX1 x6_tmp2_reg_16_ ( .D(N1109), .CK(clk), .RN(rstn), .Q(x6_tmp2[16])
         );
  DFFRHQX1 x7_tmp2_reg_20_ ( .D(N1186), .CK(clk), .RN(rstn), .Q(x7_tmp2[20])
         );
  DFFRHQX1 x7_tmp2_reg_19_ ( .D(N1185), .CK(clk), .RN(rstn), .Q(x7_tmp2[19])
         );
  DFFRHQX1 x7_tmp2_reg_18_ ( .D(N1184), .CK(clk), .RN(rstn), .Q(x7_tmp2[18])
         );
  DFFRHQX1 x7_tmp2_reg_17_ ( .D(N1183), .CK(clk), .RN(rstn), .Q(x7_tmp2[17])
         );
  DFFRHQX1 x7_tmp2_reg_16_ ( .D(N1182), .CK(clk), .RN(rstn), .Q(x7_tmp2[16])
         );
  DFFRHQX1 y0_tmp_reg_22_ ( .D(N1237), .CK(clk), .RN(rstn), .Q(y0_tmp[22]) );
  DFFRHQX1 y1_tmp_reg_22_ ( .D(N1263), .CK(clk), .RN(rstn), .Q(y1_tmp[22]) );
  DFFRHQX1 y2_tmp_reg_22_ ( .D(N1289), .CK(clk), .RN(rstn), .Q(y2_tmp[22]) );
  DFFRHQX1 y3_tmp_reg_22_ ( .D(N1315), .CK(clk), .RN(rstn), .Q(y3_tmp[22]) );
  DFFRHQX1 x5_18_reg_20_ ( .D(N534), .CK(clk), .RN(rstn), .Q(x5_18[20]) );
  DFFRHQX1 x6_18_reg_20_ ( .D(N623), .CK(clk), .RN(rstn), .Q(x6_18[20]) );
  DFFRHQX1 x4_18_reg_20_ ( .D(N445), .CK(clk), .RN(rstn), .Q(x4_18[20]) );
  DFFRHQX1 x7_tmp_reg_18_ ( .D(N1208), .CK(clk), .RN(rstn), .Q(x7_tmp[18]) );
  DFFRHQX1 x7_tmp_reg_19_ ( .D(N1209), .CK(clk), .RN(rstn), .Q(x7_tmp[19]) );
  DFFRHQX1 x7_tmp_reg_20_ ( .D(N1210), .CK(clk), .RN(rstn), .Q(x7_tmp[20]) );
  DFFRHQX1 x7_tmp_reg_21_ ( .D(N1211), .CK(clk), .RN(rstn), .Q(x7_tmp[21]) );
  DFFRHQX1 x7_tmp_reg_22_ ( .D(N1212), .CK(clk), .RN(rstn), .Q(x7_tmp[22]) );
  DFFRHQX1 x5_tmp_reg_22_ ( .D(N996), .CK(clk), .RN(rstn), .Q(x5_tmp[22]) );
  DFFRHQX1 x5_tmp_reg_21_ ( .D(N995), .CK(clk), .RN(rstn), .Q(x5_tmp[21]) );
  DFFRHQX1 x5_tmp_reg_20_ ( .D(N994), .CK(clk), .RN(rstn), .Q(x5_tmp[20]) );
  DFFRHQX1 x5_tmp_reg_19_ ( .D(N993), .CK(clk), .RN(rstn), .Q(x5_tmp[19]) );
  DFFRHQX1 x5_tmp_reg_18_ ( .D(N992), .CK(clk), .RN(rstn), .Q(x5_tmp[18]) );
  DFFRHQX1 x6_tmp_reg_22_ ( .D(N1139), .CK(clk), .RN(rstn), .Q(x6_tmp[22]) );
  DFFRHQX1 x6_tmp_reg_21_ ( .D(N1138), .CK(clk), .RN(rstn), .Q(x6_tmp[21]) );
  DFFRHQX1 x6_tmp_reg_20_ ( .D(N1137), .CK(clk), .RN(rstn), .Q(x6_tmp[20]) );
  DFFRHQX1 x6_tmp_reg_19_ ( .D(N1136), .CK(clk), .RN(rstn), .Q(x6_tmp[19]) );
  DFFRHQX1 x6_tmp_reg_18_ ( .D(N1135), .CK(clk), .RN(rstn), .Q(x6_tmp[18]) );
  DFFRHQX1 x4_tmp_reg_18_ ( .D(N872), .CK(clk), .RN(rstn), .Q(x4_tmp[18]) );
  DFFRHQX1 x4_tmp_reg_19_ ( .D(N873), .CK(clk), .RN(rstn), .Q(x4_tmp[19]) );
  DFFRHQX1 x4_tmp_reg_20_ ( .D(N874), .CK(clk), .RN(rstn), .Q(x4_tmp[20]) );
  DFFRHQX1 x4_tmp_reg_21_ ( .D(N875), .CK(clk), .RN(rstn), .Q(x4_tmp[21]) );
  DFFRHQX1 x4_tmp_reg_22_ ( .D(N876), .CK(clk), .RN(rstn), .Q(x4_tmp[22]) );
  DFFRHQX1 y6_tmp_reg_20_ ( .D(N1544), .CK(clk), .RN(rstn), .Q(y6_tmp[20]) );
  DFFRHQX1 y6_tmp_reg_19_ ( .D(N1543), .CK(clk), .RN(rstn), .Q(y6_tmp[19]) );
  DFFRHQX1 y6_tmp_reg_18_ ( .D(N1542), .CK(clk), .RN(rstn), .Q(y6_tmp[18]) );
  DFFRHQX1 y6_tmp_reg_17_ ( .D(N1541), .CK(clk), .RN(rstn), .Q(y6_tmp[17]) );
  DFFRHQX1 y6_tmp_reg_16_ ( .D(N1540), .CK(clk), .RN(rstn), .Q(y6_tmp[16]) );
  DFFRHQX1 y6_tmp_reg_15_ ( .D(N1539), .CK(clk), .RN(rstn), .Q(y6_tmp[15]) );
  DFFRHQX1 y7_tmp_reg_20_ ( .D(N1621), .CK(clk), .RN(rstn), .Q(y7_tmp[20]) );
  DFFRHQX1 y7_tmp_reg_19_ ( .D(N1620), .CK(clk), .RN(rstn), .Q(y7_tmp[19]) );
  DFFRHQX1 y7_tmp_reg_18_ ( .D(N1619), .CK(clk), .RN(rstn), .Q(y7_tmp[18]) );
  DFFRHQX1 y7_tmp_reg_17_ ( .D(N1618), .CK(clk), .RN(rstn), .Q(y7_tmp[17]) );
  DFFRHQX1 y7_tmp_reg_16_ ( .D(N1617), .CK(clk), .RN(rstn), .Q(y7_tmp[16]) );
  DFFRHQX1 y7_tmp_reg_15_ ( .D(N1616), .CK(clk), .RN(rstn), .Q(y7_tmp[15]) );
  DFFRHQX1 y0_tmp_reg_21_ ( .D(N1236), .CK(clk), .RN(rstn), .Q(y0_tmp[21]) );
  DFFRHQX1 y0_tmp_reg_20_ ( .D(N1235), .CK(clk), .RN(rstn), .Q(y0_tmp[20]) );
  DFFRHQX1 y0_tmp_reg_19_ ( .D(N1234), .CK(clk), .RN(rstn), .Q(y0_tmp[19]) );
  DFFRHQX1 y0_tmp_reg_18_ ( .D(N1233), .CK(clk), .RN(rstn), .Q(y0_tmp[18]) );
  DFFRHQX1 y0_tmp_reg_17_ ( .D(N1232), .CK(clk), .RN(rstn), .Q(y0_tmp[17]) );
  DFFRHQX1 y1_tmp_reg_21_ ( .D(N1262), .CK(clk), .RN(rstn), .Q(y1_tmp[21]) );
  DFFRHQX1 y1_tmp_reg_20_ ( .D(N1261), .CK(clk), .RN(rstn), .Q(y1_tmp[20]) );
  DFFRHQX1 y1_tmp_reg_19_ ( .D(N1260), .CK(clk), .RN(rstn), .Q(y1_tmp[19]) );
  DFFRHQX1 y1_tmp_reg_18_ ( .D(N1259), .CK(clk), .RN(rstn), .Q(y1_tmp[18]) );
  DFFRHQX1 y1_tmp_reg_17_ ( .D(N1258), .CK(clk), .RN(rstn), .Q(y1_tmp[17]) );
  DFFRHQX1 y2_tmp_reg_21_ ( .D(N1288), .CK(clk), .RN(rstn), .Q(y2_tmp[21]) );
  DFFRHQX1 y2_tmp_reg_20_ ( .D(N1287), .CK(clk), .RN(rstn), .Q(y2_tmp[20]) );
  DFFRHQX1 y2_tmp_reg_19_ ( .D(N1286), .CK(clk), .RN(rstn), .Q(y2_tmp[19]) );
  DFFRHQX1 y2_tmp_reg_18_ ( .D(N1285), .CK(clk), .RN(rstn), .Q(y2_tmp[18]) );
  DFFRHQX1 y2_tmp_reg_17_ ( .D(N1284), .CK(clk), .RN(rstn), .Q(y2_tmp[17]) );
  DFFRHQX1 y3_tmp_reg_21_ ( .D(N1314), .CK(clk), .RN(rstn), .Q(y3_tmp[21]) );
  DFFRHQX1 y3_tmp_reg_20_ ( .D(N1313), .CK(clk), .RN(rstn), .Q(y3_tmp[20]) );
  DFFRHQX1 y3_tmp_reg_19_ ( .D(N1312), .CK(clk), .RN(rstn), .Q(y3_tmp[19]) );
  DFFRHQX1 y3_tmp_reg_18_ ( .D(N1311), .CK(clk), .RN(rstn), .Q(y3_tmp[18]) );
  DFFRHQX1 y3_tmp_reg_17_ ( .D(N1310), .CK(clk), .RN(rstn), .Q(y3_tmp[17]) );
  DFFRHQX1 y4_tmp_reg_20_ ( .D(N1390), .CK(clk), .RN(rstn), .Q(y4_tmp[20]) );
  DFFRHQX1 y4_tmp_reg_19_ ( .D(N1389), .CK(clk), .RN(rstn), .Q(y4_tmp[19]) );
  DFFRHQX1 y4_tmp_reg_18_ ( .D(N1388), .CK(clk), .RN(rstn), .Q(y4_tmp[18]) );
  DFFRHQX1 y4_tmp_reg_17_ ( .D(N1387), .CK(clk), .RN(rstn), .Q(y4_tmp[17]) );
  DFFRHQX1 y4_tmp_reg_16_ ( .D(N1386), .CK(clk), .RN(rstn), .Q(y4_tmp[16]) );
  DFFRHQX1 y4_tmp_reg_15_ ( .D(N1385), .CK(clk), .RN(rstn), .Q(y4_tmp[15]) );
  DFFRHQX1 y5_tmp_reg_20_ ( .D(N1467), .CK(clk), .RN(rstn), .Q(y5_tmp[20]) );
  DFFRHQX1 y5_tmp_reg_19_ ( .D(N1466), .CK(clk), .RN(rstn), .Q(y5_tmp[19]) );
  DFFRHQX1 y5_tmp_reg_18_ ( .D(N1465), .CK(clk), .RN(rstn), .Q(y5_tmp[18]) );
  DFFRHQX1 y5_tmp_reg_17_ ( .D(N1464), .CK(clk), .RN(rstn), .Q(y5_tmp[17]) );
  DFFRHQX1 y5_tmp_reg_16_ ( .D(N1463), .CK(clk), .RN(rstn), .Q(y5_tmp[16]) );
  DFFRHQX1 y5_tmp_reg_15_ ( .D(N1462), .CK(clk), .RN(rstn), .Q(y5_tmp[15]) );
  DFFRHQX1 x4_75_tmp2_reg_19_ ( .D(N80), .CK(clk), .RN(rstn), .Q(
        x4_75_tmp2[19]) );
  DFFRHQX1 x5_75_tmp2_reg_19_ ( .D(N165), .CK(clk), .RN(rstn), .Q(
        x5_75_tmp2[19]) );
  DFFRHQX1 x6_75_tmp2_reg_19_ ( .D(N250), .CK(clk), .RN(rstn), .Q(
        x6_75_tmp2[19]) );
  DFFRHQX1 x7_75_tmp2_reg_19_ ( .D(N335), .CK(clk), .RN(rstn), .Q(
        x7_75_tmp2[19]) );
  DFFRHQX1 x7_18_reg_20_ ( .D(N712), .CK(clk), .RN(rstn), .Q(x7_18[20]) );
  DFFRHQX1 x4_18_tmp2_reg_16_ ( .D(x4[15]), .CK(clk), .RN(rstn), .Q(
        x4_18_tmp2[16]) );
  DFFRHQX1 x6_18_tmp2_reg_16_ ( .D(x6[15]), .CK(clk), .RN(rstn), .Q(
        x6_18_tmp2[16]) );
  DFFRHQX1 x5_18_tmp2_reg_16_ ( .D(x5[15]), .CK(clk), .RN(rstn), .Q(
        x5_18_tmp2[16]) );
  DFFRHQX1 x7_18_tmp2_reg_16_ ( .D(x7[15]), .CK(clk), .RN(rstn), .Q(
        x7_18_tmp2[16]) );
  DFFRHQX1 mode_delay2_reg_1_ ( .D(mode_delay1[1]), .CK(clk), .RN(rstn), .Q(
        mode_delay2[1]) );
  DFFRHQX1 x7_89_tmp1_reg_14_ ( .D(N286), .CK(clk), .RN(rstn), .Q(
        x7_89_tmp1[14]) );
  DFFRHQX1 x7_89_tmp1_reg_13_ ( .D(N285), .CK(clk), .RN(rstn), .Q(
        x7_89_tmp1[13]) );
  DFFRHQX1 x7_89_tmp1_reg_12_ ( .D(N284), .CK(clk), .RN(rstn), .Q(
        x7_89_tmp1[12]) );
  DFFRHQX1 x7_89_tmp1_reg_11_ ( .D(N283), .CK(clk), .RN(rstn), .Q(
        x7_89_tmp1[11]) );
  DFFRHQX1 x7_89_tmp1_reg_10_ ( .D(N282), .CK(clk), .RN(rstn), .Q(
        x7_89_tmp1[10]) );
  DFFRHQX1 x6_89_tmp1_reg_14_ ( .D(N201), .CK(clk), .RN(rstn), .Q(
        x6_89_tmp1[14]) );
  DFFRHQX1 x6_89_tmp1_reg_13_ ( .D(N200), .CK(clk), .RN(rstn), .Q(
        x6_89_tmp1[13]) );
  DFFRHQX1 x6_89_tmp1_reg_12_ ( .D(N199), .CK(clk), .RN(rstn), .Q(
        x6_89_tmp1[12]) );
  DFFRHQX1 x6_89_tmp1_reg_11_ ( .D(N198), .CK(clk), .RN(rstn), .Q(
        x6_89_tmp1[11]) );
  DFFRHQX1 x6_89_tmp1_reg_10_ ( .D(N197), .CK(clk), .RN(rstn), .Q(
        x6_89_tmp1[10]) );
  DFFRHQX1 x5_89_tmp1_reg_14_ ( .D(N116), .CK(clk), .RN(rstn), .Q(
        x5_89_tmp1[14]) );
  DFFRHQX1 x5_89_tmp1_reg_13_ ( .D(N115), .CK(clk), .RN(rstn), .Q(
        x5_89_tmp1[13]) );
  DFFRHQX1 x5_89_tmp1_reg_12_ ( .D(N114), .CK(clk), .RN(rstn), .Q(
        x5_89_tmp1[12]) );
  DFFRHQX1 x5_89_tmp1_reg_11_ ( .D(N113), .CK(clk), .RN(rstn), .Q(
        x5_89_tmp1[11]) );
  DFFRHQX1 x5_89_tmp1_reg_10_ ( .D(N112), .CK(clk), .RN(rstn), .Q(
        x5_89_tmp1[10]) );
  DFFRHQX1 x5_75_tmp1_reg_14_ ( .D(N116), .CK(clk), .RN(rstn), .Q(
        x5_75_tmp1[14]) );
  DFFRHQX1 x5_75_tmp1_reg_13_ ( .D(N115), .CK(clk), .RN(rstn), .Q(
        x5_75_tmp1[13]) );
  DFFRHQX1 x5_75_tmp1_reg_12_ ( .D(N114), .CK(clk), .RN(rstn), .Q(
        x5_75_tmp1[12]) );
  DFFRHQX1 x5_75_tmp1_reg_11_ ( .D(N113), .CK(clk), .RN(rstn), .Q(
        x5_75_tmp1[11]) );
  DFFRHQX1 x5_75_tmp1_reg_10_ ( .D(N112), .CK(clk), .RN(rstn), .Q(
        x5_75_tmp1[10]) );
  DFFRHQX1 x4_75_tmp1_reg_14_ ( .D(N31), .CK(clk), .RN(rstn), .Q(
        x4_75_tmp1[14]) );
  DFFRHQX1 x4_75_tmp1_reg_13_ ( .D(N30), .CK(clk), .RN(rstn), .Q(
        x4_75_tmp1[13]) );
  DFFRHQX1 x4_75_tmp1_reg_12_ ( .D(N29), .CK(clk), .RN(rstn), .Q(
        x4_75_tmp1[12]) );
  DFFRHQX1 x4_75_tmp1_reg_11_ ( .D(N28), .CK(clk), .RN(rstn), .Q(
        x4_75_tmp1[11]) );
  DFFRHQX1 x4_75_tmp1_reg_10_ ( .D(N27), .CK(clk), .RN(rstn), .Q(
        x4_75_tmp1[10]) );
  DFFRHQX1 x7_75_tmp1_reg_14_ ( .D(N286), .CK(clk), .RN(rstn), .Q(
        x7_75_tmp1[14]) );
  DFFRHQX1 x7_75_tmp1_reg_13_ ( .D(N285), .CK(clk), .RN(rstn), .Q(
        x7_75_tmp1[13]) );
  DFFRHQX1 x7_75_tmp1_reg_12_ ( .D(N284), .CK(clk), .RN(rstn), .Q(
        x7_75_tmp1[12]) );
  DFFRHQX1 x7_75_tmp1_reg_11_ ( .D(N283), .CK(clk), .RN(rstn), .Q(
        x7_75_tmp1[11]) );
  DFFRHQX1 x7_75_tmp1_reg_10_ ( .D(N282), .CK(clk), .RN(rstn), .Q(
        x7_75_tmp1[10]) );
  DFFRHQX1 x6_75_tmp1_reg_14_ ( .D(N201), .CK(clk), .RN(rstn), .Q(
        x6_75_tmp1[14]) );
  DFFRHQX1 x6_75_tmp1_reg_13_ ( .D(N200), .CK(clk), .RN(rstn), .Q(
        x6_75_tmp1[13]) );
  DFFRHQX1 x6_75_tmp1_reg_12_ ( .D(N199), .CK(clk), .RN(rstn), .Q(
        x6_75_tmp1[12]) );
  DFFRHQX1 x6_75_tmp1_reg_11_ ( .D(N198), .CK(clk), .RN(rstn), .Q(
        x6_75_tmp1[11]) );
  DFFRHQX1 x6_75_tmp1_reg_10_ ( .D(N197), .CK(clk), .RN(rstn), .Q(
        x6_75_tmp1[10]) );
  DFFRHQX1 x4_50_tmp1_reg_13_ ( .D(n82), .CK(clk), .RN(rstn), .Q(
        x4_50_tmp1[13]) );
  DFFRHQX1 x4_50_tmp1_reg_12_ ( .D(n81), .CK(clk), .RN(rstn), .Q(
        x4_50_tmp1[12]) );
  DFFRHQX1 x4_50_tmp1_reg_11_ ( .D(n80), .CK(clk), .RN(rstn), .Q(
        x4_50_tmp1[11]) );
  DFFRHQX1 x4_50_tmp1_reg_10_ ( .D(n79), .CK(clk), .RN(rstn), .Q(
        x4_50_tmp1[10]) );
  DFFRHQX1 x4_50_tmp1_reg_9_ ( .D(n78), .CK(clk), .RN(rstn), .Q(x4_50_tmp1[9])
         );
  DFFRHQX1 x6_50_tmp1_reg_13_ ( .D(n56), .CK(clk), .RN(rstn), .Q(
        x6_50_tmp1[13]) );
  DFFRHQX1 x6_50_tmp1_reg_12_ ( .D(n55), .CK(clk), .RN(rstn), .Q(
        x6_50_tmp1[12]) );
  DFFRHQX1 x6_50_tmp1_reg_11_ ( .D(n54), .CK(clk), .RN(rstn), .Q(
        x6_50_tmp1[11]) );
  DFFRHQX1 x6_50_tmp1_reg_10_ ( .D(n53), .CK(clk), .RN(rstn), .Q(
        x6_50_tmp1[10]) );
  DFFRHQX1 x6_50_tmp1_reg_9_ ( .D(n52), .CK(clk), .RN(rstn), .Q(x6_50_tmp1[9])
         );
  DFFRHQX1 x5_50_tmp1_reg_13_ ( .D(n69), .CK(clk), .RN(rstn), .Q(
        x5_50_tmp1[13]) );
  DFFRHQX1 x5_50_tmp1_reg_12_ ( .D(n68), .CK(clk), .RN(rstn), .Q(
        x5_50_tmp1[12]) );
  DFFRHQX1 x5_50_tmp1_reg_11_ ( .D(n67), .CK(clk), .RN(rstn), .Q(
        x5_50_tmp1[11]) );
  DFFRHQX1 x5_50_tmp1_reg_10_ ( .D(n66), .CK(clk), .RN(rstn), .Q(
        x5_50_tmp1[10]) );
  DFFRHQX1 x5_50_tmp1_reg_9_ ( .D(n65), .CK(clk), .RN(rstn), .Q(x5_50_tmp1[9])
         );
  DFFRHQX1 x7_50_tmp1_reg_13_ ( .D(n43), .CK(clk), .RN(rstn), .Q(
        x7_50_tmp1[13]) );
  DFFRHQX1 x7_50_tmp1_reg_12_ ( .D(n42), .CK(clk), .RN(rstn), .Q(
        x7_50_tmp1[12]) );
  DFFRHQX1 x7_50_tmp1_reg_11_ ( .D(n41), .CK(clk), .RN(rstn), .Q(
        x7_50_tmp1[11]) );
  DFFRHQX1 x7_50_tmp1_reg_10_ ( .D(n40), .CK(clk), .RN(rstn), .Q(
        x7_50_tmp1[10]) );
  DFFRHQX1 x7_50_tmp1_reg_9_ ( .D(n39), .CK(clk), .RN(rstn), .Q(x7_50_tmp1[9])
         );
  DFFRHQX1 x4_18_tmp1_reg_12_ ( .D(n82), .CK(clk), .RN(rstn), .Q(
        x4_18_tmp1[12]) );
  DFFRHQX1 x4_18_tmp1_reg_11_ ( .D(n81), .CK(clk), .RN(rstn), .Q(
        x4_18_tmp1[11]) );
  DFFRHQX1 x4_18_tmp1_reg_10_ ( .D(n80), .CK(clk), .RN(rstn), .Q(
        x4_18_tmp1[10]) );
  DFFRHQX1 x4_18_tmp1_reg_9_ ( .D(n79), .CK(clk), .RN(rstn), .Q(x4_18_tmp1[9])
         );
  DFFRHQX1 x4_18_tmp1_reg_8_ ( .D(n78), .CK(clk), .RN(rstn), .Q(x4_18_tmp1[8])
         );
  DFFRHQX1 x5_18_tmp1_reg_12_ ( .D(n69), .CK(clk), .RN(rstn), .Q(
        x5_18_tmp1[12]) );
  DFFRHQX1 x5_18_tmp1_reg_11_ ( .D(n68), .CK(clk), .RN(rstn), .Q(
        x5_18_tmp1[11]) );
  DFFRHQX1 x5_18_tmp1_reg_10_ ( .D(n67), .CK(clk), .RN(rstn), .Q(
        x5_18_tmp1[10]) );
  DFFRHQX1 x5_18_tmp1_reg_9_ ( .D(n66), .CK(clk), .RN(rstn), .Q(x5_18_tmp1[9])
         );
  DFFRHQX1 x5_18_tmp1_reg_8_ ( .D(n65), .CK(clk), .RN(rstn), .Q(x5_18_tmp1[8])
         );
  DFFRHQX1 x6_18_tmp1_reg_12_ ( .D(n56), .CK(clk), .RN(rstn), .Q(
        x6_18_tmp1[12]) );
  DFFRHQX1 x6_18_tmp1_reg_11_ ( .D(n55), .CK(clk), .RN(rstn), .Q(
        x6_18_tmp1[11]) );
  DFFRHQX1 x6_18_tmp1_reg_10_ ( .D(n54), .CK(clk), .RN(rstn), .Q(
        x6_18_tmp1[10]) );
  DFFRHQX1 x6_18_tmp1_reg_9_ ( .D(n53), .CK(clk), .RN(rstn), .Q(x6_18_tmp1[9])
         );
  DFFRHQX1 x6_18_tmp1_reg_8_ ( .D(n52), .CK(clk), .RN(rstn), .Q(x6_18_tmp1[8])
         );
  DFFRHQX1 x7_18_tmp1_reg_12_ ( .D(n43), .CK(clk), .RN(rstn), .Q(
        x7_18_tmp1[12]) );
  DFFRHQX1 x7_18_tmp1_reg_11_ ( .D(n42), .CK(clk), .RN(rstn), .Q(
        x7_18_tmp1[11]) );
  DFFRHQX1 x7_18_tmp1_reg_10_ ( .D(n41), .CK(clk), .RN(rstn), .Q(
        x7_18_tmp1[10]) );
  DFFRHQX1 x7_18_tmp1_reg_9_ ( .D(n40), .CK(clk), .RN(rstn), .Q(x7_18_tmp1[9])
         );
  DFFRHQX1 x7_18_tmp1_reg_8_ ( .D(n39), .CK(clk), .RN(rstn), .Q(x7_18_tmp1[8])
         );
  DFFRHQX1 x5_18_reg_16_ ( .D(N530), .CK(clk), .RN(rstn), .Q(x5_18[16]) );
  DFFRHQX1 x5_18_reg_15_ ( .D(N529), .CK(clk), .RN(rstn), .Q(x5_18[15]) );
  DFFRHQX1 x5_18_reg_14_ ( .D(N528), .CK(clk), .RN(rstn), .Q(x5_18[14]) );
  DFFRHQX1 x5_18_reg_13_ ( .D(N527), .CK(clk), .RN(rstn), .Q(x5_18[13]) );
  DFFRHQX1 x6_18_reg_15_ ( .D(N618), .CK(clk), .RN(rstn), .Q(x6_18[15]) );
  DFFRHQX1 x6_18_reg_14_ ( .D(N617), .CK(clk), .RN(rstn), .Q(x6_18[14]) );
  DFFRHQX1 x6_18_reg_13_ ( .D(N616), .CK(clk), .RN(rstn), .Q(x6_18[13]) );
  DFFRHQX1 x6_18_reg_12_ ( .D(N615), .CK(clk), .RN(rstn), .Q(x6_18[12]) );
  DFFRHQX1 x6_18_reg_11_ ( .D(N614), .CK(clk), .RN(rstn), .Q(x6_18[11]) );
  DFFRHQX1 x4_18_reg_15_ ( .D(N440), .CK(clk), .RN(rstn), .Q(x4_18[15]) );
  DFFRHQX1 x4_18_reg_14_ ( .D(N439), .CK(clk), .RN(rstn), .Q(x4_18[14]) );
  DFFRHQX1 x4_18_reg_13_ ( .D(N438), .CK(clk), .RN(rstn), .Q(x4_18[13]) );
  DFFRHQX1 x4_18_reg_12_ ( .D(N437), .CK(clk), .RN(rstn), .Q(x4_18[12]) );
  DFFRHQX1 x4_18_reg_11_ ( .D(N436), .CK(clk), .RN(rstn), .Q(x4_18[11]) );
  DFFRHQX1 x4_89_tmp1_reg_14_ ( .D(N31), .CK(clk), .RN(rstn), .Q(
        x4_89_tmp1[14]) );
  DFFRHQX1 x4_89_tmp1_reg_13_ ( .D(N30), .CK(clk), .RN(rstn), .Q(
        x4_89_tmp1[13]) );
  DFFRHQX1 x4_89_tmp1_reg_12_ ( .D(N29), .CK(clk), .RN(rstn), .Q(
        x4_89_tmp1[12]) );
  DFFRHQX1 x4_89_tmp1_reg_11_ ( .D(N28), .CK(clk), .RN(rstn), .Q(
        x4_89_tmp1[11]) );
  DFFRHQX1 x4_89_tmp1_reg_10_ ( .D(N27), .CK(clk), .RN(rstn), .Q(
        x4_89_tmp1[10]) );
  DFFRHQX1 x4_89_reg_15_ ( .D(N372), .CK(clk), .RN(rstn), .Q(x4_89[15]) );
  DFFRHQX1 x4_89_reg_14_ ( .D(N371), .CK(clk), .RN(rstn), .Q(x4_89[14]) );
  DFFRHQX1 x4_89_reg_13_ ( .D(N370), .CK(clk), .RN(rstn), .Q(x4_89[13]) );
  DFFRHQX1 x4_89_reg_12_ ( .D(N369), .CK(clk), .RN(rstn), .Q(x4_89[12]) );
  DFFRHQX1 x4_89_reg_11_ ( .D(N368), .CK(clk), .RN(rstn), .Q(x4_89[11]) );
  DFFRHQX1 x4_75_reg_15_ ( .D(N395), .CK(clk), .RN(rstn), .Q(x4_75[15]) );
  DFFRHQX1 x4_75_reg_14_ ( .D(N394), .CK(clk), .RN(rstn), .Q(x4_75[14]) );
  DFFRHQX1 x4_75_reg_13_ ( .D(N393), .CK(clk), .RN(rstn), .Q(x4_75[13]) );
  DFFRHQX1 x4_75_reg_12_ ( .D(N392), .CK(clk), .RN(rstn), .Q(x4_75[12]) );
  DFFRHQX1 x4_75_reg_11_ ( .D(N391), .CK(clk), .RN(rstn), .Q(x4_75[11]) );
  DFFRHQX1 x5_75_reg_15_ ( .D(N484), .CK(clk), .RN(rstn), .Q(x5_75[15]) );
  DFFRHQX1 x5_75_reg_14_ ( .D(N483), .CK(clk), .RN(rstn), .Q(x5_75[14]) );
  DFFRHQX1 x5_75_reg_13_ ( .D(N482), .CK(clk), .RN(rstn), .Q(x5_75[13]) );
  DFFRHQX1 x5_75_reg_12_ ( .D(N481), .CK(clk), .RN(rstn), .Q(x5_75[12]) );
  DFFRHQX1 x5_75_reg_11_ ( .D(N480), .CK(clk), .RN(rstn), .Q(x5_75[11]) );
  DFFRHQX1 x6_75_reg_15_ ( .D(N573), .CK(clk), .RN(rstn), .Q(x6_75[15]) );
  DFFRHQX1 x6_75_reg_14_ ( .D(N572), .CK(clk), .RN(rstn), .Q(x6_75[14]) );
  DFFRHQX1 x6_75_reg_13_ ( .D(N571), .CK(clk), .RN(rstn), .Q(x6_75[13]) );
  DFFRHQX1 x6_75_reg_12_ ( .D(N570), .CK(clk), .RN(rstn), .Q(x6_75[12]) );
  DFFRHQX1 x6_75_reg_11_ ( .D(N569), .CK(clk), .RN(rstn), .Q(x6_75[11]) );
  DFFRHQX1 x4_50_reg_15_ ( .D(N418), .CK(clk), .RN(rstn), .Q(x4_50[15]) );
  DFFRHQX1 x4_50_reg_14_ ( .D(N417), .CK(clk), .RN(rstn), .Q(x4_50[14]) );
  DFFRHQX1 x4_50_reg_13_ ( .D(N416), .CK(clk), .RN(rstn), .Q(x4_50[13]) );
  DFFRHQX1 x4_50_reg_12_ ( .D(N415), .CK(clk), .RN(rstn), .Q(x4_50[12]) );
  DFFRHQX1 x4_50_reg_11_ ( .D(N414), .CK(clk), .RN(rstn), .Q(x4_50[11]) );
  DFFRHQX1 x5_tmp1_reg_16_ ( .D(N895), .CK(clk), .RN(rstn), .Q(x5_tmp1[16]) );
  DFFRHQX1 x5_tmp1_reg_15_ ( .D(N894), .CK(clk), .RN(rstn), .Q(x5_tmp1[15]) );
  DFFRHQX1 x5_tmp1_reg_14_ ( .D(N893), .CK(clk), .RN(rstn), .Q(x5_tmp1[14]) );
  DFFRHQX1 x5_tmp1_reg_13_ ( .D(N892), .CK(clk), .RN(rstn), .Q(x5_tmp1[13]) );
  DFFRHQX1 x5_tmp1_reg_12_ ( .D(N891), .CK(clk), .RN(rstn), .Q(x5_tmp1[12]) );
  DFFRHQX1 x6_tmp1_reg_16_ ( .D(N1061), .CK(clk), .RN(rstn), .Q(x6_tmp1[16])
         );
  DFFRHQX1 x6_tmp1_reg_15_ ( .D(N1060), .CK(clk), .RN(rstn), .Q(x6_tmp1[15])
         );
  DFFRHQX1 x6_tmp1_reg_14_ ( .D(N1059), .CK(clk), .RN(rstn), .Q(x6_tmp1[14])
         );
  DFFRHQX1 x6_tmp1_reg_13_ ( .D(N1058), .CK(clk), .RN(rstn), .Q(x6_tmp1[13])
         );
  DFFRHQX1 x6_tmp1_reg_12_ ( .D(N1057), .CK(clk), .RN(rstn), .Q(x6_tmp1[12])
         );
  DFFRHQX1 x7_tmp1_reg_16_ ( .D(N1158), .CK(clk), .RN(rstn), .Q(x7_tmp1[16])
         );
  DFFRHQX1 x7_tmp1_reg_15_ ( .D(N1157), .CK(clk), .RN(rstn), .Q(x7_tmp1[15])
         );
  DFFRHQX1 x7_tmp1_reg_14_ ( .D(N1156), .CK(clk), .RN(rstn), .Q(x7_tmp1[14])
         );
  DFFRHQX1 x7_tmp1_reg_13_ ( .D(N1155), .CK(clk), .RN(rstn), .Q(x7_tmp1[13])
         );
  DFFRHQX1 x7_tmp1_reg_12_ ( .D(N1154), .CK(clk), .RN(rstn), .Q(x7_tmp1[12])
         );
  DFFRHQX1 x4_tmp1_reg_16_ ( .D(N776), .CK(clk), .RN(rstn), .Q(x4_tmp1[16]) );
  DFFRHQX1 x4_tmp1_reg_15_ ( .D(N775), .CK(clk), .RN(rstn), .Q(x4_tmp1[15]) );
  DFFRHQX1 x4_tmp1_reg_14_ ( .D(N774), .CK(clk), .RN(rstn), .Q(x4_tmp1[14]) );
  DFFRHQX1 x4_tmp1_reg_13_ ( .D(N773), .CK(clk), .RN(rstn), .Q(x4_tmp1[13]) );
  DFFRHQX1 x4_tmp1_reg_12_ ( .D(N772), .CK(clk), .RN(rstn), .Q(x4_tmp1[12]) );
  DFFRHQX1 mode_delay2_reg_0_ ( .D(mode_delay1[0]), .CK(clk), .RN(rstn), .Q(
        mode_delay2[0]) );
  DFFRHQX1 x7_50_reg_15_ ( .D(N685), .CK(clk), .RN(rstn), .Q(x7_50[15]) );
  DFFRHQX1 x7_50_reg_14_ ( .D(N684), .CK(clk), .RN(rstn), .Q(x7_50[14]) );
  DFFRHQX1 x7_50_reg_13_ ( .D(N683), .CK(clk), .RN(rstn), .Q(x7_50[13]) );
  DFFRHQX1 x7_50_reg_12_ ( .D(N682), .CK(clk), .RN(rstn), .Q(x7_50[12]) );
  DFFRHQX1 x5_89_reg_15_ ( .D(N461), .CK(clk), .RN(rstn), .Q(x5_89[15]) );
  DFFRHQX1 x5_89_reg_14_ ( .D(N460), .CK(clk), .RN(rstn), .Q(x5_89[14]) );
  DFFRHQX1 x5_89_reg_13_ ( .D(N459), .CK(clk), .RN(rstn), .Q(x5_89[13]) );
  DFFRHQX1 x5_89_reg_12_ ( .D(N458), .CK(clk), .RN(rstn), .Q(x5_89[12]) );
  DFFRHQX1 x7_89_reg_15_ ( .D(N639), .CK(clk), .RN(rstn), .Q(x7_89[15]) );
  DFFRHQX1 x7_89_reg_14_ ( .D(N638), .CK(clk), .RN(rstn), .Q(x7_89[14]) );
  DFFRHQX1 x7_89_reg_13_ ( .D(N637), .CK(clk), .RN(rstn), .Q(x7_89[13]) );
  DFFRHQX1 x7_89_reg_12_ ( .D(N636), .CK(clk), .RN(rstn), .Q(x7_89[12]) );
  DFFRHQX1 x5_50_reg_15_ ( .D(N507), .CK(clk), .RN(rstn), .Q(x5_50[15]) );
  DFFRHQX1 x5_50_reg_14_ ( .D(N506), .CK(clk), .RN(rstn), .Q(x5_50[14]) );
  DFFRHQX1 x5_50_reg_13_ ( .D(N505), .CK(clk), .RN(rstn), .Q(x5_50[13]) );
  DFFRHQX1 x5_50_reg_12_ ( .D(N504), .CK(clk), .RN(rstn), .Q(x5_50[12]) );
  DFFRHQX1 x6_89_tmp2_reg_13_ ( .D(N223), .CK(clk), .RN(rstn), .Q(
        x6_89_tmp2[13]) );
  DFFRHQX1 x6_89_tmp2_reg_12_ ( .D(N222), .CK(clk), .RN(rstn), .Q(
        x6_89_tmp2[12]) );
  DFFRHQX1 x6_89_tmp2_reg_11_ ( .D(N221), .CK(clk), .RN(rstn), .Q(
        x6_89_tmp2[11]) );
  DFFRHQX1 x6_89_tmp2_reg_10_ ( .D(N220), .CK(clk), .RN(rstn), .Q(
        x6_89_tmp2[10]) );
  DFFRHQX1 x5_89_tmp2_reg_13_ ( .D(N138), .CK(clk), .RN(rstn), .Q(
        x5_89_tmp2[13]) );
  DFFRHQX1 x5_89_tmp2_reg_12_ ( .D(N137), .CK(clk), .RN(rstn), .Q(
        x5_89_tmp2[12]) );
  DFFRHQX1 x5_89_tmp2_reg_11_ ( .D(N136), .CK(clk), .RN(rstn), .Q(
        x5_89_tmp2[11]) );
  DFFRHQX1 x5_89_tmp2_reg_10_ ( .D(N135), .CK(clk), .RN(rstn), .Q(
        x5_89_tmp2[10]) );
  DFFRHQX1 x4_89_tmp2_reg_13_ ( .D(N53), .CK(clk), .RN(rstn), .Q(
        x4_89_tmp2[13]) );
  DFFRHQX1 x4_89_tmp2_reg_12_ ( .D(N52), .CK(clk), .RN(rstn), .Q(
        x4_89_tmp2[12]) );
  DFFRHQX1 x4_89_tmp2_reg_11_ ( .D(N51), .CK(clk), .RN(rstn), .Q(
        x4_89_tmp2[11]) );
  DFFRHQX1 x4_89_tmp2_reg_10_ ( .D(N50), .CK(clk), .RN(rstn), .Q(
        x4_89_tmp2[10]) );
  DFFRHQX1 x7_89_tmp2_reg_13_ ( .D(N308), .CK(clk), .RN(rstn), .Q(
        x7_89_tmp2[13]) );
  DFFRHQX1 x7_89_tmp2_reg_12_ ( .D(N307), .CK(clk), .RN(rstn), .Q(
        x7_89_tmp2[12]) );
  DFFRHQX1 x7_89_tmp2_reg_11_ ( .D(N306), .CK(clk), .RN(rstn), .Q(
        x7_89_tmp2[11]) );
  DFFRHQX1 x7_89_tmp2_reg_10_ ( .D(N305), .CK(clk), .RN(rstn), .Q(
        x7_89_tmp2[10]) );
  DFFRHQX1 x4_75_tmp2_reg_13_ ( .D(N74), .CK(clk), .RN(rstn), .Q(
        x4_75_tmp2[13]) );
  DFFRHQX1 x4_75_tmp2_reg_12_ ( .D(N73), .CK(clk), .RN(rstn), .Q(
        x4_75_tmp2[12]) );
  DFFRHQX1 x4_75_tmp2_reg_11_ ( .D(N72), .CK(clk), .RN(rstn), .Q(
        x4_75_tmp2[11]) );
  DFFRHQX1 x4_75_tmp2_reg_10_ ( .D(N71), .CK(clk), .RN(rstn), .Q(
        x4_75_tmp2[10]) );
  DFFRHQX1 x5_75_tmp2_reg_13_ ( .D(N159), .CK(clk), .RN(rstn), .Q(
        x5_75_tmp2[13]) );
  DFFRHQX1 x5_75_tmp2_reg_12_ ( .D(N158), .CK(clk), .RN(rstn), .Q(
        x5_75_tmp2[12]) );
  DFFRHQX1 x5_75_tmp2_reg_11_ ( .D(N157), .CK(clk), .RN(rstn), .Q(
        x5_75_tmp2[11]) );
  DFFRHQX1 x5_75_tmp2_reg_10_ ( .D(N156), .CK(clk), .RN(rstn), .Q(
        x5_75_tmp2[10]) );
  DFFRHQX1 x6_75_tmp2_reg_13_ ( .D(N244), .CK(clk), .RN(rstn), .Q(
        x6_75_tmp2[13]) );
  DFFRHQX1 x6_75_tmp2_reg_12_ ( .D(N243), .CK(clk), .RN(rstn), .Q(
        x6_75_tmp2[12]) );
  DFFRHQX1 x6_75_tmp2_reg_11_ ( .D(N242), .CK(clk), .RN(rstn), .Q(
        x6_75_tmp2[11]) );
  DFFRHQX1 x6_75_tmp2_reg_10_ ( .D(N241), .CK(clk), .RN(rstn), .Q(
        x6_75_tmp2[10]) );
  DFFRHQX1 x7_75_tmp2_reg_13_ ( .D(N329), .CK(clk), .RN(rstn), .Q(
        x7_75_tmp2[13]) );
  DFFRHQX1 x7_75_tmp2_reg_12_ ( .D(N328), .CK(clk), .RN(rstn), .Q(
        x7_75_tmp2[12]) );
  DFFRHQX1 x7_75_tmp2_reg_11_ ( .D(N327), .CK(clk), .RN(rstn), .Q(
        x7_75_tmp2[11]) );
  DFFRHQX1 x7_75_tmp2_reg_10_ ( .D(N326), .CK(clk), .RN(rstn), .Q(
        x7_75_tmp2[10]) );
  DFFRHQX1 x4_50_tmp2_reg_12_ ( .D(N93), .CK(clk), .RN(rstn), .Q(
        x4_50_tmp2[12]) );
  DFFRHQX1 x4_50_tmp2_reg_11_ ( .D(N92), .CK(clk), .RN(rstn), .Q(
        x4_50_tmp2[11]) );
  DFFRHQX1 x4_50_tmp2_reg_10_ ( .D(N91), .CK(clk), .RN(rstn), .Q(
        x4_50_tmp2[10]) );
  DFFRHQX1 x4_50_tmp2_reg_9_ ( .D(N90), .CK(clk), .RN(rstn), .Q(x4_50_tmp2[9])
         );
  DFFRHQX1 x6_50_tmp2_reg_12_ ( .D(N263), .CK(clk), .RN(rstn), .Q(
        x6_50_tmp2[12]) );
  DFFRHQX1 x6_50_tmp2_reg_11_ ( .D(N262), .CK(clk), .RN(rstn), .Q(
        x6_50_tmp2[11]) );
  DFFRHQX1 x6_50_tmp2_reg_10_ ( .D(N261), .CK(clk), .RN(rstn), .Q(
        x6_50_tmp2[10]) );
  DFFRHQX1 x6_50_tmp2_reg_9_ ( .D(N260), .CK(clk), .RN(rstn), .Q(x6_50_tmp2[9]) );
  DFFRHQX1 x6_50_reg_11_ ( .D(N592), .CK(clk), .RN(rstn), .Q(x6_50[11]) );
  DFFRHQX1 x6_50_reg_12_ ( .D(N593), .CK(clk), .RN(rstn), .Q(x6_50[12]) );
  DFFRHQX1 x6_50_reg_13_ ( .D(N594), .CK(clk), .RN(rstn), .Q(x6_50[13]) );
  DFFRHQX1 x6_50_reg_14_ ( .D(N595), .CK(clk), .RN(rstn), .Q(x6_50[14]) );
  DFFRHQX1 x5_50_tmp2_reg_12_ ( .D(N178), .CK(clk), .RN(rstn), .Q(
        x5_50_tmp2[12]) );
  DFFRHQX1 x5_50_tmp2_reg_11_ ( .D(N177), .CK(clk), .RN(rstn), .Q(
        x5_50_tmp2[11]) );
  DFFRHQX1 x5_50_tmp2_reg_10_ ( .D(N176), .CK(clk), .RN(rstn), .Q(
        x5_50_tmp2[10]) );
  DFFRHQX1 x5_50_tmp2_reg_9_ ( .D(N175), .CK(clk), .RN(rstn), .Q(x5_50_tmp2[9]) );
  DFFRHQX1 x7_50_tmp2_reg_12_ ( .D(N348), .CK(clk), .RN(rstn), .Q(
        x7_50_tmp2[12]) );
  DFFRHQX1 x7_50_tmp2_reg_11_ ( .D(N347), .CK(clk), .RN(rstn), .Q(
        x7_50_tmp2[11]) );
  DFFRHQX1 x7_50_tmp2_reg_10_ ( .D(N346), .CK(clk), .RN(rstn), .Q(
        x7_50_tmp2[10]) );
  DFFRHQX1 x7_50_tmp2_reg_9_ ( .D(N345), .CK(clk), .RN(rstn), .Q(x7_50_tmp2[9]) );
  DFFRHQX1 x4_18_tmp2_reg_11_ ( .D(n84), .CK(clk), .RN(rstn), .Q(
        x4_18_tmp2[11]) );
  DFFRHQX1 x4_18_tmp2_reg_10_ ( .D(n83), .CK(clk), .RN(rstn), .Q(
        x4_18_tmp2[10]) );
  DFFRHQX1 x4_18_tmp2_reg_9_ ( .D(n82), .CK(clk), .RN(rstn), .Q(x4_18_tmp2[9])
         );
  DFFRHQX1 x4_18_tmp2_reg_8_ ( .D(n81), .CK(clk), .RN(rstn), .Q(x4_18_tmp2[8])
         );
  DFFRHQX1 x6_18_tmp2_reg_11_ ( .D(n58), .CK(clk), .RN(rstn), .Q(
        x6_18_tmp2[11]) );
  DFFRHQX1 x6_18_tmp2_reg_10_ ( .D(n57), .CK(clk), .RN(rstn), .Q(
        x6_18_tmp2[10]) );
  DFFRHQX1 x6_18_tmp2_reg_9_ ( .D(n56), .CK(clk), .RN(rstn), .Q(x6_18_tmp2[9])
         );
  DFFRHQX1 x6_18_tmp2_reg_8_ ( .D(n55), .CK(clk), .RN(rstn), .Q(x6_18_tmp2[8])
         );
  DFFRHQX1 x5_18_tmp2_reg_11_ ( .D(n71), .CK(clk), .RN(rstn), .Q(
        x5_18_tmp2[11]) );
  DFFRHQX1 x5_18_tmp2_reg_10_ ( .D(n70), .CK(clk), .RN(rstn), .Q(
        x5_18_tmp2[10]) );
  DFFRHQX1 x5_18_tmp2_reg_9_ ( .D(n69), .CK(clk), .RN(rstn), .Q(x5_18_tmp2[9])
         );
  DFFRHQX1 x5_18_tmp2_reg_8_ ( .D(n68), .CK(clk), .RN(rstn), .Q(x5_18_tmp2[8])
         );
  DFFRHQX1 x7_18_tmp2_reg_11_ ( .D(n45), .CK(clk), .RN(rstn), .Q(
        x7_18_tmp2[11]) );
  DFFRHQX1 x7_18_tmp2_reg_10_ ( .D(n44), .CK(clk), .RN(rstn), .Q(
        x7_18_tmp2[10]) );
  DFFRHQX1 x7_18_tmp2_reg_9_ ( .D(n43), .CK(clk), .RN(rstn), .Q(x7_18_tmp2[9])
         );
  DFFRHQX1 x7_18_tmp2_reg_8_ ( .D(n42), .CK(clk), .RN(rstn), .Q(x7_18_tmp2[8])
         );
  DFFRHQX1 x7_18_reg_14_ ( .D(N706), .CK(clk), .RN(rstn), .Q(x7_18[14]) );
  DFFRHQX1 x7_18_reg_13_ ( .D(N705), .CK(clk), .RN(rstn), .Q(x7_18[13]) );
  DFFRHQX1 x7_18_reg_12_ ( .D(N704), .CK(clk), .RN(rstn), .Q(x7_18[12]) );
  DFFRHQX1 x7_18_reg_11_ ( .D(N703), .CK(clk), .RN(rstn), .Q(x7_18[11]) );
  DFFRHQX1 x6_89_reg_16_ ( .D(N551), .CK(clk), .RN(rstn), .Q(x6_89[16]) );
  DFFRHQX1 x6_89_reg_15_ ( .D(N550), .CK(clk), .RN(rstn), .Q(x6_89[15]) );
  DFFRHQX1 x6_89_reg_14_ ( .D(N549), .CK(clk), .RN(rstn), .Q(x6_89[14]) );
  DFFRHQX1 x6_89_reg_13_ ( .D(N548), .CK(clk), .RN(rstn), .Q(x6_89[13]) );
  DFFRHQX1 x6_89_reg_12_ ( .D(N547), .CK(clk), .RN(rstn), .Q(x6_89[12]) );
  DFFRHQX1 x7_75_reg_14_ ( .D(N661), .CK(clk), .RN(rstn), .Q(x7_75[14]) );
  DFFRHQX1 x7_75_reg_13_ ( .D(N660), .CK(clk), .RN(rstn), .Q(x7_75[13]) );
  DFFRHQX1 x7_75_reg_12_ ( .D(N659), .CK(clk), .RN(rstn), .Q(x7_75[12]) );
  DFFRHQX1 x7_75_reg_11_ ( .D(N658), .CK(clk), .RN(rstn), .Q(x7_75[11]) );
  DFFRHQX1 x4_tmp2_reg_15_ ( .D(N845), .CK(clk), .RN(rstn), .Q(x4_tmp2[15]) );
  DFFRHQX1 x4_tmp2_reg_14_ ( .D(N844), .CK(clk), .RN(rstn), .Q(x4_tmp2[14]) );
  DFFRHQX1 x4_tmp2_reg_13_ ( .D(N843), .CK(clk), .RN(rstn), .Q(x4_tmp2[13]) );
  DFFRHQX1 x4_tmp2_reg_12_ ( .D(N842), .CK(clk), .RN(rstn), .Q(x4_tmp2[12]) );
  DFFRHQX1 x5_tmp2_reg_15_ ( .D(N965), .CK(clk), .RN(rstn), .Q(x5_tmp2[15]) );
  DFFRHQX1 x5_tmp2_reg_14_ ( .D(N964), .CK(clk), .RN(rstn), .Q(x5_tmp2[14]) );
  DFFRHQX1 x5_tmp2_reg_13_ ( .D(N963), .CK(clk), .RN(rstn), .Q(x5_tmp2[13]) );
  DFFRHQX1 x5_tmp2_reg_12_ ( .D(N962), .CK(clk), .RN(rstn), .Q(x5_tmp2[12]) );
  DFFRHQX1 x6_tmp2_reg_15_ ( .D(N1108), .CK(clk), .RN(rstn), .Q(x6_tmp2[15])
         );
  DFFRHQX1 x6_tmp2_reg_14_ ( .D(N1107), .CK(clk), .RN(rstn), .Q(x6_tmp2[14])
         );
  DFFRHQX1 x6_tmp2_reg_13_ ( .D(N1106), .CK(clk), .RN(rstn), .Q(x6_tmp2[13])
         );
  DFFRHQX1 x6_tmp2_reg_12_ ( .D(N1105), .CK(clk), .RN(rstn), .Q(x6_tmp2[12])
         );
  DFFRHQX1 x7_tmp2_reg_15_ ( .D(N1181), .CK(clk), .RN(rstn), .Q(x7_tmp2[15])
         );
  DFFRHQX1 x7_tmp2_reg_14_ ( .D(N1180), .CK(clk), .RN(rstn), .Q(x7_tmp2[14])
         );
  DFFRHQX1 x7_tmp2_reg_13_ ( .D(N1179), .CK(clk), .RN(rstn), .Q(x7_tmp2[13])
         );
  DFFRHQX1 x7_tmp2_reg_12_ ( .D(N1178), .CK(clk), .RN(rstn), .Q(x7_tmp2[12])
         );
  DFFRHQX1 x7_tmp_reg_14_ ( .D(N1204), .CK(clk), .RN(rstn), .Q(x7_tmp[14]) );
  DFFRHQX1 x7_tmp_reg_15_ ( .D(N1205), .CK(clk), .RN(rstn), .Q(x7_tmp[15]) );
  DFFRHQX1 x7_tmp_reg_16_ ( .D(N1206), .CK(clk), .RN(rstn), .Q(x7_tmp[16]) );
  DFFRHQX1 x7_tmp_reg_17_ ( .D(N1207), .CK(clk), .RN(rstn), .Q(x7_tmp[17]) );
  DFFRHQX1 x5_tmp_reg_17_ ( .D(N991), .CK(clk), .RN(rstn), .Q(x5_tmp[17]) );
  DFFRHQX1 x5_tmp_reg_16_ ( .D(N990), .CK(clk), .RN(rstn), .Q(x5_tmp[16]) );
  DFFRHQX1 x5_tmp_reg_15_ ( .D(N989), .CK(clk), .RN(rstn), .Q(x5_tmp[15]) );
  DFFRHQX1 x5_tmp_reg_14_ ( .D(N988), .CK(clk), .RN(rstn), .Q(x5_tmp[14]) );
  DFFRHQX1 x6_tmp_reg_17_ ( .D(N1134), .CK(clk), .RN(rstn), .Q(x6_tmp[17]) );
  DFFRHQX1 x6_tmp_reg_16_ ( .D(N1133), .CK(clk), .RN(rstn), .Q(x6_tmp[16]) );
  DFFRHQX1 x6_tmp_reg_15_ ( .D(N1132), .CK(clk), .RN(rstn), .Q(x6_tmp[15]) );
  DFFRHQX1 x6_tmp_reg_14_ ( .D(N1131), .CK(clk), .RN(rstn), .Q(x6_tmp[14]) );
  DFFRHQX1 x4_tmp_reg_14_ ( .D(N868), .CK(clk), .RN(rstn), .Q(x4_tmp[14]) );
  DFFRHQX1 x4_tmp_reg_15_ ( .D(N869), .CK(clk), .RN(rstn), .Q(x4_tmp[15]) );
  DFFRHQX1 x4_tmp_reg_16_ ( .D(N870), .CK(clk), .RN(rstn), .Q(x4_tmp[16]) );
  DFFRHQX1 x4_tmp_reg_17_ ( .D(N871), .CK(clk), .RN(rstn), .Q(x4_tmp[17]) );
  DFFRHQX1 y6_tmp_reg_14_ ( .D(N1538), .CK(clk), .RN(rstn), .Q(y6_tmp[14]) );
  DFFRHQX1 y6_tmp_reg_13_ ( .D(N1537), .CK(clk), .RN(rstn), .Q(y6_tmp[13]) );
  DFFRHQX1 y6_tmp_reg_12_ ( .D(N1536), .CK(clk), .RN(rstn), .Q(y6_tmp[12]) );
  DFFRHQX1 y6_tmp_reg_11_ ( .D(N1535), .CK(clk), .RN(rstn), .Q(y6_tmp[11]) );
  DFFRHQX1 y6_tmp_reg_10_ ( .D(N1534), .CK(clk), .RN(rstn), .Q(y6_tmp[10]) );
  DFFRHQX1 y7_tmp_reg_14_ ( .D(N1615), .CK(clk), .RN(rstn), .Q(y7_tmp[14]) );
  DFFRHQX1 y7_tmp_reg_13_ ( .D(N1614), .CK(clk), .RN(rstn), .Q(y7_tmp[13]) );
  DFFRHQX1 y7_tmp_reg_12_ ( .D(N1613), .CK(clk), .RN(rstn), .Q(y7_tmp[12]) );
  DFFRHQX1 y7_tmp_reg_11_ ( .D(N1612), .CK(clk), .RN(rstn), .Q(y7_tmp[11]) );
  DFFRHQX1 y7_tmp_reg_10_ ( .D(N1611), .CK(clk), .RN(rstn), .Q(y7_tmp[10]) );
  DFFRHQX1 y0_tmp_reg_16_ ( .D(N1231), .CK(clk), .RN(rstn), .Q(y0_tmp[16]) );
  DFFRHQX1 y0_tmp_reg_15_ ( .D(N1230), .CK(clk), .RN(rstn), .Q(y0_tmp[15]) );
  DFFRHQX1 y0_tmp_reg_14_ ( .D(N1229), .CK(clk), .RN(rstn), .Q(y0_tmp[14]) );
  DFFRHQX1 y0_tmp_reg_13_ ( .D(N1228), .CK(clk), .RN(rstn), .Q(y0_tmp[13]) );
  DFFRHQX1 y0_tmp_reg_12_ ( .D(N1227), .CK(clk), .RN(rstn), .Q(y0_tmp[12]) );
  DFFRHQX1 y1_tmp_reg_16_ ( .D(N1257), .CK(clk), .RN(rstn), .Q(y1_tmp[16]) );
  DFFRHQX1 y1_tmp_reg_15_ ( .D(N1256), .CK(clk), .RN(rstn), .Q(y1_tmp[15]) );
  DFFRHQX1 y1_tmp_reg_14_ ( .D(N1255), .CK(clk), .RN(rstn), .Q(y1_tmp[14]) );
  DFFRHQX1 y1_tmp_reg_13_ ( .D(N1254), .CK(clk), .RN(rstn), .Q(y1_tmp[13]) );
  DFFRHQX1 y1_tmp_reg_12_ ( .D(N1253), .CK(clk), .RN(rstn), .Q(y1_tmp[12]) );
  DFFRHQX1 y2_tmp_reg_16_ ( .D(N1283), .CK(clk), .RN(rstn), .Q(y2_tmp[16]) );
  DFFRHQX1 y2_tmp_reg_15_ ( .D(N1282), .CK(clk), .RN(rstn), .Q(y2_tmp[15]) );
  DFFRHQX1 y2_tmp_reg_14_ ( .D(N1281), .CK(clk), .RN(rstn), .Q(y2_tmp[14]) );
  DFFRHQX1 y2_tmp_reg_13_ ( .D(N1280), .CK(clk), .RN(rstn), .Q(y2_tmp[13]) );
  DFFRHQX1 y2_tmp_reg_12_ ( .D(N1279), .CK(clk), .RN(rstn), .Q(y2_tmp[12]) );
  DFFRHQX1 y3_tmp_reg_16_ ( .D(N1309), .CK(clk), .RN(rstn), .Q(y3_tmp[16]) );
  DFFRHQX1 y3_tmp_reg_15_ ( .D(N1308), .CK(clk), .RN(rstn), .Q(y3_tmp[15]) );
  DFFRHQX1 y3_tmp_reg_14_ ( .D(N1307), .CK(clk), .RN(rstn), .Q(y3_tmp[14]) );
  DFFRHQX1 y3_tmp_reg_13_ ( .D(N1306), .CK(clk), .RN(rstn), .Q(y3_tmp[13]) );
  DFFRHQX1 y3_tmp_reg_12_ ( .D(N1305), .CK(clk), .RN(rstn), .Q(y3_tmp[12]) );
  DFFRHQX1 y4_tmp_reg_14_ ( .D(N1384), .CK(clk), .RN(rstn), .Q(y4_tmp[14]) );
  DFFRHQX1 y4_tmp_reg_13_ ( .D(N1383), .CK(clk), .RN(rstn), .Q(y4_tmp[13]) );
  DFFRHQX1 y4_tmp_reg_12_ ( .D(N1382), .CK(clk), .RN(rstn), .Q(y4_tmp[12]) );
  DFFRHQX1 y4_tmp_reg_11_ ( .D(N1381), .CK(clk), .RN(rstn), .Q(y4_tmp[11]) );
  DFFRHQX1 y4_tmp_reg_10_ ( .D(N1380), .CK(clk), .RN(rstn), .Q(y4_tmp[10]) );
  DFFRHQX1 y5_tmp_reg_14_ ( .D(N1461), .CK(clk), .RN(rstn), .Q(y5_tmp[14]) );
  DFFRHQX1 y5_tmp_reg_13_ ( .D(N1460), .CK(clk), .RN(rstn), .Q(y5_tmp[13]) );
  DFFRHQX1 y5_tmp_reg_12_ ( .D(N1459), .CK(clk), .RN(rstn), .Q(y5_tmp[12]) );
  DFFRHQX1 y5_tmp_reg_11_ ( .D(N1458), .CK(clk), .RN(rstn), .Q(y5_tmp[11]) );
  DFFRHQX1 y5_tmp_reg_10_ ( .D(N1457), .CK(clk), .RN(rstn), .Q(y5_tmp[10]) );
  DFFRHQX1 x7_89_tmp1_reg_9_ ( .D(N281), .CK(clk), .RN(rstn), .Q(x7_89_tmp1[9]) );
  DFFRHQX1 x7_89_tmp1_reg_8_ ( .D(N280), .CK(clk), .RN(rstn), .Q(x7_89_tmp1[8]) );
  DFFRHQX1 x7_89_tmp1_reg_7_ ( .D(N279), .CK(clk), .RN(rstn), .Q(x7_89_tmp1[7]) );
  DFFRHQX1 x7_89_tmp1_reg_6_ ( .D(N278), .CK(clk), .RN(rstn), .Q(x7_89_tmp1[6]) );
  DFFRHQX1 x6_89_tmp1_reg_9_ ( .D(N196), .CK(clk), .RN(rstn), .Q(x6_89_tmp1[9]) );
  DFFRHQX1 x6_89_tmp1_reg_8_ ( .D(N195), .CK(clk), .RN(rstn), .Q(x6_89_tmp1[8]) );
  DFFRHQX1 x6_89_tmp1_reg_7_ ( .D(N194), .CK(clk), .RN(rstn), .Q(x6_89_tmp1[7]) );
  DFFRHQX1 x6_89_tmp1_reg_6_ ( .D(N193), .CK(clk), .RN(rstn), .Q(x6_89_tmp1[6]) );
  DFFRHQX1 x5_89_tmp1_reg_9_ ( .D(N111), .CK(clk), .RN(rstn), .Q(x5_89_tmp1[9]) );
  DFFRHQX1 x5_89_tmp1_reg_8_ ( .D(N110), .CK(clk), .RN(rstn), .Q(x5_89_tmp1[8]) );
  DFFRHQX1 x5_89_tmp1_reg_7_ ( .D(N109), .CK(clk), .RN(rstn), .Q(x5_89_tmp1[7]) );
  DFFRHQX1 x5_89_tmp1_reg_6_ ( .D(N108), .CK(clk), .RN(rstn), .Q(x5_89_tmp1[6]) );
  DFFRHQX1 x5_75_tmp1_reg_9_ ( .D(N111), .CK(clk), .RN(rstn), .Q(x5_75_tmp1[9]) );
  DFFRHQX1 x5_75_tmp1_reg_8_ ( .D(N110), .CK(clk), .RN(rstn), .Q(x5_75_tmp1[8]) );
  DFFRHQX1 x5_75_tmp1_reg_7_ ( .D(N109), .CK(clk), .RN(rstn), .Q(x5_75_tmp1[7]) );
  DFFRHQX1 x5_75_tmp1_reg_6_ ( .D(N108), .CK(clk), .RN(rstn), .Q(x5_75_tmp1[6]) );
  DFFRHQX1 x4_75_tmp1_reg_9_ ( .D(N26), .CK(clk), .RN(rstn), .Q(x4_75_tmp1[9])
         );
  DFFRHQX1 x4_75_tmp1_reg_8_ ( .D(N25), .CK(clk), .RN(rstn), .Q(x4_75_tmp1[8])
         );
  DFFRHQX1 x4_75_tmp1_reg_7_ ( .D(N24), .CK(clk), .RN(rstn), .Q(x4_75_tmp1[7])
         );
  DFFRHQX1 x4_75_tmp1_reg_6_ ( .D(N23), .CK(clk), .RN(rstn), .Q(x4_75_tmp1[6])
         );
  DFFRHQX1 x7_75_tmp1_reg_9_ ( .D(N281), .CK(clk), .RN(rstn), .Q(x7_75_tmp1[9]) );
  DFFRHQX1 x7_75_tmp1_reg_8_ ( .D(N280), .CK(clk), .RN(rstn), .Q(x7_75_tmp1[8]) );
  DFFRHQX1 x7_75_tmp1_reg_7_ ( .D(N279), .CK(clk), .RN(rstn), .Q(x7_75_tmp1[7]) );
  DFFRHQX1 x7_75_tmp1_reg_6_ ( .D(N278), .CK(clk), .RN(rstn), .Q(x7_75_tmp1[6]) );
  DFFRHQX1 x6_75_tmp1_reg_9_ ( .D(N196), .CK(clk), .RN(rstn), .Q(x6_75_tmp1[9]) );
  DFFRHQX1 x6_75_tmp1_reg_8_ ( .D(N195), .CK(clk), .RN(rstn), .Q(x6_75_tmp1[8]) );
  DFFRHQX1 x6_75_tmp1_reg_7_ ( .D(N194), .CK(clk), .RN(rstn), .Q(x6_75_tmp1[7]) );
  DFFRHQX1 x6_75_tmp1_reg_6_ ( .D(N193), .CK(clk), .RN(rstn), .Q(x6_75_tmp1[6]) );
  DFFRHQX1 x4_50_tmp1_reg_8_ ( .D(n77), .CK(clk), .RN(rstn), .Q(x4_50_tmp1[8])
         );
  DFFRHQX1 x4_50_tmp1_reg_7_ ( .D(n76), .CK(clk), .RN(rstn), .Q(x4_50_tmp1[7])
         );
  DFFRHQX1 x4_50_tmp1_reg_6_ ( .D(x4[1]), .CK(clk), .RN(rstn), .Q(
        x4_50_tmp1[6]) );
  DFFRHQX1 x6_50_tmp1_reg_8_ ( .D(n51), .CK(clk), .RN(rstn), .Q(x6_50_tmp1[8])
         );
  DFFRHQX1 x6_50_tmp1_reg_7_ ( .D(n50), .CK(clk), .RN(rstn), .Q(x6_50_tmp1[7])
         );
  DFFRHQX1 x6_50_tmp1_reg_6_ ( .D(x6[1]), .CK(clk), .RN(rstn), .Q(
        x6_50_tmp1[6]) );
  DFFRHQX1 x5_50_tmp1_reg_8_ ( .D(n64), .CK(clk), .RN(rstn), .Q(x5_50_tmp1[8])
         );
  DFFRHQX1 x5_50_tmp1_reg_7_ ( .D(n63), .CK(clk), .RN(rstn), .Q(x5_50_tmp1[7])
         );
  DFFRHQX1 x5_50_tmp1_reg_6_ ( .D(x5[1]), .CK(clk), .RN(rstn), .Q(
        x5_50_tmp1[6]) );
  DFFRHQX1 x7_50_tmp1_reg_8_ ( .D(n38), .CK(clk), .RN(rstn), .Q(x7_50_tmp1[8])
         );
  DFFRHQX1 x7_50_tmp1_reg_7_ ( .D(n37), .CK(clk), .RN(rstn), .Q(x7_50_tmp1[7])
         );
  DFFRHQX1 x7_50_tmp1_reg_6_ ( .D(x7[1]), .CK(clk), .RN(rstn), .Q(
        x7_50_tmp1[6]) );
  DFFRHQX1 x4_18_tmp1_reg_7_ ( .D(n77), .CK(clk), .RN(rstn), .Q(x4_18_tmp1[7])
         );
  DFFRHQX1 x4_18_tmp1_reg_6_ ( .D(n76), .CK(clk), .RN(rstn), .Q(x4_18_tmp1[6])
         );
  DFFRHQX1 x4_18_tmp1_reg_5_ ( .D(x4[1]), .CK(clk), .RN(rstn), .Q(
        x4_18_tmp1[5]) );
  DFFRHQX1 x5_18_tmp1_reg_7_ ( .D(n64), .CK(clk), .RN(rstn), .Q(x5_18_tmp1[7])
         );
  DFFRHQX1 x5_18_tmp1_reg_6_ ( .D(n63), .CK(clk), .RN(rstn), .Q(x5_18_tmp1[6])
         );
  DFFRHQX1 x5_18_tmp1_reg_5_ ( .D(x5[1]), .CK(clk), .RN(rstn), .Q(
        x5_18_tmp1[5]) );
  DFFRHQX1 x6_18_tmp1_reg_7_ ( .D(n51), .CK(clk), .RN(rstn), .Q(x6_18_tmp1[7])
         );
  DFFRHQX1 x6_18_tmp1_reg_6_ ( .D(n50), .CK(clk), .RN(rstn), .Q(x6_18_tmp1[6])
         );
  DFFRHQX1 x6_18_tmp1_reg_5_ ( .D(x6[1]), .CK(clk), .RN(rstn), .Q(
        x6_18_tmp1[5]) );
  DFFRHQX1 x7_18_tmp1_reg_7_ ( .D(n38), .CK(clk), .RN(rstn), .Q(x7_18_tmp1[7])
         );
  DFFRHQX1 x7_18_tmp1_reg_6_ ( .D(n37), .CK(clk), .RN(rstn), .Q(x7_18_tmp1[6])
         );
  DFFRHQX1 x7_18_tmp1_reg_5_ ( .D(x7[1]), .CK(clk), .RN(rstn), .Q(
        x7_18_tmp1[5]) );
  DFFRHQX1 x5_18_reg_12_ ( .D(N526), .CK(clk), .RN(rstn), .Q(x5_18[12]) );
  DFFRHQX1 x5_18_reg_11_ ( .D(N525), .CK(clk), .RN(rstn), .Q(x5_18[11]) );
  DFFRHQX1 x5_18_reg_10_ ( .D(N524), .CK(clk), .RN(rstn), .Q(x5_18[10]) );
  DFFRHQX1 x5_18_reg_9_ ( .D(N523), .CK(clk), .RN(rstn), .Q(x5_18[9]) );
  DFFRHQX1 x5_18_reg_8_ ( .D(N522), .CK(clk), .RN(rstn), .Q(x5_18[8]) );
  DFFRHQX1 x6_18_reg_10_ ( .D(N613), .CK(clk), .RN(rstn), .Q(x6_18[10]) );
  DFFRHQX1 x6_18_reg_9_ ( .D(N612), .CK(clk), .RN(rstn), .Q(x6_18[9]) );
  DFFRHQX1 x6_18_reg_8_ ( .D(N611), .CK(clk), .RN(rstn), .Q(x6_18[8]) );
  DFFRHQX1 x6_18_reg_7_ ( .D(N610), .CK(clk), .RN(rstn), .Q(x6_18[7]) );
  DFFRHQX1 x4_18_reg_10_ ( .D(N435), .CK(clk), .RN(rstn), .Q(x4_18[10]) );
  DFFRHQX1 x4_18_reg_9_ ( .D(N434), .CK(clk), .RN(rstn), .Q(x4_18[9]) );
  DFFRHQX1 x4_18_reg_8_ ( .D(N433), .CK(clk), .RN(rstn), .Q(x4_18[8]) );
  DFFRHQX1 x4_18_reg_7_ ( .D(N432), .CK(clk), .RN(rstn), .Q(x4_18[7]) );
  DFFRHQX1 x4_89_tmp1_reg_9_ ( .D(N26), .CK(clk), .RN(rstn), .Q(x4_89_tmp1[9])
         );
  DFFRHQX1 x4_89_tmp1_reg_8_ ( .D(N25), .CK(clk), .RN(rstn), .Q(x4_89_tmp1[8])
         );
  DFFRHQX1 x4_89_tmp1_reg_7_ ( .D(N24), .CK(clk), .RN(rstn), .Q(x4_89_tmp1[7])
         );
  DFFRHQX1 x4_89_tmp1_reg_6_ ( .D(N23), .CK(clk), .RN(rstn), .Q(x4_89_tmp1[6])
         );
  DFFRHQX1 x4_89_reg_10_ ( .D(N367), .CK(clk), .RN(rstn), .Q(x4_89[10]) );
  DFFRHQX1 x4_89_reg_9_ ( .D(N366), .CK(clk), .RN(rstn), .Q(x4_89[9]) );
  DFFRHQX1 x4_89_reg_8_ ( .D(N365), .CK(clk), .RN(rstn), .Q(x4_89[8]) );
  DFFRHQX1 x4_89_reg_7_ ( .D(N364), .CK(clk), .RN(rstn), .Q(x4_89[7]) );
  DFFRHQX1 x4_75_reg_10_ ( .D(N390), .CK(clk), .RN(rstn), .Q(x4_75[10]) );
  DFFRHQX1 x4_75_reg_9_ ( .D(N389), .CK(clk), .RN(rstn), .Q(x4_75[9]) );
  DFFRHQX1 x4_75_reg_8_ ( .D(N388), .CK(clk), .RN(rstn), .Q(x4_75[8]) );
  DFFRHQX1 x4_75_reg_7_ ( .D(N387), .CK(clk), .RN(rstn), .Q(x4_75[7]) );
  DFFRHQX1 x5_75_reg_10_ ( .D(N479), .CK(clk), .RN(rstn), .Q(x5_75[10]) );
  DFFRHQX1 x5_75_reg_9_ ( .D(N478), .CK(clk), .RN(rstn), .Q(x5_75[9]) );
  DFFRHQX1 x5_75_reg_8_ ( .D(N477), .CK(clk), .RN(rstn), .Q(x5_75[8]) );
  DFFRHQX1 x5_75_reg_7_ ( .D(N476), .CK(clk), .RN(rstn), .Q(x5_75[7]) );
  DFFRHQX1 x6_75_reg_10_ ( .D(N568), .CK(clk), .RN(rstn), .Q(x6_75[10]) );
  DFFRHQX1 x6_75_reg_9_ ( .D(N567), .CK(clk), .RN(rstn), .Q(x6_75[9]) );
  DFFRHQX1 x6_75_reg_8_ ( .D(N566), .CK(clk), .RN(rstn), .Q(x6_75[8]) );
  DFFRHQX1 x6_75_reg_7_ ( .D(N565), .CK(clk), .RN(rstn), .Q(x6_75[7]) );
  DFFRHQX1 x4_50_reg_10_ ( .D(N413), .CK(clk), .RN(rstn), .Q(x4_50[10]) );
  DFFRHQX1 x4_50_reg_9_ ( .D(N412), .CK(clk), .RN(rstn), .Q(x4_50[9]) );
  DFFRHQX1 x4_50_reg_8_ ( .D(N411), .CK(clk), .RN(rstn), .Q(x4_50[8]) );
  DFFRHQX1 x4_50_reg_7_ ( .D(N410), .CK(clk), .RN(rstn), .Q(x4_50[7]) );
  DFFRHQX1 x5_tmp1_reg_11_ ( .D(N890), .CK(clk), .RN(rstn), .Q(x5_tmp1[11]) );
  DFFRHQX1 x5_tmp1_reg_10_ ( .D(N889), .CK(clk), .RN(rstn), .Q(x5_tmp1[10]) );
  DFFRHQX1 x5_tmp1_reg_9_ ( .D(N888), .CK(clk), .RN(rstn), .Q(x5_tmp1[9]) );
  DFFRHQX1 x5_tmp1_reg_8_ ( .D(N887), .CK(clk), .RN(rstn), .Q(x5_tmp1[8]) );
  DFFRHQX1 x6_tmp1_reg_11_ ( .D(N1056), .CK(clk), .RN(rstn), .Q(x6_tmp1[11])
         );
  DFFRHQX1 x6_tmp1_reg_10_ ( .D(N1055), .CK(clk), .RN(rstn), .Q(x6_tmp1[10])
         );
  DFFRHQX1 x6_tmp1_reg_9_ ( .D(N1054), .CK(clk), .RN(rstn), .Q(x6_tmp1[9]) );
  DFFRHQX1 x6_tmp1_reg_8_ ( .D(N1053), .CK(clk), .RN(rstn), .Q(x6_tmp1[8]) );
  DFFRHQX1 x7_tmp1_reg_11_ ( .D(N1153), .CK(clk), .RN(rstn), .Q(x7_tmp1[11])
         );
  DFFRHQX1 x7_tmp1_reg_10_ ( .D(N1152), .CK(clk), .RN(rstn), .Q(x7_tmp1[10])
         );
  DFFRHQX1 x7_tmp1_reg_9_ ( .D(N1151), .CK(clk), .RN(rstn), .Q(x7_tmp1[9]) );
  DFFRHQX1 x7_tmp1_reg_8_ ( .D(N1150), .CK(clk), .RN(rstn), .Q(x7_tmp1[8]) );
  DFFRHQX1 x4_tmp1_reg_11_ ( .D(N771), .CK(clk), .RN(rstn), .Q(x4_tmp1[11]) );
  DFFRHQX1 x4_tmp1_reg_10_ ( .D(N770), .CK(clk), .RN(rstn), .Q(x4_tmp1[10]) );
  DFFRHQX1 x4_tmp1_reg_9_ ( .D(N769), .CK(clk), .RN(rstn), .Q(x4_tmp1[9]) );
  DFFRHQX1 x4_tmp1_reg_8_ ( .D(N768), .CK(clk), .RN(rstn), .Q(x4_tmp1[8]) );
  DFFRHQX1 idct8_ready_reg ( .D(start), .CK(clk), .RN(rstn), .Q(idct8_ready)
         );
  DFFRHQX1 x7_50_reg_11_ ( .D(N681), .CK(clk), .RN(rstn), .Q(x7_50[11]) );
  DFFRHQX1 x7_50_reg_10_ ( .D(N680), .CK(clk), .RN(rstn), .Q(x7_50[10]) );
  DFFRHQX1 x7_50_reg_9_ ( .D(N679), .CK(clk), .RN(rstn), .Q(x7_50[9]) );
  DFFRHQX1 x7_50_reg_8_ ( .D(N678), .CK(clk), .RN(rstn), .Q(x7_50[8]) );
  DFFRHQX1 x7_50_reg_7_ ( .D(N677), .CK(clk), .RN(rstn), .Q(x7_50[7]) );
  DFFRHQX1 x5_89_reg_11_ ( .D(N457), .CK(clk), .RN(rstn), .Q(x5_89[11]) );
  DFFRHQX1 x5_89_reg_10_ ( .D(N456), .CK(clk), .RN(rstn), .Q(x5_89[10]) );
  DFFRHQX1 x5_89_reg_9_ ( .D(N455), .CK(clk), .RN(rstn), .Q(x5_89[9]) );
  DFFRHQX1 x5_89_reg_8_ ( .D(N454), .CK(clk), .RN(rstn), .Q(x5_89[8]) );
  DFFRHQX1 x5_89_reg_7_ ( .D(N453), .CK(clk), .RN(rstn), .Q(x5_89[7]) );
  DFFRHQX1 x7_89_reg_11_ ( .D(N635), .CK(clk), .RN(rstn), .Q(x7_89[11]) );
  DFFRHQX1 x7_89_reg_10_ ( .D(N634), .CK(clk), .RN(rstn), .Q(x7_89[10]) );
  DFFRHQX1 x7_89_reg_9_ ( .D(N633), .CK(clk), .RN(rstn), .Q(x7_89[9]) );
  DFFRHQX1 x7_89_reg_8_ ( .D(N632), .CK(clk), .RN(rstn), .Q(x7_89[8]) );
  DFFRHQX1 x7_89_reg_7_ ( .D(N631), .CK(clk), .RN(rstn), .Q(x7_89[7]) );
  DFFRHQX1 x5_50_reg_11_ ( .D(N503), .CK(clk), .RN(rstn), .Q(x5_50[11]) );
  DFFRHQX1 x5_50_reg_10_ ( .D(N502), .CK(clk), .RN(rstn), .Q(x5_50[10]) );
  DFFRHQX1 x5_50_reg_9_ ( .D(N501), .CK(clk), .RN(rstn), .Q(x5_50[9]) );
  DFFRHQX1 x5_50_reg_8_ ( .D(N500), .CK(clk), .RN(rstn), .Q(x5_50[8]) );
  DFFRHQX1 x5_50_reg_7_ ( .D(N499), .CK(clk), .RN(rstn), .Q(x5_50[7]) );
  DFFRHQX1 x6_89_tmp2_reg_9_ ( .D(N219), .CK(clk), .RN(rstn), .Q(x6_89_tmp2[9]) );
  DFFRHQX1 x6_89_tmp2_reg_8_ ( .D(N218), .CK(clk), .RN(rstn), .Q(x6_89_tmp2[8]) );
  DFFRHQX1 x6_89_tmp2_reg_7_ ( .D(N217), .CK(clk), .RN(rstn), .Q(x6_89_tmp2[7]) );
  DFFRHQX1 x6_89_tmp2_reg_6_ ( .D(N216), .CK(clk), .RN(rstn), .Q(x6_89_tmp2[6]) );
  DFFRHQX1 x5_89_tmp2_reg_9_ ( .D(N134), .CK(clk), .RN(rstn), .Q(x5_89_tmp2[9]) );
  DFFRHQX1 x5_89_tmp2_reg_8_ ( .D(N133), .CK(clk), .RN(rstn), .Q(x5_89_tmp2[8]) );
  DFFRHQX1 x5_89_tmp2_reg_7_ ( .D(N132), .CK(clk), .RN(rstn), .Q(x5_89_tmp2[7]) );
  DFFRHQX1 x5_89_tmp2_reg_6_ ( .D(N131), .CK(clk), .RN(rstn), .Q(x5_89_tmp2[6]) );
  DFFRHQX1 x4_89_tmp2_reg_9_ ( .D(N49), .CK(clk), .RN(rstn), .Q(x4_89_tmp2[9])
         );
  DFFRHQX1 x4_89_tmp2_reg_8_ ( .D(N48), .CK(clk), .RN(rstn), .Q(x4_89_tmp2[8])
         );
  DFFRHQX1 x4_89_tmp2_reg_7_ ( .D(N47), .CK(clk), .RN(rstn), .Q(x4_89_tmp2[7])
         );
  DFFRHQX1 x4_89_tmp2_reg_6_ ( .D(N46), .CK(clk), .RN(rstn), .Q(x4_89_tmp2[6])
         );
  DFFRHQX1 x7_89_tmp2_reg_9_ ( .D(N304), .CK(clk), .RN(rstn), .Q(x7_89_tmp2[9]) );
  DFFRHQX1 x7_89_tmp2_reg_8_ ( .D(N303), .CK(clk), .RN(rstn), .Q(x7_89_tmp2[8]) );
  DFFRHQX1 x7_89_tmp2_reg_7_ ( .D(N302), .CK(clk), .RN(rstn), .Q(x7_89_tmp2[7]) );
  DFFRHQX1 x7_89_tmp2_reg_6_ ( .D(N301), .CK(clk), .RN(rstn), .Q(x7_89_tmp2[6]) );
  DFFRHQX1 x4_75_tmp2_reg_9_ ( .D(N70), .CK(clk), .RN(rstn), .Q(x4_75_tmp2[9])
         );
  DFFRHQX1 x4_75_tmp2_reg_8_ ( .D(N69), .CK(clk), .RN(rstn), .Q(x4_75_tmp2[8])
         );
  DFFRHQX1 x4_75_tmp2_reg_7_ ( .D(N68), .CK(clk), .RN(rstn), .Q(x4_75_tmp2[7])
         );
  DFFRHQX1 x4_75_tmp2_reg_6_ ( .D(N67), .CK(clk), .RN(rstn), .Q(x4_75_tmp2[6])
         );
  DFFRHQX1 x5_75_tmp2_reg_9_ ( .D(N155), .CK(clk), .RN(rstn), .Q(x5_75_tmp2[9]) );
  DFFRHQX1 x5_75_tmp2_reg_8_ ( .D(N154), .CK(clk), .RN(rstn), .Q(x5_75_tmp2[8]) );
  DFFRHQX1 x5_75_tmp2_reg_7_ ( .D(N153), .CK(clk), .RN(rstn), .Q(x5_75_tmp2[7]) );
  DFFRHQX1 x5_75_tmp2_reg_6_ ( .D(N152), .CK(clk), .RN(rstn), .Q(x5_75_tmp2[6]) );
  DFFRHQX1 x6_75_tmp2_reg_9_ ( .D(N240), .CK(clk), .RN(rstn), .Q(x6_75_tmp2[9]) );
  DFFRHQX1 x6_75_tmp2_reg_8_ ( .D(N239), .CK(clk), .RN(rstn), .Q(x6_75_tmp2[8]) );
  DFFRHQX1 x6_75_tmp2_reg_7_ ( .D(N238), .CK(clk), .RN(rstn), .Q(x6_75_tmp2[7]) );
  DFFRHQX1 x6_75_tmp2_reg_6_ ( .D(N237), .CK(clk), .RN(rstn), .Q(x6_75_tmp2[6]) );
  DFFRHQX1 x7_75_tmp2_reg_9_ ( .D(N325), .CK(clk), .RN(rstn), .Q(x7_75_tmp2[9]) );
  DFFRHQX1 x7_75_tmp2_reg_8_ ( .D(N324), .CK(clk), .RN(rstn), .Q(x7_75_tmp2[8]) );
  DFFRHQX1 x7_75_tmp2_reg_7_ ( .D(N323), .CK(clk), .RN(rstn), .Q(x7_75_tmp2[7]) );
  DFFRHQX1 x7_75_tmp2_reg_6_ ( .D(N322), .CK(clk), .RN(rstn), .Q(x7_75_tmp2[6]) );
  DFFRHQX1 x4_50_tmp2_reg_8_ ( .D(N89), .CK(clk), .RN(rstn), .Q(x4_50_tmp2[8])
         );
  DFFRHQX1 x4_50_tmp2_reg_7_ ( .D(N88), .CK(clk), .RN(rstn), .Q(x4_50_tmp2[7])
         );
  DFFRHQX1 x4_50_tmp2_reg_6_ ( .D(N87), .CK(clk), .RN(rstn), .Q(x4_50_tmp2[6])
         );
  DFFRHQX1 x6_50_tmp2_reg_8_ ( .D(N259), .CK(clk), .RN(rstn), .Q(x6_50_tmp2[8]) );
  DFFRHQX1 x6_50_tmp2_reg_7_ ( .D(N258), .CK(clk), .RN(rstn), .Q(x6_50_tmp2[7]) );
  DFFRHQX1 x6_50_tmp2_reg_6_ ( .D(N257), .CK(clk), .RN(rstn), .Q(x6_50_tmp2[6]) );
  DFFRHQX1 x6_50_reg_7_ ( .D(N588), .CK(clk), .RN(rstn), .Q(x6_50[7]) );
  DFFRHQX1 x6_50_reg_8_ ( .D(N589), .CK(clk), .RN(rstn), .Q(x6_50[8]) );
  DFFRHQX1 x6_50_reg_9_ ( .D(N590), .CK(clk), .RN(rstn), .Q(x6_50[9]) );
  DFFRHQX1 x6_50_reg_10_ ( .D(N591), .CK(clk), .RN(rstn), .Q(x6_50[10]) );
  DFFRHQX1 x5_50_tmp2_reg_8_ ( .D(N174), .CK(clk), .RN(rstn), .Q(x5_50_tmp2[8]) );
  DFFRHQX1 x5_50_tmp2_reg_7_ ( .D(N173), .CK(clk), .RN(rstn), .Q(x5_50_tmp2[7]) );
  DFFRHQX1 x5_50_tmp2_reg_6_ ( .D(N172), .CK(clk), .RN(rstn), .Q(x5_50_tmp2[6]) );
  DFFRHQX1 x7_50_tmp2_reg_8_ ( .D(N344), .CK(clk), .RN(rstn), .Q(x7_50_tmp2[8]) );
  DFFRHQX1 x7_50_tmp2_reg_7_ ( .D(N343), .CK(clk), .RN(rstn), .Q(x7_50_tmp2[7]) );
  DFFRHQX1 x7_50_tmp2_reg_6_ ( .D(N342), .CK(clk), .RN(rstn), .Q(x7_50_tmp2[6]) );
  DFFRHQX1 x4_18_tmp2_reg_7_ ( .D(n80), .CK(clk), .RN(rstn), .Q(x4_18_tmp2[7])
         );
  DFFRHQX1 x4_18_tmp2_reg_6_ ( .D(n79), .CK(clk), .RN(rstn), .Q(x4_18_tmp2[6])
         );
  DFFRHQX1 x4_18_tmp2_reg_5_ ( .D(n78), .CK(clk), .RN(rstn), .Q(x4_18_tmp2[5])
         );
  DFFRHQX1 x6_18_tmp2_reg_7_ ( .D(n54), .CK(clk), .RN(rstn), .Q(x6_18_tmp2[7])
         );
  DFFRHQX1 x6_18_tmp2_reg_6_ ( .D(n53), .CK(clk), .RN(rstn), .Q(x6_18_tmp2[6])
         );
  DFFRHQX1 x6_18_tmp2_reg_5_ ( .D(n52), .CK(clk), .RN(rstn), .Q(x6_18_tmp2[5])
         );
  DFFRHQX1 x5_18_tmp2_reg_7_ ( .D(n67), .CK(clk), .RN(rstn), .Q(x5_18_tmp2[7])
         );
  DFFRHQX1 x5_18_tmp2_reg_6_ ( .D(n66), .CK(clk), .RN(rstn), .Q(x5_18_tmp2[6])
         );
  DFFRHQX1 x5_18_tmp2_reg_5_ ( .D(n65), .CK(clk), .RN(rstn), .Q(x5_18_tmp2[5])
         );
  DFFRHQX1 x7_18_tmp2_reg_7_ ( .D(n41), .CK(clk), .RN(rstn), .Q(x7_18_tmp2[7])
         );
  DFFRHQX1 x7_18_tmp2_reg_6_ ( .D(n40), .CK(clk), .RN(rstn), .Q(x7_18_tmp2[6])
         );
  DFFRHQX1 x7_18_tmp2_reg_5_ ( .D(n39), .CK(clk), .RN(rstn), .Q(x7_18_tmp2[5])
         );
  DFFRHQX1 x7_18_reg_10_ ( .D(N702), .CK(clk), .RN(rstn), .Q(x7_18[10]) );
  DFFRHQX1 x7_18_reg_9_ ( .D(N701), .CK(clk), .RN(rstn), .Q(x7_18[9]) );
  DFFRHQX1 x7_18_reg_8_ ( .D(N700), .CK(clk), .RN(rstn), .Q(x7_18[8]) );
  DFFRHQX1 x7_18_reg_7_ ( .D(N699), .CK(clk), .RN(rstn), .Q(x7_18[7]) );
  DFFRHQX1 x6_89_reg_11_ ( .D(N546), .CK(clk), .RN(rstn), .Q(x6_89[11]) );
  DFFRHQX1 x6_89_reg_10_ ( .D(N545), .CK(clk), .RN(rstn), .Q(x6_89[10]) );
  DFFRHQX1 x6_89_reg_9_ ( .D(N544), .CK(clk), .RN(rstn), .Q(x6_89[9]) );
  DFFRHQX1 x6_89_reg_8_ ( .D(N543), .CK(clk), .RN(rstn), .Q(x6_89[8]) );
  DFFRHQX1 x7_75_reg_10_ ( .D(N657), .CK(clk), .RN(rstn), .Q(x7_75[10]) );
  DFFRHQX1 x7_75_reg_9_ ( .D(N656), .CK(clk), .RN(rstn), .Q(x7_75[9]) );
  DFFRHQX1 x7_75_reg_8_ ( .D(N655), .CK(clk), .RN(rstn), .Q(x7_75[8]) );
  DFFRHQX1 x7_75_reg_7_ ( .D(N654), .CK(clk), .RN(rstn), .Q(x7_75[7]) );
  DFFRHQX1 x4_tmp2_reg_11_ ( .D(N841), .CK(clk), .RN(rstn), .Q(x4_tmp2[11]) );
  DFFRHQX1 x4_tmp2_reg_10_ ( .D(N840), .CK(clk), .RN(rstn), .Q(x4_tmp2[10]) );
  DFFRHQX1 x4_tmp2_reg_9_ ( .D(N839), .CK(clk), .RN(rstn), .Q(x4_tmp2[9]) );
  DFFRHQX1 x4_tmp2_reg_8_ ( .D(N838), .CK(clk), .RN(rstn), .Q(x4_tmp2[8]) );
  DFFRHQX1 x5_tmp2_reg_11_ ( .D(N961), .CK(clk), .RN(rstn), .Q(x5_tmp2[11]) );
  DFFRHQX1 x5_tmp2_reg_10_ ( .D(N960), .CK(clk), .RN(rstn), .Q(x5_tmp2[10]) );
  DFFRHQX1 x5_tmp2_reg_9_ ( .D(N959), .CK(clk), .RN(rstn), .Q(x5_tmp2[9]) );
  DFFRHQX1 x5_tmp2_reg_8_ ( .D(N958), .CK(clk), .RN(rstn), .Q(x5_tmp2[8]) );
  DFFRHQX1 x6_tmp2_reg_11_ ( .D(N1104), .CK(clk), .RN(rstn), .Q(x6_tmp2[11])
         );
  DFFRHQX1 x6_tmp2_reg_10_ ( .D(N1103), .CK(clk), .RN(rstn), .Q(x6_tmp2[10])
         );
  DFFRHQX1 x6_tmp2_reg_9_ ( .D(N1102), .CK(clk), .RN(rstn), .Q(x6_tmp2[9]) );
  DFFRHQX1 x6_tmp2_reg_8_ ( .D(N1101), .CK(clk), .RN(rstn), .Q(x6_tmp2[8]) );
  DFFRHQX1 x7_tmp2_reg_11_ ( .D(N1177), .CK(clk), .RN(rstn), .Q(x7_tmp2[11])
         );
  DFFRHQX1 x7_tmp2_reg_10_ ( .D(N1176), .CK(clk), .RN(rstn), .Q(x7_tmp2[10])
         );
  DFFRHQX1 x7_tmp2_reg_9_ ( .D(N1175), .CK(clk), .RN(rstn), .Q(x7_tmp2[9]) );
  DFFRHQX1 x7_tmp2_reg_8_ ( .D(N1174), .CK(clk), .RN(rstn), .Q(x7_tmp2[8]) );
  DFFRHQX1 x4_50_tmp2_reg_5_ ( .D(N86), .CK(clk), .RN(rstn), .Q(x4_50_tmp2[5])
         );
  DFFRHQX1 x6_50_tmp2_reg_5_ ( .D(N256), .CK(clk), .RN(rstn), .Q(x6_50_tmp2[5]) );
  DFFRHQX1 x5_50_tmp2_reg_5_ ( .D(N171), .CK(clk), .RN(rstn), .Q(x5_50_tmp2[5]) );
  DFFRHQX1 x7_50_tmp2_reg_5_ ( .D(N341), .CK(clk), .RN(rstn), .Q(x7_50_tmp2[5]) );
  DFFRHQX1 x4_18_tmp2_reg_4_ ( .D(n77), .CK(clk), .RN(rstn), .Q(x4_18_tmp2[4])
         );
  DFFRHQX1 x6_18_tmp2_reg_4_ ( .D(n51), .CK(clk), .RN(rstn), .Q(x6_18_tmp2[4])
         );
  DFFRHQX1 x5_18_tmp2_reg_4_ ( .D(n64), .CK(clk), .RN(rstn), .Q(x5_18_tmp2[4])
         );
  DFFRHQX1 x7_18_tmp2_reg_4_ ( .D(n38), .CK(clk), .RN(rstn), .Q(x7_18_tmp2[4])
         );
  DFFRHQX1 x4_50_tmp1_reg_5_ ( .D(x4[0]), .CK(clk), .RN(rstn), .Q(
        x4_50_tmp1[5]) );
  DFFRHQX1 x6_50_tmp1_reg_5_ ( .D(x6[0]), .CK(clk), .RN(rstn), .Q(
        x6_50_tmp1[5]) );
  DFFRHQX1 x5_50_tmp1_reg_5_ ( .D(x5[0]), .CK(clk), .RN(rstn), .Q(
        x5_50_tmp1[5]) );
  DFFRHQX1 x7_50_tmp1_reg_5_ ( .D(x7[0]), .CK(clk), .RN(rstn), .Q(
        x7_50_tmp1[5]) );
  DFFRHQX1 x4_18_tmp1_reg_4_ ( .D(x4[0]), .CK(clk), .RN(rstn), .Q(
        x4_18_tmp1[4]) );
  DFFRHQX1 x5_18_tmp1_reg_4_ ( .D(x5[0]), .CK(clk), .RN(rstn), .Q(
        x5_18_tmp1[4]) );
  DFFRHQX1 x6_18_tmp1_reg_4_ ( .D(x6[0]), .CK(clk), .RN(rstn), .Q(
        x6_18_tmp1[4]) );
  DFFRHQX1 x7_18_tmp1_reg_4_ ( .D(x7[0]), .CK(clk), .RN(rstn), .Q(
        x7_18_tmp1[4]) );
  DFFRHQX1 x7_tmp_reg_10_ ( .D(N1200), .CK(clk), .RN(rstn), .Q(x7_tmp[10]) );
  DFFRHQX1 x7_tmp_reg_11_ ( .D(N1201), .CK(clk), .RN(rstn), .Q(x7_tmp[11]) );
  DFFRHQX1 x7_tmp_reg_12_ ( .D(N1202), .CK(clk), .RN(rstn), .Q(x7_tmp[12]) );
  DFFRHQX1 x7_tmp_reg_13_ ( .D(N1203), .CK(clk), .RN(rstn), .Q(x7_tmp[13]) );
  DFFRHQX1 x5_tmp_reg_13_ ( .D(N987), .CK(clk), .RN(rstn), .Q(x5_tmp[13]) );
  DFFRHQX1 x5_tmp_reg_12_ ( .D(N986), .CK(clk), .RN(rstn), .Q(x5_tmp[12]) );
  DFFRHQX1 x5_tmp_reg_11_ ( .D(N985), .CK(clk), .RN(rstn), .Q(x5_tmp[11]) );
  DFFRHQX1 x5_tmp_reg_10_ ( .D(N984), .CK(clk), .RN(rstn), .Q(x5_tmp[10]) );
  DFFRHQX1 x6_tmp_reg_13_ ( .D(N1130), .CK(clk), .RN(rstn), .Q(x6_tmp[13]) );
  DFFRHQX1 x6_tmp_reg_12_ ( .D(N1129), .CK(clk), .RN(rstn), .Q(x6_tmp[12]) );
  DFFRHQX1 x6_tmp_reg_11_ ( .D(N1128), .CK(clk), .RN(rstn), .Q(x6_tmp[11]) );
  DFFRHQX1 x6_tmp_reg_10_ ( .D(N1127), .CK(clk), .RN(rstn), .Q(x6_tmp[10]) );
  DFFRHQX1 x4_tmp_reg_10_ ( .D(N864), .CK(clk), .RN(rstn), .Q(x4_tmp[10]) );
  DFFRHQX1 x4_tmp_reg_11_ ( .D(N865), .CK(clk), .RN(rstn), .Q(x4_tmp[11]) );
  DFFRHQX1 x4_tmp_reg_12_ ( .D(N866), .CK(clk), .RN(rstn), .Q(x4_tmp[12]) );
  DFFRHQX1 x4_tmp_reg_13_ ( .D(N867), .CK(clk), .RN(rstn), .Q(x4_tmp[13]) );
  DFFRHQX1 y6_tmp_reg_9_ ( .D(N1533), .CK(clk), .RN(rstn), .Q(y6_tmp[9]) );
  DFFRHQX1 y6_tmp_reg_8_ ( .D(N1532), .CK(clk), .RN(rstn), .Q(y6_tmp[8]) );
  DFFRHQX1 y6_tmp_reg_7_ ( .D(N1531), .CK(clk), .RN(rstn), .Q(y6_tmp[7]) );
  DFFRHQX1 y7_tmp_reg_9_ ( .D(N1610), .CK(clk), .RN(rstn), .Q(y7_tmp[9]) );
  DFFRHQX1 y7_tmp_reg_8_ ( .D(N1609), .CK(clk), .RN(rstn), .Q(y7_tmp[8]) );
  DFFRHQX1 y7_tmp_reg_7_ ( .D(N1608), .CK(clk), .RN(rstn), .Q(y7_tmp[7]) );
  DFFRHQX1 y0_tmp_reg_11_ ( .D(N1226), .CK(clk), .RN(rstn), .Q(y0_tmp[11]) );
  DFFRHQX1 y0_tmp_reg_10_ ( .D(N1225), .CK(clk), .RN(rstn), .Q(y0_tmp[10]) );
  DFFRHQX1 y0_tmp_reg_9_ ( .D(N1224), .CK(clk), .RN(rstn), .Q(y0_tmp[9]) );
  DFFRHQX1 y0_tmp_reg_8_ ( .D(N1223), .CK(clk), .RN(rstn), .Q(y0_tmp[8]) );
  DFFRHQX1 y0_tmp_reg_7_ ( .D(N1222), .CK(clk), .RN(rstn), .Q(y0_tmp[7]) );
  DFFRHQX1 y1_tmp_reg_11_ ( .D(N1252), .CK(clk), .RN(rstn), .Q(y1_tmp[11]) );
  DFFRHQX1 y1_tmp_reg_10_ ( .D(N1251), .CK(clk), .RN(rstn), .Q(y1_tmp[10]) );
  DFFRHQX1 y1_tmp_reg_9_ ( .D(N1250), .CK(clk), .RN(rstn), .Q(y1_tmp[9]) );
  DFFRHQX1 y1_tmp_reg_8_ ( .D(N1249), .CK(clk), .RN(rstn), .Q(y1_tmp[8]) );
  DFFRHQX1 y1_tmp_reg_7_ ( .D(N1248), .CK(clk), .RN(rstn), .Q(y1_tmp[7]) );
  DFFRHQX1 y2_tmp_reg_11_ ( .D(N1278), .CK(clk), .RN(rstn), .Q(y2_tmp[11]) );
  DFFRHQX1 y2_tmp_reg_10_ ( .D(N1277), .CK(clk), .RN(rstn), .Q(y2_tmp[10]) );
  DFFRHQX1 y2_tmp_reg_9_ ( .D(N1276), .CK(clk), .RN(rstn), .Q(y2_tmp[9]) );
  DFFRHQX1 y2_tmp_reg_8_ ( .D(N1275), .CK(clk), .RN(rstn), .Q(y2_tmp[8]) );
  DFFRHQX1 y2_tmp_reg_7_ ( .D(N1274), .CK(clk), .RN(rstn), .Q(y2_tmp[7]) );
  DFFRHQX1 y3_tmp_reg_11_ ( .D(N1304), .CK(clk), .RN(rstn), .Q(y3_tmp[11]) );
  DFFRHQX1 y3_tmp_reg_10_ ( .D(N1303), .CK(clk), .RN(rstn), .Q(y3_tmp[10]) );
  DFFRHQX1 y3_tmp_reg_9_ ( .D(N1302), .CK(clk), .RN(rstn), .Q(y3_tmp[9]) );
  DFFRHQX1 y3_tmp_reg_8_ ( .D(N1301), .CK(clk), .RN(rstn), .Q(y3_tmp[8]) );
  DFFRHQX1 y3_tmp_reg_7_ ( .D(N1300), .CK(clk), .RN(rstn), .Q(y3_tmp[7]) );
  DFFRHQX1 y4_tmp_reg_9_ ( .D(N1379), .CK(clk), .RN(rstn), .Q(y4_tmp[9]) );
  DFFRHQX1 y4_tmp_reg_8_ ( .D(N1378), .CK(clk), .RN(rstn), .Q(y4_tmp[8]) );
  DFFRHQX1 y4_tmp_reg_7_ ( .D(N1377), .CK(clk), .RN(rstn), .Q(y4_tmp[7]) );
  DFFRHQX1 y5_tmp_reg_9_ ( .D(N1456), .CK(clk), .RN(rstn), .Q(y5_tmp[9]) );
  DFFRHQX1 y5_tmp_reg_8_ ( .D(N1455), .CK(clk), .RN(rstn), .Q(y5_tmp[8]) );
  DFFRHQX1 y5_tmp_reg_7_ ( .D(N1454), .CK(clk), .RN(rstn), .Q(y5_tmp[7]) );
  DFFRHQX1 y6_tmp_reg_6_ ( .D(N1530), .CK(clk), .RN(rstn), .Q(y6_tmp[6]) );
  DFFRHQX1 y7_tmp_reg_6_ ( .D(N1607), .CK(clk), .RN(rstn), .Q(y7_tmp[6]) );
  DFFRHQX1 y0_tmp_reg_6_ ( .D(N1221), .CK(clk), .RN(rstn), .Q(y0_tmp[6]) );
  DFFRHQX1 y1_tmp_reg_6_ ( .D(N1247), .CK(clk), .RN(rstn), .Q(y1_tmp[6]) );
  DFFRHQX1 y2_tmp_reg_6_ ( .D(N1273), .CK(clk), .RN(rstn), .Q(y2_tmp[6]) );
  DFFRHQX1 y3_tmp_reg_6_ ( .D(N1299), .CK(clk), .RN(rstn), .Q(y3_tmp[6]) );
  DFFRHQX1 y4_tmp_reg_6_ ( .D(N1376), .CK(clk), .RN(rstn), .Q(y4_tmp[6]) );
  DFFRHQX1 y5_tmp_reg_6_ ( .D(N1453), .CK(clk), .RN(rstn), .Q(y5_tmp[6]) );
  DFFRHQX1 x7_89_tmp1_reg_5_ ( .D(n40), .CK(clk), .RN(rstn), .Q(x7_89_tmp1[5])
         );
  DFFRHQX1 x7_89_tmp1_reg_4_ ( .D(n39), .CK(clk), .RN(rstn), .Q(x7_89_tmp1[4])
         );
  DFFRHQX1 x7_89_tmp1_reg_3_ ( .D(n38), .CK(clk), .RN(rstn), .Q(x7_89_tmp1[3])
         );
  DFFRHQX1 x7_89_tmp1_reg_2_ ( .D(n37), .CK(clk), .RN(rstn), .Q(x7_89_tmp1[2])
         );
  DFFRHQX1 x6_89_tmp1_reg_5_ ( .D(n53), .CK(clk), .RN(rstn), .Q(x6_89_tmp1[5])
         );
  DFFRHQX1 x6_89_tmp1_reg_4_ ( .D(n52), .CK(clk), .RN(rstn), .Q(x6_89_tmp1[4])
         );
  DFFRHQX1 x6_89_tmp1_reg_3_ ( .D(n51), .CK(clk), .RN(rstn), .Q(x6_89_tmp1[3])
         );
  DFFRHQX1 x6_89_tmp1_reg_2_ ( .D(n50), .CK(clk), .RN(rstn), .Q(x6_89_tmp1[2])
         );
  DFFRHQX1 x5_89_tmp1_reg_5_ ( .D(n66), .CK(clk), .RN(rstn), .Q(x5_89_tmp1[5])
         );
  DFFRHQX1 x5_89_tmp1_reg_4_ ( .D(n65), .CK(clk), .RN(rstn), .Q(x5_89_tmp1[4])
         );
  DFFRHQX1 x5_89_tmp1_reg_3_ ( .D(n64), .CK(clk), .RN(rstn), .Q(x5_89_tmp1[3])
         );
  DFFRHQX1 x5_89_tmp1_reg_2_ ( .D(n63), .CK(clk), .RN(rstn), .Q(x5_89_tmp1[2])
         );
  DFFRHQX1 x5_75_tmp1_reg_5_ ( .D(n66), .CK(clk), .RN(rstn), .Q(x5_75_tmp1[5])
         );
  DFFRHQX1 x5_75_tmp1_reg_4_ ( .D(n65), .CK(clk), .RN(rstn), .Q(x5_75_tmp1[4])
         );
  DFFRHQX1 x5_75_tmp1_reg_3_ ( .D(n64), .CK(clk), .RN(rstn), .Q(x5_75_tmp1[3])
         );
  DFFRHQX1 x5_75_tmp1_reg_2_ ( .D(n63), .CK(clk), .RN(rstn), .Q(x5_75_tmp1[2])
         );
  DFFRHQX1 x4_75_tmp1_reg_5_ ( .D(n79), .CK(clk), .RN(rstn), .Q(x4_75_tmp1[5])
         );
  DFFRHQX1 x4_75_tmp1_reg_4_ ( .D(n78), .CK(clk), .RN(rstn), .Q(x4_75_tmp1[4])
         );
  DFFRHQX1 x4_75_tmp1_reg_3_ ( .D(n77), .CK(clk), .RN(rstn), .Q(x4_75_tmp1[3])
         );
  DFFRHQX1 x4_75_tmp1_reg_2_ ( .D(n76), .CK(clk), .RN(rstn), .Q(x4_75_tmp1[2])
         );
  DFFRHQX1 x7_75_tmp1_reg_5_ ( .D(n40), .CK(clk), .RN(rstn), .Q(x7_75_tmp1[5])
         );
  DFFRHQX1 x7_75_tmp1_reg_4_ ( .D(n39), .CK(clk), .RN(rstn), .Q(x7_75_tmp1[4])
         );
  DFFRHQX1 x7_75_tmp1_reg_3_ ( .D(n38), .CK(clk), .RN(rstn), .Q(x7_75_tmp1[3])
         );
  DFFRHQX1 x7_75_tmp1_reg_2_ ( .D(n37), .CK(clk), .RN(rstn), .Q(x7_75_tmp1[2])
         );
  DFFRHQX1 x6_75_tmp1_reg_5_ ( .D(n53), .CK(clk), .RN(rstn), .Q(x6_75_tmp1[5])
         );
  DFFRHQX1 x6_75_tmp1_reg_4_ ( .D(n52), .CK(clk), .RN(rstn), .Q(x6_75_tmp1[4])
         );
  DFFRHQX1 x6_75_tmp1_reg_3_ ( .D(n51), .CK(clk), .RN(rstn), .Q(x6_75_tmp1[3])
         );
  DFFRHQX1 x6_75_tmp1_reg_2_ ( .D(n50), .CK(clk), .RN(rstn), .Q(x6_75_tmp1[2])
         );
  DFFRHQX1 x5_18_reg_7_ ( .D(N521), .CK(clk), .RN(rstn), .Q(x5_18[7]) );
  DFFRHQX1 x5_18_reg_6_ ( .D(N520), .CK(clk), .RN(rstn), .Q(x5_18[6]) );
  DFFRHQX1 x5_18_reg_5_ ( .D(N519), .CK(clk), .RN(rstn), .Q(x5_18[5]) );
  DFFRHQX1 x5_18_reg_4_ ( .D(N518), .CK(clk), .RN(rstn), .Q(x5_18[4]) );
  DFFRHQX1 x6_18_reg_6_ ( .D(N609), .CK(clk), .RN(rstn), .Q(x6_18[6]) );
  DFFRHQX1 x6_18_reg_5_ ( .D(N608), .CK(clk), .RN(rstn), .Q(x6_18[5]) );
  DFFRHQX1 x6_18_reg_4_ ( .D(N607), .CK(clk), .RN(rstn), .Q(x6_18[4]) );
  DFFRHQX1 x6_18_reg_3_ ( .D(N606), .CK(clk), .RN(rstn), .Q(x6_18[3]) );
  DFFRHQX1 x4_18_reg_6_ ( .D(N431), .CK(clk), .RN(rstn), .Q(x4_18[6]) );
  DFFRHQX1 x4_18_reg_5_ ( .D(N430), .CK(clk), .RN(rstn), .Q(x4_18[5]) );
  DFFRHQX1 x4_18_reg_4_ ( .D(N429), .CK(clk), .RN(rstn), .Q(x4_18[4]) );
  DFFRHQX1 x4_18_reg_3_ ( .D(N428), .CK(clk), .RN(rstn), .Q(x4_18[3]) );
  DFFRHQX1 x4_89_tmp1_reg_5_ ( .D(n79), .CK(clk), .RN(rstn), .Q(x4_89_tmp1[5])
         );
  DFFRHQX1 x4_89_tmp1_reg_4_ ( .D(n78), .CK(clk), .RN(rstn), .Q(x4_89_tmp1[4])
         );
  DFFRHQX1 x4_89_tmp1_reg_3_ ( .D(n77), .CK(clk), .RN(rstn), .Q(x4_89_tmp1[3])
         );
  DFFRHQX1 x4_89_tmp1_reg_2_ ( .D(n76), .CK(clk), .RN(rstn), .Q(x4_89_tmp1[2])
         );
  DFFRHQX1 x4_89_reg_6_ ( .D(N363), .CK(clk), .RN(rstn), .Q(x4_89[6]) );
  DFFRHQX1 x4_89_reg_5_ ( .D(N362), .CK(clk), .RN(rstn), .Q(x4_89[5]) );
  DFFRHQX1 x4_89_reg_4_ ( .D(N361), .CK(clk), .RN(rstn), .Q(x4_89[4]) );
  DFFRHQX1 x4_89_reg_3_ ( .D(N360), .CK(clk), .RN(rstn), .Q(x4_89[3]) );
  DFFRHQX1 x4_75_reg_6_ ( .D(N386), .CK(clk), .RN(rstn), .Q(x4_75[6]) );
  DFFRHQX1 x4_75_reg_5_ ( .D(N385), .CK(clk), .RN(rstn), .Q(x4_75[5]) );
  DFFRHQX1 x4_75_reg_4_ ( .D(N384), .CK(clk), .RN(rstn), .Q(x4_75[4]) );
  DFFRHQX1 x4_75_reg_3_ ( .D(N383), .CK(clk), .RN(rstn), .Q(x4_75[3]) );
  DFFRHQX1 x5_75_reg_6_ ( .D(N475), .CK(clk), .RN(rstn), .Q(x5_75[6]) );
  DFFRHQX1 x5_75_reg_5_ ( .D(N474), .CK(clk), .RN(rstn), .Q(x5_75[5]) );
  DFFRHQX1 x5_75_reg_4_ ( .D(N473), .CK(clk), .RN(rstn), .Q(x5_75[4]) );
  DFFRHQX1 x5_75_reg_3_ ( .D(N472), .CK(clk), .RN(rstn), .Q(x5_75[3]) );
  DFFRHQX1 x6_75_reg_6_ ( .D(N564), .CK(clk), .RN(rstn), .Q(x6_75[6]) );
  DFFRHQX1 x6_75_reg_5_ ( .D(N563), .CK(clk), .RN(rstn), .Q(x6_75[5]) );
  DFFRHQX1 x6_75_reg_4_ ( .D(N562), .CK(clk), .RN(rstn), .Q(x6_75[4]) );
  DFFRHQX1 x6_75_reg_3_ ( .D(N561), .CK(clk), .RN(rstn), .Q(x6_75[3]) );
  DFFRHQX1 x4_50_reg_6_ ( .D(N409), .CK(clk), .RN(rstn), .Q(x4_50[6]) );
  DFFRHQX1 x4_50_reg_5_ ( .D(N408), .CK(clk), .RN(rstn), .Q(x4_50[5]) );
  DFFRHQX1 x4_50_reg_4_ ( .D(N407), .CK(clk), .RN(rstn), .Q(x4_50[4]) );
  DFFRHQX1 x4_50_reg_3_ ( .D(N406), .CK(clk), .RN(rstn), .Q(x4_50[3]) );
  DFFRHQX1 x5_tmp1_reg_7_ ( .D(N886), .CK(clk), .RN(rstn), .Q(x5_tmp1[7]) );
  DFFRHQX1 x5_tmp1_reg_6_ ( .D(N885), .CK(clk), .RN(rstn), .Q(x5_tmp1[6]) );
  DFFRHQX1 x5_tmp1_reg_5_ ( .D(N884), .CK(clk), .RN(rstn), .Q(x5_tmp1[5]) );
  DFFRHQX1 x5_tmp1_reg_4_ ( .D(N883), .CK(clk), .RN(rstn), .Q(x5_tmp1[4]) );
  DFFRHQX1 x6_tmp1_reg_7_ ( .D(N1052), .CK(clk), .RN(rstn), .Q(x6_tmp1[7]) );
  DFFRHQX1 x6_tmp1_reg_6_ ( .D(N1051), .CK(clk), .RN(rstn), .Q(x6_tmp1[6]) );
  DFFRHQX1 x6_tmp1_reg_5_ ( .D(N1050), .CK(clk), .RN(rstn), .Q(x6_tmp1[5]) );
  DFFRHQX1 x6_tmp1_reg_4_ ( .D(N1049), .CK(clk), .RN(rstn), .Q(x6_tmp1[4]) );
  DFFRHQX1 x7_tmp1_reg_7_ ( .D(N1149), .CK(clk), .RN(rstn), .Q(x7_tmp1[7]) );
  DFFRHQX1 x7_tmp1_reg_6_ ( .D(N1148), .CK(clk), .RN(rstn), .Q(x7_tmp1[6]) );
  DFFRHQX1 x7_tmp1_reg_5_ ( .D(N1147), .CK(clk), .RN(rstn), .Q(x7_tmp1[5]) );
  DFFRHQX1 x7_tmp1_reg_4_ ( .D(N1146), .CK(clk), .RN(rstn), .Q(x7_tmp1[4]) );
  DFFRHQX1 x4_tmp1_reg_7_ ( .D(N767), .CK(clk), .RN(rstn), .Q(x4_tmp1[7]) );
  DFFRHQX1 x4_tmp1_reg_6_ ( .D(N766), .CK(clk), .RN(rstn), .Q(x4_tmp1[6]) );
  DFFRHQX1 x4_tmp1_reg_5_ ( .D(N765), .CK(clk), .RN(rstn), .Q(x4_tmp1[5]) );
  DFFRHQX1 x4_tmp1_reg_4_ ( .D(N764), .CK(clk), .RN(rstn), .Q(x4_tmp1[4]) );
  DFFRHQX1 x6_89_reg_0_ ( .D(N535), .CK(clk), .RN(rstn), .Q(x6_89[0]) );
  DFFRHQX1 x7_50_reg_6_ ( .D(N676), .CK(clk), .RN(rstn), .Q(x7_50[6]) );
  DFFRHQX1 x7_50_reg_5_ ( .D(N675), .CK(clk), .RN(rstn), .Q(x7_50[5]) );
  DFFRHQX1 x7_50_reg_4_ ( .D(N674), .CK(clk), .RN(rstn), .Q(x7_50[4]) );
  DFFRHQX1 x7_50_reg_3_ ( .D(N673), .CK(clk), .RN(rstn), .Q(x7_50[3]) );
  DFFRHQX1 x5_89_reg_6_ ( .D(N452), .CK(clk), .RN(rstn), .Q(x5_89[6]) );
  DFFRHQX1 x5_89_reg_5_ ( .D(N451), .CK(clk), .RN(rstn), .Q(x5_89[5]) );
  DFFRHQX1 x5_89_reg_4_ ( .D(N450), .CK(clk), .RN(rstn), .Q(x5_89[4]) );
  DFFRHQX1 x5_89_reg_3_ ( .D(N449), .CK(clk), .RN(rstn), .Q(x5_89[3]) );
  DFFRHQX1 x7_89_reg_6_ ( .D(N630), .CK(clk), .RN(rstn), .Q(x7_89[6]) );
  DFFRHQX1 x7_89_reg_5_ ( .D(N629), .CK(clk), .RN(rstn), .Q(x7_89[5]) );
  DFFRHQX1 x7_89_reg_4_ ( .D(N628), .CK(clk), .RN(rstn), .Q(x7_89[4]) );
  DFFRHQX1 x7_89_reg_3_ ( .D(N627), .CK(clk), .RN(rstn), .Q(x7_89[3]) );
  DFFRHQX1 x5_50_reg_6_ ( .D(N498), .CK(clk), .RN(rstn), .Q(x5_50[6]) );
  DFFRHQX1 x5_50_reg_5_ ( .D(N497), .CK(clk), .RN(rstn), .Q(x5_50[5]) );
  DFFRHQX1 x5_50_reg_4_ ( .D(N496), .CK(clk), .RN(rstn), .Q(x5_50[4]) );
  DFFRHQX1 x5_50_reg_3_ ( .D(N495), .CK(clk), .RN(rstn), .Q(x5_50[3]) );
  DFFRHQX1 x6_89_tmp2_reg_5_ ( .D(N215), .CK(clk), .RN(rstn), .Q(x6_89_tmp2[5]) );
  DFFRHQX1 x6_89_tmp2_reg_4_ ( .D(N214), .CK(clk), .RN(rstn), .Q(x6_89_tmp2[4]) );
  DFFRHQX1 x6_89_tmp2_reg_3_ ( .D(x6[0]), .CK(clk), .RN(rstn), .Q(
        x6_89_tmp2[3]) );
  DFFRHQX1 x5_89_tmp2_reg_5_ ( .D(N130), .CK(clk), .RN(rstn), .Q(x5_89_tmp2[5]) );
  DFFRHQX1 x5_89_tmp2_reg_4_ ( .D(N129), .CK(clk), .RN(rstn), .Q(x5_89_tmp2[4]) );
  DFFRHQX1 x5_89_tmp2_reg_3_ ( .D(x5[0]), .CK(clk), .RN(rstn), .Q(
        x5_89_tmp2[3]) );
  DFFRHQX1 x4_89_tmp2_reg_5_ ( .D(N45), .CK(clk), .RN(rstn), .Q(x4_89_tmp2[5])
         );
  DFFRHQX1 x4_89_tmp2_reg_4_ ( .D(N44), .CK(clk), .RN(rstn), .Q(x4_89_tmp2[4])
         );
  DFFRHQX1 x4_89_tmp2_reg_3_ ( .D(x4[0]), .CK(clk), .RN(rstn), .Q(
        x4_89_tmp2[3]) );
  DFFRHQX1 x7_89_tmp2_reg_5_ ( .D(N300), .CK(clk), .RN(rstn), .Q(x7_89_tmp2[5]) );
  DFFRHQX1 x7_89_tmp2_reg_4_ ( .D(N299), .CK(clk), .RN(rstn), .Q(x7_89_tmp2[4]) );
  DFFRHQX1 x7_89_tmp2_reg_3_ ( .D(x7[0]), .CK(clk), .RN(rstn), .Q(
        x7_89_tmp2[3]) );
  DFFRHQX1 x4_75_tmp2_reg_5_ ( .D(N66), .CK(clk), .RN(rstn), .Q(x4_75_tmp2[5])
         );
  DFFRHQX1 x4_75_tmp2_reg_4_ ( .D(N65), .CK(clk), .RN(rstn), .Q(x4_75_tmp2[4])
         );
  DFFRHQX1 x4_75_tmp2_reg_3_ ( .D(N64), .CK(clk), .RN(rstn), .Q(x4_75_tmp2[3])
         );
  DFFRHQX1 x4_75_tmp2_reg_2_ ( .D(x4[1]), .CK(clk), .RN(rstn), .Q(
        x4_75_tmp2[2]) );
  DFFRHQX1 x4_75_tmp2_reg_1_ ( .D(x4[0]), .CK(clk), .RN(rstn), .Q(
        x4_75_tmp2[1]) );
  DFFRHQX1 x5_75_tmp2_reg_5_ ( .D(N151), .CK(clk), .RN(rstn), .Q(x5_75_tmp2[5]) );
  DFFRHQX1 x5_75_tmp2_reg_4_ ( .D(N150), .CK(clk), .RN(rstn), .Q(x5_75_tmp2[4]) );
  DFFRHQX1 x5_75_tmp2_reg_3_ ( .D(N149), .CK(clk), .RN(rstn), .Q(x5_75_tmp2[3]) );
  DFFRHQX1 x5_75_tmp2_reg_2_ ( .D(x5[1]), .CK(clk), .RN(rstn), .Q(
        x5_75_tmp2[2]) );
  DFFRHQX1 x5_75_tmp2_reg_1_ ( .D(x5[0]), .CK(clk), .RN(rstn), .Q(
        x5_75_tmp2[1]) );
  DFFRHQX1 x6_75_tmp2_reg_5_ ( .D(N236), .CK(clk), .RN(rstn), .Q(x6_75_tmp2[5]) );
  DFFRHQX1 x6_75_tmp2_reg_4_ ( .D(N235), .CK(clk), .RN(rstn), .Q(x6_75_tmp2[4]) );
  DFFRHQX1 x6_75_tmp2_reg_3_ ( .D(N234), .CK(clk), .RN(rstn), .Q(x6_75_tmp2[3]) );
  DFFRHQX1 x6_75_tmp2_reg_2_ ( .D(x6[1]), .CK(clk), .RN(rstn), .Q(
        x6_75_tmp2[2]) );
  DFFRHQX1 x6_75_tmp2_reg_1_ ( .D(x6[0]), .CK(clk), .RN(rstn), .Q(
        x6_75_tmp2[1]) );
  DFFRHQX1 x7_75_tmp2_reg_5_ ( .D(N321), .CK(clk), .RN(rstn), .Q(x7_75_tmp2[5]) );
  DFFRHQX1 x7_75_tmp2_reg_4_ ( .D(N320), .CK(clk), .RN(rstn), .Q(x7_75_tmp2[4]) );
  DFFRHQX1 x7_75_tmp2_reg_3_ ( .D(N319), .CK(clk), .RN(rstn), .Q(x7_75_tmp2[3]) );
  DFFRHQX1 x7_75_tmp2_reg_2_ ( .D(x7[1]), .CK(clk), .RN(rstn), .Q(
        x7_75_tmp2[2]) );
  DFFRHQX1 x7_75_tmp2_reg_1_ ( .D(x7[0]), .CK(clk), .RN(rstn), .Q(
        x7_75_tmp2[1]) );
  DFFRHQX1 x6_50_reg_2_ ( .D(N583), .CK(clk), .RN(rstn), .Q(x6_50[2]) );
  DFFRHQX1 x6_50_reg_3_ ( .D(N584), .CK(clk), .RN(rstn), .Q(x6_50[3]) );
  DFFRHQX1 x6_50_reg_4_ ( .D(N585), .CK(clk), .RN(rstn), .Q(x6_50[4]) );
  DFFRHQX1 x6_50_reg_5_ ( .D(N586), .CK(clk), .RN(rstn), .Q(x6_50[5]) );
  DFFRHQX1 x6_50_reg_6_ ( .D(N587), .CK(clk), .RN(rstn), .Q(x6_50[6]) );
  DFFRHQX1 x7_18_reg_6_ ( .D(N698), .CK(clk), .RN(rstn), .Q(x7_18[6]) );
  DFFRHQX1 x7_18_reg_5_ ( .D(N697), .CK(clk), .RN(rstn), .Q(x7_18[5]) );
  DFFRHQX1 x7_18_reg_4_ ( .D(N696), .CK(clk), .RN(rstn), .Q(x7_18[4]) );
  DFFRHQX1 x7_18_reg_3_ ( .D(N695), .CK(clk), .RN(rstn), .Q(x7_18[3]) );
  DFFRHQX1 x7_18_reg_2_ ( .D(N694), .CK(clk), .RN(rstn), .Q(x7_18[2]) );
  DFFRHQX1 x6_89_reg_7_ ( .D(N542), .CK(clk), .RN(rstn), .Q(x6_89[7]) );
  DFFRHQX1 x6_89_reg_6_ ( .D(N541), .CK(clk), .RN(rstn), .Q(x6_89[6]) );
  DFFRHQX1 x6_89_reg_5_ ( .D(N540), .CK(clk), .RN(rstn), .Q(x6_89[5]) );
  DFFRHQX1 x6_89_reg_4_ ( .D(N539), .CK(clk), .RN(rstn), .Q(x6_89[4]) );
  DFFRHQX1 x7_75_reg_6_ ( .D(N653), .CK(clk), .RN(rstn), .Q(x7_75[6]) );
  DFFRHQX1 x7_75_reg_5_ ( .D(N652), .CK(clk), .RN(rstn), .Q(x7_75[5]) );
  DFFRHQX1 x7_75_reg_4_ ( .D(N651), .CK(clk), .RN(rstn), .Q(x7_75[4]) );
  DFFRHQX1 x7_75_reg_3_ ( .D(N650), .CK(clk), .RN(rstn), .Q(x7_75[3]) );
  DFFRHQX1 x7_75_reg_2_ ( .D(N649), .CK(clk), .RN(rstn), .Q(x7_75[2]) );
  DFFRHQX1 x4_tmp2_reg_7_ ( .D(N837), .CK(clk), .RN(rstn), .Q(x4_tmp2[7]) );
  DFFRHQX1 x4_tmp2_reg_6_ ( .D(N836), .CK(clk), .RN(rstn), .Q(x4_tmp2[6]) );
  DFFRHQX1 x4_tmp2_reg_5_ ( .D(N835), .CK(clk), .RN(rstn), .Q(x4_tmp2[5]) );
  DFFRHQX1 x4_tmp2_reg_4_ ( .D(N834), .CK(clk), .RN(rstn), .Q(x4_tmp2[4]) );
  DFFRHQX1 x4_tmp2_reg_3_ ( .D(N833), .CK(clk), .RN(rstn), .Q(x4_tmp2[3]) );
  DFFRHQX1 x5_tmp2_reg_7_ ( .D(N957), .CK(clk), .RN(rstn), .Q(x5_tmp2[7]) );
  DFFRHQX1 x5_tmp2_reg_6_ ( .D(N956), .CK(clk), .RN(rstn), .Q(x5_tmp2[6]) );
  DFFRHQX1 x5_tmp2_reg_5_ ( .D(N955), .CK(clk), .RN(rstn), .Q(x5_tmp2[5]) );
  DFFRHQX1 x5_tmp2_reg_4_ ( .D(N954), .CK(clk), .RN(rstn), .Q(x5_tmp2[4]) );
  DFFRHQX1 x5_tmp2_reg_3_ ( .D(N953), .CK(clk), .RN(rstn), .Q(x5_tmp2[3]) );
  DFFRHQX1 x6_tmp2_reg_7_ ( .D(N1100), .CK(clk), .RN(rstn), .Q(x6_tmp2[7]) );
  DFFRHQX1 x6_tmp2_reg_6_ ( .D(N1099), .CK(clk), .RN(rstn), .Q(x6_tmp2[6]) );
  DFFRHQX1 x6_tmp2_reg_5_ ( .D(N1098), .CK(clk), .RN(rstn), .Q(x6_tmp2[5]) );
  DFFRHQX1 x6_tmp2_reg_4_ ( .D(N1097), .CK(clk), .RN(rstn), .Q(x6_tmp2[4]) );
  DFFRHQX1 x6_tmp2_reg_3_ ( .D(N1096), .CK(clk), .RN(rstn), .Q(x6_tmp2[3]) );
  DFFRHQX1 x7_tmp2_reg_7_ ( .D(N1173), .CK(clk), .RN(rstn), .Q(x7_tmp2[7]) );
  DFFRHQX1 x7_tmp2_reg_6_ ( .D(N1172), .CK(clk), .RN(rstn), .Q(x7_tmp2[6]) );
  DFFRHQX1 x7_tmp2_reg_5_ ( .D(N1171), .CK(clk), .RN(rstn), .Q(x7_tmp2[5]) );
  DFFRHQX1 x7_tmp2_reg_4_ ( .D(N1170), .CK(clk), .RN(rstn), .Q(x7_tmp2[4]) );
  DFFRHQX1 x7_tmp2_reg_3_ ( .D(N1169), .CK(clk), .RN(rstn), .Q(x7_tmp2[3]) );
  DFFRHQX1 x7_tmp_reg_5_ ( .D(N1195), .CK(clk), .RN(rstn), .Q(x7_tmp[5]) );
  DFFRHQX1 x7_tmp_reg_6_ ( .D(N1196), .CK(clk), .RN(rstn), .Q(x7_tmp[6]) );
  DFFRHQX1 x7_tmp_reg_7_ ( .D(N1197), .CK(clk), .RN(rstn), .Q(x7_tmp[7]) );
  DFFRHQX1 x7_tmp_reg_8_ ( .D(N1198), .CK(clk), .RN(rstn), .Q(x7_tmp[8]) );
  DFFRHQX1 x7_tmp_reg_9_ ( .D(N1199), .CK(clk), .RN(rstn), .Q(x7_tmp[9]) );
  DFFRHQX1 x5_tmp_reg_9_ ( .D(N983), .CK(clk), .RN(rstn), .Q(x5_tmp[9]) );
  DFFRHQX1 x5_tmp_reg_8_ ( .D(N982), .CK(clk), .RN(rstn), .Q(x5_tmp[8]) );
  DFFRHQX1 x5_tmp_reg_7_ ( .D(N981), .CK(clk), .RN(rstn), .Q(x5_tmp[7]) );
  DFFRHQX1 x5_tmp_reg_6_ ( .D(N980), .CK(clk), .RN(rstn), .Q(x5_tmp[6]) );
  DFFRHQX1 x5_tmp_reg_5_ ( .D(N979), .CK(clk), .RN(rstn), .Q(x5_tmp[5]) );
  DFFRHQX1 x6_tmp_reg_9_ ( .D(N1126), .CK(clk), .RN(rstn), .Q(x6_tmp[9]) );
  DFFRHQX1 x6_tmp_reg_8_ ( .D(N1125), .CK(clk), .RN(rstn), .Q(x6_tmp[8]) );
  DFFRHQX1 x6_tmp_reg_7_ ( .D(N1124), .CK(clk), .RN(rstn), .Q(x6_tmp[7]) );
  DFFRHQX1 x6_tmp_reg_6_ ( .D(N1123), .CK(clk), .RN(rstn), .Q(x6_tmp[6]) );
  DFFRHQX1 x6_tmp_reg_5_ ( .D(N1122), .CK(clk), .RN(rstn), .Q(x6_tmp[5]) );
  DFFRHQX1 x4_tmp_reg_5_ ( .D(N859), .CK(clk), .RN(rstn), .Q(x4_tmp[5]) );
  DFFRHQX1 x4_tmp_reg_6_ ( .D(N860), .CK(clk), .RN(rstn), .Q(x4_tmp[6]) );
  DFFRHQX1 x4_tmp_reg_7_ ( .D(N861), .CK(clk), .RN(rstn), .Q(x4_tmp[7]) );
  DFFRHQX1 x4_tmp_reg_8_ ( .D(N862), .CK(clk), .RN(rstn), .Q(x4_tmp[8]) );
  DFFRHQX1 x4_tmp_reg_9_ ( .D(N863), .CK(clk), .RN(rstn), .Q(x4_tmp[9]) );
  DFFRHQX1 x7_89_tmp1_reg_1_ ( .D(x7[1]), .CK(clk), .RN(rstn), .Q(
        x7_89_tmp1[1]) );
  DFFRHQX1 x6_89_tmp1_reg_1_ ( .D(x6[1]), .CK(clk), .RN(rstn), .Q(
        x6_89_tmp1[1]) );
  DFFRHQX1 x5_89_tmp1_reg_1_ ( .D(x5[1]), .CK(clk), .RN(rstn), .Q(
        x5_89_tmp1[1]) );
  DFFRHQX1 x5_75_tmp1_reg_1_ ( .D(x5[1]), .CK(clk), .RN(rstn), .Q(
        x5_75_tmp1[1]) );
  DFFRHQX1 x4_75_tmp1_reg_1_ ( .D(x4[1]), .CK(clk), .RN(rstn), .Q(
        x4_75_tmp1[1]) );
  DFFRHQX1 x7_75_tmp1_reg_1_ ( .D(x7[1]), .CK(clk), .RN(rstn), .Q(
        x7_75_tmp1[1]) );
  DFFRHQX1 x6_75_tmp1_reg_1_ ( .D(x6[1]), .CK(clk), .RN(rstn), .Q(
        x6_75_tmp1[1]) );
  DFFRHQX1 x5_18_reg_3_ ( .D(N517), .CK(clk), .RN(rstn), .Q(x5_18[3]) );
  DFFRHQX1 x5_18_reg_2_ ( .D(N516), .CK(clk), .RN(rstn), .Q(x5_18[2]) );
  DFFRHQX1 x5_18_reg_1_ ( .D(N515), .CK(clk), .RN(rstn), .Q(x5_18[1]) );
  DFFRHQX1 x6_18_reg_2_ ( .D(N605), .CK(clk), .RN(rstn), .Q(x6_18[2]) );
  DFFRHQX1 x6_18_reg_1_ ( .D(N604), .CK(clk), .RN(rstn), .Q(x6_18[1]) );
  DFFRHQX1 x4_18_reg_2_ ( .D(N427), .CK(clk), .RN(rstn), .Q(x4_18[2]) );
  DFFRHQX1 x4_18_reg_1_ ( .D(N426), .CK(clk), .RN(rstn), .Q(x4_18[1]) );
  DFFRHQX1 x4_89_tmp1_reg_1_ ( .D(x4[1]), .CK(clk), .RN(rstn), .Q(
        x4_89_tmp1[1]) );
  DFFRHQX1 x4_89_reg_2_ ( .D(N359), .CK(clk), .RN(rstn), .Q(x4_89[2]) );
  DFFRHQX1 x4_89_reg_1_ ( .D(N358), .CK(clk), .RN(rstn), .Q(x4_89[1]) );
  DFFRHQX1 x4_75_reg_2_ ( .D(N382), .CK(clk), .RN(rstn), .Q(x4_75[2]) );
  DFFRHQX1 x4_75_reg_1_ ( .D(N381), .CK(clk), .RN(rstn), .Q(x4_75[1]) );
  DFFRHQX1 x5_75_reg_2_ ( .D(N471), .CK(clk), .RN(rstn), .Q(x5_75[2]) );
  DFFRHQX1 x5_75_reg_1_ ( .D(N470), .CK(clk), .RN(rstn), .Q(x5_75[1]) );
  DFFRHQX1 x6_75_reg_2_ ( .D(N560), .CK(clk), .RN(rstn), .Q(x6_75[2]) );
  DFFRHQX1 x6_75_reg_1_ ( .D(N559), .CK(clk), .RN(rstn), .Q(x6_75[1]) );
  DFFRHQX1 x4_50_reg_2_ ( .D(N405), .CK(clk), .RN(rstn), .Q(x4_50[2]) );
  DFFRHQX1 x4_50_reg_1_ ( .D(N404), .CK(clk), .RN(rstn), .Q(x4_50[1]) );
  DFFRHQX1 x5_tmp1_reg_3_ ( .D(N882), .CK(clk), .RN(rstn), .Q(x5_tmp1[3]) );
  DFFRHQX1 x5_tmp1_reg_2_ ( .D(N881), .CK(clk), .RN(rstn), .Q(x5_tmp1[2]) );
  DFFRHQX1 x5_tmp1_reg_1_ ( .D(N880), .CK(clk), .RN(rstn), .Q(x5_tmp1[1]) );
  DFFRHQX1 x6_tmp1_reg_3_ ( .D(N1048), .CK(clk), .RN(rstn), .Q(x6_tmp1[3]) );
  DFFRHQX1 x6_tmp1_reg_2_ ( .D(N1047), .CK(clk), .RN(rstn), .Q(x6_tmp1[2]) );
  DFFRHQX1 x6_tmp1_reg_1_ ( .D(N1046), .CK(clk), .RN(rstn), .Q(x6_tmp1[1]) );
  DFFRHQX1 x7_tmp1_reg_3_ ( .D(N1145), .CK(clk), .RN(rstn), .Q(x7_tmp1[3]) );
  DFFRHQX1 x7_tmp1_reg_2_ ( .D(N1144), .CK(clk), .RN(rstn), .Q(x7_tmp1[2]) );
  DFFRHQX1 x7_tmp1_reg_1_ ( .D(N1143), .CK(clk), .RN(rstn), .Q(x7_tmp1[1]) );
  DFFRHQX1 x4_tmp1_reg_3_ ( .D(N763), .CK(clk), .RN(rstn), .Q(x4_tmp1[3]) );
  DFFRHQX1 x4_tmp1_reg_2_ ( .D(N762), .CK(clk), .RN(rstn), .Q(x4_tmp1[2]) );
  DFFRHQX1 x4_tmp1_reg_1_ ( .D(N761), .CK(clk), .RN(rstn), .Q(x4_tmp1[1]) );
  DFFRHQX1 x7_50_reg_2_ ( .D(N672), .CK(clk), .RN(rstn), .Q(x7_50[2]) );
  DFFRHQX1 x7_50_reg_1_ ( .D(N671), .CK(clk), .RN(rstn), .Q(x7_50[1]) );
  DFFRHQX1 x7_50_reg_0_ ( .D(1'b0), .CK(clk), .RN(rstn), .Q(x7_50[0]) );
  DFFRHQX1 x5_89_reg_2_ ( .D(N448), .CK(clk), .RN(rstn), .Q(x5_89[2]) );
  DFFRHQX1 x5_89_reg_1_ ( .D(N447), .CK(clk), .RN(rstn), .Q(x5_89[1]) );
  DFFRHQX1 x5_89_reg_0_ ( .D(N446), .CK(clk), .RN(rstn), .Q(x5_89[0]) );
  DFFRHQX1 x7_89_reg_2_ ( .D(N626), .CK(clk), .RN(rstn), .Q(x7_89[2]) );
  DFFRHQX1 x7_89_reg_1_ ( .D(N625), .CK(clk), .RN(rstn), .Q(x7_89[1]) );
  DFFRHQX1 x7_89_reg_0_ ( .D(N624), .CK(clk), .RN(rstn), .Q(x7_89[0]) );
  DFFRHQX1 x5_50_reg_2_ ( .D(N494), .CK(clk), .RN(rstn), .Q(x5_50[2]) );
  DFFRHQX1 x5_50_reg_1_ ( .D(N493), .CK(clk), .RN(rstn), .Q(x5_50[1]) );
  DFFRHQX1 x5_50_reg_0_ ( .D(1'b0), .CK(clk), .RN(rstn), .Q(x5_50[0]) );
  DFFRHQX1 x6_50_reg_1_ ( .D(N582), .CK(clk), .RN(rstn), .Q(x6_50[1]) );
  DFFRHQX1 x7_18_reg_1_ ( .D(N693), .CK(clk), .RN(rstn), .Q(x7_18[1]) );
  DFFRHQX1 x6_89_reg_3_ ( .D(N538), .CK(clk), .RN(rstn), .Q(x6_89[3]) );
  DFFRHQX1 x6_89_reg_2_ ( .D(N537), .CK(clk), .RN(rstn), .Q(x6_89[2]) );
  DFFRHQX1 x6_89_reg_1_ ( .D(N536), .CK(clk), .RN(rstn), .Q(x6_89[1]) );
  DFFRHQX1 x7_75_reg_1_ ( .D(N648), .CK(clk), .RN(rstn), .Q(x7_75[1]) );
  DFFRHQX1 x4_tmp2_reg_2_ ( .D(N832), .CK(clk), .RN(rstn), .Q(x4_tmp2[2]) );
  DFFRHQX1 x4_tmp2_reg_1_ ( .D(N831), .CK(clk), .RN(rstn), .Q(x4_tmp2[1]) );
  DFFRHQX1 x5_tmp2_reg_2_ ( .D(N952), .CK(clk), .RN(rstn), .Q(x5_tmp2[2]) );
  DFFRHQX1 x5_tmp2_reg_1_ ( .D(N951), .CK(clk), .RN(rstn), .Q(x5_tmp2[1]) );
  DFFRHQX1 x6_tmp2_reg_2_ ( .D(N1095), .CK(clk), .RN(rstn), .Q(x6_tmp2[2]) );
  DFFRHQX1 x6_tmp2_reg_1_ ( .D(N1094), .CK(clk), .RN(rstn), .Q(x6_tmp2[1]) );
  DFFRHQX1 x7_tmp2_reg_2_ ( .D(N1168), .CK(clk), .RN(rstn), .Q(x7_tmp2[2]) );
  DFFRHQX1 x7_tmp2_reg_1_ ( .D(N1167), .CK(clk), .RN(rstn), .Q(x7_tmp2[1]) );
  DFFRHQX1 x6_50_reg_0_ ( .D(1'b0), .CK(clk), .RN(rstn), .Q(x6_50[0]) );
  DFFRHQX1 x7_75_reg_0_ ( .D(N647), .CK(clk), .RN(rstn), .Q(x7_75[0]) );
  DFFRHQX1 x4_tmp2_reg_0_ ( .D(N830), .CK(clk), .RN(rstn), .Q(x4_tmp2[0]) );
  DFFRHQX1 x5_tmp2_reg_0_ ( .D(N950), .CK(clk), .RN(rstn), .Q(x5_tmp2[0]) );
  DFFRHQX1 x6_tmp2_reg_0_ ( .D(N1093), .CK(clk), .RN(rstn), .Q(x6_tmp2[0]) );
  DFFRHQX1 x7_tmp2_reg_0_ ( .D(N1166), .CK(clk), .RN(rstn), .Q(x7_tmp2[0]) );
  DFFRHQX1 x5_75_reg_0_ ( .D(N469), .CK(clk), .RN(rstn), .Q(x5_75[0]) );
  DFFRHQX1 x4_50_reg_0_ ( .D(1'b0), .CK(clk), .RN(rstn), .Q(x4_50[0]) );
  DFFRHQX1 x5_tmp1_reg_0_ ( .D(N879), .CK(clk), .RN(rstn), .Q(x5_tmp1[0]) );
  DFFRHQX1 x6_tmp1_reg_0_ ( .D(N1045), .CK(clk), .RN(rstn), .Q(x6_tmp1[0]) );
  DFFRHQX1 x7_tmp1_reg_0_ ( .D(N1142), .CK(clk), .RN(rstn), .Q(x7_tmp1[0]) );
  DFFRHQX1 x4_tmp1_reg_0_ ( .D(N760), .CK(clk), .RN(rstn), .Q(x4_tmp1[0]) );
  DFFRHQX1 x7_tmp_reg_1_ ( .D(N1191), .CK(clk), .RN(rstn), .Q(x7_tmp[1]) );
  DFFRHQX1 x7_tmp_reg_2_ ( .D(N1192), .CK(clk), .RN(rstn), .Q(x7_tmp[2]) );
  DFFRHQX1 x7_tmp_reg_3_ ( .D(N1193), .CK(clk), .RN(rstn), .Q(x7_tmp[3]) );
  DFFRHQX1 x7_tmp_reg_4_ ( .D(N1194), .CK(clk), .RN(rstn), .Q(x7_tmp[4]) );
  DFFRHQX1 x5_tmp_reg_4_ ( .D(N978), .CK(clk), .RN(rstn), .Q(x5_tmp[4]) );
  DFFRHQX1 x5_tmp_reg_3_ ( .D(N977), .CK(clk), .RN(rstn), .Q(x5_tmp[3]) );
  DFFRHQX1 x5_tmp_reg_2_ ( .D(N976), .CK(clk), .RN(rstn), .Q(x5_tmp[2]) );
  DFFRHQX1 x5_tmp_reg_1_ ( .D(N975), .CK(clk), .RN(rstn), .Q(x5_tmp[1]) );
  DFFRHQX1 x6_tmp_reg_4_ ( .D(N1121), .CK(clk), .RN(rstn), .Q(x6_tmp[4]) );
  DFFRHQX1 x6_tmp_reg_3_ ( .D(N1120), .CK(clk), .RN(rstn), .Q(x6_tmp[3]) );
  DFFRHQX1 x6_tmp_reg_2_ ( .D(N1119), .CK(clk), .RN(rstn), .Q(x6_tmp[2]) );
  DFFRHQX1 x6_tmp_reg_1_ ( .D(N1118), .CK(clk), .RN(rstn), .Q(x6_tmp[1]) );
  DFFRHQX1 x4_tmp_reg_1_ ( .D(N855), .CK(clk), .RN(rstn), .Q(x4_tmp[1]) );
  DFFRHQX1 x4_tmp_reg_2_ ( .D(N856), .CK(clk), .RN(rstn), .Q(x4_tmp[2]) );
  DFFRHQX1 x4_tmp_reg_3_ ( .D(N857), .CK(clk), .RN(rstn), .Q(x4_tmp[3]) );
  DFFRHQX1 x4_tmp_reg_4_ ( .D(N858), .CK(clk), .RN(rstn), .Q(x4_tmp[4]) );
  DFFRHQX1 x4_75_reg_0_ ( .D(N380), .CK(clk), .RN(rstn), .Q(x4_75[0]) );
  DFFRHQX1 x6_75_reg_0_ ( .D(N558), .CK(clk), .RN(rstn), .Q(x6_75[0]) );
  DFFRHQX1 x7_tmp_reg_0_ ( .D(N1190), .CK(clk), .RN(rstn), .Q(x7_tmp[0]) );
  DFFRHQX1 x5_tmp_reg_0_ ( .D(N974), .CK(clk), .RN(rstn), .Q(x5_tmp[0]) );
  DFFRHQX1 x6_tmp_reg_0_ ( .D(N1117), .CK(clk), .RN(rstn), .Q(x6_tmp[0]) );
  DFFRHQX1 x4_tmp_reg_0_ ( .D(N854), .CK(clk), .RN(rstn), .Q(x4_tmp[0]) );
  DFFRHQX1 mode_delay1_reg_1_ ( .D(mode[1]), .CK(clk), .RN(rstn), .Q(
        mode_delay1[1]) );
  DFFRHQX1 mode_delay1_reg_0_ ( .D(mode[0]), .CK(clk), .RN(rstn), .Q(
        mode_delay1[0]) );
  INVX1 U48 ( .A(n177), .Y(n89) );
  INVX1 U49 ( .A(n177), .Y(n92) );
  INVX1 U50 ( .A(n177), .Y(n90) );
  INVX1 U51 ( .A(n177), .Y(n91) );
  AND2X2 U52 ( .A(y0_tmp[25]), .B(n202), .Y(y0[25]) );
  AND2X2 U53 ( .A(y1_tmp[25]), .B(n209), .Y(y1[25]) );
  AND2X2 U54 ( .A(y2_tmp[25]), .B(n210), .Y(y2[25]) );
  AND2X2 U55 ( .A(y3_tmp[25]), .B(n211), .Y(y3[25]) );
  AND2X2 U56 ( .A(y4_tmp[25]), .B(n202), .Y(y4[25]) );
  AND2X2 U57 ( .A(y5_tmp[25]), .B(n103), .Y(y5[25]) );
  AND2X2 U58 ( .A(y6_tmp[25]), .B(n199), .Y(y6[25]) );
  AND2X2 U59 ( .A(y7_tmp[25]), .B(n198), .Y(y7[25]) );
  AND2X2 U60 ( .A(y1_tmp[22]), .B(n103), .Y(y1[22]) );
  AND2X2 U61 ( .A(y1_tmp[23]), .B(n103), .Y(y1[23]) );
  AND2X2 U62 ( .A(y1_tmp[24]), .B(n103), .Y(y1[24]) );
  AND2X2 U94 ( .A(y2_tmp[22]), .B(n103), .Y(y2[22]) );
  AND2X2 U95 ( .A(y2_tmp[24]), .B(n103), .Y(y2[24]) );
  AND2X2 U96 ( .A(y4_tmp[22]), .B(n103), .Y(y4[22]) );
  AND2X2 U97 ( .A(y4_tmp[24]), .B(n103), .Y(y4[24]) );
  AND2X2 U98 ( .A(y5_tmp[22]), .B(n103), .Y(y5[22]) );
  AND2X2 U99 ( .A(y5_tmp[23]), .B(n103), .Y(y5[23]) );
  AND2X2 U100 ( .A(y5_tmp[24]), .B(n103), .Y(y5[24]) );
  AND2X2 U101 ( .A(y6_tmp[22]), .B(n103), .Y(y6[22]) );
  AND2X2 U102 ( .A(y0_tmp[22]), .B(n205), .Y(y0[22]) );
  AND2X2 U103 ( .A(y0_tmp[23]), .B(n206), .Y(y0[23]) );
  AND2X2 U104 ( .A(y0_tmp[24]), .B(n209), .Y(y0[24]) );
  AND2X2 U105 ( .A(y2_tmp[23]), .B(n210), .Y(y2[23]) );
  AND2X2 U106 ( .A(y3_tmp[22]), .B(n211), .Y(y3[22]) );
  AND2X2 U107 ( .A(y3_tmp[23]), .B(n208), .Y(y3[23]) );
  AND2X2 U108 ( .A(y3_tmp[24]), .B(n202), .Y(y3[24]) );
  AND2X2 U109 ( .A(y4_tmp[23]), .B(n199), .Y(y4[23]) );
  AND2X2 U110 ( .A(y6_tmp[23]), .B(n198), .Y(y6[23]) );
  AND2X2 U111 ( .A(y6_tmp[24]), .B(n205), .Y(y6[24]) );
  AND2X2 U112 ( .A(y7_tmp[22]), .B(n206), .Y(y7[22]) );
  AND2X2 U113 ( .A(y7_tmp[23]), .B(n209), .Y(y7[23]) );
  AND2X2 U114 ( .A(y7_tmp[24]), .B(n210), .Y(y7[24]) );
  INVX1 U115 ( .A(n180), .Y(n103) );
  INVX1 U116 ( .A(n179), .Y(n98) );
  INVX1 U117 ( .A(n179), .Y(n99) );
  INVX1 U118 ( .A(n179), .Y(n100) );
  INVX1 U119 ( .A(n180), .Y(n102) );
  INVX1 U120 ( .A(n178), .Y(n96) );
  INVX1 U121 ( .A(n179), .Y(n97) );
  INVX1 U122 ( .A(n180), .Y(n101) );
  INVX1 U123 ( .A(n182), .Y(n177) );
  INVX1 U124 ( .A(n178), .Y(n95) );
  INVX1 U125 ( .A(n178), .Y(n94) );
  INVX1 U126 ( .A(n178), .Y(n93) );
  INVX1 U127 ( .A(n211), .Y(n105) );
  INVX1 U128 ( .A(n211), .Y(n104) );
  INVX1 U129 ( .A(n184), .Y(n171) );
  INVX1 U130 ( .A(n184), .Y(n170) );
  INVX1 U131 ( .A(n185), .Y(n169) );
  INVX1 U132 ( .A(n185), .Y(n168) );
  INVX1 U133 ( .A(n185), .Y(n167) );
  INVX1 U134 ( .A(n182), .Y(n176) );
  INVX1 U135 ( .A(n182), .Y(n175) );
  INVX1 U136 ( .A(n183), .Y(n174) );
  INVX1 U137 ( .A(n183), .Y(n173) );
  INVX1 U138 ( .A(n187), .Y(n162) );
  INVX1 U139 ( .A(n188), .Y(n161) );
  INVX1 U140 ( .A(n188), .Y(n160) );
  INVX1 U141 ( .A(n189), .Y(n159) );
  INVX1 U142 ( .A(n189), .Y(n158) );
  INVX1 U143 ( .A(n186), .Y(n166) );
  INVX1 U144 ( .A(n186), .Y(n165) );
  INVX1 U145 ( .A(n186), .Y(n164) );
  INVX1 U146 ( .A(n187), .Y(n163) );
  INVX1 U147 ( .A(n191), .Y(n153) );
  INVX1 U148 ( .A(n192), .Y(n152) );
  INVX1 U149 ( .A(n192), .Y(n151) );
  INVX1 U150 ( .A(n192), .Y(n150) );
  INVX1 U151 ( .A(n193), .Y(n149) );
  INVX1 U152 ( .A(n189), .Y(n157) );
  INVX1 U153 ( .A(n190), .Y(n156) );
  INVX1 U154 ( .A(n190), .Y(n155) );
  INVX1 U155 ( .A(n190), .Y(n154) );
  INVX1 U156 ( .A(n195), .Y(n144) );
  INVX1 U157 ( .A(n195), .Y(n143) );
  INVX1 U158 ( .A(n196), .Y(n142) );
  INVX1 U159 ( .A(n196), .Y(n141) );
  INVX1 U160 ( .A(n196), .Y(n140) );
  INVX1 U161 ( .A(n193), .Y(n148) );
  INVX1 U162 ( .A(n193), .Y(n147) );
  INVX1 U163 ( .A(n194), .Y(n146) );
  INVX1 U164 ( .A(n194), .Y(n145) );
  INVX1 U165 ( .A(n198), .Y(n135) );
  INVX1 U166 ( .A(n199), .Y(n134) );
  INVX1 U167 ( .A(n199), .Y(n133) );
  INVX1 U168 ( .A(n200), .Y(n132) );
  INVX1 U169 ( .A(n200), .Y(n131) );
  INVX1 U170 ( .A(n197), .Y(n139) );
  INVX1 U171 ( .A(n197), .Y(n138) );
  INVX1 U172 ( .A(n197), .Y(n137) );
  INVX1 U173 ( .A(n198), .Y(n136) );
  INVX1 U174 ( .A(n202), .Y(n126) );
  INVX1 U175 ( .A(n203), .Y(n125) );
  INVX1 U176 ( .A(n203), .Y(n124) );
  INVX1 U177 ( .A(n203), .Y(n123) );
  INVX1 U178 ( .A(n204), .Y(n122) );
  INVX1 U179 ( .A(n200), .Y(n130) );
  INVX1 U180 ( .A(n201), .Y(n129) );
  INVX1 U181 ( .A(n201), .Y(n128) );
  INVX1 U182 ( .A(n201), .Y(n127) );
  INVX1 U183 ( .A(n206), .Y(n117) );
  INVX1 U184 ( .A(n206), .Y(n116) );
  INVX1 U185 ( .A(n207), .Y(n115) );
  INVX1 U186 ( .A(n207), .Y(n114) );
  INVX1 U187 ( .A(n207), .Y(n113) );
  INVX1 U188 ( .A(n204), .Y(n121) );
  INVX1 U189 ( .A(n204), .Y(n120) );
  INVX1 U190 ( .A(n205), .Y(n119) );
  INVX1 U191 ( .A(n205), .Y(n118) );
  INVX1 U192 ( .A(n209), .Y(n108) );
  INVX1 U193 ( .A(n210), .Y(n107) );
  INVX1 U194 ( .A(n210), .Y(n106) );
  INVX1 U195 ( .A(n208), .Y(n112) );
  INVX1 U196 ( .A(n208), .Y(n111) );
  INVX1 U197 ( .A(n208), .Y(n110) );
  INVX1 U198 ( .A(n209), .Y(n109) );
  INVX1 U199 ( .A(n183), .Y(n172) );
  ADDFX2 U200 ( .A(x7[15]), .B(x7[15]), .CI(N355), .CO(N356) );
  ADDFX2 U201 ( .A(x5[15]), .B(x5[15]), .CI(N185), .CO(N186) );
  ADDFX2 U202 ( .A(x6[15]), .B(x6[15]), .CI(N270), .CO(N271) );
  ADDFX2 U203 ( .A(x4[15]), .B(x4[15]), .CI(N100), .CO(N101) );
  ADDFX2 U204 ( .A(x7[15]), .B(x7[15]), .CI(N334), .CO(N335) );
  ADDFX2 U205 ( .A(x6[15]), .B(x6[15]), .CI(N249), .CO(N250) );
  ADDFX2 U206 ( .A(x5[15]), .B(x5[15]), .CI(N164), .CO(N165) );
  ADDFX2 U207 ( .A(x4[15]), .B(x4[15]), .CI(N79), .CO(N80) );
  ADDFX2 U208 ( .A(x7[15]), .B(x7[15]), .CI(N314), .CO(N315) );
  ADDFX2 U209 ( .A(x4[15]), .B(x4[15]), .CI(N59), .CO(N60) );
  ADDFX2 U210 ( .A(x5[15]), .B(x5[15]), .CI(N144), .CO(N145) );
  ADDFX2 U211 ( .A(x6[15]), .B(x6[15]), .CI(N229), .CO(N230) );
  INVX1 U212 ( .A(n181), .Y(n179) );
  INVX1 U213 ( .A(n181), .Y(n178) );
  INVX1 U214 ( .A(n181), .Y(n180) );
  INVX1 U215 ( .A(n221), .Y(n182) );
  INVX1 U216 ( .A(n221), .Y(n184) );
  INVX1 U217 ( .A(n220), .Y(n185) );
  INVX1 U218 ( .A(n221), .Y(n183) );
  INVX1 U219 ( .A(n219), .Y(n188) );
  INVX1 U220 ( .A(n220), .Y(n186) );
  INVX1 U221 ( .A(n220), .Y(n187) );
  INVX1 U222 ( .A(n218), .Y(n192) );
  INVX1 U223 ( .A(n219), .Y(n189) );
  INVX1 U224 ( .A(n219), .Y(n190) );
  INVX1 U225 ( .A(n217), .Y(n195) );
  INVX1 U226 ( .A(n217), .Y(n196) );
  INVX1 U227 ( .A(n218), .Y(n193) );
  INVX1 U228 ( .A(n217), .Y(n194) );
  INVX1 U229 ( .A(n216), .Y(n199) );
  INVX1 U230 ( .A(n216), .Y(n197) );
  INVX1 U231 ( .A(n216), .Y(n198) );
  INVX1 U232 ( .A(n214), .Y(n203) );
  INVX1 U233 ( .A(n215), .Y(n200) );
  INVX1 U234 ( .A(n215), .Y(n201) );
  INVX1 U235 ( .A(n213), .Y(n206) );
  INVX1 U236 ( .A(n213), .Y(n207) );
  INVX1 U237 ( .A(n214), .Y(n204) );
  INVX1 U238 ( .A(n214), .Y(n205) );
  INVX1 U239 ( .A(n212), .Y(n210) );
  INVX1 U240 ( .A(n213), .Y(n208) );
  INVX1 U241 ( .A(n212), .Y(n209) );
  INVX1 U242 ( .A(n218), .Y(n191) );
  INVX1 U243 ( .A(n215), .Y(n202) );
  INVX1 U244 ( .A(n212), .Y(n211) );
  ADDFX2 U245 ( .A(n49), .B(x7[15]), .CI(add_104_carry_18_), .CO(N355), .S(
        N354) );
  ADDFX2 U246 ( .A(n75), .B(x5[15]), .CI(add_86_carry_18_), .CO(N185), .S(N184) );
  ADDFX2 U247 ( .A(n62), .B(x6[15]), .CI(add_95_carry_18_), .CO(N270), .S(N269) );
  ADDFX2 U248 ( .A(n88), .B(x4[15]), .CI(add_77_carry_18_), .CO(N100), .S(N99)
         );
  ADDFX2 U249 ( .A(n49), .B(x7[15]), .CI(add_102_carry_17_), .CO(N334), .S(
        N333) );
  ADDFX2 U250 ( .A(n62), .B(x6[15]), .CI(add_93_carry_17_), .CO(N249), .S(N248) );
  ADDFX2 U251 ( .A(n75), .B(x5[15]), .CI(add_84_carry_17_), .CO(N164), .S(N163) );
  ADDFX2 U252 ( .A(n88), .B(x4[15]), .CI(add_75_carry_17_), .CO(N79), .S(N78)
         );
  ADDFX2 U253 ( .A(n49), .B(x7[15]), .CI(add_100_carry_18_), .CO(N314), .S(
        N313) );
  ADDFX2 U254 ( .A(n88), .B(x4[15]), .CI(add_73_carry_18_), .CO(N59), .S(N58)
         );
  ADDFX2 U255 ( .A(n75), .B(x5[15]), .CI(add_82_carry_18_), .CO(N144), .S(N143) );
  ADDFX2 U256 ( .A(n62), .B(x6[15]), .CI(add_91_carry_18_), .CO(N229), .S(N228) );
  ADDFX2 U257 ( .A(n88), .B(x4[15]), .CI(add_72_carry_20_), .CO(N38), .S(N37)
         );
  ADDFX2 U258 ( .A(n75), .B(x5[15]), .CI(add_81_carry_20_), .CO(N123), .S(N122) );
  ADDFX2 U259 ( .A(n62), .B(x6[15]), .CI(add_90_carry_20_), .CO(N208), .S(N207) );
  ADDFX2 U260 ( .A(n49), .B(x7[15]), .CI(add_99_carry_20_), .CO(N293), .S(N292) );
  ADDFX2 U261 ( .A(n37), .B(n40), .CI(add_104_carry_6_), .CO(add_104_carry_7_), 
        .S(N342) );
  ADDFX2 U262 ( .A(n38), .B(n41), .CI(add_104_carry_7_), .CO(add_104_carry_8_), 
        .S(N343) );
  ADDFX2 U263 ( .A(n39), .B(n42), .CI(add_104_carry_8_), .CO(add_104_carry_9_), 
        .S(N344) );
  ADDFX2 U264 ( .A(n40), .B(n43), .CI(add_104_carry_9_), .CO(add_104_carry_10_), .S(N345) );
  ADDFX2 U265 ( .A(n41), .B(n44), .CI(add_104_carry_10_), .CO(
        add_104_carry_11_), .S(N346) );
  ADDFX2 U266 ( .A(n42), .B(n45), .CI(add_104_carry_11_), .CO(
        add_104_carry_12_), .S(N347) );
  ADDFX2 U267 ( .A(n43), .B(n46), .CI(add_104_carry_12_), .CO(
        add_104_carry_13_), .S(N348) );
  ADDFX2 U268 ( .A(n44), .B(n47), .CI(add_104_carry_13_), .CO(
        add_104_carry_14_), .S(N349) );
  ADDFX2 U269 ( .A(n45), .B(n48), .CI(add_104_carry_14_), .CO(
        add_104_carry_15_), .S(N350) );
  ADDFX2 U270 ( .A(n46), .B(n49), .CI(add_104_carry_15_), .CO(
        add_104_carry_16_), .S(N351) );
  ADDFX2 U271 ( .A(n47), .B(x7[15]), .CI(add_104_carry_16_), .CO(
        add_104_carry_17_), .S(N352) );
  ADDFX2 U272 ( .A(n48), .B(x7[15]), .CI(add_104_carry_17_), .CO(
        add_104_carry_18_), .S(N353) );
  ADDFX2 U273 ( .A(n63), .B(n66), .CI(add_86_carry_6_), .CO(add_86_carry_7_), 
        .S(N172) );
  ADDFX2 U274 ( .A(n64), .B(n67), .CI(add_86_carry_7_), .CO(add_86_carry_8_), 
        .S(N173) );
  ADDFX2 U275 ( .A(n65), .B(n68), .CI(add_86_carry_8_), .CO(add_86_carry_9_), 
        .S(N174) );
  ADDFX2 U276 ( .A(n66), .B(n69), .CI(add_86_carry_9_), .CO(add_86_carry_10_), 
        .S(N175) );
  ADDFX2 U277 ( .A(n67), .B(n70), .CI(add_86_carry_10_), .CO(add_86_carry_11_), 
        .S(N176) );
  ADDFX2 U278 ( .A(n68), .B(n71), .CI(add_86_carry_11_), .CO(add_86_carry_12_), 
        .S(N177) );
  ADDFX2 U279 ( .A(n69), .B(n72), .CI(add_86_carry_12_), .CO(add_86_carry_13_), 
        .S(N178) );
  ADDFX2 U280 ( .A(n70), .B(n73), .CI(add_86_carry_13_), .CO(add_86_carry_14_), 
        .S(N179) );
  ADDFX2 U281 ( .A(n71), .B(n74), .CI(add_86_carry_14_), .CO(add_86_carry_15_), 
        .S(N180) );
  ADDFX2 U282 ( .A(n72), .B(n75), .CI(add_86_carry_15_), .CO(add_86_carry_16_), 
        .S(N181) );
  ADDFX2 U283 ( .A(n73), .B(x5[15]), .CI(add_86_carry_16_), .CO(
        add_86_carry_17_), .S(N182) );
  ADDFX2 U284 ( .A(n74), .B(x5[15]), .CI(add_86_carry_17_), .CO(
        add_86_carry_18_), .S(N183) );
  ADDFX2 U285 ( .A(n50), .B(n53), .CI(add_95_carry_6_), .CO(add_95_carry_7_), 
        .S(N257) );
  ADDFX2 U286 ( .A(n51), .B(n54), .CI(add_95_carry_7_), .CO(add_95_carry_8_), 
        .S(N258) );
  ADDFX2 U287 ( .A(n52), .B(n55), .CI(add_95_carry_8_), .CO(add_95_carry_9_), 
        .S(N259) );
  ADDFX2 U288 ( .A(n53), .B(n56), .CI(add_95_carry_9_), .CO(add_95_carry_10_), 
        .S(N260) );
  ADDFX2 U289 ( .A(n54), .B(n57), .CI(add_95_carry_10_), .CO(add_95_carry_11_), 
        .S(N261) );
  ADDFX2 U290 ( .A(n55), .B(n58), .CI(add_95_carry_11_), .CO(add_95_carry_12_), 
        .S(N262) );
  ADDFX2 U291 ( .A(n56), .B(n59), .CI(add_95_carry_12_), .CO(add_95_carry_13_), 
        .S(N263) );
  ADDFX2 U292 ( .A(n57), .B(n60), .CI(add_95_carry_13_), .CO(add_95_carry_14_), 
        .S(N264) );
  ADDFX2 U293 ( .A(n58), .B(n61), .CI(add_95_carry_14_), .CO(add_95_carry_15_), 
        .S(N265) );
  ADDFX2 U294 ( .A(n59), .B(n62), .CI(add_95_carry_15_), .CO(add_95_carry_16_), 
        .S(N266) );
  ADDFX2 U295 ( .A(n60), .B(x6[15]), .CI(add_95_carry_16_), .CO(
        add_95_carry_17_), .S(N267) );
  ADDFX2 U296 ( .A(n61), .B(x6[15]), .CI(add_95_carry_17_), .CO(
        add_95_carry_18_), .S(N268) );
  ADDFX2 U297 ( .A(n76), .B(n79), .CI(add_77_carry_6_), .CO(add_77_carry_7_), 
        .S(N87) );
  ADDFX2 U298 ( .A(n77), .B(n80), .CI(add_77_carry_7_), .CO(add_77_carry_8_), 
        .S(N88) );
  ADDFX2 U299 ( .A(n78), .B(n81), .CI(add_77_carry_8_), .CO(add_77_carry_9_), 
        .S(N89) );
  ADDFX2 U300 ( .A(n79), .B(n82), .CI(add_77_carry_9_), .CO(add_77_carry_10_), 
        .S(N90) );
  ADDFX2 U301 ( .A(n80), .B(n83), .CI(add_77_carry_10_), .CO(add_77_carry_11_), 
        .S(N91) );
  ADDFX2 U302 ( .A(n81), .B(n84), .CI(add_77_carry_11_), .CO(add_77_carry_12_), 
        .S(N92) );
  ADDFX2 U303 ( .A(n82), .B(n85), .CI(add_77_carry_12_), .CO(add_77_carry_13_), 
        .S(N93) );
  ADDFX2 U304 ( .A(n83), .B(n86), .CI(add_77_carry_13_), .CO(add_77_carry_14_), 
        .S(N94) );
  ADDFX2 U305 ( .A(n84), .B(n87), .CI(add_77_carry_14_), .CO(add_77_carry_15_), 
        .S(N95) );
  ADDFX2 U306 ( .A(n85), .B(n88), .CI(add_77_carry_15_), .CO(add_77_carry_16_), 
        .S(N96) );
  ADDFX2 U307 ( .A(n86), .B(x4[15]), .CI(add_77_carry_16_), .CO(
        add_77_carry_17_), .S(N97) );
  ADDFX2 U308 ( .A(n87), .B(x4[15]), .CI(add_77_carry_17_), .CO(
        add_77_carry_18_), .S(N98) );
  ADDFX2 U309 ( .A(n37), .B(n39), .CI(add_102_carry_5_), .CO(add_102_carry_6_), 
        .S(N321) );
  ADDFX2 U310 ( .A(n38), .B(n40), .CI(add_102_carry_6_), .CO(add_102_carry_7_), 
        .S(N322) );
  ADDFX2 U311 ( .A(n39), .B(n41), .CI(add_102_carry_7_), .CO(add_102_carry_8_), 
        .S(N323) );
  ADDFX2 U312 ( .A(n40), .B(n42), .CI(add_102_carry_8_), .CO(add_102_carry_9_), 
        .S(N324) );
  ADDFX2 U313 ( .A(n41), .B(n43), .CI(add_102_carry_9_), .CO(add_102_carry_10_), .S(N325) );
  ADDFX2 U314 ( .A(n42), .B(n44), .CI(add_102_carry_10_), .CO(
        add_102_carry_11_), .S(N326) );
  ADDFX2 U315 ( .A(n43), .B(n45), .CI(add_102_carry_11_), .CO(
        add_102_carry_12_), .S(N327) );
  ADDFX2 U316 ( .A(n44), .B(n46), .CI(add_102_carry_12_), .CO(
        add_102_carry_13_), .S(N328) );
  ADDFX2 U317 ( .A(n45), .B(n47), .CI(add_102_carry_13_), .CO(
        add_102_carry_14_), .S(N329) );
  ADDFX2 U318 ( .A(n46), .B(n48), .CI(add_102_carry_14_), .CO(
        add_102_carry_15_), .S(N330) );
  ADDFX2 U319 ( .A(n47), .B(n49), .CI(add_102_carry_15_), .CO(
        add_102_carry_16_), .S(N331) );
  ADDFX2 U320 ( .A(n48), .B(x7[15]), .CI(add_102_carry_16_), .CO(
        add_102_carry_17_), .S(N332) );
  ADDFX2 U321 ( .A(n50), .B(n52), .CI(add_93_carry_5_), .CO(add_93_carry_6_), 
        .S(N236) );
  ADDFX2 U322 ( .A(n51), .B(n53), .CI(add_93_carry_6_), .CO(add_93_carry_7_), 
        .S(N237) );
  ADDFX2 U323 ( .A(n52), .B(n54), .CI(add_93_carry_7_), .CO(add_93_carry_8_), 
        .S(N238) );
  ADDFX2 U324 ( .A(n53), .B(n55), .CI(add_93_carry_8_), .CO(add_93_carry_9_), 
        .S(N239) );
  ADDFX2 U325 ( .A(n54), .B(n56), .CI(add_93_carry_9_), .CO(add_93_carry_10_), 
        .S(N240) );
  ADDFX2 U326 ( .A(n55), .B(n57), .CI(add_93_carry_10_), .CO(add_93_carry_11_), 
        .S(N241) );
  ADDFX2 U327 ( .A(n56), .B(n58), .CI(add_93_carry_11_), .CO(add_93_carry_12_), 
        .S(N242) );
  ADDFX2 U328 ( .A(n57), .B(n59), .CI(add_93_carry_12_), .CO(add_93_carry_13_), 
        .S(N243) );
  ADDFX2 U329 ( .A(n58), .B(n60), .CI(add_93_carry_13_), .CO(add_93_carry_14_), 
        .S(N244) );
  ADDFX2 U330 ( .A(n59), .B(n61), .CI(add_93_carry_14_), .CO(add_93_carry_15_), 
        .S(N245) );
  ADDFX2 U331 ( .A(n60), .B(n62), .CI(add_93_carry_15_), .CO(add_93_carry_16_), 
        .S(N246) );
  ADDFX2 U332 ( .A(n61), .B(x6[15]), .CI(add_93_carry_16_), .CO(
        add_93_carry_17_), .S(N247) );
  ADDFX2 U333 ( .A(n63), .B(n65), .CI(add_84_carry_5_), .CO(add_84_carry_6_), 
        .S(N151) );
  ADDFX2 U334 ( .A(n64), .B(n66), .CI(add_84_carry_6_), .CO(add_84_carry_7_), 
        .S(N152) );
  ADDFX2 U335 ( .A(n65), .B(n67), .CI(add_84_carry_7_), .CO(add_84_carry_8_), 
        .S(N153) );
  ADDFX2 U336 ( .A(n66), .B(n68), .CI(add_84_carry_8_), .CO(add_84_carry_9_), 
        .S(N154) );
  ADDFX2 U337 ( .A(n67), .B(n69), .CI(add_84_carry_9_), .CO(add_84_carry_10_), 
        .S(N155) );
  ADDFX2 U338 ( .A(n68), .B(n70), .CI(add_84_carry_10_), .CO(add_84_carry_11_), 
        .S(N156) );
  ADDFX2 U339 ( .A(n69), .B(n71), .CI(add_84_carry_11_), .CO(add_84_carry_12_), 
        .S(N157) );
  ADDFX2 U340 ( .A(n70), .B(n72), .CI(add_84_carry_12_), .CO(add_84_carry_13_), 
        .S(N158) );
  ADDFX2 U341 ( .A(n71), .B(n73), .CI(add_84_carry_13_), .CO(add_84_carry_14_), 
        .S(N159) );
  ADDFX2 U342 ( .A(n72), .B(n74), .CI(add_84_carry_14_), .CO(add_84_carry_15_), 
        .S(N160) );
  ADDFX2 U343 ( .A(n73), .B(n75), .CI(add_84_carry_15_), .CO(add_84_carry_16_), 
        .S(N161) );
  ADDFX2 U344 ( .A(n74), .B(x5[15]), .CI(add_84_carry_16_), .CO(
        add_84_carry_17_), .S(N162) );
  ADDFX2 U345 ( .A(n76), .B(n78), .CI(add_75_carry_5_), .CO(add_75_carry_6_), 
        .S(N66) );
  ADDFX2 U346 ( .A(n77), .B(n79), .CI(add_75_carry_6_), .CO(add_75_carry_7_), 
        .S(N67) );
  ADDFX2 U347 ( .A(n78), .B(n80), .CI(add_75_carry_7_), .CO(add_75_carry_8_), 
        .S(N68) );
  ADDFX2 U348 ( .A(n79), .B(n81), .CI(add_75_carry_8_), .CO(add_75_carry_9_), 
        .S(N69) );
  ADDFX2 U349 ( .A(n80), .B(n82), .CI(add_75_carry_9_), .CO(add_75_carry_10_), 
        .S(N70) );
  ADDFX2 U350 ( .A(n81), .B(n83), .CI(add_75_carry_10_), .CO(add_75_carry_11_), 
        .S(N71) );
  ADDFX2 U351 ( .A(n82), .B(n84), .CI(add_75_carry_11_), .CO(add_75_carry_12_), 
        .S(N72) );
  ADDFX2 U352 ( .A(n83), .B(n85), .CI(add_75_carry_12_), .CO(add_75_carry_13_), 
        .S(N73) );
  ADDFX2 U353 ( .A(n84), .B(n86), .CI(add_75_carry_13_), .CO(add_75_carry_14_), 
        .S(N74) );
  ADDFX2 U354 ( .A(n85), .B(n87), .CI(add_75_carry_14_), .CO(add_75_carry_15_), 
        .S(N75) );
  ADDFX2 U355 ( .A(n86), .B(n88), .CI(add_75_carry_15_), .CO(add_75_carry_16_), 
        .S(N76) );
  ADDFX2 U356 ( .A(n87), .B(x4[15]), .CI(add_75_carry_16_), .CO(
        add_75_carry_17_), .S(N77) );
  ADDFX2 U357 ( .A(n37), .B(n38), .CI(add_100_carry_6_), .CO(add_100_carry_7_), 
        .S(N301) );
  ADDFX2 U358 ( .A(n38), .B(n39), .CI(add_100_carry_7_), .CO(add_100_carry_8_), 
        .S(N302) );
  ADDFX2 U359 ( .A(n39), .B(n40), .CI(add_100_carry_8_), .CO(add_100_carry_9_), 
        .S(N303) );
  ADDFX2 U360 ( .A(n40), .B(n41), .CI(add_100_carry_9_), .CO(add_100_carry_10_), .S(N304) );
  ADDFX2 U361 ( .A(n41), .B(n42), .CI(add_100_carry_10_), .CO(
        add_100_carry_11_), .S(N305) );
  ADDFX2 U362 ( .A(n42), .B(n43), .CI(add_100_carry_11_), .CO(
        add_100_carry_12_), .S(N306) );
  ADDFX2 U363 ( .A(n43), .B(n44), .CI(add_100_carry_12_), .CO(
        add_100_carry_13_), .S(N307) );
  ADDFX2 U364 ( .A(n44), .B(n45), .CI(add_100_carry_13_), .CO(
        add_100_carry_14_), .S(N308) );
  ADDFX2 U365 ( .A(n45), .B(n46), .CI(add_100_carry_14_), .CO(
        add_100_carry_15_), .S(N309) );
  ADDFX2 U366 ( .A(n46), .B(n47), .CI(add_100_carry_15_), .CO(
        add_100_carry_16_), .S(N310) );
  ADDFX2 U367 ( .A(n47), .B(n48), .CI(add_100_carry_16_), .CO(
        add_100_carry_17_), .S(N311) );
  ADDFX2 U368 ( .A(n48), .B(n49), .CI(add_100_carry_17_), .CO(
        add_100_carry_18_), .S(N312) );
  ADDFX2 U369 ( .A(n76), .B(n82), .CI(add_72_carry_8_), .CO(add_72_carry_9_), 
        .S(N25) );
  ADDFX2 U370 ( .A(n77), .B(n83), .CI(add_72_carry_9_), .CO(add_72_carry_10_), 
        .S(N26) );
  ADDFX2 U371 ( .A(n78), .B(n84), .CI(add_72_carry_10_), .CO(add_72_carry_11_), 
        .S(N27) );
  ADDFX2 U372 ( .A(n79), .B(n85), .CI(add_72_carry_11_), .CO(add_72_carry_12_), 
        .S(N28) );
  ADDFX2 U373 ( .A(n80), .B(n86), .CI(add_72_carry_12_), .CO(add_72_carry_13_), 
        .S(N29) );
  ADDFX2 U374 ( .A(n81), .B(n87), .CI(add_72_carry_13_), .CO(add_72_carry_14_), 
        .S(N30) );
  ADDFX2 U375 ( .A(n82), .B(n88), .CI(add_72_carry_14_), .CO(add_72_carry_15_), 
        .S(N31) );
  ADDFX2 U376 ( .A(n83), .B(x4[15]), .CI(add_72_carry_15_), .CO(
        add_72_carry_16_), .S(N32) );
  ADDFX2 U377 ( .A(n84), .B(x4[15]), .CI(add_72_carry_16_), .CO(
        add_72_carry_17_), .S(N33) );
  ADDFX2 U378 ( .A(n85), .B(x4[15]), .CI(add_72_carry_17_), .CO(
        add_72_carry_18_), .S(N34) );
  ADDFX2 U379 ( .A(n86), .B(x4[15]), .CI(add_72_carry_18_), .CO(
        add_72_carry_19_), .S(N35) );
  ADDFX2 U380 ( .A(n87), .B(x4[15]), .CI(add_72_carry_19_), .CO(
        add_72_carry_20_), .S(N36) );
  ADDFX2 U381 ( .A(n76), .B(n77), .CI(add_73_carry_6_), .CO(add_73_carry_7_), 
        .S(N46) );
  ADDFX2 U382 ( .A(n77), .B(n78), .CI(add_73_carry_7_), .CO(add_73_carry_8_), 
        .S(N47) );
  ADDFX2 U383 ( .A(n78), .B(n79), .CI(add_73_carry_8_), .CO(add_73_carry_9_), 
        .S(N48) );
  ADDFX2 U384 ( .A(n79), .B(n80), .CI(add_73_carry_9_), .CO(add_73_carry_10_), 
        .S(N49) );
  ADDFX2 U385 ( .A(n80), .B(n81), .CI(add_73_carry_10_), .CO(add_73_carry_11_), 
        .S(N50) );
  ADDFX2 U386 ( .A(n81), .B(n82), .CI(add_73_carry_11_), .CO(add_73_carry_12_), 
        .S(N51) );
  ADDFX2 U387 ( .A(n82), .B(n83), .CI(add_73_carry_12_), .CO(add_73_carry_13_), 
        .S(N52) );
  ADDFX2 U388 ( .A(n83), .B(n84), .CI(add_73_carry_13_), .CO(add_73_carry_14_), 
        .S(N53) );
  ADDFX2 U389 ( .A(n84), .B(n85), .CI(add_73_carry_14_), .CO(add_73_carry_15_), 
        .S(N54) );
  ADDFX2 U390 ( .A(n85), .B(n86), .CI(add_73_carry_15_), .CO(add_73_carry_16_), 
        .S(N55) );
  ADDFX2 U391 ( .A(n86), .B(n87), .CI(add_73_carry_16_), .CO(add_73_carry_17_), 
        .S(N56) );
  ADDFX2 U392 ( .A(n87), .B(n88), .CI(add_73_carry_17_), .CO(add_73_carry_18_), 
        .S(N57) );
  ADDFX2 U393 ( .A(n63), .B(n64), .CI(add_82_carry_6_), .CO(add_82_carry_7_), 
        .S(N131) );
  ADDFX2 U394 ( .A(n64), .B(n65), .CI(add_82_carry_7_), .CO(add_82_carry_8_), 
        .S(N132) );
  ADDFX2 U395 ( .A(n65), .B(n66), .CI(add_82_carry_8_), .CO(add_82_carry_9_), 
        .S(N133) );
  ADDFX2 U396 ( .A(n66), .B(n67), .CI(add_82_carry_9_), .CO(add_82_carry_10_), 
        .S(N134) );
  ADDFX2 U397 ( .A(n67), .B(n68), .CI(add_82_carry_10_), .CO(add_82_carry_11_), 
        .S(N135) );
  ADDFX2 U398 ( .A(n68), .B(n69), .CI(add_82_carry_11_), .CO(add_82_carry_12_), 
        .S(N136) );
  ADDFX2 U399 ( .A(n69), .B(n70), .CI(add_82_carry_12_), .CO(add_82_carry_13_), 
        .S(N137) );
  ADDFX2 U400 ( .A(n70), .B(n71), .CI(add_82_carry_13_), .CO(add_82_carry_14_), 
        .S(N138) );
  ADDFX2 U401 ( .A(n71), .B(n72), .CI(add_82_carry_14_), .CO(add_82_carry_15_), 
        .S(N139) );
  ADDFX2 U402 ( .A(n72), .B(n73), .CI(add_82_carry_15_), .CO(add_82_carry_16_), 
        .S(N140) );
  ADDFX2 U403 ( .A(n73), .B(n74), .CI(add_82_carry_16_), .CO(add_82_carry_17_), 
        .S(N141) );
  ADDFX2 U404 ( .A(n74), .B(n75), .CI(add_82_carry_17_), .CO(add_82_carry_18_), 
        .S(N142) );
  ADDFX2 U405 ( .A(n50), .B(n51), .CI(add_91_carry_6_), .CO(add_91_carry_7_), 
        .S(N216) );
  ADDFX2 U406 ( .A(n51), .B(n52), .CI(add_91_carry_7_), .CO(add_91_carry_8_), 
        .S(N217) );
  ADDFX2 U407 ( .A(n52), .B(n53), .CI(add_91_carry_8_), .CO(add_91_carry_9_), 
        .S(N218) );
  ADDFX2 U408 ( .A(n53), .B(n54), .CI(add_91_carry_9_), .CO(add_91_carry_10_), 
        .S(N219) );
  ADDFX2 U409 ( .A(n54), .B(n55), .CI(add_91_carry_10_), .CO(add_91_carry_11_), 
        .S(N220) );
  ADDFX2 U410 ( .A(n55), .B(n56), .CI(add_91_carry_11_), .CO(add_91_carry_12_), 
        .S(N221) );
  ADDFX2 U411 ( .A(n56), .B(n57), .CI(add_91_carry_12_), .CO(add_91_carry_13_), 
        .S(N222) );
  ADDFX2 U412 ( .A(n57), .B(n58), .CI(add_91_carry_13_), .CO(add_91_carry_14_), 
        .S(N223) );
  ADDFX2 U413 ( .A(n58), .B(n59), .CI(add_91_carry_14_), .CO(add_91_carry_15_), 
        .S(N224) );
  ADDFX2 U414 ( .A(n59), .B(n60), .CI(add_91_carry_15_), .CO(add_91_carry_16_), 
        .S(N225) );
  ADDFX2 U415 ( .A(n60), .B(n61), .CI(add_91_carry_16_), .CO(add_91_carry_17_), 
        .S(N226) );
  ADDFX2 U416 ( .A(n61), .B(n62), .CI(add_91_carry_17_), .CO(add_91_carry_18_), 
        .S(N227) );
  ADDFX2 U417 ( .A(n63), .B(n69), .CI(add_81_carry_8_), .CO(add_81_carry_9_), 
        .S(N110) );
  ADDFX2 U418 ( .A(n64), .B(n70), .CI(add_81_carry_9_), .CO(add_81_carry_10_), 
        .S(N111) );
  ADDFX2 U419 ( .A(n65), .B(n71), .CI(add_81_carry_10_), .CO(add_81_carry_11_), 
        .S(N112) );
  ADDFX2 U420 ( .A(n66), .B(n72), .CI(add_81_carry_11_), .CO(add_81_carry_12_), 
        .S(N113) );
  ADDFX2 U421 ( .A(n67), .B(n73), .CI(add_81_carry_12_), .CO(add_81_carry_13_), 
        .S(N114) );
  ADDFX2 U422 ( .A(n68), .B(n74), .CI(add_81_carry_13_), .CO(add_81_carry_14_), 
        .S(N115) );
  ADDFX2 U423 ( .A(n69), .B(n75), .CI(add_81_carry_14_), .CO(add_81_carry_15_), 
        .S(N116) );
  ADDFX2 U424 ( .A(n70), .B(x5[15]), .CI(add_81_carry_15_), .CO(
        add_81_carry_16_), .S(N117) );
  ADDFX2 U425 ( .A(n71), .B(x5[15]), .CI(add_81_carry_16_), .CO(
        add_81_carry_17_), .S(N118) );
  ADDFX2 U426 ( .A(n72), .B(x5[15]), .CI(add_81_carry_17_), .CO(
        add_81_carry_18_), .S(N119) );
  ADDFX2 U427 ( .A(n73), .B(x5[15]), .CI(add_81_carry_18_), .CO(
        add_81_carry_19_), .S(N120) );
  ADDFX2 U428 ( .A(n74), .B(x5[15]), .CI(add_81_carry_19_), .CO(
        add_81_carry_20_), .S(N121) );
  ADDFX2 U429 ( .A(n50), .B(n56), .CI(add_90_carry_8_), .CO(add_90_carry_9_), 
        .S(N195) );
  ADDFX2 U430 ( .A(n51), .B(n57), .CI(add_90_carry_9_), .CO(add_90_carry_10_), 
        .S(N196) );
  ADDFX2 U431 ( .A(n52), .B(n58), .CI(add_90_carry_10_), .CO(add_90_carry_11_), 
        .S(N197) );
  ADDFX2 U432 ( .A(n53), .B(n59), .CI(add_90_carry_11_), .CO(add_90_carry_12_), 
        .S(N198) );
  ADDFX2 U433 ( .A(n54), .B(n60), .CI(add_90_carry_12_), .CO(add_90_carry_13_), 
        .S(N199) );
  ADDFX2 U434 ( .A(n55), .B(n61), .CI(add_90_carry_13_), .CO(add_90_carry_14_), 
        .S(N200) );
  ADDFX2 U435 ( .A(n56), .B(n62), .CI(add_90_carry_14_), .CO(add_90_carry_15_), 
        .S(N201) );
  ADDFX2 U436 ( .A(n57), .B(x6[15]), .CI(add_90_carry_15_), .CO(
        add_90_carry_16_), .S(N202) );
  ADDFX2 U437 ( .A(n58), .B(x6[15]), .CI(add_90_carry_16_), .CO(
        add_90_carry_17_), .S(N203) );
  ADDFX2 U438 ( .A(n59), .B(x6[15]), .CI(add_90_carry_17_), .CO(
        add_90_carry_18_), .S(N204) );
  ADDFX2 U439 ( .A(n60), .B(x6[15]), .CI(add_90_carry_18_), .CO(
        add_90_carry_19_), .S(N205) );
  ADDFX2 U440 ( .A(n61), .B(x6[15]), .CI(add_90_carry_19_), .CO(
        add_90_carry_20_), .S(N206) );
  ADDFX2 U441 ( .A(n37), .B(n43), .CI(add_99_carry_8_), .CO(add_99_carry_9_), 
        .S(N280) );
  ADDFX2 U442 ( .A(n38), .B(n44), .CI(add_99_carry_9_), .CO(add_99_carry_10_), 
        .S(N281) );
  ADDFX2 U443 ( .A(n39), .B(n45), .CI(add_99_carry_10_), .CO(add_99_carry_11_), 
        .S(N282) );
  ADDFX2 U444 ( .A(n40), .B(n46), .CI(add_99_carry_11_), .CO(add_99_carry_12_), 
        .S(N283) );
  ADDFX2 U445 ( .A(n41), .B(n47), .CI(add_99_carry_12_), .CO(add_99_carry_13_), 
        .S(N284) );
  ADDFX2 U446 ( .A(n42), .B(n48), .CI(add_99_carry_13_), .CO(add_99_carry_14_), 
        .S(N285) );
  ADDFX2 U447 ( .A(n43), .B(n49), .CI(add_99_carry_14_), .CO(add_99_carry_15_), 
        .S(N286) );
  ADDFX2 U448 ( .A(n44), .B(x7[15]), .CI(add_99_carry_15_), .CO(
        add_99_carry_16_), .S(N287) );
  ADDFX2 U449 ( .A(n45), .B(x7[15]), .CI(add_99_carry_16_), .CO(
        add_99_carry_17_), .S(N288) );
  ADDFX2 U450 ( .A(n46), .B(x7[15]), .CI(add_99_carry_17_), .CO(
        add_99_carry_18_), .S(N289) );
  ADDFX2 U451 ( .A(n47), .B(x7[15]), .CI(add_99_carry_18_), .CO(
        add_99_carry_19_), .S(N290) );
  ADDFX2 U452 ( .A(n48), .B(x7[15]), .CI(add_99_carry_19_), .CO(
        add_99_carry_20_), .S(N291) );
  INVX1 U453 ( .A(n414), .Y(n221) );
  INVX1 U454 ( .A(n222), .Y(n181) );
  INVX1 U455 ( .A(n414), .Y(n222) );
  INVX1 U456 ( .A(n414), .Y(n220) );
  INVX1 U457 ( .A(n414), .Y(n219) );
  INVX1 U458 ( .A(n414), .Y(n218) );
  INVX1 U459 ( .A(n414), .Y(n217) );
  INVX1 U460 ( .A(n414), .Y(n216) );
  INVX1 U461 ( .A(n414), .Y(n215) );
  INVX1 U462 ( .A(n414), .Y(n214) );
  INVX1 U463 ( .A(n414), .Y(n213) );
  INVX1 U464 ( .A(n414), .Y(n212) );
  INVX1 U465 ( .A(n582), .Y(y0[16]) );
  INVX1 U466 ( .A(n581), .Y(y0[17]) );
  INVX1 U467 ( .A(n580), .Y(y0[18]) );
  INVX1 U468 ( .A(n579), .Y(y0[19]) );
  INVX1 U469 ( .A(n577), .Y(y0[20]) );
  INVX1 U470 ( .A(n576), .Y(y0[21]) );
  INVX1 U471 ( .A(n560), .Y(y1[16]) );
  INVX1 U472 ( .A(n559), .Y(y1[17]) );
  INVX1 U473 ( .A(n558), .Y(y1[18]) );
  INVX1 U474 ( .A(n557), .Y(y1[19]) );
  INVX1 U475 ( .A(n555), .Y(y1[20]) );
  INVX1 U476 ( .A(n554), .Y(y1[21]) );
  INVX1 U477 ( .A(n538), .Y(y2[16]) );
  INVX1 U478 ( .A(n537), .Y(y2[17]) );
  INVX1 U479 ( .A(n536), .Y(y2[18]) );
  INVX1 U480 ( .A(n535), .Y(y2[19]) );
  INVX1 U481 ( .A(n533), .Y(y2[20]) );
  INVX1 U482 ( .A(n532), .Y(y2[21]) );
  INVX1 U483 ( .A(n516), .Y(y3[16]) );
  INVX1 U484 ( .A(n515), .Y(y3[17]) );
  INVX1 U485 ( .A(n514), .Y(y3[18]) );
  INVX1 U486 ( .A(n513), .Y(y3[19]) );
  INVX1 U487 ( .A(n511), .Y(y3[20]) );
  INVX1 U488 ( .A(n510), .Y(y3[21]) );
  INVX1 U489 ( .A(n494), .Y(y4[16]) );
  INVX1 U490 ( .A(n493), .Y(y4[17]) );
  INVX1 U491 ( .A(n492), .Y(y4[18]) );
  INVX1 U492 ( .A(n491), .Y(y4[19]) );
  INVX1 U493 ( .A(n489), .Y(y4[20]) );
  INVX1 U494 ( .A(n488), .Y(y4[21]) );
  INVX1 U495 ( .A(n472), .Y(y5[16]) );
  INVX1 U496 ( .A(n471), .Y(y5[17]) );
  INVX1 U497 ( .A(n470), .Y(y5[18]) );
  INVX1 U498 ( .A(n469), .Y(y5[19]) );
  INVX1 U499 ( .A(n467), .Y(y5[20]) );
  INVX1 U500 ( .A(n466), .Y(y5[21]) );
  INVX1 U501 ( .A(n450), .Y(y6[16]) );
  INVX1 U502 ( .A(n449), .Y(y6[17]) );
  INVX1 U503 ( .A(n448), .Y(y6[18]) );
  INVX1 U504 ( .A(n447), .Y(y6[19]) );
  INVX1 U505 ( .A(n445), .Y(y6[20]) );
  INVX1 U506 ( .A(n444), .Y(y6[21]) );
  INVX1 U507 ( .A(n428), .Y(y7[16]) );
  INVX1 U508 ( .A(n427), .Y(y7[17]) );
  INVX1 U509 ( .A(n426), .Y(y7[18]) );
  INVX1 U510 ( .A(n425), .Y(y7[19]) );
  INVX1 U511 ( .A(n423), .Y(y7[20]) );
  INVX1 U512 ( .A(n422), .Y(y7[21]) );
  INVX1 U513 ( .A(x5_tmp[2]), .Y(n363) );
  INVX1 U514 ( .A(x5_tmp[3]), .Y(n362) );
  INVX1 U515 ( .A(x5_tmp[4]), .Y(n361) );
  INVX1 U516 ( .A(x5_tmp[5]), .Y(n360) );
  INVX1 U517 ( .A(x5_tmp[6]), .Y(n359) );
  INVX1 U518 ( .A(x5_tmp[7]), .Y(n358) );
  INVX1 U519 ( .A(x5_tmp[8]), .Y(n357) );
  INVX1 U520 ( .A(x5_tmp[9]), .Y(n356) );
  INVX1 U521 ( .A(x5_tmp[10]), .Y(n355) );
  INVX1 U522 ( .A(x5_tmp[11]), .Y(n354) );
  INVX1 U523 ( .A(x5_tmp[12]), .Y(n353) );
  INVX1 U524 ( .A(x5_tmp[13]), .Y(n352) );
  INVX1 U525 ( .A(x5_tmp[14]), .Y(n351) );
  INVX1 U526 ( .A(x5_tmp[15]), .Y(n350) );
  INVX1 U527 ( .A(x5_tmp[16]), .Y(n349) );
  INVX1 U528 ( .A(x5_tmp[17]), .Y(n348) );
  INVX1 U529 ( .A(x5_tmp[18]), .Y(n347) );
  INVX1 U530 ( .A(x5_tmp[19]), .Y(n346) );
  INVX1 U531 ( .A(x5_tmp[20]), .Y(n345) );
  INVX1 U532 ( .A(x5_tmp[21]), .Y(n344) );
  INVX1 U533 ( .A(x5_tmp[22]), .Y(n343) );
  INVX1 U534 ( .A(x5_tmp[23]), .Y(n342) );
  INVX1 U535 ( .A(x4_tmp[2]), .Y(n393) );
  INVX1 U536 ( .A(x4_tmp[3]), .Y(n394) );
  INVX1 U537 ( .A(x4_tmp[4]), .Y(n395) );
  INVX1 U538 ( .A(x4_tmp[5]), .Y(n396) );
  INVX1 U539 ( .A(x4_tmp[6]), .Y(n397) );
  INVX1 U540 ( .A(x4_tmp[7]), .Y(n398) );
  INVX1 U541 ( .A(x4_tmp[8]), .Y(n399) );
  INVX1 U542 ( .A(x4_tmp[9]), .Y(n400) );
  INVX1 U543 ( .A(x4_tmp[10]), .Y(n401) );
  INVX1 U544 ( .A(x4_tmp[11]), .Y(n402) );
  INVX1 U545 ( .A(x4_tmp[12]), .Y(n403) );
  INVX1 U546 ( .A(x4_tmp[13]), .Y(n404) );
  INVX1 U547 ( .A(x4_tmp[14]), .Y(n405) );
  INVX1 U548 ( .A(x4_tmp[15]), .Y(n406) );
  INVX1 U549 ( .A(x4_tmp[16]), .Y(n407) );
  INVX1 U550 ( .A(x4_tmp[17]), .Y(n408) );
  INVX1 U551 ( .A(x4_tmp[18]), .Y(n409) );
  INVX1 U552 ( .A(x4_tmp[19]), .Y(n410) );
  INVX1 U553 ( .A(x4_tmp[20]), .Y(n411) );
  INVX1 U554 ( .A(x4_tmp[21]), .Y(n412) );
  INVX1 U555 ( .A(x4_tmp[22]), .Y(n590) );
  INVX1 U556 ( .A(x4_tmp[23]), .Y(n591) );
  INVX1 U557 ( .A(x7_tmp[2]), .Y(n318) );
  INVX1 U558 ( .A(x7_tmp[3]), .Y(n319) );
  INVX1 U559 ( .A(x7_tmp[4]), .Y(n320) );
  INVX1 U560 ( .A(x7_tmp[5]), .Y(n321) );
  INVX1 U561 ( .A(x7_tmp[6]), .Y(n322) );
  INVX1 U562 ( .A(x7_tmp[7]), .Y(n323) );
  INVX1 U563 ( .A(x7_tmp[8]), .Y(n324) );
  INVX1 U564 ( .A(x7_tmp[9]), .Y(n325) );
  INVX1 U565 ( .A(x7_tmp[10]), .Y(n326) );
  INVX1 U566 ( .A(x7_tmp[11]), .Y(n327) );
  INVX1 U567 ( .A(x7_tmp[12]), .Y(n328) );
  INVX1 U568 ( .A(x7_tmp[13]), .Y(n329) );
  INVX1 U569 ( .A(x7_tmp[14]), .Y(n330) );
  INVX1 U570 ( .A(x7_tmp[15]), .Y(n331) );
  INVX1 U571 ( .A(x7_tmp[16]), .Y(n332) );
  INVX1 U572 ( .A(x7_tmp[17]), .Y(n333) );
  INVX1 U573 ( .A(x7_tmp[18]), .Y(n334) );
  INVX1 U574 ( .A(x7_tmp[19]), .Y(n335) );
  INVX1 U575 ( .A(x7_tmp[20]), .Y(n336) );
  INVX1 U576 ( .A(x7_tmp[21]), .Y(n337) );
  INVX1 U577 ( .A(x7_tmp[22]), .Y(n338) );
  INVX1 U578 ( .A(x7_tmp[23]), .Y(n339) );
  INVX1 U579 ( .A(x6_tmp[2]), .Y(n388) );
  INVX1 U580 ( .A(x6_tmp[3]), .Y(n387) );
  INVX1 U581 ( .A(x6_tmp[4]), .Y(n386) );
  INVX1 U582 ( .A(x6_tmp[5]), .Y(n385) );
  INVX1 U583 ( .A(x6_tmp[6]), .Y(n384) );
  INVX1 U584 ( .A(x6_tmp[7]), .Y(n383) );
  INVX1 U585 ( .A(x6_tmp[8]), .Y(n382) );
  INVX1 U586 ( .A(x6_tmp[9]), .Y(n381) );
  INVX1 U587 ( .A(x6_tmp[10]), .Y(n380) );
  INVX1 U588 ( .A(x6_tmp[11]), .Y(n379) );
  INVX1 U589 ( .A(x6_tmp[12]), .Y(n378) );
  INVX1 U590 ( .A(x6_tmp[13]), .Y(n377) );
  INVX1 U591 ( .A(x6_tmp[14]), .Y(n376) );
  INVX1 U592 ( .A(x6_tmp[15]), .Y(n375) );
  INVX1 U593 ( .A(x6_tmp[16]), .Y(n374) );
  INVX1 U594 ( .A(x6_tmp[17]), .Y(n373) );
  INVX1 U595 ( .A(x6_tmp[18]), .Y(n372) );
  INVX1 U596 ( .A(x6_tmp[19]), .Y(n371) );
  INVX1 U597 ( .A(x6_tmp[20]), .Y(n370) );
  INVX1 U598 ( .A(x6_tmp[21]), .Y(n369) );
  INVX1 U599 ( .A(x6_tmp[22]), .Y(n368) );
  INVX1 U600 ( .A(x6_tmp[23]), .Y(n367) );
  INVX1 U601 ( .A(x5_tmp[1]), .Y(n364) );
  INVX1 U602 ( .A(x4_tmp[1]), .Y(n392) );
  INVX1 U603 ( .A(x7_tmp[1]), .Y(n317) );
  INVX1 U604 ( .A(x6_tmp[1]), .Y(n389) );
  INVX1 U605 ( .A(x5_tmp[0]), .Y(n365) );
  INVX1 U606 ( .A(x4_tmp[0]), .Y(n391) );
  INVX1 U607 ( .A(x7_tmp[0]), .Y(n316) );
  INVX1 U608 ( .A(x6_tmp[0]), .Y(n390) );
  INVX1 U609 ( .A(x7_89[0]), .Y(n293) );
  INVX1 U610 ( .A(x5_89[0]), .Y(n270) );
  INVX1 U611 ( .A(x7_50[0]), .Y(n247) );
  INVX1 U612 ( .A(x5_50[0]), .Y(n315) );
  INVX1 U613 ( .A(x7_89[2]), .Y(n291) );
  INVX1 U614 ( .A(x7_89[3]), .Y(n290) );
  INVX1 U615 ( .A(x7_89[4]), .Y(n289) );
  INVX1 U616 ( .A(x7_89[5]), .Y(n288) );
  INVX1 U617 ( .A(x7_89[6]), .Y(n287) );
  INVX1 U618 ( .A(x7_89[7]), .Y(n286) );
  INVX1 U619 ( .A(x7_89[8]), .Y(n285) );
  INVX1 U620 ( .A(x7_89[9]), .Y(n284) );
  INVX1 U621 ( .A(x7_89[10]), .Y(n283) );
  INVX1 U622 ( .A(x7_89[11]), .Y(n282) );
  INVX1 U623 ( .A(x7_89[12]), .Y(n281) );
  INVX1 U624 ( .A(x7_89[13]), .Y(n280) );
  INVX1 U625 ( .A(x7_89[14]), .Y(n279) );
  INVX1 U626 ( .A(x7_89[15]), .Y(n278) );
  INVX1 U627 ( .A(x7_89[16]), .Y(n277) );
  INVX1 U628 ( .A(x7_89[17]), .Y(n276) );
  INVX1 U629 ( .A(x7_89[18]), .Y(n275) );
  INVX1 U630 ( .A(x7_89[19]), .Y(n274) );
  INVX1 U631 ( .A(x7_89[20]), .Y(n273) );
  INVX1 U632 ( .A(x7_89[21]), .Y(n272) );
  INVX1 U633 ( .A(x5_89[2]), .Y(n268) );
  INVX1 U634 ( .A(x5_89[3]), .Y(n267) );
  INVX1 U635 ( .A(x5_89[4]), .Y(n266) );
  INVX1 U636 ( .A(x5_89[5]), .Y(n265) );
  INVX1 U637 ( .A(x5_89[6]), .Y(n264) );
  INVX1 U638 ( .A(x5_89[7]), .Y(n263) );
  INVX1 U639 ( .A(x5_89[8]), .Y(n262) );
  INVX1 U640 ( .A(x5_89[9]), .Y(n261) );
  INVX1 U641 ( .A(x5_89[10]), .Y(n260) );
  INVX1 U642 ( .A(x5_89[11]), .Y(n259) );
  INVX1 U643 ( .A(x5_89[12]), .Y(n258) );
  INVX1 U644 ( .A(x5_89[13]), .Y(n257) );
  INVX1 U645 ( .A(x5_89[14]), .Y(n256) );
  INVX1 U646 ( .A(x5_89[15]), .Y(n255) );
  INVX1 U647 ( .A(x5_89[16]), .Y(n254) );
  INVX1 U648 ( .A(x5_89[17]), .Y(n253) );
  INVX1 U649 ( .A(x5_89[18]), .Y(n252) );
  INVX1 U650 ( .A(x5_89[19]), .Y(n251) );
  INVX1 U651 ( .A(x5_89[20]), .Y(n250) );
  INVX1 U652 ( .A(x5_89[21]), .Y(n249) );
  INVX1 U653 ( .A(x7_50[2]), .Y(n245) );
  INVX1 U654 ( .A(x7_50[3]), .Y(n244) );
  INVX1 U655 ( .A(x7_50[4]), .Y(n243) );
  INVX1 U656 ( .A(x7_50[5]), .Y(n242) );
  INVX1 U657 ( .A(x7_50[6]), .Y(n241) );
  INVX1 U658 ( .A(x7_50[7]), .Y(n240) );
  INVX1 U659 ( .A(x7_50[8]), .Y(n239) );
  INVX1 U660 ( .A(x7_50[9]), .Y(n238) );
  INVX1 U661 ( .A(x7_50[10]), .Y(n237) );
  INVX1 U662 ( .A(x7_50[11]), .Y(n236) );
  INVX1 U663 ( .A(x7_50[12]), .Y(n235) );
  INVX1 U664 ( .A(x7_50[13]), .Y(n234) );
  INVX1 U665 ( .A(x7_50[14]), .Y(n233) );
  INVX1 U666 ( .A(x7_50[15]), .Y(n232) );
  INVX1 U667 ( .A(x7_50[16]), .Y(n231) );
  INVX1 U668 ( .A(x7_50[17]), .Y(n230) );
  INVX1 U669 ( .A(x7_50[18]), .Y(n229) );
  INVX1 U670 ( .A(x7_50[19]), .Y(n228) );
  INVX1 U671 ( .A(x7_50[20]), .Y(n227) );
  INVX1 U672 ( .A(x5_50[2]), .Y(n313) );
  INVX1 U673 ( .A(x5_50[3]), .Y(n312) );
  INVX1 U674 ( .A(x5_50[4]), .Y(n311) );
  INVX1 U675 ( .A(x5_50[5]), .Y(n310) );
  INVX1 U676 ( .A(x5_50[6]), .Y(n309) );
  INVX1 U677 ( .A(x5_50[7]), .Y(n308) );
  INVX1 U678 ( .A(x5_50[8]), .Y(n307) );
  INVX1 U679 ( .A(x5_50[9]), .Y(n306) );
  INVX1 U680 ( .A(x5_50[10]), .Y(n305) );
  INVX1 U681 ( .A(x5_50[11]), .Y(n304) );
  INVX1 U682 ( .A(x5_50[12]), .Y(n303) );
  INVX1 U683 ( .A(x5_50[13]), .Y(n302) );
  INVX1 U684 ( .A(x5_50[14]), .Y(n301) );
  INVX1 U685 ( .A(x5_50[15]), .Y(n300) );
  INVX1 U686 ( .A(x5_50[16]), .Y(n299) );
  INVX1 U687 ( .A(x5_50[17]), .Y(n298) );
  INVX1 U688 ( .A(x5_50[18]), .Y(n297) );
  INVX1 U689 ( .A(x5_50[19]), .Y(n296) );
  INVX1 U690 ( .A(x5_50[20]), .Y(n295) );
  INVX1 U691 ( .A(x7_50[1]), .Y(n246) );
  INVX1 U692 ( .A(x5_50[1]), .Y(n314) );
  INVX1 U693 ( .A(x7_89[1]), .Y(n292) );
  INVX1 U694 ( .A(x5_89[1]), .Y(n269) );
  INVX1 U695 ( .A(n585), .Y(y0[13]) );
  AOI22X1 U696 ( .A0(N1640), .A1(n174), .B0(y0_tmp[13]), .B1(n97), .Y(n585) );
  INVX1 U697 ( .A(n584), .Y(y0[14]) );
  AOI22X1 U698 ( .A0(N1641), .A1(n174), .B0(y0_tmp[14]), .B1(n97), .Y(n584) );
  INVX1 U699 ( .A(n563), .Y(y1[13]) );
  AOI22X1 U700 ( .A0(N1662), .A1(n164), .B0(y1_tmp[13]), .B1(n99), .Y(n563) );
  INVX1 U701 ( .A(n562), .Y(y1[14]) );
  AOI22X1 U702 ( .A0(N1663), .A1(n164), .B0(y1_tmp[14]), .B1(n99), .Y(n562) );
  INVX1 U703 ( .A(n541), .Y(y2[13]) );
  AOI22X1 U704 ( .A0(N1684), .A1(n155), .B0(y2_tmp[13]), .B1(n101), .Y(n541)
         );
  INVX1 U705 ( .A(n540), .Y(y2[14]) );
  AOI22X1 U706 ( .A0(N1685), .A1(n155), .B0(y2_tmp[14]), .B1(n101), .Y(n540)
         );
  INVX1 U707 ( .A(n519), .Y(y3[13]) );
  AOI22X1 U708 ( .A0(N1706), .A1(n146), .B0(y3_tmp[13]), .B1(n103), .Y(n519)
         );
  INVX1 U709 ( .A(n518), .Y(y3[14]) );
  AOI22X1 U710 ( .A0(N1707), .A1(n146), .B0(y3_tmp[14]), .B1(n102), .Y(n518)
         );
  INVX1 U711 ( .A(n583), .Y(y0[15]) );
  AOI22X1 U712 ( .A0(N1642), .A1(n173), .B0(y0_tmp[15]), .B1(n97), .Y(n583) );
  INVX1 U713 ( .A(n561), .Y(y1[15]) );
  AOI22X1 U714 ( .A0(N1664), .A1(n163), .B0(y1_tmp[15]), .B1(n99), .Y(n561) );
  INVX1 U715 ( .A(n539), .Y(y2[15]) );
  AOI22X1 U716 ( .A0(N1686), .A1(n154), .B0(y2_tmp[15]), .B1(n101), .Y(n539)
         );
  INVX1 U717 ( .A(n517), .Y(y3[15]) );
  AOI22X1 U718 ( .A0(N1708), .A1(n145), .B0(y3_tmp[15]), .B1(n102), .Y(n517)
         );
  AOI22X1 U719 ( .A0(N1728), .A1(n137), .B0(y4_tmp[13]), .B1(n95), .Y(n497) );
  AOI22X1 U720 ( .A0(N1729), .A1(n137), .B0(y4_tmp[14]), .B1(n95), .Y(n496) );
  AOI22X1 U721 ( .A0(N1730), .A1(n136), .B0(y4_tmp[15]), .B1(n95), .Y(n495) );
  AOI22X1 U722 ( .A0(N1750), .A1(n128), .B0(y5_tmp[13]), .B1(n94), .Y(n475) );
  AOI22X1 U723 ( .A0(N1751), .A1(n128), .B0(y5_tmp[14]), .B1(n94), .Y(n474) );
  AOI22X1 U724 ( .A0(N1752), .A1(n127), .B0(y5_tmp[15]), .B1(n93), .Y(n473) );
  AOI22X1 U725 ( .A0(N1772), .A1(n119), .B0(y6_tmp[13]), .B1(n92), .Y(n453) );
  AOI22X1 U726 ( .A0(N1773), .A1(n119), .B0(y6_tmp[14]), .B1(n92), .Y(n452) );
  AOI22X1 U727 ( .A0(N1774), .A1(n118), .B0(y6_tmp[15]), .B1(n92), .Y(n451) );
  AOI22X1 U728 ( .A0(N1794), .A1(n110), .B0(y7_tmp[13]), .B1(n90), .Y(n431) );
  AOI22X1 U729 ( .A0(N1795), .A1(n110), .B0(y7_tmp[14]), .B1(n90), .Y(n430) );
  AOI22X1 U730 ( .A0(N1796), .A1(n109), .B0(y7_tmp[15]), .B1(n90), .Y(n429) );
  INVX1 U731 ( .A(n569), .Y(y0[8]) );
  AOI22X1 U732 ( .A0(N1635), .A1(n167), .B0(y0_tmp[8]), .B1(n98), .Y(n569) );
  INVX1 U733 ( .A(n568), .Y(y0[9]) );
  AOI22X1 U734 ( .A0(N1636), .A1(n167), .B0(y0_tmp[9]), .B1(n98), .Y(n568) );
  INVX1 U735 ( .A(n588), .Y(y0[10]) );
  AOI22X1 U736 ( .A0(N1637), .A1(n176), .B0(y0_tmp[10]), .B1(n100), .Y(n588)
         );
  INVX1 U737 ( .A(n587), .Y(y0[11]) );
  AOI22X1 U738 ( .A0(N1638), .A1(n175), .B0(y0_tmp[11]), .B1(n97), .Y(n587) );
  INVX1 U739 ( .A(n547), .Y(y1[8]) );
  AOI22X1 U740 ( .A0(N1657), .A1(n158), .B0(y1_tmp[8]), .B1(n100), .Y(n547) );
  INVX1 U741 ( .A(n546), .Y(y1[9]) );
  AOI22X1 U742 ( .A0(N1658), .A1(n158), .B0(y1_tmp[9]), .B1(n100), .Y(n546) );
  INVX1 U743 ( .A(n566), .Y(y1[10]) );
  AOI22X1 U744 ( .A0(N1659), .A1(n166), .B0(y1_tmp[10]), .B1(n98), .Y(n566) );
  INVX1 U745 ( .A(n565), .Y(y1[11]) );
  AOI22X1 U746 ( .A0(N1660), .A1(n165), .B0(y1_tmp[11]), .B1(n98), .Y(n565) );
  INVX1 U747 ( .A(n525), .Y(y2[8]) );
  AOI22X1 U748 ( .A0(N1679), .A1(n149), .B0(y2_tmp[8]), .B1(n103), .Y(n525) );
  INVX1 U749 ( .A(n524), .Y(y2[9]) );
  AOI22X1 U750 ( .A0(N1680), .A1(n149), .B0(y2_tmp[9]), .B1(n102), .Y(n524) );
  INVX1 U751 ( .A(n544), .Y(y2[10]) );
  AOI22X1 U752 ( .A0(N1681), .A1(n157), .B0(y2_tmp[10]), .B1(n100), .Y(n544)
         );
  INVX1 U753 ( .A(n543), .Y(y2[11]) );
  AOI22X1 U754 ( .A0(N1682), .A1(n156), .B0(y2_tmp[11]), .B1(n100), .Y(n543)
         );
  INVX1 U755 ( .A(n522), .Y(y3[10]) );
  AOI22X1 U756 ( .A0(N1703), .A1(n148), .B0(y3_tmp[10]), .B1(n102), .Y(n522)
         );
  INVX1 U757 ( .A(n521), .Y(y3[11]) );
  AOI22X1 U758 ( .A0(N1704), .A1(n147), .B0(y3_tmp[11]), .B1(n103), .Y(n521)
         );
  INVX1 U759 ( .A(n431), .Y(y7[13]) );
  INVX1 U760 ( .A(n503), .Y(y3[8]) );
  AOI22X1 U761 ( .A0(N1701), .A1(n140), .B0(y3_tmp[8]), .B1(n96), .Y(n503) );
  INVX1 U762 ( .A(n502), .Y(y3[9]) );
  AOI22X1 U763 ( .A0(N1702), .A1(n140), .B0(y3_tmp[9]), .B1(n96), .Y(n502) );
  INVX1 U764 ( .A(n496), .Y(y4[14]) );
  INVX1 U765 ( .A(n495), .Y(y4[15]) );
  INVX1 U766 ( .A(n474), .Y(y5[14]) );
  INVX1 U767 ( .A(n473), .Y(y5[15]) );
  INVX1 U768 ( .A(n452), .Y(y6[14]) );
  INVX1 U769 ( .A(n451), .Y(y6[15]) );
  ADDFX2 U770 ( .A(x4[1]), .B(n81), .CI(add_72_carry_7_), .CO(add_72_carry_8_), 
        .S(N24) );
  ADDFX2 U771 ( .A(x5[1]), .B(n68), .CI(add_81_carry_7_), .CO(add_81_carry_8_), 
        .S(N109) );
  ADDFX2 U772 ( .A(x6[1]), .B(n55), .CI(add_90_carry_7_), .CO(add_90_carry_8_), 
        .S(N194) );
  BUFX3 U773 ( .A(x5[7]), .Y(n68) );
  BUFX3 U774 ( .A(x5[8]), .Y(n69) );
  BUFX3 U775 ( .A(x6[7]), .Y(n55) );
  BUFX3 U776 ( .A(x6[8]), .Y(n56) );
  BUFX3 U777 ( .A(x4[7]), .Y(n81) );
  BUFX3 U778 ( .A(x4[8]), .Y(n82) );
  BUFX3 U779 ( .A(x7[7]), .Y(n42) );
  BUFX3 U780 ( .A(x7[8]), .Y(n43) );
  BUFX3 U781 ( .A(x4[4]), .Y(n78) );
  BUFX3 U782 ( .A(x4[5]), .Y(n79) );
  BUFX3 U783 ( .A(x5[4]), .Y(n65) );
  BUFX3 U784 ( .A(x5[5]), .Y(n66) );
  BUFX3 U785 ( .A(x6[4]), .Y(n52) );
  BUFX3 U786 ( .A(x6[5]), .Y(n53) );
  BUFX3 U787 ( .A(x5[6]), .Y(n67) );
  BUFX3 U788 ( .A(x6[6]), .Y(n54) );
  BUFX3 U789 ( .A(x4[6]), .Y(n80) );
  BUFX3 U790 ( .A(x7[4]), .Y(n39) );
  BUFX3 U791 ( .A(x7[5]), .Y(n40) );
  BUFX3 U792 ( .A(x7[6]), .Y(n41) );
  INVX1 U793 ( .A(n430), .Y(y7[14]) );
  INVX1 U794 ( .A(n429), .Y(y7[15]) );
  INVX1 U795 ( .A(n586), .Y(y0[12]) );
  AOI22X1 U796 ( .A0(N1639), .A1(n175), .B0(y0_tmp[12]), .B1(n97), .Y(n586) );
  INVX1 U797 ( .A(n564), .Y(y1[12]) );
  AOI22X1 U798 ( .A0(N1661), .A1(n165), .B0(y1_tmp[12]), .B1(n99), .Y(n564) );
  INVX1 U799 ( .A(n542), .Y(y2[12]) );
  AOI22X1 U800 ( .A0(N1683), .A1(n156), .B0(y2_tmp[12]), .B1(n100), .Y(n542)
         );
  INVX1 U801 ( .A(n520), .Y(y3[12]) );
  AOI22X1 U802 ( .A0(N1705), .A1(n147), .B0(y3_tmp[12]), .B1(n102), .Y(n520)
         );
  BUFX3 U803 ( .A(x4[3]), .Y(n77) );
  BUFX3 U804 ( .A(x5[3]), .Y(n64) );
  BUFX3 U805 ( .A(x6[3]), .Y(n51) );
  BUFX3 U806 ( .A(x7[3]), .Y(n38) );
  BUFX3 U807 ( .A(x4[2]), .Y(n76) );
  BUFX3 U808 ( .A(x5[2]), .Y(n63) );
  BUFX3 U809 ( .A(x6[2]), .Y(n50) );
  INVX1 U810 ( .A(n497), .Y(y4[13]) );
  INVX1 U811 ( .A(n475), .Y(y5[13]) );
  INVX1 U812 ( .A(n453), .Y(y6[13]) );
  ADDFX2 U813 ( .A(x4[1]), .B(n76), .CI(add_73_carry_5_), .CO(add_73_carry_6_), 
        .S(N45) );
  ADDFX2 U814 ( .A(x5[1]), .B(n63), .CI(add_82_carry_5_), .CO(add_82_carry_6_), 
        .S(N130) );
  ADDFX2 U815 ( .A(x6[1]), .B(n50), .CI(add_91_carry_5_), .CO(add_91_carry_6_), 
        .S(N215) );
  ADDFX2 U816 ( .A(x7[1]), .B(n39), .CI(add_104_carry_5_), .CO(
        add_104_carry_6_), .S(N341) );
  ADDFX2 U817 ( .A(x5[1]), .B(n65), .CI(add_86_carry_5_), .CO(add_86_carry_6_), 
        .S(N171) );
  ADDFX2 U818 ( .A(x6[1]), .B(n52), .CI(add_95_carry_5_), .CO(add_95_carry_6_), 
        .S(N256) );
  ADDFX2 U819 ( .A(x4[1]), .B(n78), .CI(add_77_carry_5_), .CO(add_77_carry_6_), 
        .S(N86) );
  ADDFX2 U820 ( .A(x7[1]), .B(n38), .CI(add_102_carry_4_), .CO(
        add_102_carry_5_), .S(N320) );
  ADDFX2 U821 ( .A(x6[1]), .B(n51), .CI(add_93_carry_4_), .CO(add_93_carry_5_), 
        .S(N235) );
  ADDFX2 U822 ( .A(x5[1]), .B(n64), .CI(add_84_carry_4_), .CO(add_84_carry_5_), 
        .S(N150) );
  ADDFX2 U823 ( .A(x4[1]), .B(n77), .CI(add_75_carry_4_), .CO(add_75_carry_5_), 
        .S(N65) );
  ADDFX2 U824 ( .A(x7[1]), .B(n37), .CI(add_100_carry_5_), .CO(
        add_100_carry_6_), .S(N300) );
  ADDFX2 U825 ( .A(x7[1]), .B(n42), .CI(add_99_carry_7_), .CO(add_99_carry_8_), 
        .S(N279) );
  BUFX3 U826 ( .A(x7[2]), .Y(n37) );
  NAND2BX1 U827 ( .AN(mode_delay2[1]), .B(mode_delay2[0]), .Y(n414) );
  AOI22X1 U828 ( .A0(N1723), .A1(n131), .B0(y4_tmp[8]), .B1(n94), .Y(n481) );
  AOI22X1 U829 ( .A0(N1724), .A1(n131), .B0(y4_tmp[9]), .B1(n94), .Y(n480) );
  AOI22X1 U830 ( .A0(N1725), .A1(n139), .B0(y4_tmp[10]), .B1(n96), .Y(n500) );
  AOI22X1 U831 ( .A0(N1726), .A1(n138), .B0(y4_tmp[11]), .B1(n96), .Y(n499) );
  AOI22X1 U832 ( .A0(N1727), .A1(n138), .B0(y4_tmp[12]), .B1(n96), .Y(n498) );
  AOI22X1 U833 ( .A0(N1745), .A1(n122), .B0(y5_tmp[8]), .B1(n92), .Y(n459) );
  AOI22X1 U834 ( .A0(N1746), .A1(n122), .B0(y5_tmp[9]), .B1(n92), .Y(n458) );
  AOI22X1 U835 ( .A0(N1747), .A1(n130), .B0(y5_tmp[10]), .B1(n94), .Y(n478) );
  AOI22X1 U836 ( .A0(N1748), .A1(n129), .B0(y5_tmp[11]), .B1(n94), .Y(n477) );
  AOI22X1 U837 ( .A0(N1749), .A1(n129), .B0(y5_tmp[12]), .B1(n94), .Y(n476) );
  AOI22X1 U838 ( .A0(N1767), .A1(n113), .B0(y6_tmp[8]), .B1(n90), .Y(n437) );
  AOI22X1 U839 ( .A0(N1768), .A1(n113), .B0(y6_tmp[9]), .B1(n90), .Y(n436) );
  AOI22X1 U840 ( .A0(N1769), .A1(n121), .B0(y6_tmp[10]), .B1(n92), .Y(n456) );
  AOI22X1 U841 ( .A0(N1770), .A1(n120), .B0(y6_tmp[11]), .B1(n92), .Y(n455) );
  AOI22X1 U842 ( .A0(N1771), .A1(n120), .B0(y6_tmp[12]), .B1(n92), .Y(n454) );
  AOI22X1 U843 ( .A0(N1789), .A1(n104), .B0(y7_tmp[8]), .B1(n89), .Y(n415) );
  AOI22X1 U844 ( .A0(N1790), .A1(n104), .B0(y7_tmp[9]), .B1(n97), .Y(n413) );
  AOI22X1 U845 ( .A0(N1791), .A1(n112), .B0(y7_tmp[10]), .B1(n90), .Y(n434) );
  AOI22X1 U846 ( .A0(N1792), .A1(n111), .B0(y7_tmp[11]), .B1(n90), .Y(n433) );
  AOI22X1 U847 ( .A0(N1793), .A1(n111), .B0(y7_tmp[12]), .B1(n90), .Y(n432) );
  INVX1 U848 ( .A(n589), .Y(y0[0]) );
  AOI22X1 U849 ( .A0(N1627), .A1(n176), .B0(y0_tmp[0]), .B1(n89), .Y(n589) );
  INVX1 U850 ( .A(n573), .Y(y0[4]) );
  AOI22X1 U851 ( .A0(N1631), .A1(n169), .B0(y0_tmp[4]), .B1(n98), .Y(n573) );
  INVX1 U852 ( .A(n571), .Y(y0[6]) );
  AOI22X1 U853 ( .A0(N1633), .A1(n168), .B0(y0_tmp[6]), .B1(n98), .Y(n571) );
  INVX1 U854 ( .A(n551), .Y(y1[4]) );
  AOI22X1 U855 ( .A0(N1653), .A1(n160), .B0(y1_tmp[4]), .B1(n100), .Y(n551) );
  INVX1 U856 ( .A(n549), .Y(y1[6]) );
  AOI22X1 U857 ( .A0(N1655), .A1(n159), .B0(y1_tmp[6]), .B1(n100), .Y(n549) );
  INVX1 U858 ( .A(n529), .Y(y2[4]) );
  AOI22X1 U859 ( .A0(N1675), .A1(n151), .B0(y2_tmp[4]), .B1(n102), .Y(n529) );
  INVX1 U860 ( .A(n527), .Y(y2[6]) );
  AOI22X1 U861 ( .A0(N1677), .A1(n150), .B0(y2_tmp[6]), .B1(n102), .Y(n527) );
  INVX1 U862 ( .A(n507), .Y(y3[4]) );
  AOI22X1 U863 ( .A0(N1697), .A1(n142), .B0(y3_tmp[4]), .B1(n96), .Y(n507) );
  INVX1 U864 ( .A(n506), .Y(y3[5]) );
  AOI22X1 U865 ( .A0(N1698), .A1(n142), .B0(y3_tmp[5]), .B1(n96), .Y(n506) );
  INVX1 U866 ( .A(n505), .Y(y3[6]) );
  AOI22X1 U867 ( .A0(N1699), .A1(n141), .B0(y3_tmp[6]), .B1(n96), .Y(n505) );
  INVX1 U868 ( .A(n504), .Y(y3[7]) );
  AOI22X1 U869 ( .A0(N1700), .A1(n141), .B0(y3_tmp[7]), .B1(n96), .Y(n504) );
  BUFX3 U870 ( .A(x5[9]), .Y(n70) );
  BUFX3 U871 ( .A(x5[10]), .Y(n71) );
  BUFX3 U872 ( .A(x5[11]), .Y(n72) );
  BUFX3 U873 ( .A(x5[12]), .Y(n73) );
  BUFX3 U874 ( .A(x6[9]), .Y(n57) );
  BUFX3 U875 ( .A(x6[10]), .Y(n58) );
  BUFX3 U876 ( .A(x6[11]), .Y(n59) );
  BUFX3 U877 ( .A(x6[12]), .Y(n60) );
  BUFX3 U878 ( .A(x4[9]), .Y(n83) );
  BUFX3 U879 ( .A(x4[10]), .Y(n84) );
  BUFX3 U880 ( .A(x4[11]), .Y(n85) );
  BUFX3 U881 ( .A(x4[12]), .Y(n86) );
  BUFX3 U882 ( .A(x7[9]), .Y(n44) );
  BUFX3 U883 ( .A(x7[10]), .Y(n45) );
  BUFX3 U884 ( .A(x7[11]), .Y(n46) );
  BUFX3 U885 ( .A(x7[12]), .Y(n47) );
  INVX1 U886 ( .A(n572), .Y(y0[5]) );
  AOI22X1 U887 ( .A0(N1632), .A1(n169), .B0(y0_tmp[5]), .B1(n98), .Y(n572) );
  INVX1 U888 ( .A(n570), .Y(y0[7]) );
  AOI22X1 U889 ( .A0(N1634), .A1(n168), .B0(y0_tmp[7]), .B1(n98), .Y(n570) );
  INVX1 U890 ( .A(n550), .Y(y1[5]) );
  AOI22X1 U891 ( .A0(N1654), .A1(n160), .B0(y1_tmp[5]), .B1(n100), .Y(n550) );
  INVX1 U892 ( .A(n548), .Y(y1[7]) );
  AOI22X1 U893 ( .A0(N1656), .A1(n159), .B0(y1_tmp[7]), .B1(n100), .Y(n548) );
  INVX1 U894 ( .A(n528), .Y(y2[5]) );
  AOI22X1 U895 ( .A0(N1676), .A1(n151), .B0(y2_tmp[5]), .B1(n102), .Y(n528) );
  INVX1 U896 ( .A(n526), .Y(y2[7]) );
  AOI22X1 U897 ( .A0(N1678), .A1(n150), .B0(y2_tmp[7]), .B1(n102), .Y(n526) );
  INVX1 U898 ( .A(n512), .Y(y3[1]) );
  AOI22X1 U899 ( .A0(N1694), .A1(n144), .B0(y3_tmp[1]), .B1(n103), .Y(n512) );
  INVX1 U900 ( .A(n485), .Y(y4[4]) );
  INVX1 U901 ( .A(n484), .Y(y4[5]) );
  INVX1 U902 ( .A(n483), .Y(y4[6]) );
  INVX1 U903 ( .A(n482), .Y(y4[7]) );
  INVX1 U904 ( .A(n481), .Y(y4[8]) );
  INVX1 U905 ( .A(n480), .Y(y4[9]) );
  INVX1 U906 ( .A(n500), .Y(y4[10]) );
  INVX1 U907 ( .A(n499), .Y(y4[11]) );
  INVX1 U908 ( .A(n498), .Y(y4[12]) );
  INVX1 U909 ( .A(n479), .Y(y5[0]) );
  INVX1 U910 ( .A(n468), .Y(y5[1]) );
  INVX1 U911 ( .A(n465), .Y(y5[2]) );
  INVX1 U912 ( .A(n464), .Y(y5[3]) );
  INVX1 U913 ( .A(n463), .Y(y5[4]) );
  INVX1 U914 ( .A(n462), .Y(y5[5]) );
  INVX1 U915 ( .A(n461), .Y(y5[6]) );
  INVX1 U916 ( .A(n460), .Y(y5[7]) );
  INVX1 U917 ( .A(n459), .Y(y5[8]) );
  INVX1 U918 ( .A(n458), .Y(y5[9]) );
  INVX1 U919 ( .A(n478), .Y(y5[10]) );
  INVX1 U920 ( .A(n477), .Y(y5[11]) );
  INVX1 U921 ( .A(n476), .Y(y5[12]) );
  INVX1 U922 ( .A(n457), .Y(y6[0]) );
  INVX1 U923 ( .A(n446), .Y(y6[1]) );
  INVX1 U924 ( .A(n443), .Y(y6[2]) );
  INVX1 U925 ( .A(n442), .Y(y6[3]) );
  INVX1 U926 ( .A(n441), .Y(y6[4]) );
  INVX1 U927 ( .A(n440), .Y(y6[5]) );
  INVX1 U928 ( .A(n439), .Y(y6[6]) );
  INVX1 U929 ( .A(n438), .Y(y6[7]) );
  INVX1 U930 ( .A(n437), .Y(y6[8]) );
  INVX1 U931 ( .A(n436), .Y(y6[9]) );
  INVX1 U932 ( .A(n456), .Y(y6[10]) );
  INVX1 U933 ( .A(n455), .Y(y6[11]) );
  INVX1 U934 ( .A(n454), .Y(y6[12]) );
  INVX1 U935 ( .A(n501), .Y(y4[0]) );
  INVX1 U936 ( .A(n490), .Y(y4[1]) );
  INVX1 U937 ( .A(n487), .Y(y4[2]) );
  INVX1 U938 ( .A(n486), .Y(y4[3]) );
  INVX1 U939 ( .A(n578), .Y(y0[1]) );
  AOI22X1 U940 ( .A0(N1628), .A1(n171), .B0(y0_tmp[1]), .B1(n97), .Y(n578) );
  INVX1 U941 ( .A(n575), .Y(y0[2]) );
  AOI22X1 U942 ( .A0(N1629), .A1(n170), .B0(y0_tmp[2]), .B1(n98), .Y(n575) );
  INVX1 U943 ( .A(n574), .Y(y0[3]) );
  AOI22X1 U944 ( .A0(N1630), .A1(n170), .B0(y0_tmp[3]), .B1(n98), .Y(n574) );
  INVX1 U945 ( .A(n567), .Y(y1[0]) );
  AOI22X1 U946 ( .A0(N1649), .A1(n166), .B0(y1_tmp[0]), .B1(n98), .Y(n567) );
  INVX1 U947 ( .A(n556), .Y(y1[1]) );
  AOI22X1 U948 ( .A0(N1650), .A1(n162), .B0(y1_tmp[1]), .B1(n99), .Y(n556) );
  INVX1 U949 ( .A(n553), .Y(y1[2]) );
  AOI22X1 U950 ( .A0(N1651), .A1(n161), .B0(y1_tmp[2]), .B1(n99), .Y(n553) );
  INVX1 U951 ( .A(n552), .Y(y1[3]) );
  AOI22X1 U952 ( .A0(N1652), .A1(n161), .B0(y1_tmp[3]), .B1(n100), .Y(n552) );
  INVX1 U953 ( .A(n545), .Y(y2[0]) );
  AOI22X1 U954 ( .A0(N1671), .A1(n157), .B0(y2_tmp[0]), .B1(n100), .Y(n545) );
  INVX1 U955 ( .A(n534), .Y(y2[1]) );
  AOI22X1 U956 ( .A0(N1672), .A1(n153), .B0(y2_tmp[1]), .B1(n101), .Y(n534) );
  INVX1 U957 ( .A(n531), .Y(y2[2]) );
  AOI22X1 U958 ( .A0(N1673), .A1(n152), .B0(y2_tmp[2]), .B1(n102), .Y(n531) );
  INVX1 U959 ( .A(n530), .Y(y2[3]) );
  AOI22X1 U960 ( .A0(N1674), .A1(n152), .B0(y2_tmp[3]), .B1(n101), .Y(n530) );
  INVX1 U961 ( .A(n523), .Y(y3[0]) );
  AOI22X1 U962 ( .A0(N1693), .A1(n148), .B0(y3_tmp[0]), .B1(n101), .Y(n523) );
  INVX1 U963 ( .A(n509), .Y(y3[2]) );
  AOI22X1 U964 ( .A0(N1695), .A1(n143), .B0(y3_tmp[2]), .B1(n96), .Y(n509) );
  INVX1 U965 ( .A(n508), .Y(y3[3]) );
  AOI22X1 U966 ( .A0(N1696), .A1(n143), .B0(y3_tmp[3]), .B1(n96), .Y(n508) );
  INVX1 U967 ( .A(n435), .Y(y7[0]) );
  INVX1 U968 ( .A(n424), .Y(y7[1]) );
  INVX1 U969 ( .A(n421), .Y(y7[2]) );
  INVX1 U970 ( .A(n420), .Y(y7[3]) );
  INVX1 U971 ( .A(n419), .Y(y7[4]) );
  INVX1 U972 ( .A(n418), .Y(y7[5]) );
  INVX1 U973 ( .A(n417), .Y(y7[6]) );
  INVX1 U974 ( .A(n416), .Y(y7[7]) );
  INVX1 U975 ( .A(n415), .Y(y7[8]) );
  INVX1 U976 ( .A(n413), .Y(y7[9]) );
  INVX1 U977 ( .A(n434), .Y(y7[10]) );
  INVX1 U978 ( .A(n433), .Y(y7[11]) );
  INVX1 U979 ( .A(n432), .Y(y7[12]) );
  AOI22X1 U980 ( .A0(N1715), .A1(n139), .B0(y4_tmp[0]), .B1(n96), .Y(n501) );
  AOI22X1 U981 ( .A0(N1716), .A1(n135), .B0(y4_tmp[1]), .B1(n95), .Y(n490) );
  AOI22X1 U982 ( .A0(N1717), .A1(n134), .B0(y4_tmp[2]), .B1(n95), .Y(n487) );
  AOI22X1 U983 ( .A0(N1718), .A1(n134), .B0(y4_tmp[3]), .B1(n95), .Y(n486) );
  AOI22X1 U984 ( .A0(N1719), .A1(n133), .B0(y4_tmp[4]), .B1(n94), .Y(n485) );
  AOI22X1 U985 ( .A0(N1720), .A1(n133), .B0(y4_tmp[5]), .B1(n94), .Y(n484) );
  AOI22X1 U986 ( .A0(N1721), .A1(n132), .B0(y4_tmp[6]), .B1(n94), .Y(n483) );
  AOI22X1 U987 ( .A0(N1722), .A1(n132), .B0(y4_tmp[7]), .B1(n94), .Y(n482) );
  AOI22X1 U988 ( .A0(N1737), .A1(n130), .B0(y5_tmp[0]), .B1(n94), .Y(n479) );
  AOI22X1 U989 ( .A0(N1738), .A1(n126), .B0(y5_tmp[1]), .B1(n93), .Y(n468) );
  AOI22X1 U990 ( .A0(N1739), .A1(n125), .B0(y5_tmp[2]), .B1(n93), .Y(n465) );
  AOI22X1 U991 ( .A0(N1740), .A1(n125), .B0(y5_tmp[3]), .B1(n93), .Y(n464) );
  AOI22X1 U992 ( .A0(N1741), .A1(n124), .B0(y5_tmp[4]), .B1(n93), .Y(n463) );
  AOI22X1 U993 ( .A0(N1742), .A1(n124), .B0(y5_tmp[5]), .B1(n93), .Y(n462) );
  AOI22X1 U994 ( .A0(N1743), .A1(n123), .B0(y5_tmp[6]), .B1(n92), .Y(n461) );
  AOI22X1 U995 ( .A0(N1744), .A1(n123), .B0(y5_tmp[7]), .B1(n92), .Y(n460) );
  AOI22X1 U996 ( .A0(N1759), .A1(n121), .B0(y6_tmp[0]), .B1(n92), .Y(n457) );
  AOI22X1 U997 ( .A0(N1760), .A1(n117), .B0(y6_tmp[1]), .B1(n91), .Y(n446) );
  AOI22X1 U998 ( .A0(N1761), .A1(n116), .B0(y6_tmp[2]), .B1(n91), .Y(n443) );
  AOI22X1 U999 ( .A0(N1762), .A1(n116), .B0(y6_tmp[3]), .B1(n91), .Y(n442) );
  AOI22X1 U1000 ( .A0(N1763), .A1(n115), .B0(y6_tmp[4]), .B1(n91), .Y(n441) );
  AOI22X1 U1001 ( .A0(N1764), .A1(n115), .B0(y6_tmp[5]), .B1(n91), .Y(n440) );
  AOI22X1 U1002 ( .A0(N1765), .A1(n114), .B0(y6_tmp[6]), .B1(n91), .Y(n439) );
  AOI22X1 U1003 ( .A0(N1766), .A1(n114), .B0(y6_tmp[7]), .B1(n91), .Y(n438) );
  AOI22X1 U1004 ( .A0(N1781), .A1(n112), .B0(y7_tmp[0]), .B1(n90), .Y(n435) );
  AOI22X1 U1005 ( .A0(N1782), .A1(n108), .B0(y7_tmp[1]), .B1(n89), .Y(n424) );
  AOI22X1 U1006 ( .A0(N1783), .A1(n107), .B0(y7_tmp[2]), .B1(n89), .Y(n421) );
  AOI22X1 U1007 ( .A0(N1784), .A1(n107), .B0(y7_tmp[3]), .B1(n89), .Y(n420) );
  AOI22X1 U1008 ( .A0(N1785), .A1(n106), .B0(y7_tmp[4]), .B1(n89), .Y(n419) );
  AOI22X1 U1009 ( .A0(N1786), .A1(n106), .B0(y7_tmp[5]), .B1(n89), .Y(n418) );
  AOI22X1 U1010 ( .A0(N1787), .A1(n105), .B0(y7_tmp[6]), .B1(n89), .Y(n417) );
  AOI22X1 U1011 ( .A0(N1788), .A1(n105), .B0(y7_tmp[7]), .B1(n89), .Y(n416) );
  BUFX3 U1012 ( .A(x5[13]), .Y(n74) );
  BUFX3 U1013 ( .A(x5[14]), .Y(n75) );
  BUFX3 U1014 ( .A(x6[13]), .Y(n61) );
  BUFX3 U1015 ( .A(x6[14]), .Y(n62) );
  BUFX3 U1016 ( .A(x4[13]), .Y(n87) );
  BUFX3 U1017 ( .A(x4[14]), .Y(n88) );
  BUFX3 U1018 ( .A(x7[13]), .Y(n48) );
  BUFX3 U1019 ( .A(x7[14]), .Y(n49) );
  INVX1 U1020 ( .A(x7_50[21]), .Y(n226) );
  INVX1 U1021 ( .A(x5_50[21]), .Y(n294) );
  INVX1 U1022 ( .A(x5_tmp[24]), .Y(n341) );
  INVX1 U1023 ( .A(x4_tmp[24]), .Y(n592) );
  INVX1 U1024 ( .A(x7_tmp[24]), .Y(n340) );
  INVX1 U1025 ( .A(x6_tmp[24]), .Y(n366) );
  INVX1 U1026 ( .A(x7_89[22]), .Y(n271) );
  INVX1 U1027 ( .A(x5_89[22]), .Y(n248) );
  AOI22X1 U1028 ( .A0(N1643), .A1(n173), .B0(y0_tmp[16]), .B1(n97), .Y(n582)
         );
  AOI22X1 U1029 ( .A0(N1644), .A1(n172), .B0(y0_tmp[17]), .B1(n97), .Y(n581)
         );
  AOI22X1 U1030 ( .A0(N1645), .A1(n172), .B0(y0_tmp[18]), .B1(n97), .Y(n580)
         );
  AOI22X1 U1031 ( .A0(N1646), .A1(n171), .B0(y0_tmp[19]), .B1(n97), .Y(n579)
         );
  AOI22X1 U1032 ( .A0(N1647), .A1(n172), .B0(y0_tmp[20]), .B1(n97), .Y(n577)
         );
  AOI22X1 U1033 ( .A0(N1648), .A1(n172), .B0(y0_tmp[21]), .B1(n98), .Y(n576)
         );
  AOI22X1 U1034 ( .A0(N1665), .A1(n163), .B0(y1_tmp[16]), .B1(n99), .Y(n560)
         );
  AOI22X1 U1035 ( .A0(N1666), .A1(n172), .B0(y1_tmp[17]), .B1(n99), .Y(n559)
         );
  AOI22X1 U1036 ( .A0(N1667), .A1(n172), .B0(y1_tmp[18]), .B1(n99), .Y(n558)
         );
  AOI22X1 U1037 ( .A0(N1668), .A1(n162), .B0(y1_tmp[19]), .B1(n99), .Y(n557)
         );
  AOI22X1 U1038 ( .A0(N1669), .A1(n172), .B0(y1_tmp[20]), .B1(n99), .Y(n555)
         );
  AOI22X1 U1039 ( .A0(N1670), .A1(n172), .B0(y1_tmp[21]), .B1(n99), .Y(n554)
         );
  AOI22X1 U1040 ( .A0(N1687), .A1(n154), .B0(y2_tmp[16]), .B1(n101), .Y(n538)
         );
  AOI22X1 U1041 ( .A0(N1688), .A1(n172), .B0(y2_tmp[17]), .B1(n101), .Y(n537)
         );
  AOI22X1 U1042 ( .A0(N1689), .A1(n172), .B0(y2_tmp[18]), .B1(n101), .Y(n536)
         );
  AOI22X1 U1043 ( .A0(N1690), .A1(n153), .B0(y2_tmp[19]), .B1(n101), .Y(n535)
         );
  AOI22X1 U1044 ( .A0(N1691), .A1(n172), .B0(y2_tmp[20]), .B1(n101), .Y(n533)
         );
  AOI22X1 U1045 ( .A0(N1692), .A1(n172), .B0(y2_tmp[21]), .B1(n101), .Y(n532)
         );
  AOI22X1 U1046 ( .A0(N1709), .A1(n145), .B0(y3_tmp[16]), .B1(n102), .Y(n516)
         );
  AOI22X1 U1047 ( .A0(N1710), .A1(n172), .B0(y3_tmp[17]), .B1(n103), .Y(n515)
         );
  AOI22X1 U1048 ( .A0(N1711), .A1(n172), .B0(y3_tmp[18]), .B1(n103), .Y(n514)
         );
  AOI22X1 U1049 ( .A0(N1712), .A1(n144), .B0(y3_tmp[19]), .B1(n103), .Y(n513)
         );
  AOI22X1 U1050 ( .A0(N1713), .A1(n172), .B0(y3_tmp[20]), .B1(n102), .Y(n511)
         );
  AOI22X1 U1051 ( .A0(N1714), .A1(n172), .B0(y3_tmp[21]), .B1(n103), .Y(n510)
         );
  AOI22X1 U1052 ( .A0(N1731), .A1(n136), .B0(y4_tmp[16]), .B1(n95), .Y(n494)
         );
  AOI22X1 U1053 ( .A0(N1732), .A1(n172), .B0(y4_tmp[17]), .B1(n95), .Y(n493)
         );
  AOI22X1 U1054 ( .A0(N1733), .A1(n172), .B0(y4_tmp[18]), .B1(n95), .Y(n492)
         );
  AOI22X1 U1055 ( .A0(N1734), .A1(n135), .B0(y4_tmp[19]), .B1(n95), .Y(n491)
         );
  AOI22X1 U1056 ( .A0(N1735), .A1(n172), .B0(y4_tmp[20]), .B1(n95), .Y(n489)
         );
  AOI22X1 U1057 ( .A0(N1736), .A1(n172), .B0(y4_tmp[21]), .B1(n95), .Y(n488)
         );
  AOI22X1 U1058 ( .A0(N1753), .A1(n127), .B0(y5_tmp[16]), .B1(n93), .Y(n472)
         );
  AOI22X1 U1059 ( .A0(N1754), .A1(n172), .B0(y5_tmp[17]), .B1(n93), .Y(n471)
         );
  AOI22X1 U1060 ( .A0(N1755), .A1(n172), .B0(y5_tmp[18]), .B1(n93), .Y(n470)
         );
  AOI22X1 U1061 ( .A0(N1756), .A1(n126), .B0(y5_tmp[19]), .B1(n93), .Y(n469)
         );
  AOI22X1 U1062 ( .A0(N1757), .A1(n172), .B0(y5_tmp[20]), .B1(n93), .Y(n467)
         );
  AOI22X1 U1063 ( .A0(N1758), .A1(n172), .B0(y5_tmp[21]), .B1(n93), .Y(n466)
         );
  AOI22X1 U1064 ( .A0(N1775), .A1(n118), .B0(y6_tmp[16]), .B1(n92), .Y(n450)
         );
  AOI22X1 U1065 ( .A0(N1776), .A1(n172), .B0(y6_tmp[17]), .B1(n91), .Y(n449)
         );
  AOI22X1 U1066 ( .A0(N1777), .A1(n172), .B0(y6_tmp[18]), .B1(n91), .Y(n448)
         );
  AOI22X1 U1067 ( .A0(N1778), .A1(n117), .B0(y6_tmp[19]), .B1(n91), .Y(n447)
         );
  AOI22X1 U1068 ( .A0(N1779), .A1(n172), .B0(y6_tmp[20]), .B1(n91), .Y(n445)
         );
  AOI22X1 U1069 ( .A0(N1780), .A1(n172), .B0(y6_tmp[21]), .B1(n91), .Y(n444)
         );
  AOI22X1 U1070 ( .A0(N1797), .A1(n109), .B0(y7_tmp[16]), .B1(n90), .Y(n428)
         );
  AOI22X1 U1071 ( .A0(N1798), .A1(n172), .B0(y7_tmp[17]), .B1(n90), .Y(n427)
         );
  AOI22X1 U1072 ( .A0(N1799), .A1(n172), .B0(y7_tmp[18]), .B1(n90), .Y(n426)
         );
  AOI22X1 U1073 ( .A0(N1800), .A1(n108), .B0(y7_tmp[19]), .B1(n89), .Y(n425)
         );
  AOI22X1 U1074 ( .A0(N1801), .A1(n172), .B0(y7_tmp[20]), .B1(n89), .Y(n423)
         );
  AOI22X1 U1075 ( .A0(N1802), .A1(n172), .B0(y7_tmp[21]), .B1(n89), .Y(n422)
         );
  AND2X1 U1100 ( .A(x7[0]), .B(n38), .Y(add_104_carry_5_) );
  XOR2X1 U1101 ( .A(n38), .B(x7[0]), .Y(N340) );
  AND2X1 U1102 ( .A(x5[0]), .B(n64), .Y(add_86_carry_5_) );
  XOR2X1 U1103 ( .A(n64), .B(x5[0]), .Y(N170) );
  AND2X1 U1104 ( .A(x6[0]), .B(n51), .Y(add_95_carry_5_) );
  XOR2X1 U1105 ( .A(n51), .B(x6[0]), .Y(N255) );
  AND2X1 U1106 ( .A(x4[0]), .B(n77), .Y(add_77_carry_5_) );
  XOR2X1 U1107 ( .A(n77), .B(x4[0]), .Y(N85) );
  AND2X1 U1108 ( .A(x7[0]), .B(n37), .Y(add_102_carry_4_) );
  XOR2X1 U1109 ( .A(n37), .B(x7[0]), .Y(N319) );
  AND2X1 U1110 ( .A(x6[0]), .B(n50), .Y(add_93_carry_4_) );
  XOR2X1 U1111 ( .A(n50), .B(x6[0]), .Y(N234) );
  AND2X1 U1112 ( .A(x5[0]), .B(n63), .Y(add_84_carry_4_) );
  XOR2X1 U1113 ( .A(n63), .B(x5[0]), .Y(N149) );
  AND2X1 U1114 ( .A(x4[0]), .B(n76), .Y(add_75_carry_4_) );
  XOR2X1 U1115 ( .A(n76), .B(x4[0]), .Y(N64) );
  AND2X1 U1116 ( .A(x7[0]), .B(x7[1]), .Y(add_100_carry_5_) );
  XOR2X1 U1117 ( .A(x7[1]), .B(x7[0]), .Y(N299) );
  AND2X1 U1118 ( .A(x4[0]), .B(n80), .Y(add_72_carry_7_) );
  XOR2X1 U1119 ( .A(n80), .B(x4[0]), .Y(N23) );
  AND2X1 U1120 ( .A(x4[0]), .B(x4[1]), .Y(add_73_carry_5_) );
  XOR2X1 U1121 ( .A(x4[1]), .B(x4[0]), .Y(N44) );
  AND2X1 U1122 ( .A(x5[0]), .B(x5[1]), .Y(add_82_carry_5_) );
  XOR2X1 U1123 ( .A(x5[1]), .B(x5[0]), .Y(N129) );
  AND2X1 U1124 ( .A(x6[0]), .B(x6[1]), .Y(add_91_carry_5_) );
  XOR2X1 U1125 ( .A(x6[1]), .B(x6[0]), .Y(N214) );
  AND2X1 U1126 ( .A(x5[0]), .B(n67), .Y(add_81_carry_7_) );
  XOR2X1 U1127 ( .A(n67), .B(x5[0]), .Y(N108) );
  AND2X1 U1128 ( .A(x6[0]), .B(n54), .Y(add_90_carry_7_) );
  XOR2X1 U1129 ( .A(n54), .B(x6[0]), .Y(N193) );
  AND2X1 U1130 ( .A(x7[0]), .B(n41), .Y(add_99_carry_7_) );
  XOR2X1 U1131 ( .A(n41), .B(x7[0]), .Y(N278) );
endmodule


module idct_cal_shift7_add64 ( clk, rstn, mode, start, x0, x1, x2, x3, x4, x5, 
        x6, x7, y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, 
        y14, y15, idct_ready, mode_out );
  input [1:0] mode;
  input [15:0] x0;
  input [15:0] x1;
  input [15:0] x2;
  input [15:0] x3;
  input [15:0] x4;
  input [15:0] x5;
  input [15:0] x6;
  input [15:0] x7;
  output [15:0] y0;
  output [15:0] y1;
  output [15:0] y2;
  output [15:0] y3;
  output [15:0] y4;
  output [15:0] y5;
  output [15:0] y6;
  output [15:0] y7;
  output [15:0] y8;
  output [15:0] y9;
  output [15:0] y10;
  output [15:0] y11;
  output [15:0] y12;
  output [15:0] y13;
  output [15:0] y14;
  output [15:0] y15;
  output [1:0] mode_out;
  input clk, rstn, start;
  output idct_ready;
  wire   idct4_ready, idct8_ready, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n325, n326, n327, n328, n329, n330, n331, n332;
  wire   [1:0] mode_delay2;
  wire   [1:0] mode_delay1;
  wire   [24:0] y0_idct4;
  wire   [24:0] y1_idct4;
  wire   [24:0] y2_idct4;
  wire   [24:0] y3_idct4;
  wire   [15:0] y0_idct8;
  wire   [15:0] y1_idct8;
  wire   [15:0] y2_idct8;
  wire   [15:0] y3_idct8;
  wire   [15:0] y4_idct8;
  wire   [15:0] y5_idct8;
  wire   [15:0] y6_idct8;
  wire   [15:0] y7_idct8;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75, 
        SYNOPSYS_UNCONNECTED__76, SYNOPSYS_UNCONNECTED__77, 
        SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79;

  CLKINVX8 U3 ( .A(n2), .Y(mode_out[0]) );
  AOI22X4 U4 ( .A0(idct_ready), .A1(mode_delay2[0]), .B0(n3), .B1(mode_out[0]), 
        .Y(n2) );
  NOR2BX4 U5 ( .AN(mode_out[1]), .B(idct_ready), .Y(mode_out[1]) );
  idct4_shift7_add64 idct4_cal ( .clk(clk), .rstn(rstn), .mode(mode), .start(
        start), .x0(x0), .x1(x1), .x2(x2), .x3(x3), .y0(y0_idct4), .y1(
        y1_idct4), .y2(y2_idct4), .y3(y3_idct4), .idct4_ready(idct4_ready) );
  idct8_shift7_add64 idct8_cal ( .clk(clk), .rstn(rstn), .mode(mode), .start(
        idct4_ready), .x0(y0_idct4), .x1(y1_idct4), .x2(y2_idct4), .x3(
        y3_idct4), .x4(x4), .x5(x5), .x6(x6), .x7(x7), .y0({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, y0_idct8}), .y1({
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, y1_idct8}), .y2({
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, y2_idct8}), .y3({
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, y3_idct8}), .y4({
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, y4_idct8}), .y5({
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, y5_idct8}), .y6({
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, y6_idct8}), .y7({
        SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75, 
        SYNOPSYS_UNCONNECTED__76, SYNOPSYS_UNCONNECTED__77, 
        SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79, y7_idct8}), 
        .idct8_ready(idct8_ready) );
  DFFRHQX1 mode_delay2_reg_1_ ( .D(mode_delay1[1]), .CK(clk), .RN(rstn), .Q(
        mode_delay2[1]) );
  DFFRHQX1 mode_delay2_reg_0_ ( .D(mode_delay1[0]), .CK(clk), .RN(rstn), .Q(
        mode_delay2[0]) );
  DFFRHQX1 mode_delay1_reg_1_ ( .D(mode[1]), .CK(clk), .RN(rstn), .Q(
        mode_delay1[1]) );
  DFFRHQX1 mode_delay1_reg_0_ ( .D(mode[0]), .CK(clk), .RN(rstn), .Q(
        mode_delay1[0]) );
  INVX1 U6 ( .A(1'b1), .Y(y15[0]) );
  INVX1 U8 ( .A(1'b1), .Y(y15[1]) );
  INVX1 U10 ( .A(1'b1), .Y(y15[2]) );
  INVX1 U12 ( .A(1'b1), .Y(y15[3]) );
  INVX1 U14 ( .A(1'b1), .Y(y15[4]) );
  INVX1 U16 ( .A(1'b1), .Y(y15[5]) );
  INVX1 U18 ( .A(1'b1), .Y(y15[6]) );
  INVX1 U20 ( .A(1'b1), .Y(y15[7]) );
  INVX1 U22 ( .A(1'b1), .Y(y15[8]) );
  INVX1 U24 ( .A(1'b1), .Y(y15[9]) );
  INVX1 U26 ( .A(1'b1), .Y(y15[10]) );
  INVX1 U28 ( .A(1'b1), .Y(y15[11]) );
  INVX1 U30 ( .A(1'b1), .Y(y15[12]) );
  INVX1 U32 ( .A(1'b1), .Y(y15[13]) );
  INVX1 U34 ( .A(1'b1), .Y(y15[14]) );
  INVX1 U36 ( .A(1'b1), .Y(y15[15]) );
  INVX1 U38 ( .A(1'b1), .Y(y14[0]) );
  INVX1 U40 ( .A(1'b1), .Y(y14[1]) );
  INVX1 U42 ( .A(1'b1), .Y(y14[2]) );
  INVX1 U44 ( .A(1'b1), .Y(y14[3]) );
  INVX1 U46 ( .A(1'b1), .Y(y14[4]) );
  INVX1 U48 ( .A(1'b1), .Y(y14[5]) );
  INVX1 U50 ( .A(1'b1), .Y(y14[6]) );
  INVX1 U52 ( .A(1'b1), .Y(y14[7]) );
  INVX1 U54 ( .A(1'b1), .Y(y14[8]) );
  INVX1 U56 ( .A(1'b1), .Y(y14[9]) );
  INVX1 U58 ( .A(1'b1), .Y(y14[10]) );
  INVX1 U60 ( .A(1'b1), .Y(y14[11]) );
  INVX1 U62 ( .A(1'b1), .Y(y14[12]) );
  INVX1 U64 ( .A(1'b1), .Y(y14[13]) );
  INVX1 U66 ( .A(1'b1), .Y(y14[14]) );
  INVX1 U68 ( .A(1'b1), .Y(y14[15]) );
  INVX1 U70 ( .A(1'b1), .Y(y13[0]) );
  INVX1 U72 ( .A(1'b1), .Y(y13[1]) );
  INVX1 U74 ( .A(1'b1), .Y(y13[2]) );
  INVX1 U76 ( .A(1'b1), .Y(y13[3]) );
  INVX1 U78 ( .A(1'b1), .Y(y13[4]) );
  INVX1 U80 ( .A(1'b1), .Y(y13[5]) );
  INVX1 U82 ( .A(1'b1), .Y(y13[6]) );
  INVX1 U84 ( .A(1'b1), .Y(y13[7]) );
  INVX1 U86 ( .A(1'b1), .Y(y13[8]) );
  INVX1 U88 ( .A(1'b1), .Y(y13[9]) );
  INVX1 U90 ( .A(1'b1), .Y(y13[10]) );
  INVX1 U92 ( .A(1'b1), .Y(y13[11]) );
  INVX1 U94 ( .A(1'b1), .Y(y13[12]) );
  INVX1 U96 ( .A(1'b1), .Y(y13[13]) );
  INVX1 U98 ( .A(1'b1), .Y(y13[14]) );
  INVX1 U100 ( .A(1'b1), .Y(y13[15]) );
  INVX1 U102 ( .A(1'b1), .Y(y12[0]) );
  INVX1 U104 ( .A(1'b1), .Y(y12[1]) );
  INVX1 U106 ( .A(1'b1), .Y(y12[2]) );
  INVX1 U108 ( .A(1'b1), .Y(y12[3]) );
  INVX1 U110 ( .A(1'b1), .Y(y12[4]) );
  INVX1 U112 ( .A(1'b1), .Y(y12[5]) );
  INVX1 U114 ( .A(1'b1), .Y(y12[6]) );
  INVX1 U116 ( .A(1'b1), .Y(y12[7]) );
  INVX1 U118 ( .A(1'b1), .Y(y12[8]) );
  INVX1 U120 ( .A(1'b1), .Y(y12[9]) );
  INVX1 U122 ( .A(1'b1), .Y(y12[10]) );
  INVX1 U124 ( .A(1'b1), .Y(y12[11]) );
  INVX1 U126 ( .A(1'b1), .Y(y12[12]) );
  INVX1 U128 ( .A(1'b1), .Y(y12[13]) );
  INVX1 U130 ( .A(1'b1), .Y(y12[14]) );
  INVX1 U132 ( .A(1'b1), .Y(y12[15]) );
  INVX1 U134 ( .A(1'b1), .Y(y11[0]) );
  INVX1 U136 ( .A(1'b1), .Y(y11[1]) );
  INVX1 U138 ( .A(1'b1), .Y(y11[2]) );
  INVX1 U140 ( .A(1'b1), .Y(y11[3]) );
  INVX1 U142 ( .A(1'b1), .Y(y11[4]) );
  INVX1 U144 ( .A(1'b1), .Y(y11[5]) );
  INVX1 U146 ( .A(1'b1), .Y(y11[6]) );
  INVX1 U148 ( .A(1'b1), .Y(y11[7]) );
  INVX1 U150 ( .A(1'b1), .Y(y11[8]) );
  INVX1 U152 ( .A(1'b1), .Y(y11[9]) );
  INVX1 U154 ( .A(1'b1), .Y(y11[10]) );
  INVX1 U156 ( .A(1'b1), .Y(y11[11]) );
  INVX1 U158 ( .A(1'b1), .Y(y11[12]) );
  INVX1 U160 ( .A(1'b1), .Y(y11[13]) );
  INVX1 U162 ( .A(1'b1), .Y(y11[14]) );
  INVX1 U164 ( .A(1'b1), .Y(y11[15]) );
  INVX1 U166 ( .A(1'b1), .Y(y10[0]) );
  INVX1 U168 ( .A(1'b1), .Y(y10[1]) );
  INVX1 U170 ( .A(1'b1), .Y(y10[2]) );
  INVX1 U172 ( .A(1'b1), .Y(y10[3]) );
  INVX1 U174 ( .A(1'b1), .Y(y10[4]) );
  INVX1 U176 ( .A(1'b1), .Y(y10[5]) );
  INVX1 U178 ( .A(1'b1), .Y(y10[6]) );
  INVX1 U180 ( .A(1'b1), .Y(y10[7]) );
  INVX1 U182 ( .A(1'b1), .Y(y10[8]) );
  INVX1 U184 ( .A(1'b1), .Y(y10[9]) );
  INVX1 U186 ( .A(1'b1), .Y(y10[10]) );
  INVX1 U188 ( .A(1'b1), .Y(y10[11]) );
  INVX1 U190 ( .A(1'b1), .Y(y10[12]) );
  INVX1 U192 ( .A(1'b1), .Y(y10[13]) );
  INVX1 U194 ( .A(1'b1), .Y(y10[14]) );
  INVX1 U196 ( .A(1'b1), .Y(y10[15]) );
  INVX1 U198 ( .A(1'b1), .Y(y9[0]) );
  INVX1 U200 ( .A(1'b1), .Y(y9[1]) );
  INVX1 U202 ( .A(1'b1), .Y(y9[2]) );
  INVX1 U204 ( .A(1'b1), .Y(y9[3]) );
  INVX1 U206 ( .A(1'b1), .Y(y9[4]) );
  INVX1 U208 ( .A(1'b1), .Y(y9[5]) );
  INVX1 U210 ( .A(1'b1), .Y(y9[6]) );
  INVX1 U212 ( .A(1'b1), .Y(y9[7]) );
  INVX1 U214 ( .A(1'b1), .Y(y9[8]) );
  INVX1 U216 ( .A(1'b1), .Y(y9[9]) );
  INVX1 U218 ( .A(1'b1), .Y(y9[10]) );
  INVX1 U220 ( .A(1'b1), .Y(y9[11]) );
  INVX1 U222 ( .A(1'b1), .Y(y9[12]) );
  INVX1 U224 ( .A(1'b1), .Y(y9[13]) );
  INVX1 U226 ( .A(1'b1), .Y(y9[14]) );
  INVX1 U228 ( .A(1'b1), .Y(y9[15]) );
  INVX1 U230 ( .A(1'b1), .Y(y8[0]) );
  INVX1 U232 ( .A(1'b1), .Y(y8[1]) );
  INVX1 U234 ( .A(1'b1), .Y(y8[2]) );
  INVX1 U236 ( .A(1'b1), .Y(y8[3]) );
  INVX1 U238 ( .A(1'b1), .Y(y8[4]) );
  INVX1 U240 ( .A(1'b1), .Y(y8[5]) );
  INVX1 U242 ( .A(1'b1), .Y(y8[6]) );
  INVX1 U244 ( .A(1'b1), .Y(y8[7]) );
  INVX1 U246 ( .A(1'b1), .Y(y8[8]) );
  INVX1 U248 ( .A(1'b1), .Y(y8[9]) );
  INVX1 U250 ( .A(1'b1), .Y(y8[10]) );
  INVX1 U252 ( .A(1'b1), .Y(y8[11]) );
  INVX1 U254 ( .A(1'b1), .Y(y8[12]) );
  INVX1 U256 ( .A(1'b1), .Y(y8[13]) );
  INVX1 U258 ( .A(1'b1), .Y(y8[14]) );
  INVX1 U260 ( .A(1'b1), .Y(y8[15]) );
  INVX1 U262 ( .A(n327), .Y(n325) );
  INVX1 U263 ( .A(n332), .Y(n329) );
  INVX1 U264 ( .A(n332), .Y(n330) );
  INVX1 U265 ( .A(n327), .Y(n326) );
  INVX1 U266 ( .A(n332), .Y(n331) );
  INVX1 U267 ( .A(n3), .Y(idct_ready) );
  INVX1 U268 ( .A(n6), .Y(n327) );
  INVX1 U269 ( .A(n332), .Y(n328) );
  INVX1 U270 ( .A(n4), .Y(n332) );
  INVX1 U271 ( .A(n65), .Y(y0[13]) );
  AOI22X1 U272 ( .A0(y0_idct8[13]), .A1(n328), .B0(y0_idct4[13]), .B1(n325), 
        .Y(n65) );
  INVX1 U273 ( .A(n64), .Y(y0[14]) );
  AOI22X1 U274 ( .A0(y0_idct8[14]), .A1(n328), .B0(y0_idct4[14]), .B1(n325), 
        .Y(n64) );
  INVX1 U275 ( .A(n49), .Y(y1[13]) );
  AOI22X1 U276 ( .A0(y1_idct8[13]), .A1(n329), .B0(y1_idct4[13]), .B1(n326), 
        .Y(n49) );
  INVX1 U277 ( .A(n48), .Y(y1[14]) );
  AOI22X1 U278 ( .A0(y1_idct8[14]), .A1(n330), .B0(y1_idct4[14]), .B1(n326), 
        .Y(n48) );
  INVX1 U279 ( .A(n33), .Y(y2[13]) );
  AOI22X1 U280 ( .A0(y2_idct8[13]), .A1(n329), .B0(y2_idct4[13]), .B1(n326), 
        .Y(n33) );
  INVX1 U281 ( .A(n32), .Y(y2[14]) );
  AOI22X1 U282 ( .A0(y2_idct8[14]), .A1(n330), .B0(y2_idct4[14]), .B1(n326), 
        .Y(n32) );
  INVX1 U283 ( .A(n17), .Y(y3[13]) );
  AOI22X1 U284 ( .A0(y3_idct8[13]), .A1(n330), .B0(y3_idct4[13]), .B1(n326), 
        .Y(n17) );
  INVX1 U285 ( .A(n16), .Y(y3[14]) );
  AOI22X1 U286 ( .A0(y3_idct8[14]), .A1(n330), .B0(y3_idct4[14]), .B1(n6), .Y(
        n16) );
  INVX1 U287 ( .A(n63), .Y(y0[15]) );
  AOI22X1 U288 ( .A0(y0_idct8[15]), .A1(n328), .B0(y0_idct4[15]), .B1(n325), 
        .Y(n63) );
  INVX1 U289 ( .A(n47), .Y(y1[15]) );
  AOI22X1 U290 ( .A0(y1_idct8[15]), .A1(n329), .B0(y1_idct4[15]), .B1(n326), 
        .Y(n47) );
  INVX1 U291 ( .A(n31), .Y(y2[15]) );
  AOI22X1 U292 ( .A0(y2_idct8[15]), .A1(n329), .B0(y2_idct4[15]), .B1(n326), 
        .Y(n31) );
  INVX1 U293 ( .A(n15), .Y(y3[15]) );
  AOI22X1 U294 ( .A0(y3_idct8[15]), .A1(n330), .B0(y3_idct4[15]), .B1(n326), 
        .Y(n15) );
  AOI22X1 U295 ( .A0(idct8_ready), .A1(n328), .B0(idct4_ready), .B1(n325), .Y(
        n3) );
  INVX1 U296 ( .A(n55), .Y(y0[8]) );
  AOI22X1 U297 ( .A0(y0_idct8[8]), .A1(n330), .B0(y0_idct4[8]), .B1(n326), .Y(
        n55) );
  INVX1 U298 ( .A(n54), .Y(y0[9]) );
  AOI22X1 U299 ( .A0(y0_idct8[9]), .A1(n329), .B0(y0_idct4[9]), .B1(n326), .Y(
        n54) );
  INVX1 U300 ( .A(n68), .Y(y0[10]) );
  AOI22X1 U301 ( .A0(y0_idct8[10]), .A1(n328), .B0(y0_idct4[10]), .B1(n325), 
        .Y(n68) );
  INVX1 U302 ( .A(n67), .Y(y0[11]) );
  AOI22X1 U303 ( .A0(y0_idct8[11]), .A1(n328), .B0(y0_idct4[11]), .B1(n325), 
        .Y(n67) );
  INVX1 U304 ( .A(n39), .Y(y1[8]) );
  AOI22X1 U305 ( .A0(y1_idct8[8]), .A1(n330), .B0(y1_idct4[8]), .B1(n6), .Y(
        n39) );
  INVX1 U306 ( .A(n38), .Y(y1[9]) );
  AOI22X1 U307 ( .A0(y1_idct8[9]), .A1(n330), .B0(y1_idct4[9]), .B1(n6), .Y(
        n38) );
  INVX1 U308 ( .A(n52), .Y(y1[10]) );
  AOI22X1 U309 ( .A0(y1_idct8[10]), .A1(n330), .B0(y1_idct4[10]), .B1(n326), 
        .Y(n52) );
  INVX1 U310 ( .A(n51), .Y(y1[11]) );
  AOI22X1 U311 ( .A0(y1_idct8[11]), .A1(n329), .B0(y1_idct4[11]), .B1(n326), 
        .Y(n51) );
  INVX1 U312 ( .A(n23), .Y(y2[8]) );
  AOI22X1 U313 ( .A0(y2_idct8[8]), .A1(n329), .B0(y2_idct4[8]), .B1(n326), .Y(
        n23) );
  INVX1 U314 ( .A(n22), .Y(y2[9]) );
  AOI22X1 U315 ( .A0(y2_idct8[9]), .A1(n329), .B0(y2_idct4[9]), .B1(n326), .Y(
        n22) );
  INVX1 U316 ( .A(n36), .Y(y2[10]) );
  AOI22X1 U317 ( .A0(y2_idct8[10]), .A1(n329), .B0(y2_idct4[10]), .B1(n6), .Y(
        n36) );
  INVX1 U318 ( .A(n35), .Y(y2[11]) );
  AOI22X1 U319 ( .A0(y2_idct8[11]), .A1(n329), .B0(y2_idct4[11]), .B1(n6), .Y(
        n35) );
  INVX1 U320 ( .A(n20), .Y(y3[10]) );
  AOI22X1 U321 ( .A0(y3_idct8[10]), .A1(n329), .B0(y3_idct4[10]), .B1(n326), 
        .Y(n20) );
  INVX1 U322 ( .A(n19), .Y(y3[11]) );
  AOI22X1 U323 ( .A0(y3_idct8[11]), .A1(n329), .B0(y3_idct4[11]), .B1(n6), .Y(
        n19) );
  AND2X2 U324 ( .A(y7_idct8[13]), .B(n4), .Y(y7[13]) );
  INVX1 U325 ( .A(n7), .Y(y3[8]) );
  AOI22X1 U326 ( .A0(y3_idct8[8]), .A1(n330), .B0(y3_idct4[8]), .B1(n6), .Y(n7) );
  INVX1 U327 ( .A(n5), .Y(y3[9]) );
  AOI22X1 U328 ( .A0(y3_idct8[9]), .A1(n330), .B0(y3_idct4[9]), .B1(n6), .Y(n5) );
  NOR2BX1 U329 ( .AN(mode_delay2[0]), .B(mode_delay2[1]), .Y(n4) );
  AND2X2 U330 ( .A(y4_idct8[14]), .B(n331), .Y(y4[14]) );
  AND2X2 U331 ( .A(y4_idct8[15]), .B(n331), .Y(y4[15]) );
  AND2X2 U332 ( .A(y5_idct8[14]), .B(n331), .Y(y5[14]) );
  AND2X2 U333 ( .A(y5_idct8[15]), .B(n331), .Y(y5[15]) );
  AND2X2 U334 ( .A(y6_idct8[14]), .B(n330), .Y(y6[14]) );
  AND2X2 U335 ( .A(y6_idct8[15]), .B(n329), .Y(y6[15]) );
  NOR2X1 U336 ( .A(mode_delay2[0]), .B(mode_delay2[1]), .Y(n6) );
  AND2X2 U337 ( .A(y7_idct8[14]), .B(n4), .Y(y7[14]) );
  AND2X2 U338 ( .A(y7_idct8[15]), .B(n4), .Y(y7[15]) );
  INVX1 U339 ( .A(n66), .Y(y0[12]) );
  AOI22X1 U340 ( .A0(y0_idct8[12]), .A1(n328), .B0(y0_idct4[12]), .B1(n325), 
        .Y(n66) );
  INVX1 U341 ( .A(n50), .Y(y1[12]) );
  AOI22X1 U342 ( .A0(y1_idct8[12]), .A1(n330), .B0(y1_idct4[12]), .B1(n326), 
        .Y(n50) );
  INVX1 U343 ( .A(n34), .Y(y2[12]) );
  AOI22X1 U344 ( .A0(y2_idct8[12]), .A1(n330), .B0(y2_idct4[12]), .B1(n326), 
        .Y(n34) );
  INVX1 U345 ( .A(n18), .Y(y3[12]) );
  AOI22X1 U346 ( .A0(y3_idct8[12]), .A1(n330), .B0(y3_idct4[12]), .B1(n6), .Y(
        n18) );
  AND2X2 U347 ( .A(y4_idct8[13]), .B(n331), .Y(y4[13]) );
  AND2X2 U348 ( .A(y5_idct8[13]), .B(n331), .Y(y5[13]) );
  AND2X2 U349 ( .A(y6_idct8[13]), .B(n330), .Y(y6[13]) );
  INVX1 U350 ( .A(n69), .Y(y0[0]) );
  AOI22X1 U351 ( .A0(y0_idct8[0]), .A1(n328), .B0(y0_idct4[0]), .B1(n325), .Y(
        n69) );
  INVX1 U352 ( .A(n59), .Y(y0[4]) );
  AOI22X1 U353 ( .A0(y0_idct8[4]), .A1(n328), .B0(y0_idct4[4]), .B1(n325), .Y(
        n59) );
  INVX1 U354 ( .A(n57), .Y(y0[6]) );
  AOI22X1 U355 ( .A0(y0_idct8[6]), .A1(n330), .B0(y0_idct4[6]), .B1(n326), .Y(
        n57) );
  INVX1 U356 ( .A(n43), .Y(y1[4]) );
  AOI22X1 U357 ( .A0(y1_idct8[4]), .A1(n329), .B0(y1_idct4[4]), .B1(n6), .Y(
        n43) );
  INVX1 U358 ( .A(n41), .Y(y1[6]) );
  AOI22X1 U359 ( .A0(y1_idct8[6]), .A1(n330), .B0(y1_idct4[6]), .B1(n6), .Y(
        n41) );
  INVX1 U360 ( .A(n27), .Y(y2[4]) );
  AOI22X1 U361 ( .A0(y2_idct8[4]), .A1(n329), .B0(y2_idct4[4]), .B1(n326), .Y(
        n27) );
  INVX1 U362 ( .A(n25), .Y(y2[6]) );
  AOI22X1 U363 ( .A0(y2_idct8[6]), .A1(n329), .B0(y2_idct4[6]), .B1(n326), .Y(
        n25) );
  INVX1 U364 ( .A(n11), .Y(y3[4]) );
  AOI22X1 U365 ( .A0(y3_idct8[4]), .A1(n330), .B0(y3_idct4[4]), .B1(n326), .Y(
        n11) );
  INVX1 U366 ( .A(n10), .Y(y3[5]) );
  AOI22X1 U367 ( .A0(y3_idct8[5]), .A1(n330), .B0(y3_idct4[5]), .B1(n326), .Y(
        n10) );
  INVX1 U368 ( .A(n9), .Y(y3[6]) );
  AOI22X1 U369 ( .A0(y3_idct8[6]), .A1(n330), .B0(y3_idct4[6]), .B1(n6), .Y(n9) );
  INVX1 U370 ( .A(n8), .Y(y3[7]) );
  AOI22X1 U371 ( .A0(y3_idct8[7]), .A1(n330), .B0(y3_idct4[7]), .B1(n326), .Y(
        n8) );
  INVX1 U372 ( .A(n58), .Y(y0[5]) );
  AOI22X1 U373 ( .A0(y0_idct8[5]), .A1(n328), .B0(y0_idct4[5]), .B1(n326), .Y(
        n58) );
  INVX1 U374 ( .A(n56), .Y(y0[7]) );
  AOI22X1 U375 ( .A0(y0_idct8[7]), .A1(n329), .B0(y0_idct4[7]), .B1(n326), .Y(
        n56) );
  INVX1 U376 ( .A(n42), .Y(y1[5]) );
  AOI22X1 U377 ( .A0(y1_idct8[5]), .A1(n330), .B0(y1_idct4[5]), .B1(n6), .Y(
        n42) );
  INVX1 U378 ( .A(n40), .Y(y1[7]) );
  AOI22X1 U379 ( .A0(y1_idct8[7]), .A1(n329), .B0(y1_idct4[7]), .B1(n6), .Y(
        n40) );
  INVX1 U380 ( .A(n26), .Y(y2[5]) );
  AOI22X1 U381 ( .A0(y2_idct8[5]), .A1(n329), .B0(y2_idct4[5]), .B1(n326), .Y(
        n26) );
  INVX1 U382 ( .A(n24), .Y(y2[7]) );
  AOI22X1 U383 ( .A0(y2_idct8[7]), .A1(n329), .B0(y2_idct4[7]), .B1(n326), .Y(
        n24) );
  INVX1 U384 ( .A(n14), .Y(y3[1]) );
  AOI22X1 U385 ( .A0(y3_idct8[1]), .A1(n330), .B0(y3_idct4[1]), .B1(n6), .Y(
        n14) );
  AND2X2 U386 ( .A(y4_idct8[4]), .B(n331), .Y(y4[4]) );
  AND2X2 U387 ( .A(y4_idct8[5]), .B(n331), .Y(y4[5]) );
  AND2X2 U388 ( .A(y4_idct8[6]), .B(n331), .Y(y4[6]) );
  AND2X2 U389 ( .A(y4_idct8[7]), .B(n331), .Y(y4[7]) );
  AND2X2 U390 ( .A(y4_idct8[8]), .B(n331), .Y(y4[8]) );
  AND2X2 U391 ( .A(y4_idct8[9]), .B(n331), .Y(y4[9]) );
  AND2X2 U392 ( .A(y4_idct8[10]), .B(n331), .Y(y4[10]) );
  AND2X2 U393 ( .A(y4_idct8[11]), .B(n331), .Y(y4[11]) );
  AND2X2 U394 ( .A(y4_idct8[12]), .B(n331), .Y(y4[12]) );
  AND2X2 U395 ( .A(y5_idct8[0]), .B(n331), .Y(y5[0]) );
  AND2X2 U396 ( .A(y5_idct8[1]), .B(n331), .Y(y5[1]) );
  AND2X2 U397 ( .A(y5_idct8[2]), .B(n331), .Y(y5[2]) );
  AND2X2 U398 ( .A(y5_idct8[3]), .B(n331), .Y(y5[3]) );
  AND2X2 U399 ( .A(y5_idct8[4]), .B(n331), .Y(y5[4]) );
  AND2X2 U400 ( .A(y5_idct8[5]), .B(n331), .Y(y5[5]) );
  AND2X2 U401 ( .A(y5_idct8[6]), .B(n331), .Y(y5[6]) );
  AND2X2 U402 ( .A(y5_idct8[7]), .B(n331), .Y(y5[7]) );
  AND2X2 U403 ( .A(y5_idct8[8]), .B(n331), .Y(y5[8]) );
  AND2X2 U404 ( .A(y5_idct8[9]), .B(n331), .Y(y5[9]) );
  AND2X2 U405 ( .A(y5_idct8[10]), .B(n331), .Y(y5[10]) );
  AND2X2 U406 ( .A(y5_idct8[11]), .B(n331), .Y(y5[11]) );
  AND2X2 U407 ( .A(y5_idct8[12]), .B(n331), .Y(y5[12]) );
  AND2X2 U408 ( .A(y6_idct8[0]), .B(n330), .Y(y6[0]) );
  AND2X2 U409 ( .A(y6_idct8[1]), .B(n329), .Y(y6[1]) );
  AND2X2 U410 ( .A(y6_idct8[2]), .B(n329), .Y(y6[2]) );
  AND2X2 U411 ( .A(y6_idct8[3]), .B(n330), .Y(y6[3]) );
  AND2X2 U412 ( .A(y6_idct8[4]), .B(n330), .Y(y6[4]) );
  AND2X2 U413 ( .A(y6_idct8[5]), .B(n329), .Y(y6[5]) );
  AND2X2 U414 ( .A(y6_idct8[6]), .B(n328), .Y(y6[6]) );
  AND2X2 U415 ( .A(y6_idct8[7]), .B(n4), .Y(y6[7]) );
  AND2X2 U416 ( .A(y6_idct8[8]), .B(n329), .Y(y6[8]) );
  AND2X2 U417 ( .A(y6_idct8[9]), .B(n4), .Y(y6[9]) );
  AND2X2 U418 ( .A(y6_idct8[10]), .B(n329), .Y(y6[10]) );
  AND2X2 U419 ( .A(y6_idct8[11]), .B(n4), .Y(y6[11]) );
  AND2X2 U420 ( .A(y6_idct8[12]), .B(n330), .Y(y6[12]) );
  AND2X2 U421 ( .A(y4_idct8[0]), .B(n331), .Y(y4[0]) );
  AND2X2 U422 ( .A(y4_idct8[1]), .B(n331), .Y(y4[1]) );
  AND2X2 U423 ( .A(y4_idct8[2]), .B(n331), .Y(y4[2]) );
  AND2X2 U424 ( .A(y4_idct8[3]), .B(n331), .Y(y4[3]) );
  INVX1 U425 ( .A(n62), .Y(y0[1]) );
  AOI22X1 U426 ( .A0(y0_idct8[1]), .A1(n328), .B0(y0_idct4[1]), .B1(n325), .Y(
        n62) );
  INVX1 U427 ( .A(n61), .Y(y0[2]) );
  AOI22X1 U428 ( .A0(y0_idct8[2]), .A1(n328), .B0(y0_idct4[2]), .B1(n325), .Y(
        n61) );
  INVX1 U429 ( .A(n60), .Y(y0[3]) );
  AOI22X1 U430 ( .A0(y0_idct8[3]), .A1(n328), .B0(y0_idct4[3]), .B1(n325), .Y(
        n60) );
  INVX1 U431 ( .A(n53), .Y(y1[0]) );
  AOI22X1 U432 ( .A0(y1_idct8[0]), .A1(n329), .B0(y1_idct4[0]), .B1(n326), .Y(
        n53) );
  INVX1 U433 ( .A(n46), .Y(y1[1]) );
  AOI22X1 U434 ( .A0(y1_idct8[1]), .A1(n330), .B0(y1_idct4[1]), .B1(n6), .Y(
        n46) );
  INVX1 U435 ( .A(n45), .Y(y1[2]) );
  AOI22X1 U436 ( .A0(y1_idct8[2]), .A1(n329), .B0(y1_idct4[2]), .B1(n6), .Y(
        n45) );
  INVX1 U437 ( .A(n44), .Y(y1[3]) );
  AOI22X1 U438 ( .A0(y1_idct8[3]), .A1(n329), .B0(y1_idct4[3]), .B1(n6), .Y(
        n44) );
  INVX1 U439 ( .A(n37), .Y(y2[0]) );
  AOI22X1 U440 ( .A0(y2_idct8[0]), .A1(n330), .B0(y2_idct4[0]), .B1(n6), .Y(
        n37) );
  INVX1 U441 ( .A(n30), .Y(y2[1]) );
  AOI22X1 U442 ( .A0(y2_idct8[1]), .A1(n329), .B0(y2_idct4[1]), .B1(n326), .Y(
        n30) );
  INVX1 U443 ( .A(n29), .Y(y2[2]) );
  AOI22X1 U444 ( .A0(y2_idct8[2]), .A1(n329), .B0(y2_idct4[2]), .B1(n326), .Y(
        n29) );
  INVX1 U445 ( .A(n28), .Y(y2[3]) );
  AOI22X1 U446 ( .A0(y2_idct8[3]), .A1(n329), .B0(y2_idct4[3]), .B1(n325), .Y(
        n28) );
  INVX1 U447 ( .A(n21), .Y(y3[0]) );
  AOI22X1 U448 ( .A0(y3_idct8[0]), .A1(n329), .B0(y3_idct4[0]), .B1(n326), .Y(
        n21) );
  INVX1 U449 ( .A(n13), .Y(y3[2]) );
  AOI22X1 U450 ( .A0(y3_idct8[2]), .A1(n330), .B0(y3_idct4[2]), .B1(n326), .Y(
        n13) );
  INVX1 U451 ( .A(n12), .Y(y3[3]) );
  AOI22X1 U452 ( .A0(y3_idct8[3]), .A1(n330), .B0(y3_idct4[3]), .B1(n6), .Y(
        n12) );
  AND2X2 U453 ( .A(y7_idct8[0]), .B(n4), .Y(y7[0]) );
  AND2X2 U454 ( .A(y7_idct8[1]), .B(n4), .Y(y7[1]) );
  AND2X2 U455 ( .A(y7_idct8[2]), .B(n4), .Y(y7[2]) );
  AND2X2 U456 ( .A(y7_idct8[3]), .B(n4), .Y(y7[3]) );
  AND2X2 U457 ( .A(y7_idct8[4]), .B(n4), .Y(y7[4]) );
  AND2X2 U458 ( .A(y7_idct8[5]), .B(n4), .Y(y7[5]) );
  AND2X2 U459 ( .A(y7_idct8[6]), .B(n4), .Y(y7[6]) );
  AND2X2 U460 ( .A(y7_idct8[7]), .B(n4), .Y(y7[7]) );
  AND2X2 U461 ( .A(y7_idct8[8]), .B(n4), .Y(y7[8]) );
  AND2X2 U462 ( .A(y7_idct8[9]), .B(n4), .Y(y7[9]) );
  AND2X2 U463 ( .A(y7_idct8[10]), .B(n4), .Y(y7[10]) );
  AND2X2 U464 ( .A(y7_idct8[11]), .B(n4), .Y(y7[11]) );
  AND2X2 U465 ( .A(y7_idct8[12]), .B(n4), .Y(y7[12]) );
endmodule


module p2s_0 ( clk, rstn, start, mode, cal_result, dout, p2s_ready, mode_out
 );
  input [1:0] mode;
  input [127:0] cal_result;
  output [15:0] dout;
  output [1:0] mode_out;
  input clk, rstn, start;
  output p2s_ready;
  wire   ready8, mode_reg_0_, shift4_flag, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n215, n221,
         n286, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n308, n309,
         n310, n311, n312, n313, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n209, n210,
         n211, n212, n213, n214, n216, n217, n218, n219, n220, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n287, n307, n314, n447,
         n448, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745;
  wire   [5:0] start_reg4;
  wire   [143:0] result_reg4;
  wire   [127:0] result_reg8;

  AND2X4 U4 ( .A(mode_out[1]), .B(n286), .Y(mode_out[1]) );
  OAI2BB1X4 U5 ( .A0N(n680), .A1N(mode_out[0]), .B0(n674), .Y(mode_out[0]) );
  DFFRHQX1 result_reg8_reg_111_ ( .D(n533), .CK(clk), .RN(rstn), .Q(
        result_reg8[111]) );
  DFFRHQX1 result_reg8_reg_110_ ( .D(n534), .CK(clk), .RN(rstn), .Q(
        result_reg8[110]) );
  DFFRHQX1 result_reg8_reg_109_ ( .D(n535), .CK(clk), .RN(rstn), .Q(
        result_reg8[109]) );
  DFFRHQX1 result_reg8_reg_108_ ( .D(n536), .CK(clk), .RN(rstn), .Q(
        result_reg8[108]) );
  DFFRHQX1 result_reg8_reg_107_ ( .D(n537), .CK(clk), .RN(rstn), .Q(
        result_reg8[107]) );
  DFFRHQX1 result_reg8_reg_106_ ( .D(n538), .CK(clk), .RN(rstn), .Q(
        result_reg8[106]) );
  DFFRHQX1 result_reg8_reg_105_ ( .D(n539), .CK(clk), .RN(rstn), .Q(
        result_reg8[105]) );
  DFFRHQX1 result_reg8_reg_104_ ( .D(n540), .CK(clk), .RN(rstn), .Q(
        result_reg8[104]) );
  DFFRHQX1 result_reg8_reg_103_ ( .D(n541), .CK(clk), .RN(rstn), .Q(
        result_reg8[103]) );
  DFFRHQX1 result_reg8_reg_102_ ( .D(n542), .CK(clk), .RN(rstn), .Q(
        result_reg8[102]) );
  DFFRHQX1 result_reg8_reg_101_ ( .D(n543), .CK(clk), .RN(rstn), .Q(
        result_reg8[101]) );
  DFFRHQX1 result_reg8_reg_100_ ( .D(n544), .CK(clk), .RN(rstn), .Q(
        result_reg8[100]) );
  DFFRHQX1 result_reg8_reg_99_ ( .D(n545), .CK(clk), .RN(rstn), .Q(
        result_reg8[99]) );
  DFFRHQX1 result_reg8_reg_98_ ( .D(n546), .CK(clk), .RN(rstn), .Q(
        result_reg8[98]) );
  DFFRHQX1 result_reg8_reg_97_ ( .D(n547), .CK(clk), .RN(rstn), .Q(
        result_reg8[97]) );
  DFFRHQX1 result_reg8_reg_96_ ( .D(n548), .CK(clk), .RN(rstn), .Q(
        result_reg8[96]) );
  DFFRHQX1 result_reg8_reg_95_ ( .D(n549), .CK(clk), .RN(rstn), .Q(
        result_reg8[95]) );
  DFFRHQX1 result_reg8_reg_94_ ( .D(n550), .CK(clk), .RN(rstn), .Q(
        result_reg8[94]) );
  DFFRHQX1 result_reg8_reg_93_ ( .D(n551), .CK(clk), .RN(rstn), .Q(
        result_reg8[93]) );
  DFFRHQX1 result_reg8_reg_92_ ( .D(n552), .CK(clk), .RN(rstn), .Q(
        result_reg8[92]) );
  DFFRHQX1 result_reg8_reg_91_ ( .D(n553), .CK(clk), .RN(rstn), .Q(
        result_reg8[91]) );
  DFFRHQX1 result_reg8_reg_90_ ( .D(n554), .CK(clk), .RN(rstn), .Q(
        result_reg8[90]) );
  DFFRHQX1 result_reg8_reg_89_ ( .D(n555), .CK(clk), .RN(rstn), .Q(
        result_reg8[89]) );
  DFFRHQX1 result_reg8_reg_88_ ( .D(n556), .CK(clk), .RN(rstn), .Q(
        result_reg8[88]) );
  DFFRHQX1 result_reg8_reg_87_ ( .D(n557), .CK(clk), .RN(rstn), .Q(
        result_reg8[87]) );
  DFFRHQX1 result_reg8_reg_86_ ( .D(n558), .CK(clk), .RN(rstn), .Q(
        result_reg8[86]) );
  DFFRHQX1 result_reg8_reg_85_ ( .D(n559), .CK(clk), .RN(rstn), .Q(
        result_reg8[85]) );
  DFFRHQX1 result_reg8_reg_84_ ( .D(n560), .CK(clk), .RN(rstn), .Q(
        result_reg8[84]) );
  DFFRHQX1 result_reg8_reg_83_ ( .D(n561), .CK(clk), .RN(rstn), .Q(
        result_reg8[83]) );
  DFFRHQX1 result_reg8_reg_82_ ( .D(n562), .CK(clk), .RN(rstn), .Q(
        result_reg8[82]) );
  DFFRHQX1 result_reg8_reg_81_ ( .D(n563), .CK(clk), .RN(rstn), .Q(
        result_reg8[81]) );
  DFFRHQX1 result_reg8_reg_80_ ( .D(n564), .CK(clk), .RN(rstn), .Q(
        result_reg8[80]) );
  DFFRHQX1 start_reg4_reg_5_ ( .D(n667), .CK(clk), .RN(rstn), .Q(start_reg4[5]) );
  DFFRHQX1 start_reg4_reg_4_ ( .D(n666), .CK(clk), .RN(rstn), .Q(start_reg4[4]) );
  DFFRHQX1 start_reg4_reg_3_ ( .D(n665), .CK(clk), .RN(rstn), .Q(start_reg4[3]) );
  DFFRHQX1 start_reg4_reg_2_ ( .D(n664), .CK(clk), .RN(rstn), .Q(start_reg4[2]) );
  DFFRHQX1 start_reg4_reg_1_ ( .D(n663), .CK(clk), .RN(rstn), .Q(start_reg4[1]) );
  DFFRHQX1 result_reg4_reg_95_ ( .D(n630), .CK(clk), .RN(rstn), .Q(
        result_reg4[95]) );
  DFFRHQX1 result_reg4_reg_94_ ( .D(n632), .CK(clk), .RN(rstn), .Q(
        result_reg4[94]) );
  DFFRHQX1 result_reg4_reg_93_ ( .D(n634), .CK(clk), .RN(rstn), .Q(
        result_reg4[93]) );
  DFFRHQX1 result_reg4_reg_92_ ( .D(n636), .CK(clk), .RN(rstn), .Q(
        result_reg4[92]) );
  DFFRHQX1 result_reg4_reg_91_ ( .D(n638), .CK(clk), .RN(rstn), .Q(
        result_reg4[91]) );
  DFFRHQX1 result_reg4_reg_90_ ( .D(n640), .CK(clk), .RN(rstn), .Q(
        result_reg4[90]) );
  DFFRHQX1 result_reg4_reg_89_ ( .D(n642), .CK(clk), .RN(rstn), .Q(
        result_reg4[89]) );
  DFFRHQX1 result_reg4_reg_88_ ( .D(n644), .CK(clk), .RN(rstn), .Q(
        result_reg4[88]) );
  DFFRHQX1 result_reg4_reg_87_ ( .D(n646), .CK(clk), .RN(rstn), .Q(
        result_reg4[87]) );
  DFFRHQX1 result_reg4_reg_86_ ( .D(n648), .CK(clk), .RN(rstn), .Q(
        result_reg4[86]) );
  DFFRHQX1 result_reg4_reg_85_ ( .D(n650), .CK(clk), .RN(rstn), .Q(
        result_reg4[85]) );
  DFFRHQX1 result_reg4_reg_84_ ( .D(n652), .CK(clk), .RN(rstn), .Q(
        result_reg4[84]) );
  DFFRHQX1 result_reg4_reg_83_ ( .D(n654), .CK(clk), .RN(rstn), .Q(
        result_reg4[83]) );
  DFFRHQX1 result_reg4_reg_82_ ( .D(n656), .CK(clk), .RN(rstn), .Q(
        result_reg4[82]) );
  DFFRHQX1 result_reg4_reg_81_ ( .D(n658), .CK(clk), .RN(rstn), .Q(
        result_reg4[81]) );
  DFFRHQX1 result_reg4_reg_80_ ( .D(n660), .CK(clk), .RN(rstn), .Q(
        result_reg4[80]) );
  DFFRHQX1 result_reg4_reg_79_ ( .D(n629), .CK(clk), .RN(rstn), .Q(
        result_reg4[79]) );
  DFFRHQX1 result_reg4_reg_78_ ( .D(n631), .CK(clk), .RN(rstn), .Q(
        result_reg4[78]) );
  DFFRHQX1 result_reg4_reg_77_ ( .D(n633), .CK(clk), .RN(rstn), .Q(
        result_reg4[77]) );
  DFFRHQX1 result_reg4_reg_76_ ( .D(n635), .CK(clk), .RN(rstn), .Q(
        result_reg4[76]) );
  DFFRHQX1 result_reg4_reg_75_ ( .D(n637), .CK(clk), .RN(rstn), .Q(
        result_reg4[75]) );
  DFFRHQX1 result_reg4_reg_74_ ( .D(n639), .CK(clk), .RN(rstn), .Q(
        result_reg4[74]) );
  DFFRHQX1 result_reg4_reg_73_ ( .D(n641), .CK(clk), .RN(rstn), .Q(
        result_reg4[73]) );
  DFFRHQX1 result_reg4_reg_72_ ( .D(n643), .CK(clk), .RN(rstn), .Q(
        result_reg4[72]) );
  DFFRHQX1 result_reg4_reg_71_ ( .D(n645), .CK(clk), .RN(rstn), .Q(
        result_reg4[71]) );
  DFFRHQX1 result_reg4_reg_70_ ( .D(n647), .CK(clk), .RN(rstn), .Q(
        result_reg4[70]) );
  DFFRHQX1 result_reg4_reg_69_ ( .D(n649), .CK(clk), .RN(rstn), .Q(
        result_reg4[69]) );
  DFFRHQX1 result_reg4_reg_68_ ( .D(n651), .CK(clk), .RN(rstn), .Q(
        result_reg4[68]) );
  DFFRHQX1 result_reg4_reg_67_ ( .D(n653), .CK(clk), .RN(rstn), .Q(
        result_reg4[67]) );
  DFFRHQX1 result_reg4_reg_66_ ( .D(n655), .CK(clk), .RN(rstn), .Q(
        result_reg4[66]) );
  DFFRHQX1 result_reg4_reg_65_ ( .D(n657), .CK(clk), .RN(rstn), .Q(
        result_reg4[65]) );
  DFFRHQX1 result_reg4_reg_64_ ( .D(n659), .CK(clk), .RN(rstn), .Q(
        result_reg4[64]) );
  DFFRHQX1 result_reg8_reg_63_ ( .D(n17), .CK(clk), .RN(rstn), .Q(
        result_reg8[63]) );
  DFFRHQX1 result_reg8_reg_62_ ( .D(n18), .CK(clk), .RN(rstn), .Q(
        result_reg8[62]) );
  DFFRHQX1 result_reg8_reg_61_ ( .D(n19), .CK(clk), .RN(rstn), .Q(
        result_reg8[61]) );
  DFFRHQX1 result_reg8_reg_60_ ( .D(n20), .CK(clk), .RN(rstn), .Q(
        result_reg8[60]) );
  DFFRHQX1 result_reg8_reg_59_ ( .D(n21), .CK(clk), .RN(rstn), .Q(
        result_reg8[59]) );
  DFFRHQX1 result_reg8_reg_58_ ( .D(n22), .CK(clk), .RN(rstn), .Q(
        result_reg8[58]) );
  DFFRHQX1 result_reg8_reg_57_ ( .D(n23), .CK(clk), .RN(rstn), .Q(
        result_reg8[57]) );
  DFFRHQX1 result_reg8_reg_56_ ( .D(n24), .CK(clk), .RN(rstn), .Q(
        result_reg8[56]) );
  DFFRHQX1 result_reg8_reg_55_ ( .D(n25), .CK(clk), .RN(rstn), .Q(
        result_reg8[55]) );
  DFFRHQX1 result_reg8_reg_54_ ( .D(n26), .CK(clk), .RN(rstn), .Q(
        result_reg8[54]) );
  DFFRHQX1 result_reg8_reg_53_ ( .D(n27), .CK(clk), .RN(rstn), .Q(
        result_reg8[53]) );
  DFFRHQX1 result_reg8_reg_52_ ( .D(n28), .CK(clk), .RN(rstn), .Q(
        result_reg8[52]) );
  DFFRHQX1 result_reg8_reg_51_ ( .D(n29), .CK(clk), .RN(rstn), .Q(
        result_reg8[51]) );
  DFFRHQX1 result_reg8_reg_50_ ( .D(n30), .CK(clk), .RN(rstn), .Q(
        result_reg8[50]) );
  DFFRHQX1 result_reg8_reg_49_ ( .D(n31), .CK(clk), .RN(rstn), .Q(
        result_reg8[49]) );
  DFFRHQX1 result_reg8_reg_48_ ( .D(n32), .CK(clk), .RN(rstn), .Q(
        result_reg8[48]) );
  DFFRHQX1 result_reg8_reg_47_ ( .D(n33), .CK(clk), .RN(rstn), .Q(
        result_reg8[47]) );
  DFFRHQX1 result_reg8_reg_46_ ( .D(n34), .CK(clk), .RN(rstn), .Q(
        result_reg8[46]) );
  DFFRHQX1 result_reg8_reg_45_ ( .D(n35), .CK(clk), .RN(rstn), .Q(
        result_reg8[45]) );
  DFFRHQX1 result_reg8_reg_44_ ( .D(n36), .CK(clk), .RN(rstn), .Q(
        result_reg8[44]) );
  DFFRHQX1 result_reg8_reg_43_ ( .D(n37), .CK(clk), .RN(rstn), .Q(
        result_reg8[43]) );
  DFFRHQX1 result_reg8_reg_42_ ( .D(n38), .CK(clk), .RN(rstn), .Q(
        result_reg8[42]) );
  DFFRHQX1 result_reg8_reg_41_ ( .D(n39), .CK(clk), .RN(rstn), .Q(
        result_reg8[41]) );
  DFFRHQX1 result_reg8_reg_40_ ( .D(n40), .CK(clk), .RN(rstn), .Q(
        result_reg8[40]) );
  DFFRHQX1 result_reg8_reg_39_ ( .D(n41), .CK(clk), .RN(rstn), .Q(
        result_reg8[39]) );
  DFFRHQX1 result_reg8_reg_38_ ( .D(n42), .CK(clk), .RN(rstn), .Q(
        result_reg8[38]) );
  DFFRHQX1 result_reg8_reg_37_ ( .D(n43), .CK(clk), .RN(rstn), .Q(
        result_reg8[37]) );
  DFFRHQX1 result_reg8_reg_36_ ( .D(n44), .CK(clk), .RN(rstn), .Q(
        result_reg8[36]) );
  DFFRHQX1 result_reg8_reg_35_ ( .D(n45), .CK(clk), .RN(rstn), .Q(
        result_reg8[35]) );
  DFFRHQX1 result_reg8_reg_34_ ( .D(n46), .CK(clk), .RN(rstn), .Q(
        result_reg8[34]) );
  DFFRHQX1 result_reg8_reg_33_ ( .D(n47), .CK(clk), .RN(rstn), .Q(
        result_reg8[33]) );
  DFFRHQX1 result_reg8_reg_32_ ( .D(n48), .CK(clk), .RN(rstn), .Q(
        result_reg8[32]) );
  DFFRHQX1 result_reg8_reg_31_ ( .D(n49), .CK(clk), .RN(rstn), .Q(
        result_reg8[31]) );
  DFFRHQX1 result_reg8_reg_30_ ( .D(n50), .CK(clk), .RN(rstn), .Q(
        result_reg8[30]) );
  DFFRHQX1 result_reg8_reg_29_ ( .D(n51), .CK(clk), .RN(rstn), .Q(
        result_reg8[29]) );
  DFFRHQX1 result_reg8_reg_28_ ( .D(n52), .CK(clk), .RN(rstn), .Q(
        result_reg8[28]) );
  DFFRHQX1 result_reg8_reg_27_ ( .D(n53), .CK(clk), .RN(rstn), .Q(
        result_reg8[27]) );
  DFFRHQX1 result_reg8_reg_26_ ( .D(n54), .CK(clk), .RN(rstn), .Q(
        result_reg8[26]) );
  DFFRHQX1 result_reg8_reg_25_ ( .D(n55), .CK(clk), .RN(rstn), .Q(
        result_reg8[25]) );
  DFFRHQX1 result_reg8_reg_24_ ( .D(n56), .CK(clk), .RN(rstn), .Q(
        result_reg8[24]) );
  DFFRHQX1 result_reg8_reg_23_ ( .D(n57), .CK(clk), .RN(rstn), .Q(
        result_reg8[23]) );
  DFFRHQX1 result_reg8_reg_22_ ( .D(n58), .CK(clk), .RN(rstn), .Q(
        result_reg8[22]) );
  DFFRHQX1 result_reg8_reg_21_ ( .D(n59), .CK(clk), .RN(rstn), .Q(
        result_reg8[21]) );
  DFFRHQX1 result_reg8_reg_20_ ( .D(n60), .CK(clk), .RN(rstn), .Q(
        result_reg8[20]) );
  DFFRHQX1 result_reg8_reg_19_ ( .D(n61), .CK(clk), .RN(rstn), .Q(
        result_reg8[19]) );
  DFFRHQX1 result_reg8_reg_18_ ( .D(n62), .CK(clk), .RN(rstn), .Q(
        result_reg8[18]) );
  DFFRHQX1 result_reg8_reg_17_ ( .D(n63), .CK(clk), .RN(rstn), .Q(
        result_reg8[17]) );
  DFFRHQX1 result_reg8_reg_16_ ( .D(n64), .CK(clk), .RN(rstn), .Q(
        result_reg8[16]) );
  DFFRHQX1 result_reg8_reg_79_ ( .D(n565), .CK(clk), .RN(rstn), .Q(
        result_reg8[79]) );
  DFFRHQX1 result_reg8_reg_78_ ( .D(n566), .CK(clk), .RN(rstn), .Q(
        result_reg8[78]) );
  DFFRHQX1 result_reg8_reg_77_ ( .D(n567), .CK(clk), .RN(rstn), .Q(
        result_reg8[77]) );
  DFFRHQX1 result_reg8_reg_76_ ( .D(n568), .CK(clk), .RN(rstn), .Q(
        result_reg8[76]) );
  DFFRHQX1 result_reg8_reg_75_ ( .D(n569), .CK(clk), .RN(rstn), .Q(
        result_reg8[75]) );
  DFFRHQX1 result_reg8_reg_74_ ( .D(n570), .CK(clk), .RN(rstn), .Q(
        result_reg8[74]) );
  DFFRHQX1 result_reg8_reg_73_ ( .D(n571), .CK(clk), .RN(rstn), .Q(
        result_reg8[73]) );
  DFFRHQX1 result_reg8_reg_72_ ( .D(n572), .CK(clk), .RN(rstn), .Q(
        result_reg8[72]) );
  DFFRHQX1 result_reg8_reg_71_ ( .D(n573), .CK(clk), .RN(rstn), .Q(
        result_reg8[71]) );
  DFFRHQX1 result_reg8_reg_70_ ( .D(n574), .CK(clk), .RN(rstn), .Q(
        result_reg8[70]) );
  DFFRHQX1 result_reg8_reg_69_ ( .D(n575), .CK(clk), .RN(rstn), .Q(
        result_reg8[69]) );
  DFFRHQX1 result_reg8_reg_68_ ( .D(n576), .CK(clk), .RN(rstn), .Q(
        result_reg8[68]) );
  DFFRHQX1 result_reg8_reg_67_ ( .D(n577), .CK(clk), .RN(rstn), .Q(
        result_reg8[67]) );
  DFFRHQX1 result_reg8_reg_66_ ( .D(n578), .CK(clk), .RN(rstn), .Q(
        result_reg8[66]) );
  DFFRHQX1 result_reg8_reg_65_ ( .D(n579), .CK(clk), .RN(rstn), .Q(
        result_reg8[65]) );
  DFFRHQX1 result_reg8_reg_64_ ( .D(n580), .CK(clk), .RN(rstn), .Q(
        result_reg8[64]) );
  DFFRHQX1 result_reg8_reg_15_ ( .D(n65), .CK(clk), .RN(rstn), .Q(
        result_reg8[15]) );
  DFFRHQX1 result_reg8_reg_14_ ( .D(n66), .CK(clk), .RN(rstn), .Q(
        result_reg8[14]) );
  DFFRHQX1 result_reg8_reg_13_ ( .D(n67), .CK(clk), .RN(rstn), .Q(
        result_reg8[13]) );
  DFFRHQX1 result_reg8_reg_12_ ( .D(n68), .CK(clk), .RN(rstn), .Q(
        result_reg8[12]) );
  DFFRHQX1 result_reg8_reg_11_ ( .D(n69), .CK(clk), .RN(rstn), .Q(
        result_reg8[11]) );
  DFFRHQX1 result_reg8_reg_10_ ( .D(n70), .CK(clk), .RN(rstn), .Q(
        result_reg8[10]) );
  DFFRHQX1 result_reg8_reg_9_ ( .D(n71), .CK(clk), .RN(rstn), .Q(
        result_reg8[9]) );
  DFFRHQX1 result_reg8_reg_8_ ( .D(n72), .CK(clk), .RN(rstn), .Q(
        result_reg8[8]) );
  DFFRHQX1 result_reg8_reg_7_ ( .D(n73), .CK(clk), .RN(rstn), .Q(
        result_reg8[7]) );
  DFFRHQX1 result_reg8_reg_6_ ( .D(n74), .CK(clk), .RN(rstn), .Q(
        result_reg8[6]) );
  DFFRHQX1 result_reg8_reg_5_ ( .D(n75), .CK(clk), .RN(rstn), .Q(
        result_reg8[5]) );
  DFFRHQX1 result_reg8_reg_4_ ( .D(n76), .CK(clk), .RN(rstn), .Q(
        result_reg8[4]) );
  DFFRHQX1 result_reg8_reg_3_ ( .D(n77), .CK(clk), .RN(rstn), .Q(
        result_reg8[3]) );
  DFFRHQX1 result_reg8_reg_2_ ( .D(n78), .CK(clk), .RN(rstn), .Q(
        result_reg8[2]) );
  DFFRHQX1 result_reg8_reg_1_ ( .D(n79), .CK(clk), .RN(rstn), .Q(
        result_reg8[1]) );
  DFFRHQX1 result_reg8_reg_0_ ( .D(n80), .CK(clk), .RN(rstn), .Q(
        result_reg8[0]) );
  DFFRHQX1 result_reg4_reg_143_ ( .D(n581), .CK(clk), .RN(rstn), .Q(
        result_reg4[143]) );
  DFFRHQX1 result_reg4_reg_142_ ( .D(n582), .CK(clk), .RN(rstn), .Q(
        result_reg4[142]) );
  DFFRHQX1 result_reg4_reg_141_ ( .D(n583), .CK(clk), .RN(rstn), .Q(
        result_reg4[141]) );
  DFFRHQX1 result_reg4_reg_140_ ( .D(n584), .CK(clk), .RN(rstn), .Q(
        result_reg4[140]) );
  DFFRHQX1 result_reg4_reg_139_ ( .D(n585), .CK(clk), .RN(rstn), .Q(
        result_reg4[139]) );
  DFFRHQX1 result_reg4_reg_138_ ( .D(n586), .CK(clk), .RN(rstn), .Q(
        result_reg4[138]) );
  DFFRHQX1 result_reg4_reg_137_ ( .D(n587), .CK(clk), .RN(rstn), .Q(
        result_reg4[137]) );
  DFFRHQX1 result_reg4_reg_136_ ( .D(n588), .CK(clk), .RN(rstn), .Q(
        result_reg4[136]) );
  DFFRHQX1 result_reg4_reg_135_ ( .D(n589), .CK(clk), .RN(rstn), .Q(
        result_reg4[135]) );
  DFFRHQX1 result_reg4_reg_134_ ( .D(n590), .CK(clk), .RN(rstn), .Q(
        result_reg4[134]) );
  DFFRHQX1 result_reg4_reg_133_ ( .D(n591), .CK(clk), .RN(rstn), .Q(
        result_reg4[133]) );
  DFFRHQX1 result_reg4_reg_132_ ( .D(n592), .CK(clk), .RN(rstn), .Q(
        result_reg4[132]) );
  DFFRHQX1 result_reg4_reg_131_ ( .D(n593), .CK(clk), .RN(rstn), .Q(
        result_reg4[131]) );
  DFFRHQX1 result_reg4_reg_130_ ( .D(n594), .CK(clk), .RN(rstn), .Q(
        result_reg4[130]) );
  DFFRHQX1 result_reg4_reg_129_ ( .D(n595), .CK(clk), .RN(rstn), .Q(
        result_reg4[129]) );
  DFFRHQX1 result_reg4_reg_128_ ( .D(n596), .CK(clk), .RN(rstn), .Q(
        result_reg4[128]) );
  DFFRHQX1 result_reg4_reg_127_ ( .D(n597), .CK(clk), .RN(rstn), .Q(
        result_reg4[127]) );
  DFFRHQX1 result_reg4_reg_126_ ( .D(n598), .CK(clk), .RN(rstn), .Q(
        result_reg4[126]) );
  DFFRHQX1 result_reg4_reg_125_ ( .D(n599), .CK(clk), .RN(rstn), .Q(
        result_reg4[125]) );
  DFFRHQX1 result_reg4_reg_124_ ( .D(n600), .CK(clk), .RN(rstn), .Q(
        result_reg4[124]) );
  DFFRHQX1 result_reg4_reg_123_ ( .D(n601), .CK(clk), .RN(rstn), .Q(
        result_reg4[123]) );
  DFFRHQX1 result_reg4_reg_122_ ( .D(n602), .CK(clk), .RN(rstn), .Q(
        result_reg4[122]) );
  DFFRHQX1 result_reg4_reg_121_ ( .D(n603), .CK(clk), .RN(rstn), .Q(
        result_reg4[121]) );
  DFFRHQX1 result_reg4_reg_120_ ( .D(n604), .CK(clk), .RN(rstn), .Q(
        result_reg4[120]) );
  DFFRHQX1 result_reg4_reg_119_ ( .D(n605), .CK(clk), .RN(rstn), .Q(
        result_reg4[119]) );
  DFFRHQX1 result_reg4_reg_118_ ( .D(n606), .CK(clk), .RN(rstn), .Q(
        result_reg4[118]) );
  DFFRHQX1 result_reg4_reg_117_ ( .D(n607), .CK(clk), .RN(rstn), .Q(
        result_reg4[117]) );
  DFFRHQX1 result_reg4_reg_116_ ( .D(n608), .CK(clk), .RN(rstn), .Q(
        result_reg4[116]) );
  DFFRHQX1 result_reg4_reg_115_ ( .D(n609), .CK(clk), .RN(rstn), .Q(
        result_reg4[115]) );
  DFFRHQX1 result_reg4_reg_114_ ( .D(n610), .CK(clk), .RN(rstn), .Q(
        result_reg4[114]) );
  DFFRHQX1 result_reg4_reg_113_ ( .D(n611), .CK(clk), .RN(rstn), .Q(
        result_reg4[113]) );
  DFFRHQX1 result_reg4_reg_112_ ( .D(n612), .CK(clk), .RN(rstn), .Q(
        result_reg4[112]) );
  DFFRHQX1 result_reg4_reg_111_ ( .D(n613), .CK(clk), .RN(rstn), .Q(
        result_reg4[111]) );
  DFFRHQX1 result_reg4_reg_110_ ( .D(n614), .CK(clk), .RN(rstn), .Q(
        result_reg4[110]) );
  DFFRHQX1 result_reg4_reg_109_ ( .D(n615), .CK(clk), .RN(rstn), .Q(
        result_reg4[109]) );
  DFFRHQX1 result_reg4_reg_108_ ( .D(n616), .CK(clk), .RN(rstn), .Q(
        result_reg4[108]) );
  DFFRHQX1 result_reg4_reg_107_ ( .D(n617), .CK(clk), .RN(rstn), .Q(
        result_reg4[107]) );
  DFFRHQX1 result_reg4_reg_106_ ( .D(n618), .CK(clk), .RN(rstn), .Q(
        result_reg4[106]) );
  DFFRHQX1 result_reg4_reg_105_ ( .D(n619), .CK(clk), .RN(rstn), .Q(
        result_reg4[105]) );
  DFFRHQX1 result_reg4_reg_104_ ( .D(n620), .CK(clk), .RN(rstn), .Q(
        result_reg4[104]) );
  DFFRHQX1 result_reg4_reg_103_ ( .D(n621), .CK(clk), .RN(rstn), .Q(
        result_reg4[103]) );
  DFFRHQX1 result_reg4_reg_102_ ( .D(n622), .CK(clk), .RN(rstn), .Q(
        result_reg4[102]) );
  DFFRHQX1 result_reg4_reg_101_ ( .D(n623), .CK(clk), .RN(rstn), .Q(
        result_reg4[101]) );
  DFFRHQX1 result_reg4_reg_100_ ( .D(n624), .CK(clk), .RN(rstn), .Q(
        result_reg4[100]) );
  DFFRHQX1 result_reg4_reg_99_ ( .D(n625), .CK(clk), .RN(rstn), .Q(
        result_reg4[99]) );
  DFFRHQX1 result_reg4_reg_98_ ( .D(n626), .CK(clk), .RN(rstn), .Q(
        result_reg4[98]) );
  DFFRHQX1 result_reg4_reg_97_ ( .D(n627), .CK(clk), .RN(rstn), .Q(
        result_reg4[97]) );
  DFFRHQX1 result_reg4_reg_96_ ( .D(n628), .CK(clk), .RN(rstn), .Q(
        result_reg4[96]) );
  DFFRHQX1 result_reg4_reg_15_ ( .D(n193), .CK(clk), .RN(rstn), .Q(
        result_reg4[15]) );
  DFFRHQX1 result_reg4_reg_14_ ( .D(n194), .CK(clk), .RN(rstn), .Q(
        result_reg4[14]) );
  DFFRHQX1 result_reg4_reg_13_ ( .D(n195), .CK(clk), .RN(rstn), .Q(
        result_reg4[13]) );
  DFFRHQX1 result_reg4_reg_12_ ( .D(n196), .CK(clk), .RN(rstn), .Q(
        result_reg4[12]) );
  DFFRHQX1 result_reg4_reg_11_ ( .D(n197), .CK(clk), .RN(rstn), .Q(
        result_reg4[11]) );
  DFFRHQX1 result_reg4_reg_10_ ( .D(n198), .CK(clk), .RN(rstn), .Q(
        result_reg4[10]) );
  DFFRHQX1 result_reg4_reg_9_ ( .D(n199), .CK(clk), .RN(rstn), .Q(
        result_reg4[9]) );
  DFFRHQX1 result_reg4_reg_8_ ( .D(n200), .CK(clk), .RN(rstn), .Q(
        result_reg4[8]) );
  DFFRHQX1 result_reg4_reg_7_ ( .D(n201), .CK(clk), .RN(rstn), .Q(
        result_reg4[7]) );
  DFFRHQX1 result_reg4_reg_6_ ( .D(n202), .CK(clk), .RN(rstn), .Q(
        result_reg4[6]) );
  DFFRHQX1 result_reg4_reg_5_ ( .D(n203), .CK(clk), .RN(rstn), .Q(
        result_reg4[5]) );
  DFFRHQX1 result_reg4_reg_4_ ( .D(n204), .CK(clk), .RN(rstn), .Q(
        result_reg4[4]) );
  DFFRHQX1 result_reg4_reg_3_ ( .D(n205), .CK(clk), .RN(rstn), .Q(
        result_reg4[3]) );
  DFFRHQX1 result_reg4_reg_2_ ( .D(n206), .CK(clk), .RN(rstn), .Q(
        result_reg4[2]) );
  DFFRHQX1 result_reg4_reg_1_ ( .D(n207), .CK(clk), .RN(rstn), .Q(
        result_reg4[1]) );
  DFFRHQX1 result_reg4_reg_0_ ( .D(n208), .CK(clk), .RN(rstn), .Q(
        result_reg4[0]) );
  DFFRHQX1 result_reg4_reg_63_ ( .D(n145), .CK(clk), .RN(rstn), .Q(
        result_reg4[63]) );
  DFFRHQX1 result_reg4_reg_47_ ( .D(n161), .CK(clk), .RN(rstn), .Q(
        result_reg4[47]) );
  DFFRHQX1 result_reg4_reg_31_ ( .D(n177), .CK(clk), .RN(rstn), .Q(
        result_reg4[31]) );
  DFFRHQX1 result_reg4_reg_62_ ( .D(n146), .CK(clk), .RN(rstn), .Q(
        result_reg4[62]) );
  DFFRHQX1 result_reg4_reg_46_ ( .D(n162), .CK(clk), .RN(rstn), .Q(
        result_reg4[46]) );
  DFFRHQX1 result_reg4_reg_30_ ( .D(n178), .CK(clk), .RN(rstn), .Q(
        result_reg4[30]) );
  DFFRHQX1 result_reg4_reg_61_ ( .D(n147), .CK(clk), .RN(rstn), .Q(
        result_reg4[61]) );
  DFFRHQX1 result_reg4_reg_45_ ( .D(n163), .CK(clk), .RN(rstn), .Q(
        result_reg4[45]) );
  DFFRHQX1 result_reg4_reg_29_ ( .D(n179), .CK(clk), .RN(rstn), .Q(
        result_reg4[29]) );
  DFFRHQX1 result_reg4_reg_60_ ( .D(n148), .CK(clk), .RN(rstn), .Q(
        result_reg4[60]) );
  DFFRHQX1 result_reg4_reg_44_ ( .D(n164), .CK(clk), .RN(rstn), .Q(
        result_reg4[44]) );
  DFFRHQX1 result_reg4_reg_28_ ( .D(n180), .CK(clk), .RN(rstn), .Q(
        result_reg4[28]) );
  DFFRHQX1 result_reg4_reg_59_ ( .D(n149), .CK(clk), .RN(rstn), .Q(
        result_reg4[59]) );
  DFFRHQX1 result_reg4_reg_43_ ( .D(n165), .CK(clk), .RN(rstn), .Q(
        result_reg4[43]) );
  DFFRHQX1 result_reg4_reg_27_ ( .D(n181), .CK(clk), .RN(rstn), .Q(
        result_reg4[27]) );
  DFFRHQX1 result_reg4_reg_58_ ( .D(n150), .CK(clk), .RN(rstn), .Q(
        result_reg4[58]) );
  DFFRHQX1 result_reg4_reg_42_ ( .D(n166), .CK(clk), .RN(rstn), .Q(
        result_reg4[42]) );
  DFFRHQX1 result_reg4_reg_26_ ( .D(n182), .CK(clk), .RN(rstn), .Q(
        result_reg4[26]) );
  DFFRHQX1 result_reg4_reg_57_ ( .D(n151), .CK(clk), .RN(rstn), .Q(
        result_reg4[57]) );
  DFFRHQX1 result_reg4_reg_41_ ( .D(n167), .CK(clk), .RN(rstn), .Q(
        result_reg4[41]) );
  DFFRHQX1 result_reg4_reg_25_ ( .D(n183), .CK(clk), .RN(rstn), .Q(
        result_reg4[25]) );
  DFFRHQX1 result_reg4_reg_56_ ( .D(n152), .CK(clk), .RN(rstn), .Q(
        result_reg4[56]) );
  DFFRHQX1 result_reg4_reg_40_ ( .D(n168), .CK(clk), .RN(rstn), .Q(
        result_reg4[40]) );
  DFFRHQX1 result_reg4_reg_24_ ( .D(n184), .CK(clk), .RN(rstn), .Q(
        result_reg4[24]) );
  DFFRHQX1 result_reg4_reg_55_ ( .D(n153), .CK(clk), .RN(rstn), .Q(
        result_reg4[55]) );
  DFFRHQX1 result_reg4_reg_39_ ( .D(n169), .CK(clk), .RN(rstn), .Q(
        result_reg4[39]) );
  DFFRHQX1 result_reg4_reg_23_ ( .D(n185), .CK(clk), .RN(rstn), .Q(
        result_reg4[23]) );
  DFFRHQX1 result_reg4_reg_54_ ( .D(n154), .CK(clk), .RN(rstn), .Q(
        result_reg4[54]) );
  DFFRHQX1 result_reg4_reg_38_ ( .D(n170), .CK(clk), .RN(rstn), .Q(
        result_reg4[38]) );
  DFFRHQX1 result_reg4_reg_22_ ( .D(n186), .CK(clk), .RN(rstn), .Q(
        result_reg4[22]) );
  DFFRHQX1 result_reg4_reg_53_ ( .D(n155), .CK(clk), .RN(rstn), .Q(
        result_reg4[53]) );
  DFFRHQX1 result_reg4_reg_37_ ( .D(n171), .CK(clk), .RN(rstn), .Q(
        result_reg4[37]) );
  DFFRHQX1 result_reg4_reg_21_ ( .D(n187), .CK(clk), .RN(rstn), .Q(
        result_reg4[21]) );
  DFFRHQX1 result_reg4_reg_52_ ( .D(n156), .CK(clk), .RN(rstn), .Q(
        result_reg4[52]) );
  DFFRHQX1 result_reg4_reg_36_ ( .D(n172), .CK(clk), .RN(rstn), .Q(
        result_reg4[36]) );
  DFFRHQX1 result_reg4_reg_20_ ( .D(n188), .CK(clk), .RN(rstn), .Q(
        result_reg4[20]) );
  DFFRHQX1 result_reg4_reg_51_ ( .D(n157), .CK(clk), .RN(rstn), .Q(
        result_reg4[51]) );
  DFFRHQX1 result_reg4_reg_35_ ( .D(n173), .CK(clk), .RN(rstn), .Q(
        result_reg4[35]) );
  DFFRHQX1 result_reg4_reg_19_ ( .D(n189), .CK(clk), .RN(rstn), .Q(
        result_reg4[19]) );
  DFFRHQX1 result_reg4_reg_50_ ( .D(n158), .CK(clk), .RN(rstn), .Q(
        result_reg4[50]) );
  DFFRHQX1 result_reg4_reg_34_ ( .D(n174), .CK(clk), .RN(rstn), .Q(
        result_reg4[34]) );
  DFFRHQX1 result_reg4_reg_18_ ( .D(n190), .CK(clk), .RN(rstn), .Q(
        result_reg4[18]) );
  DFFRHQX1 result_reg4_reg_49_ ( .D(n159), .CK(clk), .RN(rstn), .Q(
        result_reg4[49]) );
  DFFRHQX1 result_reg4_reg_33_ ( .D(n175), .CK(clk), .RN(rstn), .Q(
        result_reg4[33]) );
  DFFRHQX1 result_reg4_reg_17_ ( .D(n191), .CK(clk), .RN(rstn), .Q(
        result_reg4[17]) );
  DFFRHQX1 result_reg4_reg_48_ ( .D(n160), .CK(clk), .RN(rstn), .Q(
        result_reg4[48]) );
  DFFRHQX1 result_reg4_reg_32_ ( .D(n176), .CK(clk), .RN(rstn), .Q(
        result_reg4[32]) );
  DFFRHQX1 result_reg4_reg_16_ ( .D(n192), .CK(clk), .RN(rstn), .Q(
        result_reg4[16]) );
  DFFRHQX1 result_reg8_reg_127_ ( .D(n1), .CK(clk), .RN(rstn), .Q(
        result_reg8[127]) );
  DFFRHQX1 result_reg8_reg_126_ ( .D(n2), .CK(clk), .RN(rstn), .Q(
        result_reg8[126]) );
  DFFRHQX1 result_reg8_reg_125_ ( .D(n3), .CK(clk), .RN(rstn), .Q(
        result_reg8[125]) );
  DFFRHQX1 result_reg8_reg_124_ ( .D(n4), .CK(clk), .RN(rstn), .Q(
        result_reg8[124]) );
  DFFRHQX1 result_reg8_reg_123_ ( .D(n5), .CK(clk), .RN(rstn), .Q(
        result_reg8[123]) );
  DFFRHQX1 result_reg8_reg_122_ ( .D(n6), .CK(clk), .RN(rstn), .Q(
        result_reg8[122]) );
  DFFRHQX1 result_reg8_reg_121_ ( .D(n7), .CK(clk), .RN(rstn), .Q(
        result_reg8[121]) );
  DFFRHQX1 result_reg8_reg_120_ ( .D(n8), .CK(clk), .RN(rstn), .Q(
        result_reg8[120]) );
  DFFRHQX1 result_reg8_reg_119_ ( .D(n9), .CK(clk), .RN(rstn), .Q(
        result_reg8[119]) );
  DFFRHQX1 result_reg8_reg_118_ ( .D(n10), .CK(clk), .RN(rstn), .Q(
        result_reg8[118]) );
  DFFRHQX1 result_reg8_reg_117_ ( .D(n11), .CK(clk), .RN(rstn), .Q(
        result_reg8[117]) );
  DFFRHQX1 result_reg8_reg_116_ ( .D(n12), .CK(clk), .RN(rstn), .Q(
        result_reg8[116]) );
  DFFRHQX1 result_reg8_reg_115_ ( .D(n13), .CK(clk), .RN(rstn), .Q(
        result_reg8[115]) );
  DFFRHQX1 result_reg8_reg_114_ ( .D(n14), .CK(clk), .RN(rstn), .Q(
        result_reg8[114]) );
  DFFRHQX1 result_reg8_reg_113_ ( .D(n15), .CK(clk), .RN(rstn), .Q(
        result_reg8[113]) );
  DFFRHQX1 result_reg8_reg_112_ ( .D(n16), .CK(clk), .RN(rstn), .Q(
        result_reg8[112]) );
  DFFRHQX1 mode_reg_reg_0_ ( .D(n532), .CK(clk), .RN(rstn), .Q(mode_reg_0_) );
  DFFRHQX1 dout_reg_15_ ( .D(n531), .CK(clk), .RN(rstn), .Q(dout[15]) );
  DFFRHQX1 dout_reg_14_ ( .D(n530), .CK(clk), .RN(rstn), .Q(dout[14]) );
  DFFRHQX1 dout_reg_13_ ( .D(n529), .CK(clk), .RN(rstn), .Q(dout[13]) );
  DFFRHQX1 dout_reg_12_ ( .D(n528), .CK(clk), .RN(rstn), .Q(dout[12]) );
  DFFRHQX1 dout_reg_11_ ( .D(n527), .CK(clk), .RN(rstn), .Q(dout[11]) );
  DFFRHQX1 dout_reg_10_ ( .D(n526), .CK(clk), .RN(rstn), .Q(dout[10]) );
  DFFRHQX1 dout_reg_9_ ( .D(n525), .CK(clk), .RN(rstn), .Q(dout[9]) );
  DFFRHQX1 dout_reg_8_ ( .D(n524), .CK(clk), .RN(rstn), .Q(dout[8]) );
  DFFRHQX1 dout_reg_7_ ( .D(n523), .CK(clk), .RN(rstn), .Q(dout[7]) );
  DFFRHQX1 dout_reg_6_ ( .D(n522), .CK(clk), .RN(rstn), .Q(dout[6]) );
  DFFRHQX1 dout_reg_5_ ( .D(n521), .CK(clk), .RN(rstn), .Q(dout[5]) );
  DFFRHQX1 dout_reg_4_ ( .D(n520), .CK(clk), .RN(rstn), .Q(dout[4]) );
  DFFRHQX1 dout_reg_3_ ( .D(n519), .CK(clk), .RN(rstn), .Q(dout[3]) );
  DFFRHQX1 dout_reg_2_ ( .D(n518), .CK(clk), .RN(rstn), .Q(dout[2]) );
  DFFRHQX1 dout_reg_1_ ( .D(n517), .CK(clk), .RN(rstn), .Q(dout[1]) );
  DFFRHQX1 dout_reg_0_ ( .D(n516), .CK(clk), .RN(rstn), .Q(dout[0]) );
  DFFRHQX1 shift4_flag_reg ( .D(n661), .CK(clk), .RN(rstn), .Q(shift4_flag) );
  DFFRHQX1 start_reg4_reg_0_ ( .D(n662), .CK(clk), .RN(rstn), .Q(start_reg4[0]) );
  DFFRHQX1 ready8_reg ( .D(n668), .CK(clk), .RN(rstn), .Q(ready8) );
  OR3XL U3 ( .A(n221), .B(n225), .C(n672), .Y(n81) );
  AND2X2 U6 ( .A(n309), .B(n225), .Y(n82) );
  AND2X2 U7 ( .A(start), .B(n97), .Y(n83) );
  INVX1 U8 ( .A(n133), .Y(n92) );
  INVX1 U9 ( .A(n133), .Y(n93) );
  INVX1 U10 ( .A(n134), .Y(n94) );
  INVX1 U11 ( .A(n134), .Y(n95) );
  INVX1 U12 ( .A(n134), .Y(n96) );
  INVX1 U13 ( .A(n135), .Y(n98) );
  INVX1 U14 ( .A(n134), .Y(n97) );
  INVX1 U15 ( .A(n133), .Y(n91) );
  INVX1 U16 ( .A(n133), .Y(n99) );
  INVX1 U17 ( .A(n138), .Y(n134) );
  INVX1 U18 ( .A(n138), .Y(n133) );
  INVX1 U19 ( .A(n138), .Y(n135) );
  INVX1 U20 ( .A(n139), .Y(n112) );
  INVX1 U21 ( .A(n144), .Y(n108) );
  INVX1 U22 ( .A(n144), .Y(n110) );
  INVX1 U23 ( .A(n144), .Y(n109) );
  INVX1 U24 ( .A(n139), .Y(n111) );
  INVX1 U25 ( .A(n141), .Y(n122) );
  INVX1 U26 ( .A(n139), .Y(n129) );
  INVX1 U27 ( .A(n139), .Y(n130) );
  INVX1 U28 ( .A(n141), .Y(n123) );
  INVX1 U29 ( .A(n139), .Y(n131) );
  INVX1 U30 ( .A(n140), .Y(n125) );
  INVX1 U31 ( .A(n139), .Y(n132) );
  INVX1 U32 ( .A(n141), .Y(n124) );
  INVX1 U33 ( .A(n139), .Y(n128) );
  INVX1 U34 ( .A(n140), .Y(n127) );
  INVX1 U35 ( .A(n140), .Y(n126) );
  INVX1 U36 ( .A(n141), .Y(n120) );
  INVX1 U37 ( .A(n143), .Y(n116) );
  INVX1 U38 ( .A(n142), .Y(n113) );
  INVX1 U39 ( .A(n140), .Y(n121) );
  INVX1 U40 ( .A(n143), .Y(n115) );
  INVX1 U41 ( .A(n142), .Y(n117) );
  INVX1 U42 ( .A(n142), .Y(n118) );
  INVX1 U43 ( .A(n143), .Y(n114) );
  INVX1 U44 ( .A(n142), .Y(n119) );
  INVX1 U45 ( .A(n144), .Y(n107) );
  INVX1 U46 ( .A(n210), .Y(n103) );
  INVX1 U47 ( .A(n210), .Y(n101) );
  INVX1 U48 ( .A(n210), .Y(n102) );
  INVX1 U49 ( .A(n209), .Y(n105) );
  INVX1 U50 ( .A(n209), .Y(n106) );
  INVX1 U51 ( .A(n209), .Y(n104) );
  INVX1 U52 ( .A(n83), .Y(n89) );
  INVX1 U53 ( .A(n83), .Y(n90) );
  INVX1 U54 ( .A(n211), .Y(n136) );
  INVX1 U55 ( .A(n211), .Y(n137) );
  INVX1 U56 ( .A(n214), .Y(n138) );
  INVX1 U57 ( .A(n214), .Y(n139) );
  INVX1 U58 ( .A(n213), .Y(n141) );
  INVX1 U59 ( .A(n212), .Y(n140) );
  INVX1 U60 ( .A(n212), .Y(n144) );
  INVX1 U61 ( .A(n213), .Y(n142) );
  INVX1 U62 ( .A(n213), .Y(n143) );
  INVX1 U63 ( .A(n211), .Y(n100) );
  INVX1 U64 ( .A(n212), .Y(n211) );
  INVX1 U65 ( .A(n212), .Y(n210) );
  INVX1 U66 ( .A(n212), .Y(n209) );
  INVX1 U67 ( .A(n229), .Y(n225) );
  INVX1 U68 ( .A(n81), .Y(n223) );
  INVX1 U69 ( .A(n81), .Y(n224) );
  INVX1 U70 ( .A(n219), .Y(n217) );
  INVX1 U71 ( .A(n219), .Y(n218) );
  INVX1 U72 ( .A(n446), .Y(n214) );
  INVX1 U73 ( .A(n446), .Y(n213) );
  INVX1 U74 ( .A(n219), .Y(n216) );
  INVX1 U75 ( .A(n81), .Y(n222) );
  INVX1 U76 ( .A(n81), .Y(n220) );
  INVX1 U77 ( .A(n229), .Y(n226) );
  INVX1 U78 ( .A(n229), .Y(n227) );
  INVX1 U79 ( .A(n229), .Y(n228) );
  INVX1 U80 ( .A(n446), .Y(n212) );
  NAND2X1 U81 ( .A(n513), .B(n87), .Y(n446) );
  INVX1 U82 ( .A(start), .Y(n672) );
  INVX1 U83 ( .A(n84), .Y(n87) );
  INVX1 U84 ( .A(n331), .Y(n219) );
  INVX1 U85 ( .A(n514), .Y(n215) );
  INVX1 U86 ( .A(n84), .Y(n88) );
  INVX1 U87 ( .A(n311), .Y(n229) );
  OAI222XL U88 ( .A0(n231), .A1(n89), .B0(n87), .B1(n714), .C0(n98), .C1(n730), 
        .Y(n632) );
  INVX1 U89 ( .A(cal_result[14]), .Y(n231) );
  OAI222XL U90 ( .A0(n230), .A1(n89), .B0(n87), .B1(n713), .C0(n98), .C1(n729), 
        .Y(n630) );
  INVX1 U91 ( .A(cal_result[15]), .Y(n230) );
  OAI222XL U92 ( .A0(n247), .A1(n89), .B0(n88), .B1(n698), .C0(n97), .C1(n714), 
        .Y(n614) );
  INVX1 U93 ( .A(cal_result[30]), .Y(n247) );
  OAI222XL U94 ( .A0(n246), .A1(n90), .B0(n88), .B1(n697), .C0(n97), .C1(n713), 
        .Y(n613) );
  INVX1 U95 ( .A(cal_result[31]), .Y(n246) );
  OAI222XL U96 ( .A0(n263), .A1(n89), .B0(n88), .B1(n682), .C0(n98), .C1(n698), 
        .Y(n598) );
  INVX1 U97 ( .A(cal_result[46]), .Y(n263) );
  OAI222XL U98 ( .A0(n262), .A1(n89), .B0(n88), .B1(n681), .C0(n98), .C1(n697), 
        .Y(n597) );
  INVX1 U99 ( .A(cal_result[47]), .Y(n262) );
  OAI22X1 U100 ( .A0(n91), .A1(n681), .B0(n278), .B1(n90), .Y(n581) );
  INVX1 U101 ( .A(cal_result[63]), .Y(n278) );
  OAI222XL U102 ( .A0(n245), .A1(n90), .B0(n87), .B1(n728), .C0(n99), .C1(n744), .Y(n660) );
  INVX1 U103 ( .A(cal_result[0]), .Y(n245) );
  OAI222XL U104 ( .A0(n244), .A1(n90), .B0(n87), .B1(n727), .C0(n99), .C1(n743), .Y(n658) );
  INVX1 U105 ( .A(cal_result[1]), .Y(n244) );
  OAI222XL U106 ( .A0(n243), .A1(n90), .B0(n87), .B1(n726), .C0(n99), .C1(n742), .Y(n656) );
  INVX1 U107 ( .A(cal_result[2]), .Y(n243) );
  OAI222XL U108 ( .A0(n242), .A1(n90), .B0(n87), .B1(n725), .C0(n99), .C1(n741), .Y(n654) );
  INVX1 U109 ( .A(cal_result[3]), .Y(n242) );
  OAI222XL U110 ( .A0(n241), .A1(n90), .B0(n87), .B1(n724), .C0(n99), .C1(n740), .Y(n652) );
  INVX1 U111 ( .A(cal_result[4]), .Y(n241) );
  OAI222XL U112 ( .A0(n240), .A1(n90), .B0(n87), .B1(n723), .C0(n99), .C1(n739), .Y(n650) );
  INVX1 U113 ( .A(cal_result[5]), .Y(n240) );
  OAI222XL U114 ( .A0(n239), .A1(n90), .B0(n87), .B1(n722), .C0(n99), .C1(n738), .Y(n648) );
  INVX1 U115 ( .A(cal_result[6]), .Y(n239) );
  OAI222XL U116 ( .A0(n238), .A1(n90), .B0(n87), .B1(n721), .C0(n99), .C1(n737), .Y(n646) );
  INVX1 U117 ( .A(cal_result[7]), .Y(n238) );
  OAI222XL U118 ( .A0(n237), .A1(n90), .B0(n87), .B1(n720), .C0(n99), .C1(n736), .Y(n644) );
  INVX1 U119 ( .A(cal_result[8]), .Y(n237) );
  OAI222XL U120 ( .A0(n236), .A1(n89), .B0(n87), .B1(n719), .C0(n98), .C1(n735), .Y(n642) );
  INVX1 U121 ( .A(cal_result[9]), .Y(n236) );
  OAI222XL U122 ( .A0(n235), .A1(n89), .B0(n87), .B1(n718), .C0(n98), .C1(n734), .Y(n640) );
  INVX1 U123 ( .A(cal_result[10]), .Y(n235) );
  OAI222XL U124 ( .A0(n234), .A1(n89), .B0(n87), .B1(n717), .C0(n98), .C1(n733), .Y(n638) );
  INVX1 U125 ( .A(cal_result[11]), .Y(n234) );
  OAI222XL U126 ( .A0(n233), .A1(n89), .B0(n87), .B1(n716), .C0(n98), .C1(n732), .Y(n636) );
  INVX1 U127 ( .A(cal_result[12]), .Y(n233) );
  OAI222XL U128 ( .A0(n232), .A1(n89), .B0(n87), .B1(n715), .C0(n98), .C1(n731), .Y(n634) );
  INVX1 U129 ( .A(cal_result[13]), .Y(n232) );
  OAI222XL U130 ( .A0(n261), .A1(n89), .B0(n87), .B1(n712), .C0(n97), .C1(n728), .Y(n628) );
  INVX1 U131 ( .A(cal_result[16]), .Y(n261) );
  OAI222XL U132 ( .A0(n260), .A1(n89), .B0(n87), .B1(n711), .C0(n97), .C1(n727), .Y(n627) );
  INVX1 U133 ( .A(cal_result[17]), .Y(n260) );
  OAI222XL U134 ( .A0(n259), .A1(n89), .B0(n88), .B1(n710), .C0(n97), .C1(n726), .Y(n626) );
  INVX1 U135 ( .A(cal_result[18]), .Y(n259) );
  OAI222XL U136 ( .A0(n258), .A1(n89), .B0(n88), .B1(n709), .C0(n97), .C1(n725), .Y(n625) );
  INVX1 U137 ( .A(cal_result[19]), .Y(n258) );
  OAI222XL U138 ( .A0(n257), .A1(n89), .B0(n88), .B1(n708), .C0(n97), .C1(n724), .Y(n624) );
  INVX1 U139 ( .A(cal_result[20]), .Y(n257) );
  OAI222XL U140 ( .A0(n256), .A1(n89), .B0(n88), .B1(n707), .C0(n97), .C1(n723), .Y(n623) );
  INVX1 U141 ( .A(cal_result[21]), .Y(n256) );
  OAI222XL U142 ( .A0(n255), .A1(n89), .B0(n88), .B1(n706), .C0(n97), .C1(n722), .Y(n622) );
  INVX1 U143 ( .A(cal_result[22]), .Y(n255) );
  OAI222XL U144 ( .A0(n254), .A1(n89), .B0(n88), .B1(n705), .C0(n97), .C1(n721), .Y(n621) );
  INVX1 U145 ( .A(cal_result[23]), .Y(n254) );
  OAI222XL U146 ( .A0(n253), .A1(n89), .B0(n88), .B1(n704), .C0(n97), .C1(n720), .Y(n620) );
  INVX1 U147 ( .A(cal_result[24]), .Y(n253) );
  OAI222XL U148 ( .A0(n252), .A1(n89), .B0(n88), .B1(n703), .C0(n97), .C1(n719), .Y(n619) );
  INVX1 U149 ( .A(cal_result[25]), .Y(n252) );
  OAI222XL U150 ( .A0(n251), .A1(n89), .B0(n88), .B1(n702), .C0(n97), .C1(n718), .Y(n618) );
  INVX1 U151 ( .A(cal_result[26]), .Y(n251) );
  OAI222XL U152 ( .A0(n250), .A1(n89), .B0(n88), .B1(n701), .C0(n97), .C1(n717), .Y(n617) );
  INVX1 U153 ( .A(cal_result[27]), .Y(n250) );
  OAI222XL U154 ( .A0(n249), .A1(n89), .B0(n88), .B1(n700), .C0(n97), .C1(n716), .Y(n616) );
  INVX1 U155 ( .A(cal_result[28]), .Y(n249) );
  OAI222XL U156 ( .A0(n248), .A1(n89), .B0(n88), .B1(n699), .C0(n97), .C1(n715), .Y(n615) );
  INVX1 U157 ( .A(cal_result[29]), .Y(n248) );
  OAI222XL U158 ( .A0(n277), .A1(n90), .B0(n88), .B1(n696), .C0(n98), .C1(n712), .Y(n612) );
  INVX1 U159 ( .A(cal_result[32]), .Y(n277) );
  OAI222XL U160 ( .A0(n276), .A1(n89), .B0(n88), .B1(n695), .C0(n98), .C1(n711), .Y(n611) );
  INVX1 U161 ( .A(cal_result[33]), .Y(n276) );
  OAI222XL U162 ( .A0(n275), .A1(n90), .B0(n88), .B1(n694), .C0(n98), .C1(n710), .Y(n610) );
  INVX1 U163 ( .A(cal_result[34]), .Y(n275) );
  OAI222XL U164 ( .A0(n274), .A1(n89), .B0(n88), .B1(n693), .C0(n98), .C1(n709), .Y(n609) );
  INVX1 U165 ( .A(cal_result[35]), .Y(n274) );
  OAI222XL U166 ( .A0(n273), .A1(n90), .B0(n88), .B1(n692), .C0(n98), .C1(n708), .Y(n608) );
  INVX1 U167 ( .A(cal_result[36]), .Y(n273) );
  OAI222XL U168 ( .A0(n272), .A1(n89), .B0(n88), .B1(n691), .C0(n98), .C1(n707), .Y(n607) );
  INVX1 U169 ( .A(cal_result[37]), .Y(n272) );
  OAI222XL U170 ( .A0(n271), .A1(n90), .B0(n88), .B1(n690), .C0(n98), .C1(n706), .Y(n606) );
  INVX1 U171 ( .A(cal_result[38]), .Y(n271) );
  OAI222XL U172 ( .A0(n270), .A1(n89), .B0(n88), .B1(n689), .C0(n98), .C1(n705), .Y(n605) );
  INVX1 U173 ( .A(cal_result[39]), .Y(n270) );
  OAI222XL U174 ( .A0(n269), .A1(n90), .B0(n88), .B1(n688), .C0(n98), .C1(n704), .Y(n604) );
  INVX1 U175 ( .A(cal_result[40]), .Y(n269) );
  OAI222XL U176 ( .A0(n268), .A1(n89), .B0(n88), .B1(n687), .C0(n98), .C1(n703), .Y(n603) );
  INVX1 U177 ( .A(cal_result[41]), .Y(n268) );
  OAI222XL U178 ( .A0(n267), .A1(n90), .B0(n88), .B1(n686), .C0(n98), .C1(n702), .Y(n602) );
  INVX1 U179 ( .A(cal_result[42]), .Y(n267) );
  OAI222XL U180 ( .A0(n266), .A1(n89), .B0(n88), .B1(n685), .C0(n98), .C1(n701), .Y(n601) );
  INVX1 U181 ( .A(cal_result[43]), .Y(n266) );
  OAI222XL U182 ( .A0(n265), .A1(n90), .B0(n88), .B1(n684), .C0(n98), .C1(n700), .Y(n600) );
  INVX1 U183 ( .A(cal_result[44]), .Y(n265) );
  OAI222XL U184 ( .A0(n264), .A1(n89), .B0(n88), .B1(n683), .C0(n98), .C1(n699), .Y(n599) );
  INVX1 U185 ( .A(cal_result[45]), .Y(n264) );
  OAI22X1 U186 ( .A0(n91), .A1(n696), .B0(n671), .B1(n90), .Y(n596) );
  INVX1 U187 ( .A(cal_result[48]), .Y(n671) );
  OAI22X1 U188 ( .A0(n92), .A1(n695), .B0(n670), .B1(n90), .Y(n595) );
  INVX1 U189 ( .A(cal_result[49]), .Y(n670) );
  OAI22X1 U190 ( .A0(n92), .A1(n693), .B0(n448), .B1(n90), .Y(n593) );
  INVX1 U191 ( .A(cal_result[51]), .Y(n448) );
  OAI22X1 U192 ( .A0(n91), .A1(n692), .B0(n447), .B1(n90), .Y(n592) );
  INVX1 U193 ( .A(cal_result[52]), .Y(n447) );
  OAI22X1 U194 ( .A0(n92), .A1(n691), .B0(n314), .B1(n90), .Y(n591) );
  INVX1 U195 ( .A(cal_result[53]), .Y(n314) );
  OAI22X1 U196 ( .A0(n91), .A1(n690), .B0(n307), .B1(n90), .Y(n590) );
  INVX1 U197 ( .A(cal_result[54]), .Y(n307) );
  OAI22X1 U198 ( .A0(n92), .A1(n689), .B0(n287), .B1(n90), .Y(n589) );
  INVX1 U199 ( .A(cal_result[55]), .Y(n287) );
  OAI22X1 U200 ( .A0(n91), .A1(n688), .B0(n285), .B1(n90), .Y(n588) );
  INVX1 U201 ( .A(cal_result[56]), .Y(n285) );
  OAI22X1 U202 ( .A0(n91), .A1(n687), .B0(n284), .B1(n90), .Y(n587) );
  INVX1 U203 ( .A(cal_result[57]), .Y(n284) );
  OAI22X1 U204 ( .A0(n91), .A1(n686), .B0(n283), .B1(n90), .Y(n586) );
  INVX1 U205 ( .A(cal_result[58]), .Y(n283) );
  OAI22X1 U206 ( .A0(n91), .A1(n684), .B0(n281), .B1(n90), .Y(n584) );
  INVX1 U207 ( .A(cal_result[60]), .Y(n281) );
  OAI22X1 U208 ( .A0(n91), .A1(n683), .B0(n280), .B1(n90), .Y(n583) );
  INVX1 U209 ( .A(cal_result[61]), .Y(n280) );
  OAI22X1 U210 ( .A0(n91), .A1(n682), .B0(n279), .B1(n90), .Y(n582) );
  INVX1 U211 ( .A(cal_result[62]), .Y(n279) );
  OAI22X1 U212 ( .A0(n91), .A1(n694), .B0(n669), .B1(n90), .Y(n594) );
  INVX1 U213 ( .A(cal_result[50]), .Y(n669) );
  OAI22X1 U214 ( .A0(n91), .A1(n685), .B0(n282), .B1(n89), .Y(n585) );
  INVX1 U215 ( .A(cal_result[59]), .Y(n282) );
  NAND2X1 U216 ( .A(n444), .B(n221), .Y(n513) );
  NOR2X1 U217 ( .A(n443), .B(n444), .Y(n311) );
  AOI2BB1X1 U218 ( .A0N(n221), .A1N(n443), .B0(n225), .Y(n331) );
  NAND2X1 U219 ( .A(n308), .B(n310), .Y(n443) );
  NAND3X1 U220 ( .A(n673), .B(n672), .C(n286), .Y(n445) );
  INVX1 U221 ( .A(n286), .Y(p2s_ready) );
  AND2X2 U222 ( .A(n312), .B(n445), .Y(n308) );
  NAND3X1 U223 ( .A(n310), .B(n309), .C(n445), .Y(n84) );
  NAND3X1 U224 ( .A(n310), .B(n309), .C(n513), .Y(n514) );
  OAI22X1 U225 ( .A0(n215), .A1(n678), .B0(n514), .B1(n679), .Y(n663) );
  OAI22X1 U226 ( .A0(n215), .A1(n677), .B0(n514), .B1(n678), .Y(n664) );
  OAI22X1 U227 ( .A0(n215), .A1(n676), .B0(n514), .B1(n677), .Y(n665) );
  OAI22X1 U228 ( .A0(n215), .A1(n675), .B0(n514), .B1(n676), .Y(n666) );
  OAI22X1 U229 ( .A0(n215), .A1(n672), .B0(n514), .B1(n675), .Y(n667) );
  OAI22X1 U230 ( .A0(n215), .A1(n679), .B0(n680), .B1(n514), .Y(n662) );
  AND2X2 U231 ( .A(n310), .B(n672), .Y(n306) );
  OAI21XL U232 ( .A0(n444), .A1(n673), .B0(n513), .Y(n661) );
  NOR2X1 U233 ( .A(start_reg4[0]), .B(ready8), .Y(n286) );
  INVX1 U234 ( .A(n429), .Y(n67) );
  AOI222X1 U235 ( .A0(n224), .A1(cal_result[13]), .B0(n218), .B1(
        result_reg8[29]), .C0(n228), .C1(result_reg8[13]), .Y(n429) );
  INVX1 U236 ( .A(n428), .Y(n66) );
  AOI222X1 U237 ( .A0(n224), .A1(cal_result[14]), .B0(n218), .B1(
        result_reg8[30]), .C0(n228), .C1(result_reg8[14]), .Y(n428) );
  INVX1 U238 ( .A(n427), .Y(n65) );
  AOI222X1 U239 ( .A0(n224), .A1(cal_result[15]), .B0(n218), .B1(
        result_reg8[31]), .C0(n228), .C1(result_reg8[15]), .Y(n427) );
  INVX1 U240 ( .A(n413), .Y(n51) );
  AOI222X1 U241 ( .A0(n224), .A1(cal_result[29]), .B0(n217), .B1(
        result_reg8[45]), .C0(n228), .C1(result_reg8[29]), .Y(n413) );
  INVX1 U242 ( .A(n412), .Y(n50) );
  AOI222X1 U243 ( .A0(n224), .A1(cal_result[30]), .B0(n217), .B1(
        result_reg8[46]), .C0(n226), .C1(result_reg8[30]), .Y(n412) );
  INVX1 U244 ( .A(n411), .Y(n49) );
  AOI222X1 U245 ( .A0(n224), .A1(cal_result[31]), .B0(n217), .B1(
        result_reg8[47]), .C0(n227), .C1(result_reg8[31]), .Y(n411) );
  INVX1 U246 ( .A(n397), .Y(n35) );
  AOI222X1 U247 ( .A0(n223), .A1(cal_result[45]), .B0(n217), .B1(
        result_reg8[61]), .C0(n227), .C1(result_reg8[45]), .Y(n397) );
  INVX1 U248 ( .A(n396), .Y(n34) );
  AOI222X1 U249 ( .A0(n223), .A1(cal_result[46]), .B0(n217), .B1(
        result_reg8[62]), .C0(n227), .C1(result_reg8[46]), .Y(n396) );
  INVX1 U250 ( .A(n395), .Y(n33) );
  AOI222X1 U251 ( .A0(n223), .A1(cal_result[47]), .B0(n217), .B1(
        result_reg8[63]), .C0(n227), .C1(result_reg8[47]), .Y(n395) );
  INVX1 U252 ( .A(n381), .Y(n19) );
  AOI222X1 U253 ( .A0(n223), .A1(cal_result[61]), .B0(n218), .B1(
        result_reg8[77]), .C0(n227), .C1(result_reg8[61]), .Y(n381) );
  INVX1 U254 ( .A(n380), .Y(n18) );
  AOI222X1 U255 ( .A0(n223), .A1(cal_result[62]), .B0(n218), .B1(
        result_reg8[78]), .C0(n227), .C1(result_reg8[62]), .Y(n380) );
  INVX1 U256 ( .A(n379), .Y(n17) );
  AOI222X1 U257 ( .A0(n223), .A1(cal_result[63]), .B0(n218), .B1(
        result_reg8[79]), .C0(n226), .C1(result_reg8[63]), .Y(n379) );
  NOR2X1 U258 ( .A(mode[1]), .B(n672), .Y(n444) );
  NAND3X1 U259 ( .A(n674), .B(n672), .C(start_reg4[0]), .Y(n309) );
  NAND3X1 U260 ( .A(n286), .B(n672), .C(shift4_flag), .Y(n310) );
  INVX1 U261 ( .A(n316), .Y(n3) );
  AOI22X1 U262 ( .A0(n228), .A1(result_reg8[125]), .B0(cal_result[125]), .B1(
        n222), .Y(n316) );
  OAI2BB1X1 U263 ( .A0N(n226), .A1N(result_reg8[78]), .B0(n364), .Y(n566) );
  AOI22X1 U264 ( .A0(result_reg8[94]), .A1(n216), .B0(cal_result[78]), .B1(
        n222), .Y(n364) );
  OAI2BB1X1 U265 ( .A0N(n226), .A1N(result_reg8[79]), .B0(n363), .Y(n565) );
  AOI22X1 U266 ( .A0(result_reg8[95]), .A1(n216), .B0(cal_result[79]), .B1(
        n220), .Y(n363) );
  OAI2BB1X1 U267 ( .A0N(n225), .A1N(result_reg8[94]), .B0(n348), .Y(n550) );
  AOI22X1 U268 ( .A0(result_reg8[110]), .A1(n216), .B0(cal_result[94]), .B1(
        n222), .Y(n348) );
  OAI2BB1X1 U269 ( .A0N(n225), .A1N(result_reg8[95]), .B0(n347), .Y(n549) );
  AOI22X1 U270 ( .A0(result_reg8[111]), .A1(n216), .B0(cal_result[95]), .B1(
        n222), .Y(n347) );
  OAI2BB1X1 U271 ( .A0N(n225), .A1N(result_reg8[110]), .B0(n332), .Y(n534) );
  AOI22X1 U272 ( .A0(n218), .A1(result_reg8[126]), .B0(cal_result[110]), .B1(
        n220), .Y(n332) );
  OAI2BB1X1 U273 ( .A0N(n225), .A1N(result_reg8[111]), .B0(n330), .Y(n533) );
  AOI22X1 U274 ( .A0(n331), .A1(result_reg8[127]), .B0(cal_result[111]), .B1(
        n220), .Y(n330) );
  NAND2X1 U275 ( .A(ready8), .B(n672), .Y(n312) );
  OAI2BB2X1 U276 ( .B0(n106), .B1(n744), .A0N(n135), .A1N(result_reg4[64]), 
        .Y(n659) );
  OAI2BB2X1 U277 ( .B0(n105), .B1(n743), .A0N(n136), .A1N(result_reg4[65]), 
        .Y(n657) );
  OAI2BB2X1 U278 ( .B0(n103), .B1(n742), .A0N(n136), .A1N(result_reg4[66]), 
        .Y(n655) );
  OAI2BB2X1 U279 ( .B0(n100), .B1(n741), .A0N(n136), .A1N(result_reg4[67]), 
        .Y(n653) );
  OAI2BB2X1 U280 ( .B0(n107), .B1(n740), .A0N(n136), .A1N(result_reg4[68]), 
        .Y(n651) );
  OAI2BB2X1 U281 ( .B0(n100), .B1(n739), .A0N(n137), .A1N(result_reg4[69]), 
        .Y(n649) );
  OAI2BB2X1 U282 ( .B0(n101), .B1(n738), .A0N(n135), .A1N(result_reg4[70]), 
        .Y(n647) );
  OAI2BB2X1 U283 ( .B0(n104), .B1(n737), .A0N(n135), .A1N(result_reg4[71]), 
        .Y(n645) );
  OAI2BB2X1 U284 ( .B0(n107), .B1(n736), .A0N(n136), .A1N(result_reg4[72]), 
        .Y(n643) );
  OAI2BB2X1 U285 ( .B0(n103), .B1(n735), .A0N(n135), .A1N(result_reg4[73]), 
        .Y(n641) );
  OAI2BB2X1 U286 ( .B0(n102), .B1(n734), .A0N(n137), .A1N(result_reg4[74]), 
        .Y(n639) );
  OAI2BB2X1 U287 ( .B0(n101), .B1(n733), .A0N(n136), .A1N(result_reg4[75]), 
        .Y(n637) );
  OAI2BB2X1 U288 ( .B0(n102), .B1(n732), .A0N(n137), .A1N(result_reg4[76]), 
        .Y(n635) );
  OAI2BB2X1 U289 ( .B0(n105), .B1(n731), .A0N(n137), .A1N(result_reg4[77]), 
        .Y(n633) );
  OAI2BB2X1 U290 ( .B0(n106), .B1(n730), .A0N(n137), .A1N(result_reg4[78]), 
        .Y(n631) );
  OAI2BB2X1 U291 ( .B0(n104), .B1(n729), .A0N(n137), .A1N(result_reg4[79]), 
        .Y(n629) );
  INVX1 U292 ( .A(ready8), .Y(n674) );
  INVX1 U293 ( .A(start_reg4[0]), .Y(n680) );
  INVX1 U294 ( .A(mode[0]), .Y(n221) );
  INVX1 U295 ( .A(n315), .Y(n2) );
  AOI22X1 U296 ( .A0(n228), .A1(result_reg8[126]), .B0(cal_result[126]), .B1(
        n220), .Y(n315) );
  INVX1 U297 ( .A(n313), .Y(n1) );
  AOI22X1 U298 ( .A0(n228), .A1(result_reg8[127]), .B0(cal_result[127]), .B1(
        n222), .Y(n313) );
  OAI2BB1X1 U299 ( .A0N(n226), .A1N(result_reg8[77]), .B0(n365), .Y(n567) );
  AOI22X1 U300 ( .A0(result_reg8[93]), .A1(n216), .B0(cal_result[77]), .B1(
        n222), .Y(n365) );
  OAI2BB1X1 U301 ( .A0N(n226), .A1N(result_reg8[93]), .B0(n349), .Y(n551) );
  AOI22X1 U302 ( .A0(result_reg8[109]), .A1(n216), .B0(cal_result[93]), .B1(
        n222), .Y(n349) );
  OAI2BB1X1 U303 ( .A0N(n225), .A1N(result_reg8[109]), .B0(n333), .Y(n535) );
  AOI22X1 U304 ( .A0(n331), .A1(result_reg8[125]), .B0(cal_result[109]), .B1(
        n220), .Y(n333) );
  INVX1 U305 ( .A(n510), .Y(n192) );
  AOI22X1 U306 ( .A0(n92), .A1(result_reg4[32]), .B0(n121), .B1(
        result_reg4[16]), .Y(n510) );
  INVX1 U307 ( .A(n511), .Y(n176) );
  AOI22X1 U308 ( .A0(n92), .A1(result_reg4[48]), .B0(n116), .B1(
        result_reg4[32]), .Y(n511) );
  INVX1 U309 ( .A(n512), .Y(n160) );
  AOI22X1 U310 ( .A0(n92), .A1(result_reg4[64]), .B0(n114), .B1(
        result_reg4[48]), .Y(n512) );
  INVX1 U311 ( .A(n506), .Y(n191) );
  AOI22X1 U312 ( .A0(n93), .A1(result_reg4[33]), .B0(n122), .B1(
        result_reg4[17]), .Y(n506) );
  INVX1 U313 ( .A(n507), .Y(n175) );
  AOI22X1 U314 ( .A0(n92), .A1(result_reg4[49]), .B0(n122), .B1(
        result_reg4[33]), .Y(n507) );
  INVX1 U315 ( .A(n508), .Y(n159) );
  AOI22X1 U316 ( .A0(n93), .A1(result_reg4[65]), .B0(n131), .B1(
        result_reg4[49]), .Y(n508) );
  INVX1 U317 ( .A(n502), .Y(n190) );
  AOI22X1 U318 ( .A0(n92), .A1(result_reg4[34]), .B0(n127), .B1(
        result_reg4[18]), .Y(n502) );
  INVX1 U319 ( .A(n503), .Y(n174) );
  AOI22X1 U320 ( .A0(n93), .A1(result_reg4[50]), .B0(n118), .B1(
        result_reg4[34]), .Y(n503) );
  INVX1 U321 ( .A(n504), .Y(n158) );
  AOI22X1 U322 ( .A0(n92), .A1(result_reg4[66]), .B0(n119), .B1(
        result_reg4[50]), .Y(n504) );
  INVX1 U323 ( .A(n498), .Y(n189) );
  AOI22X1 U324 ( .A0(n94), .A1(result_reg4[35]), .B0(n126), .B1(
        result_reg4[19]), .Y(n498) );
  INVX1 U325 ( .A(n499), .Y(n173) );
  AOI22X1 U326 ( .A0(n92), .A1(result_reg4[51]), .B0(n129), .B1(
        result_reg4[35]), .Y(n499) );
  INVX1 U327 ( .A(n500), .Y(n157) );
  AOI22X1 U328 ( .A0(n93), .A1(result_reg4[67]), .B0(n124), .B1(
        result_reg4[51]), .Y(n500) );
  INVX1 U329 ( .A(n494), .Y(n188) );
  AOI22X1 U330 ( .A0(n93), .A1(result_reg4[36]), .B0(n129), .B1(
        result_reg4[20]), .Y(n494) );
  INVX1 U331 ( .A(n495), .Y(n172) );
  AOI22X1 U332 ( .A0(n93), .A1(result_reg4[52]), .B0(n131), .B1(
        result_reg4[36]), .Y(n495) );
  INVX1 U333 ( .A(n496), .Y(n156) );
  AOI22X1 U334 ( .A0(n93), .A1(result_reg4[68]), .B0(n132), .B1(
        result_reg4[52]), .Y(n496) );
  INVX1 U335 ( .A(n490), .Y(n187) );
  AOI22X1 U336 ( .A0(n94), .A1(result_reg4[37]), .B0(n130), .B1(
        result_reg4[21]), .Y(n490) );
  INVX1 U337 ( .A(n491), .Y(n171) );
  AOI22X1 U338 ( .A0(n93), .A1(result_reg4[53]), .B0(n123), .B1(
        result_reg4[37]), .Y(n491) );
  INVX1 U339 ( .A(n492), .Y(n155) );
  AOI22X1 U340 ( .A0(n93), .A1(result_reg4[69]), .B0(n130), .B1(
        result_reg4[53]), .Y(n492) );
  INVX1 U341 ( .A(n486), .Y(n186) );
  AOI22X1 U342 ( .A0(n94), .A1(result_reg4[38]), .B0(n123), .B1(
        result_reg4[22]), .Y(n486) );
  INVX1 U343 ( .A(n487), .Y(n170) );
  AOI22X1 U344 ( .A0(n94), .A1(result_reg4[54]), .B0(n125), .B1(
        result_reg4[38]), .Y(n487) );
  INVX1 U345 ( .A(n488), .Y(n154) );
  AOI22X1 U346 ( .A0(n93), .A1(result_reg4[70]), .B0(n131), .B1(
        result_reg4[54]), .Y(n488) );
  INVX1 U347 ( .A(n482), .Y(n185) );
  AOI22X1 U348 ( .A0(n94), .A1(result_reg4[39]), .B0(n125), .B1(
        result_reg4[23]), .Y(n482) );
  INVX1 U349 ( .A(n483), .Y(n169) );
  AOI22X1 U350 ( .A0(n94), .A1(result_reg4[55]), .B0(n132), .B1(
        result_reg4[39]), .Y(n483) );
  INVX1 U351 ( .A(n484), .Y(n153) );
  AOI22X1 U352 ( .A0(n94), .A1(result_reg4[71]), .B0(n124), .B1(
        result_reg4[55]), .Y(n484) );
  INVX1 U353 ( .A(n478), .Y(n184) );
  AOI22X1 U354 ( .A0(n94), .A1(result_reg4[40]), .B0(n128), .B1(
        result_reg4[24]), .Y(n478) );
  INVX1 U355 ( .A(n479), .Y(n168) );
  AOI22X1 U356 ( .A0(n95), .A1(result_reg4[56]), .B0(n128), .B1(
        result_reg4[40]), .Y(n479) );
  INVX1 U357 ( .A(n480), .Y(n152) );
  AOI22X1 U358 ( .A0(n94), .A1(result_reg4[72]), .B0(n127), .B1(
        result_reg4[56]), .Y(n480) );
  INVX1 U359 ( .A(n474), .Y(n183) );
  AOI22X1 U360 ( .A0(n95), .A1(result_reg4[41]), .B0(n115), .B1(
        result_reg4[25]), .Y(n474) );
  INVX1 U361 ( .A(n475), .Y(n167) );
  AOI22X1 U362 ( .A0(n94), .A1(result_reg4[57]), .B0(n117), .B1(
        result_reg4[41]), .Y(n475) );
  INVX1 U363 ( .A(n476), .Y(n151) );
  AOI22X1 U364 ( .A0(n95), .A1(result_reg4[73]), .B0(n126), .B1(
        result_reg4[57]), .Y(n476) );
  INVX1 U365 ( .A(n470), .Y(n182) );
  AOI22X1 U366 ( .A0(n95), .A1(result_reg4[42]), .B0(n120), .B1(
        result_reg4[26]), .Y(n470) );
  INVX1 U367 ( .A(n471), .Y(n166) );
  AOI22X1 U368 ( .A0(n95), .A1(result_reg4[58]), .B0(n120), .B1(
        result_reg4[42]), .Y(n471) );
  INVX1 U369 ( .A(n472), .Y(n150) );
  AOI22X1 U370 ( .A0(n95), .A1(result_reg4[74]), .B0(n116), .B1(
        result_reg4[58]), .Y(n472) );
  INVX1 U371 ( .A(n466), .Y(n181) );
  AOI22X1 U372 ( .A0(n95), .A1(result_reg4[43]), .B0(n129), .B1(
        result_reg4[27]), .Y(n466) );
  INVX1 U373 ( .A(n467), .Y(n165) );
  AOI22X1 U374 ( .A0(n95), .A1(result_reg4[59]), .B0(n128), .B1(
        result_reg4[43]), .Y(n467) );
  INVX1 U375 ( .A(n468), .Y(n149) );
  AOI22X1 U376 ( .A0(n95), .A1(result_reg4[75]), .B0(n120), .B1(
        result_reg4[59]), .Y(n468) );
  INVX1 U377 ( .A(n462), .Y(n180) );
  AOI22X1 U378 ( .A0(n96), .A1(result_reg4[44]), .B0(n113), .B1(
        result_reg4[28]), .Y(n462) );
  INVX1 U379 ( .A(n463), .Y(n164) );
  AOI22X1 U380 ( .A0(n96), .A1(result_reg4[60]), .B0(n116), .B1(
        result_reg4[44]), .Y(n463) );
  INVX1 U381 ( .A(n464), .Y(n148) );
  AOI22X1 U382 ( .A0(n95), .A1(result_reg4[76]), .B0(n113), .B1(
        result_reg4[60]), .Y(n464) );
  INVX1 U383 ( .A(n458), .Y(n179) );
  AOI22X1 U384 ( .A0(n96), .A1(result_reg4[45]), .B0(n121), .B1(
        result_reg4[29]), .Y(n458) );
  INVX1 U385 ( .A(n459), .Y(n163) );
  AOI22X1 U386 ( .A0(n96), .A1(result_reg4[61]), .B0(n115), .B1(
        result_reg4[45]), .Y(n459) );
  INVX1 U387 ( .A(n460), .Y(n147) );
  AOI22X1 U388 ( .A0(n96), .A1(result_reg4[77]), .B0(n121), .B1(
        result_reg4[61]), .Y(n460) );
  INVX1 U389 ( .A(n454), .Y(n178) );
  AOI22X1 U390 ( .A0(n96), .A1(result_reg4[46]), .B0(n117), .B1(
        result_reg4[30]), .Y(n454) );
  INVX1 U391 ( .A(n455), .Y(n162) );
  AOI22X1 U392 ( .A0(n96), .A1(result_reg4[62]), .B0(n118), .B1(
        result_reg4[46]), .Y(n455) );
  INVX1 U393 ( .A(n456), .Y(n146) );
  AOI22X1 U394 ( .A0(n96), .A1(result_reg4[78]), .B0(n114), .B1(
        result_reg4[62]), .Y(n456) );
  INVX1 U395 ( .A(n450), .Y(n177) );
  AOI22X1 U396 ( .A0(n97), .A1(result_reg4[47]), .B0(n119), .B1(
        result_reg4[31]), .Y(n450) );
  INVX1 U397 ( .A(n451), .Y(n161) );
  AOI22X1 U398 ( .A0(n97), .A1(result_reg4[63]), .B0(n114), .B1(
        result_reg4[47]), .Y(n451) );
  INVX1 U399 ( .A(n452), .Y(n145) );
  AOI22X1 U400 ( .A0(n97), .A1(result_reg4[79]), .B0(n130), .B1(
        result_reg4[63]), .Y(n452) );
  INVX1 U401 ( .A(n509), .Y(n208) );
  AOI22X1 U402 ( .A0(n92), .A1(result_reg4[16]), .B0(result_reg4[0]), .B1(n112), .Y(n509) );
  INVX1 U403 ( .A(n505), .Y(n207) );
  AOI22X1 U404 ( .A0(n92), .A1(result_reg4[17]), .B0(result_reg4[1]), .B1(n111), .Y(n505) );
  INVX1 U405 ( .A(n501), .Y(n206) );
  AOI22X1 U406 ( .A0(n93), .A1(result_reg4[18]), .B0(result_reg4[2]), .B1(n112), .Y(n501) );
  INVX1 U407 ( .A(n497), .Y(n205) );
  AOI22X1 U408 ( .A0(n93), .A1(result_reg4[19]), .B0(result_reg4[3]), .B1(n132), .Y(n497) );
  INVX1 U409 ( .A(n493), .Y(n204) );
  AOI22X1 U410 ( .A0(n94), .A1(result_reg4[20]), .B0(result_reg4[4]), .B1(n110), .Y(n493) );
  INVX1 U411 ( .A(n489), .Y(n203) );
  AOI22X1 U412 ( .A0(n93), .A1(result_reg4[21]), .B0(result_reg4[5]), .B1(n108), .Y(n489) );
  INVX1 U413 ( .A(n485), .Y(n202) );
  AOI22X1 U414 ( .A0(n94), .A1(result_reg4[22]), .B0(result_reg4[6]), .B1(n109), .Y(n485) );
  INVX1 U415 ( .A(n481), .Y(n201) );
  AOI22X1 U416 ( .A0(n94), .A1(result_reg4[23]), .B0(result_reg4[7]), .B1(n112), .Y(n481) );
  INVX1 U417 ( .A(n477), .Y(n200) );
  AOI22X1 U418 ( .A0(n95), .A1(result_reg4[24]), .B0(result_reg4[8]), .B1(n110), .Y(n477) );
  INVX1 U419 ( .A(n473), .Y(n199) );
  AOI22X1 U420 ( .A0(n95), .A1(result_reg4[25]), .B0(result_reg4[9]), .B1(n108), .Y(n473) );
  INVX1 U421 ( .A(n469), .Y(n198) );
  AOI22X1 U422 ( .A0(n96), .A1(result_reg4[26]), .B0(result_reg4[10]), .B1(
        n111), .Y(n469) );
  INVX1 U423 ( .A(n465), .Y(n197) );
  AOI22X1 U424 ( .A0(n95), .A1(result_reg4[27]), .B0(result_reg4[11]), .B1(
        n110), .Y(n465) );
  INVX1 U425 ( .A(n461), .Y(n196) );
  AOI22X1 U426 ( .A0(n96), .A1(result_reg4[28]), .B0(result_reg4[12]), .B1(
        n109), .Y(n461) );
  INVX1 U427 ( .A(n457), .Y(n195) );
  AOI22X1 U428 ( .A0(n96), .A1(result_reg4[29]), .B0(result_reg4[13]), .B1(
        n112), .Y(n457) );
  INVX1 U429 ( .A(n453), .Y(n194) );
  AOI22X1 U430 ( .A0(n96), .A1(result_reg4[30]), .B0(result_reg4[14]), .B1(
        n111), .Y(n453) );
  INVX1 U431 ( .A(n449), .Y(n193) );
  AOI22X1 U432 ( .A0(n96), .A1(result_reg4[31]), .B0(result_reg4[15]), .B1(
        n111), .Y(n449) );
  INVX1 U433 ( .A(n442), .Y(n80) );
  AOI222X1 U434 ( .A0(n220), .A1(cal_result[0]), .B0(n331), .B1(
        result_reg8[16]), .C0(n226), .C1(result_reg8[0]), .Y(n442) );
  INVX1 U435 ( .A(n441), .Y(n79) );
  AOI222X1 U436 ( .A0(n220), .A1(cal_result[1]), .B0(n331), .B1(
        result_reg8[17]), .C0(n228), .C1(result_reg8[1]), .Y(n441) );
  INVX1 U437 ( .A(n440), .Y(n78) );
  AOI222X1 U438 ( .A0(n222), .A1(cal_result[2]), .B0(n218), .B1(
        result_reg8[18]), .C0(n228), .C1(result_reg8[2]), .Y(n440) );
  INVX1 U439 ( .A(n439), .Y(n77) );
  AOI222X1 U440 ( .A0(n220), .A1(cal_result[3]), .B0(n218), .B1(
        result_reg8[19]), .C0(n228), .C1(result_reg8[3]), .Y(n439) );
  INVX1 U441 ( .A(n438), .Y(n76) );
  AOI222X1 U442 ( .A0(n224), .A1(cal_result[4]), .B0(n218), .B1(
        result_reg8[20]), .C0(n228), .C1(result_reg8[4]), .Y(n438) );
  INVX1 U443 ( .A(n437), .Y(n75) );
  AOI222X1 U444 ( .A0(n224), .A1(cal_result[5]), .B0(n218), .B1(
        result_reg8[21]), .C0(n228), .C1(result_reg8[5]), .Y(n437) );
  INVX1 U445 ( .A(n436), .Y(n74) );
  AOI222X1 U446 ( .A0(n224), .A1(cal_result[6]), .B0(n218), .B1(
        result_reg8[22]), .C0(n228), .C1(result_reg8[6]), .Y(n436) );
  INVX1 U447 ( .A(n435), .Y(n73) );
  AOI222X1 U448 ( .A0(n224), .A1(cal_result[7]), .B0(n218), .B1(
        result_reg8[23]), .C0(n228), .C1(result_reg8[7]), .Y(n435) );
  INVX1 U449 ( .A(n434), .Y(n72) );
  AOI222X1 U450 ( .A0(n224), .A1(cal_result[8]), .B0(n218), .B1(
        result_reg8[24]), .C0(n228), .C1(result_reg8[8]), .Y(n434) );
  INVX1 U451 ( .A(n433), .Y(n71) );
  AOI222X1 U452 ( .A0(n224), .A1(cal_result[9]), .B0(n218), .B1(
        result_reg8[25]), .C0(n228), .C1(result_reg8[9]), .Y(n433) );
  INVX1 U453 ( .A(n432), .Y(n70) );
  AOI222X1 U454 ( .A0(n224), .A1(cal_result[10]), .B0(n218), .B1(
        result_reg8[26]), .C0(n228), .C1(result_reg8[10]), .Y(n432) );
  INVX1 U455 ( .A(n431), .Y(n69) );
  AOI222X1 U456 ( .A0(n224), .A1(cal_result[11]), .B0(n218), .B1(
        result_reg8[27]), .C0(n228), .C1(result_reg8[11]), .Y(n431) );
  INVX1 U457 ( .A(n430), .Y(n68) );
  AOI222X1 U458 ( .A0(n224), .A1(cal_result[12]), .B0(n218), .B1(
        result_reg8[28]), .C0(n228), .C1(result_reg8[12]), .Y(n430) );
  INVX1 U459 ( .A(n426), .Y(n64) );
  AOI222X1 U460 ( .A0(n224), .A1(cal_result[16]), .B0(n217), .B1(
        result_reg8[32]), .C0(n228), .C1(result_reg8[16]), .Y(n426) );
  INVX1 U461 ( .A(n425), .Y(n63) );
  AOI222X1 U462 ( .A0(n224), .A1(cal_result[17]), .B0(n217), .B1(
        result_reg8[33]), .C0(n228), .C1(result_reg8[17]), .Y(n425) );
  INVX1 U463 ( .A(n424), .Y(n62) );
  AOI222X1 U464 ( .A0(n224), .A1(cal_result[18]), .B0(n217), .B1(
        result_reg8[34]), .C0(n228), .C1(result_reg8[18]), .Y(n424) );
  INVX1 U465 ( .A(n423), .Y(n61) );
  AOI222X1 U466 ( .A0(n224), .A1(cal_result[19]), .B0(n217), .B1(
        result_reg8[35]), .C0(n228), .C1(result_reg8[19]), .Y(n423) );
  INVX1 U467 ( .A(n422), .Y(n60) );
  AOI222X1 U468 ( .A0(n224), .A1(cal_result[20]), .B0(n217), .B1(
        result_reg8[36]), .C0(n228), .C1(result_reg8[20]), .Y(n422) );
  INVX1 U469 ( .A(n421), .Y(n59) );
  AOI222X1 U470 ( .A0(n224), .A1(cal_result[21]), .B0(n217), .B1(
        result_reg8[37]), .C0(n228), .C1(result_reg8[21]), .Y(n421) );
  INVX1 U471 ( .A(n420), .Y(n58) );
  AOI222X1 U472 ( .A0(n224), .A1(cal_result[22]), .B0(n217), .B1(
        result_reg8[38]), .C0(n228), .C1(result_reg8[22]), .Y(n420) );
  INVX1 U473 ( .A(n419), .Y(n57) );
  AOI222X1 U474 ( .A0(n224), .A1(cal_result[23]), .B0(n217), .B1(
        result_reg8[39]), .C0(n228), .C1(result_reg8[23]), .Y(n419) );
  INVX1 U475 ( .A(n418), .Y(n56) );
  AOI222X1 U476 ( .A0(n224), .A1(cal_result[24]), .B0(n217), .B1(
        result_reg8[40]), .C0(n228), .C1(result_reg8[24]), .Y(n418) );
  INVX1 U477 ( .A(n417), .Y(n55) );
  AOI222X1 U478 ( .A0(n224), .A1(cal_result[25]), .B0(n217), .B1(
        result_reg8[41]), .C0(n228), .C1(result_reg8[25]), .Y(n417) );
  INVX1 U479 ( .A(n416), .Y(n54) );
  AOI222X1 U480 ( .A0(n224), .A1(cal_result[26]), .B0(n217), .B1(
        result_reg8[42]), .C0(n228), .C1(result_reg8[26]), .Y(n416) );
  INVX1 U481 ( .A(n415), .Y(n53) );
  AOI222X1 U482 ( .A0(n224), .A1(cal_result[27]), .B0(n217), .B1(
        result_reg8[43]), .C0(n228), .C1(result_reg8[27]), .Y(n415) );
  INVX1 U483 ( .A(n414), .Y(n52) );
  AOI222X1 U484 ( .A0(n224), .A1(cal_result[28]), .B0(n217), .B1(
        result_reg8[44]), .C0(n228), .C1(result_reg8[28]), .Y(n414) );
  INVX1 U485 ( .A(n410), .Y(n48) );
  AOI222X1 U486 ( .A0(n224), .A1(cal_result[32]), .B0(n217), .B1(
        result_reg8[48]), .C0(n227), .C1(result_reg8[32]), .Y(n410) );
  INVX1 U487 ( .A(n409), .Y(n47) );
  AOI222X1 U488 ( .A0(n224), .A1(cal_result[33]), .B0(n217), .B1(
        result_reg8[49]), .C0(n227), .C1(result_reg8[33]), .Y(n409) );
  INVX1 U489 ( .A(n408), .Y(n46) );
  AOI222X1 U490 ( .A0(n224), .A1(cal_result[34]), .B0(n217), .B1(
        result_reg8[50]), .C0(n227), .C1(result_reg8[34]), .Y(n408) );
  INVX1 U491 ( .A(n407), .Y(n45) );
  AOI222X1 U492 ( .A0(n224), .A1(cal_result[35]), .B0(n217), .B1(
        result_reg8[51]), .C0(n227), .C1(result_reg8[35]), .Y(n407) );
  INVX1 U493 ( .A(n406), .Y(n44) );
  AOI222X1 U494 ( .A0(n223), .A1(cal_result[36]), .B0(n217), .B1(
        result_reg8[52]), .C0(n227), .C1(result_reg8[36]), .Y(n406) );
  INVX1 U495 ( .A(n405), .Y(n43) );
  AOI222X1 U496 ( .A0(n223), .A1(cal_result[37]), .B0(n217), .B1(
        result_reg8[53]), .C0(n227), .C1(result_reg8[37]), .Y(n405) );
  INVX1 U497 ( .A(n404), .Y(n42) );
  AOI222X1 U498 ( .A0(n223), .A1(cal_result[38]), .B0(n217), .B1(
        result_reg8[54]), .C0(n227), .C1(result_reg8[38]), .Y(n404) );
  INVX1 U499 ( .A(n403), .Y(n41) );
  AOI222X1 U500 ( .A0(n223), .A1(cal_result[39]), .B0(n217), .B1(
        result_reg8[55]), .C0(n227), .C1(result_reg8[39]), .Y(n403) );
  INVX1 U501 ( .A(n402), .Y(n40) );
  AOI222X1 U502 ( .A0(n223), .A1(cal_result[40]), .B0(n217), .B1(
        result_reg8[56]), .C0(n227), .C1(result_reg8[40]), .Y(n402) );
  INVX1 U503 ( .A(n401), .Y(n39) );
  AOI222X1 U504 ( .A0(n223), .A1(cal_result[41]), .B0(n217), .B1(
        result_reg8[57]), .C0(n227), .C1(result_reg8[41]), .Y(n401) );
  INVX1 U505 ( .A(n400), .Y(n38) );
  AOI222X1 U506 ( .A0(n223), .A1(cal_result[42]), .B0(n217), .B1(
        result_reg8[58]), .C0(n227), .C1(result_reg8[42]), .Y(n400) );
  INVX1 U507 ( .A(n399), .Y(n37) );
  AOI222X1 U508 ( .A0(n223), .A1(cal_result[43]), .B0(n217), .B1(
        result_reg8[59]), .C0(n227), .C1(result_reg8[43]), .Y(n399) );
  INVX1 U509 ( .A(n398), .Y(n36) );
  AOI222X1 U510 ( .A0(n223), .A1(cal_result[44]), .B0(n217), .B1(
        result_reg8[60]), .C0(n227), .C1(result_reg8[44]), .Y(n398) );
  INVX1 U511 ( .A(n394), .Y(n32) );
  AOI222X1 U512 ( .A0(n223), .A1(cal_result[48]), .B0(n216), .B1(
        result_reg8[64]), .C0(n227), .C1(result_reg8[48]), .Y(n394) );
  INVX1 U513 ( .A(n393), .Y(n31) );
  AOI222X1 U514 ( .A0(n223), .A1(cal_result[49]), .B0(n218), .B1(
        result_reg8[65]), .C0(n227), .C1(result_reg8[49]), .Y(n393) );
  INVX1 U515 ( .A(n392), .Y(n30) );
  AOI222X1 U516 ( .A0(n223), .A1(cal_result[50]), .B0(n216), .B1(
        result_reg8[66]), .C0(n227), .C1(result_reg8[50]), .Y(n392) );
  INVX1 U517 ( .A(n391), .Y(n29) );
  AOI222X1 U518 ( .A0(n223), .A1(cal_result[51]), .B0(n218), .B1(
        result_reg8[67]), .C0(n227), .C1(result_reg8[51]), .Y(n391) );
  INVX1 U519 ( .A(n390), .Y(n28) );
  AOI222X1 U520 ( .A0(n223), .A1(cal_result[52]), .B0(n216), .B1(
        result_reg8[68]), .C0(n227), .C1(result_reg8[52]), .Y(n390) );
  INVX1 U521 ( .A(n389), .Y(n27) );
  AOI222X1 U522 ( .A0(n223), .A1(cal_result[53]), .B0(n218), .B1(
        result_reg8[69]), .C0(n227), .C1(result_reg8[53]), .Y(n389) );
  INVX1 U523 ( .A(n388), .Y(n26) );
  AOI222X1 U524 ( .A0(n223), .A1(cal_result[54]), .B0(n216), .B1(
        result_reg8[70]), .C0(n227), .C1(result_reg8[54]), .Y(n388) );
  INVX1 U525 ( .A(n387), .Y(n25) );
  AOI222X1 U526 ( .A0(n223), .A1(cal_result[55]), .B0(n218), .B1(
        result_reg8[71]), .C0(n227), .C1(result_reg8[55]), .Y(n387) );
  INVX1 U527 ( .A(n386), .Y(n24) );
  AOI222X1 U528 ( .A0(n223), .A1(cal_result[56]), .B0(n331), .B1(
        result_reg8[72]), .C0(n227), .C1(result_reg8[56]), .Y(n386) );
  INVX1 U529 ( .A(n385), .Y(n23) );
  AOI222X1 U530 ( .A0(n223), .A1(cal_result[57]), .B0(n331), .B1(
        result_reg8[73]), .C0(n227), .C1(result_reg8[57]), .Y(n385) );
  INVX1 U531 ( .A(n384), .Y(n22) );
  AOI222X1 U532 ( .A0(n223), .A1(cal_result[58]), .B0(n331), .B1(
        result_reg8[74]), .C0(n227), .C1(result_reg8[58]), .Y(n384) );
  INVX1 U533 ( .A(n383), .Y(n21) );
  AOI222X1 U534 ( .A0(n223), .A1(cal_result[59]), .B0(n331), .B1(
        result_reg8[75]), .C0(n227), .C1(result_reg8[59]), .Y(n383) );
  INVX1 U535 ( .A(n382), .Y(n20) );
  AOI222X1 U536 ( .A0(n223), .A1(cal_result[60]), .B0(n331), .B1(
        result_reg8[76]), .C0(n227), .C1(result_reg8[60]), .Y(n382) );
  BUFX3 U537 ( .A(n289), .Y(n86) );
  OAI21XL U538 ( .A0(n306), .A1(mode_reg_0_), .B0(n309), .Y(n289) );
  OAI2BB2X1 U539 ( .B0(n82), .B1(n288), .A0N(dout[0]), .A1N(n82), .Y(n516) );
  AOI22X1 U540 ( .A0(result_reg4[0]), .A1(n86), .B0(result_reg8[0]), .B1(n85), 
        .Y(n288) );
  OAI2BB2X1 U541 ( .B0(n82), .B1(n291), .A0N(dout[1]), .A1N(n82), .Y(n517) );
  AOI22X1 U542 ( .A0(result_reg4[1]), .A1(n86), .B0(result_reg8[1]), .B1(n85), 
        .Y(n291) );
  OAI2BB2X1 U543 ( .B0(n82), .B1(n292), .A0N(dout[2]), .A1N(n82), .Y(n518) );
  AOI22X1 U544 ( .A0(result_reg4[2]), .A1(n86), .B0(result_reg8[2]), .B1(n85), 
        .Y(n292) );
  OAI2BB2X1 U545 ( .B0(n82), .B1(n293), .A0N(dout[3]), .A1N(n82), .Y(n519) );
  AOI22X1 U546 ( .A0(result_reg4[3]), .A1(n86), .B0(result_reg8[3]), .B1(n85), 
        .Y(n293) );
  OAI2BB2X1 U547 ( .B0(n82), .B1(n294), .A0N(dout[4]), .A1N(n82), .Y(n520) );
  AOI22X1 U548 ( .A0(result_reg4[4]), .A1(n86), .B0(result_reg8[4]), .B1(n85), 
        .Y(n294) );
  OAI2BB2X1 U549 ( .B0(n82), .B1(n295), .A0N(dout[5]), .A1N(n82), .Y(n521) );
  AOI22X1 U550 ( .A0(result_reg4[5]), .A1(n86), .B0(result_reg8[5]), .B1(n85), 
        .Y(n295) );
  OAI2BB2X1 U551 ( .B0(n82), .B1(n296), .A0N(dout[6]), .A1N(n82), .Y(n522) );
  AOI22X1 U552 ( .A0(result_reg4[6]), .A1(n86), .B0(result_reg8[6]), .B1(n85), 
        .Y(n296) );
  OAI2BB2X1 U553 ( .B0(n82), .B1(n297), .A0N(dout[7]), .A1N(n82), .Y(n523) );
  AOI22X1 U554 ( .A0(result_reg4[7]), .A1(n86), .B0(result_reg8[7]), .B1(n85), 
        .Y(n297) );
  OAI2BB2X1 U555 ( .B0(n82), .B1(n298), .A0N(dout[8]), .A1N(n82), .Y(n524) );
  AOI22X1 U556 ( .A0(result_reg4[8]), .A1(n86), .B0(result_reg8[8]), .B1(n85), 
        .Y(n298) );
  OAI2BB2X1 U557 ( .B0(n82), .B1(n299), .A0N(dout[9]), .A1N(n82), .Y(n525) );
  AOI22X1 U558 ( .A0(result_reg4[9]), .A1(n86), .B0(result_reg8[9]), .B1(n85), 
        .Y(n299) );
  OAI2BB2X1 U559 ( .B0(n82), .B1(n300), .A0N(dout[10]), .A1N(n82), .Y(n526) );
  AOI22X1 U560 ( .A0(result_reg4[10]), .A1(n86), .B0(result_reg8[10]), .B1(n85), .Y(n300) );
  OAI2BB2X1 U561 ( .B0(n82), .B1(n301), .A0N(dout[11]), .A1N(n82), .Y(n527) );
  AOI22X1 U562 ( .A0(result_reg4[11]), .A1(n86), .B0(result_reg8[11]), .B1(n85), .Y(n301) );
  OAI2BB2X1 U563 ( .B0(n82), .B1(n302), .A0N(dout[12]), .A1N(n82), .Y(n528) );
  AOI22X1 U564 ( .A0(result_reg4[12]), .A1(n86), .B0(result_reg8[12]), .B1(n85), .Y(n302) );
  OAI2BB2X1 U565 ( .B0(n82), .B1(n303), .A0N(dout[13]), .A1N(n82), .Y(n529) );
  AOI22X1 U566 ( .A0(result_reg4[13]), .A1(n86), .B0(result_reg8[13]), .B1(n85), .Y(n303) );
  OAI2BB2X1 U567 ( .B0(n82), .B1(n304), .A0N(dout[14]), .A1N(n82), .Y(n530) );
  AOI22X1 U568 ( .A0(result_reg4[14]), .A1(n86), .B0(result_reg8[14]), .B1(n85), .Y(n304) );
  OAI2BB2X1 U569 ( .B0(n82), .B1(n305), .A0N(dout[15]), .A1N(n82), .Y(n531) );
  AOI22X1 U570 ( .A0(result_reg4[15]), .A1(n86), .B0(result_reg8[15]), .B1(n85), .Y(n305) );
  BUFX3 U571 ( .A(n290), .Y(n85) );
  OAI21XL U572 ( .A0(n306), .A1(n745), .B0(n308), .Y(n290) );
  INVX1 U573 ( .A(mode_reg_0_), .Y(n745) );
  INVX1 U574 ( .A(shift4_flag), .Y(n673) );
  OAI2BB1X1 U575 ( .A0N(n226), .A1N(result_reg8[68]), .B0(n374), .Y(n576) );
  AOI22X1 U576 ( .A0(result_reg8[84]), .A1(n218), .B0(cal_result[68]), .B1(
        n222), .Y(n374) );
  OAI2BB1X1 U577 ( .A0N(n226), .A1N(result_reg8[69]), .B0(n373), .Y(n575) );
  AOI22X1 U578 ( .A0(result_reg8[85]), .A1(n216), .B0(cal_result[69]), .B1(
        n220), .Y(n373) );
  OAI2BB1X1 U579 ( .A0N(n226), .A1N(result_reg8[70]), .B0(n372), .Y(n574) );
  AOI22X1 U580 ( .A0(result_reg8[86]), .A1(n216), .B0(cal_result[70]), .B1(
        n222), .Y(n372) );
  OAI2BB1X1 U581 ( .A0N(n226), .A1N(result_reg8[71]), .B0(n371), .Y(n573) );
  AOI22X1 U582 ( .A0(result_reg8[87]), .A1(n218), .B0(cal_result[71]), .B1(
        n220), .Y(n371) );
  OAI2BB1X1 U583 ( .A0N(n226), .A1N(result_reg8[72]), .B0(n370), .Y(n572) );
  AOI22X1 U584 ( .A0(result_reg8[88]), .A1(n216), .B0(cal_result[72]), .B1(
        n220), .Y(n370) );
  OAI2BB1X1 U585 ( .A0N(n226), .A1N(result_reg8[73]), .B0(n369), .Y(n571) );
  AOI22X1 U586 ( .A0(result_reg8[89]), .A1(n216), .B0(cal_result[73]), .B1(
        n222), .Y(n369) );
  OAI2BB1X1 U587 ( .A0N(n226), .A1N(result_reg8[74]), .B0(n368), .Y(n570) );
  AOI22X1 U588 ( .A0(result_reg8[90]), .A1(n216), .B0(cal_result[74]), .B1(
        n220), .Y(n368) );
  OAI2BB1X1 U589 ( .A0N(n226), .A1N(result_reg8[75]), .B0(n367), .Y(n569) );
  AOI22X1 U590 ( .A0(result_reg8[91]), .A1(n218), .B0(cal_result[75]), .B1(
        n222), .Y(n367) );
  OAI2BB1X1 U591 ( .A0N(n226), .A1N(result_reg8[76]), .B0(n366), .Y(n568) );
  AOI22X1 U592 ( .A0(result_reg8[92]), .A1(n218), .B0(cal_result[76]), .B1(
        n220), .Y(n366) );
  OAI2BB1X1 U593 ( .A0N(n226), .A1N(result_reg8[80]), .B0(n362), .Y(n564) );
  AOI22X1 U594 ( .A0(result_reg8[96]), .A1(n216), .B0(cal_result[80]), .B1(
        n220), .Y(n362) );
  OAI2BB1X1 U595 ( .A0N(n226), .A1N(result_reg8[81]), .B0(n361), .Y(n563) );
  AOI22X1 U596 ( .A0(result_reg8[97]), .A1(n218), .B0(cal_result[81]), .B1(
        n220), .Y(n361) );
  OAI2BB1X1 U597 ( .A0N(n226), .A1N(result_reg8[82]), .B0(n360), .Y(n562) );
  AOI22X1 U598 ( .A0(result_reg8[98]), .A1(n216), .B0(cal_result[82]), .B1(
        n220), .Y(n360) );
  OAI2BB1X1 U599 ( .A0N(n226), .A1N(result_reg8[83]), .B0(n359), .Y(n561) );
  AOI22X1 U600 ( .A0(result_reg8[99]), .A1(n216), .B0(cal_result[83]), .B1(
        n222), .Y(n359) );
  OAI2BB1X1 U601 ( .A0N(n226), .A1N(result_reg8[84]), .B0(n358), .Y(n560) );
  AOI22X1 U602 ( .A0(result_reg8[100]), .A1(n216), .B0(cal_result[84]), .B1(
        n222), .Y(n358) );
  OAI2BB1X1 U603 ( .A0N(n226), .A1N(result_reg8[85]), .B0(n357), .Y(n559) );
  AOI22X1 U604 ( .A0(result_reg8[101]), .A1(n216), .B0(cal_result[85]), .B1(
        n222), .Y(n357) );
  OAI2BB1X1 U605 ( .A0N(n226), .A1N(result_reg8[86]), .B0(n356), .Y(n558) );
  AOI22X1 U606 ( .A0(result_reg8[102]), .A1(n218), .B0(cal_result[86]), .B1(
        n222), .Y(n356) );
  OAI2BB1X1 U607 ( .A0N(n226), .A1N(result_reg8[87]), .B0(n355), .Y(n557) );
  AOI22X1 U608 ( .A0(result_reg8[103]), .A1(n216), .B0(cal_result[87]), .B1(
        n220), .Y(n355) );
  OAI2BB1X1 U609 ( .A0N(n226), .A1N(result_reg8[88]), .B0(n354), .Y(n556) );
  AOI22X1 U610 ( .A0(result_reg8[104]), .A1(n216), .B0(cal_result[88]), .B1(
        n222), .Y(n354) );
  OAI2BB1X1 U611 ( .A0N(n226), .A1N(result_reg8[89]), .B0(n353), .Y(n555) );
  AOI22X1 U612 ( .A0(result_reg8[105]), .A1(n216), .B0(cal_result[89]), .B1(
        n222), .Y(n353) );
  OAI2BB1X1 U613 ( .A0N(n225), .A1N(result_reg8[90]), .B0(n352), .Y(n554) );
  AOI22X1 U614 ( .A0(result_reg8[106]), .A1(n216), .B0(cal_result[90]), .B1(
        n222), .Y(n352) );
  OAI2BB1X1 U615 ( .A0N(n226), .A1N(result_reg8[91]), .B0(n351), .Y(n553) );
  AOI22X1 U616 ( .A0(result_reg8[107]), .A1(n216), .B0(cal_result[91]), .B1(
        n220), .Y(n351) );
  OAI2BB1X1 U617 ( .A0N(n226), .A1N(result_reg8[92]), .B0(n350), .Y(n552) );
  AOI22X1 U618 ( .A0(result_reg8[108]), .A1(n216), .B0(cal_result[92]), .B1(
        n222), .Y(n350) );
  OAI2BB1X1 U619 ( .A0N(n225), .A1N(result_reg8[96]), .B0(n346), .Y(n548) );
  AOI22X1 U620 ( .A0(n216), .A1(result_reg8[112]), .B0(cal_result[96]), .B1(
        n222), .Y(n346) );
  OAI2BB1X1 U621 ( .A0N(n225), .A1N(result_reg8[97]), .B0(n345), .Y(n547) );
  AOI22X1 U622 ( .A0(n331), .A1(result_reg8[113]), .B0(cal_result[97]), .B1(
        n222), .Y(n345) );
  OAI2BB1X1 U623 ( .A0N(n225), .A1N(result_reg8[98]), .B0(n344), .Y(n546) );
  AOI22X1 U624 ( .A0(n216), .A1(result_reg8[114]), .B0(cal_result[98]), .B1(
        n222), .Y(n344) );
  OAI2BB1X1 U625 ( .A0N(n225), .A1N(result_reg8[99]), .B0(n343), .Y(n545) );
  AOI22X1 U626 ( .A0(n331), .A1(result_reg8[115]), .B0(cal_result[99]), .B1(
        n222), .Y(n343) );
  OAI2BB1X1 U627 ( .A0N(n225), .A1N(result_reg8[100]), .B0(n342), .Y(n544) );
  AOI22X1 U628 ( .A0(n216), .A1(result_reg8[116]), .B0(cal_result[100]), .B1(
        n222), .Y(n342) );
  OAI2BB1X1 U629 ( .A0N(n225), .A1N(result_reg8[101]), .B0(n341), .Y(n543) );
  AOI22X1 U630 ( .A0(n331), .A1(result_reg8[117]), .B0(cal_result[101]), .B1(
        n222), .Y(n341) );
  OAI2BB1X1 U631 ( .A0N(n225), .A1N(result_reg8[102]), .B0(n340), .Y(n542) );
  AOI22X1 U632 ( .A0(n331), .A1(result_reg8[118]), .B0(cal_result[102]), .B1(
        n222), .Y(n340) );
  OAI2BB1X1 U633 ( .A0N(n225), .A1N(result_reg8[103]), .B0(n339), .Y(n541) );
  AOI22X1 U634 ( .A0(n331), .A1(result_reg8[119]), .B0(cal_result[103]), .B1(
        n222), .Y(n339) );
  OAI2BB1X1 U635 ( .A0N(n225), .A1N(result_reg8[104]), .B0(n338), .Y(n540) );
  AOI22X1 U636 ( .A0(n216), .A1(result_reg8[120]), .B0(cal_result[104]), .B1(
        n220), .Y(n338) );
  OAI2BB1X1 U637 ( .A0N(n225), .A1N(result_reg8[105]), .B0(n337), .Y(n539) );
  AOI22X1 U638 ( .A0(n331), .A1(result_reg8[121]), .B0(cal_result[105]), .B1(
        n220), .Y(n337) );
  OAI2BB1X1 U639 ( .A0N(n225), .A1N(result_reg8[106]), .B0(n336), .Y(n538) );
  AOI22X1 U640 ( .A0(n218), .A1(result_reg8[122]), .B0(cal_result[106]), .B1(
        n220), .Y(n336) );
  OAI2BB1X1 U641 ( .A0N(n225), .A1N(result_reg8[107]), .B0(n335), .Y(n537) );
  AOI22X1 U642 ( .A0(n331), .A1(result_reg8[123]), .B0(cal_result[107]), .B1(
        n220), .Y(n335) );
  OAI2BB1X1 U643 ( .A0N(n225), .A1N(result_reg8[108]), .B0(n334), .Y(n536) );
  AOI22X1 U644 ( .A0(n216), .A1(result_reg8[124]), .B0(cal_result[108]), .B1(
        n220), .Y(n334) );
  OAI2BB1X1 U645 ( .A0N(n226), .A1N(result_reg8[64]), .B0(n378), .Y(n580) );
  AOI22X1 U646 ( .A0(result_reg8[80]), .A1(n216), .B0(cal_result[64]), .B1(
        n223), .Y(n378) );
  OAI2BB1X1 U647 ( .A0N(n226), .A1N(result_reg8[65]), .B0(n377), .Y(n579) );
  AOI22X1 U648 ( .A0(result_reg8[81]), .A1(n218), .B0(cal_result[65]), .B1(
        n223), .Y(n377) );
  OAI2BB1X1 U649 ( .A0N(n226), .A1N(result_reg8[66]), .B0(n376), .Y(n578) );
  AOI22X1 U650 ( .A0(result_reg8[82]), .A1(n218), .B0(cal_result[66]), .B1(
        n223), .Y(n376) );
  OAI2BB1X1 U651 ( .A0N(n226), .A1N(result_reg8[67]), .B0(n375), .Y(n577) );
  AOI22X1 U652 ( .A0(result_reg8[83]), .A1(n218), .B0(cal_result[67]), .B1(
        n223), .Y(n375) );
  INVX1 U653 ( .A(n329), .Y(n16) );
  AOI22X1 U654 ( .A0(n225), .A1(result_reg8[112]), .B0(cal_result[112]), .B1(
        n220), .Y(n329) );
  INVX1 U655 ( .A(n328), .Y(n15) );
  AOI22X1 U656 ( .A0(n225), .A1(result_reg8[113]), .B0(cal_result[113]), .B1(
        n220), .Y(n328) );
  INVX1 U657 ( .A(n327), .Y(n14) );
  AOI22X1 U658 ( .A0(n225), .A1(result_reg8[114]), .B0(cal_result[114]), .B1(
        n220), .Y(n327) );
  INVX1 U659 ( .A(n326), .Y(n13) );
  AOI22X1 U660 ( .A0(n225), .A1(result_reg8[115]), .B0(cal_result[115]), .B1(
        n220), .Y(n326) );
  INVX1 U661 ( .A(n325), .Y(n12) );
  AOI22X1 U662 ( .A0(n225), .A1(result_reg8[116]), .B0(cal_result[116]), .B1(
        n220), .Y(n325) );
  INVX1 U663 ( .A(n324), .Y(n11) );
  AOI22X1 U664 ( .A0(n311), .A1(result_reg8[117]), .B0(cal_result[117]), .B1(
        n220), .Y(n324) );
  INVX1 U665 ( .A(n323), .Y(n10) );
  AOI22X1 U666 ( .A0(n311), .A1(result_reg8[118]), .B0(cal_result[118]), .B1(
        n222), .Y(n323) );
  INVX1 U667 ( .A(n322), .Y(n9) );
  AOI22X1 U668 ( .A0(n311), .A1(result_reg8[119]), .B0(cal_result[119]), .B1(
        n222), .Y(n322) );
  INVX1 U669 ( .A(n321), .Y(n8) );
  AOI22X1 U670 ( .A0(n311), .A1(result_reg8[120]), .B0(cal_result[120]), .B1(
        n220), .Y(n321) );
  INVX1 U671 ( .A(n320), .Y(n7) );
  AOI22X1 U672 ( .A0(n311), .A1(result_reg8[121]), .B0(cal_result[121]), .B1(
        n222), .Y(n320) );
  INVX1 U673 ( .A(n319), .Y(n6) );
  AOI22X1 U674 ( .A0(n311), .A1(result_reg8[122]), .B0(cal_result[122]), .B1(
        n220), .Y(n319) );
  INVX1 U675 ( .A(n318), .Y(n5) );
  AOI22X1 U676 ( .A0(n311), .A1(result_reg8[123]), .B0(cal_result[123]), .B1(
        n220), .Y(n318) );
  INVX1 U677 ( .A(n317), .Y(n4) );
  AOI22X1 U678 ( .A0(n311), .A1(result_reg8[124]), .B0(cal_result[124]), .B1(
        n222), .Y(n317) );
  OAI2BB2X1 U679 ( .B0(n674), .B1(n515), .A0N(n515), .A1N(start), .Y(n668) );
  OAI2BB1X1 U680 ( .A0N(mode[0]), .A1N(n444), .B0(n312), .Y(n515) );
  OAI2BB1X1 U681 ( .A0N(n309), .A1N(mode_reg_0_), .B0(n312), .Y(n532) );
  INVX1 U682 ( .A(result_reg4[128]), .Y(n696) );
  INVX1 U683 ( .A(result_reg4[129]), .Y(n695) );
  INVX1 U684 ( .A(result_reg4[130]), .Y(n694) );
  INVX1 U685 ( .A(result_reg4[131]), .Y(n693) );
  INVX1 U686 ( .A(result_reg4[132]), .Y(n692) );
  INVX1 U687 ( .A(result_reg4[133]), .Y(n691) );
  INVX1 U688 ( .A(result_reg4[134]), .Y(n690) );
  INVX1 U689 ( .A(result_reg4[135]), .Y(n689) );
  INVX1 U690 ( .A(result_reg4[136]), .Y(n688) );
  INVX1 U691 ( .A(result_reg4[137]), .Y(n687) );
  INVX1 U692 ( .A(result_reg4[138]), .Y(n686) );
  INVX1 U693 ( .A(result_reg4[139]), .Y(n685) );
  INVX1 U694 ( .A(result_reg4[140]), .Y(n684) );
  INVX1 U695 ( .A(result_reg4[141]), .Y(n683) );
  INVX1 U696 ( .A(result_reg4[142]), .Y(n682) );
  INVX1 U697 ( .A(result_reg4[143]), .Y(n681) );
  INVX1 U698 ( .A(result_reg4[96]), .Y(n728) );
  INVX1 U699 ( .A(result_reg4[97]), .Y(n727) );
  INVX1 U700 ( .A(result_reg4[98]), .Y(n726) );
  INVX1 U701 ( .A(result_reg4[99]), .Y(n725) );
  INVX1 U702 ( .A(result_reg4[100]), .Y(n724) );
  INVX1 U703 ( .A(result_reg4[101]), .Y(n723) );
  INVX1 U704 ( .A(result_reg4[102]), .Y(n722) );
  INVX1 U705 ( .A(result_reg4[103]), .Y(n721) );
  INVX1 U706 ( .A(result_reg4[104]), .Y(n720) );
  INVX1 U707 ( .A(result_reg4[105]), .Y(n719) );
  INVX1 U708 ( .A(result_reg4[106]), .Y(n718) );
  INVX1 U709 ( .A(result_reg4[107]), .Y(n717) );
  INVX1 U710 ( .A(result_reg4[108]), .Y(n716) );
  INVX1 U711 ( .A(result_reg4[109]), .Y(n715) );
  INVX1 U712 ( .A(result_reg4[110]), .Y(n714) );
  INVX1 U713 ( .A(result_reg4[111]), .Y(n713) );
  INVX1 U714 ( .A(result_reg4[112]), .Y(n712) );
  INVX1 U715 ( .A(result_reg4[113]), .Y(n711) );
  INVX1 U716 ( .A(result_reg4[114]), .Y(n710) );
  INVX1 U717 ( .A(result_reg4[115]), .Y(n709) );
  INVX1 U718 ( .A(result_reg4[116]), .Y(n708) );
  INVX1 U719 ( .A(result_reg4[117]), .Y(n707) );
  INVX1 U720 ( .A(result_reg4[118]), .Y(n706) );
  INVX1 U721 ( .A(result_reg4[119]), .Y(n705) );
  INVX1 U722 ( .A(result_reg4[120]), .Y(n704) );
  INVX1 U723 ( .A(result_reg4[121]), .Y(n703) );
  INVX1 U724 ( .A(result_reg4[122]), .Y(n702) );
  INVX1 U725 ( .A(result_reg4[123]), .Y(n701) );
  INVX1 U726 ( .A(result_reg4[124]), .Y(n700) );
  INVX1 U727 ( .A(result_reg4[125]), .Y(n699) );
  INVX1 U728 ( .A(result_reg4[126]), .Y(n698) );
  INVX1 U729 ( .A(result_reg4[127]), .Y(n697) );
  INVX1 U730 ( .A(start_reg4[1]), .Y(n679) );
  INVX1 U731 ( .A(start_reg4[2]), .Y(n678) );
  INVX1 U732 ( .A(start_reg4[3]), .Y(n677) );
  INVX1 U733 ( .A(start_reg4[4]), .Y(n676) );
  INVX1 U734 ( .A(start_reg4[5]), .Y(n675) );
  INVX1 U735 ( .A(result_reg4[80]), .Y(n744) );
  INVX1 U736 ( .A(result_reg4[81]), .Y(n743) );
  INVX1 U737 ( .A(result_reg4[82]), .Y(n742) );
  INVX1 U738 ( .A(result_reg4[83]), .Y(n741) );
  INVX1 U739 ( .A(result_reg4[84]), .Y(n740) );
  INVX1 U740 ( .A(result_reg4[85]), .Y(n739) );
  INVX1 U741 ( .A(result_reg4[86]), .Y(n738) );
  INVX1 U742 ( .A(result_reg4[87]), .Y(n737) );
  INVX1 U743 ( .A(result_reg4[88]), .Y(n736) );
  INVX1 U744 ( .A(result_reg4[89]), .Y(n735) );
  INVX1 U745 ( .A(result_reg4[90]), .Y(n734) );
  INVX1 U746 ( .A(result_reg4[91]), .Y(n733) );
  INVX1 U747 ( .A(result_reg4[92]), .Y(n732) );
  INVX1 U748 ( .A(result_reg4[93]), .Y(n731) );
  INVX1 U749 ( .A(result_reg4[94]), .Y(n730) );
  INVX1 U750 ( .A(result_reg4[95]), .Y(n729) );
endmodule


module mem_ctrl_tran_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  XOR2X1 U1 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module mem_ctrl_tran_DW01_inc_5 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  ADDHXL U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  XOR2X1 U1 ( .A(carry[8]), .B(A[8]), .Y(SUM[8]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module mem_ctrl_tran_DW01_inc_4 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  ADDHXL U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  XOR2X1 U1 ( .A(carry[8]), .B(A[8]), .Y(SUM[8]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module mem_ctrl_tran_DW01_inc_3 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  ADDHXL U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  XOR2X1 U1 ( .A(carry[8]), .B(A[8]), .Y(SUM[8]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module mem_ctrl_tran_DW01_inc_2 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  ADDHXL U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  XOR2X1 U1 ( .A(carry[8]), .B(A[8]), .Y(SUM[8]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module mem_ctrl_tran_DW01_inc_1 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  ADDHXL U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  XOR2X1 U1 ( .A(carry[8]), .B(A[8]), .Y(SUM[8]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module mem_ctrl_tran ( clk, rstn, start, mode, en_ram8x8_1, wr_rd_ram8x8_1, 
        addr_ram8x8_1, en_ram8x8_2, wr_rd_ram8x8_2, addr_ram8x8_2, en_ram4x4_1, 
        wr_rd_ram4x4_1, addr_ram4x4_1, en_ram4x4_2, wr_rd_ram4x4_2, 
        addr_ram4x4_2, en_ram4x4_3, wr_rd_ram4x4_3, addr_ram4x4_3, en_ram4x4_4, 
        wr_rd_ram4x4_4, addr_ram4x4_4, ram8x8_1_ready, ram8x8_2_ready, 
        ram4x4_1_ready, ram4x4_2_ready, ram4x4_3_ready, ram4x4_4_ready, 
        mode_out );
  input [1:0] mode;
  output [5:0] addr_ram8x8_1;
  output [5:0] addr_ram8x8_2;
  output [3:0] addr_ram4x4_1;
  output [3:0] addr_ram4x4_2;
  output [3:0] addr_ram4x4_3;
  output [3:0] addr_ram4x4_4;
  output [1:0] mode_out;
  input clk, rstn, start;
  output en_ram8x8_1, wr_rd_ram8x8_1, en_ram8x8_2, wr_rd_ram8x8_2, en_ram4x4_1,
         wr_rd_ram4x4_1, en_ram4x4_2, wr_rd_ram4x4_2, en_ram4x4_3,
         wr_rd_ram4x4_3, en_ram4x4_4, wr_rd_ram4x4_4, ram8x8_1_ready,
         ram8x8_2_ready, ram4x4_1_ready, ram4x4_2_ready, ram4x4_3_ready,
         ram4x4_4_ready;
  wire   coeff_shift_w_0_, mode_r_0_, coeff_shift_r_0_, ram_write_reg,
         ram_write, ram, ram8x8_w_ready, en_ram8x8_w, wr_rd_ram8x8_w,
         ram8x8_r_ready, en_ram8x8_r, count_r2_3_, ram8_4, N329, N330, N331,
         N593, N716, N717, N718, N724, N725, N726, N727, N728, N729, N730,
         N731, N732, N737, N738, N739, N749, N750, N751, N752, N758, N760,
         N761, N762, N763, N764, N765, N766, N767, N780, N782, N783, N805,
         N807, N808, N824, N825, N826, N827, N828, N830, N831, N832, N833,
         N834, N835, N836, N837, N851, N852, N853, N854, N855, N856, N857,
         N858, N859, N979, N980, N981, N982, N983, N984, N985, N986, N987,
         N1067, N1068, N1069, N1070, N1071, N1074, N1075, N1076, N1077, N1078,
         N1079, N1361, N1362, N1363, N1364, N1365, N1366, N1367, N1368, N1369,
         N1399, N1400, N1401, N1402, N1403, N1404, N1405, N1406, N1407, N1838,
         N1888, n139, n141, n142, n143, n144, n145, n148, n149, n600, n601,
         n602, n603, n604, n605, n606, n607, n610, n611, n612, n613, n614,
         n615, n616, n617, n624, n625, n627, n628, n629, n630, n631, n632,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, r616_carry_3_, r616_carry_4_, r616_carry_5_,
         r616_carry_6_, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n19, n20,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n140,
         n146, n147, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490;
  wire   [1:0] mode_w;
  wire   [3:2] coeff_num_w;
  wire   [3:2] coeff_num_r;
  wire   [7:0] addr_ram8x8_w;
  wire   [8:0] state;
  wire   [7:2] next_state;
  wire   [8:0] count_w;
  wire   [3:0] count_r1;
  wire   [3:0] full;
  wire   [2:0] rd_cnt;
  wire   [2:0] rd_num;
  wire   [1:0] count_r1_ram4x4;
  wire   [1:0] count_r2_ram4x4;
  wire   [6:4] r620_carry;
  wire   [5:3] r619_carry;

  mem_ctrl_tran_DW01_inc_0 r608 ( .A(addr_ram8x8_w), .SUM({N767, N766, N765, 
        N764, N763, N762, N761, N760}) );
  mem_ctrl_tran_DW01_inc_5 add_620_aco ( .A({n10, n3, n9, n8, n7, n6, n4, n5, 
        n1}), .SUM({N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, 
        N1399}) );
  mem_ctrl_tran_DW01_inc_4 add_612_aco ( .A({n10, n3, n9, n8, n7, n6, n4, n5, 
        n1}), .SUM({N1369, N1368, N1367, N1366, N1365, N1364, N1363, N1362, 
        N1361}) );
  mem_ctrl_tran_DW01_inc_3 add_415_aco ( .A({n10, n3, n9, n8, n7, n6, n4, n5, 
        n1}), .SUM({N732, N731, N730, N729, N728, N727, N726, N725, N724}) );
  mem_ctrl_tran_DW01_inc_2 add_455_aco ( .A({n10, n3, n9, n8, n7, n6, n4, n5, 
        n1}), .SUM({N859, N858, N857, N856, N855, N854, N853, N852, N851}) );
  mem_ctrl_tran_DW01_inc_1 add_484_aco ( .A({n10, n3, n9, n8, n7, n6, n4, n5, 
        n1}), .SUM({N987, N986, N985, N984, N983, N982, N981, N980, N979}) );
  TLATNX1 coeff_num_r_reg_3_ ( .D(mode_r_0_), .GN(n141), .Q(coeff_num_r[3]) );
  TLATX1 mode_r_reg_1_ ( .G(N593), .D(mode_w[1]), .Q(n141), .QN(n610) );
  TLATNX1 coeff_num_w_reg_2_ ( .D(n490), .GN(mode_w[1]), .Q(coeff_num_w[2]), 
        .QN(n20) );
  TLATNX1 coeff_num_w_reg_3_ ( .D(mode_w[0]), .GN(mode_w[1]), .Q(
        coeff_num_w[3]) );
  TLATX1 mode_r_reg_0_ ( .G(N593), .D(mode_w[0]), .Q(mode_r_0_), .QN(n611) );
  TLATNX1 coeff_shift_r_reg_0_ ( .D(mode_r_0_), .GN(n141), .Q(coeff_shift_r_0_) );
  TLATNX1 coeff_num_r_reg_2_ ( .D(n611), .GN(n141), .Q(coeff_num_r[2]), .QN(
        n11) );
  TLATNX1 coeff_shift_w_reg_0_ ( .D(mode_w[0]), .GN(mode_w[1]), .Q(
        coeff_shift_w_0_) );
  DFFRHQX1 count_r2_ram4x4_reg_1_ ( .D(n700), .CK(clk), .RN(rstn), .Q(
        count_r2_ram4x4[1]) );
  DFFRHQX1 count_r1_ram4x4_reg_1_ ( .D(n677), .CK(clk), .RN(rstn), .Q(
        count_r1_ram4x4[1]) );
  DFFRHQX1 count_r1_ram4x4_reg_0_ ( .D(n676), .CK(clk), .RN(rstn), .Q(
        count_r1_ram4x4[0]) );
  DFFRHQX1 count_r2_ram4x4_reg_0_ ( .D(n678), .CK(clk), .RN(rstn), .Q(
        count_r2_ram4x4[0]) );
  DFFRHQX1 en_ram8x8_r_reg ( .D(n664), .CK(clk), .RN(rstn), .Q(en_ram8x8_r) );
  DFFRHQX1 wr_rd_ram8x8_w_reg ( .D(n679), .CK(clk), .RN(rstn), .Q(
        wr_rd_ram8x8_w) );
  DFFRHQX1 en_ram8x8_w_reg ( .D(N1838), .CK(clk), .RN(rstn), .Q(en_ram8x8_w)
         );
  DFFRHQX1 rd_num_reg_2_ ( .D(n701), .CK(clk), .RN(rstn), .Q(rd_num[2]) );
  DFFRHQX1 wr_rd_ram4x4_2_reg ( .D(n686), .CK(clk), .RN(rstn), .Q(
        wr_rd_ram4x4_2) );
  DFFRHQX1 wr_rd_ram4x4_1_reg ( .D(n683), .CK(clk), .RN(rstn), .Q(
        wr_rd_ram4x4_1) );
  DFFRHQX1 wr_rd_ram4x4_3_reg ( .D(n687), .CK(clk), .RN(rstn), .Q(
        wr_rd_ram4x4_3) );
  DFFRHQX1 wr_rd_ram4x4_4_reg ( .D(n685), .CK(clk), .RN(rstn), .Q(
        wr_rd_ram4x4_4) );
  DFFRHQX1 rd_num_reg_1_ ( .D(n690), .CK(clk), .RN(rstn), .Q(rd_num[1]) );
  DFFRHQX1 rd_num_reg_0_ ( .D(n691), .CK(clk), .RN(rstn), .Q(rd_num[0]) );
  DFFRHQX1 en_ram4x4_2_reg ( .D(n661), .CK(clk), .RN(rstn), .Q(en_ram4x4_2) );
  DFFRHQX1 en_ram4x4_3_reg ( .D(n660), .CK(clk), .RN(rstn), .Q(en_ram4x4_3) );
  DFFRHQX1 en_ram4x4_1_reg ( .D(n662), .CK(clk), .RN(rstn), .Q(en_ram4x4_1) );
  DFFRHQX1 en_ram4x4_4_reg ( .D(n659), .CK(clk), .RN(rstn), .Q(en_ram4x4_4) );
  DFFRHQX1 ram4x4_4_ready_reg ( .D(n655), .CK(clk), .RN(rstn), .Q(
        ram4x4_4_ready) );
  DFFRHQX1 ram4x4_2_ready_reg ( .D(n657), .CK(clk), .RN(rstn), .Q(
        ram4x4_2_ready) );
  DFFRHQX1 ram4x4_3_ready_reg ( .D(n656), .CK(clk), .RN(rstn), .Q(
        ram4x4_3_ready) );
  DFFRHQX1 ram4x4_1_ready_reg ( .D(n658), .CK(clk), .RN(rstn), .Q(
        ram4x4_1_ready) );
  DFFRHQX1 mode_out_reg_1_ ( .D(n654), .CK(clk), .RN(rstn), .Q(mode_out[1]) );
  DFFRHQX1 mode_out_reg_0_ ( .D(n653), .CK(clk), .RN(rstn), .Q(mode_out[0]) );
  DFFRHQX1 ram8x8_r_ready_reg ( .D(n663), .CK(clk), .RN(rstn), .Q(
        ram8x8_r_ready) );
  DFFRHQX1 ram8x8_w_ready_reg ( .D(N1888), .CK(clk), .RN(rstn), .Q(
        ram8x8_w_ready) );
  DFFRHQX1 rd_cnt_reg_2_ ( .D(n712), .CK(clk), .RN(rstn), .Q(rd_cnt[2]) );
  DFFRHQX1 ram8_4_reg ( .D(n709), .CK(clk), .RN(rstn), .Q(ram8_4) );
  DFFRHQX1 ram_write_reg_reg ( .D(ram_write), .CK(clk), .RN(rstn), .Q(
        ram_write_reg) );
  DFFRHQX1 state_reg_8_ ( .D(n605), .CK(clk), .RN(rstn), .Q(state[8]) );
  DFFRHQX1 state_reg_6_ ( .D(next_state[6]), .CK(clk), .RN(rstn), .Q(state[6])
         );
  DFFRHQX1 state_reg_1_ ( .D(n607), .CK(clk), .RN(rstn), .Q(state[1]) );
  DFFRHQX1 state_reg_3_ ( .D(next_state[3]), .CK(clk), .RN(rstn), .Q(state[3])
         );
  DFFRHQX1 state_reg_7_ ( .D(n26), .CK(clk), .RN(rstn), .Q(state[7]) );
  DFFRHQX1 rd_cnt_reg_0_ ( .D(n711), .CK(clk), .RN(rstn), .Q(rd_cnt[0]) );
  DFFRHQX1 state_reg_5_ ( .D(n606), .CK(clk), .RN(rstn), .Q(state[5]) );
  DFFRHQX1 rd_cnt_reg_1_ ( .D(n710), .CK(clk), .RN(rstn), .Q(rd_cnt[1]) );
  DFFRHQX1 full_reg_3_ ( .D(n698), .CK(clk), .RN(rstn), .Q(full[3]) );
  DFFRHQX1 state_reg_4_ ( .D(next_state[4]), .CK(clk), .RN(rstn), .Q(state[4])
         );
  DFFRHQX1 state_reg_2_ ( .D(next_state[2]), .CK(clk), .RN(rstn), .Q(state[2])
         );
  DFFRHQX1 full_reg_2_ ( .D(n689), .CK(clk), .RN(rstn), .Q(full[2]) );
  DFFRHQX1 full_reg_1_ ( .D(n688), .CK(clk), .RN(rstn), .Q(full[1]) );
  DFFRHQX1 full_reg_0_ ( .D(n684), .CK(clk), .RN(rstn), .Q(full[0]) );
  DFFRHQX1 ram_reg ( .D(ram_write), .CK(clk), .RN(rstn), .Q(ram) );
  DFFRHQX1 mode_w_reg_1_ ( .D(n601), .CK(clk), .RN(rstn), .Q(mode_w[1]) );
  DFFRHQX1 count_r1_reg_3_ ( .D(n603), .CK(clk), .RN(rstn), .Q(count_r1[3]) );
  DFFRHQX1 count_r2_reg_2_ ( .D(n695), .CK(clk), .RN(rstn), .Q(N1074) );
  DFFRHQX1 mode_w_reg_0_ ( .D(n600), .CK(clk), .RN(rstn), .Q(mode_w[0]) );
  DFFRHQX1 count_r1_reg_2_ ( .D(n693), .CK(clk), .RN(rstn), .Q(count_r1[2]) );
  DFFRHQX1 count_r2_reg_1_ ( .D(n696), .CK(clk), .RN(rstn), .Q(N831) );
  DFFRHQX1 count_r2_reg_0_ ( .D(n697), .CK(clk), .RN(rstn), .Q(N830) );
  DFFRHQX1 count_r1_reg_1_ ( .D(n694), .CK(clk), .RN(rstn), .Q(count_r1[1]) );
  DFFRHQX1 count_r2_reg_3_ ( .D(n714), .CK(clk), .RN(rstn), .Q(count_r2_3_) );
  DFFRHQX1 count_w_reg_8_ ( .D(n645), .CK(clk), .RN(rstn), .Q(count_w[8]) );
  DFFRHQX1 count_w_reg_7_ ( .D(n646), .CK(clk), .RN(rstn), .Q(count_w[7]) );
  DFFRHQX1 count_w_reg_3_ ( .D(n650), .CK(clk), .RN(rstn), .Q(count_w[3]) );
  DFFRHQX1 count_w_reg_0_ ( .D(n715), .CK(clk), .RN(rstn), .Q(count_w[0]) );
  DFFRHQX1 count_w_reg_2_ ( .D(n651), .CK(clk), .RN(rstn), .Q(count_w[2]) );
  DFFRHQX1 count_w_reg_1_ ( .D(n652), .CK(clk), .RN(rstn), .Q(count_w[1]) );
  DFFRHQX1 count_w_reg_6_ ( .D(n647), .CK(clk), .RN(rstn), .Q(count_w[6]) );
  DFFRHQX1 count_w_reg_5_ ( .D(n648), .CK(clk), .RN(rstn), .Q(count_w[5]) );
  DFFRHQX1 count_w_reg_4_ ( .D(n649), .CK(clk), .RN(rstn), .Q(count_w[4]) );
  DFFSXL addr_ram4x4_4_reg_0_ ( .D(n602), .CK(clk), .SN(rstn), .Q(
        addr_ram4x4_4[0]), .QN(n142) );
  DFFSXL addr_ram4x4_4_reg_1_ ( .D(n675), .CK(clk), .SN(rstn), .Q(
        addr_ram4x4_4[1]), .QN(n613) );
  DFFSXL addr_ram4x4_1_reg_1_ ( .D(n681), .CK(clk), .SN(rstn), .Q(
        addr_ram4x4_1[1]), .QN(n624) );
  DFFSXL addr_ram4x4_3_reg_0_ ( .D(n672), .CK(clk), .SN(rstn), .Q(
        addr_ram4x4_3[0]), .QN(n617) );
  DFFSXL addr_ram4x4_2_reg_1_ ( .D(n667), .CK(clk), .SN(rstn), .Q(
        addr_ram4x4_2[1]), .QN(n144) );
  DFFSXL addr_ram4x4_1_reg_2_ ( .D(n680), .CK(clk), .SN(rstn), .Q(
        addr_ram4x4_1[2]), .QN(n143) );
  DFFSXL addr_ram4x4_4_reg_2_ ( .D(n674), .CK(clk), .SN(rstn), .Q(
        addr_ram4x4_4[2]), .QN(n612) );
  DFFSXL addr_ram4x4_1_reg_3_ ( .D(n699), .CK(clk), .SN(rstn), .Q(
        addr_ram4x4_1[3]), .QN(n139) );
  DFFSXL addr_ram4x4_2_reg_2_ ( .D(n666), .CK(clk), .SN(rstn), .Q(
        addr_ram4x4_2[2]), .QN(n627) );
  DFFSXL addr_ram4x4_4_reg_3_ ( .D(n673), .CK(clk), .SN(rstn), .Q(
        addr_ram4x4_4[3]), .QN(n145) );
  DFFSXL addr_ram4x4_2_reg_3_ ( .D(n665), .CK(clk), .SN(rstn), .Q(
        addr_ram4x4_2[3]) );
  DFFSXL addr_ram4x4_3_reg_1_ ( .D(n671), .CK(clk), .SN(rstn), .Q(
        addr_ram4x4_3[1]), .QN(n616) );
  DFFSXL addr_ram4x4_3_reg_2_ ( .D(n670), .CK(clk), .SN(rstn), .Q(
        addr_ram4x4_3[2]), .QN(n615) );
  DFFSXL addr_ram4x4_3_reg_3_ ( .D(n669), .CK(clk), .SN(rstn), .Q(
        addr_ram4x4_3[3]), .QN(n614) );
  DFFSXL addr_ram8x8_w_reg_7_ ( .D(n637), .CK(clk), .SN(rstn), .Q(
        addr_ram8x8_w[7]), .QN(n149) );
  DFFSXL addr_ram8x8_w_reg_6_ ( .D(n638), .CK(clk), .SN(rstn), .Q(
        addr_ram8x8_w[6]), .QN(n148) );
  DFFSXL addr_ram8x8_w_reg_5_ ( .D(n639), .CK(clk), .SN(rstn), .Q(
        addr_ram8x8_w[5]), .QN(n629) );
  DFFSXL addr_ram8x8_w_reg_4_ ( .D(n640), .CK(clk), .SN(rstn), .Q(
        addr_ram8x8_w[4]), .QN(n630) );
  DFFSXL addr_ram8x8_w_reg_3_ ( .D(n641), .CK(clk), .SN(rstn), .Q(
        addr_ram8x8_w[3]), .QN(n631) );
  DFFSXL addr_ram8x8_w_reg_2_ ( .D(n642), .CK(clk), .SN(rstn), .Q(
        addr_ram8x8_w[2]), .QN(n632) );
  DFFSXL addr_ram8x8_w_reg_1_ ( .D(n643), .CK(clk), .SN(rstn), .Q(
        addr_ram8x8_w[1]), .QN(n36) );
  DFFSXL addr_ram8x8_w_reg_0_ ( .D(n644), .CK(clk), .SN(rstn), .Q(
        addr_ram8x8_w[0]), .QN(n37) );
  JKFFRXL count_r1_reg_0_ ( .J(n604), .K(n636), .CK(clk), .RN(rstn), .Q(
        count_r1[0]), .QN(n635) );
  DFFSXL state_reg_0_ ( .D(n25), .CK(clk), .SN(rstn), .Q(state[0]) );
  DFFSXL finish_reg ( .D(n692), .CK(clk), .SN(rstn), .Q(n489), .QN(n196) );
  DFFSXL addr_ram8x8_r_reg_7_ ( .D(n713), .CK(clk), .SN(rstn), .QN(n63) );
  DFFSXL addr_ram8x8_r_reg_6_ ( .D(n702), .CK(clk), .SN(rstn), .QN(n117) );
  DFFSXL addr_ram8x8_r_reg_5_ ( .D(n703), .CK(clk), .SN(rstn), .QN(n114) );
  DFFSXL addr_ram8x8_r_reg_4_ ( .D(n704), .CK(clk), .SN(rstn), .QN(n111) );
  DFFSXL addr_ram8x8_r_reg_3_ ( .D(n705), .CK(clk), .SN(rstn), .Q(n486), .QN(
        n108) );
  DFFSXL addr_ram8x8_r_reg_2_ ( .D(n706), .CK(clk), .SN(rstn), .Q(n487), .QN(
        n105) );
  DFFSXL addr_ram8x8_r_reg_1_ ( .D(n707), .CK(clk), .SN(rstn), .Q(n488), .QN(
        n102) );
  DFFSXL addr_ram8x8_r_reg_0_ ( .D(n708), .CK(clk), .SN(rstn), .QN(n98) );
  DFFSX1 addr_ram4x4_1_reg_0_ ( .D(n682), .CK(clk), .SN(rstn), .Q(
        addr_ram4x4_1[0]), .QN(n625) );
  DFFSX1 addr_ram4x4_2_reg_0_ ( .D(n668), .CK(clk), .SN(rstn), .Q(
        addr_ram4x4_2[0]), .QN(n628) );
  AND2X2 U3 ( .A(count_w[0]), .B(n2), .Y(n1) );
  NAND4X1 U4 ( .A(n442), .B(n443), .C(n444), .D(n445), .Y(n2) );
  AND2X2 U5 ( .A(count_w[7]), .B(n2), .Y(n3) );
  AND2X2 U6 ( .A(count_w[2]), .B(n2), .Y(n4) );
  AND2X2 U7 ( .A(count_w[1]), .B(n2), .Y(n5) );
  AND2X2 U8 ( .A(count_w[3]), .B(n2), .Y(n6) );
  AND2X2 U9 ( .A(count_w[4]), .B(n2), .Y(n7) );
  AND2X2 U10 ( .A(count_w[5]), .B(n2), .Y(n8) );
  AND2X2 U11 ( .A(count_w[6]), .B(n2), .Y(n9) );
  AND2X2 U12 ( .A(n2), .B(count_w[8]), .Y(n10) );
  INVX1 U13 ( .A(n25), .Y(n64) );
  NAND2X1 U14 ( .A(n332), .B(n64), .Y(n62) );
  INVX1 U15 ( .A(n181), .Y(n66) );
  OR2X2 U16 ( .A(next_state[3]), .B(next_state[6]), .Y(n53) );
  NOR2X1 U17 ( .A(n417), .B(n87), .Y(n67) );
  OR2X2 U18 ( .A(n606), .B(n607), .Y(n54) );
  AND3X2 U19 ( .A(n64), .B(n197), .C(n368), .Y(n51) );
  INVX1 U20 ( .A(n26), .Y(n197) );
  NOR2X1 U21 ( .A(n409), .B(n87), .Y(n50) );
  INVX1 U22 ( .A(n28), .Y(N752) );
  NOR3X1 U23 ( .A(N807), .B(n43), .C(n42), .Y(N808) );
  NAND4X1 U24 ( .A(n368), .B(n386), .C(n199), .D(n64), .Y(n258) );
  INVX1 U25 ( .A(n214), .Y(n165) );
  INVX1 U26 ( .A(n605), .Y(n87) );
  OAI221XL U27 ( .A0(n429), .A1(n430), .B0(n423), .B1(n431), .C0(n432), .Y(n25) );
  BUFX3 U28 ( .A(next_state[7]), .Y(n26) );
  OAI22X1 U29 ( .A0(n405), .A1(n436), .B0(n465), .B1(n462), .Y(next_state[7])
         );
  NAND2X1 U30 ( .A(n28), .B(n29), .Y(n35) );
  NOR2X1 U31 ( .A(n37), .B(n36), .Y(n29) );
  INVX1 U32 ( .A(N737), .Y(N749) );
  OAI21XL U33 ( .A0(n436), .A1(n407), .B0(n464), .Y(n605) );
  NOR3X1 U34 ( .A(n489), .B(start), .C(n87), .Y(n52) );
  INVX1 U35 ( .A(ram), .Y(n44) );
  AND3X2 U36 ( .A(n19), .B(addr_ram8x8_w[2]), .C(addr_ram8x8_w[3]), .Y(n30) );
  XNOR2X1 U37 ( .A(N749), .B(addr_ram8x8_w[4]), .Y(n19) );
  NOR3X1 U38 ( .A(N782), .B(n40), .C(n39), .Y(N783) );
  NOR2X1 U39 ( .A(n635), .B(coeff_shift_r_0_), .Y(N824) );
  MX2X1 U40 ( .A(count_r1[2]), .B(count_r1[1]), .S0(coeff_shift_r_0_), .Y(N826) );
  ADDFX2 U41 ( .A(count_r1[1]), .B(count_r2_3_), .CI(r619_carry[3]), .CO(
        r619_carry[4]), .S(N1068) );
  ADDFX2 U42 ( .A(N825), .B(count_r2_3_), .CI(r616_carry_3_), .CO(
        r616_carry_4_), .S(N833) );
  MX2X1 U43 ( .A(count_r1[1]), .B(count_r1[0]), .S0(coeff_shift_r_0_), .Y(N825) );
  MX2X1 U44 ( .A(count_r1[3]), .B(count_r1[2]), .S0(coeff_shift_r_0_), .Y(N827) );
  NOR2X1 U45 ( .A(n20), .B(coeff_shift_w_0_), .Y(N737) );
  NOR2BX1 U46 ( .AN(N805), .B(coeff_num_r[2]), .Y(N807) );
  NOR2X1 U47 ( .A(n20), .B(coeff_shift_w_0_), .Y(N716) );
  NOR2X1 U48 ( .A(n20), .B(coeff_shift_w_0_), .Y(N329) );
  MX2X1 U49 ( .A(coeff_num_w[3]), .B(coeff_num_w[2]), .S0(coeff_shift_w_0_), 
        .Y(N717) );
  MX2X1 U50 ( .A(coeff_num_w[3]), .B(coeff_num_w[2]), .S0(coeff_shift_w_0_), 
        .Y(N330) );
  MX2X1 U51 ( .A(coeff_num_w[3]), .B(coeff_num_w[2]), .S0(coeff_shift_w_0_), 
        .Y(N738) );
  AND2X1 U52 ( .A(r620_carry[6]), .B(count_r1[3]), .Y(N1079) );
  XOR2X1 U53 ( .A(count_r1[3]), .B(r620_carry[6]), .Y(N1078) );
  AND2X1 U54 ( .A(r616_carry_6_), .B(N828), .Y(N837) );
  XOR2X1 U55 ( .A(N828), .B(r616_carry_6_), .Y(N836) );
  AND2X1 U56 ( .A(r620_carry[5]), .B(count_r1[2]), .Y(r620_carry[6]) );
  XOR2X1 U57 ( .A(count_r1[2]), .B(r620_carry[5]), .Y(N1077) );
  AND2X1 U58 ( .A(r616_carry_5_), .B(N827), .Y(r616_carry_6_) );
  XOR2X1 U59 ( .A(N827), .B(r616_carry_5_), .Y(N835) );
  AND2X1 U60 ( .A(r619_carry[5]), .B(count_r1[3]), .Y(N1071) );
  XOR2X1 U61 ( .A(count_r1[3]), .B(r619_carry[5]), .Y(N1070) );
  AND2X1 U62 ( .A(r620_carry[4]), .B(count_r1[1]), .Y(r620_carry[5]) );
  XOR2X1 U63 ( .A(count_r1[1]), .B(r620_carry[4]), .Y(N1076) );
  AND2X1 U64 ( .A(r616_carry_4_), .B(N826), .Y(r616_carry_5_) );
  XOR2X1 U65 ( .A(N826), .B(r616_carry_4_), .Y(N834) );
  AND2X1 U66 ( .A(r619_carry[4]), .B(count_r1[2]), .Y(r619_carry[5]) );
  XOR2X1 U67 ( .A(count_r1[2]), .B(r619_carry[4]), .Y(N1069) );
  AND2X1 U68 ( .A(count_r1[0]), .B(count_r2_3_), .Y(r620_carry[4]) );
  XOR2X1 U69 ( .A(count_r2_3_), .B(count_r1[0]), .Y(N1075) );
  AND2X1 U70 ( .A(N824), .B(N1074), .Y(r616_carry_3_) );
  XOR2X1 U71 ( .A(N1074), .B(N824), .Y(N832) );
  AND2X1 U72 ( .A(count_r1[0]), .B(N1074), .Y(r619_carry[3]) );
  XOR2X1 U73 ( .A(N1074), .B(count_r1[0]), .Y(N1067) );
  AND2X1 U74 ( .A(coeff_num_w[3]), .B(coeff_shift_w_0_), .Y(N331) );
  AND2X1 U75 ( .A(coeff_num_w[3]), .B(coeff_shift_w_0_), .Y(N718) );
  AND2X1 U76 ( .A(coeff_num_w[3]), .B(coeff_shift_w_0_), .Y(N739) );
  OR2X1 U77 ( .A(N737), .B(N738), .Y(n27) );
  OR2X1 U78 ( .A(n27), .B(N739), .Y(n28) );
  OAI2BB1X1 U79 ( .A0N(N737), .A1N(N738), .B0(n27), .Y(N750) );
  OAI2BB1X1 U80 ( .A0N(n27), .A1N(N739), .B0(n28), .Y(N751) );
  XNOR2X1 U81 ( .A(coeff_num_r[2]), .B(coeff_num_r[3]), .Y(N780) );
  AND2X1 U82 ( .A(N780), .B(n11), .Y(N782) );
  XNOR2X1 U83 ( .A(coeff_num_r[2]), .B(coeff_num_r[3]), .Y(N805) );
  AND2X1 U84 ( .A(count_r1[3]), .B(coeff_shift_r_0_), .Y(N828) );
  XNOR2X1 U85 ( .A(N751), .B(addr_ram8x8_w[6]), .Y(n33) );
  XNOR2X1 U86 ( .A(N750), .B(addr_ram8x8_w[5]), .Y(n32) );
  XNOR2X1 U87 ( .A(N752), .B(addr_ram8x8_w[7]), .Y(n31) );
  NAND4X1 U88 ( .A(n33), .B(n32), .C(n31), .D(n30), .Y(n34) );
  NOR2X1 U89 ( .A(n35), .B(n34), .Y(N758) );
  XNOR2X1 U90 ( .A(N780), .B(count_r1[3]), .Y(n38) );
  NAND3X1 U91 ( .A(count_r1[1]), .B(n38), .C(count_r1[0]), .Y(n40) );
  XOR2X1 U92 ( .A(n11), .B(count_r1[2]), .Y(n39) );
  XNOR2X1 U93 ( .A(N805), .B(count_r2_3_), .Y(n41) );
  NAND3X1 U94 ( .A(N831), .B(n41), .C(N830), .Y(n43) );
  XOR2X1 U95 ( .A(n11), .B(N1074), .Y(n42) );
  NOR2X1 U96 ( .A(n44), .B(n45), .Y(wr_rd_ram8x8_2) );
  NOR2X1 U97 ( .A(ram), .B(n45), .Y(wr_rd_ram8x8_1) );
  MXI2X1 U98 ( .A(n46), .B(n47), .S0(n44), .Y(ram8x8_2_ready) );
  MXI2X1 U99 ( .A(n47), .B(n46), .S0(n44), .Y(ram8x8_1_ready) );
  INVX1 U100 ( .A(ram8x8_w_ready), .Y(n46) );
  NAND2X1 U101 ( .A(n48), .B(n49), .Y(n715) );
  AOI222X1 U102 ( .A0(N1361), .A1(n50), .B0(count_w[0]), .B1(n51), .C0(N1399), 
        .C1(n52), .Y(n49) );
  AOI222X1 U103 ( .A0(N979), .A1(n26), .B0(N851), .B1(n53), .C0(N724), .C1(n54), .Y(n48) );
  OAI22X1 U104 ( .A0(n55), .A1(n56), .B0(n57), .B1(n58), .Y(n714) );
  AOI21X1 U105 ( .A0(n59), .A1(n60), .B0(n61), .Y(n57) );
  OAI211X1 U106 ( .A0(n62), .A1(n63), .B0(n64), .C0(n65), .Y(n713) );
  AOI22X1 U107 ( .A0(N837), .A1(n66), .B0(N1079), .B1(n67), .Y(n65) );
  OAI22X1 U108 ( .A0(n68), .A1(n69), .B0(n70), .B1(n71), .Y(n712) );
  XNOR2X1 U109 ( .A(n72), .B(n69), .Y(n70) );
  NAND2X1 U110 ( .A(rd_cnt[1]), .B(rd_cnt[0]), .Y(n72) );
  MXI2X1 U111 ( .A(n68), .B(n71), .S0(n73), .Y(n711) );
  OAI22X1 U112 ( .A0(n68), .A1(n74), .B0(n75), .B1(n71), .Y(n710) );
  NAND2X1 U113 ( .A(n76), .B(n77), .Y(n71) );
  OAI211X1 U114 ( .A0(n78), .A1(n79), .B0(n80), .C0(n81), .Y(n77) );
  AOI22X1 U115 ( .A0(n82), .A1(n83), .B0(n84), .B1(n85), .Y(n81) );
  INVX1 U116 ( .A(n86), .Y(n82) );
  XNOR2X1 U117 ( .A(rd_cnt[0]), .B(rd_cnt[1]), .Y(n75) );
  AOI2BB1X1 U118 ( .A0N(n87), .A1N(n88), .B0(n89), .Y(n68) );
  MXI2X1 U119 ( .A(n90), .B(n91), .S0(n92), .Y(n709) );
  NOR2X1 U120 ( .A(n93), .B(n94), .Y(n92) );
  AOI21X1 U121 ( .A0(n95), .A1(n605), .B0(n26), .Y(n90) );
  NAND4X1 U122 ( .A(n88), .B(rd_cnt[1]), .C(rd_cnt[0]), .D(n69), .Y(n95) );
  INVX1 U123 ( .A(rd_cnt[2]), .Y(n69) );
  AOI21X1 U124 ( .A0(n78), .A1(n96), .B0(n97), .Y(n88) );
  OAI211X1 U125 ( .A0(n62), .A1(n98), .B0(n99), .C0(n100), .Y(n708) );
  AOI22X1 U126 ( .A0(N830), .A1(n66), .B0(n67), .B1(N830), .Y(n100) );
  AOI21X1 U127 ( .A0(N830), .A1(n101), .B0(n25), .Y(n99) );
  OAI211X1 U128 ( .A0(n62), .A1(n102), .B0(n103), .C0(n104), .Y(n707) );
  AOI22X1 U129 ( .A0(N831), .A1(n66), .B0(n67), .B1(N831), .Y(n104) );
  AOI21X1 U130 ( .A0(N831), .A1(n101), .B0(n25), .Y(n103) );
  OAI211X1 U131 ( .A0(n62), .A1(n105), .B0(n106), .C0(n107), .Y(n706) );
  AOI22X1 U132 ( .A0(N832), .A1(n66), .B0(n67), .B1(N1074), .Y(n107) );
  AOI21X1 U133 ( .A0(N1067), .A1(n101), .B0(n25), .Y(n106) );
  OAI211X1 U134 ( .A0(n62), .A1(n108), .B0(n109), .C0(n110), .Y(n705) );
  AOI22X1 U135 ( .A0(N833), .A1(n66), .B0(N1075), .B1(n67), .Y(n110) );
  AOI21X1 U136 ( .A0(N1068), .A1(n101), .B0(n25), .Y(n109) );
  OAI211X1 U137 ( .A0(n62), .A1(n111), .B0(n112), .C0(n113), .Y(n704) );
  AOI22X1 U138 ( .A0(N834), .A1(n66), .B0(N1076), .B1(n67), .Y(n113) );
  AOI21X1 U139 ( .A0(N1069), .A1(n101), .B0(n25), .Y(n112) );
  OAI211X1 U140 ( .A0(n62), .A1(n114), .B0(n115), .C0(n116), .Y(n703) );
  AOI22X1 U141 ( .A0(N835), .A1(n66), .B0(N1077), .B1(n67), .Y(n116) );
  AOI21X1 U142 ( .A0(N1070), .A1(n101), .B0(n25), .Y(n115) );
  OAI211X1 U143 ( .A0(n62), .A1(n117), .B0(n118), .C0(n119), .Y(n702) );
  AOI22X1 U144 ( .A0(N836), .A1(n66), .B0(N1078), .B1(n67), .Y(n119) );
  AOI21X1 U145 ( .A0(N1071), .A1(n101), .B0(n25), .Y(n118) );
  NOR2BX1 U146 ( .AN(n62), .B(n120), .Y(n101) );
  OAI21XL U147 ( .A0(n121), .A1(n122), .B0(n123), .Y(n701) );
  AOI31X1 U148 ( .A0(n96), .A1(n124), .A2(n76), .B0(n125), .Y(n123) );
  AND4X1 U149 ( .A(n126), .B(n127), .C(n128), .D(n129), .Y(n121) );
  AOI221X1 U150 ( .A0(n97), .A1(n605), .B0(n130), .B1(n131), .C0(n89), .Y(n126) );
  OAI211X1 U151 ( .A0(n132), .A1(n133), .B0(n134), .C0(n135), .Y(n97) );
  AOI22X1 U152 ( .A0(n136), .A1(n137), .B0(n83), .B1(n86), .Y(n135) );
  NAND4X1 U153 ( .A(n486), .B(n488), .C(n138), .D(n140), .Y(n86) );
  AND4X1 U154 ( .A(n117), .B(n63), .C(n114), .D(n111), .Y(n140) );
  NOR2X1 U155 ( .A(n487), .B(n98), .Y(n138) );
  MXI2X1 U156 ( .A(n146), .B(n147), .S0(n150), .Y(n700) );
  NAND3X1 U157 ( .A(n151), .B(n152), .C(count_r2_ram4x4[0]), .Y(n147) );
  NOR2X1 U158 ( .A(n153), .B(n154), .Y(n146) );
  AOI21X1 U159 ( .A0(count_r2_ram4x4[0]), .A1(n151), .B0(n155), .Y(n153) );
  OAI211X1 U160 ( .A0(n156), .A1(n157), .B0(n158), .C0(n159), .Y(n699) );
  AOI31X1 U161 ( .A0(n160), .A1(addr_ram4x4_1[2]), .A2(n161), .B0(n25), .Y(
        n159) );
  OAI21XL U162 ( .A0(n161), .A1(n162), .B0(addr_ram4x4_1[3]), .Y(n158) );
  OAI32X1 U163 ( .A0(n164), .A1(n165), .A2(addr_ram4x4_1[0]), .B0(n166), .B1(
        n167), .Y(n698) );
  AOI21X1 U164 ( .A0(n168), .A1(n137), .B0(n169), .Y(n166) );
  NAND3BX1 U165 ( .AN(n624), .B(addr_ram4x4_1[2]), .C(addr_ram4x4_1[3]), .Y(
        n164) );
  MXI2X1 U166 ( .A(n56), .B(n170), .S0(N830), .Y(n697) );
  MXI2X1 U167 ( .A(n171), .B(n172), .S0(N831), .Y(n696) );
  NAND2X1 U168 ( .A(n173), .B(N830), .Y(n171) );
  MXI2X1 U169 ( .A(n174), .B(n175), .S0(n60), .Y(n695) );
  NAND3X1 U170 ( .A(N831), .B(N830), .C(n173), .Y(n175) );
  INVX1 U171 ( .A(n56), .Y(n173) );
  NAND2X1 U172 ( .A(n59), .B(n636), .Y(n56) );
  INVX1 U173 ( .A(n61), .Y(n174) );
  OAI21XL U174 ( .A0(N831), .A1(n176), .B0(n172), .Y(n61) );
  INVX1 U175 ( .A(n177), .Y(n172) );
  OAI21XL U176 ( .A0(N830), .A1(n176), .B0(n170), .Y(n177) );
  NOR2X1 U177 ( .A(n178), .B(n179), .Y(n170) );
  INVX1 U178 ( .A(n59), .Y(n176) );
  OAI31X1 U179 ( .A0(n180), .A1(N808), .A2(n181), .B0(n182), .Y(n59) );
  AOI31X1 U180 ( .A0(n183), .A1(n55), .A2(n184), .B0(n185), .Y(n182) );
  AOI211X1 U181 ( .A0(n186), .A1(n60), .B0(n187), .C0(n188), .Y(n185) );
  INVX1 U182 ( .A(n189), .Y(n187) );
  INVX1 U183 ( .A(N1074), .Y(n60) );
  NAND2X1 U184 ( .A(N1074), .B(n186), .Y(n55) );
  AND3X1 U185 ( .A(N830), .B(n58), .C(N831), .Y(n186) );
  INVX1 U186 ( .A(n190), .Y(n183) );
  INVX1 U187 ( .A(N783), .Y(n180) );
  MXI2X1 U188 ( .A(n191), .B(n192), .S0(count_r1[1]), .Y(n694) );
  NAND2X1 U189 ( .A(n604), .B(count_r1[0]), .Y(n191) );
  OAI2BB2X1 U190 ( .B0(n193), .B1(n194), .A0N(n195), .A1N(count_r1[2]), .Y(
        n693) );
  OAI211X1 U191 ( .A0(n50), .A1(n196), .B0(n64), .C0(n197), .Y(n692) );
  NAND3X1 U192 ( .A(n198), .B(n199), .C(n200), .Y(n691) );
  AOI22X1 U193 ( .A0(rd_num[0]), .A1(n201), .B0(n76), .B1(n202), .Y(n200) );
  INVX1 U194 ( .A(n80), .Y(n202) );
  AOI22X1 U195 ( .A0(n132), .A1(n203), .B0(n204), .B1(n136), .Y(n80) );
  INVX1 U196 ( .A(n137), .Y(n204) );
  NAND2X1 U197 ( .A(n143), .B(n205), .Y(n137) );
  OAI211X1 U198 ( .A0(n87), .A1(n134), .B0(n128), .C0(n206), .Y(n201) );
  INVX1 U199 ( .A(n207), .Y(n206) );
  NAND2X1 U200 ( .A(n84), .B(n208), .Y(n134) );
  OAI221XL U201 ( .A0(n209), .A1(n210), .B0(n211), .B1(n165), .C0(n212), .Y(
        n690) );
  AOI31X1 U202 ( .A0(n84), .A1(n85), .A2(n76), .B0(n213), .Y(n212) );
  NOR2X1 U203 ( .A(n87), .B(n89), .Y(n76) );
  INVX1 U204 ( .A(n208), .Y(n85) );
  NOR2X1 U205 ( .A(n214), .B(n207), .Y(n209) );
  OAI211X1 U206 ( .A0(n215), .A1(n216), .B0(n217), .C0(n218), .Y(n207) );
  AOI211X1 U207 ( .A0(n219), .A1(n605), .B0(n89), .C0(n220), .Y(n218) );
  NOR2X1 U208 ( .A(n94), .B(n26), .Y(n89) );
  NAND2X1 U209 ( .A(n221), .B(n64), .Y(n94) );
  OAI21XL U210 ( .A0(n83), .A1(n222), .B0(n223), .Y(n221) );
  INVX1 U211 ( .A(n224), .Y(n222) );
  OAI21XL U212 ( .A0(n124), .A1(n79), .B0(n133), .Y(n219) );
  INVX1 U213 ( .A(n203), .Y(n133) );
  OAI32X1 U214 ( .A0(n225), .A1(n217), .A2(addr_ram4x4_2[0]), .B0(n226), .B1(
        n211), .Y(n689) );
  AOI21X1 U215 ( .A0(n227), .A1(n208), .B0(n228), .Y(n226) );
  NAND2X1 U216 ( .A(n627), .B(n229), .Y(n208) );
  NAND2X1 U217 ( .A(n165), .B(n87), .Y(n227) );
  NAND3BX1 U218 ( .AN(n144), .B(addr_ram4x4_2[3]), .C(addr_ram4x4_2[2]), .Y(
        n225) );
  OAI21XL U219 ( .A0(n132), .A1(n198), .B0(n231), .Y(n688) );
  AOI32X1 U220 ( .A0(n617), .A1(n232), .A2(n233), .B0(full[1]), .B1(n234), .Y(
        n231) );
  OAI21XL U221 ( .A0(n87), .A1(n132), .B0(n235), .Y(n234) );
  NOR3X1 U222 ( .A(n614), .B(n616), .C(n615), .Y(n233) );
  NOR2X1 U223 ( .A(addr_ram4x4_3[2]), .B(n236), .Y(n132) );
  OAI21XL U224 ( .A0(n237), .A1(n235), .B0(n129), .Y(n687) );
  INVX1 U225 ( .A(wr_rd_ram4x4_3), .Y(n237) );
  OAI2BB1X1 U226 ( .A0N(wr_rd_ram4x4_2), .A1N(n228), .B0(n217), .Y(n686) );
  OAI21XL U227 ( .A0(n238), .A1(n239), .B0(n216), .Y(n685) );
  INVX1 U228 ( .A(wr_rd_ram4x4_4), .Y(n238) );
  OAI21XL U229 ( .A0(n124), .A1(n240), .B0(n241), .Y(n684) );
  AOI32X1 U230 ( .A0(n142), .A1(n131), .A2(n242), .B0(full[0]), .B1(n243), .Y(
        n241) );
  OAI21XL U231 ( .A0(n124), .A1(n87), .B0(n239), .Y(n243) );
  NOR3X1 U232 ( .A(n145), .B(n613), .C(n612), .Y(n242) );
  INVX1 U233 ( .A(n78), .Y(n124) );
  NAND3X1 U234 ( .A(n244), .B(addr_ram4x4_4[3]), .C(n612), .Y(n78) );
  OAI2BB1X1 U235 ( .A0N(wr_rd_ram4x4_1), .A1N(n169), .B0(n165), .Y(n683) );
  OAI211X1 U236 ( .A0(n245), .A1(n157), .B0(n64), .C0(n246), .Y(n682) );
  MXI2X1 U237 ( .A(n161), .B(n169), .S0(addr_ram4x4_1[0]), .Y(n246) );
  INVX1 U238 ( .A(n247), .Y(n169) );
  OAI211X1 U239 ( .A0(n150), .A1(n157), .B0(n64), .C0(n248), .Y(n681) );
  MXI2X1 U240 ( .A(n249), .B(n250), .S0(n624), .Y(n248) );
  NOR2X1 U241 ( .A(n625), .B(n251), .Y(n250) );
  OAI21XL U242 ( .A0(n251), .A1(addr_ram4x4_1[0]), .B0(n247), .Y(n249) );
  OAI211X1 U243 ( .A0(n252), .A1(n157), .B0(n64), .C0(n253), .Y(n680) );
  MXI2X1 U244 ( .A(n254), .B(n162), .S0(addr_ram4x4_1[2]), .Y(n253) );
  OAI21XL U245 ( .A0(n160), .A1(n251), .B0(n247), .Y(n162) );
  NOR2X1 U246 ( .A(n255), .B(n251), .Y(n254) );
  INVX1 U247 ( .A(n161), .Y(n251) );
  AOI21X1 U248 ( .A0(addr_ram4x4_1[2]), .A1(n205), .B0(n165), .Y(n161) );
  NOR2X1 U249 ( .A(n255), .B(n139), .Y(n205) );
  INVX1 U250 ( .A(n160), .Y(n255) );
  NOR2X1 U251 ( .A(n625), .B(n624), .Y(n160) );
  NAND2X1 U252 ( .A(n247), .B(n168), .Y(n157) );
  NAND3X1 U253 ( .A(n165), .B(n64), .C(n256), .Y(n247) );
  MXI2X1 U254 ( .A(n45), .B(n257), .S0(n258), .Y(n679) );
  NOR2X1 U255 ( .A(n259), .B(n168), .Y(n257) );
  NAND2X1 U256 ( .A(n199), .B(n87), .Y(n168) );
  INVX1 U257 ( .A(wr_rd_ram8x8_w), .Y(n45) );
  MXI2X1 U258 ( .A(n260), .B(n261), .S0(n245), .Y(n678) );
  NAND2X1 U259 ( .A(n151), .B(n152), .Y(n261) );
  AOI211X1 U260 ( .A0(n262), .A1(n605), .B0(n263), .C0(n264), .Y(n260) );
  AOI2BB1X1 U261 ( .A0N(n262), .A1N(n265), .B0(n197), .Y(n264) );
  INVX1 U262 ( .A(n151), .Y(n262) );
  NOR2X1 U263 ( .A(n156), .B(n252), .Y(n151) );
  MXI2X1 U264 ( .A(n266), .B(n267), .S0(n156), .Y(n677) );
  NAND2X1 U265 ( .A(count_r1_ram4x4[0]), .B(n152), .Y(n267) );
  AOI21X1 U266 ( .A0(n152), .A1(n252), .B0(n154), .Y(n266) );
  NAND4X1 U267 ( .A(n268), .B(n269), .C(n127), .D(n270), .Y(n154) );
  NAND2X1 U268 ( .A(n265), .B(n26), .Y(n268) );
  INVX1 U269 ( .A(n155), .Y(n152) );
  MXI2X1 U270 ( .A(n271), .B(n155), .S0(n252), .Y(n676) );
  AOI2BB2X1 U271 ( .B0(n269), .B1(n605), .A0N(n272), .A1N(n197), .Y(n155) );
  AOI211X1 U272 ( .A0(n273), .A1(full[1]), .B0(n274), .C0(n275), .Y(n272) );
  NOR2X1 U273 ( .A(n276), .B(n263), .Y(n271) );
  OAI211X1 U274 ( .A0(full[2]), .A1(n277), .B0(n269), .C0(n270), .Y(n263) );
  OAI211X1 U275 ( .A0(n224), .A1(n278), .B0(n279), .C0(n280), .Y(n269) );
  AOI32X1 U276 ( .A0(n605), .A1(n281), .A2(n282), .B0(n283), .B1(n26), .Y(n280) );
  NOR4BX1 U277 ( .AN(n79), .B(n203), .C(n136), .D(n84), .Y(n224) );
  OAI211X1 U278 ( .A0(n150), .A1(n284), .B0(n64), .C0(n285), .Y(n675) );
  MXI2X1 U279 ( .A(n286), .B(n287), .S0(n613), .Y(n285) );
  NOR2BX1 U280 ( .AN(n288), .B(n142), .Y(n287) );
  OAI2BB1X1 U281 ( .A0N(n142), .A1N(n288), .B0(n289), .Y(n286) );
  OAI211X1 U282 ( .A0(n252), .A1(n284), .B0(n64), .C0(n290), .Y(n674) );
  MXI2X1 U283 ( .A(n291), .B(n292), .S0(addr_ram4x4_4[2]), .Y(n290) );
  AND2X1 U284 ( .A(n244), .B(n288), .Y(n291) );
  OAI211X1 U285 ( .A0(n156), .A1(n284), .B0(n293), .C0(n294), .Y(n673) );
  AOI31X1 U286 ( .A0(n244), .A1(addr_ram4x4_4[2]), .A2(n288), .B0(n25), .Y(
        n294) );
  OAI21XL U287 ( .A0(n288), .A1(n292), .B0(addr_ram4x4_4[3]), .Y(n293) );
  OAI21XL U288 ( .A0(n244), .A1(n216), .B0(n289), .Y(n292) );
  INVX1 U289 ( .A(n295), .Y(n289) );
  OAI211X1 U290 ( .A0(n245), .A1(n296), .B0(n64), .C0(n297), .Y(n672) );
  MXI2X1 U291 ( .A(n298), .B(n299), .S0(n617), .Y(n297) );
  OAI211X1 U292 ( .A0(n150), .A1(n296), .B0(n64), .C0(n300), .Y(n671) );
  MXI2X1 U293 ( .A(n301), .B(n302), .S0(n616), .Y(n300) );
  NOR2X1 U294 ( .A(n617), .B(n303), .Y(n302) );
  OAI2BB1X1 U295 ( .A0N(n617), .A1N(n299), .B0(n304), .Y(n301) );
  OAI211X1 U296 ( .A0(n252), .A1(n296), .B0(n64), .C0(n305), .Y(n670) );
  MXI2X1 U297 ( .A(n306), .B(n307), .S0(addr_ram4x4_3[2]), .Y(n305) );
  NOR2BX1 U298 ( .AN(n308), .B(n303), .Y(n306) );
  OAI211X1 U299 ( .A0(n156), .A1(n296), .B0(n309), .C0(n310), .Y(n669) );
  AOI31X1 U300 ( .A0(n308), .A1(addr_ram4x4_3[2]), .A2(n299), .B0(n25), .Y(
        n310) );
  OAI21XL U301 ( .A0(n299), .A1(n307), .B0(addr_ram4x4_3[3]), .Y(n309) );
  OAI21XL U302 ( .A0(n308), .A1(n129), .B0(n304), .Y(n307) );
  INVX1 U303 ( .A(n298), .Y(n304) );
  NAND2X1 U304 ( .A(n235), .B(n127), .Y(n298) );
  OR2X1 U305 ( .A(n217), .B(full[1]), .Y(n127) );
  INVX1 U306 ( .A(n303), .Y(n299) );
  OAI21XL U307 ( .A0(n615), .A1(n236), .B0(n232), .Y(n303) );
  NAND2X1 U308 ( .A(n308), .B(addr_ram4x4_3[3]), .Y(n236) );
  NOR2X1 U309 ( .A(n616), .B(n617), .Y(n308) );
  OAI21XL U310 ( .A0(n605), .A1(n213), .B0(n235), .Y(n296) );
  NAND3X1 U311 ( .A(n279), .B(n217), .C(n311), .Y(n235) );
  OAI211X1 U312 ( .A0(n245), .A1(n312), .B0(n64), .C0(n313), .Y(n668) );
  MX2X1 U313 ( .A(n314), .B(n315), .S0(n628), .Y(n313) );
  OAI211X1 U314 ( .A0(n150), .A1(n312), .B0(n64), .C0(n316), .Y(n667) );
  MXI2X1 U315 ( .A(n317), .B(n318), .S0(n144), .Y(n316) );
  NOR2X1 U316 ( .A(n628), .B(n315), .Y(n318) );
  OAI21XL U317 ( .A0(addr_ram4x4_2[0]), .A1(n315), .B0(n314), .Y(n317) );
  INVX1 U318 ( .A(count_r2_ram4x4[1]), .Y(n150) );
  OAI211X1 U319 ( .A0(n252), .A1(n312), .B0(n64), .C0(n319), .Y(n666) );
  MXI2X1 U320 ( .A(n320), .B(n321), .S0(addr_ram4x4_2[2]), .Y(n319) );
  NOR2BX1 U321 ( .AN(n322), .B(n315), .Y(n320) );
  INVX1 U322 ( .A(count_r1_ram4x4[0]), .Y(n252) );
  OAI211X1 U323 ( .A0(n156), .A1(n312), .B0(n323), .C0(n324), .Y(n665) );
  AOI31X1 U324 ( .A0(n322), .A1(addr_ram4x4_2[2]), .A2(n325), .B0(n25), .Y(
        n324) );
  OAI21XL U325 ( .A0(n325), .A1(n321), .B0(addr_ram4x4_2[3]), .Y(n323) );
  OAI21XL U326 ( .A0(n322), .A1(n315), .B0(n314), .Y(n321) );
  NOR2X1 U327 ( .A(n276), .B(n228), .Y(n314) );
  INVX1 U328 ( .A(n326), .Y(n228) );
  INVX1 U329 ( .A(n325), .Y(n315) );
  AOI21X1 U330 ( .A0(addr_ram4x4_2[2]), .A1(n229), .B0(n217), .Y(n325) );
  AND2X1 U331 ( .A(n322), .B(addr_ram4x4_2[3]), .Y(n229) );
  NOR2X1 U332 ( .A(n144), .B(n628), .Y(n322) );
  NAND2X1 U333 ( .A(n326), .B(n327), .Y(n312) );
  OAI21XL U334 ( .A0(n211), .A1(n165), .B0(n87), .Y(n327) );
  OAI221XL U335 ( .A0(n328), .A1(n87), .B0(n329), .B1(n197), .C0(n64), .Y(n326) );
  INVX1 U336 ( .A(count_r1_ram4x4[1]), .Y(n156) );
  OAI21XL U337 ( .A0(n330), .A1(n331), .B0(n332), .Y(n664) );
  OAI21XL U338 ( .A0(n47), .A1(n330), .B0(n332), .Y(n663) );
  INVX1 U339 ( .A(ram8x8_r_ready), .Y(n47) );
  NAND3X1 U340 ( .A(n333), .B(n165), .C(n256), .Y(n662) );
  NAND2X1 U341 ( .A(en_ram4x4_1), .B(n334), .Y(n333) );
  NAND3X1 U342 ( .A(n335), .B(n217), .C(n336), .Y(n661) );
  NAND2X1 U343 ( .A(en_ram4x4_2), .B(n334), .Y(n335) );
  NAND4X1 U344 ( .A(n311), .B(n337), .C(n198), .D(n129), .Y(n660) );
  NAND2X1 U345 ( .A(en_ram4x4_3), .B(n334), .Y(n337) );
  NAND4X1 U346 ( .A(n338), .B(n339), .C(n216), .D(n240), .Y(n659) );
  NAND2X1 U347 ( .A(en_ram4x4_4), .B(n334), .Y(n339) );
  OAI2BB1X1 U348 ( .A0N(ram4x4_1_ready), .A1N(n334), .B0(n256), .Y(n658) );
  AOI2BB1X1 U349 ( .A0N(n340), .A1N(n87), .B0(n93), .Y(n256) );
  AOI22X1 U350 ( .A0(n136), .A1(n341), .B0(n282), .B1(full[3]), .Y(n340) );
  NOR3X1 U351 ( .A(rd_num[1]), .B(rd_num[2]), .C(rd_num[0]), .Y(n136) );
  OAI2BB1X1 U352 ( .A0N(ram4x4_2_ready), .A1N(n334), .B0(n336), .Y(n657) );
  AOI2BB2X1 U353 ( .B0(full[2]), .B1(n214), .A0N(n328), .A1N(n87), .Y(n336) );
  AOI22X1 U354 ( .A0(n282), .A1(n275), .B0(n341), .B1(n84), .Y(n328) );
  AND3X1 U355 ( .A(n210), .B(n122), .C(rd_num[0]), .Y(n84) );
  NAND3X1 U356 ( .A(n342), .B(n198), .C(n311), .Y(n656) );
  AOI21X1 U357 ( .A0(n223), .A1(n203), .B0(n343), .Y(n311) );
  NOR4BX1 U358 ( .AN(n265), .B(n344), .C(n345), .D(n87), .Y(n343) );
  NOR3X1 U359 ( .A(rd_num[0]), .B(rd_num[2]), .C(n210), .Y(n203) );
  INVX1 U360 ( .A(rd_num[1]), .Y(n210) );
  INVX1 U361 ( .A(n213), .Y(n198) );
  NOR2X1 U362 ( .A(n217), .B(n345), .Y(n213) );
  NAND2X1 U363 ( .A(n273), .B(n26), .Y(n217) );
  NAND2X1 U364 ( .A(ram4x4_3_ready), .B(n334), .Y(n342) );
  NAND3X1 U365 ( .A(n346), .B(n240), .C(n338), .Y(n655) );
  INVX1 U366 ( .A(n125), .Y(n240) );
  NAND2X1 U367 ( .A(ram4x4_4_ready), .B(n334), .Y(n346) );
  INVX1 U368 ( .A(n330), .Y(n334) );
  NAND2X1 U369 ( .A(n347), .B(n348), .Y(n330) );
  OAI2BB2X1 U370 ( .B0(n610), .B1(n181), .A0N(mode_out[1]), .A1N(n347), .Y(
        n654) );
  NAND2X1 U371 ( .A(n349), .B(n350), .Y(n653) );
  AOI31X1 U372 ( .A0(n26), .A1(n91), .A2(n351), .B0(n67), .Y(n350) );
  AOI22X1 U373 ( .A0(mode_out[0]), .A1(n347), .B0(n66), .B1(mode_r_0_), .Y(
        n349) );
  OAI31X1 U374 ( .A0(n120), .A1(n282), .A2(n341), .B0(n348), .Y(n347) );
  NOR2X1 U375 ( .A(n54), .B(n25), .Y(n348) );
  NAND2X1 U376 ( .A(n352), .B(n353), .Y(n652) );
  AOI222X1 U377 ( .A0(N1362), .A1(n50), .B0(count_w[1]), .B1(n51), .C0(N1400), 
        .C1(n52), .Y(n353) );
  AOI222X1 U378 ( .A0(N980), .A1(n26), .B0(N852), .B1(n53), .C0(N725), .C1(n54), .Y(n352) );
  NAND2X1 U379 ( .A(n354), .B(n355), .Y(n651) );
  AOI222X1 U380 ( .A0(N1363), .A1(n50), .B0(count_w[2]), .B1(n51), .C0(N1401), 
        .C1(n52), .Y(n355) );
  AOI222X1 U381 ( .A0(N981), .A1(n26), .B0(N853), .B1(n53), .C0(N726), .C1(n54), .Y(n354) );
  NAND2X1 U382 ( .A(n356), .B(n357), .Y(n650) );
  AOI222X1 U383 ( .A0(N1364), .A1(n50), .B0(count_w[3]), .B1(n51), .C0(N1402), 
        .C1(n52), .Y(n357) );
  AOI222X1 U384 ( .A0(N982), .A1(n26), .B0(N854), .B1(n53), .C0(N727), .C1(n54), .Y(n356) );
  NAND2X1 U385 ( .A(n358), .B(n359), .Y(n649) );
  AOI222X1 U386 ( .A0(N1365), .A1(n50), .B0(n51), .B1(count_w[4]), .C0(N1403), 
        .C1(n52), .Y(n359) );
  AOI222X1 U387 ( .A0(N983), .A1(n26), .B0(N855), .B1(n53), .C0(N728), .C1(n54), .Y(n358) );
  NAND2X1 U388 ( .A(n360), .B(n361), .Y(n648) );
  AOI222X1 U389 ( .A0(N1366), .A1(n50), .B0(n51), .B1(count_w[5]), .C0(N1404), 
        .C1(n52), .Y(n361) );
  AOI222X1 U390 ( .A0(N984), .A1(n26), .B0(N856), .B1(n53), .C0(N729), .C1(n54), .Y(n360) );
  NAND2X1 U391 ( .A(n362), .B(n363), .Y(n647) );
  AOI222X1 U392 ( .A0(N1367), .A1(n50), .B0(n51), .B1(count_w[6]), .C0(N1405), 
        .C1(n52), .Y(n363) );
  AOI222X1 U393 ( .A0(N985), .A1(n26), .B0(N857), .B1(n53), .C0(N730), .C1(n54), .Y(n362) );
  NAND2X1 U394 ( .A(n364), .B(n365), .Y(n646) );
  AOI222X1 U395 ( .A0(N1368), .A1(n50), .B0(count_w[7]), .B1(n51), .C0(N1406), 
        .C1(n52), .Y(n365) );
  AOI222X1 U396 ( .A0(N986), .A1(n26), .B0(N858), .B1(n53), .C0(N731), .C1(n54), .Y(n364) );
  NAND2X1 U397 ( .A(n366), .B(n367), .Y(n645) );
  AOI222X1 U398 ( .A0(N1369), .A1(n50), .B0(count_w[8]), .B1(n51), .C0(N1407), 
        .C1(n52), .Y(n367) );
  AOI222X1 U399 ( .A0(N987), .A1(n26), .B0(N859), .B1(n53), .C0(N732), .C1(n54), .Y(n366) );
  OAI211X1 U400 ( .A0(n37), .A1(n258), .B0(n369), .C0(n370), .Y(n644) );
  AOI22X1 U401 ( .A0(N760), .A1(n371), .B0(N830), .B1(n372), .Y(n370) );
  AOI21X1 U402 ( .A0(n373), .A1(N830), .B0(n25), .Y(n369) );
  OAI211X1 U403 ( .A0(n36), .A1(n258), .B0(n374), .C0(n375), .Y(n643) );
  AOI22X1 U404 ( .A0(N761), .A1(n371), .B0(N831), .B1(n372), .Y(n375) );
  AOI21X1 U405 ( .A0(n373), .A1(N831), .B0(n25), .Y(n374) );
  OAI211X1 U406 ( .A0(n632), .A1(n258), .B0(n376), .C0(n377), .Y(n642) );
  AOI22X1 U407 ( .A0(N762), .A1(n371), .B0(N1074), .B1(n372), .Y(n377) );
  AOI21X1 U408 ( .A0(n373), .A1(N1067), .B0(n25), .Y(n376) );
  OAI211X1 U409 ( .A0(n631), .A1(n258), .B0(n378), .C0(n379), .Y(n641) );
  AOI22X1 U410 ( .A0(N763), .A1(n371), .B0(n372), .B1(N1075), .Y(n379) );
  AOI21X1 U411 ( .A0(n373), .A1(N1068), .B0(n25), .Y(n378) );
  OAI211X1 U412 ( .A0(n630), .A1(n258), .B0(n380), .C0(n381), .Y(n640) );
  AOI22X1 U413 ( .A0(N764), .A1(n371), .B0(n372), .B1(N1076), .Y(n381) );
  AOI21X1 U414 ( .A0(n373), .A1(N1069), .B0(n25), .Y(n380) );
  OAI211X1 U415 ( .A0(n629), .A1(n258), .B0(n382), .C0(n383), .Y(n639) );
  AOI22X1 U416 ( .A0(N765), .A1(n371), .B0(n372), .B1(N1077), .Y(n383) );
  AOI21X1 U417 ( .A0(n373), .A1(N1070), .B0(n25), .Y(n382) );
  OAI211X1 U418 ( .A0(n148), .A1(n258), .B0(n384), .C0(n385), .Y(n638) );
  AOI22X1 U419 ( .A0(N766), .A1(n371), .B0(n372), .B1(N1078), .Y(n385) );
  AOI21X1 U420 ( .A0(n373), .A1(N1071), .B0(n25), .Y(n384) );
  NOR2X1 U421 ( .A(n386), .B(n130), .Y(n373) );
  OAI211X1 U422 ( .A0(n149), .A1(n258), .B0(n64), .C0(n387), .Y(n637) );
  AOI22X1 U423 ( .A0(N767), .A1(n371), .B0(n372), .B1(N1079), .Y(n387) );
  NOR2X1 U424 ( .A(n386), .B(n215), .Y(n372) );
  OAI22X1 U425 ( .A0(n388), .A1(n389), .B0(N758), .B1(n390), .Y(n371) );
  AOI211X1 U426 ( .A0(n50), .A1(n391), .B0(n52), .C0(n392), .Y(n389) );
  AOI31X1 U427 ( .A0(n630), .A1(n629), .A2(n393), .B0(n199), .Y(n392) );
  NOR3X1 U428 ( .A(addr_ram8x8_w[7]), .B(n394), .C(addr_ram8x8_w[6]), .Y(n393)
         );
  XNOR2X1 U429 ( .A(ram), .B(ram_write), .Y(n391) );
  OAI211X1 U430 ( .A0(n395), .A1(n396), .B0(n397), .C0(n398), .Y(ram_write) );
  AOI21X1 U431 ( .A0(n399), .A1(n400), .B0(n401), .Y(n398) );
  MXI2X1 U432 ( .A(n402), .B(n403), .S0(n404), .Y(n401) );
  NAND2X1 U433 ( .A(n405), .B(n406), .Y(n403) );
  AOI21X1 U434 ( .A0(n406), .A1(n407), .B0(n408), .Y(n402) );
  INVX1 U435 ( .A(next_state[2]), .Y(n397) );
  NOR3X1 U436 ( .A(n410), .B(addr_ram8x8_w[6]), .C(addr_ram8x8_w[7]), .Y(n388)
         );
  OR3XL U437 ( .A(n629), .B(n630), .C(n394), .Y(n410) );
  OR4X1 U438 ( .A(n631), .B(n632), .C(n36), .D(n37), .Y(n394) );
  INVX1 U439 ( .A(n93), .Y(n199) );
  NOR2X1 U440 ( .A(n351), .B(n197), .Y(n93) );
  NAND2X1 U441 ( .A(n274), .B(full[1]), .Y(n351) );
  INVX1 U442 ( .A(n411), .Y(n274) );
  OAI22X1 U443 ( .A0(n412), .A1(n194), .B0(n413), .B1(n414), .Y(n603) );
  AOI21X1 U444 ( .A0(n604), .A1(n415), .B0(n195), .Y(n413) );
  OAI21XL U445 ( .A0(count_r1[1]), .A1(n194), .B0(n192), .Y(n195) );
  AOI21X1 U446 ( .A0(n635), .A1(n604), .B0(n178), .Y(n192) );
  INVX1 U447 ( .A(n636), .Y(n178) );
  INVX1 U448 ( .A(n194), .Y(n604) );
  NAND2X1 U449 ( .A(n636), .B(n179), .Y(n194) );
  OAI222XL U450 ( .A0(n184), .A1(n190), .B0(n189), .B1(n188), .C0(N783), .C1(
        n181), .Y(n179) );
  INVX1 U451 ( .A(n416), .Y(n188) );
  OAI21XL U452 ( .A0(n197), .A1(n130), .B0(n120), .Y(n416) );
  NAND2X1 U453 ( .A(n605), .B(n417), .Y(n120) );
  NOR2X1 U454 ( .A(n193), .B(count_r1[3]), .Y(n189) );
  NAND3X1 U455 ( .A(n415), .B(count_r1[0]), .C(count_r1[1]), .Y(n193) );
  INVX1 U456 ( .A(count_r1[2]), .Y(n415) );
  AOI21X1 U457 ( .A0(n26), .A1(n130), .B0(n67), .Y(n190) );
  INVX1 U458 ( .A(n215), .Y(n130) );
  NOR3X1 U459 ( .A(n345), .B(n91), .C(n283), .Y(n215) );
  INVX1 U460 ( .A(n412), .Y(n184) );
  NAND2BX1 U461 ( .AN(n62), .B(n386), .Y(n636) );
  NAND3X1 U462 ( .A(n26), .B(n411), .C(n418), .Y(n386) );
  OAI211X1 U463 ( .A0(n273), .A1(n275), .B0(full[0]), .C0(full[1]), .Y(n418)
         );
  NOR2X1 U464 ( .A(n211), .B(full[3]), .Y(n275) );
  NOR2X1 U465 ( .A(n167), .B(full[2]), .Y(n273) );
  NAND2X1 U466 ( .A(full[0]), .B(n329), .Y(n411) );
  AOI211X1 U467 ( .A0(n223), .A1(n83), .B0(n67), .C0(n66), .Y(n332) );
  NOR3X1 U468 ( .A(next_state[2]), .B(next_state[4]), .C(n53), .Y(n181) );
  OAI21XL U469 ( .A0(n419), .A1(n420), .B0(n421), .Y(next_state[4]) );
  NAND4BXL U470 ( .AN(state[2]), .B(state[4]), .C(n422), .D(n423), .Y(n421) );
  OAI21XL U471 ( .A0(n395), .A1(n420), .B0(n424), .Y(next_state[2]) );
  NAND4BXL U472 ( .AN(state[4]), .B(state[2]), .C(n422), .D(n423), .Y(n424) );
  NOR3X1 U473 ( .A(rd_num[0]), .B(rd_num[1]), .C(n122), .Y(n83) );
  NAND4X1 U474 ( .A(count_r1[2]), .B(count_r1[1]), .C(n414), .D(count_r1[0]), 
        .Y(n412) );
  INVX1 U475 ( .A(count_r1[3]), .Y(n414) );
  OAI211X1 U476 ( .A0(n245), .A1(n284), .B0(n64), .C0(n425), .Y(n602) );
  MXI2X1 U477 ( .A(n295), .B(n288), .S0(n142), .Y(n425) );
  AOI31X1 U478 ( .A0(n244), .A1(addr_ram4x4_4[2]), .A2(addr_ram4x4_4[3]), .B0(
        n216), .Y(n288) );
  NOR2X1 U479 ( .A(n142), .B(n613), .Y(n244) );
  NAND2X1 U480 ( .A(n239), .B(n270), .Y(n295) );
  INVX1 U481 ( .A(n220), .Y(n270) );
  NOR2X1 U482 ( .A(n129), .B(full[0]), .Y(n220) );
  OAI21XL U483 ( .A0(n605), .A1(n125), .B0(n239), .Y(n284) );
  NAND3X1 U484 ( .A(n279), .B(n216), .C(n338), .Y(n239) );
  AOI32X1 U485 ( .A0(n426), .A1(full[0]), .A2(n282), .B0(n223), .B1(n96), .Y(
        n338) );
  INVX1 U486 ( .A(n79), .Y(n96) );
  NAND3X1 U487 ( .A(rd_num[0]), .B(n122), .C(rd_num[1]), .Y(n79) );
  INVX1 U488 ( .A(rd_num[2]), .Y(n122) );
  INVX1 U489 ( .A(n278), .Y(n223) );
  NAND2X1 U490 ( .A(n341), .B(n605), .Y(n278) );
  AND3X1 U491 ( .A(n344), .B(n427), .C(n417), .Y(n341) );
  NAND2X1 U492 ( .A(n423), .B(n91), .Y(n417) );
  INVX1 U493 ( .A(n282), .Y(n344) );
  NOR2X1 U494 ( .A(n423), .B(ram8_4), .Y(n282) );
  AND3X1 U495 ( .A(n605), .B(n345), .C(n265), .Y(n426) );
  INVX1 U496 ( .A(n131), .Y(n216) );
  NOR3X1 U497 ( .A(n345), .B(n197), .C(n283), .Y(n131) );
  NAND2X1 U498 ( .A(n329), .B(n428), .Y(n283) );
  NOR2X1 U499 ( .A(n232), .B(n25), .Y(n279) );
  MXI2X1 U500 ( .A(n409), .B(n433), .S0(n434), .Y(n432) );
  NOR4BX1 U501 ( .AN(n431), .B(n435), .C(n400), .D(n406), .Y(n433) );
  INVX1 U502 ( .A(n436), .Y(n406) );
  NAND3X1 U503 ( .A(n437), .B(n438), .C(n429), .Y(n435) );
  NAND2X1 U504 ( .A(n422), .B(n439), .Y(n431) );
  XOR2X1 U505 ( .A(state[4]), .B(state[2]), .Y(n439) );
  NOR4BX1 U506 ( .AN(n440), .B(state[0]), .C(state[1]), .D(state[3]), .Y(n422)
         );
  INVX1 U507 ( .A(n129), .Y(n232) );
  NOR2X1 U508 ( .A(n129), .B(n428), .Y(n125) );
  NAND2BX1 U509 ( .AN(n277), .B(n329), .Y(n129) );
  INVX1 U510 ( .A(count_r2_ram4x4[0]), .Y(n245) );
  MX2X1 U511 ( .A(mode_w[1]), .B(mode[1]), .S0(start), .Y(n601) );
  MX2X1 U512 ( .A(mode_w[0]), .B(mode[0]), .S0(start), .Y(n600) );
  MXI2X1 U513 ( .A(n441), .B(n331), .S0(n44), .Y(en_ram8x8_2) );
  MXI2X1 U514 ( .A(n331), .B(n441), .S0(n44), .Y(en_ram8x8_1) );
  INVX1 U515 ( .A(en_ram8x8_w), .Y(n441) );
  INVX1 U516 ( .A(en_ram8x8_r), .Y(n331) );
  MXI2X1 U517 ( .A(n629), .B(n114), .S0(n44), .Y(addr_ram8x8_2[5]) );
  MXI2X1 U518 ( .A(n630), .B(n111), .S0(n44), .Y(addr_ram8x8_2[4]) );
  MXI2X1 U519 ( .A(n631), .B(n108), .S0(n44), .Y(addr_ram8x8_2[3]) );
  MXI2X1 U520 ( .A(n632), .B(n105), .S0(n44), .Y(addr_ram8x8_2[2]) );
  MXI2X1 U521 ( .A(n36), .B(n102), .S0(n44), .Y(addr_ram8x8_2[1]) );
  MXI2X1 U522 ( .A(n37), .B(n98), .S0(n44), .Y(addr_ram8x8_2[0]) );
  MXI2X1 U523 ( .A(n114), .B(n629), .S0(n44), .Y(addr_ram8x8_1[5]) );
  MXI2X1 U524 ( .A(n111), .B(n630), .S0(n44), .Y(addr_ram8x8_1[4]) );
  MXI2X1 U525 ( .A(n108), .B(n631), .S0(n44), .Y(addr_ram8x8_1[3]) );
  MXI2X1 U526 ( .A(n105), .B(n632), .S0(n44), .Y(addr_ram8x8_1[2]) );
  MXI2X1 U527 ( .A(n102), .B(n36), .S0(n44), .Y(addr_ram8x8_1[1]) );
  MXI2X1 U528 ( .A(n98), .B(n37), .S0(n44), .Y(addr_ram8x8_1[0]) );
  XNOR2X1 U529 ( .A(count_w[4]), .B(N716), .Y(n444) );
  XNOR2X1 U530 ( .A(count_w[5]), .B(N717), .Y(n443) );
  XNOR2X1 U531 ( .A(count_w[6]), .B(N718), .Y(n442) );
  AOI31X1 U532 ( .A0(n446), .A1(n437), .A2(n447), .B0(n399), .Y(N593) );
  NOR2X1 U533 ( .A(n448), .B(n449), .Y(n447) );
  INVX1 U534 ( .A(n400), .Y(n446) );
  NAND3BX1 U535 ( .AN(N1888), .B(n450), .C(n368), .Y(N1838) );
  AOI2BB1X1 U536 ( .A0N(n451), .A1N(n87), .B0(n259), .Y(n368) );
  INVX1 U537 ( .A(n390), .Y(n259) );
  NOR2X1 U538 ( .A(n54), .B(n53), .Y(n390) );
  OAI32X1 U539 ( .A0(n452), .A1(n453), .A2(n437), .B0(n419), .B1(n396), .Y(
        next_state[6]) );
  AOI21X1 U540 ( .A0(n448), .A1(ram_write_reg), .B0(n400), .Y(n419) );
  NAND2X1 U541 ( .A(n454), .B(n455), .Y(n400) );
  OAI32X1 U542 ( .A0(n455), .A1(n453), .A2(n452), .B0(n395), .B1(n396), .Y(
        next_state[3]) );
  AOI211X1 U543 ( .A0(n404), .A1(n448), .B0(n456), .C0(n449), .Y(n395) );
  INVX1 U544 ( .A(n438), .Y(n449) );
  INVX1 U545 ( .A(n437), .Y(n456) );
  NOR2X1 U546 ( .A(n429), .B(n489), .Y(n448) );
  INVX1 U547 ( .A(ram_write_reg), .Y(n404) );
  OAI222XL U548 ( .A0(n452), .A1(n438), .B0(n437), .B1(n457), .C0(n409), .C1(
        n434), .Y(n607) );
  NAND3X1 U549 ( .A(n458), .B(n440), .C(state[0]), .Y(n434) );
  OAI22X1 U550 ( .A0(n452), .A1(n454), .B0(n455), .B1(n457), .Y(n606) );
  INVX1 U551 ( .A(n453), .Y(n457) );
  NOR2X1 U552 ( .A(n423), .B(n459), .Y(n453) );
  NAND4BXL U553 ( .AN(count_r1[1]), .B(n635), .C(n460), .D(n461), .Y(n423) );
  NOR4BX1 U554 ( .AN(n58), .B(N1074), .C(N831), .D(N830), .Y(n461) );
  INVX1 U555 ( .A(count_r2_3_), .Y(n58) );
  NOR2X1 U556 ( .A(count_r1[3]), .B(count_r1[2]), .Y(n460) );
  NAND2X1 U557 ( .A(n399), .B(n462), .Y(n452) );
  INVX1 U558 ( .A(n463), .Y(n399) );
  OAI21XL U559 ( .A0(n489), .A1(n462), .B0(n408), .Y(n464) );
  INVX1 U560 ( .A(n405), .Y(n407) );
  NOR2X1 U561 ( .A(start), .B(n196), .Y(n451) );
  NAND3X1 U562 ( .A(n329), .B(n26), .C(full[1]), .Y(n450) );
  OAI221XL U563 ( .A0(n329), .A1(n277), .B0(full[0]), .B1(n197), .C0(n128), 
        .Y(N1888) );
  INVX1 U564 ( .A(n276), .Y(n128) );
  NOR2X1 U565 ( .A(n165), .B(full[2]), .Y(n276) );
  NOR2X1 U566 ( .A(full[3]), .B(n197), .Y(n214) );
  NAND2X1 U567 ( .A(n26), .B(n345), .Y(n277) );
  NAND3X1 U568 ( .A(n459), .B(n466), .C(start), .Y(n462) );
  AOI211X1 U569 ( .A0(n408), .A1(n196), .B0(n467), .C0(n468), .Y(n465) );
  INVX1 U570 ( .A(n455), .Y(n468) );
  NAND3BX1 U571 ( .AN(state[1]), .B(n469), .C(state[3]), .Y(n455) );
  NAND3X1 U572 ( .A(n437), .B(n438), .C(n454), .Y(n467) );
  NAND4X1 U573 ( .A(state[5]), .B(n470), .C(n471), .D(n472), .Y(n454) );
  NAND3BX1 U574 ( .AN(state[3]), .B(n469), .C(state[1]), .Y(n438) );
  NOR4BX1 U575 ( .AN(n440), .B(state[0]), .C(state[2]), .D(state[4]), .Y(n469)
         );
  NOR4BX1 U576 ( .AN(n471), .B(state[5]), .C(state[7]), .D(state[8]), .Y(n440)
         );
  NAND4X1 U577 ( .A(state[6]), .B(n470), .C(n473), .D(n472), .Y(n437) );
  INVX1 U578 ( .A(state[7]), .Y(n472) );
  AOI211X1 U579 ( .A0(n463), .A1(n196), .B0(n474), .C0(n429), .Y(n408) );
  NAND4BXL U580 ( .AN(state[0]), .B(n458), .C(state[8]), .D(n475), .Y(n429) );
  NOR3X1 U581 ( .A(state[5]), .B(state[7]), .C(state[6]), .Y(n475) );
  INVX1 U582 ( .A(n430), .Y(n474) );
  NAND2X1 U583 ( .A(n476), .B(n489), .Y(n430) );
  MXI2X1 U584 ( .A(n427), .B(n281), .S0(n91), .Y(n476) );
  INVX1 U585 ( .A(ram8_4), .Y(n91) );
  NAND3X1 U586 ( .A(n428), .B(n345), .C(n265), .Y(n281) );
  NOR2X1 U587 ( .A(full[2]), .B(full[3]), .Y(n265) );
  INVX1 U588 ( .A(full[1]), .Y(n345) );
  INVX1 U589 ( .A(full[0]), .Y(n428) );
  NAND3X1 U590 ( .A(n73), .B(n74), .C(rd_cnt[2]), .Y(n427) );
  INVX1 U591 ( .A(rd_cnt[1]), .Y(n74) );
  INVX1 U592 ( .A(rd_cnt[0]), .Y(n73) );
  NAND2X1 U593 ( .A(n396), .B(n420), .Y(n463) );
  NAND2X1 U594 ( .A(n459), .B(n409), .Y(n420) );
  INVX1 U595 ( .A(start), .Y(n409) );
  NAND3BX1 U596 ( .AN(n466), .B(n459), .C(start), .Y(n396) );
  INVX1 U597 ( .A(n477), .Y(n459) );
  OAI31X1 U598 ( .A0(n478), .A1(mode[0]), .A2(n490), .B0(n479), .Y(n466) );
  NAND4X1 U599 ( .A(state[7]), .B(n470), .C(n473), .D(n471), .Y(n436) );
  INVX1 U600 ( .A(state[6]), .Y(n471) );
  INVX1 U601 ( .A(state[5]), .Y(n473) );
  NOR3BX1 U602 ( .AN(n458), .B(state[0]), .C(state[8]), .Y(n470) );
  NOR4X1 U603 ( .A(state[3]), .B(state[1]), .C(state[2]), .D(state[4]), .Y(
        n458) );
  AOI21X1 U604 ( .A0(n480), .A1(start), .B0(n477), .Y(n405) );
  NAND4X1 U605 ( .A(n481), .B(n482), .C(n483), .D(n445), .Y(n477) );
  NOR4BX1 U606 ( .AN(n484), .B(count_w[1]), .C(count_w[2]), .D(count_w[0]), 
        .Y(n445) );
  NOR3X1 U607 ( .A(count_w[3]), .B(count_w[8]), .C(count_w[7]), .Y(n484) );
  XNOR2X1 U608 ( .A(count_w[4]), .B(N329), .Y(n483) );
  XNOR2X1 U609 ( .A(count_w[5]), .B(N330), .Y(n482) );
  XNOR2X1 U610 ( .A(count_w[6]), .B(N331), .Y(n481) );
  AOI31X1 U611 ( .A0(n479), .A1(n490), .A2(mode[0]), .B0(n478), .Y(n480) );
  NOR2X1 U612 ( .A(n485), .B(mode_w[1]), .Y(n478) );
  INVX1 U613 ( .A(mode_w[0]), .Y(n490) );
  NAND2X1 U614 ( .A(mode_w[1]), .B(n485), .Y(n479) );
  INVX1 U615 ( .A(mode[1]), .Y(n485) );
  NOR2X1 U616 ( .A(n167), .B(n211), .Y(n329) );
  INVX1 U617 ( .A(full[2]), .Y(n211) );
  INVX1 U618 ( .A(full[3]), .Y(n167) );
endmodule


module mem8x8_0 ( clk, rstn, en, wr_rd, addr, din, dout );
  input [5:0] addr;
  input [15:0] din;
  output [15:0] dout;
  input clk, rstn, en, wr_rd;
  wire   N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98,
         N99, N100, n23, n24, n26, n28, n30, n32, n34, n36, n38, n39, n41, n50,
         n59, n68, n77, n86, n95, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
         n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
         n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
         n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
         n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
         n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
         n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
         n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n25, n27, n29, n31, n33, n35, n37, n40, n42, n43, n44, n45,
         n46, n47, n48, n49, n51, n52, n53, n54, n55, n56, n57, n58, n60, n61,
         n62, n63, n64, n65, n66, n67, n69, n70, n71, n72, n73, n74, n75, n76,
         n78, n79, n80, n81, n82, n83, n84, n85, n87, n88, n89, n90, n91, n92,
         n93, n94, n96, n97, n98, n99, n100, n101, n102, n1128, n1129, n1130,
         n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
         n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
         n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
         n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
         n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
         n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
         n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
         n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
         n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
         n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
         n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
         n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
         n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
         n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
         n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
         n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
         n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
         n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
         n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
         n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
         n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
         n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
         n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
         n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
         n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
         n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
         n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
         n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
         n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
         n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
         n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
         n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
         n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
         n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
         n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
         n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
         n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
         n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
         n1511, n1512;
  wire   [1023:0] memory;

  DFFRHQX1 memory_reg_1__15_ ( .D(n1111), .CK(clk), .RN(rstn), .Q(memory[1007]) );
  DFFRHQX1 memory_reg_1__14_ ( .D(n1110), .CK(clk), .RN(rstn), .Q(memory[1006]) );
  DFFRHQX1 memory_reg_1__13_ ( .D(n1109), .CK(clk), .RN(rstn), .Q(memory[1005]) );
  DFFRHQX1 memory_reg_1__12_ ( .D(n1108), .CK(clk), .RN(rstn), .Q(memory[1004]) );
  DFFRHQX1 memory_reg_1__11_ ( .D(n1107), .CK(clk), .RN(rstn), .Q(memory[1003]) );
  DFFRHQX1 memory_reg_1__10_ ( .D(n1106), .CK(clk), .RN(rstn), .Q(memory[1002]) );
  DFFRHQX1 memory_reg_1__9_ ( .D(n1105), .CK(clk), .RN(rstn), .Q(memory[1001])
         );
  DFFRHQX1 memory_reg_1__8_ ( .D(n1104), .CK(clk), .RN(rstn), .Q(memory[1000])
         );
  DFFRHQX1 memory_reg_1__7_ ( .D(n1103), .CK(clk), .RN(rstn), .Q(memory[999])
         );
  DFFRHQX1 memory_reg_1__6_ ( .D(n1102), .CK(clk), .RN(rstn), .Q(memory[998])
         );
  DFFRHQX1 memory_reg_1__5_ ( .D(n1101), .CK(clk), .RN(rstn), .Q(memory[997])
         );
  DFFRHQX1 memory_reg_1__4_ ( .D(n1100), .CK(clk), .RN(rstn), .Q(memory[996])
         );
  DFFRHQX1 memory_reg_1__3_ ( .D(n1099), .CK(clk), .RN(rstn), .Q(memory[995])
         );
  DFFRHQX1 memory_reg_1__2_ ( .D(n1098), .CK(clk), .RN(rstn), .Q(memory[994])
         );
  DFFRHQX1 memory_reg_1__1_ ( .D(n1097), .CK(clk), .RN(rstn), .Q(memory[993])
         );
  DFFRHQX1 memory_reg_1__0_ ( .D(n1096), .CK(clk), .RN(rstn), .Q(memory[992])
         );
  DFFRHQX1 memory_reg_5__15_ ( .D(n1047), .CK(clk), .RN(rstn), .Q(memory[943])
         );
  DFFRHQX1 memory_reg_5__14_ ( .D(n1046), .CK(clk), .RN(rstn), .Q(memory[942])
         );
  DFFRHQX1 memory_reg_5__13_ ( .D(n1045), .CK(clk), .RN(rstn), .Q(memory[941])
         );
  DFFRHQX1 memory_reg_5__12_ ( .D(n1044), .CK(clk), .RN(rstn), .Q(memory[940])
         );
  DFFRHQX1 memory_reg_5__11_ ( .D(n1043), .CK(clk), .RN(rstn), .Q(memory[939])
         );
  DFFRHQX1 memory_reg_5__10_ ( .D(n1042), .CK(clk), .RN(rstn), .Q(memory[938])
         );
  DFFRHQX1 memory_reg_5__9_ ( .D(n1041), .CK(clk), .RN(rstn), .Q(memory[937])
         );
  DFFRHQX1 memory_reg_5__8_ ( .D(n1040), .CK(clk), .RN(rstn), .Q(memory[936])
         );
  DFFRHQX1 memory_reg_5__7_ ( .D(n1039), .CK(clk), .RN(rstn), .Q(memory[935])
         );
  DFFRHQX1 memory_reg_5__6_ ( .D(n1038), .CK(clk), .RN(rstn), .Q(memory[934])
         );
  DFFRHQX1 memory_reg_5__5_ ( .D(n1037), .CK(clk), .RN(rstn), .Q(memory[933])
         );
  DFFRHQX1 memory_reg_5__4_ ( .D(n1036), .CK(clk), .RN(rstn), .Q(memory[932])
         );
  DFFRHQX1 memory_reg_5__3_ ( .D(n1035), .CK(clk), .RN(rstn), .Q(memory[931])
         );
  DFFRHQX1 memory_reg_5__2_ ( .D(n1034), .CK(clk), .RN(rstn), .Q(memory[930])
         );
  DFFRHQX1 memory_reg_5__1_ ( .D(n1033), .CK(clk), .RN(rstn), .Q(memory[929])
         );
  DFFRHQX1 memory_reg_5__0_ ( .D(n1032), .CK(clk), .RN(rstn), .Q(memory[928])
         );
  DFFRHQX1 memory_reg_9__15_ ( .D(n983), .CK(clk), .RN(rstn), .Q(memory[879])
         );
  DFFRHQX1 memory_reg_9__14_ ( .D(n982), .CK(clk), .RN(rstn), .Q(memory[878])
         );
  DFFRHQX1 memory_reg_9__13_ ( .D(n981), .CK(clk), .RN(rstn), .Q(memory[877])
         );
  DFFRHQX1 memory_reg_9__12_ ( .D(n980), .CK(clk), .RN(rstn), .Q(memory[876])
         );
  DFFRHQX1 memory_reg_9__11_ ( .D(n979), .CK(clk), .RN(rstn), .Q(memory[875])
         );
  DFFRHQX1 memory_reg_9__10_ ( .D(n978), .CK(clk), .RN(rstn), .Q(memory[874])
         );
  DFFRHQX1 memory_reg_9__9_ ( .D(n977), .CK(clk), .RN(rstn), .Q(memory[873])
         );
  DFFRHQX1 memory_reg_9__8_ ( .D(n976), .CK(clk), .RN(rstn), .Q(memory[872])
         );
  DFFRHQX1 memory_reg_9__7_ ( .D(n975), .CK(clk), .RN(rstn), .Q(memory[871])
         );
  DFFRHQX1 memory_reg_9__6_ ( .D(n974), .CK(clk), .RN(rstn), .Q(memory[870])
         );
  DFFRHQX1 memory_reg_9__5_ ( .D(n973), .CK(clk), .RN(rstn), .Q(memory[869])
         );
  DFFRHQX1 memory_reg_9__4_ ( .D(n972), .CK(clk), .RN(rstn), .Q(memory[868])
         );
  DFFRHQX1 memory_reg_9__3_ ( .D(n971), .CK(clk), .RN(rstn), .Q(memory[867])
         );
  DFFRHQX1 memory_reg_9__2_ ( .D(n970), .CK(clk), .RN(rstn), .Q(memory[866])
         );
  DFFRHQX1 memory_reg_9__1_ ( .D(n969), .CK(clk), .RN(rstn), .Q(memory[865])
         );
  DFFRHQX1 memory_reg_9__0_ ( .D(n968), .CK(clk), .RN(rstn), .Q(memory[864])
         );
  DFFRHQX1 memory_reg_13__15_ ( .D(n919), .CK(clk), .RN(rstn), .Q(memory[815])
         );
  DFFRHQX1 memory_reg_13__14_ ( .D(n918), .CK(clk), .RN(rstn), .Q(memory[814])
         );
  DFFRHQX1 memory_reg_13__13_ ( .D(n917), .CK(clk), .RN(rstn), .Q(memory[813])
         );
  DFFRHQX1 memory_reg_13__12_ ( .D(n916), .CK(clk), .RN(rstn), .Q(memory[812])
         );
  DFFRHQX1 memory_reg_13__11_ ( .D(n915), .CK(clk), .RN(rstn), .Q(memory[811])
         );
  DFFRHQX1 memory_reg_13__10_ ( .D(n914), .CK(clk), .RN(rstn), .Q(memory[810])
         );
  DFFRHQX1 memory_reg_13__9_ ( .D(n913), .CK(clk), .RN(rstn), .Q(memory[809])
         );
  DFFRHQX1 memory_reg_13__8_ ( .D(n912), .CK(clk), .RN(rstn), .Q(memory[808])
         );
  DFFRHQX1 memory_reg_13__7_ ( .D(n911), .CK(clk), .RN(rstn), .Q(memory[807])
         );
  DFFRHQX1 memory_reg_13__6_ ( .D(n910), .CK(clk), .RN(rstn), .Q(memory[806])
         );
  DFFRHQX1 memory_reg_13__5_ ( .D(n909), .CK(clk), .RN(rstn), .Q(memory[805])
         );
  DFFRHQX1 memory_reg_13__4_ ( .D(n908), .CK(clk), .RN(rstn), .Q(memory[804])
         );
  DFFRHQX1 memory_reg_13__3_ ( .D(n907), .CK(clk), .RN(rstn), .Q(memory[803])
         );
  DFFRHQX1 memory_reg_13__2_ ( .D(n906), .CK(clk), .RN(rstn), .Q(memory[802])
         );
  DFFRHQX1 memory_reg_13__1_ ( .D(n905), .CK(clk), .RN(rstn), .Q(memory[801])
         );
  DFFRHQX1 memory_reg_13__0_ ( .D(n904), .CK(clk), .RN(rstn), .Q(memory[800])
         );
  DFFRHQX1 memory_reg_17__15_ ( .D(n855), .CK(clk), .RN(rstn), .Q(memory[751])
         );
  DFFRHQX1 memory_reg_17__14_ ( .D(n854), .CK(clk), .RN(rstn), .Q(memory[750])
         );
  DFFRHQX1 memory_reg_17__13_ ( .D(n853), .CK(clk), .RN(rstn), .Q(memory[749])
         );
  DFFRHQX1 memory_reg_17__12_ ( .D(n852), .CK(clk), .RN(rstn), .Q(memory[748])
         );
  DFFRHQX1 memory_reg_17__11_ ( .D(n851), .CK(clk), .RN(rstn), .Q(memory[747])
         );
  DFFRHQX1 memory_reg_17__10_ ( .D(n850), .CK(clk), .RN(rstn), .Q(memory[746])
         );
  DFFRHQX1 memory_reg_17__9_ ( .D(n849), .CK(clk), .RN(rstn), .Q(memory[745])
         );
  DFFRHQX1 memory_reg_17__8_ ( .D(n848), .CK(clk), .RN(rstn), .Q(memory[744])
         );
  DFFRHQX1 memory_reg_17__7_ ( .D(n847), .CK(clk), .RN(rstn), .Q(memory[743])
         );
  DFFRHQX1 memory_reg_17__6_ ( .D(n846), .CK(clk), .RN(rstn), .Q(memory[742])
         );
  DFFRHQX1 memory_reg_17__5_ ( .D(n845), .CK(clk), .RN(rstn), .Q(memory[741])
         );
  DFFRHQX1 memory_reg_17__4_ ( .D(n844), .CK(clk), .RN(rstn), .Q(memory[740])
         );
  DFFRHQX1 memory_reg_17__3_ ( .D(n843), .CK(clk), .RN(rstn), .Q(memory[739])
         );
  DFFRHQX1 memory_reg_17__2_ ( .D(n842), .CK(clk), .RN(rstn), .Q(memory[738])
         );
  DFFRHQX1 memory_reg_17__1_ ( .D(n841), .CK(clk), .RN(rstn), .Q(memory[737])
         );
  DFFRHQX1 memory_reg_17__0_ ( .D(n840), .CK(clk), .RN(rstn), .Q(memory[736])
         );
  DFFRHQX1 memory_reg_21__15_ ( .D(n791), .CK(clk), .RN(rstn), .Q(memory[687])
         );
  DFFRHQX1 memory_reg_21__14_ ( .D(n790), .CK(clk), .RN(rstn), .Q(memory[686])
         );
  DFFRHQX1 memory_reg_21__13_ ( .D(n789), .CK(clk), .RN(rstn), .Q(memory[685])
         );
  DFFRHQX1 memory_reg_21__12_ ( .D(n788), .CK(clk), .RN(rstn), .Q(memory[684])
         );
  DFFRHQX1 memory_reg_21__11_ ( .D(n787), .CK(clk), .RN(rstn), .Q(memory[683])
         );
  DFFRHQX1 memory_reg_21__10_ ( .D(n786), .CK(clk), .RN(rstn), .Q(memory[682])
         );
  DFFRHQX1 memory_reg_21__9_ ( .D(n785), .CK(clk), .RN(rstn), .Q(memory[681])
         );
  DFFRHQX1 memory_reg_21__8_ ( .D(n784), .CK(clk), .RN(rstn), .Q(memory[680])
         );
  DFFRHQX1 memory_reg_21__7_ ( .D(n783), .CK(clk), .RN(rstn), .Q(memory[679])
         );
  DFFRHQX1 memory_reg_21__6_ ( .D(n782), .CK(clk), .RN(rstn), .Q(memory[678])
         );
  DFFRHQX1 memory_reg_21__5_ ( .D(n781), .CK(clk), .RN(rstn), .Q(memory[677])
         );
  DFFRHQX1 memory_reg_21__4_ ( .D(n780), .CK(clk), .RN(rstn), .Q(memory[676])
         );
  DFFRHQX1 memory_reg_21__3_ ( .D(n779), .CK(clk), .RN(rstn), .Q(memory[675])
         );
  DFFRHQX1 memory_reg_21__2_ ( .D(n778), .CK(clk), .RN(rstn), .Q(memory[674])
         );
  DFFRHQX1 memory_reg_21__1_ ( .D(n777), .CK(clk), .RN(rstn), .Q(memory[673])
         );
  DFFRHQX1 memory_reg_21__0_ ( .D(n776), .CK(clk), .RN(rstn), .Q(memory[672])
         );
  DFFRHQX1 memory_reg_25__15_ ( .D(n727), .CK(clk), .RN(rstn), .Q(memory[623])
         );
  DFFRHQX1 memory_reg_25__14_ ( .D(n726), .CK(clk), .RN(rstn), .Q(memory[622])
         );
  DFFRHQX1 memory_reg_25__13_ ( .D(n725), .CK(clk), .RN(rstn), .Q(memory[621])
         );
  DFFRHQX1 memory_reg_25__12_ ( .D(n724), .CK(clk), .RN(rstn), .Q(memory[620])
         );
  DFFRHQX1 memory_reg_25__11_ ( .D(n723), .CK(clk), .RN(rstn), .Q(memory[619])
         );
  DFFRHQX1 memory_reg_25__10_ ( .D(n722), .CK(clk), .RN(rstn), .Q(memory[618])
         );
  DFFRHQX1 memory_reg_25__9_ ( .D(n721), .CK(clk), .RN(rstn), .Q(memory[617])
         );
  DFFRHQX1 memory_reg_25__8_ ( .D(n720), .CK(clk), .RN(rstn), .Q(memory[616])
         );
  DFFRHQX1 memory_reg_25__7_ ( .D(n719), .CK(clk), .RN(rstn), .Q(memory[615])
         );
  DFFRHQX1 memory_reg_25__6_ ( .D(n718), .CK(clk), .RN(rstn), .Q(memory[614])
         );
  DFFRHQX1 memory_reg_25__5_ ( .D(n717), .CK(clk), .RN(rstn), .Q(memory[613])
         );
  DFFRHQX1 memory_reg_25__4_ ( .D(n716), .CK(clk), .RN(rstn), .Q(memory[612])
         );
  DFFRHQX1 memory_reg_25__3_ ( .D(n715), .CK(clk), .RN(rstn), .Q(memory[611])
         );
  DFFRHQX1 memory_reg_25__2_ ( .D(n714), .CK(clk), .RN(rstn), .Q(memory[610])
         );
  DFFRHQX1 memory_reg_25__1_ ( .D(n713), .CK(clk), .RN(rstn), .Q(memory[609])
         );
  DFFRHQX1 memory_reg_25__0_ ( .D(n712), .CK(clk), .RN(rstn), .Q(memory[608])
         );
  DFFRHQX1 memory_reg_29__15_ ( .D(n663), .CK(clk), .RN(rstn), .Q(memory[559])
         );
  DFFRHQX1 memory_reg_29__14_ ( .D(n662), .CK(clk), .RN(rstn), .Q(memory[558])
         );
  DFFRHQX1 memory_reg_29__13_ ( .D(n661), .CK(clk), .RN(rstn), .Q(memory[557])
         );
  DFFRHQX1 memory_reg_29__12_ ( .D(n660), .CK(clk), .RN(rstn), .Q(memory[556])
         );
  DFFRHQX1 memory_reg_29__11_ ( .D(n659), .CK(clk), .RN(rstn), .Q(memory[555])
         );
  DFFRHQX1 memory_reg_29__10_ ( .D(n658), .CK(clk), .RN(rstn), .Q(memory[554])
         );
  DFFRHQX1 memory_reg_29__9_ ( .D(n657), .CK(clk), .RN(rstn), .Q(memory[553])
         );
  DFFRHQX1 memory_reg_29__8_ ( .D(n656), .CK(clk), .RN(rstn), .Q(memory[552])
         );
  DFFRHQX1 memory_reg_29__7_ ( .D(n655), .CK(clk), .RN(rstn), .Q(memory[551])
         );
  DFFRHQX1 memory_reg_29__6_ ( .D(n654), .CK(clk), .RN(rstn), .Q(memory[550])
         );
  DFFRHQX1 memory_reg_29__5_ ( .D(n653), .CK(clk), .RN(rstn), .Q(memory[549])
         );
  DFFRHQX1 memory_reg_29__4_ ( .D(n652), .CK(clk), .RN(rstn), .Q(memory[548])
         );
  DFFRHQX1 memory_reg_29__3_ ( .D(n651), .CK(clk), .RN(rstn), .Q(memory[547])
         );
  DFFRHQX1 memory_reg_29__2_ ( .D(n650), .CK(clk), .RN(rstn), .Q(memory[546])
         );
  DFFRHQX1 memory_reg_29__1_ ( .D(n649), .CK(clk), .RN(rstn), .Q(memory[545])
         );
  DFFRHQX1 memory_reg_29__0_ ( .D(n648), .CK(clk), .RN(rstn), .Q(memory[544])
         );
  DFFRHQX1 memory_reg_33__15_ ( .D(n599), .CK(clk), .RN(rstn), .Q(memory[495])
         );
  DFFRHQX1 memory_reg_33__14_ ( .D(n598), .CK(clk), .RN(rstn), .Q(memory[494])
         );
  DFFRHQX1 memory_reg_33__13_ ( .D(n597), .CK(clk), .RN(rstn), .Q(memory[493])
         );
  DFFRHQX1 memory_reg_33__12_ ( .D(n596), .CK(clk), .RN(rstn), .Q(memory[492])
         );
  DFFRHQX1 memory_reg_33__11_ ( .D(n595), .CK(clk), .RN(rstn), .Q(memory[491])
         );
  DFFRHQX1 memory_reg_33__10_ ( .D(n594), .CK(clk), .RN(rstn), .Q(memory[490])
         );
  DFFRHQX1 memory_reg_33__9_ ( .D(n593), .CK(clk), .RN(rstn), .Q(memory[489])
         );
  DFFRHQX1 memory_reg_33__8_ ( .D(n592), .CK(clk), .RN(rstn), .Q(memory[488])
         );
  DFFRHQX1 memory_reg_33__7_ ( .D(n591), .CK(clk), .RN(rstn), .Q(memory[487])
         );
  DFFRHQX1 memory_reg_33__6_ ( .D(n590), .CK(clk), .RN(rstn), .Q(memory[486])
         );
  DFFRHQX1 memory_reg_33__5_ ( .D(n589), .CK(clk), .RN(rstn), .Q(memory[485])
         );
  DFFRHQX1 memory_reg_33__4_ ( .D(n588), .CK(clk), .RN(rstn), .Q(memory[484])
         );
  DFFRHQX1 memory_reg_33__3_ ( .D(n587), .CK(clk), .RN(rstn), .Q(memory[483])
         );
  DFFRHQX1 memory_reg_33__2_ ( .D(n586), .CK(clk), .RN(rstn), .Q(memory[482])
         );
  DFFRHQX1 memory_reg_33__1_ ( .D(n585), .CK(clk), .RN(rstn), .Q(memory[481])
         );
  DFFRHQX1 memory_reg_33__0_ ( .D(n584), .CK(clk), .RN(rstn), .Q(memory[480])
         );
  DFFRHQX1 memory_reg_37__15_ ( .D(n535), .CK(clk), .RN(rstn), .Q(memory[431])
         );
  DFFRHQX1 memory_reg_37__14_ ( .D(n534), .CK(clk), .RN(rstn), .Q(memory[430])
         );
  DFFRHQX1 memory_reg_37__13_ ( .D(n533), .CK(clk), .RN(rstn), .Q(memory[429])
         );
  DFFRHQX1 memory_reg_37__12_ ( .D(n532), .CK(clk), .RN(rstn), .Q(memory[428])
         );
  DFFRHQX1 memory_reg_37__11_ ( .D(n531), .CK(clk), .RN(rstn), .Q(memory[427])
         );
  DFFRHQX1 memory_reg_37__10_ ( .D(n530), .CK(clk), .RN(rstn), .Q(memory[426])
         );
  DFFRHQX1 memory_reg_37__9_ ( .D(n529), .CK(clk), .RN(rstn), .Q(memory[425])
         );
  DFFRHQX1 memory_reg_37__8_ ( .D(n528), .CK(clk), .RN(rstn), .Q(memory[424])
         );
  DFFRHQX1 memory_reg_37__7_ ( .D(n527), .CK(clk), .RN(rstn), .Q(memory[423])
         );
  DFFRHQX1 memory_reg_37__6_ ( .D(n526), .CK(clk), .RN(rstn), .Q(memory[422])
         );
  DFFRHQX1 memory_reg_37__5_ ( .D(n525), .CK(clk), .RN(rstn), .Q(memory[421])
         );
  DFFRHQX1 memory_reg_37__4_ ( .D(n524), .CK(clk), .RN(rstn), .Q(memory[420])
         );
  DFFRHQX1 memory_reg_37__3_ ( .D(n523), .CK(clk), .RN(rstn), .Q(memory[419])
         );
  DFFRHQX1 memory_reg_37__2_ ( .D(n522), .CK(clk), .RN(rstn), .Q(memory[418])
         );
  DFFRHQX1 memory_reg_37__1_ ( .D(n521), .CK(clk), .RN(rstn), .Q(memory[417])
         );
  DFFRHQX1 memory_reg_37__0_ ( .D(n520), .CK(clk), .RN(rstn), .Q(memory[416])
         );
  DFFRHQX1 memory_reg_41__15_ ( .D(n471), .CK(clk), .RN(rstn), .Q(memory[367])
         );
  DFFRHQX1 memory_reg_41__14_ ( .D(n470), .CK(clk), .RN(rstn), .Q(memory[366])
         );
  DFFRHQX1 memory_reg_41__13_ ( .D(n469), .CK(clk), .RN(rstn), .Q(memory[365])
         );
  DFFRHQX1 memory_reg_41__12_ ( .D(n468), .CK(clk), .RN(rstn), .Q(memory[364])
         );
  DFFRHQX1 memory_reg_41__11_ ( .D(n467), .CK(clk), .RN(rstn), .Q(memory[363])
         );
  DFFRHQX1 memory_reg_41__10_ ( .D(n466), .CK(clk), .RN(rstn), .Q(memory[362])
         );
  DFFRHQX1 memory_reg_41__9_ ( .D(n465), .CK(clk), .RN(rstn), .Q(memory[361])
         );
  DFFRHQX1 memory_reg_41__8_ ( .D(n464), .CK(clk), .RN(rstn), .Q(memory[360])
         );
  DFFRHQX1 memory_reg_41__7_ ( .D(n463), .CK(clk), .RN(rstn), .Q(memory[359])
         );
  DFFRHQX1 memory_reg_41__6_ ( .D(n462), .CK(clk), .RN(rstn), .Q(memory[358])
         );
  DFFRHQX1 memory_reg_41__5_ ( .D(n461), .CK(clk), .RN(rstn), .Q(memory[357])
         );
  DFFRHQX1 memory_reg_41__4_ ( .D(n460), .CK(clk), .RN(rstn), .Q(memory[356])
         );
  DFFRHQX1 memory_reg_41__3_ ( .D(n459), .CK(clk), .RN(rstn), .Q(memory[355])
         );
  DFFRHQX1 memory_reg_41__2_ ( .D(n458), .CK(clk), .RN(rstn), .Q(memory[354])
         );
  DFFRHQX1 memory_reg_41__1_ ( .D(n457), .CK(clk), .RN(rstn), .Q(memory[353])
         );
  DFFRHQX1 memory_reg_41__0_ ( .D(n456), .CK(clk), .RN(rstn), .Q(memory[352])
         );
  DFFRHQX1 memory_reg_45__15_ ( .D(n407), .CK(clk), .RN(rstn), .Q(memory[303])
         );
  DFFRHQX1 memory_reg_45__14_ ( .D(n406), .CK(clk), .RN(rstn), .Q(memory[302])
         );
  DFFRHQX1 memory_reg_45__13_ ( .D(n405), .CK(clk), .RN(rstn), .Q(memory[301])
         );
  DFFRHQX1 memory_reg_45__12_ ( .D(n404), .CK(clk), .RN(rstn), .Q(memory[300])
         );
  DFFRHQX1 memory_reg_45__11_ ( .D(n403), .CK(clk), .RN(rstn), .Q(memory[299])
         );
  DFFRHQX1 memory_reg_45__10_ ( .D(n402), .CK(clk), .RN(rstn), .Q(memory[298])
         );
  DFFRHQX1 memory_reg_45__9_ ( .D(n401), .CK(clk), .RN(rstn), .Q(memory[297])
         );
  DFFRHQX1 memory_reg_45__8_ ( .D(n400), .CK(clk), .RN(rstn), .Q(memory[296])
         );
  DFFRHQX1 memory_reg_45__7_ ( .D(n399), .CK(clk), .RN(rstn), .Q(memory[295])
         );
  DFFRHQX1 memory_reg_45__6_ ( .D(n398), .CK(clk), .RN(rstn), .Q(memory[294])
         );
  DFFRHQX1 memory_reg_45__5_ ( .D(n397), .CK(clk), .RN(rstn), .Q(memory[293])
         );
  DFFRHQX1 memory_reg_45__4_ ( .D(n396), .CK(clk), .RN(rstn), .Q(memory[292])
         );
  DFFRHQX1 memory_reg_45__3_ ( .D(n395), .CK(clk), .RN(rstn), .Q(memory[291])
         );
  DFFRHQX1 memory_reg_45__2_ ( .D(n394), .CK(clk), .RN(rstn), .Q(memory[290])
         );
  DFFRHQX1 memory_reg_45__1_ ( .D(n393), .CK(clk), .RN(rstn), .Q(memory[289])
         );
  DFFRHQX1 memory_reg_45__0_ ( .D(n392), .CK(clk), .RN(rstn), .Q(memory[288])
         );
  DFFRHQX1 memory_reg_49__15_ ( .D(n343), .CK(clk), .RN(rstn), .Q(memory[239])
         );
  DFFRHQX1 memory_reg_49__14_ ( .D(n342), .CK(clk), .RN(rstn), .Q(memory[238])
         );
  DFFRHQX1 memory_reg_49__13_ ( .D(n341), .CK(clk), .RN(rstn), .Q(memory[237])
         );
  DFFRHQX1 memory_reg_49__12_ ( .D(n340), .CK(clk), .RN(rstn), .Q(memory[236])
         );
  DFFRHQX1 memory_reg_49__11_ ( .D(n339), .CK(clk), .RN(rstn), .Q(memory[235])
         );
  DFFRHQX1 memory_reg_49__10_ ( .D(n338), .CK(clk), .RN(rstn), .Q(memory[234])
         );
  DFFRHQX1 memory_reg_49__9_ ( .D(n337), .CK(clk), .RN(rstn), .Q(memory[233])
         );
  DFFRHQX1 memory_reg_49__8_ ( .D(n336), .CK(clk), .RN(rstn), .Q(memory[232])
         );
  DFFRHQX1 memory_reg_49__7_ ( .D(n335), .CK(clk), .RN(rstn), .Q(memory[231])
         );
  DFFRHQX1 memory_reg_49__6_ ( .D(n334), .CK(clk), .RN(rstn), .Q(memory[230])
         );
  DFFRHQX1 memory_reg_49__5_ ( .D(n333), .CK(clk), .RN(rstn), .Q(memory[229])
         );
  DFFRHQX1 memory_reg_49__4_ ( .D(n332), .CK(clk), .RN(rstn), .Q(memory[228])
         );
  DFFRHQX1 memory_reg_49__3_ ( .D(n331), .CK(clk), .RN(rstn), .Q(memory[227])
         );
  DFFRHQX1 memory_reg_49__2_ ( .D(n330), .CK(clk), .RN(rstn), .Q(memory[226])
         );
  DFFRHQX1 memory_reg_49__1_ ( .D(n329), .CK(clk), .RN(rstn), .Q(memory[225])
         );
  DFFRHQX1 memory_reg_49__0_ ( .D(n328), .CK(clk), .RN(rstn), .Q(memory[224])
         );
  DFFRHQX1 memory_reg_53__15_ ( .D(n279), .CK(clk), .RN(rstn), .Q(memory[175])
         );
  DFFRHQX1 memory_reg_53__14_ ( .D(n278), .CK(clk), .RN(rstn), .Q(memory[174])
         );
  DFFRHQX1 memory_reg_53__13_ ( .D(n277), .CK(clk), .RN(rstn), .Q(memory[173])
         );
  DFFRHQX1 memory_reg_53__12_ ( .D(n276), .CK(clk), .RN(rstn), .Q(memory[172])
         );
  DFFRHQX1 memory_reg_53__11_ ( .D(n275), .CK(clk), .RN(rstn), .Q(memory[171])
         );
  DFFRHQX1 memory_reg_53__10_ ( .D(n274), .CK(clk), .RN(rstn), .Q(memory[170])
         );
  DFFRHQX1 memory_reg_53__9_ ( .D(n273), .CK(clk), .RN(rstn), .Q(memory[169])
         );
  DFFRHQX1 memory_reg_53__8_ ( .D(n272), .CK(clk), .RN(rstn), .Q(memory[168])
         );
  DFFRHQX1 memory_reg_53__7_ ( .D(n271), .CK(clk), .RN(rstn), .Q(memory[167])
         );
  DFFRHQX1 memory_reg_53__6_ ( .D(n270), .CK(clk), .RN(rstn), .Q(memory[166])
         );
  DFFRHQX1 memory_reg_53__5_ ( .D(n269), .CK(clk), .RN(rstn), .Q(memory[165])
         );
  DFFRHQX1 memory_reg_53__4_ ( .D(n268), .CK(clk), .RN(rstn), .Q(memory[164])
         );
  DFFRHQX1 memory_reg_53__3_ ( .D(n267), .CK(clk), .RN(rstn), .Q(memory[163])
         );
  DFFRHQX1 memory_reg_53__2_ ( .D(n266), .CK(clk), .RN(rstn), .Q(memory[162])
         );
  DFFRHQX1 memory_reg_53__1_ ( .D(n265), .CK(clk), .RN(rstn), .Q(memory[161])
         );
  DFFRHQX1 memory_reg_53__0_ ( .D(n264), .CK(clk), .RN(rstn), .Q(memory[160])
         );
  DFFRHQX1 memory_reg_57__15_ ( .D(n215), .CK(clk), .RN(rstn), .Q(memory[111])
         );
  DFFRHQX1 memory_reg_57__14_ ( .D(n214), .CK(clk), .RN(rstn), .Q(memory[110])
         );
  DFFRHQX1 memory_reg_57__13_ ( .D(n213), .CK(clk), .RN(rstn), .Q(memory[109])
         );
  DFFRHQX1 memory_reg_57__12_ ( .D(n212), .CK(clk), .RN(rstn), .Q(memory[108])
         );
  DFFRHQX1 memory_reg_57__11_ ( .D(n211), .CK(clk), .RN(rstn), .Q(memory[107])
         );
  DFFRHQX1 memory_reg_57__10_ ( .D(n210), .CK(clk), .RN(rstn), .Q(memory[106])
         );
  DFFRHQX1 memory_reg_57__9_ ( .D(n209), .CK(clk), .RN(rstn), .Q(memory[105])
         );
  DFFRHQX1 memory_reg_57__8_ ( .D(n208), .CK(clk), .RN(rstn), .Q(memory[104])
         );
  DFFRHQX1 memory_reg_57__7_ ( .D(n207), .CK(clk), .RN(rstn), .Q(memory[103])
         );
  DFFRHQX1 memory_reg_57__6_ ( .D(n206), .CK(clk), .RN(rstn), .Q(memory[102])
         );
  DFFRHQX1 memory_reg_57__5_ ( .D(n205), .CK(clk), .RN(rstn), .Q(memory[101])
         );
  DFFRHQX1 memory_reg_57__4_ ( .D(n204), .CK(clk), .RN(rstn), .Q(memory[100])
         );
  DFFRHQX1 memory_reg_57__3_ ( .D(n203), .CK(clk), .RN(rstn), .Q(memory[99])
         );
  DFFRHQX1 memory_reg_57__2_ ( .D(n202), .CK(clk), .RN(rstn), .Q(memory[98])
         );
  DFFRHQX1 memory_reg_57__1_ ( .D(n201), .CK(clk), .RN(rstn), .Q(memory[97])
         );
  DFFRHQX1 memory_reg_57__0_ ( .D(n200), .CK(clk), .RN(rstn), .Q(memory[96])
         );
  DFFRHQX1 memory_reg_61__15_ ( .D(n151), .CK(clk), .RN(rstn), .Q(memory[47])
         );
  DFFRHQX1 memory_reg_61__14_ ( .D(n150), .CK(clk), .RN(rstn), .Q(memory[46])
         );
  DFFRHQX1 memory_reg_61__13_ ( .D(n149), .CK(clk), .RN(rstn), .Q(memory[45])
         );
  DFFRHQX1 memory_reg_61__12_ ( .D(n148), .CK(clk), .RN(rstn), .Q(memory[44])
         );
  DFFRHQX1 memory_reg_61__11_ ( .D(n147), .CK(clk), .RN(rstn), .Q(memory[43])
         );
  DFFRHQX1 memory_reg_61__10_ ( .D(n146), .CK(clk), .RN(rstn), .Q(memory[42])
         );
  DFFRHQX1 memory_reg_61__9_ ( .D(n145), .CK(clk), .RN(rstn), .Q(memory[41])
         );
  DFFRHQX1 memory_reg_61__8_ ( .D(n144), .CK(clk), .RN(rstn), .Q(memory[40])
         );
  DFFRHQX1 memory_reg_61__7_ ( .D(n143), .CK(clk), .RN(rstn), .Q(memory[39])
         );
  DFFRHQX1 memory_reg_61__6_ ( .D(n142), .CK(clk), .RN(rstn), .Q(memory[38])
         );
  DFFRHQX1 memory_reg_61__5_ ( .D(n141), .CK(clk), .RN(rstn), .Q(memory[37])
         );
  DFFRHQX1 memory_reg_61__4_ ( .D(n140), .CK(clk), .RN(rstn), .Q(memory[36])
         );
  DFFRHQX1 memory_reg_61__3_ ( .D(n139), .CK(clk), .RN(rstn), .Q(memory[35])
         );
  DFFRHQX1 memory_reg_61__2_ ( .D(n138), .CK(clk), .RN(rstn), .Q(memory[34])
         );
  DFFRHQX1 memory_reg_61__1_ ( .D(n137), .CK(clk), .RN(rstn), .Q(memory[33])
         );
  DFFRHQX1 memory_reg_61__0_ ( .D(n136), .CK(clk), .RN(rstn), .Q(memory[32])
         );
  DFFRHQX1 memory_reg_3__15_ ( .D(n1079), .CK(clk), .RN(rstn), .Q(memory[975])
         );
  DFFRHQX1 memory_reg_3__14_ ( .D(n1078), .CK(clk), .RN(rstn), .Q(memory[974])
         );
  DFFRHQX1 memory_reg_3__13_ ( .D(n1077), .CK(clk), .RN(rstn), .Q(memory[973])
         );
  DFFRHQX1 memory_reg_3__12_ ( .D(n1076), .CK(clk), .RN(rstn), .Q(memory[972])
         );
  DFFRHQX1 memory_reg_3__11_ ( .D(n1075), .CK(clk), .RN(rstn), .Q(memory[971])
         );
  DFFRHQX1 memory_reg_3__10_ ( .D(n1074), .CK(clk), .RN(rstn), .Q(memory[970])
         );
  DFFRHQX1 memory_reg_3__9_ ( .D(n1073), .CK(clk), .RN(rstn), .Q(memory[969])
         );
  DFFRHQX1 memory_reg_3__8_ ( .D(n1072), .CK(clk), .RN(rstn), .Q(memory[968])
         );
  DFFRHQX1 memory_reg_3__7_ ( .D(n1071), .CK(clk), .RN(rstn), .Q(memory[967])
         );
  DFFRHQX1 memory_reg_3__6_ ( .D(n1070), .CK(clk), .RN(rstn), .Q(memory[966])
         );
  DFFRHQX1 memory_reg_3__5_ ( .D(n1069), .CK(clk), .RN(rstn), .Q(memory[965])
         );
  DFFRHQX1 memory_reg_3__4_ ( .D(n1068), .CK(clk), .RN(rstn), .Q(memory[964])
         );
  DFFRHQX1 memory_reg_3__3_ ( .D(n1067), .CK(clk), .RN(rstn), .Q(memory[963])
         );
  DFFRHQX1 memory_reg_3__2_ ( .D(n1066), .CK(clk), .RN(rstn), .Q(memory[962])
         );
  DFFRHQX1 memory_reg_3__1_ ( .D(n1065), .CK(clk), .RN(rstn), .Q(memory[961])
         );
  DFFRHQX1 memory_reg_3__0_ ( .D(n1064), .CK(clk), .RN(rstn), .Q(memory[960])
         );
  DFFRHQX1 memory_reg_7__15_ ( .D(n1015), .CK(clk), .RN(rstn), .Q(memory[911])
         );
  DFFRHQX1 memory_reg_7__14_ ( .D(n1014), .CK(clk), .RN(rstn), .Q(memory[910])
         );
  DFFRHQX1 memory_reg_7__13_ ( .D(n1013), .CK(clk), .RN(rstn), .Q(memory[909])
         );
  DFFRHQX1 memory_reg_7__12_ ( .D(n1012), .CK(clk), .RN(rstn), .Q(memory[908])
         );
  DFFRHQX1 memory_reg_7__11_ ( .D(n1011), .CK(clk), .RN(rstn), .Q(memory[907])
         );
  DFFRHQX1 memory_reg_7__10_ ( .D(n1010), .CK(clk), .RN(rstn), .Q(memory[906])
         );
  DFFRHQX1 memory_reg_7__9_ ( .D(n1009), .CK(clk), .RN(rstn), .Q(memory[905])
         );
  DFFRHQX1 memory_reg_7__8_ ( .D(n1008), .CK(clk), .RN(rstn), .Q(memory[904])
         );
  DFFRHQX1 memory_reg_7__7_ ( .D(n1007), .CK(clk), .RN(rstn), .Q(memory[903])
         );
  DFFRHQX1 memory_reg_7__6_ ( .D(n1006), .CK(clk), .RN(rstn), .Q(memory[902])
         );
  DFFRHQX1 memory_reg_7__5_ ( .D(n1005), .CK(clk), .RN(rstn), .Q(memory[901])
         );
  DFFRHQX1 memory_reg_7__4_ ( .D(n1004), .CK(clk), .RN(rstn), .Q(memory[900])
         );
  DFFRHQX1 memory_reg_7__3_ ( .D(n1003), .CK(clk), .RN(rstn), .Q(memory[899])
         );
  DFFRHQX1 memory_reg_7__2_ ( .D(n1002), .CK(clk), .RN(rstn), .Q(memory[898])
         );
  DFFRHQX1 memory_reg_7__1_ ( .D(n1001), .CK(clk), .RN(rstn), .Q(memory[897])
         );
  DFFRHQX1 memory_reg_7__0_ ( .D(n1000), .CK(clk), .RN(rstn), .Q(memory[896])
         );
  DFFRHQX1 memory_reg_11__15_ ( .D(n951), .CK(clk), .RN(rstn), .Q(memory[847])
         );
  DFFRHQX1 memory_reg_11__14_ ( .D(n950), .CK(clk), .RN(rstn), .Q(memory[846])
         );
  DFFRHQX1 memory_reg_11__13_ ( .D(n949), .CK(clk), .RN(rstn), .Q(memory[845])
         );
  DFFRHQX1 memory_reg_11__12_ ( .D(n948), .CK(clk), .RN(rstn), .Q(memory[844])
         );
  DFFRHQX1 memory_reg_11__11_ ( .D(n947), .CK(clk), .RN(rstn), .Q(memory[843])
         );
  DFFRHQX1 memory_reg_11__10_ ( .D(n946), .CK(clk), .RN(rstn), .Q(memory[842])
         );
  DFFRHQX1 memory_reg_11__9_ ( .D(n945), .CK(clk), .RN(rstn), .Q(memory[841])
         );
  DFFRHQX1 memory_reg_11__8_ ( .D(n944), .CK(clk), .RN(rstn), .Q(memory[840])
         );
  DFFRHQX1 memory_reg_11__7_ ( .D(n943), .CK(clk), .RN(rstn), .Q(memory[839])
         );
  DFFRHQX1 memory_reg_11__6_ ( .D(n942), .CK(clk), .RN(rstn), .Q(memory[838])
         );
  DFFRHQX1 memory_reg_11__5_ ( .D(n941), .CK(clk), .RN(rstn), .Q(memory[837])
         );
  DFFRHQX1 memory_reg_11__4_ ( .D(n940), .CK(clk), .RN(rstn), .Q(memory[836])
         );
  DFFRHQX1 memory_reg_11__3_ ( .D(n939), .CK(clk), .RN(rstn), .Q(memory[835])
         );
  DFFRHQX1 memory_reg_11__2_ ( .D(n938), .CK(clk), .RN(rstn), .Q(memory[834])
         );
  DFFRHQX1 memory_reg_11__1_ ( .D(n937), .CK(clk), .RN(rstn), .Q(memory[833])
         );
  DFFRHQX1 memory_reg_11__0_ ( .D(n936), .CK(clk), .RN(rstn), .Q(memory[832])
         );
  DFFRHQX1 memory_reg_15__15_ ( .D(n887), .CK(clk), .RN(rstn), .Q(memory[783])
         );
  DFFRHQX1 memory_reg_15__14_ ( .D(n886), .CK(clk), .RN(rstn), .Q(memory[782])
         );
  DFFRHQX1 memory_reg_15__13_ ( .D(n885), .CK(clk), .RN(rstn), .Q(memory[781])
         );
  DFFRHQX1 memory_reg_15__12_ ( .D(n884), .CK(clk), .RN(rstn), .Q(memory[780])
         );
  DFFRHQX1 memory_reg_15__11_ ( .D(n883), .CK(clk), .RN(rstn), .Q(memory[779])
         );
  DFFRHQX1 memory_reg_15__10_ ( .D(n882), .CK(clk), .RN(rstn), .Q(memory[778])
         );
  DFFRHQX1 memory_reg_15__9_ ( .D(n881), .CK(clk), .RN(rstn), .Q(memory[777])
         );
  DFFRHQX1 memory_reg_15__8_ ( .D(n880), .CK(clk), .RN(rstn), .Q(memory[776])
         );
  DFFRHQX1 memory_reg_15__7_ ( .D(n879), .CK(clk), .RN(rstn), .Q(memory[775])
         );
  DFFRHQX1 memory_reg_15__6_ ( .D(n878), .CK(clk), .RN(rstn), .Q(memory[774])
         );
  DFFRHQX1 memory_reg_15__5_ ( .D(n877), .CK(clk), .RN(rstn), .Q(memory[773])
         );
  DFFRHQX1 memory_reg_15__4_ ( .D(n876), .CK(clk), .RN(rstn), .Q(memory[772])
         );
  DFFRHQX1 memory_reg_15__3_ ( .D(n875), .CK(clk), .RN(rstn), .Q(memory[771])
         );
  DFFRHQX1 memory_reg_15__2_ ( .D(n874), .CK(clk), .RN(rstn), .Q(memory[770])
         );
  DFFRHQX1 memory_reg_15__1_ ( .D(n873), .CK(clk), .RN(rstn), .Q(memory[769])
         );
  DFFRHQX1 memory_reg_15__0_ ( .D(n872), .CK(clk), .RN(rstn), .Q(memory[768])
         );
  DFFRHQX1 memory_reg_19__15_ ( .D(n823), .CK(clk), .RN(rstn), .Q(memory[719])
         );
  DFFRHQX1 memory_reg_19__14_ ( .D(n822), .CK(clk), .RN(rstn), .Q(memory[718])
         );
  DFFRHQX1 memory_reg_19__13_ ( .D(n821), .CK(clk), .RN(rstn), .Q(memory[717])
         );
  DFFRHQX1 memory_reg_19__12_ ( .D(n820), .CK(clk), .RN(rstn), .Q(memory[716])
         );
  DFFRHQX1 memory_reg_19__11_ ( .D(n819), .CK(clk), .RN(rstn), .Q(memory[715])
         );
  DFFRHQX1 memory_reg_19__10_ ( .D(n818), .CK(clk), .RN(rstn), .Q(memory[714])
         );
  DFFRHQX1 memory_reg_19__9_ ( .D(n817), .CK(clk), .RN(rstn), .Q(memory[713])
         );
  DFFRHQX1 memory_reg_19__8_ ( .D(n816), .CK(clk), .RN(rstn), .Q(memory[712])
         );
  DFFRHQX1 memory_reg_19__7_ ( .D(n815), .CK(clk), .RN(rstn), .Q(memory[711])
         );
  DFFRHQX1 memory_reg_19__6_ ( .D(n814), .CK(clk), .RN(rstn), .Q(memory[710])
         );
  DFFRHQX1 memory_reg_19__5_ ( .D(n813), .CK(clk), .RN(rstn), .Q(memory[709])
         );
  DFFRHQX1 memory_reg_19__4_ ( .D(n812), .CK(clk), .RN(rstn), .Q(memory[708])
         );
  DFFRHQX1 memory_reg_19__3_ ( .D(n811), .CK(clk), .RN(rstn), .Q(memory[707])
         );
  DFFRHQX1 memory_reg_19__2_ ( .D(n810), .CK(clk), .RN(rstn), .Q(memory[706])
         );
  DFFRHQX1 memory_reg_19__1_ ( .D(n809), .CK(clk), .RN(rstn), .Q(memory[705])
         );
  DFFRHQX1 memory_reg_19__0_ ( .D(n808), .CK(clk), .RN(rstn), .Q(memory[704])
         );
  DFFRHQX1 memory_reg_23__15_ ( .D(n759), .CK(clk), .RN(rstn), .Q(memory[655])
         );
  DFFRHQX1 memory_reg_23__14_ ( .D(n758), .CK(clk), .RN(rstn), .Q(memory[654])
         );
  DFFRHQX1 memory_reg_23__13_ ( .D(n757), .CK(clk), .RN(rstn), .Q(memory[653])
         );
  DFFRHQX1 memory_reg_23__12_ ( .D(n756), .CK(clk), .RN(rstn), .Q(memory[652])
         );
  DFFRHQX1 memory_reg_23__11_ ( .D(n755), .CK(clk), .RN(rstn), .Q(memory[651])
         );
  DFFRHQX1 memory_reg_23__10_ ( .D(n754), .CK(clk), .RN(rstn), .Q(memory[650])
         );
  DFFRHQX1 memory_reg_23__9_ ( .D(n753), .CK(clk), .RN(rstn), .Q(memory[649])
         );
  DFFRHQX1 memory_reg_23__8_ ( .D(n752), .CK(clk), .RN(rstn), .Q(memory[648])
         );
  DFFRHQX1 memory_reg_23__7_ ( .D(n751), .CK(clk), .RN(rstn), .Q(memory[647])
         );
  DFFRHQX1 memory_reg_23__6_ ( .D(n750), .CK(clk), .RN(rstn), .Q(memory[646])
         );
  DFFRHQX1 memory_reg_23__5_ ( .D(n749), .CK(clk), .RN(rstn), .Q(memory[645])
         );
  DFFRHQX1 memory_reg_23__4_ ( .D(n748), .CK(clk), .RN(rstn), .Q(memory[644])
         );
  DFFRHQX1 memory_reg_23__3_ ( .D(n747), .CK(clk), .RN(rstn), .Q(memory[643])
         );
  DFFRHQX1 memory_reg_23__2_ ( .D(n746), .CK(clk), .RN(rstn), .Q(memory[642])
         );
  DFFRHQX1 memory_reg_23__1_ ( .D(n745), .CK(clk), .RN(rstn), .Q(memory[641])
         );
  DFFRHQX1 memory_reg_23__0_ ( .D(n744), .CK(clk), .RN(rstn), .Q(memory[640])
         );
  DFFRHQX1 memory_reg_27__15_ ( .D(n695), .CK(clk), .RN(rstn), .Q(memory[591])
         );
  DFFRHQX1 memory_reg_27__14_ ( .D(n694), .CK(clk), .RN(rstn), .Q(memory[590])
         );
  DFFRHQX1 memory_reg_27__13_ ( .D(n693), .CK(clk), .RN(rstn), .Q(memory[589])
         );
  DFFRHQX1 memory_reg_27__12_ ( .D(n692), .CK(clk), .RN(rstn), .Q(memory[588])
         );
  DFFRHQX1 memory_reg_27__11_ ( .D(n691), .CK(clk), .RN(rstn), .Q(memory[587])
         );
  DFFRHQX1 memory_reg_27__10_ ( .D(n690), .CK(clk), .RN(rstn), .Q(memory[586])
         );
  DFFRHQX1 memory_reg_27__9_ ( .D(n689), .CK(clk), .RN(rstn), .Q(memory[585])
         );
  DFFRHQX1 memory_reg_27__8_ ( .D(n688), .CK(clk), .RN(rstn), .Q(memory[584])
         );
  DFFRHQX1 memory_reg_27__7_ ( .D(n687), .CK(clk), .RN(rstn), .Q(memory[583])
         );
  DFFRHQX1 memory_reg_27__6_ ( .D(n686), .CK(clk), .RN(rstn), .Q(memory[582])
         );
  DFFRHQX1 memory_reg_27__5_ ( .D(n685), .CK(clk), .RN(rstn), .Q(memory[581])
         );
  DFFRHQX1 memory_reg_27__4_ ( .D(n684), .CK(clk), .RN(rstn), .Q(memory[580])
         );
  DFFRHQX1 memory_reg_27__3_ ( .D(n683), .CK(clk), .RN(rstn), .Q(memory[579])
         );
  DFFRHQX1 memory_reg_27__2_ ( .D(n682), .CK(clk), .RN(rstn), .Q(memory[578])
         );
  DFFRHQX1 memory_reg_27__1_ ( .D(n681), .CK(clk), .RN(rstn), .Q(memory[577])
         );
  DFFRHQX1 memory_reg_27__0_ ( .D(n680), .CK(clk), .RN(rstn), .Q(memory[576])
         );
  DFFRHQX1 memory_reg_31__15_ ( .D(n631), .CK(clk), .RN(rstn), .Q(memory[527])
         );
  DFFRHQX1 memory_reg_31__14_ ( .D(n630), .CK(clk), .RN(rstn), .Q(memory[526])
         );
  DFFRHQX1 memory_reg_31__13_ ( .D(n629), .CK(clk), .RN(rstn), .Q(memory[525])
         );
  DFFRHQX1 memory_reg_31__12_ ( .D(n628), .CK(clk), .RN(rstn), .Q(memory[524])
         );
  DFFRHQX1 memory_reg_31__11_ ( .D(n627), .CK(clk), .RN(rstn), .Q(memory[523])
         );
  DFFRHQX1 memory_reg_31__10_ ( .D(n626), .CK(clk), .RN(rstn), .Q(memory[522])
         );
  DFFRHQX1 memory_reg_31__9_ ( .D(n625), .CK(clk), .RN(rstn), .Q(memory[521])
         );
  DFFRHQX1 memory_reg_31__8_ ( .D(n624), .CK(clk), .RN(rstn), .Q(memory[520])
         );
  DFFRHQX1 memory_reg_31__7_ ( .D(n623), .CK(clk), .RN(rstn), .Q(memory[519])
         );
  DFFRHQX1 memory_reg_31__6_ ( .D(n622), .CK(clk), .RN(rstn), .Q(memory[518])
         );
  DFFRHQX1 memory_reg_31__5_ ( .D(n621), .CK(clk), .RN(rstn), .Q(memory[517])
         );
  DFFRHQX1 memory_reg_31__4_ ( .D(n620), .CK(clk), .RN(rstn), .Q(memory[516])
         );
  DFFRHQX1 memory_reg_31__3_ ( .D(n619), .CK(clk), .RN(rstn), .Q(memory[515])
         );
  DFFRHQX1 memory_reg_31__2_ ( .D(n618), .CK(clk), .RN(rstn), .Q(memory[514])
         );
  DFFRHQX1 memory_reg_31__1_ ( .D(n617), .CK(clk), .RN(rstn), .Q(memory[513])
         );
  DFFRHQX1 memory_reg_31__0_ ( .D(n616), .CK(clk), .RN(rstn), .Q(memory[512])
         );
  DFFRHQX1 memory_reg_35__15_ ( .D(n567), .CK(clk), .RN(rstn), .Q(memory[463])
         );
  DFFRHQX1 memory_reg_35__14_ ( .D(n566), .CK(clk), .RN(rstn), .Q(memory[462])
         );
  DFFRHQX1 memory_reg_35__13_ ( .D(n565), .CK(clk), .RN(rstn), .Q(memory[461])
         );
  DFFRHQX1 memory_reg_35__12_ ( .D(n564), .CK(clk), .RN(rstn), .Q(memory[460])
         );
  DFFRHQX1 memory_reg_35__11_ ( .D(n563), .CK(clk), .RN(rstn), .Q(memory[459])
         );
  DFFRHQX1 memory_reg_35__10_ ( .D(n562), .CK(clk), .RN(rstn), .Q(memory[458])
         );
  DFFRHQX1 memory_reg_35__9_ ( .D(n561), .CK(clk), .RN(rstn), .Q(memory[457])
         );
  DFFRHQX1 memory_reg_35__8_ ( .D(n560), .CK(clk), .RN(rstn), .Q(memory[456])
         );
  DFFRHQX1 memory_reg_35__7_ ( .D(n559), .CK(clk), .RN(rstn), .Q(memory[455])
         );
  DFFRHQX1 memory_reg_35__6_ ( .D(n558), .CK(clk), .RN(rstn), .Q(memory[454])
         );
  DFFRHQX1 memory_reg_35__5_ ( .D(n557), .CK(clk), .RN(rstn), .Q(memory[453])
         );
  DFFRHQX1 memory_reg_35__4_ ( .D(n556), .CK(clk), .RN(rstn), .Q(memory[452])
         );
  DFFRHQX1 memory_reg_35__3_ ( .D(n555), .CK(clk), .RN(rstn), .Q(memory[451])
         );
  DFFRHQX1 memory_reg_35__2_ ( .D(n554), .CK(clk), .RN(rstn), .Q(memory[450])
         );
  DFFRHQX1 memory_reg_35__1_ ( .D(n553), .CK(clk), .RN(rstn), .Q(memory[449])
         );
  DFFRHQX1 memory_reg_35__0_ ( .D(n552), .CK(clk), .RN(rstn), .Q(memory[448])
         );
  DFFRHQX1 memory_reg_39__15_ ( .D(n503), .CK(clk), .RN(rstn), .Q(memory[399])
         );
  DFFRHQX1 memory_reg_39__14_ ( .D(n502), .CK(clk), .RN(rstn), .Q(memory[398])
         );
  DFFRHQX1 memory_reg_39__13_ ( .D(n501), .CK(clk), .RN(rstn), .Q(memory[397])
         );
  DFFRHQX1 memory_reg_39__12_ ( .D(n500), .CK(clk), .RN(rstn), .Q(memory[396])
         );
  DFFRHQX1 memory_reg_39__11_ ( .D(n499), .CK(clk), .RN(rstn), .Q(memory[395])
         );
  DFFRHQX1 memory_reg_39__10_ ( .D(n498), .CK(clk), .RN(rstn), .Q(memory[394])
         );
  DFFRHQX1 memory_reg_39__9_ ( .D(n497), .CK(clk), .RN(rstn), .Q(memory[393])
         );
  DFFRHQX1 memory_reg_39__8_ ( .D(n496), .CK(clk), .RN(rstn), .Q(memory[392])
         );
  DFFRHQX1 memory_reg_39__7_ ( .D(n495), .CK(clk), .RN(rstn), .Q(memory[391])
         );
  DFFRHQX1 memory_reg_39__6_ ( .D(n494), .CK(clk), .RN(rstn), .Q(memory[390])
         );
  DFFRHQX1 memory_reg_39__5_ ( .D(n493), .CK(clk), .RN(rstn), .Q(memory[389])
         );
  DFFRHQX1 memory_reg_39__4_ ( .D(n492), .CK(clk), .RN(rstn), .Q(memory[388])
         );
  DFFRHQX1 memory_reg_39__3_ ( .D(n491), .CK(clk), .RN(rstn), .Q(memory[387])
         );
  DFFRHQX1 memory_reg_39__2_ ( .D(n490), .CK(clk), .RN(rstn), .Q(memory[386])
         );
  DFFRHQX1 memory_reg_39__1_ ( .D(n489), .CK(clk), .RN(rstn), .Q(memory[385])
         );
  DFFRHQX1 memory_reg_39__0_ ( .D(n488), .CK(clk), .RN(rstn), .Q(memory[384])
         );
  DFFRHQX1 memory_reg_43__15_ ( .D(n439), .CK(clk), .RN(rstn), .Q(memory[335])
         );
  DFFRHQX1 memory_reg_43__14_ ( .D(n438), .CK(clk), .RN(rstn), .Q(memory[334])
         );
  DFFRHQX1 memory_reg_43__13_ ( .D(n437), .CK(clk), .RN(rstn), .Q(memory[333])
         );
  DFFRHQX1 memory_reg_43__12_ ( .D(n436), .CK(clk), .RN(rstn), .Q(memory[332])
         );
  DFFRHQX1 memory_reg_43__11_ ( .D(n435), .CK(clk), .RN(rstn), .Q(memory[331])
         );
  DFFRHQX1 memory_reg_43__10_ ( .D(n434), .CK(clk), .RN(rstn), .Q(memory[330])
         );
  DFFRHQX1 memory_reg_43__9_ ( .D(n433), .CK(clk), .RN(rstn), .Q(memory[329])
         );
  DFFRHQX1 memory_reg_43__8_ ( .D(n432), .CK(clk), .RN(rstn), .Q(memory[328])
         );
  DFFRHQX1 memory_reg_43__7_ ( .D(n431), .CK(clk), .RN(rstn), .Q(memory[327])
         );
  DFFRHQX1 memory_reg_43__6_ ( .D(n430), .CK(clk), .RN(rstn), .Q(memory[326])
         );
  DFFRHQX1 memory_reg_43__5_ ( .D(n429), .CK(clk), .RN(rstn), .Q(memory[325])
         );
  DFFRHQX1 memory_reg_43__4_ ( .D(n428), .CK(clk), .RN(rstn), .Q(memory[324])
         );
  DFFRHQX1 memory_reg_43__3_ ( .D(n427), .CK(clk), .RN(rstn), .Q(memory[323])
         );
  DFFRHQX1 memory_reg_43__2_ ( .D(n426), .CK(clk), .RN(rstn), .Q(memory[322])
         );
  DFFRHQX1 memory_reg_43__1_ ( .D(n425), .CK(clk), .RN(rstn), .Q(memory[321])
         );
  DFFRHQX1 memory_reg_43__0_ ( .D(n424), .CK(clk), .RN(rstn), .Q(memory[320])
         );
  DFFRHQX1 memory_reg_47__15_ ( .D(n375), .CK(clk), .RN(rstn), .Q(memory[271])
         );
  DFFRHQX1 memory_reg_47__14_ ( .D(n374), .CK(clk), .RN(rstn), .Q(memory[270])
         );
  DFFRHQX1 memory_reg_47__13_ ( .D(n373), .CK(clk), .RN(rstn), .Q(memory[269])
         );
  DFFRHQX1 memory_reg_47__12_ ( .D(n372), .CK(clk), .RN(rstn), .Q(memory[268])
         );
  DFFRHQX1 memory_reg_47__11_ ( .D(n371), .CK(clk), .RN(rstn), .Q(memory[267])
         );
  DFFRHQX1 memory_reg_47__10_ ( .D(n370), .CK(clk), .RN(rstn), .Q(memory[266])
         );
  DFFRHQX1 memory_reg_47__9_ ( .D(n369), .CK(clk), .RN(rstn), .Q(memory[265])
         );
  DFFRHQX1 memory_reg_47__8_ ( .D(n368), .CK(clk), .RN(rstn), .Q(memory[264])
         );
  DFFRHQX1 memory_reg_47__7_ ( .D(n367), .CK(clk), .RN(rstn), .Q(memory[263])
         );
  DFFRHQX1 memory_reg_47__6_ ( .D(n366), .CK(clk), .RN(rstn), .Q(memory[262])
         );
  DFFRHQX1 memory_reg_47__5_ ( .D(n365), .CK(clk), .RN(rstn), .Q(memory[261])
         );
  DFFRHQX1 memory_reg_47__4_ ( .D(n364), .CK(clk), .RN(rstn), .Q(memory[260])
         );
  DFFRHQX1 memory_reg_47__3_ ( .D(n363), .CK(clk), .RN(rstn), .Q(memory[259])
         );
  DFFRHQX1 memory_reg_47__2_ ( .D(n362), .CK(clk), .RN(rstn), .Q(memory[258])
         );
  DFFRHQX1 memory_reg_47__1_ ( .D(n361), .CK(clk), .RN(rstn), .Q(memory[257])
         );
  DFFRHQX1 memory_reg_47__0_ ( .D(n360), .CK(clk), .RN(rstn), .Q(memory[256])
         );
  DFFRHQX1 memory_reg_51__15_ ( .D(n311), .CK(clk), .RN(rstn), .Q(memory[207])
         );
  DFFRHQX1 memory_reg_51__14_ ( .D(n310), .CK(clk), .RN(rstn), .Q(memory[206])
         );
  DFFRHQX1 memory_reg_51__13_ ( .D(n309), .CK(clk), .RN(rstn), .Q(memory[205])
         );
  DFFRHQX1 memory_reg_51__12_ ( .D(n308), .CK(clk), .RN(rstn), .Q(memory[204])
         );
  DFFRHQX1 memory_reg_51__11_ ( .D(n307), .CK(clk), .RN(rstn), .Q(memory[203])
         );
  DFFRHQX1 memory_reg_51__10_ ( .D(n306), .CK(clk), .RN(rstn), .Q(memory[202])
         );
  DFFRHQX1 memory_reg_51__9_ ( .D(n305), .CK(clk), .RN(rstn), .Q(memory[201])
         );
  DFFRHQX1 memory_reg_51__8_ ( .D(n304), .CK(clk), .RN(rstn), .Q(memory[200])
         );
  DFFRHQX1 memory_reg_51__7_ ( .D(n303), .CK(clk), .RN(rstn), .Q(memory[199])
         );
  DFFRHQX1 memory_reg_51__6_ ( .D(n302), .CK(clk), .RN(rstn), .Q(memory[198])
         );
  DFFRHQX1 memory_reg_51__5_ ( .D(n301), .CK(clk), .RN(rstn), .Q(memory[197])
         );
  DFFRHQX1 memory_reg_51__4_ ( .D(n300), .CK(clk), .RN(rstn), .Q(memory[196])
         );
  DFFRHQX1 memory_reg_51__3_ ( .D(n299), .CK(clk), .RN(rstn), .Q(memory[195])
         );
  DFFRHQX1 memory_reg_51__2_ ( .D(n298), .CK(clk), .RN(rstn), .Q(memory[194])
         );
  DFFRHQX1 memory_reg_51__1_ ( .D(n297), .CK(clk), .RN(rstn), .Q(memory[193])
         );
  DFFRHQX1 memory_reg_51__0_ ( .D(n296), .CK(clk), .RN(rstn), .Q(memory[192])
         );
  DFFRHQX1 memory_reg_55__15_ ( .D(n247), .CK(clk), .RN(rstn), .Q(memory[143])
         );
  DFFRHQX1 memory_reg_55__14_ ( .D(n246), .CK(clk), .RN(rstn), .Q(memory[142])
         );
  DFFRHQX1 memory_reg_55__13_ ( .D(n245), .CK(clk), .RN(rstn), .Q(memory[141])
         );
  DFFRHQX1 memory_reg_55__12_ ( .D(n244), .CK(clk), .RN(rstn), .Q(memory[140])
         );
  DFFRHQX1 memory_reg_55__11_ ( .D(n243), .CK(clk), .RN(rstn), .Q(memory[139])
         );
  DFFRHQX1 memory_reg_55__10_ ( .D(n242), .CK(clk), .RN(rstn), .Q(memory[138])
         );
  DFFRHQX1 memory_reg_55__9_ ( .D(n241), .CK(clk), .RN(rstn), .Q(memory[137])
         );
  DFFRHQX1 memory_reg_55__8_ ( .D(n240), .CK(clk), .RN(rstn), .Q(memory[136])
         );
  DFFRHQX1 memory_reg_55__7_ ( .D(n239), .CK(clk), .RN(rstn), .Q(memory[135])
         );
  DFFRHQX1 memory_reg_55__6_ ( .D(n238), .CK(clk), .RN(rstn), .Q(memory[134])
         );
  DFFRHQX1 memory_reg_55__5_ ( .D(n237), .CK(clk), .RN(rstn), .Q(memory[133])
         );
  DFFRHQX1 memory_reg_55__4_ ( .D(n236), .CK(clk), .RN(rstn), .Q(memory[132])
         );
  DFFRHQX1 memory_reg_55__3_ ( .D(n235), .CK(clk), .RN(rstn), .Q(memory[131])
         );
  DFFRHQX1 memory_reg_55__2_ ( .D(n234), .CK(clk), .RN(rstn), .Q(memory[130])
         );
  DFFRHQX1 memory_reg_55__1_ ( .D(n233), .CK(clk), .RN(rstn), .Q(memory[129])
         );
  DFFRHQX1 memory_reg_55__0_ ( .D(n232), .CK(clk), .RN(rstn), .Q(memory[128])
         );
  DFFRHQX1 memory_reg_59__15_ ( .D(n183), .CK(clk), .RN(rstn), .Q(memory[79])
         );
  DFFRHQX1 memory_reg_59__14_ ( .D(n182), .CK(clk), .RN(rstn), .Q(memory[78])
         );
  DFFRHQX1 memory_reg_59__13_ ( .D(n181), .CK(clk), .RN(rstn), .Q(memory[77])
         );
  DFFRHQX1 memory_reg_59__12_ ( .D(n180), .CK(clk), .RN(rstn), .Q(memory[76])
         );
  DFFRHQX1 memory_reg_59__11_ ( .D(n179), .CK(clk), .RN(rstn), .Q(memory[75])
         );
  DFFRHQX1 memory_reg_59__10_ ( .D(n178), .CK(clk), .RN(rstn), .Q(memory[74])
         );
  DFFRHQX1 memory_reg_59__9_ ( .D(n177), .CK(clk), .RN(rstn), .Q(memory[73])
         );
  DFFRHQX1 memory_reg_59__8_ ( .D(n176), .CK(clk), .RN(rstn), .Q(memory[72])
         );
  DFFRHQX1 memory_reg_59__7_ ( .D(n175), .CK(clk), .RN(rstn), .Q(memory[71])
         );
  DFFRHQX1 memory_reg_59__6_ ( .D(n174), .CK(clk), .RN(rstn), .Q(memory[70])
         );
  DFFRHQX1 memory_reg_59__5_ ( .D(n173), .CK(clk), .RN(rstn), .Q(memory[69])
         );
  DFFRHQX1 memory_reg_59__4_ ( .D(n172), .CK(clk), .RN(rstn), .Q(memory[68])
         );
  DFFRHQX1 memory_reg_59__3_ ( .D(n171), .CK(clk), .RN(rstn), .Q(memory[67])
         );
  DFFRHQX1 memory_reg_59__2_ ( .D(n170), .CK(clk), .RN(rstn), .Q(memory[66])
         );
  DFFRHQX1 memory_reg_59__1_ ( .D(n169), .CK(clk), .RN(rstn), .Q(memory[65])
         );
  DFFRHQX1 memory_reg_59__0_ ( .D(n168), .CK(clk), .RN(rstn), .Q(memory[64])
         );
  DFFRHQX1 memory_reg_63__15_ ( .D(n119), .CK(clk), .RN(rstn), .Q(memory[15])
         );
  DFFRHQX1 memory_reg_63__14_ ( .D(n118), .CK(clk), .RN(rstn), .Q(memory[14])
         );
  DFFRHQX1 memory_reg_63__13_ ( .D(n117), .CK(clk), .RN(rstn), .Q(memory[13])
         );
  DFFRHQX1 memory_reg_63__12_ ( .D(n116), .CK(clk), .RN(rstn), .Q(memory[12])
         );
  DFFRHQX1 memory_reg_63__11_ ( .D(n115), .CK(clk), .RN(rstn), .Q(memory[11])
         );
  DFFRHQX1 memory_reg_63__10_ ( .D(n114), .CK(clk), .RN(rstn), .Q(memory[10])
         );
  DFFRHQX1 memory_reg_63__9_ ( .D(n113), .CK(clk), .RN(rstn), .Q(memory[9]) );
  DFFRHQX1 memory_reg_63__8_ ( .D(n112), .CK(clk), .RN(rstn), .Q(memory[8]) );
  DFFRHQX1 memory_reg_63__7_ ( .D(n111), .CK(clk), .RN(rstn), .Q(memory[7]) );
  DFFRHQX1 memory_reg_63__6_ ( .D(n110), .CK(clk), .RN(rstn), .Q(memory[6]) );
  DFFRHQX1 memory_reg_63__5_ ( .D(n109), .CK(clk), .RN(rstn), .Q(memory[5]) );
  DFFRHQX1 memory_reg_63__4_ ( .D(n108), .CK(clk), .RN(rstn), .Q(memory[4]) );
  DFFRHQX1 memory_reg_63__3_ ( .D(n107), .CK(clk), .RN(rstn), .Q(memory[3]) );
  DFFRHQX1 memory_reg_63__2_ ( .D(n106), .CK(clk), .RN(rstn), .Q(memory[2]) );
  DFFRHQX1 memory_reg_63__1_ ( .D(n105), .CK(clk), .RN(rstn), .Q(memory[1]) );
  DFFRHQX1 memory_reg_63__0_ ( .D(n104), .CK(clk), .RN(rstn), .Q(memory[0]) );
  DFFRHQX1 memory_reg_0__15_ ( .D(n1127), .CK(clk), .RN(rstn), .Q(memory[1023]) );
  DFFRHQX1 memory_reg_0__14_ ( .D(n1126), .CK(clk), .RN(rstn), .Q(memory[1022]) );
  DFFRHQX1 memory_reg_0__13_ ( .D(n1125), .CK(clk), .RN(rstn), .Q(memory[1021]) );
  DFFRHQX1 memory_reg_0__12_ ( .D(n1124), .CK(clk), .RN(rstn), .Q(memory[1020]) );
  DFFRHQX1 memory_reg_0__11_ ( .D(n1123), .CK(clk), .RN(rstn), .Q(memory[1019]) );
  DFFRHQX1 memory_reg_0__10_ ( .D(n1122), .CK(clk), .RN(rstn), .Q(memory[1018]) );
  DFFRHQX1 memory_reg_0__9_ ( .D(n1121), .CK(clk), .RN(rstn), .Q(memory[1017])
         );
  DFFRHQX1 memory_reg_0__8_ ( .D(n1120), .CK(clk), .RN(rstn), .Q(memory[1016])
         );
  DFFRHQX1 memory_reg_0__7_ ( .D(n1119), .CK(clk), .RN(rstn), .Q(memory[1015])
         );
  DFFRHQX1 memory_reg_0__6_ ( .D(n1118), .CK(clk), .RN(rstn), .Q(memory[1014])
         );
  DFFRHQX1 memory_reg_0__5_ ( .D(n1117), .CK(clk), .RN(rstn), .Q(memory[1013])
         );
  DFFRHQX1 memory_reg_0__4_ ( .D(n1116), .CK(clk), .RN(rstn), .Q(memory[1012])
         );
  DFFRHQX1 memory_reg_0__3_ ( .D(n1115), .CK(clk), .RN(rstn), .Q(memory[1011])
         );
  DFFRHQX1 memory_reg_0__2_ ( .D(n1114), .CK(clk), .RN(rstn), .Q(memory[1010])
         );
  DFFRHQX1 memory_reg_0__1_ ( .D(n1113), .CK(clk), .RN(rstn), .Q(memory[1009])
         );
  DFFRHQX1 memory_reg_0__0_ ( .D(n1112), .CK(clk), .RN(rstn), .Q(memory[1008])
         );
  DFFRHQX1 memory_reg_4__15_ ( .D(n1063), .CK(clk), .RN(rstn), .Q(memory[959])
         );
  DFFRHQX1 memory_reg_4__14_ ( .D(n1062), .CK(clk), .RN(rstn), .Q(memory[958])
         );
  DFFRHQX1 memory_reg_4__13_ ( .D(n1061), .CK(clk), .RN(rstn), .Q(memory[957])
         );
  DFFRHQX1 memory_reg_4__12_ ( .D(n1060), .CK(clk), .RN(rstn), .Q(memory[956])
         );
  DFFRHQX1 memory_reg_4__11_ ( .D(n1059), .CK(clk), .RN(rstn), .Q(memory[955])
         );
  DFFRHQX1 memory_reg_4__10_ ( .D(n1058), .CK(clk), .RN(rstn), .Q(memory[954])
         );
  DFFRHQX1 memory_reg_4__9_ ( .D(n1057), .CK(clk), .RN(rstn), .Q(memory[953])
         );
  DFFRHQX1 memory_reg_4__8_ ( .D(n1056), .CK(clk), .RN(rstn), .Q(memory[952])
         );
  DFFRHQX1 memory_reg_4__7_ ( .D(n1055), .CK(clk), .RN(rstn), .Q(memory[951])
         );
  DFFRHQX1 memory_reg_4__6_ ( .D(n1054), .CK(clk), .RN(rstn), .Q(memory[950])
         );
  DFFRHQX1 memory_reg_4__5_ ( .D(n1053), .CK(clk), .RN(rstn), .Q(memory[949])
         );
  DFFRHQX1 memory_reg_4__4_ ( .D(n1052), .CK(clk), .RN(rstn), .Q(memory[948])
         );
  DFFRHQX1 memory_reg_4__3_ ( .D(n1051), .CK(clk), .RN(rstn), .Q(memory[947])
         );
  DFFRHQX1 memory_reg_4__2_ ( .D(n1050), .CK(clk), .RN(rstn), .Q(memory[946])
         );
  DFFRHQX1 memory_reg_4__1_ ( .D(n1049), .CK(clk), .RN(rstn), .Q(memory[945])
         );
  DFFRHQX1 memory_reg_4__0_ ( .D(n1048), .CK(clk), .RN(rstn), .Q(memory[944])
         );
  DFFRHQX1 memory_reg_8__15_ ( .D(n999), .CK(clk), .RN(rstn), .Q(memory[895])
         );
  DFFRHQX1 memory_reg_8__14_ ( .D(n998), .CK(clk), .RN(rstn), .Q(memory[894])
         );
  DFFRHQX1 memory_reg_8__13_ ( .D(n997), .CK(clk), .RN(rstn), .Q(memory[893])
         );
  DFFRHQX1 memory_reg_8__12_ ( .D(n996), .CK(clk), .RN(rstn), .Q(memory[892])
         );
  DFFRHQX1 memory_reg_8__11_ ( .D(n995), .CK(clk), .RN(rstn), .Q(memory[891])
         );
  DFFRHQX1 memory_reg_8__10_ ( .D(n994), .CK(clk), .RN(rstn), .Q(memory[890])
         );
  DFFRHQX1 memory_reg_8__9_ ( .D(n993), .CK(clk), .RN(rstn), .Q(memory[889])
         );
  DFFRHQX1 memory_reg_8__8_ ( .D(n992), .CK(clk), .RN(rstn), .Q(memory[888])
         );
  DFFRHQX1 memory_reg_8__7_ ( .D(n991), .CK(clk), .RN(rstn), .Q(memory[887])
         );
  DFFRHQX1 memory_reg_8__6_ ( .D(n990), .CK(clk), .RN(rstn), .Q(memory[886])
         );
  DFFRHQX1 memory_reg_8__5_ ( .D(n989), .CK(clk), .RN(rstn), .Q(memory[885])
         );
  DFFRHQX1 memory_reg_8__4_ ( .D(n988), .CK(clk), .RN(rstn), .Q(memory[884])
         );
  DFFRHQX1 memory_reg_8__3_ ( .D(n987), .CK(clk), .RN(rstn), .Q(memory[883])
         );
  DFFRHQX1 memory_reg_8__2_ ( .D(n986), .CK(clk), .RN(rstn), .Q(memory[882])
         );
  DFFRHQX1 memory_reg_8__1_ ( .D(n985), .CK(clk), .RN(rstn), .Q(memory[881])
         );
  DFFRHQX1 memory_reg_8__0_ ( .D(n984), .CK(clk), .RN(rstn), .Q(memory[880])
         );
  DFFRHQX1 memory_reg_12__15_ ( .D(n935), .CK(clk), .RN(rstn), .Q(memory[831])
         );
  DFFRHQX1 memory_reg_12__14_ ( .D(n934), .CK(clk), .RN(rstn), .Q(memory[830])
         );
  DFFRHQX1 memory_reg_12__13_ ( .D(n933), .CK(clk), .RN(rstn), .Q(memory[829])
         );
  DFFRHQX1 memory_reg_12__12_ ( .D(n932), .CK(clk), .RN(rstn), .Q(memory[828])
         );
  DFFRHQX1 memory_reg_12__11_ ( .D(n931), .CK(clk), .RN(rstn), .Q(memory[827])
         );
  DFFRHQX1 memory_reg_12__10_ ( .D(n930), .CK(clk), .RN(rstn), .Q(memory[826])
         );
  DFFRHQX1 memory_reg_12__9_ ( .D(n929), .CK(clk), .RN(rstn), .Q(memory[825])
         );
  DFFRHQX1 memory_reg_12__8_ ( .D(n928), .CK(clk), .RN(rstn), .Q(memory[824])
         );
  DFFRHQX1 memory_reg_12__7_ ( .D(n927), .CK(clk), .RN(rstn), .Q(memory[823])
         );
  DFFRHQX1 memory_reg_12__6_ ( .D(n926), .CK(clk), .RN(rstn), .Q(memory[822])
         );
  DFFRHQX1 memory_reg_12__5_ ( .D(n925), .CK(clk), .RN(rstn), .Q(memory[821])
         );
  DFFRHQX1 memory_reg_12__4_ ( .D(n924), .CK(clk), .RN(rstn), .Q(memory[820])
         );
  DFFRHQX1 memory_reg_12__3_ ( .D(n923), .CK(clk), .RN(rstn), .Q(memory[819])
         );
  DFFRHQX1 memory_reg_12__2_ ( .D(n922), .CK(clk), .RN(rstn), .Q(memory[818])
         );
  DFFRHQX1 memory_reg_12__1_ ( .D(n921), .CK(clk), .RN(rstn), .Q(memory[817])
         );
  DFFRHQX1 memory_reg_12__0_ ( .D(n920), .CK(clk), .RN(rstn), .Q(memory[816])
         );
  DFFRHQX1 memory_reg_16__15_ ( .D(n871), .CK(clk), .RN(rstn), .Q(memory[767])
         );
  DFFRHQX1 memory_reg_16__14_ ( .D(n870), .CK(clk), .RN(rstn), .Q(memory[766])
         );
  DFFRHQX1 memory_reg_16__13_ ( .D(n869), .CK(clk), .RN(rstn), .Q(memory[765])
         );
  DFFRHQX1 memory_reg_16__12_ ( .D(n868), .CK(clk), .RN(rstn), .Q(memory[764])
         );
  DFFRHQX1 memory_reg_16__11_ ( .D(n867), .CK(clk), .RN(rstn), .Q(memory[763])
         );
  DFFRHQX1 memory_reg_16__10_ ( .D(n866), .CK(clk), .RN(rstn), .Q(memory[762])
         );
  DFFRHQX1 memory_reg_16__9_ ( .D(n865), .CK(clk), .RN(rstn), .Q(memory[761])
         );
  DFFRHQX1 memory_reg_16__8_ ( .D(n864), .CK(clk), .RN(rstn), .Q(memory[760])
         );
  DFFRHQX1 memory_reg_16__7_ ( .D(n863), .CK(clk), .RN(rstn), .Q(memory[759])
         );
  DFFRHQX1 memory_reg_16__6_ ( .D(n862), .CK(clk), .RN(rstn), .Q(memory[758])
         );
  DFFRHQX1 memory_reg_16__5_ ( .D(n861), .CK(clk), .RN(rstn), .Q(memory[757])
         );
  DFFRHQX1 memory_reg_16__4_ ( .D(n860), .CK(clk), .RN(rstn), .Q(memory[756])
         );
  DFFRHQX1 memory_reg_16__3_ ( .D(n859), .CK(clk), .RN(rstn), .Q(memory[755])
         );
  DFFRHQX1 memory_reg_16__2_ ( .D(n858), .CK(clk), .RN(rstn), .Q(memory[754])
         );
  DFFRHQX1 memory_reg_16__1_ ( .D(n857), .CK(clk), .RN(rstn), .Q(memory[753])
         );
  DFFRHQX1 memory_reg_16__0_ ( .D(n856), .CK(clk), .RN(rstn), .Q(memory[752])
         );
  DFFRHQX1 memory_reg_20__15_ ( .D(n807), .CK(clk), .RN(rstn), .Q(memory[703])
         );
  DFFRHQX1 memory_reg_20__14_ ( .D(n806), .CK(clk), .RN(rstn), .Q(memory[702])
         );
  DFFRHQX1 memory_reg_20__13_ ( .D(n805), .CK(clk), .RN(rstn), .Q(memory[701])
         );
  DFFRHQX1 memory_reg_20__12_ ( .D(n804), .CK(clk), .RN(rstn), .Q(memory[700])
         );
  DFFRHQX1 memory_reg_20__11_ ( .D(n803), .CK(clk), .RN(rstn), .Q(memory[699])
         );
  DFFRHQX1 memory_reg_20__10_ ( .D(n802), .CK(clk), .RN(rstn), .Q(memory[698])
         );
  DFFRHQX1 memory_reg_20__9_ ( .D(n801), .CK(clk), .RN(rstn), .Q(memory[697])
         );
  DFFRHQX1 memory_reg_20__8_ ( .D(n800), .CK(clk), .RN(rstn), .Q(memory[696])
         );
  DFFRHQX1 memory_reg_20__7_ ( .D(n799), .CK(clk), .RN(rstn), .Q(memory[695])
         );
  DFFRHQX1 memory_reg_20__6_ ( .D(n798), .CK(clk), .RN(rstn), .Q(memory[694])
         );
  DFFRHQX1 memory_reg_20__5_ ( .D(n797), .CK(clk), .RN(rstn), .Q(memory[693])
         );
  DFFRHQX1 memory_reg_20__4_ ( .D(n796), .CK(clk), .RN(rstn), .Q(memory[692])
         );
  DFFRHQX1 memory_reg_20__3_ ( .D(n795), .CK(clk), .RN(rstn), .Q(memory[691])
         );
  DFFRHQX1 memory_reg_20__2_ ( .D(n794), .CK(clk), .RN(rstn), .Q(memory[690])
         );
  DFFRHQX1 memory_reg_20__1_ ( .D(n793), .CK(clk), .RN(rstn), .Q(memory[689])
         );
  DFFRHQX1 memory_reg_20__0_ ( .D(n792), .CK(clk), .RN(rstn), .Q(memory[688])
         );
  DFFRHQX1 memory_reg_24__15_ ( .D(n743), .CK(clk), .RN(rstn), .Q(memory[639])
         );
  DFFRHQX1 memory_reg_24__14_ ( .D(n742), .CK(clk), .RN(rstn), .Q(memory[638])
         );
  DFFRHQX1 memory_reg_24__13_ ( .D(n741), .CK(clk), .RN(rstn), .Q(memory[637])
         );
  DFFRHQX1 memory_reg_24__12_ ( .D(n740), .CK(clk), .RN(rstn), .Q(memory[636])
         );
  DFFRHQX1 memory_reg_24__11_ ( .D(n739), .CK(clk), .RN(rstn), .Q(memory[635])
         );
  DFFRHQX1 memory_reg_24__10_ ( .D(n738), .CK(clk), .RN(rstn), .Q(memory[634])
         );
  DFFRHQX1 memory_reg_24__9_ ( .D(n737), .CK(clk), .RN(rstn), .Q(memory[633])
         );
  DFFRHQX1 memory_reg_24__8_ ( .D(n736), .CK(clk), .RN(rstn), .Q(memory[632])
         );
  DFFRHQX1 memory_reg_24__7_ ( .D(n735), .CK(clk), .RN(rstn), .Q(memory[631])
         );
  DFFRHQX1 memory_reg_24__6_ ( .D(n734), .CK(clk), .RN(rstn), .Q(memory[630])
         );
  DFFRHQX1 memory_reg_24__5_ ( .D(n733), .CK(clk), .RN(rstn), .Q(memory[629])
         );
  DFFRHQX1 memory_reg_24__4_ ( .D(n732), .CK(clk), .RN(rstn), .Q(memory[628])
         );
  DFFRHQX1 memory_reg_24__3_ ( .D(n731), .CK(clk), .RN(rstn), .Q(memory[627])
         );
  DFFRHQX1 memory_reg_24__2_ ( .D(n730), .CK(clk), .RN(rstn), .Q(memory[626])
         );
  DFFRHQX1 memory_reg_24__1_ ( .D(n729), .CK(clk), .RN(rstn), .Q(memory[625])
         );
  DFFRHQX1 memory_reg_24__0_ ( .D(n728), .CK(clk), .RN(rstn), .Q(memory[624])
         );
  DFFRHQX1 memory_reg_28__15_ ( .D(n679), .CK(clk), .RN(rstn), .Q(memory[575])
         );
  DFFRHQX1 memory_reg_28__14_ ( .D(n678), .CK(clk), .RN(rstn), .Q(memory[574])
         );
  DFFRHQX1 memory_reg_28__13_ ( .D(n677), .CK(clk), .RN(rstn), .Q(memory[573])
         );
  DFFRHQX1 memory_reg_28__12_ ( .D(n676), .CK(clk), .RN(rstn), .Q(memory[572])
         );
  DFFRHQX1 memory_reg_28__11_ ( .D(n675), .CK(clk), .RN(rstn), .Q(memory[571])
         );
  DFFRHQX1 memory_reg_28__10_ ( .D(n674), .CK(clk), .RN(rstn), .Q(memory[570])
         );
  DFFRHQX1 memory_reg_28__9_ ( .D(n673), .CK(clk), .RN(rstn), .Q(memory[569])
         );
  DFFRHQX1 memory_reg_28__8_ ( .D(n672), .CK(clk), .RN(rstn), .Q(memory[568])
         );
  DFFRHQX1 memory_reg_28__7_ ( .D(n671), .CK(clk), .RN(rstn), .Q(memory[567])
         );
  DFFRHQX1 memory_reg_28__6_ ( .D(n670), .CK(clk), .RN(rstn), .Q(memory[566])
         );
  DFFRHQX1 memory_reg_28__5_ ( .D(n669), .CK(clk), .RN(rstn), .Q(memory[565])
         );
  DFFRHQX1 memory_reg_28__4_ ( .D(n668), .CK(clk), .RN(rstn), .Q(memory[564])
         );
  DFFRHQX1 memory_reg_28__3_ ( .D(n667), .CK(clk), .RN(rstn), .Q(memory[563])
         );
  DFFRHQX1 memory_reg_28__2_ ( .D(n666), .CK(clk), .RN(rstn), .Q(memory[562])
         );
  DFFRHQX1 memory_reg_28__1_ ( .D(n665), .CK(clk), .RN(rstn), .Q(memory[561])
         );
  DFFRHQX1 memory_reg_28__0_ ( .D(n664), .CK(clk), .RN(rstn), .Q(memory[560])
         );
  DFFRHQX1 memory_reg_32__15_ ( .D(n615), .CK(clk), .RN(rstn), .Q(memory[511])
         );
  DFFRHQX1 memory_reg_32__14_ ( .D(n614), .CK(clk), .RN(rstn), .Q(memory[510])
         );
  DFFRHQX1 memory_reg_32__13_ ( .D(n613), .CK(clk), .RN(rstn), .Q(memory[509])
         );
  DFFRHQX1 memory_reg_32__12_ ( .D(n612), .CK(clk), .RN(rstn), .Q(memory[508])
         );
  DFFRHQX1 memory_reg_32__11_ ( .D(n611), .CK(clk), .RN(rstn), .Q(memory[507])
         );
  DFFRHQX1 memory_reg_32__10_ ( .D(n610), .CK(clk), .RN(rstn), .Q(memory[506])
         );
  DFFRHQX1 memory_reg_32__9_ ( .D(n609), .CK(clk), .RN(rstn), .Q(memory[505])
         );
  DFFRHQX1 memory_reg_32__8_ ( .D(n608), .CK(clk), .RN(rstn), .Q(memory[504])
         );
  DFFRHQX1 memory_reg_32__7_ ( .D(n607), .CK(clk), .RN(rstn), .Q(memory[503])
         );
  DFFRHQX1 memory_reg_32__6_ ( .D(n606), .CK(clk), .RN(rstn), .Q(memory[502])
         );
  DFFRHQX1 memory_reg_32__5_ ( .D(n605), .CK(clk), .RN(rstn), .Q(memory[501])
         );
  DFFRHQX1 memory_reg_32__4_ ( .D(n604), .CK(clk), .RN(rstn), .Q(memory[500])
         );
  DFFRHQX1 memory_reg_32__3_ ( .D(n603), .CK(clk), .RN(rstn), .Q(memory[499])
         );
  DFFRHQX1 memory_reg_32__2_ ( .D(n602), .CK(clk), .RN(rstn), .Q(memory[498])
         );
  DFFRHQX1 memory_reg_32__1_ ( .D(n601), .CK(clk), .RN(rstn), .Q(memory[497])
         );
  DFFRHQX1 memory_reg_32__0_ ( .D(n600), .CK(clk), .RN(rstn), .Q(memory[496])
         );
  DFFRHQX1 memory_reg_36__15_ ( .D(n551), .CK(clk), .RN(rstn), .Q(memory[447])
         );
  DFFRHQX1 memory_reg_36__14_ ( .D(n550), .CK(clk), .RN(rstn), .Q(memory[446])
         );
  DFFRHQX1 memory_reg_36__13_ ( .D(n549), .CK(clk), .RN(rstn), .Q(memory[445])
         );
  DFFRHQX1 memory_reg_36__12_ ( .D(n548), .CK(clk), .RN(rstn), .Q(memory[444])
         );
  DFFRHQX1 memory_reg_36__11_ ( .D(n547), .CK(clk), .RN(rstn), .Q(memory[443])
         );
  DFFRHQX1 memory_reg_36__10_ ( .D(n546), .CK(clk), .RN(rstn), .Q(memory[442])
         );
  DFFRHQX1 memory_reg_36__9_ ( .D(n545), .CK(clk), .RN(rstn), .Q(memory[441])
         );
  DFFRHQX1 memory_reg_36__8_ ( .D(n544), .CK(clk), .RN(rstn), .Q(memory[440])
         );
  DFFRHQX1 memory_reg_36__7_ ( .D(n543), .CK(clk), .RN(rstn), .Q(memory[439])
         );
  DFFRHQX1 memory_reg_36__6_ ( .D(n542), .CK(clk), .RN(rstn), .Q(memory[438])
         );
  DFFRHQX1 memory_reg_36__5_ ( .D(n541), .CK(clk), .RN(rstn), .Q(memory[437])
         );
  DFFRHQX1 memory_reg_36__4_ ( .D(n540), .CK(clk), .RN(rstn), .Q(memory[436])
         );
  DFFRHQX1 memory_reg_36__3_ ( .D(n539), .CK(clk), .RN(rstn), .Q(memory[435])
         );
  DFFRHQX1 memory_reg_36__2_ ( .D(n538), .CK(clk), .RN(rstn), .Q(memory[434])
         );
  DFFRHQX1 memory_reg_36__1_ ( .D(n537), .CK(clk), .RN(rstn), .Q(memory[433])
         );
  DFFRHQX1 memory_reg_36__0_ ( .D(n536), .CK(clk), .RN(rstn), .Q(memory[432])
         );
  DFFRHQX1 memory_reg_40__15_ ( .D(n487), .CK(clk), .RN(rstn), .Q(memory[383])
         );
  DFFRHQX1 memory_reg_40__14_ ( .D(n486), .CK(clk), .RN(rstn), .Q(memory[382])
         );
  DFFRHQX1 memory_reg_40__13_ ( .D(n485), .CK(clk), .RN(rstn), .Q(memory[381])
         );
  DFFRHQX1 memory_reg_40__12_ ( .D(n484), .CK(clk), .RN(rstn), .Q(memory[380])
         );
  DFFRHQX1 memory_reg_40__11_ ( .D(n483), .CK(clk), .RN(rstn), .Q(memory[379])
         );
  DFFRHQX1 memory_reg_40__10_ ( .D(n482), .CK(clk), .RN(rstn), .Q(memory[378])
         );
  DFFRHQX1 memory_reg_40__9_ ( .D(n481), .CK(clk), .RN(rstn), .Q(memory[377])
         );
  DFFRHQX1 memory_reg_40__8_ ( .D(n480), .CK(clk), .RN(rstn), .Q(memory[376])
         );
  DFFRHQX1 memory_reg_40__7_ ( .D(n479), .CK(clk), .RN(rstn), .Q(memory[375])
         );
  DFFRHQX1 memory_reg_40__6_ ( .D(n478), .CK(clk), .RN(rstn), .Q(memory[374])
         );
  DFFRHQX1 memory_reg_40__5_ ( .D(n477), .CK(clk), .RN(rstn), .Q(memory[373])
         );
  DFFRHQX1 memory_reg_40__4_ ( .D(n476), .CK(clk), .RN(rstn), .Q(memory[372])
         );
  DFFRHQX1 memory_reg_40__3_ ( .D(n475), .CK(clk), .RN(rstn), .Q(memory[371])
         );
  DFFRHQX1 memory_reg_40__2_ ( .D(n474), .CK(clk), .RN(rstn), .Q(memory[370])
         );
  DFFRHQX1 memory_reg_40__1_ ( .D(n473), .CK(clk), .RN(rstn), .Q(memory[369])
         );
  DFFRHQX1 memory_reg_40__0_ ( .D(n472), .CK(clk), .RN(rstn), .Q(memory[368])
         );
  DFFRHQX1 memory_reg_44__15_ ( .D(n423), .CK(clk), .RN(rstn), .Q(memory[319])
         );
  DFFRHQX1 memory_reg_44__14_ ( .D(n422), .CK(clk), .RN(rstn), .Q(memory[318])
         );
  DFFRHQX1 memory_reg_44__13_ ( .D(n421), .CK(clk), .RN(rstn), .Q(memory[317])
         );
  DFFRHQX1 memory_reg_44__12_ ( .D(n420), .CK(clk), .RN(rstn), .Q(memory[316])
         );
  DFFRHQX1 memory_reg_44__11_ ( .D(n419), .CK(clk), .RN(rstn), .Q(memory[315])
         );
  DFFRHQX1 memory_reg_44__10_ ( .D(n418), .CK(clk), .RN(rstn), .Q(memory[314])
         );
  DFFRHQX1 memory_reg_44__9_ ( .D(n417), .CK(clk), .RN(rstn), .Q(memory[313])
         );
  DFFRHQX1 memory_reg_44__8_ ( .D(n416), .CK(clk), .RN(rstn), .Q(memory[312])
         );
  DFFRHQX1 memory_reg_44__7_ ( .D(n415), .CK(clk), .RN(rstn), .Q(memory[311])
         );
  DFFRHQX1 memory_reg_44__6_ ( .D(n414), .CK(clk), .RN(rstn), .Q(memory[310])
         );
  DFFRHQX1 memory_reg_44__5_ ( .D(n413), .CK(clk), .RN(rstn), .Q(memory[309])
         );
  DFFRHQX1 memory_reg_44__4_ ( .D(n412), .CK(clk), .RN(rstn), .Q(memory[308])
         );
  DFFRHQX1 memory_reg_44__3_ ( .D(n411), .CK(clk), .RN(rstn), .Q(memory[307])
         );
  DFFRHQX1 memory_reg_44__2_ ( .D(n410), .CK(clk), .RN(rstn), .Q(memory[306])
         );
  DFFRHQX1 memory_reg_44__1_ ( .D(n409), .CK(clk), .RN(rstn), .Q(memory[305])
         );
  DFFRHQX1 memory_reg_44__0_ ( .D(n408), .CK(clk), .RN(rstn), .Q(memory[304])
         );
  DFFRHQX1 memory_reg_48__15_ ( .D(n359), .CK(clk), .RN(rstn), .Q(memory[255])
         );
  DFFRHQX1 memory_reg_48__14_ ( .D(n358), .CK(clk), .RN(rstn), .Q(memory[254])
         );
  DFFRHQX1 memory_reg_48__13_ ( .D(n357), .CK(clk), .RN(rstn), .Q(memory[253])
         );
  DFFRHQX1 memory_reg_48__12_ ( .D(n356), .CK(clk), .RN(rstn), .Q(memory[252])
         );
  DFFRHQX1 memory_reg_48__11_ ( .D(n355), .CK(clk), .RN(rstn), .Q(memory[251])
         );
  DFFRHQX1 memory_reg_48__10_ ( .D(n354), .CK(clk), .RN(rstn), .Q(memory[250])
         );
  DFFRHQX1 memory_reg_48__9_ ( .D(n353), .CK(clk), .RN(rstn), .Q(memory[249])
         );
  DFFRHQX1 memory_reg_48__8_ ( .D(n352), .CK(clk), .RN(rstn), .Q(memory[248])
         );
  DFFRHQX1 memory_reg_48__7_ ( .D(n351), .CK(clk), .RN(rstn), .Q(memory[247])
         );
  DFFRHQX1 memory_reg_48__6_ ( .D(n350), .CK(clk), .RN(rstn), .Q(memory[246])
         );
  DFFRHQX1 memory_reg_48__5_ ( .D(n349), .CK(clk), .RN(rstn), .Q(memory[245])
         );
  DFFRHQX1 memory_reg_48__4_ ( .D(n348), .CK(clk), .RN(rstn), .Q(memory[244])
         );
  DFFRHQX1 memory_reg_48__3_ ( .D(n347), .CK(clk), .RN(rstn), .Q(memory[243])
         );
  DFFRHQX1 memory_reg_48__2_ ( .D(n346), .CK(clk), .RN(rstn), .Q(memory[242])
         );
  DFFRHQX1 memory_reg_48__1_ ( .D(n345), .CK(clk), .RN(rstn), .Q(memory[241])
         );
  DFFRHQX1 memory_reg_48__0_ ( .D(n344), .CK(clk), .RN(rstn), .Q(memory[240])
         );
  DFFRHQX1 memory_reg_52__15_ ( .D(n295), .CK(clk), .RN(rstn), .Q(memory[191])
         );
  DFFRHQX1 memory_reg_52__14_ ( .D(n294), .CK(clk), .RN(rstn), .Q(memory[190])
         );
  DFFRHQX1 memory_reg_52__13_ ( .D(n293), .CK(clk), .RN(rstn), .Q(memory[189])
         );
  DFFRHQX1 memory_reg_52__12_ ( .D(n292), .CK(clk), .RN(rstn), .Q(memory[188])
         );
  DFFRHQX1 memory_reg_52__11_ ( .D(n291), .CK(clk), .RN(rstn), .Q(memory[187])
         );
  DFFRHQX1 memory_reg_52__10_ ( .D(n290), .CK(clk), .RN(rstn), .Q(memory[186])
         );
  DFFRHQX1 memory_reg_52__9_ ( .D(n289), .CK(clk), .RN(rstn), .Q(memory[185])
         );
  DFFRHQX1 memory_reg_52__8_ ( .D(n288), .CK(clk), .RN(rstn), .Q(memory[184])
         );
  DFFRHQX1 memory_reg_52__7_ ( .D(n287), .CK(clk), .RN(rstn), .Q(memory[183])
         );
  DFFRHQX1 memory_reg_52__6_ ( .D(n286), .CK(clk), .RN(rstn), .Q(memory[182])
         );
  DFFRHQX1 memory_reg_52__5_ ( .D(n285), .CK(clk), .RN(rstn), .Q(memory[181])
         );
  DFFRHQX1 memory_reg_52__4_ ( .D(n284), .CK(clk), .RN(rstn), .Q(memory[180])
         );
  DFFRHQX1 memory_reg_52__3_ ( .D(n283), .CK(clk), .RN(rstn), .Q(memory[179])
         );
  DFFRHQX1 memory_reg_52__2_ ( .D(n282), .CK(clk), .RN(rstn), .Q(memory[178])
         );
  DFFRHQX1 memory_reg_52__1_ ( .D(n281), .CK(clk), .RN(rstn), .Q(memory[177])
         );
  DFFRHQX1 memory_reg_52__0_ ( .D(n280), .CK(clk), .RN(rstn), .Q(memory[176])
         );
  DFFRHQX1 memory_reg_56__15_ ( .D(n231), .CK(clk), .RN(rstn), .Q(memory[127])
         );
  DFFRHQX1 memory_reg_56__14_ ( .D(n230), .CK(clk), .RN(rstn), .Q(memory[126])
         );
  DFFRHQX1 memory_reg_56__13_ ( .D(n229), .CK(clk), .RN(rstn), .Q(memory[125])
         );
  DFFRHQX1 memory_reg_56__12_ ( .D(n228), .CK(clk), .RN(rstn), .Q(memory[124])
         );
  DFFRHQX1 memory_reg_56__11_ ( .D(n227), .CK(clk), .RN(rstn), .Q(memory[123])
         );
  DFFRHQX1 memory_reg_56__10_ ( .D(n226), .CK(clk), .RN(rstn), .Q(memory[122])
         );
  DFFRHQX1 memory_reg_56__9_ ( .D(n225), .CK(clk), .RN(rstn), .Q(memory[121])
         );
  DFFRHQX1 memory_reg_56__8_ ( .D(n224), .CK(clk), .RN(rstn), .Q(memory[120])
         );
  DFFRHQX1 memory_reg_56__7_ ( .D(n223), .CK(clk), .RN(rstn), .Q(memory[119])
         );
  DFFRHQX1 memory_reg_56__6_ ( .D(n222), .CK(clk), .RN(rstn), .Q(memory[118])
         );
  DFFRHQX1 memory_reg_56__5_ ( .D(n221), .CK(clk), .RN(rstn), .Q(memory[117])
         );
  DFFRHQX1 memory_reg_56__4_ ( .D(n220), .CK(clk), .RN(rstn), .Q(memory[116])
         );
  DFFRHQX1 memory_reg_56__3_ ( .D(n219), .CK(clk), .RN(rstn), .Q(memory[115])
         );
  DFFRHQX1 memory_reg_56__2_ ( .D(n218), .CK(clk), .RN(rstn), .Q(memory[114])
         );
  DFFRHQX1 memory_reg_56__1_ ( .D(n217), .CK(clk), .RN(rstn), .Q(memory[113])
         );
  DFFRHQX1 memory_reg_56__0_ ( .D(n216), .CK(clk), .RN(rstn), .Q(memory[112])
         );
  DFFRHQX1 memory_reg_60__15_ ( .D(n167), .CK(clk), .RN(rstn), .Q(memory[63])
         );
  DFFRHQX1 memory_reg_60__14_ ( .D(n166), .CK(clk), .RN(rstn), .Q(memory[62])
         );
  DFFRHQX1 memory_reg_60__13_ ( .D(n165), .CK(clk), .RN(rstn), .Q(memory[61])
         );
  DFFRHQX1 memory_reg_60__12_ ( .D(n164), .CK(clk), .RN(rstn), .Q(memory[60])
         );
  DFFRHQX1 memory_reg_60__11_ ( .D(n163), .CK(clk), .RN(rstn), .Q(memory[59])
         );
  DFFRHQX1 memory_reg_60__10_ ( .D(n162), .CK(clk), .RN(rstn), .Q(memory[58])
         );
  DFFRHQX1 memory_reg_60__9_ ( .D(n161), .CK(clk), .RN(rstn), .Q(memory[57])
         );
  DFFRHQX1 memory_reg_60__8_ ( .D(n160), .CK(clk), .RN(rstn), .Q(memory[56])
         );
  DFFRHQX1 memory_reg_60__7_ ( .D(n159), .CK(clk), .RN(rstn), .Q(memory[55])
         );
  DFFRHQX1 memory_reg_60__6_ ( .D(n158), .CK(clk), .RN(rstn), .Q(memory[54])
         );
  DFFRHQX1 memory_reg_60__5_ ( .D(n157), .CK(clk), .RN(rstn), .Q(memory[53])
         );
  DFFRHQX1 memory_reg_60__4_ ( .D(n156), .CK(clk), .RN(rstn), .Q(memory[52])
         );
  DFFRHQX1 memory_reg_60__3_ ( .D(n155), .CK(clk), .RN(rstn), .Q(memory[51])
         );
  DFFRHQX1 memory_reg_60__2_ ( .D(n154), .CK(clk), .RN(rstn), .Q(memory[50])
         );
  DFFRHQX1 memory_reg_60__1_ ( .D(n153), .CK(clk), .RN(rstn), .Q(memory[49])
         );
  DFFRHQX1 memory_reg_60__0_ ( .D(n152), .CK(clk), .RN(rstn), .Q(memory[48])
         );
  DFFRHQX1 memory_reg_2__15_ ( .D(n1095), .CK(clk), .RN(rstn), .Q(memory[991])
         );
  DFFRHQX1 memory_reg_2__14_ ( .D(n1094), .CK(clk), .RN(rstn), .Q(memory[990])
         );
  DFFRHQX1 memory_reg_2__13_ ( .D(n1093), .CK(clk), .RN(rstn), .Q(memory[989])
         );
  DFFRHQX1 memory_reg_2__12_ ( .D(n1092), .CK(clk), .RN(rstn), .Q(memory[988])
         );
  DFFRHQX1 memory_reg_2__11_ ( .D(n1091), .CK(clk), .RN(rstn), .Q(memory[987])
         );
  DFFRHQX1 memory_reg_2__10_ ( .D(n1090), .CK(clk), .RN(rstn), .Q(memory[986])
         );
  DFFRHQX1 memory_reg_2__9_ ( .D(n1089), .CK(clk), .RN(rstn), .Q(memory[985])
         );
  DFFRHQX1 memory_reg_2__8_ ( .D(n1088), .CK(clk), .RN(rstn), .Q(memory[984])
         );
  DFFRHQX1 memory_reg_2__7_ ( .D(n1087), .CK(clk), .RN(rstn), .Q(memory[983])
         );
  DFFRHQX1 memory_reg_2__6_ ( .D(n1086), .CK(clk), .RN(rstn), .Q(memory[982])
         );
  DFFRHQX1 memory_reg_2__5_ ( .D(n1085), .CK(clk), .RN(rstn), .Q(memory[981])
         );
  DFFRHQX1 memory_reg_2__4_ ( .D(n1084), .CK(clk), .RN(rstn), .Q(memory[980])
         );
  DFFRHQX1 memory_reg_2__3_ ( .D(n1083), .CK(clk), .RN(rstn), .Q(memory[979])
         );
  DFFRHQX1 memory_reg_2__2_ ( .D(n1082), .CK(clk), .RN(rstn), .Q(memory[978])
         );
  DFFRHQX1 memory_reg_2__1_ ( .D(n1081), .CK(clk), .RN(rstn), .Q(memory[977])
         );
  DFFRHQX1 memory_reg_2__0_ ( .D(n1080), .CK(clk), .RN(rstn), .Q(memory[976])
         );
  DFFRHQX1 memory_reg_6__15_ ( .D(n1031), .CK(clk), .RN(rstn), .Q(memory[927])
         );
  DFFRHQX1 memory_reg_6__14_ ( .D(n1030), .CK(clk), .RN(rstn), .Q(memory[926])
         );
  DFFRHQX1 memory_reg_6__13_ ( .D(n1029), .CK(clk), .RN(rstn), .Q(memory[925])
         );
  DFFRHQX1 memory_reg_6__12_ ( .D(n1028), .CK(clk), .RN(rstn), .Q(memory[924])
         );
  DFFRHQX1 memory_reg_6__11_ ( .D(n1027), .CK(clk), .RN(rstn), .Q(memory[923])
         );
  DFFRHQX1 memory_reg_6__10_ ( .D(n1026), .CK(clk), .RN(rstn), .Q(memory[922])
         );
  DFFRHQX1 memory_reg_6__9_ ( .D(n1025), .CK(clk), .RN(rstn), .Q(memory[921])
         );
  DFFRHQX1 memory_reg_6__8_ ( .D(n1024), .CK(clk), .RN(rstn), .Q(memory[920])
         );
  DFFRHQX1 memory_reg_6__7_ ( .D(n1023), .CK(clk), .RN(rstn), .Q(memory[919])
         );
  DFFRHQX1 memory_reg_6__6_ ( .D(n1022), .CK(clk), .RN(rstn), .Q(memory[918])
         );
  DFFRHQX1 memory_reg_6__5_ ( .D(n1021), .CK(clk), .RN(rstn), .Q(memory[917])
         );
  DFFRHQX1 memory_reg_6__4_ ( .D(n1020), .CK(clk), .RN(rstn), .Q(memory[916])
         );
  DFFRHQX1 memory_reg_6__3_ ( .D(n1019), .CK(clk), .RN(rstn), .Q(memory[915])
         );
  DFFRHQX1 memory_reg_6__2_ ( .D(n1018), .CK(clk), .RN(rstn), .Q(memory[914])
         );
  DFFRHQX1 memory_reg_6__1_ ( .D(n1017), .CK(clk), .RN(rstn), .Q(memory[913])
         );
  DFFRHQX1 memory_reg_6__0_ ( .D(n1016), .CK(clk), .RN(rstn), .Q(memory[912])
         );
  DFFRHQX1 memory_reg_10__15_ ( .D(n967), .CK(clk), .RN(rstn), .Q(memory[863])
         );
  DFFRHQX1 memory_reg_10__14_ ( .D(n966), .CK(clk), .RN(rstn), .Q(memory[862])
         );
  DFFRHQX1 memory_reg_10__13_ ( .D(n965), .CK(clk), .RN(rstn), .Q(memory[861])
         );
  DFFRHQX1 memory_reg_10__12_ ( .D(n964), .CK(clk), .RN(rstn), .Q(memory[860])
         );
  DFFRHQX1 memory_reg_10__11_ ( .D(n963), .CK(clk), .RN(rstn), .Q(memory[859])
         );
  DFFRHQX1 memory_reg_10__10_ ( .D(n962), .CK(clk), .RN(rstn), .Q(memory[858])
         );
  DFFRHQX1 memory_reg_10__9_ ( .D(n961), .CK(clk), .RN(rstn), .Q(memory[857])
         );
  DFFRHQX1 memory_reg_10__8_ ( .D(n960), .CK(clk), .RN(rstn), .Q(memory[856])
         );
  DFFRHQX1 memory_reg_10__7_ ( .D(n959), .CK(clk), .RN(rstn), .Q(memory[855])
         );
  DFFRHQX1 memory_reg_10__6_ ( .D(n958), .CK(clk), .RN(rstn), .Q(memory[854])
         );
  DFFRHQX1 memory_reg_10__5_ ( .D(n957), .CK(clk), .RN(rstn), .Q(memory[853])
         );
  DFFRHQX1 memory_reg_10__4_ ( .D(n956), .CK(clk), .RN(rstn), .Q(memory[852])
         );
  DFFRHQX1 memory_reg_10__3_ ( .D(n955), .CK(clk), .RN(rstn), .Q(memory[851])
         );
  DFFRHQX1 memory_reg_10__2_ ( .D(n954), .CK(clk), .RN(rstn), .Q(memory[850])
         );
  DFFRHQX1 memory_reg_10__1_ ( .D(n953), .CK(clk), .RN(rstn), .Q(memory[849])
         );
  DFFRHQX1 memory_reg_10__0_ ( .D(n952), .CK(clk), .RN(rstn), .Q(memory[848])
         );
  DFFRHQX1 memory_reg_14__15_ ( .D(n903), .CK(clk), .RN(rstn), .Q(memory[799])
         );
  DFFRHQX1 memory_reg_14__14_ ( .D(n902), .CK(clk), .RN(rstn), .Q(memory[798])
         );
  DFFRHQX1 memory_reg_14__13_ ( .D(n901), .CK(clk), .RN(rstn), .Q(memory[797])
         );
  DFFRHQX1 memory_reg_14__12_ ( .D(n900), .CK(clk), .RN(rstn), .Q(memory[796])
         );
  DFFRHQX1 memory_reg_14__11_ ( .D(n899), .CK(clk), .RN(rstn), .Q(memory[795])
         );
  DFFRHQX1 memory_reg_14__10_ ( .D(n898), .CK(clk), .RN(rstn), .Q(memory[794])
         );
  DFFRHQX1 memory_reg_14__9_ ( .D(n897), .CK(clk), .RN(rstn), .Q(memory[793])
         );
  DFFRHQX1 memory_reg_14__8_ ( .D(n896), .CK(clk), .RN(rstn), .Q(memory[792])
         );
  DFFRHQX1 memory_reg_14__7_ ( .D(n895), .CK(clk), .RN(rstn), .Q(memory[791])
         );
  DFFRHQX1 memory_reg_14__6_ ( .D(n894), .CK(clk), .RN(rstn), .Q(memory[790])
         );
  DFFRHQX1 memory_reg_14__5_ ( .D(n893), .CK(clk), .RN(rstn), .Q(memory[789])
         );
  DFFRHQX1 memory_reg_14__4_ ( .D(n892), .CK(clk), .RN(rstn), .Q(memory[788])
         );
  DFFRHQX1 memory_reg_14__3_ ( .D(n891), .CK(clk), .RN(rstn), .Q(memory[787])
         );
  DFFRHQX1 memory_reg_14__2_ ( .D(n890), .CK(clk), .RN(rstn), .Q(memory[786])
         );
  DFFRHQX1 memory_reg_14__1_ ( .D(n889), .CK(clk), .RN(rstn), .Q(memory[785])
         );
  DFFRHQX1 memory_reg_14__0_ ( .D(n888), .CK(clk), .RN(rstn), .Q(memory[784])
         );
  DFFRHQX1 memory_reg_18__15_ ( .D(n839), .CK(clk), .RN(rstn), .Q(memory[735])
         );
  DFFRHQX1 memory_reg_18__14_ ( .D(n838), .CK(clk), .RN(rstn), .Q(memory[734])
         );
  DFFRHQX1 memory_reg_18__13_ ( .D(n837), .CK(clk), .RN(rstn), .Q(memory[733])
         );
  DFFRHQX1 memory_reg_18__12_ ( .D(n836), .CK(clk), .RN(rstn), .Q(memory[732])
         );
  DFFRHQX1 memory_reg_18__11_ ( .D(n835), .CK(clk), .RN(rstn), .Q(memory[731])
         );
  DFFRHQX1 memory_reg_18__10_ ( .D(n834), .CK(clk), .RN(rstn), .Q(memory[730])
         );
  DFFRHQX1 memory_reg_18__9_ ( .D(n833), .CK(clk), .RN(rstn), .Q(memory[729])
         );
  DFFRHQX1 memory_reg_18__8_ ( .D(n832), .CK(clk), .RN(rstn), .Q(memory[728])
         );
  DFFRHQX1 memory_reg_18__7_ ( .D(n831), .CK(clk), .RN(rstn), .Q(memory[727])
         );
  DFFRHQX1 memory_reg_18__6_ ( .D(n830), .CK(clk), .RN(rstn), .Q(memory[726])
         );
  DFFRHQX1 memory_reg_18__5_ ( .D(n829), .CK(clk), .RN(rstn), .Q(memory[725])
         );
  DFFRHQX1 memory_reg_18__4_ ( .D(n828), .CK(clk), .RN(rstn), .Q(memory[724])
         );
  DFFRHQX1 memory_reg_18__3_ ( .D(n827), .CK(clk), .RN(rstn), .Q(memory[723])
         );
  DFFRHQX1 memory_reg_18__2_ ( .D(n826), .CK(clk), .RN(rstn), .Q(memory[722])
         );
  DFFRHQX1 memory_reg_18__1_ ( .D(n825), .CK(clk), .RN(rstn), .Q(memory[721])
         );
  DFFRHQX1 memory_reg_18__0_ ( .D(n824), .CK(clk), .RN(rstn), .Q(memory[720])
         );
  DFFRHQX1 memory_reg_22__15_ ( .D(n775), .CK(clk), .RN(rstn), .Q(memory[671])
         );
  DFFRHQX1 memory_reg_22__14_ ( .D(n774), .CK(clk), .RN(rstn), .Q(memory[670])
         );
  DFFRHQX1 memory_reg_22__13_ ( .D(n773), .CK(clk), .RN(rstn), .Q(memory[669])
         );
  DFFRHQX1 memory_reg_22__12_ ( .D(n772), .CK(clk), .RN(rstn), .Q(memory[668])
         );
  DFFRHQX1 memory_reg_22__11_ ( .D(n771), .CK(clk), .RN(rstn), .Q(memory[667])
         );
  DFFRHQX1 memory_reg_22__10_ ( .D(n770), .CK(clk), .RN(rstn), .Q(memory[666])
         );
  DFFRHQX1 memory_reg_22__9_ ( .D(n769), .CK(clk), .RN(rstn), .Q(memory[665])
         );
  DFFRHQX1 memory_reg_22__8_ ( .D(n768), .CK(clk), .RN(rstn), .Q(memory[664])
         );
  DFFRHQX1 memory_reg_22__7_ ( .D(n767), .CK(clk), .RN(rstn), .Q(memory[663])
         );
  DFFRHQX1 memory_reg_22__6_ ( .D(n766), .CK(clk), .RN(rstn), .Q(memory[662])
         );
  DFFRHQX1 memory_reg_22__5_ ( .D(n765), .CK(clk), .RN(rstn), .Q(memory[661])
         );
  DFFRHQX1 memory_reg_22__4_ ( .D(n764), .CK(clk), .RN(rstn), .Q(memory[660])
         );
  DFFRHQX1 memory_reg_22__3_ ( .D(n763), .CK(clk), .RN(rstn), .Q(memory[659])
         );
  DFFRHQX1 memory_reg_22__2_ ( .D(n762), .CK(clk), .RN(rstn), .Q(memory[658])
         );
  DFFRHQX1 memory_reg_22__1_ ( .D(n761), .CK(clk), .RN(rstn), .Q(memory[657])
         );
  DFFRHQX1 memory_reg_22__0_ ( .D(n760), .CK(clk), .RN(rstn), .Q(memory[656])
         );
  DFFRHQX1 memory_reg_26__15_ ( .D(n711), .CK(clk), .RN(rstn), .Q(memory[607])
         );
  DFFRHQX1 memory_reg_26__14_ ( .D(n710), .CK(clk), .RN(rstn), .Q(memory[606])
         );
  DFFRHQX1 memory_reg_26__13_ ( .D(n709), .CK(clk), .RN(rstn), .Q(memory[605])
         );
  DFFRHQX1 memory_reg_26__12_ ( .D(n708), .CK(clk), .RN(rstn), .Q(memory[604])
         );
  DFFRHQX1 memory_reg_26__11_ ( .D(n707), .CK(clk), .RN(rstn), .Q(memory[603])
         );
  DFFRHQX1 memory_reg_26__10_ ( .D(n706), .CK(clk), .RN(rstn), .Q(memory[602])
         );
  DFFRHQX1 memory_reg_26__9_ ( .D(n705), .CK(clk), .RN(rstn), .Q(memory[601])
         );
  DFFRHQX1 memory_reg_26__8_ ( .D(n704), .CK(clk), .RN(rstn), .Q(memory[600])
         );
  DFFRHQX1 memory_reg_26__7_ ( .D(n703), .CK(clk), .RN(rstn), .Q(memory[599])
         );
  DFFRHQX1 memory_reg_26__6_ ( .D(n702), .CK(clk), .RN(rstn), .Q(memory[598])
         );
  DFFRHQX1 memory_reg_26__5_ ( .D(n701), .CK(clk), .RN(rstn), .Q(memory[597])
         );
  DFFRHQX1 memory_reg_26__4_ ( .D(n700), .CK(clk), .RN(rstn), .Q(memory[596])
         );
  DFFRHQX1 memory_reg_26__3_ ( .D(n699), .CK(clk), .RN(rstn), .Q(memory[595])
         );
  DFFRHQX1 memory_reg_26__2_ ( .D(n698), .CK(clk), .RN(rstn), .Q(memory[594])
         );
  DFFRHQX1 memory_reg_26__1_ ( .D(n697), .CK(clk), .RN(rstn), .Q(memory[593])
         );
  DFFRHQX1 memory_reg_26__0_ ( .D(n696), .CK(clk), .RN(rstn), .Q(memory[592])
         );
  DFFRHQX1 memory_reg_30__15_ ( .D(n647), .CK(clk), .RN(rstn), .Q(memory[543])
         );
  DFFRHQX1 memory_reg_30__14_ ( .D(n646), .CK(clk), .RN(rstn), .Q(memory[542])
         );
  DFFRHQX1 memory_reg_30__13_ ( .D(n645), .CK(clk), .RN(rstn), .Q(memory[541])
         );
  DFFRHQX1 memory_reg_30__12_ ( .D(n644), .CK(clk), .RN(rstn), .Q(memory[540])
         );
  DFFRHQX1 memory_reg_30__11_ ( .D(n643), .CK(clk), .RN(rstn), .Q(memory[539])
         );
  DFFRHQX1 memory_reg_30__10_ ( .D(n642), .CK(clk), .RN(rstn), .Q(memory[538])
         );
  DFFRHQX1 memory_reg_30__9_ ( .D(n641), .CK(clk), .RN(rstn), .Q(memory[537])
         );
  DFFRHQX1 memory_reg_30__8_ ( .D(n640), .CK(clk), .RN(rstn), .Q(memory[536])
         );
  DFFRHQX1 memory_reg_30__7_ ( .D(n639), .CK(clk), .RN(rstn), .Q(memory[535])
         );
  DFFRHQX1 memory_reg_30__6_ ( .D(n638), .CK(clk), .RN(rstn), .Q(memory[534])
         );
  DFFRHQX1 memory_reg_30__5_ ( .D(n637), .CK(clk), .RN(rstn), .Q(memory[533])
         );
  DFFRHQX1 memory_reg_30__4_ ( .D(n636), .CK(clk), .RN(rstn), .Q(memory[532])
         );
  DFFRHQX1 memory_reg_30__3_ ( .D(n635), .CK(clk), .RN(rstn), .Q(memory[531])
         );
  DFFRHQX1 memory_reg_30__2_ ( .D(n634), .CK(clk), .RN(rstn), .Q(memory[530])
         );
  DFFRHQX1 memory_reg_30__1_ ( .D(n633), .CK(clk), .RN(rstn), .Q(memory[529])
         );
  DFFRHQX1 memory_reg_30__0_ ( .D(n632), .CK(clk), .RN(rstn), .Q(memory[528])
         );
  DFFRHQX1 memory_reg_34__15_ ( .D(n583), .CK(clk), .RN(rstn), .Q(memory[479])
         );
  DFFRHQX1 memory_reg_34__14_ ( .D(n582), .CK(clk), .RN(rstn), .Q(memory[478])
         );
  DFFRHQX1 memory_reg_34__13_ ( .D(n581), .CK(clk), .RN(rstn), .Q(memory[477])
         );
  DFFRHQX1 memory_reg_34__12_ ( .D(n580), .CK(clk), .RN(rstn), .Q(memory[476])
         );
  DFFRHQX1 memory_reg_34__11_ ( .D(n579), .CK(clk), .RN(rstn), .Q(memory[475])
         );
  DFFRHQX1 memory_reg_34__10_ ( .D(n578), .CK(clk), .RN(rstn), .Q(memory[474])
         );
  DFFRHQX1 memory_reg_34__9_ ( .D(n577), .CK(clk), .RN(rstn), .Q(memory[473])
         );
  DFFRHQX1 memory_reg_34__8_ ( .D(n576), .CK(clk), .RN(rstn), .Q(memory[472])
         );
  DFFRHQX1 memory_reg_34__7_ ( .D(n575), .CK(clk), .RN(rstn), .Q(memory[471])
         );
  DFFRHQX1 memory_reg_34__6_ ( .D(n574), .CK(clk), .RN(rstn), .Q(memory[470])
         );
  DFFRHQX1 memory_reg_34__5_ ( .D(n573), .CK(clk), .RN(rstn), .Q(memory[469])
         );
  DFFRHQX1 memory_reg_34__4_ ( .D(n572), .CK(clk), .RN(rstn), .Q(memory[468])
         );
  DFFRHQX1 memory_reg_34__3_ ( .D(n571), .CK(clk), .RN(rstn), .Q(memory[467])
         );
  DFFRHQX1 memory_reg_34__2_ ( .D(n570), .CK(clk), .RN(rstn), .Q(memory[466])
         );
  DFFRHQX1 memory_reg_34__1_ ( .D(n569), .CK(clk), .RN(rstn), .Q(memory[465])
         );
  DFFRHQX1 memory_reg_34__0_ ( .D(n568), .CK(clk), .RN(rstn), .Q(memory[464])
         );
  DFFRHQX1 memory_reg_38__15_ ( .D(n519), .CK(clk), .RN(rstn), .Q(memory[415])
         );
  DFFRHQX1 memory_reg_38__14_ ( .D(n518), .CK(clk), .RN(rstn), .Q(memory[414])
         );
  DFFRHQX1 memory_reg_38__13_ ( .D(n517), .CK(clk), .RN(rstn), .Q(memory[413])
         );
  DFFRHQX1 memory_reg_38__12_ ( .D(n516), .CK(clk), .RN(rstn), .Q(memory[412])
         );
  DFFRHQX1 memory_reg_38__11_ ( .D(n515), .CK(clk), .RN(rstn), .Q(memory[411])
         );
  DFFRHQX1 memory_reg_38__10_ ( .D(n514), .CK(clk), .RN(rstn), .Q(memory[410])
         );
  DFFRHQX1 memory_reg_38__9_ ( .D(n513), .CK(clk), .RN(rstn), .Q(memory[409])
         );
  DFFRHQX1 memory_reg_38__8_ ( .D(n512), .CK(clk), .RN(rstn), .Q(memory[408])
         );
  DFFRHQX1 memory_reg_38__7_ ( .D(n511), .CK(clk), .RN(rstn), .Q(memory[407])
         );
  DFFRHQX1 memory_reg_38__6_ ( .D(n510), .CK(clk), .RN(rstn), .Q(memory[406])
         );
  DFFRHQX1 memory_reg_38__5_ ( .D(n509), .CK(clk), .RN(rstn), .Q(memory[405])
         );
  DFFRHQX1 memory_reg_38__4_ ( .D(n508), .CK(clk), .RN(rstn), .Q(memory[404])
         );
  DFFRHQX1 memory_reg_38__3_ ( .D(n507), .CK(clk), .RN(rstn), .Q(memory[403])
         );
  DFFRHQX1 memory_reg_38__2_ ( .D(n506), .CK(clk), .RN(rstn), .Q(memory[402])
         );
  DFFRHQX1 memory_reg_38__1_ ( .D(n505), .CK(clk), .RN(rstn), .Q(memory[401])
         );
  DFFRHQX1 memory_reg_38__0_ ( .D(n504), .CK(clk), .RN(rstn), .Q(memory[400])
         );
  DFFRHQX1 memory_reg_42__15_ ( .D(n455), .CK(clk), .RN(rstn), .Q(memory[351])
         );
  DFFRHQX1 memory_reg_42__14_ ( .D(n454), .CK(clk), .RN(rstn), .Q(memory[350])
         );
  DFFRHQX1 memory_reg_42__13_ ( .D(n453), .CK(clk), .RN(rstn), .Q(memory[349])
         );
  DFFRHQX1 memory_reg_42__12_ ( .D(n452), .CK(clk), .RN(rstn), .Q(memory[348])
         );
  DFFRHQX1 memory_reg_42__11_ ( .D(n451), .CK(clk), .RN(rstn), .Q(memory[347])
         );
  DFFRHQX1 memory_reg_42__10_ ( .D(n450), .CK(clk), .RN(rstn), .Q(memory[346])
         );
  DFFRHQX1 memory_reg_42__9_ ( .D(n449), .CK(clk), .RN(rstn), .Q(memory[345])
         );
  DFFRHQX1 memory_reg_42__8_ ( .D(n448), .CK(clk), .RN(rstn), .Q(memory[344])
         );
  DFFRHQX1 memory_reg_42__7_ ( .D(n447), .CK(clk), .RN(rstn), .Q(memory[343])
         );
  DFFRHQX1 memory_reg_42__6_ ( .D(n446), .CK(clk), .RN(rstn), .Q(memory[342])
         );
  DFFRHQX1 memory_reg_42__5_ ( .D(n445), .CK(clk), .RN(rstn), .Q(memory[341])
         );
  DFFRHQX1 memory_reg_42__4_ ( .D(n444), .CK(clk), .RN(rstn), .Q(memory[340])
         );
  DFFRHQX1 memory_reg_42__3_ ( .D(n443), .CK(clk), .RN(rstn), .Q(memory[339])
         );
  DFFRHQX1 memory_reg_42__2_ ( .D(n442), .CK(clk), .RN(rstn), .Q(memory[338])
         );
  DFFRHQX1 memory_reg_42__1_ ( .D(n441), .CK(clk), .RN(rstn), .Q(memory[337])
         );
  DFFRHQX1 memory_reg_42__0_ ( .D(n440), .CK(clk), .RN(rstn), .Q(memory[336])
         );
  DFFRHQX1 memory_reg_46__15_ ( .D(n391), .CK(clk), .RN(rstn), .Q(memory[287])
         );
  DFFRHQX1 memory_reg_46__14_ ( .D(n390), .CK(clk), .RN(rstn), .Q(memory[286])
         );
  DFFRHQX1 memory_reg_46__13_ ( .D(n389), .CK(clk), .RN(rstn), .Q(memory[285])
         );
  DFFRHQX1 memory_reg_46__12_ ( .D(n388), .CK(clk), .RN(rstn), .Q(memory[284])
         );
  DFFRHQX1 memory_reg_46__11_ ( .D(n387), .CK(clk), .RN(rstn), .Q(memory[283])
         );
  DFFRHQX1 memory_reg_46__10_ ( .D(n386), .CK(clk), .RN(rstn), .Q(memory[282])
         );
  DFFRHQX1 memory_reg_46__9_ ( .D(n385), .CK(clk), .RN(rstn), .Q(memory[281])
         );
  DFFRHQX1 memory_reg_46__8_ ( .D(n384), .CK(clk), .RN(rstn), .Q(memory[280])
         );
  DFFRHQX1 memory_reg_46__7_ ( .D(n383), .CK(clk), .RN(rstn), .Q(memory[279])
         );
  DFFRHQX1 memory_reg_46__6_ ( .D(n382), .CK(clk), .RN(rstn), .Q(memory[278])
         );
  DFFRHQX1 memory_reg_46__5_ ( .D(n381), .CK(clk), .RN(rstn), .Q(memory[277])
         );
  DFFRHQX1 memory_reg_46__4_ ( .D(n380), .CK(clk), .RN(rstn), .Q(memory[276])
         );
  DFFRHQX1 memory_reg_46__3_ ( .D(n379), .CK(clk), .RN(rstn), .Q(memory[275])
         );
  DFFRHQX1 memory_reg_46__2_ ( .D(n378), .CK(clk), .RN(rstn), .Q(memory[274])
         );
  DFFRHQX1 memory_reg_46__1_ ( .D(n377), .CK(clk), .RN(rstn), .Q(memory[273])
         );
  DFFRHQX1 memory_reg_46__0_ ( .D(n376), .CK(clk), .RN(rstn), .Q(memory[272])
         );
  DFFRHQX1 memory_reg_50__15_ ( .D(n327), .CK(clk), .RN(rstn), .Q(memory[223])
         );
  DFFRHQX1 memory_reg_50__14_ ( .D(n326), .CK(clk), .RN(rstn), .Q(memory[222])
         );
  DFFRHQX1 memory_reg_50__13_ ( .D(n325), .CK(clk), .RN(rstn), .Q(memory[221])
         );
  DFFRHQX1 memory_reg_50__12_ ( .D(n324), .CK(clk), .RN(rstn), .Q(memory[220])
         );
  DFFRHQX1 memory_reg_50__11_ ( .D(n323), .CK(clk), .RN(rstn), .Q(memory[219])
         );
  DFFRHQX1 memory_reg_50__10_ ( .D(n322), .CK(clk), .RN(rstn), .Q(memory[218])
         );
  DFFRHQX1 memory_reg_50__9_ ( .D(n321), .CK(clk), .RN(rstn), .Q(memory[217])
         );
  DFFRHQX1 memory_reg_50__8_ ( .D(n320), .CK(clk), .RN(rstn), .Q(memory[216])
         );
  DFFRHQX1 memory_reg_50__7_ ( .D(n319), .CK(clk), .RN(rstn), .Q(memory[215])
         );
  DFFRHQX1 memory_reg_50__6_ ( .D(n318), .CK(clk), .RN(rstn), .Q(memory[214])
         );
  DFFRHQX1 memory_reg_50__5_ ( .D(n317), .CK(clk), .RN(rstn), .Q(memory[213])
         );
  DFFRHQX1 memory_reg_50__4_ ( .D(n316), .CK(clk), .RN(rstn), .Q(memory[212])
         );
  DFFRHQX1 memory_reg_50__3_ ( .D(n315), .CK(clk), .RN(rstn), .Q(memory[211])
         );
  DFFRHQX1 memory_reg_50__2_ ( .D(n314), .CK(clk), .RN(rstn), .Q(memory[210])
         );
  DFFRHQX1 memory_reg_50__1_ ( .D(n313), .CK(clk), .RN(rstn), .Q(memory[209])
         );
  DFFRHQX1 memory_reg_50__0_ ( .D(n312), .CK(clk), .RN(rstn), .Q(memory[208])
         );
  DFFRHQX1 memory_reg_54__15_ ( .D(n263), .CK(clk), .RN(rstn), .Q(memory[159])
         );
  DFFRHQX1 memory_reg_54__14_ ( .D(n262), .CK(clk), .RN(rstn), .Q(memory[158])
         );
  DFFRHQX1 memory_reg_54__13_ ( .D(n261), .CK(clk), .RN(rstn), .Q(memory[157])
         );
  DFFRHQX1 memory_reg_54__12_ ( .D(n260), .CK(clk), .RN(rstn), .Q(memory[156])
         );
  DFFRHQX1 memory_reg_54__11_ ( .D(n259), .CK(clk), .RN(rstn), .Q(memory[155])
         );
  DFFRHQX1 memory_reg_54__10_ ( .D(n258), .CK(clk), .RN(rstn), .Q(memory[154])
         );
  DFFRHQX1 memory_reg_54__9_ ( .D(n257), .CK(clk), .RN(rstn), .Q(memory[153])
         );
  DFFRHQX1 memory_reg_54__8_ ( .D(n256), .CK(clk), .RN(rstn), .Q(memory[152])
         );
  DFFRHQX1 memory_reg_54__7_ ( .D(n255), .CK(clk), .RN(rstn), .Q(memory[151])
         );
  DFFRHQX1 memory_reg_54__6_ ( .D(n254), .CK(clk), .RN(rstn), .Q(memory[150])
         );
  DFFRHQX1 memory_reg_54__5_ ( .D(n253), .CK(clk), .RN(rstn), .Q(memory[149])
         );
  DFFRHQX1 memory_reg_54__4_ ( .D(n252), .CK(clk), .RN(rstn), .Q(memory[148])
         );
  DFFRHQX1 memory_reg_54__3_ ( .D(n251), .CK(clk), .RN(rstn), .Q(memory[147])
         );
  DFFRHQX1 memory_reg_54__2_ ( .D(n250), .CK(clk), .RN(rstn), .Q(memory[146])
         );
  DFFRHQX1 memory_reg_54__1_ ( .D(n249), .CK(clk), .RN(rstn), .Q(memory[145])
         );
  DFFRHQX1 memory_reg_54__0_ ( .D(n248), .CK(clk), .RN(rstn), .Q(memory[144])
         );
  DFFRHQX1 memory_reg_58__15_ ( .D(n199), .CK(clk), .RN(rstn), .Q(memory[95])
         );
  DFFRHQX1 memory_reg_58__14_ ( .D(n198), .CK(clk), .RN(rstn), .Q(memory[94])
         );
  DFFRHQX1 memory_reg_58__13_ ( .D(n197), .CK(clk), .RN(rstn), .Q(memory[93])
         );
  DFFRHQX1 memory_reg_58__12_ ( .D(n196), .CK(clk), .RN(rstn), .Q(memory[92])
         );
  DFFRHQX1 memory_reg_58__11_ ( .D(n195), .CK(clk), .RN(rstn), .Q(memory[91])
         );
  DFFRHQX1 memory_reg_58__10_ ( .D(n194), .CK(clk), .RN(rstn), .Q(memory[90])
         );
  DFFRHQX1 memory_reg_58__9_ ( .D(n193), .CK(clk), .RN(rstn), .Q(memory[89])
         );
  DFFRHQX1 memory_reg_58__8_ ( .D(n192), .CK(clk), .RN(rstn), .Q(memory[88])
         );
  DFFRHQX1 memory_reg_58__7_ ( .D(n191), .CK(clk), .RN(rstn), .Q(memory[87])
         );
  DFFRHQX1 memory_reg_58__6_ ( .D(n190), .CK(clk), .RN(rstn), .Q(memory[86])
         );
  DFFRHQX1 memory_reg_58__5_ ( .D(n189), .CK(clk), .RN(rstn), .Q(memory[85])
         );
  DFFRHQX1 memory_reg_58__4_ ( .D(n188), .CK(clk), .RN(rstn), .Q(memory[84])
         );
  DFFRHQX1 memory_reg_58__3_ ( .D(n187), .CK(clk), .RN(rstn), .Q(memory[83])
         );
  DFFRHQX1 memory_reg_58__2_ ( .D(n186), .CK(clk), .RN(rstn), .Q(memory[82])
         );
  DFFRHQX1 memory_reg_58__1_ ( .D(n185), .CK(clk), .RN(rstn), .Q(memory[81])
         );
  DFFRHQX1 memory_reg_58__0_ ( .D(n184), .CK(clk), .RN(rstn), .Q(memory[80])
         );
  DFFRHQX1 memory_reg_62__15_ ( .D(n135), .CK(clk), .RN(rstn), .Q(memory[31])
         );
  DFFRHQX1 memory_reg_62__14_ ( .D(n134), .CK(clk), .RN(rstn), .Q(memory[30])
         );
  DFFRHQX1 memory_reg_62__13_ ( .D(n133), .CK(clk), .RN(rstn), .Q(memory[29])
         );
  DFFRHQX1 memory_reg_62__12_ ( .D(n132), .CK(clk), .RN(rstn), .Q(memory[28])
         );
  DFFRHQX1 memory_reg_62__11_ ( .D(n131), .CK(clk), .RN(rstn), .Q(memory[27])
         );
  DFFRHQX1 memory_reg_62__10_ ( .D(n130), .CK(clk), .RN(rstn), .Q(memory[26])
         );
  DFFRHQX1 memory_reg_62__9_ ( .D(n129), .CK(clk), .RN(rstn), .Q(memory[25])
         );
  DFFRHQX1 memory_reg_62__8_ ( .D(n128), .CK(clk), .RN(rstn), .Q(memory[24])
         );
  DFFRHQX1 memory_reg_62__7_ ( .D(n127), .CK(clk), .RN(rstn), .Q(memory[23])
         );
  DFFRHQX1 memory_reg_62__6_ ( .D(n126), .CK(clk), .RN(rstn), .Q(memory[22])
         );
  DFFRHQX1 memory_reg_62__5_ ( .D(n125), .CK(clk), .RN(rstn), .Q(memory[21])
         );
  DFFRHQX1 memory_reg_62__4_ ( .D(n124), .CK(clk), .RN(rstn), .Q(memory[20])
         );
  DFFRHQX1 memory_reg_62__3_ ( .D(n123), .CK(clk), .RN(rstn), .Q(memory[19])
         );
  DFFRHQX1 memory_reg_62__2_ ( .D(n122), .CK(clk), .RN(rstn), .Q(memory[18])
         );
  DFFRHQX1 memory_reg_62__1_ ( .D(n121), .CK(clk), .RN(rstn), .Q(memory[17])
         );
  DFFRHQX1 memory_reg_62__0_ ( .D(n120), .CK(clk), .RN(rstn), .Q(memory[16])
         );
  INVXL U2 ( .A(addr[2]), .Y(n1509) );
  NAND2X1 U3 ( .A(n23), .B(n24), .Y(n1) );
  NAND2X1 U4 ( .A(n26), .B(n24), .Y(n2) );
  NAND2X1 U5 ( .A(n30), .B(n24), .Y(n3) );
  NAND2X1 U6 ( .A(n34), .B(n24), .Y(n4) );
  NAND2X1 U7 ( .A(n38), .B(n24), .Y(n5) );
  NAND2X1 U8 ( .A(n41), .B(n23), .Y(n6) );
  NAND2X1 U9 ( .A(n41), .B(n26), .Y(n7) );
  NAND2X1 U10 ( .A(n41), .B(n30), .Y(n8) );
  NAND2X1 U11 ( .A(n41), .B(n34), .Y(n9) );
  NAND2X1 U12 ( .A(n41), .B(n38), .Y(n10) );
  NAND2X1 U13 ( .A(n50), .B(n23), .Y(n11) );
  NAND2X1 U14 ( .A(n50), .B(n26), .Y(n12) );
  NAND2X1 U15 ( .A(n50), .B(n30), .Y(n13) );
  NAND2X1 U16 ( .A(n50), .B(n34), .Y(n14) );
  NAND2X1 U17 ( .A(n50), .B(n38), .Y(n15) );
  NAND2X1 U18 ( .A(n59), .B(n23), .Y(n16) );
  NAND2X1 U19 ( .A(n59), .B(n26), .Y(n17) );
  NAND2X1 U20 ( .A(n59), .B(n30), .Y(n18) );
  NAND2X1 U21 ( .A(n59), .B(n34), .Y(n19) );
  NAND2X1 U22 ( .A(n59), .B(n38), .Y(n20) );
  NAND2X1 U23 ( .A(n68), .B(n23), .Y(n21) );
  NAND2X1 U24 ( .A(n68), .B(n26), .Y(n22) );
  NAND2X1 U25 ( .A(n68), .B(n28), .Y(n25) );
  NAND2X1 U26 ( .A(n68), .B(n30), .Y(n27) );
  NAND2X1 U27 ( .A(n68), .B(n32), .Y(n29) );
  NAND2X1 U28 ( .A(n68), .B(n34), .Y(n31) );
  NAND2X1 U29 ( .A(n68), .B(n36), .Y(n33) );
  NAND2X1 U30 ( .A(n68), .B(n38), .Y(n35) );
  NAND2X1 U31 ( .A(n77), .B(n23), .Y(n37) );
  NAND2X1 U32 ( .A(n77), .B(n26), .Y(n40) );
  NAND2X1 U33 ( .A(n77), .B(n28), .Y(n42) );
  NAND2X1 U34 ( .A(n77), .B(n30), .Y(n43) );
  NAND2X1 U35 ( .A(n77), .B(n32), .Y(n44) );
  NAND2X1 U36 ( .A(n77), .B(n34), .Y(n45) );
  NAND2X1 U37 ( .A(n77), .B(n36), .Y(n46) );
  NAND2X1 U38 ( .A(n77), .B(n38), .Y(n47) );
  NAND2X1 U39 ( .A(n86), .B(n23), .Y(n48) );
  NAND2X1 U40 ( .A(n86), .B(n26), .Y(n49) );
  NAND2X1 U41 ( .A(n86), .B(n28), .Y(n51) );
  NAND2X1 U42 ( .A(n86), .B(n30), .Y(n52) );
  NAND2X1 U43 ( .A(n86), .B(n32), .Y(n53) );
  NAND2X1 U44 ( .A(n86), .B(n34), .Y(n54) );
  NAND2X1 U45 ( .A(n86), .B(n36), .Y(n55) );
  NAND2X1 U46 ( .A(n86), .B(n38), .Y(n56) );
  NAND2X1 U47 ( .A(n95), .B(n23), .Y(n57) );
  NAND2X1 U48 ( .A(n95), .B(n26), .Y(n58) );
  NAND2X1 U49 ( .A(n95), .B(n28), .Y(n60) );
  NAND2X1 U50 ( .A(n95), .B(n30), .Y(n61) );
  NAND2X1 U51 ( .A(n95), .B(n32), .Y(n62) );
  NAND2X1 U52 ( .A(n95), .B(n34), .Y(n63) );
  NAND2X1 U53 ( .A(n95), .B(n36), .Y(n64) );
  NAND2X1 U54 ( .A(n95), .B(n38), .Y(n65) );
  NAND2X1 U55 ( .A(n28), .B(n24), .Y(n66) );
  NAND2X1 U56 ( .A(n32), .B(n24), .Y(n67) );
  NAND2X1 U57 ( .A(n36), .B(n24), .Y(n69) );
  NAND2X1 U58 ( .A(n41), .B(n28), .Y(n70) );
  NAND2X1 U59 ( .A(n41), .B(n32), .Y(n71) );
  NAND2X1 U60 ( .A(n41), .B(n36), .Y(n72) );
  NAND2X1 U61 ( .A(n50), .B(n28), .Y(n73) );
  NAND2X1 U62 ( .A(n50), .B(n32), .Y(n74) );
  NAND2X1 U63 ( .A(n50), .B(n36), .Y(n75) );
  NAND2X1 U64 ( .A(n59), .B(n28), .Y(n76) );
  NAND2X1 U65 ( .A(n59), .B(n32), .Y(n78) );
  NAND2X1 U66 ( .A(n59), .B(n36), .Y(n79) );
  NOR4BX1 U67 ( .AN(n39), .B(n1510), .C(addr[4]), .D(n1511), .Y(n86) );
  NOR4BX1 U68 ( .AN(n39), .B(n1429), .C(addr[4]), .D(n1511), .Y(n95) );
  NOR4BX1 U69 ( .AN(n39), .B(n1512), .C(n1510), .D(n1511), .Y(n68) );
  NOR4BX1 U70 ( .AN(n39), .B(n1512), .C(n1430), .D(n1511), .Y(n77) );
  INVX1 U71 ( .A(n1506), .Y(n1452) );
  INVX1 U72 ( .A(n1506), .Y(n1453) );
  INVX1 U73 ( .A(n1506), .Y(n1454) );
  INVX1 U74 ( .A(n1506), .Y(n1455) );
  INVX1 U75 ( .A(n1506), .Y(n1456) );
  INVX1 U76 ( .A(n1506), .Y(n1457) );
  INVX1 U77 ( .A(n1506), .Y(n1458) );
  INVX1 U78 ( .A(n1506), .Y(n1459) );
  INVX1 U79 ( .A(n1506), .Y(n1460) );
  INVX1 U80 ( .A(n1506), .Y(n1461) );
  INVX1 U81 ( .A(n1506), .Y(n1462) );
  INVX1 U82 ( .A(n1506), .Y(n1463) );
  INVX1 U83 ( .A(n1506), .Y(n1464) );
  INVX1 U84 ( .A(n1506), .Y(n1465) );
  INVX1 U85 ( .A(n1506), .Y(n1466) );
  INVX1 U86 ( .A(n1506), .Y(n1467) );
  INVX1 U87 ( .A(n1506), .Y(n1468) );
  INVX1 U88 ( .A(n1506), .Y(n1469) );
  INVX1 U89 ( .A(n1506), .Y(n1470) );
  INVX1 U90 ( .A(n1506), .Y(n1471) );
  INVX1 U91 ( .A(n1434), .Y(n1435) );
  INVX1 U92 ( .A(n1434), .Y(n1436) );
  INVX1 U93 ( .A(n1434), .Y(n1437) );
  INVX1 U94 ( .A(n1434), .Y(n1438) );
  INVX1 U95 ( .A(n1434), .Y(n1439) );
  INVX1 U96 ( .A(n1508), .Y(n1440) );
  INVX1 U97 ( .A(n1433), .Y(n1441) );
  INVX1 U98 ( .A(n1433), .Y(n1442) );
  INVX1 U99 ( .A(n1433), .Y(n1443) );
  INVX1 U100 ( .A(n1434), .Y(n1444) );
  INVX1 U101 ( .A(n1433), .Y(n1445) );
  INVX1 U102 ( .A(n1433), .Y(n1446) );
  INVX1 U103 ( .A(n1434), .Y(n1447) );
  INVX1 U104 ( .A(n1433), .Y(n1448) );
  INVX1 U105 ( .A(n1433), .Y(n1449) );
  INVX1 U106 ( .A(n1433), .Y(n1450) );
  INVX1 U107 ( .A(n1434), .Y(n1451) );
  INVX1 U108 ( .A(n1507), .Y(n1434) );
  INVX1 U109 ( .A(n1507), .Y(n1433) );
  INVX1 U110 ( .A(n1510), .Y(n1427) );
  INVX1 U111 ( .A(n1510), .Y(n1428) );
  INVX1 U112 ( .A(n1510), .Y(n1429) );
  INVX1 U113 ( .A(n1510), .Y(n1430) );
  INVX1 U114 ( .A(n1509), .Y(n1431) );
  INVX1 U115 ( .A(n1509), .Y(n1432) );
  INVX1 U116 ( .A(n1508), .Y(n1507) );
  NOR3X1 U117 ( .A(n1433), .B(n1506), .C(n1509), .Y(n23) );
  NOR3X1 U118 ( .A(n1433), .B(n1455), .C(n1509), .Y(n26) );
  NOR3X1 U119 ( .A(n1506), .B(n1507), .C(n1509), .Y(n28) );
  NOR3X1 U120 ( .A(n1459), .B(n1507), .C(n1509), .Y(n30) );
  NOR3X1 U121 ( .A(n1506), .B(addr[2]), .C(n1508), .Y(n32) );
  NOR3X1 U122 ( .A(n1458), .B(addr[2]), .C(n1508), .Y(n34) );
  NOR3X1 U123 ( .A(n1507), .B(addr[2]), .C(n1506), .Y(n36) );
  NOR3X1 U124 ( .A(n1507), .B(addr[2]), .C(n1454), .Y(n38) );
  INVX1 U125 ( .A(din[0]), .Y(n1505) );
  INVX1 U126 ( .A(din[1]), .Y(n1503) );
  INVX1 U127 ( .A(din[2]), .Y(n1501) );
  INVX1 U128 ( .A(din[3]), .Y(n1499) );
  INVX1 U129 ( .A(din[4]), .Y(n1497) );
  INVX1 U130 ( .A(din[5]), .Y(n1495) );
  INVX1 U131 ( .A(din[6]), .Y(n1493) );
  INVX1 U132 ( .A(din[7]), .Y(n1491) );
  INVX1 U133 ( .A(din[8]), .Y(n1489) );
  INVX1 U134 ( .A(din[9]), .Y(n1487) );
  INVX1 U135 ( .A(din[10]), .Y(n1485) );
  INVX1 U136 ( .A(din[11]), .Y(n1483) );
  INVX1 U137 ( .A(din[12]), .Y(n1481) );
  INVX1 U138 ( .A(din[13]), .Y(n1479) );
  INVX1 U139 ( .A(din[14]), .Y(n1477) );
  INVX1 U140 ( .A(din[15]), .Y(n1475) );
  INVX1 U141 ( .A(din[0]), .Y(n1504) );
  INVX1 U142 ( .A(din[1]), .Y(n1502) );
  INVX1 U143 ( .A(din[2]), .Y(n1500) );
  INVX1 U144 ( .A(din[3]), .Y(n1498) );
  INVX1 U145 ( .A(din[4]), .Y(n1496) );
  INVX1 U146 ( .A(din[5]), .Y(n1494) );
  INVX1 U147 ( .A(din[6]), .Y(n1492) );
  INVX1 U148 ( .A(din[7]), .Y(n1490) );
  INVX1 U149 ( .A(din[8]), .Y(n1488) );
  INVX1 U150 ( .A(din[9]), .Y(n1486) );
  INVX1 U151 ( .A(din[10]), .Y(n1484) );
  INVX1 U152 ( .A(din[11]), .Y(n1482) );
  INVX1 U153 ( .A(din[12]), .Y(n1480) );
  INVX1 U154 ( .A(din[13]), .Y(n1478) );
  INVX1 U155 ( .A(din[14]), .Y(n1476) );
  INVX1 U156 ( .A(din[15]), .Y(n1474) );
  NOR2BX1 U157 ( .AN(N99), .B(n1473), .Y(dout[1]) );
  MX4X1 U158 ( .A(n1146), .B(n1136), .C(n1141), .D(n1131), .S0(n1511), .S1(
        n1472), .Y(N99) );
  MX4X1 U159 ( .A(n1145), .B(n1143), .C(n1144), .D(n1142), .S0(n1427), .S1(
        n1431), .Y(n1146) );
  MX4X1 U160 ( .A(n1135), .B(n1133), .C(n1134), .D(n1132), .S0(n1427), .S1(
        n1431), .Y(n1136) );
  NOR2BX1 U161 ( .AN(N98), .B(n1473), .Y(dout[2]) );
  MX4X1 U162 ( .A(n1166), .B(n1156), .C(n1161), .D(n1151), .S0(n1511), .S1(
        n1472), .Y(N98) );
  MX4X1 U163 ( .A(n1165), .B(n1163), .C(n1164), .D(n1162), .S0(n1427), .S1(
        n1431), .Y(n1166) );
  MX4X1 U164 ( .A(n1155), .B(n1153), .C(n1154), .D(n1152), .S0(n1427), .S1(
        n1431), .Y(n1156) );
  NOR2BX1 U165 ( .AN(N97), .B(n1473), .Y(dout[3]) );
  MX4X1 U166 ( .A(n1186), .B(n1176), .C(n1181), .D(n1171), .S0(n1511), .S1(
        n1472), .Y(N97) );
  MX4X1 U167 ( .A(n1185), .B(n1183), .C(n1184), .D(n1182), .S0(n1427), .S1(
        n1431), .Y(n1186) );
  MX4X1 U168 ( .A(n1175), .B(n1173), .C(n1174), .D(n1172), .S0(n1427), .S1(
        n1431), .Y(n1176) );
  NOR2BX1 U169 ( .AN(N96), .B(n1473), .Y(dout[4]) );
  MX4X1 U170 ( .A(n1206), .B(n1196), .C(n1201), .D(n1191), .S0(addr[5]), .S1(
        n1472), .Y(N96) );
  MX4X1 U171 ( .A(n1205), .B(n1203), .C(n1204), .D(n1202), .S0(n1428), .S1(
        n1432), .Y(n1206) );
  MX4X1 U172 ( .A(n1195), .B(n1193), .C(n1194), .D(n1192), .S0(n1428), .S1(
        n1432), .Y(n1196) );
  NOR2BX1 U173 ( .AN(N95), .B(n1473), .Y(dout[5]) );
  MX4X1 U174 ( .A(n1226), .B(n1216), .C(n1221), .D(n1211), .S0(n1511), .S1(
        n1472), .Y(N95) );
  MX4X1 U175 ( .A(n1225), .B(n1223), .C(n1224), .D(n1222), .S0(n1428), .S1(
        n1432), .Y(n1226) );
  MX4X1 U176 ( .A(n1215), .B(n1213), .C(n1214), .D(n1212), .S0(n1428), .S1(
        n1432), .Y(n1216) );
  NOR2BX1 U177 ( .AN(N94), .B(n1473), .Y(dout[6]) );
  MX4X1 U178 ( .A(n1246), .B(n1236), .C(n1241), .D(n1231), .S0(n1511), .S1(
        n1472), .Y(N94) );
  MX4X1 U179 ( .A(n1245), .B(n1243), .C(n1244), .D(n1242), .S0(n1428), .S1(
        n1432), .Y(n1246) );
  MX4X1 U180 ( .A(n1235), .B(n1233), .C(n1234), .D(n1232), .S0(n1428), .S1(
        n1432), .Y(n1236) );
  NOR2BX1 U181 ( .AN(N93), .B(n1473), .Y(dout[7]) );
  MX4X1 U182 ( .A(n1266), .B(n1256), .C(n1261), .D(n1251), .S0(n1511), .S1(
        n1472), .Y(N93) );
  MX4X1 U183 ( .A(n1265), .B(n1263), .C(n1264), .D(n1262), .S0(n1429), .S1(
        n1431), .Y(n1266) );
  MX4X1 U184 ( .A(n1255), .B(n1253), .C(n1254), .D(n1252), .S0(n1429), .S1(
        n1431), .Y(n1256) );
  NOR2BX1 U185 ( .AN(N92), .B(n1473), .Y(dout[8]) );
  MX4X1 U186 ( .A(n1286), .B(n1276), .C(n1281), .D(n1271), .S0(n1511), .S1(
        n1472), .Y(N92) );
  MX4X1 U187 ( .A(n1285), .B(n1283), .C(n1284), .D(n1282), .S0(n1429), .S1(
        n1432), .Y(n1286) );
  MX4X1 U188 ( .A(n1275), .B(n1273), .C(n1274), .D(n1272), .S0(n1429), .S1(
        n1432), .Y(n1276) );
  NOR2BX1 U189 ( .AN(N91), .B(n1473), .Y(dout[9]) );
  MX4X1 U190 ( .A(n1306), .B(n1296), .C(n1301), .D(n1291), .S0(addr[5]), .S1(
        n1472), .Y(N91) );
  MX4X1 U191 ( .A(n1305), .B(n1303), .C(n1304), .D(n1302), .S0(n1429), .S1(
        n1432), .Y(n1306) );
  MX4X1 U192 ( .A(n1295), .B(n1293), .C(n1294), .D(n1292), .S0(n1429), .S1(
        n1431), .Y(n1296) );
  NOR2BX1 U193 ( .AN(N90), .B(n1473), .Y(dout[10]) );
  MX4X1 U194 ( .A(n1326), .B(n1316), .C(n1321), .D(n1311), .S0(addr[5]), .S1(
        n1472), .Y(N90) );
  MX4X1 U195 ( .A(n1325), .B(n1323), .C(n1324), .D(n1322), .S0(n1430), .S1(
        n1432), .Y(n1326) );
  MX4X1 U196 ( .A(n1315), .B(n1313), .C(n1314), .D(n1312), .S0(n1430), .S1(
        addr[2]), .Y(n1316) );
  NOR2BX1 U197 ( .AN(N89), .B(n1473), .Y(dout[11]) );
  MX4X1 U198 ( .A(n1346), .B(n1336), .C(n1341), .D(n1331), .S0(addr[5]), .S1(
        n1472), .Y(N89) );
  MX4X1 U199 ( .A(n1345), .B(n1343), .C(n1344), .D(n1342), .S0(n1430), .S1(
        n1431), .Y(n1346) );
  MX4X1 U200 ( .A(n1335), .B(n1333), .C(n1334), .D(n1332), .S0(n1430), .S1(
        addr[2]), .Y(n1336) );
  NOR2BX1 U201 ( .AN(N88), .B(n1473), .Y(dout[12]) );
  MX4X1 U202 ( .A(n1366), .B(n1356), .C(n1361), .D(n1351), .S0(addr[5]), .S1(
        n1472), .Y(N88) );
  MX4X1 U203 ( .A(n1365), .B(n1363), .C(n1364), .D(n1362), .S0(n1430), .S1(
        n1432), .Y(n1366) );
  MX4X1 U204 ( .A(n1355), .B(n1353), .C(n1354), .D(n1352), .S0(n1430), .S1(
        n1432), .Y(n1356) );
  NOR2BX1 U205 ( .AN(N87), .B(n1473), .Y(dout[13]) );
  MX4X1 U206 ( .A(n1386), .B(n1376), .C(n1381), .D(n1371), .S0(addr[5]), .S1(
        n1472), .Y(N87) );
  MX4X1 U207 ( .A(n1385), .B(n1383), .C(n1384), .D(n1382), .S0(addr[3]), .S1(
        addr[2]), .Y(n1386) );
  MX4X1 U208 ( .A(n1375), .B(n1373), .C(n1374), .D(n1372), .S0(addr[3]), .S1(
        addr[2]), .Y(n1376) );
  NOR2BX1 U209 ( .AN(N86), .B(n1473), .Y(dout[14]) );
  MX4X1 U210 ( .A(n1406), .B(n1396), .C(n1401), .D(n1391), .S0(addr[5]), .S1(
        n1472), .Y(N86) );
  MX4X1 U211 ( .A(n1405), .B(n1403), .C(n1404), .D(n1402), .S0(addr[3]), .S1(
        addr[2]), .Y(n1406) );
  MX4X1 U212 ( .A(n1395), .B(n1393), .C(n1394), .D(n1392), .S0(addr[3]), .S1(
        addr[2]), .Y(n1396) );
  NOR2BX1 U213 ( .AN(N85), .B(n1473), .Y(dout[15]) );
  MX4X1 U214 ( .A(n1426), .B(n1416), .C(n1421), .D(n1411), .S0(addr[5]), .S1(
        n1472), .Y(N85) );
  MX4X1 U215 ( .A(n1425), .B(n1423), .C(n1424), .D(n1422), .S0(addr[3]), .S1(
        addr[2]), .Y(n1426) );
  MX4X1 U216 ( .A(n1415), .B(n1413), .C(n1414), .D(n1412), .S0(addr[3]), .S1(
        addr[2]), .Y(n1416) );
  NOR2BX1 U217 ( .AN(N100), .B(n1473), .Y(dout[0]) );
  MX4X1 U218 ( .A(n101), .B(n90), .C(n96), .D(n84), .S0(n1511), .S1(n1472), 
        .Y(N100) );
  MX4X1 U219 ( .A(n83), .B(n81), .C(n82), .D(n80), .S0(n1427), .S1(addr[2]), 
        .Y(n84) );
  MX4X1 U220 ( .A(n100), .B(n98), .C(n99), .D(n97), .S0(n1430), .S1(addr[2]), 
        .Y(n101) );
  INVX1 U221 ( .A(addr[0]), .Y(n1506) );
  INVX1 U222 ( .A(addr[1]), .Y(n1508) );
  INVX1 U223 ( .A(addr[3]), .Y(n1510) );
  AND4X2 U224 ( .A(n39), .B(n1511), .C(addr[4]), .D(n1510), .Y(n41) );
  AND4X2 U225 ( .A(n39), .B(n1511), .C(addr[4]), .D(addr[3]), .Y(n24) );
  AND4X2 U226 ( .A(n39), .B(n1511), .C(addr[3]), .D(n1512), .Y(n50) );
  AND4X2 U227 ( .A(n39), .B(n1511), .C(n1510), .D(n1512), .Y(n59) );
  INVX1 U228 ( .A(addr[4]), .Y(n1512) );
  AND2X2 U229 ( .A(wr_rd), .B(en), .Y(n39) );
  BUFX3 U230 ( .A(addr[4]), .Y(n1472) );
  BUFX3 U231 ( .A(n103), .Y(n1473) );
  NAND2BX1 U232 ( .AN(wr_rd), .B(en), .Y(n103) );
  MX4X1 U233 ( .A(memory[944]), .B(memory[928]), .C(memory[912]), .D(
        memory[896]), .S0(n1452), .S1(n1446), .Y(n99) );
  MX4X1 U234 ( .A(memory[176]), .B(memory[160]), .C(memory[144]), .D(
        memory[128]), .S0(n1453), .S1(n1449), .Y(n82) );
  MX4X1 U235 ( .A(memory[433]), .B(memory[417]), .C(memory[401]), .D(
        memory[385]), .S0(n1453), .S1(n1435), .Y(n1134) );
  MX4X1 U236 ( .A(memory[945]), .B(memory[929]), .C(memory[913]), .D(
        memory[897]), .S0(n1454), .S1(n1436), .Y(n1144) );
  MX4X1 U237 ( .A(memory[434]), .B(memory[418]), .C(memory[402]), .D(
        memory[386]), .S0(n1454), .S1(n1436), .Y(n1154) );
  MX4X1 U238 ( .A(memory[946]), .B(memory[930]), .C(memory[914]), .D(
        memory[898]), .S0(n1455), .S1(n1437), .Y(n1164) );
  MX4X1 U239 ( .A(memory[435]), .B(memory[419]), .C(memory[403]), .D(
        memory[387]), .S0(n1456), .S1(n1438), .Y(n1174) );
  MX4X1 U240 ( .A(memory[947]), .B(memory[931]), .C(memory[915]), .D(
        memory[899]), .S0(n1456), .S1(n1438), .Y(n1184) );
  MX4X1 U241 ( .A(memory[436]), .B(memory[420]), .C(memory[404]), .D(
        memory[388]), .S0(n1457), .S1(n1439), .Y(n1194) );
  MX4X1 U242 ( .A(memory[948]), .B(memory[932]), .C(memory[916]), .D(
        memory[900]), .S0(n1458), .S1(n1440), .Y(n1204) );
  MX4X1 U243 ( .A(memory[437]), .B(memory[421]), .C(memory[405]), .D(
        memory[389]), .S0(n1458), .S1(n1440), .Y(n1214) );
  MX4X1 U244 ( .A(memory[949]), .B(memory[933]), .C(memory[917]), .D(
        memory[901]), .S0(n1459), .S1(n1440), .Y(n1224) );
  MX4X1 U245 ( .A(memory[438]), .B(memory[422]), .C(memory[406]), .D(
        memory[390]), .S0(n1460), .S1(n1441), .Y(n1234) );
  MX4X1 U246 ( .A(memory[950]), .B(memory[934]), .C(memory[918]), .D(
        memory[902]), .S0(n1460), .S1(n1441), .Y(n1244) );
  MX4X1 U247 ( .A(memory[439]), .B(memory[423]), .C(memory[407]), .D(
        memory[391]), .S0(n1461), .S1(n1442), .Y(n1254) );
  MX4X1 U248 ( .A(memory[951]), .B(memory[935]), .C(memory[919]), .D(
        memory[903]), .S0(n1462), .S1(n1443), .Y(n1264) );
  MX4X1 U249 ( .A(memory[440]), .B(memory[424]), .C(memory[408]), .D(
        memory[392]), .S0(n1462), .S1(n1443), .Y(n1274) );
  MX4X1 U250 ( .A(memory[952]), .B(memory[936]), .C(memory[920]), .D(
        memory[904]), .S0(n1463), .S1(n1444), .Y(n1284) );
  MX4X1 U251 ( .A(memory[441]), .B(memory[425]), .C(memory[409]), .D(
        memory[393]), .S0(n1464), .S1(n1445), .Y(n1294) );
  MX4X1 U252 ( .A(memory[953]), .B(memory[937]), .C(memory[921]), .D(
        memory[905]), .S0(n1464), .S1(n1445), .Y(n1304) );
  MX4X1 U253 ( .A(memory[442]), .B(memory[426]), .C(memory[410]), .D(
        memory[394]), .S0(n1465), .S1(n1446), .Y(n1314) );
  MX4X1 U254 ( .A(memory[954]), .B(memory[938]), .C(memory[922]), .D(
        memory[906]), .S0(n1466), .S1(n1447), .Y(n1324) );
  MX4X1 U255 ( .A(memory[443]), .B(memory[427]), .C(memory[411]), .D(
        memory[395]), .S0(n1466), .S1(n1447), .Y(n1334) );
  MX4X1 U256 ( .A(memory[955]), .B(memory[939]), .C(memory[923]), .D(
        memory[907]), .S0(n1467), .S1(n1448), .Y(n1344) );
  MX4X1 U257 ( .A(memory[444]), .B(memory[428]), .C(memory[412]), .D(
        memory[396]), .S0(n1468), .S1(n1447), .Y(n1354) );
  MX4X1 U258 ( .A(memory[956]), .B(memory[940]), .C(memory[924]), .D(
        memory[908]), .S0(n1468), .S1(n1441), .Y(n1364) );
  MX4X1 U259 ( .A(memory[445]), .B(memory[429]), .C(memory[413]), .D(
        memory[397]), .S0(n1469), .S1(n1449), .Y(n1374) );
  MX4X1 U260 ( .A(memory[957]), .B(memory[941]), .C(memory[925]), .D(
        memory[909]), .S0(n1470), .S1(n1450), .Y(n1384) );
  MX4X1 U261 ( .A(memory[446]), .B(memory[430]), .C(memory[414]), .D(
        memory[398]), .S0(n1470), .S1(n1450), .Y(n1394) );
  MX4X1 U262 ( .A(memory[958]), .B(memory[942]), .C(memory[926]), .D(
        memory[910]), .S0(n1471), .S1(n1442), .Y(n1404) );
  MX4X1 U263 ( .A(memory[447]), .B(memory[431]), .C(memory[415]), .D(
        memory[399]), .S0(n1468), .S1(n1451), .Y(n1414) );
  MX4X1 U264 ( .A(memory[959]), .B(memory[943]), .C(memory[927]), .D(
        memory[911]), .S0(n1466), .S1(n1451), .Y(n1424) );
  MX4X1 U265 ( .A(n94), .B(n92), .C(n93), .D(n91), .S0(n1428), .S1(addr[2]), 
        .Y(n96) );
  MX4X1 U266 ( .A(memory[752]), .B(memory[736]), .C(memory[720]), .D(
        memory[704]), .S0(n1452), .S1(n1440), .Y(n94) );
  MX4X1 U267 ( .A(memory[624]), .B(memory[608]), .C(memory[592]), .D(
        memory[576]), .S0(n1452), .S1(n1451), .Y(n92) );
  MX4X1 U268 ( .A(memory[688]), .B(memory[672]), .C(memory[656]), .D(
        memory[640]), .S0(n1452), .S1(n1440), .Y(n93) );
  MX4X1 U269 ( .A(n1140), .B(n1138), .C(n1139), .D(n1137), .S0(n1427), .S1(
        n1431), .Y(n1141) );
  MX4X1 U270 ( .A(memory[753]), .B(memory[737]), .C(memory[721]), .D(
        memory[705]), .S0(n1453), .S1(n1435), .Y(n1140) );
  MX4X1 U271 ( .A(memory[625]), .B(memory[609]), .C(memory[593]), .D(
        memory[577]), .S0(n1453), .S1(n1435), .Y(n1138) );
  MX4X1 U272 ( .A(memory[689]), .B(memory[673]), .C(memory[657]), .D(
        memory[641]), .S0(n1453), .S1(n1435), .Y(n1139) );
  MX4X1 U273 ( .A(n1160), .B(n1158), .C(n1159), .D(n1157), .S0(n1427), .S1(
        n1431), .Y(n1161) );
  MX4X1 U274 ( .A(memory[754]), .B(memory[738]), .C(memory[722]), .D(
        memory[706]), .S0(n1455), .S1(n1437), .Y(n1160) );
  MX4X1 U275 ( .A(memory[626]), .B(memory[610]), .C(memory[594]), .D(
        memory[578]), .S0(n1455), .S1(n1437), .Y(n1158) );
  MX4X1 U276 ( .A(memory[690]), .B(memory[674]), .C(memory[658]), .D(
        memory[642]), .S0(n1455), .S1(n1437), .Y(n1159) );
  MX4X1 U277 ( .A(n1180), .B(n1178), .C(n1179), .D(n1177), .S0(n1427), .S1(
        n1431), .Y(n1181) );
  MX4X1 U278 ( .A(memory[755]), .B(memory[739]), .C(memory[723]), .D(
        memory[707]), .S0(n1456), .S1(n1438), .Y(n1180) );
  MX4X1 U279 ( .A(memory[627]), .B(memory[611]), .C(memory[595]), .D(
        memory[579]), .S0(n1456), .S1(n1438), .Y(n1178) );
  MX4X1 U280 ( .A(memory[691]), .B(memory[675]), .C(memory[659]), .D(
        memory[643]), .S0(n1456), .S1(n1438), .Y(n1179) );
  MX4X1 U281 ( .A(n1200), .B(n1198), .C(n1199), .D(n1197), .S0(n1428), .S1(
        n1432), .Y(n1201) );
  MX4X1 U282 ( .A(memory[756]), .B(memory[740]), .C(memory[724]), .D(
        memory[708]), .S0(n1457), .S1(n1439), .Y(n1200) );
  MX4X1 U283 ( .A(memory[628]), .B(memory[612]), .C(memory[596]), .D(
        memory[580]), .S0(n1457), .S1(n1439), .Y(n1198) );
  MX4X1 U284 ( .A(memory[692]), .B(memory[676]), .C(memory[660]), .D(
        memory[644]), .S0(n1457), .S1(n1439), .Y(n1199) );
  MX4X1 U285 ( .A(n1220), .B(n1218), .C(n1219), .D(n1217), .S0(n1428), .S1(
        n1432), .Y(n1221) );
  MX4X1 U286 ( .A(memory[757]), .B(memory[741]), .C(memory[725]), .D(
        memory[709]), .S0(n1459), .S1(n1439), .Y(n1220) );
  MX4X1 U287 ( .A(memory[629]), .B(memory[613]), .C(memory[597]), .D(
        memory[581]), .S0(n1459), .S1(n1440), .Y(n1218) );
  MX4X1 U288 ( .A(memory[693]), .B(memory[677]), .C(memory[661]), .D(
        memory[645]), .S0(n1459), .S1(n1439), .Y(n1219) );
  MX4X1 U289 ( .A(n1240), .B(n1238), .C(n1239), .D(n1237), .S0(n1428), .S1(
        n1432), .Y(n1241) );
  MX4X1 U290 ( .A(memory[758]), .B(memory[742]), .C(memory[726]), .D(
        memory[710]), .S0(n1460), .S1(n1441), .Y(n1240) );
  MX4X1 U291 ( .A(memory[630]), .B(memory[614]), .C(memory[598]), .D(
        memory[582]), .S0(n1460), .S1(n1441), .Y(n1238) );
  MX4X1 U292 ( .A(memory[694]), .B(memory[678]), .C(memory[662]), .D(
        memory[646]), .S0(n1460), .S1(n1441), .Y(n1239) );
  MX4X1 U293 ( .A(n1260), .B(n1258), .C(n1259), .D(n1257), .S0(n1429), .S1(
        n1431), .Y(n1261) );
  MX4X1 U294 ( .A(memory[759]), .B(memory[743]), .C(memory[727]), .D(
        memory[711]), .S0(n1461), .S1(n1442), .Y(n1260) );
  MX4X1 U295 ( .A(memory[631]), .B(memory[615]), .C(memory[599]), .D(
        memory[583]), .S0(n1461), .S1(n1442), .Y(n1258) );
  MX4X1 U296 ( .A(memory[695]), .B(memory[679]), .C(memory[663]), .D(
        memory[647]), .S0(n1461), .S1(n1442), .Y(n1259) );
  MX4X1 U297 ( .A(n1280), .B(n1278), .C(n1279), .D(n1277), .S0(n1429), .S1(
        n1432), .Y(n1281) );
  MX4X1 U298 ( .A(memory[760]), .B(memory[744]), .C(memory[728]), .D(
        memory[712]), .S0(n1463), .S1(n1444), .Y(n1280) );
  MX4X1 U299 ( .A(memory[632]), .B(memory[616]), .C(memory[600]), .D(
        memory[584]), .S0(n1463), .S1(n1444), .Y(n1278) );
  MX4X1 U300 ( .A(memory[696]), .B(memory[680]), .C(memory[664]), .D(
        memory[648]), .S0(n1463), .S1(n1444), .Y(n1279) );
  MX4X1 U301 ( .A(n1300), .B(n1298), .C(n1299), .D(n1297), .S0(n1429), .S1(
        n1431), .Y(n1301) );
  MX4X1 U302 ( .A(memory[761]), .B(memory[745]), .C(memory[729]), .D(
        memory[713]), .S0(n1464), .S1(n1445), .Y(n1300) );
  MX4X1 U303 ( .A(memory[633]), .B(memory[617]), .C(memory[601]), .D(
        memory[585]), .S0(n1464), .S1(n1445), .Y(n1298) );
  MX4X1 U304 ( .A(memory[697]), .B(memory[681]), .C(memory[665]), .D(
        memory[649]), .S0(n1464), .S1(n1445), .Y(n1299) );
  MX4X1 U305 ( .A(n1320), .B(n1318), .C(n1319), .D(n1317), .S0(n1430), .S1(
        addr[2]), .Y(n1321) );
  MX4X1 U306 ( .A(memory[762]), .B(memory[746]), .C(memory[730]), .D(
        memory[714]), .S0(n1465), .S1(n1446), .Y(n1320) );
  MX4X1 U307 ( .A(memory[634]), .B(memory[618]), .C(memory[602]), .D(
        memory[586]), .S0(n1465), .S1(n1446), .Y(n1318) );
  MX4X1 U308 ( .A(memory[698]), .B(memory[682]), .C(memory[666]), .D(
        memory[650]), .S0(n1465), .S1(n1446), .Y(n1319) );
  MX4X1 U309 ( .A(n1340), .B(n1338), .C(n1339), .D(n1337), .S0(n1430), .S1(
        addr[2]), .Y(n1341) );
  MX4X1 U310 ( .A(memory[763]), .B(memory[747]), .C(memory[731]), .D(
        memory[715]), .S0(n1467), .S1(n1448), .Y(n1340) );
  MX4X1 U311 ( .A(memory[635]), .B(memory[619]), .C(memory[603]), .D(
        memory[587]), .S0(n1467), .S1(n1448), .Y(n1338) );
  MX4X1 U312 ( .A(memory[699]), .B(memory[683]), .C(memory[667]), .D(
        memory[651]), .S0(n1467), .S1(n1448), .Y(n1339) );
  MX4X1 U313 ( .A(n1360), .B(n1358), .C(n1359), .D(n1357), .S0(n1430), .S1(
        addr[2]), .Y(n1361) );
  MX4X1 U314 ( .A(memory[764]), .B(memory[748]), .C(memory[732]), .D(
        memory[716]), .S0(n1468), .S1(n1442), .Y(n1360) );
  MX4X1 U315 ( .A(memory[636]), .B(memory[620]), .C(memory[604]), .D(
        memory[588]), .S0(n1468), .S1(n1438), .Y(n1358) );
  MX4X1 U316 ( .A(memory[700]), .B(memory[684]), .C(memory[668]), .D(
        memory[652]), .S0(n1468), .S1(n1444), .Y(n1359) );
  MX4X1 U317 ( .A(n1380), .B(n1378), .C(n1379), .D(n1377), .S0(n1429), .S1(
        n1431), .Y(n1381) );
  MX4X1 U318 ( .A(memory[765]), .B(memory[749]), .C(memory[733]), .D(
        memory[717]), .S0(n1469), .S1(n1449), .Y(n1380) );
  MX4X1 U319 ( .A(memory[637]), .B(memory[621]), .C(memory[605]), .D(
        memory[589]), .S0(n1469), .S1(n1449), .Y(n1378) );
  MX4X1 U320 ( .A(memory[701]), .B(memory[685]), .C(memory[669]), .D(
        memory[653]), .S0(n1469), .S1(n1449), .Y(n1379) );
  MX4X1 U321 ( .A(n1400), .B(n1398), .C(n1399), .D(n1397), .S0(n1428), .S1(
        n1432), .Y(n1401) );
  MX4X1 U322 ( .A(memory[766]), .B(memory[750]), .C(memory[734]), .D(
        memory[718]), .S0(n1471), .S1(n1441), .Y(n1400) );
  MX4X1 U323 ( .A(memory[638]), .B(memory[622]), .C(memory[606]), .D(
        memory[590]), .S0(n1471), .S1(n1438), .Y(n1398) );
  MX4X1 U324 ( .A(memory[702]), .B(memory[686]), .C(memory[670]), .D(
        memory[654]), .S0(n1471), .S1(n1444), .Y(n1399) );
  MX4X1 U325 ( .A(n1420), .B(n1418), .C(n1419), .D(n1417), .S0(n1427), .S1(
        addr[2]), .Y(n1421) );
  MX4X1 U326 ( .A(memory[767]), .B(memory[751]), .C(memory[735]), .D(
        memory[719]), .S0(n1471), .S1(n1451), .Y(n1420) );
  MX4X1 U327 ( .A(memory[639]), .B(memory[623]), .C(memory[607]), .D(
        memory[591]), .S0(n1463), .S1(n1451), .Y(n1418) );
  MX4X1 U328 ( .A(memory[703]), .B(memory[687]), .C(memory[671]), .D(
        memory[655]), .S0(n1461), .S1(n1451), .Y(n1419) );
  MX4X1 U329 ( .A(memory[1008]), .B(memory[992]), .C(memory[976]), .D(
        memory[960]), .S0(n1452), .S1(n1451), .Y(n100) );
  MX4X1 U330 ( .A(memory[240]), .B(memory[224]), .C(memory[208]), .D(
        memory[192]), .S0(n1456), .S1(n1437), .Y(n83) );
  MX4X1 U331 ( .A(memory[497]), .B(memory[481]), .C(memory[465]), .D(
        memory[449]), .S0(n1453), .S1(n1435), .Y(n1135) );
  MX4X1 U332 ( .A(memory[1009]), .B(memory[993]), .C(memory[977]), .D(
        memory[961]), .S0(n1454), .S1(n1436), .Y(n1145) );
  MX4X1 U333 ( .A(memory[498]), .B(memory[482]), .C(memory[466]), .D(
        memory[450]), .S0(n1454), .S1(n1436), .Y(n1155) );
  MX4X1 U334 ( .A(memory[1010]), .B(memory[994]), .C(memory[978]), .D(
        memory[962]), .S0(n1455), .S1(n1437), .Y(n1165) );
  MX4X1 U335 ( .A(memory[499]), .B(memory[483]), .C(memory[467]), .D(
        memory[451]), .S0(n1456), .S1(n1438), .Y(n1175) );
  MX4X1 U336 ( .A(memory[1011]), .B(memory[995]), .C(memory[979]), .D(
        memory[963]), .S0(n1456), .S1(n1438), .Y(n1185) );
  MX4X1 U337 ( .A(memory[500]), .B(memory[484]), .C(memory[468]), .D(
        memory[452]), .S0(n1457), .S1(n1439), .Y(n1195) );
  MX4X1 U338 ( .A(memory[1012]), .B(memory[996]), .C(memory[980]), .D(
        memory[964]), .S0(n1458), .S1(n1440), .Y(n1205) );
  MX4X1 U339 ( .A(memory[501]), .B(memory[485]), .C(memory[469]), .D(
        memory[453]), .S0(n1458), .S1(n1440), .Y(n1215) );
  MX4X1 U340 ( .A(memory[1013]), .B(memory[997]), .C(memory[981]), .D(
        memory[965]), .S0(n1459), .S1(n1451), .Y(n1225) );
  MX4X1 U341 ( .A(memory[502]), .B(memory[486]), .C(memory[470]), .D(
        memory[454]), .S0(n1460), .S1(n1441), .Y(n1235) );
  MX4X1 U342 ( .A(memory[1014]), .B(memory[998]), .C(memory[982]), .D(
        memory[966]), .S0(n1460), .S1(n1441), .Y(n1245) );
  MX4X1 U343 ( .A(memory[503]), .B(memory[487]), .C(memory[471]), .D(
        memory[455]), .S0(n1461), .S1(n1442), .Y(n1255) );
  MX4X1 U344 ( .A(memory[1015]), .B(memory[999]), .C(memory[983]), .D(
        memory[967]), .S0(n1462), .S1(n1443), .Y(n1265) );
  MX4X1 U345 ( .A(memory[504]), .B(memory[488]), .C(memory[472]), .D(
        memory[456]), .S0(n1462), .S1(n1443), .Y(n1275) );
  MX4X1 U346 ( .A(memory[1016]), .B(memory[1000]), .C(memory[984]), .D(
        memory[968]), .S0(n1463), .S1(n1444), .Y(n1285) );
  MX4X1 U347 ( .A(memory[505]), .B(memory[489]), .C(memory[473]), .D(
        memory[457]), .S0(n1464), .S1(n1445), .Y(n1295) );
  MX4X1 U348 ( .A(memory[1017]), .B(memory[1001]), .C(memory[985]), .D(
        memory[969]), .S0(n1464), .S1(n1445), .Y(n1305) );
  MX4X1 U349 ( .A(memory[506]), .B(memory[490]), .C(memory[474]), .D(
        memory[458]), .S0(n1465), .S1(n1446), .Y(n1315) );
  MX4X1 U350 ( .A(memory[1018]), .B(memory[1002]), .C(memory[986]), .D(
        memory[970]), .S0(n1466), .S1(n1447), .Y(n1325) );
  MX4X1 U351 ( .A(memory[507]), .B(memory[491]), .C(memory[475]), .D(
        memory[459]), .S0(n1466), .S1(n1447), .Y(n1335) );
  MX4X1 U352 ( .A(memory[1019]), .B(memory[1003]), .C(memory[987]), .D(
        memory[971]), .S0(n1467), .S1(n1448), .Y(n1345) );
  MX4X1 U353 ( .A(memory[508]), .B(memory[492]), .C(memory[476]), .D(
        memory[460]), .S0(n1468), .S1(n1446), .Y(n1355) );
  MX4X1 U354 ( .A(memory[1020]), .B(memory[1004]), .C(memory[988]), .D(
        memory[972]), .S0(n1468), .S1(n1448), .Y(n1365) );
  MX4X1 U355 ( .A(memory[509]), .B(memory[493]), .C(memory[477]), .D(
        memory[461]), .S0(n1469), .S1(n1449), .Y(n1375) );
  MX4X1 U356 ( .A(memory[1021]), .B(memory[1005]), .C(memory[989]), .D(
        memory[973]), .S0(n1470), .S1(n1450), .Y(n1385) );
  MX4X1 U357 ( .A(memory[510]), .B(memory[494]), .C(memory[478]), .D(
        memory[462]), .S0(n1470), .S1(n1450), .Y(n1395) );
  MX4X1 U358 ( .A(memory[1022]), .B(memory[1006]), .C(memory[990]), .D(
        memory[974]), .S0(n1471), .S1(n1436), .Y(n1405) );
  MX4X1 U359 ( .A(memory[511]), .B(memory[495]), .C(memory[479]), .D(
        memory[463]), .S0(n1465), .S1(n1451), .Y(n1415) );
  MX4X1 U360 ( .A(memory[1023]), .B(memory[1007]), .C(memory[991]), .D(
        memory[975]), .S0(n1470), .S1(n1451), .Y(n1425) );
  MX4X1 U361 ( .A(memory[560]), .B(memory[544]), .C(memory[528]), .D(
        memory[512]), .S0(n1452), .S1(n1440), .Y(n91) );
  MX4X1 U362 ( .A(memory[304]), .B(memory[288]), .C(memory[272]), .D(
        memory[256]), .S0(n1452), .S1(n1440), .Y(n85) );
  MX4X1 U363 ( .A(memory[816]), .B(memory[800]), .C(memory[784]), .D(
        memory[768]), .S0(n1452), .S1(n1440), .Y(n97) );
  MX4X1 U364 ( .A(memory[48]), .B(memory[32]), .C(memory[16]), .D(memory[0]), 
        .S0(n1452), .S1(n1440), .Y(n80) );
  MX4X1 U365 ( .A(memory[49]), .B(memory[33]), .C(memory[17]), .D(memory[1]), 
        .S0(n1453), .S1(n1435), .Y(n102) );
  MX4X1 U366 ( .A(memory[561]), .B(memory[545]), .C(memory[529]), .D(
        memory[513]), .S0(n1453), .S1(n1435), .Y(n1137) );
  MX4X1 U367 ( .A(memory[305]), .B(memory[289]), .C(memory[273]), .D(
        memory[257]), .S0(n1453), .S1(n1435), .Y(n1132) );
  MX4X1 U368 ( .A(memory[817]), .B(memory[801]), .C(memory[785]), .D(
        memory[769]), .S0(n1454), .S1(n1436), .Y(n1142) );
  MX4X1 U369 ( .A(memory[50]), .B(memory[34]), .C(memory[18]), .D(memory[2]), 
        .S0(n1454), .S1(n1436), .Y(n1147) );
  MX4X1 U370 ( .A(memory[562]), .B(memory[546]), .C(memory[530]), .D(
        memory[514]), .S0(n1455), .S1(n1437), .Y(n1157) );
  MX4X1 U371 ( .A(memory[306]), .B(memory[290]), .C(memory[274]), .D(
        memory[258]), .S0(n1454), .S1(n1436), .Y(n1152) );
  MX4X1 U372 ( .A(memory[818]), .B(memory[802]), .C(memory[786]), .D(
        memory[770]), .S0(n1455), .S1(n1437), .Y(n1162) );
  MX4X1 U373 ( .A(memory[51]), .B(memory[35]), .C(memory[19]), .D(memory[3]), 
        .S0(n1455), .S1(n1437), .Y(n1167) );
  MX4X1 U374 ( .A(memory[563]), .B(memory[547]), .C(memory[531]), .D(
        memory[515]), .S0(n1456), .S1(n1438), .Y(n1177) );
  MX4X1 U375 ( .A(memory[307]), .B(memory[291]), .C(memory[275]), .D(
        memory[259]), .S0(n1456), .S1(n1438), .Y(n1172) );
  MX4X1 U376 ( .A(memory[819]), .B(memory[803]), .C(memory[787]), .D(
        memory[771]), .S0(n1456), .S1(n1438), .Y(n1182) );
  MX4X1 U377 ( .A(memory[52]), .B(memory[36]), .C(memory[20]), .D(memory[4]), 
        .S0(n1457), .S1(n1439), .Y(n1187) );
  MX4X1 U378 ( .A(memory[564]), .B(memory[548]), .C(memory[532]), .D(
        memory[516]), .S0(n1457), .S1(n1439), .Y(n1197) );
  MX4X1 U379 ( .A(memory[308]), .B(memory[292]), .C(memory[276]), .D(
        memory[260]), .S0(n1457), .S1(n1439), .Y(n1192) );
  MX4X1 U380 ( .A(memory[820]), .B(memory[804]), .C(memory[788]), .D(
        memory[772]), .S0(n1458), .S1(n1440), .Y(n1202) );
  MX4X1 U381 ( .A(memory[53]), .B(memory[37]), .C(memory[21]), .D(memory[5]), 
        .S0(n1458), .S1(n1440), .Y(n1207) );
  MX4X1 U382 ( .A(memory[565]), .B(memory[549]), .C(memory[533]), .D(
        memory[517]), .S0(n1459), .S1(n1440), .Y(n1217) );
  MX4X1 U383 ( .A(memory[309]), .B(memory[293]), .C(memory[277]), .D(
        memory[261]), .S0(n1458), .S1(n1440), .Y(n1212) );
  MX4X1 U384 ( .A(memory[821]), .B(memory[805]), .C(memory[789]), .D(
        memory[773]), .S0(n1459), .S1(n1440), .Y(n1222) );
  MX4X1 U385 ( .A(memory[54]), .B(memory[38]), .C(memory[22]), .D(memory[6]), 
        .S0(n1459), .S1(n1440), .Y(n1227) );
  MX4X1 U386 ( .A(memory[566]), .B(memory[550]), .C(memory[534]), .D(
        memory[518]), .S0(n1460), .S1(n1441), .Y(n1237) );
  MX4X1 U387 ( .A(memory[310]), .B(memory[294]), .C(memory[278]), .D(
        memory[262]), .S0(n1460), .S1(n1441), .Y(n1232) );
  MX4X1 U388 ( .A(memory[822]), .B(memory[806]), .C(memory[790]), .D(
        memory[774]), .S0(n1460), .S1(n1441), .Y(n1242) );
  MX4X1 U389 ( .A(memory[55]), .B(memory[39]), .C(memory[23]), .D(memory[7]), 
        .S0(n1461), .S1(n1442), .Y(n1247) );
  MX4X1 U390 ( .A(memory[567]), .B(memory[551]), .C(memory[535]), .D(
        memory[519]), .S0(n1461), .S1(n1442), .Y(n1257) );
  MX4X1 U391 ( .A(memory[311]), .B(memory[295]), .C(memory[279]), .D(
        memory[263]), .S0(n1461), .S1(n1442), .Y(n1252) );
  MX4X1 U392 ( .A(memory[823]), .B(memory[807]), .C(memory[791]), .D(
        memory[775]), .S0(n1462), .S1(n1443), .Y(n1262) );
  MX4X1 U393 ( .A(memory[56]), .B(memory[40]), .C(memory[24]), .D(memory[8]), 
        .S0(n1462), .S1(n1443), .Y(n1267) );
  MX4X1 U394 ( .A(memory[568]), .B(memory[552]), .C(memory[536]), .D(
        memory[520]), .S0(n1463), .S1(n1444), .Y(n1277) );
  MX4X1 U395 ( .A(memory[312]), .B(memory[296]), .C(memory[280]), .D(
        memory[264]), .S0(n1462), .S1(n1443), .Y(n1272) );
  MX4X1 U396 ( .A(memory[824]), .B(memory[808]), .C(memory[792]), .D(
        memory[776]), .S0(n1463), .S1(n1444), .Y(n1282) );
  MX4X1 U397 ( .A(memory[57]), .B(memory[41]), .C(memory[25]), .D(memory[9]), 
        .S0(n1463), .S1(n1444), .Y(n1287) );
  MX4X1 U398 ( .A(memory[569]), .B(memory[553]), .C(memory[537]), .D(
        memory[521]), .S0(n1464), .S1(n1445), .Y(n1297) );
  MX4X1 U399 ( .A(memory[313]), .B(memory[297]), .C(memory[281]), .D(
        memory[265]), .S0(n1464), .S1(n1445), .Y(n1292) );
  MX4X1 U400 ( .A(memory[825]), .B(memory[809]), .C(memory[793]), .D(
        memory[777]), .S0(n1464), .S1(n1445), .Y(n1302) );
  MX4X1 U401 ( .A(memory[58]), .B(memory[42]), .C(memory[26]), .D(memory[10]), 
        .S0(n1465), .S1(n1446), .Y(n1307) );
  MX4X1 U402 ( .A(memory[570]), .B(memory[554]), .C(memory[538]), .D(
        memory[522]), .S0(n1465), .S1(n1446), .Y(n1317) );
  MX4X1 U403 ( .A(memory[314]), .B(memory[298]), .C(memory[282]), .D(
        memory[266]), .S0(n1465), .S1(n1446), .Y(n1312) );
  MX4X1 U404 ( .A(memory[826]), .B(memory[810]), .C(memory[794]), .D(
        memory[778]), .S0(n1466), .S1(n1447), .Y(n1322) );
  MX4X1 U405 ( .A(memory[59]), .B(memory[43]), .C(memory[27]), .D(memory[11]), 
        .S0(n1466), .S1(n1447), .Y(n1327) );
  MX4X1 U406 ( .A(memory[571]), .B(memory[555]), .C(memory[539]), .D(
        memory[523]), .S0(n1467), .S1(n1448), .Y(n1337) );
  MX4X1 U407 ( .A(memory[315]), .B(memory[299]), .C(memory[283]), .D(
        memory[267]), .S0(n1466), .S1(n1447), .Y(n1332) );
  MX4X1 U408 ( .A(memory[827]), .B(memory[811]), .C(memory[795]), .D(
        memory[779]), .S0(n1467), .S1(n1448), .Y(n1342) );
  MX4X1 U409 ( .A(memory[60]), .B(memory[44]), .C(memory[28]), .D(memory[12]), 
        .S0(n1467), .S1(n1448), .Y(n1347) );
  MX4X1 U410 ( .A(memory[572]), .B(memory[556]), .C(memory[540]), .D(
        memory[524]), .S0(n1468), .S1(n1435), .Y(n1357) );
  MX4X1 U411 ( .A(memory[316]), .B(memory[300]), .C(memory[284]), .D(
        memory[268]), .S0(n1468), .S1(n1436), .Y(n1352) );
  MX4X1 U412 ( .A(memory[828]), .B(memory[812]), .C(memory[796]), .D(
        memory[780]), .S0(n1468), .S1(n1437), .Y(n1362) );
  MX4X1 U413 ( .A(memory[61]), .B(memory[45]), .C(memory[29]), .D(memory[13]), 
        .S0(n1469), .S1(n1449), .Y(n1367) );
  MX4X1 U414 ( .A(memory[573]), .B(memory[557]), .C(memory[541]), .D(
        memory[525]), .S0(n1469), .S1(n1449), .Y(n1377) );
  MX4X1 U415 ( .A(memory[317]), .B(memory[301]), .C(memory[285]), .D(
        memory[269]), .S0(n1469), .S1(n1449), .Y(n1372) );
  MX4X1 U416 ( .A(memory[829]), .B(memory[813]), .C(memory[797]), .D(
        memory[781]), .S0(n1470), .S1(n1450), .Y(n1382) );
  MX4X1 U417 ( .A(memory[62]), .B(memory[46]), .C(memory[30]), .D(memory[14]), 
        .S0(n1470), .S1(n1450), .Y(n1387) );
  MX4X1 U418 ( .A(memory[574]), .B(memory[558]), .C(memory[542]), .D(
        memory[526]), .S0(n1471), .S1(n1435), .Y(n1397) );
  MX4X1 U419 ( .A(memory[318]), .B(memory[302]), .C(memory[286]), .D(
        memory[270]), .S0(n1470), .S1(n1450), .Y(n1392) );
  MX4X1 U420 ( .A(memory[830]), .B(memory[814]), .C(memory[798]), .D(
        memory[782]), .S0(n1471), .S1(n1447), .Y(n1402) );
  MX4X1 U421 ( .A(memory[63]), .B(memory[47]), .C(memory[31]), .D(memory[15]), 
        .S0(n1471), .S1(n1436), .Y(n1407) );
  MX4X1 U422 ( .A(memory[575]), .B(memory[559]), .C(memory[543]), .D(
        memory[527]), .S0(n1464), .S1(n1451), .Y(n1417) );
  MX4X1 U423 ( .A(memory[319]), .B(memory[303]), .C(memory[287]), .D(
        memory[271]), .S0(n1462), .S1(n1451), .Y(n1412) );
  MX4X1 U424 ( .A(memory[831]), .B(memory[815]), .C(memory[799]), .D(
        memory[783]), .S0(n1457), .S1(n1451), .Y(n1422) );
  MX4X1 U425 ( .A(n1130), .B(n1128), .C(n1129), .D(n102), .S0(n1427), .S1(
        n1431), .Y(n1131) );
  MX4X1 U426 ( .A(memory[241]), .B(memory[225]), .C(memory[209]), .D(
        memory[193]), .S0(n1453), .S1(n1435), .Y(n1130) );
  MX4X1 U427 ( .A(memory[113]), .B(memory[97]), .C(memory[81]), .D(memory[65]), 
        .S0(n1453), .S1(n1435), .Y(n1128) );
  MX4X1 U428 ( .A(memory[177]), .B(memory[161]), .C(memory[145]), .D(
        memory[129]), .S0(n1453), .S1(n1435), .Y(n1129) );
  MX4X1 U429 ( .A(n1150), .B(n1148), .C(n1149), .D(n1147), .S0(n1427), .S1(
        n1431), .Y(n1151) );
  MX4X1 U430 ( .A(memory[242]), .B(memory[226]), .C(memory[210]), .D(
        memory[194]), .S0(n1454), .S1(n1436), .Y(n1150) );
  MX4X1 U431 ( .A(memory[114]), .B(memory[98]), .C(memory[82]), .D(memory[66]), 
        .S0(n1454), .S1(n1436), .Y(n1148) );
  MX4X1 U432 ( .A(memory[178]), .B(memory[162]), .C(memory[146]), .D(
        memory[130]), .S0(n1454), .S1(n1436), .Y(n1149) );
  MX4X1 U433 ( .A(n1170), .B(n1168), .C(n1169), .D(n1167), .S0(n1427), .S1(
        n1431), .Y(n1171) );
  MX4X1 U434 ( .A(memory[243]), .B(memory[227]), .C(memory[211]), .D(
        memory[195]), .S0(n1455), .S1(n1437), .Y(n1170) );
  MX4X1 U435 ( .A(memory[115]), .B(memory[99]), .C(memory[83]), .D(memory[67]), 
        .S0(n1455), .S1(n1437), .Y(n1168) );
  MX4X1 U436 ( .A(memory[179]), .B(memory[163]), .C(memory[147]), .D(
        memory[131]), .S0(n1455), .S1(n1437), .Y(n1169) );
  MX4X1 U437 ( .A(n1190), .B(n1188), .C(n1189), .D(n1187), .S0(n1428), .S1(
        n1432), .Y(n1191) );
  MX4X1 U438 ( .A(memory[244]), .B(memory[228]), .C(memory[212]), .D(
        memory[196]), .S0(n1457), .S1(n1439), .Y(n1190) );
  MX4X1 U439 ( .A(memory[116]), .B(memory[100]), .C(memory[84]), .D(memory[68]), .S0(n1457), .S1(n1439), .Y(n1188) );
  MX4X1 U440 ( .A(memory[180]), .B(memory[164]), .C(memory[148]), .D(
        memory[132]), .S0(n1457), .S1(n1439), .Y(n1189) );
  MX4X1 U441 ( .A(n1210), .B(n1208), .C(n1209), .D(n1207), .S0(n1428), .S1(
        n1432), .Y(n1211) );
  MX4X1 U442 ( .A(memory[245]), .B(memory[229]), .C(memory[213]), .D(
        memory[197]), .S0(n1458), .S1(n1440), .Y(n1210) );
  MX4X1 U443 ( .A(memory[117]), .B(memory[101]), .C(memory[85]), .D(memory[69]), .S0(n1458), .S1(n1440), .Y(n1208) );
  MX4X1 U444 ( .A(memory[181]), .B(memory[165]), .C(memory[149]), .D(
        memory[133]), .S0(n1458), .S1(n1440), .Y(n1209) );
  MX4X1 U445 ( .A(n1230), .B(n1228), .C(n1229), .D(n1227), .S0(n1428), .S1(
        n1432), .Y(n1231) );
  MX4X1 U446 ( .A(memory[246]), .B(memory[230]), .C(memory[214]), .D(
        memory[198]), .S0(n1459), .S1(n1439), .Y(n1230) );
  MX4X1 U447 ( .A(memory[118]), .B(memory[102]), .C(memory[86]), .D(memory[70]), .S0(n1459), .S1(n1440), .Y(n1228) );
  MX4X1 U448 ( .A(memory[182]), .B(memory[166]), .C(memory[150]), .D(
        memory[134]), .S0(n1459), .S1(n1439), .Y(n1229) );
  MX4X1 U449 ( .A(n1250), .B(n1248), .C(n1249), .D(n1247), .S0(n1429), .S1(
        n1431), .Y(n1251) );
  MX4X1 U450 ( .A(memory[247]), .B(memory[231]), .C(memory[215]), .D(
        memory[199]), .S0(n1461), .S1(n1442), .Y(n1250) );
  MX4X1 U451 ( .A(memory[119]), .B(memory[103]), .C(memory[87]), .D(memory[71]), .S0(n1461), .S1(n1442), .Y(n1248) );
  MX4X1 U452 ( .A(memory[183]), .B(memory[167]), .C(memory[151]), .D(
        memory[135]), .S0(n1461), .S1(n1442), .Y(n1249) );
  MX4X1 U453 ( .A(n1270), .B(n1268), .C(n1269), .D(n1267), .S0(n1429), .S1(
        n1432), .Y(n1271) );
  MX4X1 U454 ( .A(memory[248]), .B(memory[232]), .C(memory[216]), .D(
        memory[200]), .S0(n1462), .S1(n1443), .Y(n1270) );
  MX4X1 U455 ( .A(memory[120]), .B(memory[104]), .C(memory[88]), .D(memory[72]), .S0(n1462), .S1(n1443), .Y(n1268) );
  MX4X1 U456 ( .A(memory[184]), .B(memory[168]), .C(memory[152]), .D(
        memory[136]), .S0(n1462), .S1(n1443), .Y(n1269) );
  MX4X1 U457 ( .A(n1290), .B(n1288), .C(n1289), .D(n1287), .S0(n1429), .S1(
        n1432), .Y(n1291) );
  MX4X1 U458 ( .A(memory[249]), .B(memory[233]), .C(memory[217]), .D(
        memory[201]), .S0(n1463), .S1(n1444), .Y(n1290) );
  MX4X1 U459 ( .A(memory[121]), .B(memory[105]), .C(memory[89]), .D(memory[73]), .S0(n1463), .S1(n1444), .Y(n1288) );
  MX4X1 U460 ( .A(memory[185]), .B(memory[169]), .C(memory[153]), .D(
        memory[137]), .S0(n1463), .S1(n1444), .Y(n1289) );
  MX4X1 U461 ( .A(n1310), .B(n1308), .C(n1309), .D(n1307), .S0(n1430), .S1(
        n1432), .Y(n1311) );
  MX4X1 U462 ( .A(memory[250]), .B(memory[234]), .C(memory[218]), .D(
        memory[202]), .S0(n1465), .S1(n1446), .Y(n1310) );
  MX4X1 U463 ( .A(memory[122]), .B(memory[106]), .C(memory[90]), .D(memory[74]), .S0(n1465), .S1(n1446), .Y(n1308) );
  MX4X1 U464 ( .A(memory[186]), .B(memory[170]), .C(memory[154]), .D(
        memory[138]), .S0(n1465), .S1(n1446), .Y(n1309) );
  MX4X1 U465 ( .A(n1330), .B(n1328), .C(n1329), .D(n1327), .S0(n1430), .S1(
        n1431), .Y(n1331) );
  MX4X1 U466 ( .A(memory[251]), .B(memory[235]), .C(memory[219]), .D(
        memory[203]), .S0(n1466), .S1(n1447), .Y(n1330) );
  MX4X1 U467 ( .A(memory[123]), .B(memory[107]), .C(memory[91]), .D(memory[75]), .S0(n1466), .S1(n1447), .Y(n1328) );
  MX4X1 U468 ( .A(memory[187]), .B(memory[171]), .C(memory[155]), .D(
        memory[139]), .S0(n1466), .S1(n1447), .Y(n1329) );
  MX4X1 U469 ( .A(n1350), .B(n1348), .C(n1349), .D(n1347), .S0(n1430), .S1(
        addr[2]), .Y(n1351) );
  MX4X1 U470 ( .A(memory[252]), .B(memory[236]), .C(memory[220]), .D(
        memory[204]), .S0(n1467), .S1(n1448), .Y(n1350) );
  MX4X1 U471 ( .A(memory[124]), .B(memory[108]), .C(memory[92]), .D(memory[76]), .S0(n1467), .S1(n1448), .Y(n1348) );
  MX4X1 U472 ( .A(memory[188]), .B(memory[172]), .C(memory[156]), .D(
        memory[140]), .S0(n1467), .S1(n1448), .Y(n1349) );
  MX4X1 U473 ( .A(n1370), .B(n1368), .C(n1369), .D(n1367), .S0(n1428), .S1(
        n1431), .Y(n1371) );
  MX4X1 U474 ( .A(memory[253]), .B(memory[237]), .C(memory[221]), .D(
        memory[205]), .S0(n1469), .S1(n1449), .Y(n1370) );
  MX4X1 U475 ( .A(memory[125]), .B(memory[109]), .C(memory[93]), .D(memory[77]), .S0(n1469), .S1(n1449), .Y(n1368) );
  MX4X1 U476 ( .A(memory[189]), .B(memory[173]), .C(memory[157]), .D(
        memory[141]), .S0(n1469), .S1(n1449), .Y(n1369) );
  MX4X1 U477 ( .A(n1390), .B(n1388), .C(n1389), .D(n1387), .S0(n1427), .S1(
        n1431), .Y(n1391) );
  MX4X1 U478 ( .A(memory[254]), .B(memory[238]), .C(memory[222]), .D(
        memory[206]), .S0(n1470), .S1(n1450), .Y(n1390) );
  MX4X1 U479 ( .A(memory[126]), .B(memory[110]), .C(memory[94]), .D(memory[78]), .S0(n1470), .S1(n1450), .Y(n1388) );
  MX4X1 U480 ( .A(memory[190]), .B(memory[174]), .C(memory[158]), .D(
        memory[142]), .S0(n1470), .S1(n1450), .Y(n1389) );
  MX4X1 U481 ( .A(n1410), .B(n1408), .C(n1409), .D(n1407), .S0(n1430), .S1(
        addr[2]), .Y(n1411) );
  MX4X1 U482 ( .A(memory[255]), .B(memory[239]), .C(memory[223]), .D(
        memory[207]), .S0(n1471), .S1(n1445), .Y(n1410) );
  MX4X1 U483 ( .A(memory[127]), .B(memory[111]), .C(memory[95]), .D(memory[79]), .S0(n1471), .S1(n1443), .Y(n1408) );
  MX4X1 U484 ( .A(memory[191]), .B(memory[175]), .C(memory[159]), .D(
        memory[143]), .S0(n1471), .S1(n1437), .Y(n1409) );
  MX4X1 U485 ( .A(memory[880]), .B(memory[864]), .C(memory[848]), .D(
        memory[832]), .S0(n1452), .S1(n1444), .Y(n98) );
  MX4X1 U486 ( .A(memory[112]), .B(memory[96]), .C(memory[80]), .D(memory[64]), 
        .S0(n1460), .S1(n1450), .Y(n81) );
  MX4X1 U487 ( .A(memory[369]), .B(memory[353]), .C(memory[337]), .D(
        memory[321]), .S0(n1453), .S1(n1435), .Y(n1133) );
  MX4X1 U488 ( .A(memory[881]), .B(memory[865]), .C(memory[849]), .D(
        memory[833]), .S0(n1454), .S1(n1436), .Y(n1143) );
  MX4X1 U489 ( .A(memory[370]), .B(memory[354]), .C(memory[338]), .D(
        memory[322]), .S0(n1454), .S1(n1436), .Y(n1153) );
  MX4X1 U490 ( .A(memory[882]), .B(memory[866]), .C(memory[850]), .D(
        memory[834]), .S0(n1455), .S1(n1437), .Y(n1163) );
  MX4X1 U491 ( .A(memory[371]), .B(memory[355]), .C(memory[339]), .D(
        memory[323]), .S0(n1456), .S1(n1438), .Y(n1173) );
  MX4X1 U492 ( .A(memory[883]), .B(memory[867]), .C(memory[851]), .D(
        memory[835]), .S0(n1456), .S1(n1438), .Y(n1183) );
  MX4X1 U493 ( .A(memory[372]), .B(memory[356]), .C(memory[340]), .D(
        memory[324]), .S0(n1457), .S1(n1439), .Y(n1193) );
  MX4X1 U494 ( .A(memory[884]), .B(memory[868]), .C(memory[852]), .D(
        memory[836]), .S0(n1458), .S1(n1440), .Y(n1203) );
  MX4X1 U495 ( .A(memory[373]), .B(memory[357]), .C(memory[341]), .D(
        memory[325]), .S0(n1458), .S1(n1440), .Y(n1213) );
  MX4X1 U496 ( .A(memory[885]), .B(memory[869]), .C(memory[853]), .D(
        memory[837]), .S0(n1459), .S1(n1450), .Y(n1223) );
  MX4X1 U497 ( .A(memory[374]), .B(memory[358]), .C(memory[342]), .D(
        memory[326]), .S0(n1460), .S1(n1441), .Y(n1233) );
  MX4X1 U498 ( .A(memory[886]), .B(memory[870]), .C(memory[854]), .D(
        memory[838]), .S0(n1460), .S1(n1441), .Y(n1243) );
  MX4X1 U499 ( .A(memory[375]), .B(memory[359]), .C(memory[343]), .D(
        memory[327]), .S0(n1461), .S1(n1442), .Y(n1253) );
  MX4X1 U500 ( .A(memory[887]), .B(memory[871]), .C(memory[855]), .D(
        memory[839]), .S0(n1462), .S1(n1443), .Y(n1263) );
  MX4X1 U501 ( .A(memory[376]), .B(memory[360]), .C(memory[344]), .D(
        memory[328]), .S0(n1462), .S1(n1443), .Y(n1273) );
  MX4X1 U502 ( .A(memory[888]), .B(memory[872]), .C(memory[856]), .D(
        memory[840]), .S0(n1463), .S1(n1444), .Y(n1283) );
  MX4X1 U503 ( .A(memory[377]), .B(memory[361]), .C(memory[345]), .D(
        memory[329]), .S0(n1464), .S1(n1445), .Y(n1293) );
  MX4X1 U504 ( .A(memory[889]), .B(memory[873]), .C(memory[857]), .D(
        memory[841]), .S0(n1464), .S1(n1445), .Y(n1303) );
  MX4X1 U505 ( .A(memory[378]), .B(memory[362]), .C(memory[346]), .D(
        memory[330]), .S0(n1465), .S1(n1446), .Y(n1313) );
  MX4X1 U506 ( .A(memory[890]), .B(memory[874]), .C(memory[858]), .D(
        memory[842]), .S0(n1466), .S1(n1447), .Y(n1323) );
  MX4X1 U507 ( .A(memory[379]), .B(memory[363]), .C(memory[347]), .D(
        memory[331]), .S0(n1466), .S1(n1447), .Y(n1333) );
  MX4X1 U508 ( .A(memory[891]), .B(memory[875]), .C(memory[859]), .D(
        memory[843]), .S0(n1467), .S1(n1448), .Y(n1343) );
  MX4X1 U509 ( .A(memory[380]), .B(memory[364]), .C(memory[348]), .D(
        memory[332]), .S0(n1468), .S1(n1443), .Y(n1353) );
  MX4X1 U510 ( .A(memory[892]), .B(memory[876]), .C(memory[860]), .D(
        memory[844]), .S0(n1468), .S1(n1445), .Y(n1363) );
  MX4X1 U511 ( .A(memory[381]), .B(memory[365]), .C(memory[349]), .D(
        memory[333]), .S0(n1469), .S1(n1449), .Y(n1373) );
  MX4X1 U512 ( .A(memory[893]), .B(memory[877]), .C(memory[861]), .D(
        memory[845]), .S0(n1470), .S1(n1450), .Y(n1383) );
  MX4X1 U513 ( .A(memory[382]), .B(memory[366]), .C(memory[350]), .D(
        memory[334]), .S0(n1470), .S1(n1450), .Y(n1393) );
  MX4X1 U514 ( .A(memory[894]), .B(memory[878]), .C(memory[862]), .D(
        memory[846]), .S0(n1471), .S1(n1438), .Y(n1403) );
  MX4X1 U515 ( .A(memory[383]), .B(memory[367]), .C(memory[351]), .D(
        memory[335]), .S0(n1467), .S1(n1451), .Y(n1413) );
  MX4X1 U516 ( .A(memory[895]), .B(memory[879]), .C(memory[863]), .D(
        memory[847]), .S0(n1469), .S1(n1451), .Y(n1423) );
  MX4X1 U517 ( .A(n89), .B(n87), .C(n88), .D(n85), .S0(n1429), .S1(addr[2]), 
        .Y(n90) );
  MX4X1 U518 ( .A(memory[496]), .B(memory[480]), .C(memory[464]), .D(
        memory[448]), .S0(n1452), .S1(n1449), .Y(n89) );
  MX4X1 U519 ( .A(memory[368]), .B(memory[352]), .C(memory[336]), .D(
        memory[320]), .S0(n1452), .S1(n1448), .Y(n87) );
  MX4X1 U520 ( .A(memory[432]), .B(memory[416]), .C(memory[400]), .D(
        memory[384]), .S0(n1452), .S1(n1451), .Y(n88) );
  OAI2BB2X1 U521 ( .B0(n1), .B1(n1505), .A0N(memory[0]), .A1N(n1), .Y(n104) );
  OAI2BB2X1 U522 ( .B0(n1), .B1(n1503), .A0N(memory[1]), .A1N(n1), .Y(n105) );
  OAI2BB2X1 U523 ( .B0(n1), .B1(n1501), .A0N(memory[2]), .A1N(n1), .Y(n106) );
  OAI2BB2X1 U524 ( .B0(n1), .B1(n1499), .A0N(memory[3]), .A1N(n1), .Y(n107) );
  OAI2BB2X1 U525 ( .B0(n1), .B1(n1497), .A0N(memory[4]), .A1N(n1), .Y(n108) );
  OAI2BB2X1 U526 ( .B0(n1), .B1(n1495), .A0N(memory[5]), .A1N(n1), .Y(n109) );
  OAI2BB2X1 U527 ( .B0(n1), .B1(n1493), .A0N(memory[6]), .A1N(n1), .Y(n110) );
  OAI2BB2X1 U528 ( .B0(n1), .B1(n1491), .A0N(memory[7]), .A1N(n1), .Y(n111) );
  OAI2BB2X1 U529 ( .B0(n1), .B1(n1489), .A0N(memory[8]), .A1N(n1), .Y(n112) );
  OAI2BB2X1 U530 ( .B0(n1), .B1(n1487), .A0N(memory[9]), .A1N(n1), .Y(n113) );
  OAI2BB2X1 U531 ( .B0(n1), .B1(n1485), .A0N(memory[10]), .A1N(n1), .Y(n114)
         );
  OAI2BB2X1 U532 ( .B0(n1), .B1(n1483), .A0N(memory[11]), .A1N(n1), .Y(n115)
         );
  OAI2BB2X1 U533 ( .B0(n1), .B1(n1481), .A0N(memory[12]), .A1N(n1), .Y(n116)
         );
  OAI2BB2X1 U534 ( .B0(n1), .B1(n1479), .A0N(memory[13]), .A1N(n1), .Y(n117)
         );
  OAI2BB2X1 U535 ( .B0(n1), .B1(n1477), .A0N(memory[14]), .A1N(n1), .Y(n118)
         );
  OAI2BB2X1 U536 ( .B0(n1), .B1(n1475), .A0N(memory[15]), .A1N(n1), .Y(n119)
         );
  OAI2BB2X1 U537 ( .B0(n1505), .B1(n2), .A0N(memory[16]), .A1N(n2), .Y(n120)
         );
  OAI2BB2X1 U538 ( .B0(n1503), .B1(n2), .A0N(memory[17]), .A1N(n2), .Y(n121)
         );
  OAI2BB2X1 U539 ( .B0(n1501), .B1(n2), .A0N(memory[18]), .A1N(n2), .Y(n122)
         );
  OAI2BB2X1 U540 ( .B0(n1499), .B1(n2), .A0N(memory[19]), .A1N(n2), .Y(n123)
         );
  OAI2BB2X1 U541 ( .B0(n1497), .B1(n2), .A0N(memory[20]), .A1N(n2), .Y(n124)
         );
  OAI2BB2X1 U542 ( .B0(n1495), .B1(n2), .A0N(memory[21]), .A1N(n2), .Y(n125)
         );
  OAI2BB2X1 U543 ( .B0(n1493), .B1(n2), .A0N(memory[22]), .A1N(n2), .Y(n126)
         );
  OAI2BB2X1 U544 ( .B0(n1491), .B1(n2), .A0N(memory[23]), .A1N(n2), .Y(n127)
         );
  OAI2BB2X1 U545 ( .B0(n1481), .B1(n2), .A0N(memory[28]), .A1N(n2), .Y(n132)
         );
  OAI2BB2X1 U546 ( .B0(n1479), .B1(n2), .A0N(memory[29]), .A1N(n2), .Y(n133)
         );
  OAI2BB2X1 U547 ( .B0(n1477), .B1(n2), .A0N(memory[30]), .A1N(n2), .Y(n134)
         );
  OAI2BB2X1 U548 ( .B0(n1475), .B1(n2), .A0N(memory[31]), .A1N(n2), .Y(n135)
         );
  OAI2BB2X1 U549 ( .B0(n1504), .B1(n66), .A0N(memory[32]), .A1N(n66), .Y(n136)
         );
  OAI2BB2X1 U550 ( .B0(n1502), .B1(n66), .A0N(memory[33]), .A1N(n66), .Y(n137)
         );
  OAI2BB2X1 U551 ( .B0(n1500), .B1(n66), .A0N(memory[34]), .A1N(n66), .Y(n138)
         );
  OAI2BB2X1 U552 ( .B0(n1498), .B1(n66), .A0N(memory[35]), .A1N(n66), .Y(n139)
         );
  OAI2BB2X1 U553 ( .B0(n1496), .B1(n66), .A0N(memory[36]), .A1N(n66), .Y(n140)
         );
  OAI2BB2X1 U554 ( .B0(n1494), .B1(n66), .A0N(memory[37]), .A1N(n66), .Y(n141)
         );
  OAI2BB2X1 U555 ( .B0(n1492), .B1(n66), .A0N(memory[38]), .A1N(n66), .Y(n142)
         );
  OAI2BB2X1 U556 ( .B0(n1490), .B1(n66), .A0N(memory[39]), .A1N(n66), .Y(n143)
         );
  OAI2BB2X1 U557 ( .B0(n1480), .B1(n66), .A0N(memory[44]), .A1N(n66), .Y(n148)
         );
  OAI2BB2X1 U558 ( .B0(n1478), .B1(n66), .A0N(memory[45]), .A1N(n66), .Y(n149)
         );
  OAI2BB2X1 U559 ( .B0(n1476), .B1(n66), .A0N(memory[46]), .A1N(n66), .Y(n150)
         );
  OAI2BB2X1 U560 ( .B0(n1474), .B1(n66), .A0N(memory[47]), .A1N(n66), .Y(n151)
         );
  OAI2BB2X1 U561 ( .B0(n1505), .B1(n3), .A0N(memory[48]), .A1N(n3), .Y(n152)
         );
  OAI2BB2X1 U562 ( .B0(n1503), .B1(n3), .A0N(memory[49]), .A1N(n3), .Y(n153)
         );
  OAI2BB2X1 U563 ( .B0(n1501), .B1(n3), .A0N(memory[50]), .A1N(n3), .Y(n154)
         );
  OAI2BB2X1 U564 ( .B0(n1499), .B1(n3), .A0N(memory[51]), .A1N(n3), .Y(n155)
         );
  OAI2BB2X1 U565 ( .B0(n1497), .B1(n3), .A0N(memory[52]), .A1N(n3), .Y(n156)
         );
  OAI2BB2X1 U566 ( .B0(n1495), .B1(n3), .A0N(memory[53]), .A1N(n3), .Y(n157)
         );
  OAI2BB2X1 U567 ( .B0(n1493), .B1(n3), .A0N(memory[54]), .A1N(n3), .Y(n158)
         );
  OAI2BB2X1 U568 ( .B0(n1491), .B1(n3), .A0N(memory[55]), .A1N(n3), .Y(n159)
         );
  OAI2BB2X1 U569 ( .B0(n1481), .B1(n3), .A0N(memory[60]), .A1N(n3), .Y(n164)
         );
  OAI2BB2X1 U570 ( .B0(n1479), .B1(n3), .A0N(memory[61]), .A1N(n3), .Y(n165)
         );
  OAI2BB2X1 U571 ( .B0(n1477), .B1(n3), .A0N(memory[62]), .A1N(n3), .Y(n166)
         );
  OAI2BB2X1 U572 ( .B0(n1475), .B1(n3), .A0N(memory[63]), .A1N(n3), .Y(n167)
         );
  OAI2BB2X1 U573 ( .B0(n1505), .B1(n67), .A0N(memory[64]), .A1N(n67), .Y(n168)
         );
  OAI2BB2X1 U574 ( .B0(n1503), .B1(n67), .A0N(memory[65]), .A1N(n67), .Y(n169)
         );
  OAI2BB2X1 U575 ( .B0(n1501), .B1(n67), .A0N(memory[66]), .A1N(n67), .Y(n170)
         );
  OAI2BB2X1 U576 ( .B0(n1499), .B1(n67), .A0N(memory[67]), .A1N(n67), .Y(n171)
         );
  OAI2BB2X1 U577 ( .B0(n1497), .B1(n67), .A0N(memory[68]), .A1N(n67), .Y(n172)
         );
  OAI2BB2X1 U578 ( .B0(n1495), .B1(n67), .A0N(memory[69]), .A1N(n67), .Y(n173)
         );
  OAI2BB2X1 U579 ( .B0(n1493), .B1(n67), .A0N(memory[70]), .A1N(n67), .Y(n174)
         );
  OAI2BB2X1 U580 ( .B0(n1491), .B1(n67), .A0N(memory[71]), .A1N(n67), .Y(n175)
         );
  OAI2BB2X1 U581 ( .B0(n1481), .B1(n67), .A0N(memory[76]), .A1N(n67), .Y(n180)
         );
  OAI2BB2X1 U582 ( .B0(n1479), .B1(n67), .A0N(memory[77]), .A1N(n67), .Y(n181)
         );
  OAI2BB2X1 U583 ( .B0(n1477), .B1(n67), .A0N(memory[78]), .A1N(n67), .Y(n182)
         );
  OAI2BB2X1 U584 ( .B0(n1475), .B1(n67), .A0N(memory[79]), .A1N(n67), .Y(n183)
         );
  OAI2BB2X1 U585 ( .B0(n1504), .B1(n4), .A0N(memory[80]), .A1N(n4), .Y(n184)
         );
  OAI2BB2X1 U586 ( .B0(n1502), .B1(n4), .A0N(memory[81]), .A1N(n4), .Y(n185)
         );
  OAI2BB2X1 U587 ( .B0(n1500), .B1(n4), .A0N(memory[82]), .A1N(n4), .Y(n186)
         );
  OAI2BB2X1 U588 ( .B0(n1498), .B1(n4), .A0N(memory[83]), .A1N(n4), .Y(n187)
         );
  OAI2BB2X1 U589 ( .B0(n1496), .B1(n4), .A0N(memory[84]), .A1N(n4), .Y(n188)
         );
  OAI2BB2X1 U590 ( .B0(n1494), .B1(n4), .A0N(memory[85]), .A1N(n4), .Y(n189)
         );
  OAI2BB2X1 U591 ( .B0(n1492), .B1(n4), .A0N(memory[86]), .A1N(n4), .Y(n190)
         );
  OAI2BB2X1 U592 ( .B0(n1490), .B1(n4), .A0N(memory[87]), .A1N(n4), .Y(n191)
         );
  OAI2BB2X1 U593 ( .B0(n1480), .B1(n4), .A0N(memory[92]), .A1N(n4), .Y(n196)
         );
  OAI2BB2X1 U594 ( .B0(n1478), .B1(n4), .A0N(memory[93]), .A1N(n4), .Y(n197)
         );
  OAI2BB2X1 U595 ( .B0(n1476), .B1(n4), .A0N(memory[94]), .A1N(n4), .Y(n198)
         );
  OAI2BB2X1 U596 ( .B0(n1474), .B1(n4), .A0N(memory[95]), .A1N(n4), .Y(n199)
         );
  OAI2BB2X1 U597 ( .B0(n1504), .B1(n69), .A0N(memory[96]), .A1N(n69), .Y(n200)
         );
  OAI2BB2X1 U598 ( .B0(n1502), .B1(n69), .A0N(memory[97]), .A1N(n69), .Y(n201)
         );
  OAI2BB2X1 U599 ( .B0(n1500), .B1(n69), .A0N(memory[98]), .A1N(n69), .Y(n202)
         );
  OAI2BB2X1 U600 ( .B0(n1498), .B1(n69), .A0N(memory[99]), .A1N(n69), .Y(n203)
         );
  OAI2BB2X1 U601 ( .B0(n1496), .B1(n69), .A0N(memory[100]), .A1N(n69), .Y(n204) );
  OAI2BB2X1 U602 ( .B0(n1494), .B1(n69), .A0N(memory[101]), .A1N(n69), .Y(n205) );
  OAI2BB2X1 U603 ( .B0(n1492), .B1(n69), .A0N(memory[102]), .A1N(n69), .Y(n206) );
  OAI2BB2X1 U604 ( .B0(n1490), .B1(n69), .A0N(memory[103]), .A1N(n69), .Y(n207) );
  OAI2BB2X1 U605 ( .B0(n1480), .B1(n69), .A0N(memory[108]), .A1N(n69), .Y(n212) );
  OAI2BB2X1 U606 ( .B0(n1478), .B1(n69), .A0N(memory[109]), .A1N(n69), .Y(n213) );
  OAI2BB2X1 U607 ( .B0(n1476), .B1(n69), .A0N(memory[110]), .A1N(n69), .Y(n214) );
  OAI2BB2X1 U608 ( .B0(n1474), .B1(n69), .A0N(memory[111]), .A1N(n69), .Y(n215) );
  OAI2BB2X1 U609 ( .B0(n1505), .B1(n5), .A0N(memory[112]), .A1N(n5), .Y(n216)
         );
  OAI2BB2X1 U610 ( .B0(n1503), .B1(n5), .A0N(memory[113]), .A1N(n5), .Y(n217)
         );
  OAI2BB2X1 U611 ( .B0(n1501), .B1(n5), .A0N(memory[114]), .A1N(n5), .Y(n218)
         );
  OAI2BB2X1 U612 ( .B0(n1499), .B1(n5), .A0N(memory[115]), .A1N(n5), .Y(n219)
         );
  OAI2BB2X1 U613 ( .B0(n1497), .B1(n5), .A0N(memory[116]), .A1N(n5), .Y(n220)
         );
  OAI2BB2X1 U614 ( .B0(n1495), .B1(n5), .A0N(memory[117]), .A1N(n5), .Y(n221)
         );
  OAI2BB2X1 U615 ( .B0(n1493), .B1(n5), .A0N(memory[118]), .A1N(n5), .Y(n222)
         );
  OAI2BB2X1 U616 ( .B0(n1491), .B1(n5), .A0N(memory[119]), .A1N(n5), .Y(n223)
         );
  OAI2BB2X1 U617 ( .B0(n1481), .B1(n5), .A0N(memory[124]), .A1N(n5), .Y(n228)
         );
  OAI2BB2X1 U618 ( .B0(n1479), .B1(n5), .A0N(memory[125]), .A1N(n5), .Y(n229)
         );
  OAI2BB2X1 U619 ( .B0(n1477), .B1(n5), .A0N(memory[126]), .A1N(n5), .Y(n230)
         );
  OAI2BB2X1 U620 ( .B0(n1475), .B1(n5), .A0N(memory[127]), .A1N(n5), .Y(n231)
         );
  OAI2BB2X1 U621 ( .B0(n1504), .B1(n6), .A0N(memory[128]), .A1N(n6), .Y(n232)
         );
  OAI2BB2X1 U622 ( .B0(n1502), .B1(n6), .A0N(memory[129]), .A1N(n6), .Y(n233)
         );
  OAI2BB2X1 U623 ( .B0(n1500), .B1(n6), .A0N(memory[130]), .A1N(n6), .Y(n234)
         );
  OAI2BB2X1 U624 ( .B0(n1498), .B1(n6), .A0N(memory[131]), .A1N(n6), .Y(n235)
         );
  OAI2BB2X1 U625 ( .B0(n1496), .B1(n6), .A0N(memory[132]), .A1N(n6), .Y(n236)
         );
  OAI2BB2X1 U626 ( .B0(n1494), .B1(n6), .A0N(memory[133]), .A1N(n6), .Y(n237)
         );
  OAI2BB2X1 U627 ( .B0(n1492), .B1(n6), .A0N(memory[134]), .A1N(n6), .Y(n238)
         );
  OAI2BB2X1 U628 ( .B0(n1490), .B1(n6), .A0N(memory[135]), .A1N(n6), .Y(n239)
         );
  OAI2BB2X1 U629 ( .B0(n1480), .B1(n6), .A0N(memory[140]), .A1N(n6), .Y(n244)
         );
  OAI2BB2X1 U630 ( .B0(n1478), .B1(n6), .A0N(memory[141]), .A1N(n6), .Y(n245)
         );
  OAI2BB2X1 U631 ( .B0(n1476), .B1(n6), .A0N(memory[142]), .A1N(n6), .Y(n246)
         );
  OAI2BB2X1 U632 ( .B0(n1474), .B1(n6), .A0N(memory[143]), .A1N(n6), .Y(n247)
         );
  OAI2BB2X1 U633 ( .B0(n1505), .B1(n7), .A0N(memory[144]), .A1N(n7), .Y(n248)
         );
  OAI2BB2X1 U634 ( .B0(n1503), .B1(n7), .A0N(memory[145]), .A1N(n7), .Y(n249)
         );
  OAI2BB2X1 U635 ( .B0(n1501), .B1(n7), .A0N(memory[146]), .A1N(n7), .Y(n250)
         );
  OAI2BB2X1 U636 ( .B0(n1499), .B1(n7), .A0N(memory[147]), .A1N(n7), .Y(n251)
         );
  OAI2BB2X1 U637 ( .B0(n1497), .B1(n7), .A0N(memory[148]), .A1N(n7), .Y(n252)
         );
  OAI2BB2X1 U638 ( .B0(n1495), .B1(n7), .A0N(memory[149]), .A1N(n7), .Y(n253)
         );
  OAI2BB2X1 U639 ( .B0(n1493), .B1(n7), .A0N(memory[150]), .A1N(n7), .Y(n254)
         );
  OAI2BB2X1 U640 ( .B0(n1491), .B1(n7), .A0N(memory[151]), .A1N(n7), .Y(n255)
         );
  OAI2BB2X1 U641 ( .B0(n1481), .B1(n7), .A0N(memory[156]), .A1N(n7), .Y(n260)
         );
  OAI2BB2X1 U642 ( .B0(n1479), .B1(n7), .A0N(memory[157]), .A1N(n7), .Y(n261)
         );
  OAI2BB2X1 U643 ( .B0(n1477), .B1(n7), .A0N(memory[158]), .A1N(n7), .Y(n262)
         );
  OAI2BB2X1 U644 ( .B0(n1475), .B1(n7), .A0N(memory[159]), .A1N(n7), .Y(n263)
         );
  OAI2BB2X1 U645 ( .B0(n1504), .B1(n70), .A0N(memory[160]), .A1N(n70), .Y(n264) );
  OAI2BB2X1 U646 ( .B0(n1502), .B1(n70), .A0N(memory[161]), .A1N(n70), .Y(n265) );
  OAI2BB2X1 U647 ( .B0(n1500), .B1(n70), .A0N(memory[162]), .A1N(n70), .Y(n266) );
  OAI2BB2X1 U648 ( .B0(n1498), .B1(n70), .A0N(memory[163]), .A1N(n70), .Y(n267) );
  OAI2BB2X1 U649 ( .B0(n1496), .B1(n70), .A0N(memory[164]), .A1N(n70), .Y(n268) );
  OAI2BB2X1 U650 ( .B0(n1494), .B1(n70), .A0N(memory[165]), .A1N(n70), .Y(n269) );
  OAI2BB2X1 U651 ( .B0(n1492), .B1(n70), .A0N(memory[166]), .A1N(n70), .Y(n270) );
  OAI2BB2X1 U652 ( .B0(n1490), .B1(n70), .A0N(memory[167]), .A1N(n70), .Y(n271) );
  OAI2BB2X1 U653 ( .B0(n1480), .B1(n70), .A0N(memory[172]), .A1N(n70), .Y(n276) );
  OAI2BB2X1 U654 ( .B0(n1478), .B1(n70), .A0N(memory[173]), .A1N(n70), .Y(n277) );
  OAI2BB2X1 U655 ( .B0(n1476), .B1(n70), .A0N(memory[174]), .A1N(n70), .Y(n278) );
  OAI2BB2X1 U656 ( .B0(n1474), .B1(n70), .A0N(memory[175]), .A1N(n70), .Y(n279) );
  OAI2BB2X1 U657 ( .B0(n1505), .B1(n8), .A0N(memory[176]), .A1N(n8), .Y(n280)
         );
  OAI2BB2X1 U658 ( .B0(n1503), .B1(n8), .A0N(memory[177]), .A1N(n8), .Y(n281)
         );
  OAI2BB2X1 U659 ( .B0(n1501), .B1(n8), .A0N(memory[178]), .A1N(n8), .Y(n282)
         );
  OAI2BB2X1 U660 ( .B0(n1499), .B1(n8), .A0N(memory[179]), .A1N(n8), .Y(n283)
         );
  OAI2BB2X1 U661 ( .B0(n1497), .B1(n8), .A0N(memory[180]), .A1N(n8), .Y(n284)
         );
  OAI2BB2X1 U662 ( .B0(n1495), .B1(n8), .A0N(memory[181]), .A1N(n8), .Y(n285)
         );
  OAI2BB2X1 U663 ( .B0(n1493), .B1(n8), .A0N(memory[182]), .A1N(n8), .Y(n286)
         );
  OAI2BB2X1 U664 ( .B0(n1491), .B1(n8), .A0N(memory[183]), .A1N(n8), .Y(n287)
         );
  OAI2BB2X1 U665 ( .B0(n1481), .B1(n8), .A0N(memory[188]), .A1N(n8), .Y(n292)
         );
  OAI2BB2X1 U666 ( .B0(n1479), .B1(n8), .A0N(memory[189]), .A1N(n8), .Y(n293)
         );
  OAI2BB2X1 U667 ( .B0(n1477), .B1(n8), .A0N(memory[190]), .A1N(n8), .Y(n294)
         );
  OAI2BB2X1 U668 ( .B0(n1475), .B1(n8), .A0N(memory[191]), .A1N(n8), .Y(n295)
         );
  OAI2BB2X1 U669 ( .B0(n1505), .B1(n71), .A0N(memory[192]), .A1N(n71), .Y(n296) );
  OAI2BB2X1 U670 ( .B0(n1503), .B1(n71), .A0N(memory[193]), .A1N(n71), .Y(n297) );
  OAI2BB2X1 U671 ( .B0(n1501), .B1(n71), .A0N(memory[194]), .A1N(n71), .Y(n298) );
  OAI2BB2X1 U672 ( .B0(n1499), .B1(n71), .A0N(memory[195]), .A1N(n71), .Y(n299) );
  OAI2BB2X1 U673 ( .B0(n1497), .B1(n71), .A0N(memory[196]), .A1N(n71), .Y(n300) );
  OAI2BB2X1 U674 ( .B0(n1495), .B1(n71), .A0N(memory[197]), .A1N(n71), .Y(n301) );
  OAI2BB2X1 U675 ( .B0(n1493), .B1(n71), .A0N(memory[198]), .A1N(n71), .Y(n302) );
  OAI2BB2X1 U676 ( .B0(n1491), .B1(n71), .A0N(memory[199]), .A1N(n71), .Y(n303) );
  OAI2BB2X1 U677 ( .B0(n1481), .B1(n71), .A0N(memory[204]), .A1N(n71), .Y(n308) );
  OAI2BB2X1 U678 ( .B0(n1479), .B1(n71), .A0N(memory[205]), .A1N(n71), .Y(n309) );
  OAI2BB2X1 U679 ( .B0(n1477), .B1(n71), .A0N(memory[206]), .A1N(n71), .Y(n310) );
  OAI2BB2X1 U680 ( .B0(n1475), .B1(n71), .A0N(memory[207]), .A1N(n71), .Y(n311) );
  OAI2BB2X1 U681 ( .B0(n1505), .B1(n9), .A0N(memory[208]), .A1N(n9), .Y(n312)
         );
  OAI2BB2X1 U682 ( .B0(n1503), .B1(n9), .A0N(memory[209]), .A1N(n9), .Y(n313)
         );
  OAI2BB2X1 U683 ( .B0(n1501), .B1(n9), .A0N(memory[210]), .A1N(n9), .Y(n314)
         );
  OAI2BB2X1 U684 ( .B0(n1499), .B1(n9), .A0N(memory[211]), .A1N(n9), .Y(n315)
         );
  OAI2BB2X1 U685 ( .B0(n1497), .B1(n9), .A0N(memory[212]), .A1N(n9), .Y(n316)
         );
  OAI2BB2X1 U686 ( .B0(n1495), .B1(n9), .A0N(memory[213]), .A1N(n9), .Y(n317)
         );
  OAI2BB2X1 U687 ( .B0(n1493), .B1(n9), .A0N(memory[214]), .A1N(n9), .Y(n318)
         );
  OAI2BB2X1 U688 ( .B0(n1491), .B1(n9), .A0N(memory[215]), .A1N(n9), .Y(n319)
         );
  OAI2BB2X1 U689 ( .B0(n1481), .B1(n9), .A0N(memory[220]), .A1N(n9), .Y(n324)
         );
  OAI2BB2X1 U690 ( .B0(n1479), .B1(n9), .A0N(memory[221]), .A1N(n9), .Y(n325)
         );
  OAI2BB2X1 U691 ( .B0(n1477), .B1(n9), .A0N(memory[222]), .A1N(n9), .Y(n326)
         );
  OAI2BB2X1 U692 ( .B0(n1475), .B1(n9), .A0N(memory[223]), .A1N(n9), .Y(n327)
         );
  OAI2BB2X1 U693 ( .B0(n1505), .B1(n72), .A0N(memory[224]), .A1N(n72), .Y(n328) );
  OAI2BB2X1 U694 ( .B0(n1503), .B1(n72), .A0N(memory[225]), .A1N(n72), .Y(n329) );
  OAI2BB2X1 U695 ( .B0(n1501), .B1(n72), .A0N(memory[226]), .A1N(n72), .Y(n330) );
  OAI2BB2X1 U696 ( .B0(n1499), .B1(n72), .A0N(memory[227]), .A1N(n72), .Y(n331) );
  OAI2BB2X1 U697 ( .B0(n1497), .B1(n72), .A0N(memory[228]), .A1N(n72), .Y(n332) );
  OAI2BB2X1 U698 ( .B0(n1495), .B1(n72), .A0N(memory[229]), .A1N(n72), .Y(n333) );
  OAI2BB2X1 U699 ( .B0(n1493), .B1(n72), .A0N(memory[230]), .A1N(n72), .Y(n334) );
  OAI2BB2X1 U700 ( .B0(n1491), .B1(n72), .A0N(memory[231]), .A1N(n72), .Y(n335) );
  OAI2BB2X1 U701 ( .B0(n1481), .B1(n72), .A0N(memory[236]), .A1N(n72), .Y(n340) );
  OAI2BB2X1 U702 ( .B0(n1479), .B1(n72), .A0N(memory[237]), .A1N(n72), .Y(n341) );
  OAI2BB2X1 U703 ( .B0(n1477), .B1(n72), .A0N(memory[238]), .A1N(n72), .Y(n342) );
  OAI2BB2X1 U704 ( .B0(n1475), .B1(n72), .A0N(memory[239]), .A1N(n72), .Y(n343) );
  OAI2BB2X1 U705 ( .B0(n1505), .B1(n10), .A0N(memory[240]), .A1N(n10), .Y(n344) );
  OAI2BB2X1 U706 ( .B0(n1503), .B1(n10), .A0N(memory[241]), .A1N(n10), .Y(n345) );
  OAI2BB2X1 U707 ( .B0(n1501), .B1(n10), .A0N(memory[242]), .A1N(n10), .Y(n346) );
  OAI2BB2X1 U708 ( .B0(n1499), .B1(n10), .A0N(memory[243]), .A1N(n10), .Y(n347) );
  OAI2BB2X1 U709 ( .B0(n1497), .B1(n10), .A0N(memory[244]), .A1N(n10), .Y(n348) );
  OAI2BB2X1 U710 ( .B0(n1495), .B1(n10), .A0N(memory[245]), .A1N(n10), .Y(n349) );
  OAI2BB2X1 U711 ( .B0(n1493), .B1(n10), .A0N(memory[246]), .A1N(n10), .Y(n350) );
  OAI2BB2X1 U712 ( .B0(n1491), .B1(n10), .A0N(memory[247]), .A1N(n10), .Y(n351) );
  OAI2BB2X1 U713 ( .B0(n1481), .B1(n10), .A0N(memory[252]), .A1N(n10), .Y(n356) );
  OAI2BB2X1 U714 ( .B0(n1479), .B1(n10), .A0N(memory[253]), .A1N(n10), .Y(n357) );
  OAI2BB2X1 U715 ( .B0(n1477), .B1(n10), .A0N(memory[254]), .A1N(n10), .Y(n358) );
  OAI2BB2X1 U716 ( .B0(n1475), .B1(n10), .A0N(memory[255]), .A1N(n10), .Y(n359) );
  OAI2BB2X1 U717 ( .B0(n1505), .B1(n11), .A0N(memory[256]), .A1N(n11), .Y(n360) );
  OAI2BB2X1 U718 ( .B0(n1503), .B1(n11), .A0N(memory[257]), .A1N(n11), .Y(n361) );
  OAI2BB2X1 U719 ( .B0(n1501), .B1(n11), .A0N(memory[258]), .A1N(n11), .Y(n362) );
  OAI2BB2X1 U720 ( .B0(n1499), .B1(n11), .A0N(memory[259]), .A1N(n11), .Y(n363) );
  OAI2BB2X1 U721 ( .B0(n1497), .B1(n11), .A0N(memory[260]), .A1N(n11), .Y(n364) );
  OAI2BB2X1 U722 ( .B0(n1495), .B1(n11), .A0N(memory[261]), .A1N(n11), .Y(n365) );
  OAI2BB2X1 U723 ( .B0(n1493), .B1(n11), .A0N(memory[262]), .A1N(n11), .Y(n366) );
  OAI2BB2X1 U724 ( .B0(n1491), .B1(n11), .A0N(memory[263]), .A1N(n11), .Y(n367) );
  OAI2BB2X1 U725 ( .B0(n1481), .B1(n11), .A0N(memory[268]), .A1N(n11), .Y(n372) );
  OAI2BB2X1 U726 ( .B0(n1479), .B1(n11), .A0N(memory[269]), .A1N(n11), .Y(n373) );
  OAI2BB2X1 U727 ( .B0(n1477), .B1(n11), .A0N(memory[270]), .A1N(n11), .Y(n374) );
  OAI2BB2X1 U728 ( .B0(n1475), .B1(n11), .A0N(memory[271]), .A1N(n11), .Y(n375) );
  OAI2BB2X1 U729 ( .B0(n1505), .B1(n12), .A0N(memory[272]), .A1N(n12), .Y(n376) );
  OAI2BB2X1 U730 ( .B0(n1503), .B1(n12), .A0N(memory[273]), .A1N(n12), .Y(n377) );
  OAI2BB2X1 U731 ( .B0(n1501), .B1(n12), .A0N(memory[274]), .A1N(n12), .Y(n378) );
  OAI2BB2X1 U732 ( .B0(n1499), .B1(n12), .A0N(memory[275]), .A1N(n12), .Y(n379) );
  OAI2BB2X1 U733 ( .B0(n1497), .B1(n12), .A0N(memory[276]), .A1N(n12), .Y(n380) );
  OAI2BB2X1 U734 ( .B0(n1495), .B1(n12), .A0N(memory[277]), .A1N(n12), .Y(n381) );
  OAI2BB2X1 U735 ( .B0(n1493), .B1(n12), .A0N(memory[278]), .A1N(n12), .Y(n382) );
  OAI2BB2X1 U736 ( .B0(n1491), .B1(n12), .A0N(memory[279]), .A1N(n12), .Y(n383) );
  OAI2BB2X1 U737 ( .B0(n1481), .B1(n12), .A0N(memory[284]), .A1N(n12), .Y(n388) );
  OAI2BB2X1 U738 ( .B0(n1479), .B1(n12), .A0N(memory[285]), .A1N(n12), .Y(n389) );
  OAI2BB2X1 U739 ( .B0(n1477), .B1(n12), .A0N(memory[286]), .A1N(n12), .Y(n390) );
  OAI2BB2X1 U740 ( .B0(n1475), .B1(n12), .A0N(memory[287]), .A1N(n12), .Y(n391) );
  OAI2BB2X1 U741 ( .B0(n1505), .B1(n73), .A0N(memory[288]), .A1N(n73), .Y(n392) );
  OAI2BB2X1 U742 ( .B0(n1503), .B1(n73), .A0N(memory[289]), .A1N(n73), .Y(n393) );
  OAI2BB2X1 U743 ( .B0(n1501), .B1(n73), .A0N(memory[290]), .A1N(n73), .Y(n394) );
  OAI2BB2X1 U744 ( .B0(n1499), .B1(n73), .A0N(memory[291]), .A1N(n73), .Y(n395) );
  OAI2BB2X1 U745 ( .B0(n1497), .B1(n73), .A0N(memory[292]), .A1N(n73), .Y(n396) );
  OAI2BB2X1 U746 ( .B0(n1495), .B1(n73), .A0N(memory[293]), .A1N(n73), .Y(n397) );
  OAI2BB2X1 U747 ( .B0(n1493), .B1(n73), .A0N(memory[294]), .A1N(n73), .Y(n398) );
  OAI2BB2X1 U748 ( .B0(n1491), .B1(n73), .A0N(memory[295]), .A1N(n73), .Y(n399) );
  OAI2BB2X1 U749 ( .B0(n1481), .B1(n73), .A0N(memory[300]), .A1N(n73), .Y(n404) );
  OAI2BB2X1 U750 ( .B0(n1479), .B1(n73), .A0N(memory[301]), .A1N(n73), .Y(n405) );
  OAI2BB2X1 U751 ( .B0(n1477), .B1(n73), .A0N(memory[302]), .A1N(n73), .Y(n406) );
  OAI2BB2X1 U752 ( .B0(n1475), .B1(n73), .A0N(memory[303]), .A1N(n73), .Y(n407) );
  OAI2BB2X1 U753 ( .B0(n1505), .B1(n13), .A0N(memory[304]), .A1N(n13), .Y(n408) );
  OAI2BB2X1 U754 ( .B0(n1503), .B1(n13), .A0N(memory[305]), .A1N(n13), .Y(n409) );
  OAI2BB2X1 U755 ( .B0(n1501), .B1(n13), .A0N(memory[306]), .A1N(n13), .Y(n410) );
  OAI2BB2X1 U756 ( .B0(n1499), .B1(n13), .A0N(memory[307]), .A1N(n13), .Y(n411) );
  OAI2BB2X1 U757 ( .B0(n1497), .B1(n13), .A0N(memory[308]), .A1N(n13), .Y(n412) );
  OAI2BB2X1 U758 ( .B0(n1495), .B1(n13), .A0N(memory[309]), .A1N(n13), .Y(n413) );
  OAI2BB2X1 U759 ( .B0(n1493), .B1(n13), .A0N(memory[310]), .A1N(n13), .Y(n414) );
  OAI2BB2X1 U760 ( .B0(n1491), .B1(n13), .A0N(memory[311]), .A1N(n13), .Y(n415) );
  OAI2BB2X1 U761 ( .B0(n1481), .B1(n13), .A0N(memory[316]), .A1N(n13), .Y(n420) );
  OAI2BB2X1 U762 ( .B0(n1479), .B1(n13), .A0N(memory[317]), .A1N(n13), .Y(n421) );
  OAI2BB2X1 U763 ( .B0(n1477), .B1(n13), .A0N(memory[318]), .A1N(n13), .Y(n422) );
  OAI2BB2X1 U764 ( .B0(n1475), .B1(n13), .A0N(memory[319]), .A1N(n13), .Y(n423) );
  OAI2BB2X1 U765 ( .B0(n1505), .B1(n74), .A0N(memory[320]), .A1N(n74), .Y(n424) );
  OAI2BB2X1 U766 ( .B0(n1503), .B1(n74), .A0N(memory[321]), .A1N(n74), .Y(n425) );
  OAI2BB2X1 U767 ( .B0(n1501), .B1(n74), .A0N(memory[322]), .A1N(n74), .Y(n426) );
  OAI2BB2X1 U768 ( .B0(n1499), .B1(n74), .A0N(memory[323]), .A1N(n74), .Y(n427) );
  OAI2BB2X1 U769 ( .B0(n1497), .B1(n74), .A0N(memory[324]), .A1N(n74), .Y(n428) );
  OAI2BB2X1 U770 ( .B0(n1495), .B1(n74), .A0N(memory[325]), .A1N(n74), .Y(n429) );
  OAI2BB2X1 U771 ( .B0(n1493), .B1(n74), .A0N(memory[326]), .A1N(n74), .Y(n430) );
  OAI2BB2X1 U772 ( .B0(n1491), .B1(n74), .A0N(memory[327]), .A1N(n74), .Y(n431) );
  OAI2BB2X1 U773 ( .B0(n1481), .B1(n74), .A0N(memory[332]), .A1N(n74), .Y(n436) );
  OAI2BB2X1 U774 ( .B0(n1479), .B1(n74), .A0N(memory[333]), .A1N(n74), .Y(n437) );
  OAI2BB2X1 U775 ( .B0(n1477), .B1(n74), .A0N(memory[334]), .A1N(n74), .Y(n438) );
  OAI2BB2X1 U776 ( .B0(n1475), .B1(n74), .A0N(memory[335]), .A1N(n74), .Y(n439) );
  OAI2BB2X1 U777 ( .B0(n1505), .B1(n14), .A0N(memory[336]), .A1N(n14), .Y(n440) );
  OAI2BB2X1 U778 ( .B0(n1503), .B1(n14), .A0N(memory[337]), .A1N(n14), .Y(n441) );
  OAI2BB2X1 U779 ( .B0(n1501), .B1(n14), .A0N(memory[338]), .A1N(n14), .Y(n442) );
  OAI2BB2X1 U780 ( .B0(n1499), .B1(n14), .A0N(memory[339]), .A1N(n14), .Y(n443) );
  OAI2BB2X1 U781 ( .B0(n1497), .B1(n14), .A0N(memory[340]), .A1N(n14), .Y(n444) );
  OAI2BB2X1 U782 ( .B0(n1495), .B1(n14), .A0N(memory[341]), .A1N(n14), .Y(n445) );
  OAI2BB2X1 U783 ( .B0(n1493), .B1(n14), .A0N(memory[342]), .A1N(n14), .Y(n446) );
  OAI2BB2X1 U784 ( .B0(n1491), .B1(n14), .A0N(memory[343]), .A1N(n14), .Y(n447) );
  OAI2BB2X1 U785 ( .B0(n1481), .B1(n14), .A0N(memory[348]), .A1N(n14), .Y(n452) );
  OAI2BB2X1 U786 ( .B0(n1479), .B1(n14), .A0N(memory[349]), .A1N(n14), .Y(n453) );
  OAI2BB2X1 U787 ( .B0(n1477), .B1(n14), .A0N(memory[350]), .A1N(n14), .Y(n454) );
  OAI2BB2X1 U788 ( .B0(n1475), .B1(n14), .A0N(memory[351]), .A1N(n14), .Y(n455) );
  OAI2BB2X1 U789 ( .B0(n1505), .B1(n75), .A0N(memory[352]), .A1N(n75), .Y(n456) );
  OAI2BB2X1 U790 ( .B0(n1503), .B1(n75), .A0N(memory[353]), .A1N(n75), .Y(n457) );
  OAI2BB2X1 U791 ( .B0(n1501), .B1(n75), .A0N(memory[354]), .A1N(n75), .Y(n458) );
  OAI2BB2X1 U792 ( .B0(n1499), .B1(n75), .A0N(memory[355]), .A1N(n75), .Y(n459) );
  OAI2BB2X1 U793 ( .B0(n1497), .B1(n75), .A0N(memory[356]), .A1N(n75), .Y(n460) );
  OAI2BB2X1 U794 ( .B0(n1495), .B1(n75), .A0N(memory[357]), .A1N(n75), .Y(n461) );
  OAI2BB2X1 U795 ( .B0(n1493), .B1(n75), .A0N(memory[358]), .A1N(n75), .Y(n462) );
  OAI2BB2X1 U796 ( .B0(n1491), .B1(n75), .A0N(memory[359]), .A1N(n75), .Y(n463) );
  OAI2BB2X1 U797 ( .B0(n1481), .B1(n75), .A0N(memory[364]), .A1N(n75), .Y(n468) );
  OAI2BB2X1 U798 ( .B0(n1479), .B1(n75), .A0N(memory[365]), .A1N(n75), .Y(n469) );
  OAI2BB2X1 U799 ( .B0(n1477), .B1(n75), .A0N(memory[366]), .A1N(n75), .Y(n470) );
  OAI2BB2X1 U800 ( .B0(n1475), .B1(n75), .A0N(memory[367]), .A1N(n75), .Y(n471) );
  OAI2BB2X1 U801 ( .B0(n1505), .B1(n15), .A0N(memory[368]), .A1N(n15), .Y(n472) );
  OAI2BB2X1 U802 ( .B0(n1503), .B1(n15), .A0N(memory[369]), .A1N(n15), .Y(n473) );
  OAI2BB2X1 U803 ( .B0(n1501), .B1(n15), .A0N(memory[370]), .A1N(n15), .Y(n474) );
  OAI2BB2X1 U804 ( .B0(n1499), .B1(n15), .A0N(memory[371]), .A1N(n15), .Y(n475) );
  OAI2BB2X1 U805 ( .B0(n1497), .B1(n15), .A0N(memory[372]), .A1N(n15), .Y(n476) );
  OAI2BB2X1 U806 ( .B0(n1495), .B1(n15), .A0N(memory[373]), .A1N(n15), .Y(n477) );
  OAI2BB2X1 U807 ( .B0(n1493), .B1(n15), .A0N(memory[374]), .A1N(n15), .Y(n478) );
  OAI2BB2X1 U808 ( .B0(n1491), .B1(n15), .A0N(memory[375]), .A1N(n15), .Y(n479) );
  OAI2BB2X1 U809 ( .B0(n1481), .B1(n15), .A0N(memory[380]), .A1N(n15), .Y(n484) );
  OAI2BB2X1 U810 ( .B0(n1479), .B1(n15), .A0N(memory[381]), .A1N(n15), .Y(n485) );
  OAI2BB2X1 U811 ( .B0(n1477), .B1(n15), .A0N(memory[382]), .A1N(n15), .Y(n486) );
  OAI2BB2X1 U812 ( .B0(n1475), .B1(n15), .A0N(memory[383]), .A1N(n15), .Y(n487) );
  OAI2BB2X1 U813 ( .B0(n1505), .B1(n16), .A0N(memory[384]), .A1N(n16), .Y(n488) );
  OAI2BB2X1 U814 ( .B0(n1503), .B1(n16), .A0N(memory[385]), .A1N(n16), .Y(n489) );
  OAI2BB2X1 U815 ( .B0(n1501), .B1(n16), .A0N(memory[386]), .A1N(n16), .Y(n490) );
  OAI2BB2X1 U816 ( .B0(n1499), .B1(n16), .A0N(memory[387]), .A1N(n16), .Y(n491) );
  OAI2BB2X1 U817 ( .B0(n1497), .B1(n16), .A0N(memory[388]), .A1N(n16), .Y(n492) );
  OAI2BB2X1 U818 ( .B0(n1495), .B1(n16), .A0N(memory[389]), .A1N(n16), .Y(n493) );
  OAI2BB2X1 U819 ( .B0(n1493), .B1(n16), .A0N(memory[390]), .A1N(n16), .Y(n494) );
  OAI2BB2X1 U820 ( .B0(n1491), .B1(n16), .A0N(memory[391]), .A1N(n16), .Y(n495) );
  OAI2BB2X1 U821 ( .B0(n1481), .B1(n16), .A0N(memory[396]), .A1N(n16), .Y(n500) );
  OAI2BB2X1 U822 ( .B0(n1479), .B1(n16), .A0N(memory[397]), .A1N(n16), .Y(n501) );
  OAI2BB2X1 U823 ( .B0(n1477), .B1(n16), .A0N(memory[398]), .A1N(n16), .Y(n502) );
  OAI2BB2X1 U824 ( .B0(n1475), .B1(n16), .A0N(memory[399]), .A1N(n16), .Y(n503) );
  OAI2BB2X1 U825 ( .B0(n1504), .B1(n17), .A0N(memory[400]), .A1N(n17), .Y(n504) );
  OAI2BB2X1 U826 ( .B0(n1502), .B1(n17), .A0N(memory[401]), .A1N(n17), .Y(n505) );
  OAI2BB2X1 U827 ( .B0(n1500), .B1(n17), .A0N(memory[402]), .A1N(n17), .Y(n506) );
  OAI2BB2X1 U828 ( .B0(n1498), .B1(n17), .A0N(memory[403]), .A1N(n17), .Y(n507) );
  OAI2BB2X1 U829 ( .B0(n1496), .B1(n17), .A0N(memory[404]), .A1N(n17), .Y(n508) );
  OAI2BB2X1 U830 ( .B0(n1494), .B1(n17), .A0N(memory[405]), .A1N(n17), .Y(n509) );
  OAI2BB2X1 U831 ( .B0(n1492), .B1(n17), .A0N(memory[406]), .A1N(n17), .Y(n510) );
  OAI2BB2X1 U832 ( .B0(n1490), .B1(n17), .A0N(memory[407]), .A1N(n17), .Y(n511) );
  OAI2BB2X1 U833 ( .B0(n1480), .B1(n17), .A0N(memory[412]), .A1N(n17), .Y(n516) );
  OAI2BB2X1 U834 ( .B0(n1478), .B1(n17), .A0N(memory[413]), .A1N(n17), .Y(n517) );
  OAI2BB2X1 U835 ( .B0(n1476), .B1(n17), .A0N(memory[414]), .A1N(n17), .Y(n518) );
  OAI2BB2X1 U836 ( .B0(n1474), .B1(n17), .A0N(memory[415]), .A1N(n17), .Y(n519) );
  OAI2BB2X1 U837 ( .B0(n1505), .B1(n76), .A0N(memory[416]), .A1N(n76), .Y(n520) );
  OAI2BB2X1 U838 ( .B0(n1503), .B1(n76), .A0N(memory[417]), .A1N(n76), .Y(n521) );
  OAI2BB2X1 U839 ( .B0(n1501), .B1(n76), .A0N(memory[418]), .A1N(n76), .Y(n522) );
  OAI2BB2X1 U840 ( .B0(n1499), .B1(n76), .A0N(memory[419]), .A1N(n76), .Y(n523) );
  OAI2BB2X1 U841 ( .B0(n1497), .B1(n76), .A0N(memory[420]), .A1N(n76), .Y(n524) );
  OAI2BB2X1 U842 ( .B0(n1495), .B1(n76), .A0N(memory[421]), .A1N(n76), .Y(n525) );
  OAI2BB2X1 U843 ( .B0(n1493), .B1(n76), .A0N(memory[422]), .A1N(n76), .Y(n526) );
  OAI2BB2X1 U844 ( .B0(n1491), .B1(n76), .A0N(memory[423]), .A1N(n76), .Y(n527) );
  OAI2BB2X1 U845 ( .B0(n1481), .B1(n76), .A0N(memory[428]), .A1N(n76), .Y(n532) );
  OAI2BB2X1 U846 ( .B0(n1479), .B1(n76), .A0N(memory[429]), .A1N(n76), .Y(n533) );
  OAI2BB2X1 U847 ( .B0(n1477), .B1(n76), .A0N(memory[430]), .A1N(n76), .Y(n534) );
  OAI2BB2X1 U848 ( .B0(n1475), .B1(n76), .A0N(memory[431]), .A1N(n76), .Y(n535) );
  OAI2BB2X1 U849 ( .B0(n1505), .B1(n18), .A0N(memory[432]), .A1N(n18), .Y(n536) );
  OAI2BB2X1 U850 ( .B0(n1503), .B1(n18), .A0N(memory[433]), .A1N(n18), .Y(n537) );
  OAI2BB2X1 U851 ( .B0(n1501), .B1(n18), .A0N(memory[434]), .A1N(n18), .Y(n538) );
  OAI2BB2X1 U852 ( .B0(n1499), .B1(n18), .A0N(memory[435]), .A1N(n18), .Y(n539) );
  OAI2BB2X1 U853 ( .B0(n1497), .B1(n18), .A0N(memory[436]), .A1N(n18), .Y(n540) );
  OAI2BB2X1 U854 ( .B0(n1495), .B1(n18), .A0N(memory[437]), .A1N(n18), .Y(n541) );
  OAI2BB2X1 U855 ( .B0(n1493), .B1(n18), .A0N(memory[438]), .A1N(n18), .Y(n542) );
  OAI2BB2X1 U856 ( .B0(n1491), .B1(n18), .A0N(memory[439]), .A1N(n18), .Y(n543) );
  OAI2BB2X1 U857 ( .B0(n1481), .B1(n18), .A0N(memory[444]), .A1N(n18), .Y(n548) );
  OAI2BB2X1 U858 ( .B0(n1479), .B1(n18), .A0N(memory[445]), .A1N(n18), .Y(n549) );
  OAI2BB2X1 U859 ( .B0(n1477), .B1(n18), .A0N(memory[446]), .A1N(n18), .Y(n550) );
  OAI2BB2X1 U860 ( .B0(n1475), .B1(n18), .A0N(memory[447]), .A1N(n18), .Y(n551) );
  OAI2BB2X1 U861 ( .B0(n1505), .B1(n78), .A0N(memory[448]), .A1N(n78), .Y(n552) );
  OAI2BB2X1 U862 ( .B0(n1503), .B1(n78), .A0N(memory[449]), .A1N(n78), .Y(n553) );
  OAI2BB2X1 U863 ( .B0(n1501), .B1(n78), .A0N(memory[450]), .A1N(n78), .Y(n554) );
  OAI2BB2X1 U864 ( .B0(n1499), .B1(n78), .A0N(memory[451]), .A1N(n78), .Y(n555) );
  OAI2BB2X1 U865 ( .B0(n1497), .B1(n78), .A0N(memory[452]), .A1N(n78), .Y(n556) );
  OAI2BB2X1 U866 ( .B0(n1495), .B1(n78), .A0N(memory[453]), .A1N(n78), .Y(n557) );
  OAI2BB2X1 U867 ( .B0(n1493), .B1(n78), .A0N(memory[454]), .A1N(n78), .Y(n558) );
  OAI2BB2X1 U868 ( .B0(n1491), .B1(n78), .A0N(memory[455]), .A1N(n78), .Y(n559) );
  OAI2BB2X1 U869 ( .B0(n1481), .B1(n78), .A0N(memory[460]), .A1N(n78), .Y(n564) );
  OAI2BB2X1 U870 ( .B0(n1479), .B1(n78), .A0N(memory[461]), .A1N(n78), .Y(n565) );
  OAI2BB2X1 U871 ( .B0(n1477), .B1(n78), .A0N(memory[462]), .A1N(n78), .Y(n566) );
  OAI2BB2X1 U872 ( .B0(n1475), .B1(n78), .A0N(memory[463]), .A1N(n78), .Y(n567) );
  OAI2BB2X1 U873 ( .B0(n1504), .B1(n19), .A0N(memory[464]), .A1N(n19), .Y(n568) );
  OAI2BB2X1 U874 ( .B0(n1502), .B1(n19), .A0N(memory[465]), .A1N(n19), .Y(n569) );
  OAI2BB2X1 U875 ( .B0(n1500), .B1(n19), .A0N(memory[466]), .A1N(n19), .Y(n570) );
  OAI2BB2X1 U876 ( .B0(n1498), .B1(n19), .A0N(memory[467]), .A1N(n19), .Y(n571) );
  OAI2BB2X1 U877 ( .B0(n1496), .B1(n19), .A0N(memory[468]), .A1N(n19), .Y(n572) );
  OAI2BB2X1 U878 ( .B0(n1494), .B1(n19), .A0N(memory[469]), .A1N(n19), .Y(n573) );
  OAI2BB2X1 U879 ( .B0(n1492), .B1(n19), .A0N(memory[470]), .A1N(n19), .Y(n574) );
  OAI2BB2X1 U880 ( .B0(n1490), .B1(n19), .A0N(memory[471]), .A1N(n19), .Y(n575) );
  OAI2BB2X1 U881 ( .B0(n1480), .B1(n19), .A0N(memory[476]), .A1N(n19), .Y(n580) );
  OAI2BB2X1 U882 ( .B0(n1478), .B1(n19), .A0N(memory[477]), .A1N(n19), .Y(n581) );
  OAI2BB2X1 U883 ( .B0(n1476), .B1(n19), .A0N(memory[478]), .A1N(n19), .Y(n582) );
  OAI2BB2X1 U884 ( .B0(n1474), .B1(n19), .A0N(memory[479]), .A1N(n19), .Y(n583) );
  OAI2BB2X1 U885 ( .B0(n1505), .B1(n79), .A0N(memory[480]), .A1N(n79), .Y(n584) );
  OAI2BB2X1 U886 ( .B0(n1503), .B1(n79), .A0N(memory[481]), .A1N(n79), .Y(n585) );
  OAI2BB2X1 U887 ( .B0(n1501), .B1(n79), .A0N(memory[482]), .A1N(n79), .Y(n586) );
  OAI2BB2X1 U888 ( .B0(n1499), .B1(n79), .A0N(memory[483]), .A1N(n79), .Y(n587) );
  OAI2BB2X1 U889 ( .B0(n1497), .B1(n79), .A0N(memory[484]), .A1N(n79), .Y(n588) );
  OAI2BB2X1 U890 ( .B0(n1495), .B1(n79), .A0N(memory[485]), .A1N(n79), .Y(n589) );
  OAI2BB2X1 U891 ( .B0(n1493), .B1(n79), .A0N(memory[486]), .A1N(n79), .Y(n590) );
  OAI2BB2X1 U892 ( .B0(n1491), .B1(n79), .A0N(memory[487]), .A1N(n79), .Y(n591) );
  OAI2BB2X1 U893 ( .B0(n1481), .B1(n79), .A0N(memory[492]), .A1N(n79), .Y(n596) );
  OAI2BB2X1 U894 ( .B0(n1479), .B1(n79), .A0N(memory[493]), .A1N(n79), .Y(n597) );
  OAI2BB2X1 U895 ( .B0(n1477), .B1(n79), .A0N(memory[494]), .A1N(n79), .Y(n598) );
  OAI2BB2X1 U896 ( .B0(n1475), .B1(n79), .A0N(memory[495]), .A1N(n79), .Y(n599) );
  OAI2BB2X1 U897 ( .B0(n1504), .B1(n20), .A0N(memory[496]), .A1N(n20), .Y(n600) );
  OAI2BB2X1 U898 ( .B0(n1502), .B1(n20), .A0N(memory[497]), .A1N(n20), .Y(n601) );
  OAI2BB2X1 U899 ( .B0(n1500), .B1(n20), .A0N(memory[498]), .A1N(n20), .Y(n602) );
  OAI2BB2X1 U900 ( .B0(n1498), .B1(n20), .A0N(memory[499]), .A1N(n20), .Y(n603) );
  OAI2BB2X1 U901 ( .B0(n1496), .B1(n20), .A0N(memory[500]), .A1N(n20), .Y(n604) );
  OAI2BB2X1 U902 ( .B0(n1494), .B1(n20), .A0N(memory[501]), .A1N(n20), .Y(n605) );
  OAI2BB2X1 U903 ( .B0(n1492), .B1(n20), .A0N(memory[502]), .A1N(n20), .Y(n606) );
  OAI2BB2X1 U904 ( .B0(n1490), .B1(n20), .A0N(memory[503]), .A1N(n20), .Y(n607) );
  OAI2BB2X1 U905 ( .B0(n1480), .B1(n20), .A0N(memory[508]), .A1N(n20), .Y(n612) );
  OAI2BB2X1 U906 ( .B0(n1478), .B1(n20), .A0N(memory[509]), .A1N(n20), .Y(n613) );
  OAI2BB2X1 U907 ( .B0(n1476), .B1(n20), .A0N(memory[510]), .A1N(n20), .Y(n614) );
  OAI2BB2X1 U908 ( .B0(n1474), .B1(n20), .A0N(memory[511]), .A1N(n20), .Y(n615) );
  OAI2BB2X1 U909 ( .B0(n1504), .B1(n21), .A0N(memory[512]), .A1N(n21), .Y(n616) );
  OAI2BB2X1 U910 ( .B0(n1502), .B1(n21), .A0N(memory[513]), .A1N(n21), .Y(n617) );
  OAI2BB2X1 U911 ( .B0(n1500), .B1(n21), .A0N(memory[514]), .A1N(n21), .Y(n618) );
  OAI2BB2X1 U912 ( .B0(n1498), .B1(n21), .A0N(memory[515]), .A1N(n21), .Y(n619) );
  OAI2BB2X1 U913 ( .B0(n1496), .B1(n21), .A0N(memory[516]), .A1N(n21), .Y(n620) );
  OAI2BB2X1 U914 ( .B0(n1494), .B1(n21), .A0N(memory[517]), .A1N(n21), .Y(n621) );
  OAI2BB2X1 U915 ( .B0(n1492), .B1(n21), .A0N(memory[518]), .A1N(n21), .Y(n622) );
  OAI2BB2X1 U916 ( .B0(n1490), .B1(n21), .A0N(memory[519]), .A1N(n21), .Y(n623) );
  OAI2BB2X1 U917 ( .B0(n1480), .B1(n21), .A0N(memory[524]), .A1N(n21), .Y(n628) );
  OAI2BB2X1 U918 ( .B0(n1478), .B1(n21), .A0N(memory[525]), .A1N(n21), .Y(n629) );
  OAI2BB2X1 U919 ( .B0(n1476), .B1(n21), .A0N(memory[526]), .A1N(n21), .Y(n630) );
  OAI2BB2X1 U920 ( .B0(n1474), .B1(n21), .A0N(memory[527]), .A1N(n21), .Y(n631) );
  OAI2BB2X1 U921 ( .B0(n1505), .B1(n22), .A0N(memory[528]), .A1N(n22), .Y(n632) );
  OAI2BB2X1 U922 ( .B0(n1503), .B1(n22), .A0N(memory[529]), .A1N(n22), .Y(n633) );
  OAI2BB2X1 U923 ( .B0(n1501), .B1(n22), .A0N(memory[530]), .A1N(n22), .Y(n634) );
  OAI2BB2X1 U924 ( .B0(n1499), .B1(n22), .A0N(memory[531]), .A1N(n22), .Y(n635) );
  OAI2BB2X1 U925 ( .B0(n1497), .B1(n22), .A0N(memory[532]), .A1N(n22), .Y(n636) );
  OAI2BB2X1 U926 ( .B0(n1495), .B1(n22), .A0N(memory[533]), .A1N(n22), .Y(n637) );
  OAI2BB2X1 U927 ( .B0(n1493), .B1(n22), .A0N(memory[534]), .A1N(n22), .Y(n638) );
  OAI2BB2X1 U928 ( .B0(n1491), .B1(n22), .A0N(memory[535]), .A1N(n22), .Y(n639) );
  OAI2BB2X1 U929 ( .B0(n1481), .B1(n22), .A0N(memory[540]), .A1N(n22), .Y(n644) );
  OAI2BB2X1 U930 ( .B0(n1479), .B1(n22), .A0N(memory[541]), .A1N(n22), .Y(n645) );
  OAI2BB2X1 U931 ( .B0(n1477), .B1(n22), .A0N(memory[542]), .A1N(n22), .Y(n646) );
  OAI2BB2X1 U932 ( .B0(n1475), .B1(n22), .A0N(memory[543]), .A1N(n22), .Y(n647) );
  OAI2BB2X1 U933 ( .B0(n1504), .B1(n25), .A0N(memory[544]), .A1N(n25), .Y(n648) );
  OAI2BB2X1 U934 ( .B0(n1502), .B1(n25), .A0N(memory[545]), .A1N(n25), .Y(n649) );
  OAI2BB2X1 U935 ( .B0(n1500), .B1(n25), .A0N(memory[546]), .A1N(n25), .Y(n650) );
  OAI2BB2X1 U936 ( .B0(n1498), .B1(n25), .A0N(memory[547]), .A1N(n25), .Y(n651) );
  OAI2BB2X1 U937 ( .B0(n1496), .B1(n25), .A0N(memory[548]), .A1N(n25), .Y(n652) );
  OAI2BB2X1 U938 ( .B0(n1494), .B1(n25), .A0N(memory[549]), .A1N(n25), .Y(n653) );
  OAI2BB2X1 U939 ( .B0(n1492), .B1(n25), .A0N(memory[550]), .A1N(n25), .Y(n654) );
  OAI2BB2X1 U940 ( .B0(n1490), .B1(n25), .A0N(memory[551]), .A1N(n25), .Y(n655) );
  OAI2BB2X1 U941 ( .B0(n1480), .B1(n25), .A0N(memory[556]), .A1N(n25), .Y(n660) );
  OAI2BB2X1 U942 ( .B0(n1478), .B1(n25), .A0N(memory[557]), .A1N(n25), .Y(n661) );
  OAI2BB2X1 U943 ( .B0(n1476), .B1(n25), .A0N(memory[558]), .A1N(n25), .Y(n662) );
  OAI2BB2X1 U944 ( .B0(n1474), .B1(n25), .A0N(memory[559]), .A1N(n25), .Y(n663) );
  OAI2BB2X1 U945 ( .B0(n1505), .B1(n27), .A0N(memory[560]), .A1N(n27), .Y(n664) );
  OAI2BB2X1 U946 ( .B0(n1503), .B1(n27), .A0N(memory[561]), .A1N(n27), .Y(n665) );
  OAI2BB2X1 U947 ( .B0(n1501), .B1(n27), .A0N(memory[562]), .A1N(n27), .Y(n666) );
  OAI2BB2X1 U948 ( .B0(n1499), .B1(n27), .A0N(memory[563]), .A1N(n27), .Y(n667) );
  OAI2BB2X1 U949 ( .B0(n1497), .B1(n27), .A0N(memory[564]), .A1N(n27), .Y(n668) );
  OAI2BB2X1 U950 ( .B0(n1495), .B1(n27), .A0N(memory[565]), .A1N(n27), .Y(n669) );
  OAI2BB2X1 U951 ( .B0(n1493), .B1(n27), .A0N(memory[566]), .A1N(n27), .Y(n670) );
  OAI2BB2X1 U952 ( .B0(n1491), .B1(n27), .A0N(memory[567]), .A1N(n27), .Y(n671) );
  OAI2BB2X1 U953 ( .B0(n1481), .B1(n27), .A0N(memory[572]), .A1N(n27), .Y(n676) );
  OAI2BB2X1 U954 ( .B0(n1479), .B1(n27), .A0N(memory[573]), .A1N(n27), .Y(n677) );
  OAI2BB2X1 U955 ( .B0(n1477), .B1(n27), .A0N(memory[574]), .A1N(n27), .Y(n678) );
  OAI2BB2X1 U956 ( .B0(n1475), .B1(n27), .A0N(memory[575]), .A1N(n27), .Y(n679) );
  OAI2BB2X1 U957 ( .B0(n1504), .B1(n29), .A0N(memory[576]), .A1N(n29), .Y(n680) );
  OAI2BB2X1 U958 ( .B0(n1502), .B1(n29), .A0N(memory[577]), .A1N(n29), .Y(n681) );
  OAI2BB2X1 U959 ( .B0(n1500), .B1(n29), .A0N(memory[578]), .A1N(n29), .Y(n682) );
  OAI2BB2X1 U960 ( .B0(n1498), .B1(n29), .A0N(memory[579]), .A1N(n29), .Y(n683) );
  OAI2BB2X1 U961 ( .B0(n1496), .B1(n29), .A0N(memory[580]), .A1N(n29), .Y(n684) );
  OAI2BB2X1 U962 ( .B0(n1494), .B1(n29), .A0N(memory[581]), .A1N(n29), .Y(n685) );
  OAI2BB2X1 U963 ( .B0(n1492), .B1(n29), .A0N(memory[582]), .A1N(n29), .Y(n686) );
  OAI2BB2X1 U964 ( .B0(n1490), .B1(n29), .A0N(memory[583]), .A1N(n29), .Y(n687) );
  OAI2BB2X1 U965 ( .B0(n1480), .B1(n29), .A0N(memory[588]), .A1N(n29), .Y(n692) );
  OAI2BB2X1 U966 ( .B0(n1478), .B1(n29), .A0N(memory[589]), .A1N(n29), .Y(n693) );
  OAI2BB2X1 U967 ( .B0(n1476), .B1(n29), .A0N(memory[590]), .A1N(n29), .Y(n694) );
  OAI2BB2X1 U968 ( .B0(n1474), .B1(n29), .A0N(memory[591]), .A1N(n29), .Y(n695) );
  OAI2BB2X1 U969 ( .B0(n1505), .B1(n31), .A0N(memory[592]), .A1N(n31), .Y(n696) );
  OAI2BB2X1 U970 ( .B0(n1503), .B1(n31), .A0N(memory[593]), .A1N(n31), .Y(n697) );
  OAI2BB2X1 U971 ( .B0(n1501), .B1(n31), .A0N(memory[594]), .A1N(n31), .Y(n698) );
  OAI2BB2X1 U972 ( .B0(n1499), .B1(n31), .A0N(memory[595]), .A1N(n31), .Y(n699) );
  OAI2BB2X1 U973 ( .B0(n1497), .B1(n31), .A0N(memory[596]), .A1N(n31), .Y(n700) );
  OAI2BB2X1 U974 ( .B0(n1495), .B1(n31), .A0N(memory[597]), .A1N(n31), .Y(n701) );
  OAI2BB2X1 U975 ( .B0(n1493), .B1(n31), .A0N(memory[598]), .A1N(n31), .Y(n702) );
  OAI2BB2X1 U976 ( .B0(n1491), .B1(n31), .A0N(memory[599]), .A1N(n31), .Y(n703) );
  OAI2BB2X1 U977 ( .B0(n1481), .B1(n31), .A0N(memory[604]), .A1N(n31), .Y(n708) );
  OAI2BB2X1 U978 ( .B0(n1479), .B1(n31), .A0N(memory[605]), .A1N(n31), .Y(n709) );
  OAI2BB2X1 U979 ( .B0(n1477), .B1(n31), .A0N(memory[606]), .A1N(n31), .Y(n710) );
  OAI2BB2X1 U980 ( .B0(n1475), .B1(n31), .A0N(memory[607]), .A1N(n31), .Y(n711) );
  OAI2BB2X1 U981 ( .B0(n1504), .B1(n33), .A0N(memory[608]), .A1N(n33), .Y(n712) );
  OAI2BB2X1 U982 ( .B0(n1502), .B1(n33), .A0N(memory[609]), .A1N(n33), .Y(n713) );
  OAI2BB2X1 U983 ( .B0(n1500), .B1(n33), .A0N(memory[610]), .A1N(n33), .Y(n714) );
  OAI2BB2X1 U984 ( .B0(n1498), .B1(n33), .A0N(memory[611]), .A1N(n33), .Y(n715) );
  OAI2BB2X1 U985 ( .B0(n1496), .B1(n33), .A0N(memory[612]), .A1N(n33), .Y(n716) );
  OAI2BB2X1 U986 ( .B0(n1494), .B1(n33), .A0N(memory[613]), .A1N(n33), .Y(n717) );
  OAI2BB2X1 U987 ( .B0(n1492), .B1(n33), .A0N(memory[614]), .A1N(n33), .Y(n718) );
  OAI2BB2X1 U988 ( .B0(n1490), .B1(n33), .A0N(memory[615]), .A1N(n33), .Y(n719) );
  OAI2BB2X1 U989 ( .B0(n1480), .B1(n33), .A0N(memory[620]), .A1N(n33), .Y(n724) );
  OAI2BB2X1 U990 ( .B0(n1478), .B1(n33), .A0N(memory[621]), .A1N(n33), .Y(n725) );
  OAI2BB2X1 U991 ( .B0(n1476), .B1(n33), .A0N(memory[622]), .A1N(n33), .Y(n726) );
  OAI2BB2X1 U992 ( .B0(n1474), .B1(n33), .A0N(memory[623]), .A1N(n33), .Y(n727) );
  OAI2BB2X1 U993 ( .B0(n1505), .B1(n35), .A0N(memory[624]), .A1N(n35), .Y(n728) );
  OAI2BB2X1 U994 ( .B0(n1503), .B1(n35), .A0N(memory[625]), .A1N(n35), .Y(n729) );
  OAI2BB2X1 U995 ( .B0(n1501), .B1(n35), .A0N(memory[626]), .A1N(n35), .Y(n730) );
  OAI2BB2X1 U996 ( .B0(n1499), .B1(n35), .A0N(memory[627]), .A1N(n35), .Y(n731) );
  OAI2BB2X1 U997 ( .B0(n1497), .B1(n35), .A0N(memory[628]), .A1N(n35), .Y(n732) );
  OAI2BB2X1 U998 ( .B0(n1495), .B1(n35), .A0N(memory[629]), .A1N(n35), .Y(n733) );
  OAI2BB2X1 U999 ( .B0(n1493), .B1(n35), .A0N(memory[630]), .A1N(n35), .Y(n734) );
  OAI2BB2X1 U1000 ( .B0(n1491), .B1(n35), .A0N(memory[631]), .A1N(n35), .Y(
        n735) );
  OAI2BB2X1 U1001 ( .B0(n1481), .B1(n35), .A0N(memory[636]), .A1N(n35), .Y(
        n740) );
  OAI2BB2X1 U1002 ( .B0(n1479), .B1(n35), .A0N(memory[637]), .A1N(n35), .Y(
        n741) );
  OAI2BB2X1 U1003 ( .B0(n1477), .B1(n35), .A0N(memory[638]), .A1N(n35), .Y(
        n742) );
  OAI2BB2X1 U1004 ( .B0(n1475), .B1(n35), .A0N(memory[639]), .A1N(n35), .Y(
        n743) );
  OAI2BB2X1 U1005 ( .B0(n1504), .B1(n37), .A0N(memory[640]), .A1N(n37), .Y(
        n744) );
  OAI2BB2X1 U1006 ( .B0(n1502), .B1(n37), .A0N(memory[641]), .A1N(n37), .Y(
        n745) );
  OAI2BB2X1 U1007 ( .B0(n1500), .B1(n37), .A0N(memory[642]), .A1N(n37), .Y(
        n746) );
  OAI2BB2X1 U1008 ( .B0(n1498), .B1(n37), .A0N(memory[643]), .A1N(n37), .Y(
        n747) );
  OAI2BB2X1 U1009 ( .B0(n1496), .B1(n37), .A0N(memory[644]), .A1N(n37), .Y(
        n748) );
  OAI2BB2X1 U1010 ( .B0(n1494), .B1(n37), .A0N(memory[645]), .A1N(n37), .Y(
        n749) );
  OAI2BB2X1 U1011 ( .B0(n1492), .B1(n37), .A0N(memory[646]), .A1N(n37), .Y(
        n750) );
  OAI2BB2X1 U1012 ( .B0(n1490), .B1(n37), .A0N(memory[647]), .A1N(n37), .Y(
        n751) );
  OAI2BB2X1 U1013 ( .B0(n1480), .B1(n37), .A0N(memory[652]), .A1N(n37), .Y(
        n756) );
  OAI2BB2X1 U1014 ( .B0(n1478), .B1(n37), .A0N(memory[653]), .A1N(n37), .Y(
        n757) );
  OAI2BB2X1 U1015 ( .B0(n1476), .B1(n37), .A0N(memory[654]), .A1N(n37), .Y(
        n758) );
  OAI2BB2X1 U1016 ( .B0(n1474), .B1(n37), .A0N(memory[655]), .A1N(n37), .Y(
        n759) );
  OAI2BB2X1 U1017 ( .B0(n1505), .B1(n40), .A0N(memory[656]), .A1N(n40), .Y(
        n760) );
  OAI2BB2X1 U1018 ( .B0(n1503), .B1(n40), .A0N(memory[657]), .A1N(n40), .Y(
        n761) );
  OAI2BB2X1 U1019 ( .B0(n1501), .B1(n40), .A0N(memory[658]), .A1N(n40), .Y(
        n762) );
  OAI2BB2X1 U1020 ( .B0(n1499), .B1(n40), .A0N(memory[659]), .A1N(n40), .Y(
        n763) );
  OAI2BB2X1 U1021 ( .B0(n1497), .B1(n40), .A0N(memory[660]), .A1N(n40), .Y(
        n764) );
  OAI2BB2X1 U1022 ( .B0(n1495), .B1(n40), .A0N(memory[661]), .A1N(n40), .Y(
        n765) );
  OAI2BB2X1 U1023 ( .B0(n1493), .B1(n40), .A0N(memory[662]), .A1N(n40), .Y(
        n766) );
  OAI2BB2X1 U1024 ( .B0(n1491), .B1(n40), .A0N(memory[663]), .A1N(n40), .Y(
        n767) );
  OAI2BB2X1 U1025 ( .B0(n1481), .B1(n40), .A0N(memory[668]), .A1N(n40), .Y(
        n772) );
  OAI2BB2X1 U1026 ( .B0(n1479), .B1(n40), .A0N(memory[669]), .A1N(n40), .Y(
        n773) );
  OAI2BB2X1 U1027 ( .B0(n1477), .B1(n40), .A0N(memory[670]), .A1N(n40), .Y(
        n774) );
  OAI2BB2X1 U1028 ( .B0(n1475), .B1(n40), .A0N(memory[671]), .A1N(n40), .Y(
        n775) );
  OAI2BB2X1 U1029 ( .B0(n1504), .B1(n42), .A0N(memory[672]), .A1N(n42), .Y(
        n776) );
  OAI2BB2X1 U1030 ( .B0(n1502), .B1(n42), .A0N(memory[673]), .A1N(n42), .Y(
        n777) );
  OAI2BB2X1 U1031 ( .B0(n1500), .B1(n42), .A0N(memory[674]), .A1N(n42), .Y(
        n778) );
  OAI2BB2X1 U1032 ( .B0(n1498), .B1(n42), .A0N(memory[675]), .A1N(n42), .Y(
        n779) );
  OAI2BB2X1 U1033 ( .B0(n1496), .B1(n42), .A0N(memory[676]), .A1N(n42), .Y(
        n780) );
  OAI2BB2X1 U1034 ( .B0(n1494), .B1(n42), .A0N(memory[677]), .A1N(n42), .Y(
        n781) );
  OAI2BB2X1 U1035 ( .B0(n1492), .B1(n42), .A0N(memory[678]), .A1N(n42), .Y(
        n782) );
  OAI2BB2X1 U1036 ( .B0(n1490), .B1(n42), .A0N(memory[679]), .A1N(n42), .Y(
        n783) );
  OAI2BB2X1 U1037 ( .B0(n1480), .B1(n42), .A0N(memory[684]), .A1N(n42), .Y(
        n788) );
  OAI2BB2X1 U1038 ( .B0(n1478), .B1(n42), .A0N(memory[685]), .A1N(n42), .Y(
        n789) );
  OAI2BB2X1 U1039 ( .B0(n1476), .B1(n42), .A0N(memory[686]), .A1N(n42), .Y(
        n790) );
  OAI2BB2X1 U1040 ( .B0(n1474), .B1(n42), .A0N(memory[687]), .A1N(n42), .Y(
        n791) );
  OAI2BB2X1 U1041 ( .B0(n1504), .B1(n43), .A0N(memory[688]), .A1N(n43), .Y(
        n792) );
  OAI2BB2X1 U1042 ( .B0(n1502), .B1(n43), .A0N(memory[689]), .A1N(n43), .Y(
        n793) );
  OAI2BB2X1 U1043 ( .B0(n1500), .B1(n43), .A0N(memory[690]), .A1N(n43), .Y(
        n794) );
  OAI2BB2X1 U1044 ( .B0(n1498), .B1(n43), .A0N(memory[691]), .A1N(n43), .Y(
        n795) );
  OAI2BB2X1 U1045 ( .B0(n1496), .B1(n43), .A0N(memory[692]), .A1N(n43), .Y(
        n796) );
  OAI2BB2X1 U1046 ( .B0(n1494), .B1(n43), .A0N(memory[693]), .A1N(n43), .Y(
        n797) );
  OAI2BB2X1 U1047 ( .B0(n1492), .B1(n43), .A0N(memory[694]), .A1N(n43), .Y(
        n798) );
  OAI2BB2X1 U1048 ( .B0(n1490), .B1(n43), .A0N(memory[695]), .A1N(n43), .Y(
        n799) );
  OAI2BB2X1 U1049 ( .B0(n1480), .B1(n43), .A0N(memory[700]), .A1N(n43), .Y(
        n804) );
  OAI2BB2X1 U1050 ( .B0(n1478), .B1(n43), .A0N(memory[701]), .A1N(n43), .Y(
        n805) );
  OAI2BB2X1 U1051 ( .B0(n1476), .B1(n43), .A0N(memory[702]), .A1N(n43), .Y(
        n806) );
  OAI2BB2X1 U1052 ( .B0(n1474), .B1(n43), .A0N(memory[703]), .A1N(n43), .Y(
        n807) );
  OAI2BB2X1 U1053 ( .B0(n1504), .B1(n44), .A0N(memory[704]), .A1N(n44), .Y(
        n808) );
  OAI2BB2X1 U1054 ( .B0(n1502), .B1(n44), .A0N(memory[705]), .A1N(n44), .Y(
        n809) );
  OAI2BB2X1 U1055 ( .B0(n1500), .B1(n44), .A0N(memory[706]), .A1N(n44), .Y(
        n810) );
  OAI2BB2X1 U1056 ( .B0(n1498), .B1(n44), .A0N(memory[707]), .A1N(n44), .Y(
        n811) );
  OAI2BB2X1 U1057 ( .B0(n1496), .B1(n44), .A0N(memory[708]), .A1N(n44), .Y(
        n812) );
  OAI2BB2X1 U1058 ( .B0(n1494), .B1(n44), .A0N(memory[709]), .A1N(n44), .Y(
        n813) );
  OAI2BB2X1 U1059 ( .B0(n1492), .B1(n44), .A0N(memory[710]), .A1N(n44), .Y(
        n814) );
  OAI2BB2X1 U1060 ( .B0(n1490), .B1(n44), .A0N(memory[711]), .A1N(n44), .Y(
        n815) );
  OAI2BB2X1 U1061 ( .B0(n1480), .B1(n44), .A0N(memory[716]), .A1N(n44), .Y(
        n820) );
  OAI2BB2X1 U1062 ( .B0(n1478), .B1(n44), .A0N(memory[717]), .A1N(n44), .Y(
        n821) );
  OAI2BB2X1 U1063 ( .B0(n1476), .B1(n44), .A0N(memory[718]), .A1N(n44), .Y(
        n822) );
  OAI2BB2X1 U1064 ( .B0(n1474), .B1(n44), .A0N(memory[719]), .A1N(n44), .Y(
        n823) );
  OAI2BB2X1 U1065 ( .B0(n1504), .B1(n45), .A0N(memory[720]), .A1N(n45), .Y(
        n824) );
  OAI2BB2X1 U1066 ( .B0(n1502), .B1(n45), .A0N(memory[721]), .A1N(n45), .Y(
        n825) );
  OAI2BB2X1 U1067 ( .B0(n1500), .B1(n45), .A0N(memory[722]), .A1N(n45), .Y(
        n826) );
  OAI2BB2X1 U1068 ( .B0(n1498), .B1(n45), .A0N(memory[723]), .A1N(n45), .Y(
        n827) );
  OAI2BB2X1 U1069 ( .B0(n1496), .B1(n45), .A0N(memory[724]), .A1N(n45), .Y(
        n828) );
  OAI2BB2X1 U1070 ( .B0(n1494), .B1(n45), .A0N(memory[725]), .A1N(n45), .Y(
        n829) );
  OAI2BB2X1 U1071 ( .B0(n1492), .B1(n45), .A0N(memory[726]), .A1N(n45), .Y(
        n830) );
  OAI2BB2X1 U1072 ( .B0(n1490), .B1(n45), .A0N(memory[727]), .A1N(n45), .Y(
        n831) );
  OAI2BB2X1 U1073 ( .B0(n1480), .B1(n45), .A0N(memory[732]), .A1N(n45), .Y(
        n836) );
  OAI2BB2X1 U1074 ( .B0(n1478), .B1(n45), .A0N(memory[733]), .A1N(n45), .Y(
        n837) );
  OAI2BB2X1 U1075 ( .B0(n1476), .B1(n45), .A0N(memory[734]), .A1N(n45), .Y(
        n838) );
  OAI2BB2X1 U1076 ( .B0(n1474), .B1(n45), .A0N(memory[735]), .A1N(n45), .Y(
        n839) );
  OAI2BB2X1 U1077 ( .B0(n1505), .B1(n46), .A0N(memory[736]), .A1N(n46), .Y(
        n840) );
  OAI2BB2X1 U1078 ( .B0(n1503), .B1(n46), .A0N(memory[737]), .A1N(n46), .Y(
        n841) );
  OAI2BB2X1 U1079 ( .B0(n1501), .B1(n46), .A0N(memory[738]), .A1N(n46), .Y(
        n842) );
  OAI2BB2X1 U1080 ( .B0(n1499), .B1(n46), .A0N(memory[739]), .A1N(n46), .Y(
        n843) );
  OAI2BB2X1 U1081 ( .B0(n1497), .B1(n46), .A0N(memory[740]), .A1N(n46), .Y(
        n844) );
  OAI2BB2X1 U1082 ( .B0(n1495), .B1(n46), .A0N(memory[741]), .A1N(n46), .Y(
        n845) );
  OAI2BB2X1 U1083 ( .B0(n1493), .B1(n46), .A0N(memory[742]), .A1N(n46), .Y(
        n846) );
  OAI2BB2X1 U1084 ( .B0(n1491), .B1(n46), .A0N(memory[743]), .A1N(n46), .Y(
        n847) );
  OAI2BB2X1 U1085 ( .B0(n1481), .B1(n46), .A0N(memory[748]), .A1N(n46), .Y(
        n852) );
  OAI2BB2X1 U1086 ( .B0(n1479), .B1(n46), .A0N(memory[749]), .A1N(n46), .Y(
        n853) );
  OAI2BB2X1 U1087 ( .B0(n1477), .B1(n46), .A0N(memory[750]), .A1N(n46), .Y(
        n854) );
  OAI2BB2X1 U1088 ( .B0(n1475), .B1(n46), .A0N(memory[751]), .A1N(n46), .Y(
        n855) );
  OAI2BB2X1 U1089 ( .B0(n1504), .B1(n47), .A0N(memory[752]), .A1N(n47), .Y(
        n856) );
  OAI2BB2X1 U1090 ( .B0(n1502), .B1(n47), .A0N(memory[753]), .A1N(n47), .Y(
        n857) );
  OAI2BB2X1 U1091 ( .B0(n1500), .B1(n47), .A0N(memory[754]), .A1N(n47), .Y(
        n858) );
  OAI2BB2X1 U1092 ( .B0(n1498), .B1(n47), .A0N(memory[755]), .A1N(n47), .Y(
        n859) );
  OAI2BB2X1 U1093 ( .B0(n1496), .B1(n47), .A0N(memory[756]), .A1N(n47), .Y(
        n860) );
  OAI2BB2X1 U1094 ( .B0(n1494), .B1(n47), .A0N(memory[757]), .A1N(n47), .Y(
        n861) );
  OAI2BB2X1 U1095 ( .B0(n1492), .B1(n47), .A0N(memory[758]), .A1N(n47), .Y(
        n862) );
  OAI2BB2X1 U1096 ( .B0(n1490), .B1(n47), .A0N(memory[759]), .A1N(n47), .Y(
        n863) );
  OAI2BB2X1 U1097 ( .B0(n1480), .B1(n47), .A0N(memory[764]), .A1N(n47), .Y(
        n868) );
  OAI2BB2X1 U1098 ( .B0(n1478), .B1(n47), .A0N(memory[765]), .A1N(n47), .Y(
        n869) );
  OAI2BB2X1 U1099 ( .B0(n1476), .B1(n47), .A0N(memory[766]), .A1N(n47), .Y(
        n870) );
  OAI2BB2X1 U1100 ( .B0(n1474), .B1(n47), .A0N(memory[767]), .A1N(n47), .Y(
        n871) );
  OAI2BB2X1 U1101 ( .B0(n1505), .B1(n48), .A0N(memory[768]), .A1N(n48), .Y(
        n872) );
  OAI2BB2X1 U1102 ( .B0(n1503), .B1(n48), .A0N(memory[769]), .A1N(n48), .Y(
        n873) );
  OAI2BB2X1 U1103 ( .B0(n1501), .B1(n48), .A0N(memory[770]), .A1N(n48), .Y(
        n874) );
  OAI2BB2X1 U1104 ( .B0(n1499), .B1(n48), .A0N(memory[771]), .A1N(n48), .Y(
        n875) );
  OAI2BB2X1 U1105 ( .B0(n1497), .B1(n48), .A0N(memory[772]), .A1N(n48), .Y(
        n876) );
  OAI2BB2X1 U1106 ( .B0(n1495), .B1(n48), .A0N(memory[773]), .A1N(n48), .Y(
        n877) );
  OAI2BB2X1 U1107 ( .B0(n1493), .B1(n48), .A0N(memory[774]), .A1N(n48), .Y(
        n878) );
  OAI2BB2X1 U1108 ( .B0(n1491), .B1(n48), .A0N(memory[775]), .A1N(n48), .Y(
        n879) );
  OAI2BB2X1 U1109 ( .B0(n1481), .B1(n48), .A0N(memory[780]), .A1N(n48), .Y(
        n884) );
  OAI2BB2X1 U1110 ( .B0(n1479), .B1(n48), .A0N(memory[781]), .A1N(n48), .Y(
        n885) );
  OAI2BB2X1 U1111 ( .B0(n1477), .B1(n48), .A0N(memory[782]), .A1N(n48), .Y(
        n886) );
  OAI2BB2X1 U1112 ( .B0(n1475), .B1(n48), .A0N(memory[783]), .A1N(n48), .Y(
        n887) );
  OAI2BB2X1 U1113 ( .B0(n1504), .B1(n49), .A0N(memory[784]), .A1N(n49), .Y(
        n888) );
  OAI2BB2X1 U1114 ( .B0(n1502), .B1(n49), .A0N(memory[785]), .A1N(n49), .Y(
        n889) );
  OAI2BB2X1 U1115 ( .B0(n1500), .B1(n49), .A0N(memory[786]), .A1N(n49), .Y(
        n890) );
  OAI2BB2X1 U1116 ( .B0(n1498), .B1(n49), .A0N(memory[787]), .A1N(n49), .Y(
        n891) );
  OAI2BB2X1 U1117 ( .B0(n1496), .B1(n49), .A0N(memory[788]), .A1N(n49), .Y(
        n892) );
  OAI2BB2X1 U1118 ( .B0(n1494), .B1(n49), .A0N(memory[789]), .A1N(n49), .Y(
        n893) );
  OAI2BB2X1 U1119 ( .B0(n1492), .B1(n49), .A0N(memory[790]), .A1N(n49), .Y(
        n894) );
  OAI2BB2X1 U1120 ( .B0(n1490), .B1(n49), .A0N(memory[791]), .A1N(n49), .Y(
        n895) );
  OAI2BB2X1 U1121 ( .B0(n1480), .B1(n49), .A0N(memory[796]), .A1N(n49), .Y(
        n900) );
  OAI2BB2X1 U1122 ( .B0(n1478), .B1(n49), .A0N(memory[797]), .A1N(n49), .Y(
        n901) );
  OAI2BB2X1 U1123 ( .B0(n1476), .B1(n49), .A0N(memory[798]), .A1N(n49), .Y(
        n902) );
  OAI2BB2X1 U1124 ( .B0(n1474), .B1(n49), .A0N(memory[799]), .A1N(n49), .Y(
        n903) );
  OAI2BB2X1 U1125 ( .B0(n1505), .B1(n51), .A0N(memory[800]), .A1N(n51), .Y(
        n904) );
  OAI2BB2X1 U1126 ( .B0(n1503), .B1(n51), .A0N(memory[801]), .A1N(n51), .Y(
        n905) );
  OAI2BB2X1 U1127 ( .B0(n1501), .B1(n51), .A0N(memory[802]), .A1N(n51), .Y(
        n906) );
  OAI2BB2X1 U1128 ( .B0(n1499), .B1(n51), .A0N(memory[803]), .A1N(n51), .Y(
        n907) );
  OAI2BB2X1 U1129 ( .B0(n1497), .B1(n51), .A0N(memory[804]), .A1N(n51), .Y(
        n908) );
  OAI2BB2X1 U1130 ( .B0(n1495), .B1(n51), .A0N(memory[805]), .A1N(n51), .Y(
        n909) );
  OAI2BB2X1 U1131 ( .B0(n1493), .B1(n51), .A0N(memory[806]), .A1N(n51), .Y(
        n910) );
  OAI2BB2X1 U1132 ( .B0(n1491), .B1(n51), .A0N(memory[807]), .A1N(n51), .Y(
        n911) );
  OAI2BB2X1 U1133 ( .B0(n1481), .B1(n51), .A0N(memory[812]), .A1N(n51), .Y(
        n916) );
  OAI2BB2X1 U1134 ( .B0(n1479), .B1(n51), .A0N(memory[813]), .A1N(n51), .Y(
        n917) );
  OAI2BB2X1 U1135 ( .B0(n1477), .B1(n51), .A0N(memory[814]), .A1N(n51), .Y(
        n918) );
  OAI2BB2X1 U1136 ( .B0(n1475), .B1(n51), .A0N(memory[815]), .A1N(n51), .Y(
        n919) );
  OAI2BB2X1 U1137 ( .B0(n1504), .B1(n52), .A0N(memory[816]), .A1N(n52), .Y(
        n920) );
  OAI2BB2X1 U1138 ( .B0(n1502), .B1(n52), .A0N(memory[817]), .A1N(n52), .Y(
        n921) );
  OAI2BB2X1 U1139 ( .B0(n1500), .B1(n52), .A0N(memory[818]), .A1N(n52), .Y(
        n922) );
  OAI2BB2X1 U1140 ( .B0(n1498), .B1(n52), .A0N(memory[819]), .A1N(n52), .Y(
        n923) );
  OAI2BB2X1 U1141 ( .B0(n1496), .B1(n52), .A0N(memory[820]), .A1N(n52), .Y(
        n924) );
  OAI2BB2X1 U1142 ( .B0(n1494), .B1(n52), .A0N(memory[821]), .A1N(n52), .Y(
        n925) );
  OAI2BB2X1 U1143 ( .B0(n1492), .B1(n52), .A0N(memory[822]), .A1N(n52), .Y(
        n926) );
  OAI2BB2X1 U1144 ( .B0(n1490), .B1(n52), .A0N(memory[823]), .A1N(n52), .Y(
        n927) );
  OAI2BB2X1 U1145 ( .B0(n1480), .B1(n52), .A0N(memory[828]), .A1N(n52), .Y(
        n932) );
  OAI2BB2X1 U1146 ( .B0(n1478), .B1(n52), .A0N(memory[829]), .A1N(n52), .Y(
        n933) );
  OAI2BB2X1 U1147 ( .B0(n1476), .B1(n52), .A0N(memory[830]), .A1N(n52), .Y(
        n934) );
  OAI2BB2X1 U1148 ( .B0(n1474), .B1(n52), .A0N(memory[831]), .A1N(n52), .Y(
        n935) );
  OAI2BB2X1 U1149 ( .B0(n1504), .B1(n53), .A0N(memory[832]), .A1N(n53), .Y(
        n936) );
  OAI2BB2X1 U1150 ( .B0(n1502), .B1(n53), .A0N(memory[833]), .A1N(n53), .Y(
        n937) );
  OAI2BB2X1 U1151 ( .B0(n1500), .B1(n53), .A0N(memory[834]), .A1N(n53), .Y(
        n938) );
  OAI2BB2X1 U1152 ( .B0(n1498), .B1(n53), .A0N(memory[835]), .A1N(n53), .Y(
        n939) );
  OAI2BB2X1 U1153 ( .B0(n1496), .B1(n53), .A0N(memory[836]), .A1N(n53), .Y(
        n940) );
  OAI2BB2X1 U1154 ( .B0(n1494), .B1(n53), .A0N(memory[837]), .A1N(n53), .Y(
        n941) );
  OAI2BB2X1 U1155 ( .B0(n1492), .B1(n53), .A0N(memory[838]), .A1N(n53), .Y(
        n942) );
  OAI2BB2X1 U1156 ( .B0(n1490), .B1(n53), .A0N(memory[839]), .A1N(n53), .Y(
        n943) );
  OAI2BB2X1 U1157 ( .B0(n1480), .B1(n53), .A0N(memory[844]), .A1N(n53), .Y(
        n948) );
  OAI2BB2X1 U1158 ( .B0(n1478), .B1(n53), .A0N(memory[845]), .A1N(n53), .Y(
        n949) );
  OAI2BB2X1 U1159 ( .B0(n1476), .B1(n53), .A0N(memory[846]), .A1N(n53), .Y(
        n950) );
  OAI2BB2X1 U1160 ( .B0(n1474), .B1(n53), .A0N(memory[847]), .A1N(n53), .Y(
        n951) );
  OAI2BB2X1 U1161 ( .B0(n1504), .B1(n54), .A0N(memory[848]), .A1N(n54), .Y(
        n952) );
  OAI2BB2X1 U1162 ( .B0(n1502), .B1(n54), .A0N(memory[849]), .A1N(n54), .Y(
        n953) );
  OAI2BB2X1 U1163 ( .B0(n1500), .B1(n54), .A0N(memory[850]), .A1N(n54), .Y(
        n954) );
  OAI2BB2X1 U1164 ( .B0(n1498), .B1(n54), .A0N(memory[851]), .A1N(n54), .Y(
        n955) );
  OAI2BB2X1 U1165 ( .B0(n1496), .B1(n54), .A0N(memory[852]), .A1N(n54), .Y(
        n956) );
  OAI2BB2X1 U1166 ( .B0(n1494), .B1(n54), .A0N(memory[853]), .A1N(n54), .Y(
        n957) );
  OAI2BB2X1 U1167 ( .B0(n1492), .B1(n54), .A0N(memory[854]), .A1N(n54), .Y(
        n958) );
  OAI2BB2X1 U1168 ( .B0(n1490), .B1(n54), .A0N(memory[855]), .A1N(n54), .Y(
        n959) );
  OAI2BB2X1 U1169 ( .B0(n1480), .B1(n54), .A0N(memory[860]), .A1N(n54), .Y(
        n964) );
  OAI2BB2X1 U1170 ( .B0(n1478), .B1(n54), .A0N(memory[861]), .A1N(n54), .Y(
        n965) );
  OAI2BB2X1 U1171 ( .B0(n1476), .B1(n54), .A0N(memory[862]), .A1N(n54), .Y(
        n966) );
  OAI2BB2X1 U1172 ( .B0(n1474), .B1(n54), .A0N(memory[863]), .A1N(n54), .Y(
        n967) );
  OAI2BB2X1 U1173 ( .B0(n1504), .B1(n55), .A0N(memory[864]), .A1N(n55), .Y(
        n968) );
  OAI2BB2X1 U1174 ( .B0(n1502), .B1(n55), .A0N(memory[865]), .A1N(n55), .Y(
        n969) );
  OAI2BB2X1 U1175 ( .B0(n1500), .B1(n55), .A0N(memory[866]), .A1N(n55), .Y(
        n970) );
  OAI2BB2X1 U1176 ( .B0(n1498), .B1(n55), .A0N(memory[867]), .A1N(n55), .Y(
        n971) );
  OAI2BB2X1 U1177 ( .B0(n1496), .B1(n55), .A0N(memory[868]), .A1N(n55), .Y(
        n972) );
  OAI2BB2X1 U1178 ( .B0(n1494), .B1(n55), .A0N(memory[869]), .A1N(n55), .Y(
        n973) );
  OAI2BB2X1 U1179 ( .B0(n1492), .B1(n55), .A0N(memory[870]), .A1N(n55), .Y(
        n974) );
  OAI2BB2X1 U1180 ( .B0(n1490), .B1(n55), .A0N(memory[871]), .A1N(n55), .Y(
        n975) );
  OAI2BB2X1 U1181 ( .B0(n1480), .B1(n55), .A0N(memory[876]), .A1N(n55), .Y(
        n980) );
  OAI2BB2X1 U1182 ( .B0(n1478), .B1(n55), .A0N(memory[877]), .A1N(n55), .Y(
        n981) );
  OAI2BB2X1 U1183 ( .B0(n1476), .B1(n55), .A0N(memory[878]), .A1N(n55), .Y(
        n982) );
  OAI2BB2X1 U1184 ( .B0(n1474), .B1(n55), .A0N(memory[879]), .A1N(n55), .Y(
        n983) );
  OAI2BB2X1 U1185 ( .B0(n1504), .B1(n56), .A0N(memory[880]), .A1N(n56), .Y(
        n984) );
  OAI2BB2X1 U1186 ( .B0(n1502), .B1(n56), .A0N(memory[881]), .A1N(n56), .Y(
        n985) );
  OAI2BB2X1 U1187 ( .B0(n1500), .B1(n56), .A0N(memory[882]), .A1N(n56), .Y(
        n986) );
  OAI2BB2X1 U1188 ( .B0(n1498), .B1(n56), .A0N(memory[883]), .A1N(n56), .Y(
        n987) );
  OAI2BB2X1 U1189 ( .B0(n1496), .B1(n56), .A0N(memory[884]), .A1N(n56), .Y(
        n988) );
  OAI2BB2X1 U1190 ( .B0(n1494), .B1(n56), .A0N(memory[885]), .A1N(n56), .Y(
        n989) );
  OAI2BB2X1 U1191 ( .B0(n1492), .B1(n56), .A0N(memory[886]), .A1N(n56), .Y(
        n990) );
  OAI2BB2X1 U1192 ( .B0(n1490), .B1(n56), .A0N(memory[887]), .A1N(n56), .Y(
        n991) );
  OAI2BB2X1 U1193 ( .B0(n1480), .B1(n56), .A0N(memory[892]), .A1N(n56), .Y(
        n996) );
  OAI2BB2X1 U1194 ( .B0(n1478), .B1(n56), .A0N(memory[893]), .A1N(n56), .Y(
        n997) );
  OAI2BB2X1 U1195 ( .B0(n1476), .B1(n56), .A0N(memory[894]), .A1N(n56), .Y(
        n998) );
  OAI2BB2X1 U1196 ( .B0(n1474), .B1(n56), .A0N(memory[895]), .A1N(n56), .Y(
        n999) );
  OAI2BB2X1 U1197 ( .B0(n1504), .B1(n57), .A0N(memory[896]), .A1N(n57), .Y(
        n1000) );
  OAI2BB2X1 U1198 ( .B0(n1502), .B1(n57), .A0N(memory[897]), .A1N(n57), .Y(
        n1001) );
  OAI2BB2X1 U1199 ( .B0(n1500), .B1(n57), .A0N(memory[898]), .A1N(n57), .Y(
        n1002) );
  OAI2BB2X1 U1200 ( .B0(n1498), .B1(n57), .A0N(memory[899]), .A1N(n57), .Y(
        n1003) );
  OAI2BB2X1 U1201 ( .B0(n1496), .B1(n57), .A0N(memory[900]), .A1N(n57), .Y(
        n1004) );
  OAI2BB2X1 U1202 ( .B0(n1494), .B1(n57), .A0N(memory[901]), .A1N(n57), .Y(
        n1005) );
  OAI2BB2X1 U1203 ( .B0(n1492), .B1(n57), .A0N(memory[902]), .A1N(n57), .Y(
        n1006) );
  OAI2BB2X1 U1204 ( .B0(n1490), .B1(n57), .A0N(memory[903]), .A1N(n57), .Y(
        n1007) );
  OAI2BB2X1 U1205 ( .B0(n1480), .B1(n57), .A0N(memory[908]), .A1N(n57), .Y(
        n1012) );
  OAI2BB2X1 U1206 ( .B0(n1478), .B1(n57), .A0N(memory[909]), .A1N(n57), .Y(
        n1013) );
  OAI2BB2X1 U1207 ( .B0(n1476), .B1(n57), .A0N(memory[910]), .A1N(n57), .Y(
        n1014) );
  OAI2BB2X1 U1208 ( .B0(n1474), .B1(n57), .A0N(memory[911]), .A1N(n57), .Y(
        n1015) );
  OAI2BB2X1 U1209 ( .B0(n1504), .B1(n58), .A0N(memory[912]), .A1N(n58), .Y(
        n1016) );
  OAI2BB2X1 U1210 ( .B0(n1502), .B1(n58), .A0N(memory[913]), .A1N(n58), .Y(
        n1017) );
  OAI2BB2X1 U1211 ( .B0(n1500), .B1(n58), .A0N(memory[914]), .A1N(n58), .Y(
        n1018) );
  OAI2BB2X1 U1212 ( .B0(n1498), .B1(n58), .A0N(memory[915]), .A1N(n58), .Y(
        n1019) );
  OAI2BB2X1 U1213 ( .B0(n1496), .B1(n58), .A0N(memory[916]), .A1N(n58), .Y(
        n1020) );
  OAI2BB2X1 U1214 ( .B0(n1494), .B1(n58), .A0N(memory[917]), .A1N(n58), .Y(
        n1021) );
  OAI2BB2X1 U1215 ( .B0(n1492), .B1(n58), .A0N(memory[918]), .A1N(n58), .Y(
        n1022) );
  OAI2BB2X1 U1216 ( .B0(n1490), .B1(n58), .A0N(memory[919]), .A1N(n58), .Y(
        n1023) );
  OAI2BB2X1 U1217 ( .B0(n1480), .B1(n58), .A0N(memory[924]), .A1N(n58), .Y(
        n1028) );
  OAI2BB2X1 U1218 ( .B0(n1478), .B1(n58), .A0N(memory[925]), .A1N(n58), .Y(
        n1029) );
  OAI2BB2X1 U1219 ( .B0(n1476), .B1(n58), .A0N(memory[926]), .A1N(n58), .Y(
        n1030) );
  OAI2BB2X1 U1220 ( .B0(n1474), .B1(n58), .A0N(memory[927]), .A1N(n58), .Y(
        n1031) );
  OAI2BB2X1 U1221 ( .B0(n1504), .B1(n60), .A0N(memory[928]), .A1N(n60), .Y(
        n1032) );
  OAI2BB2X1 U1222 ( .B0(n1502), .B1(n60), .A0N(memory[929]), .A1N(n60), .Y(
        n1033) );
  OAI2BB2X1 U1223 ( .B0(n1500), .B1(n60), .A0N(memory[930]), .A1N(n60), .Y(
        n1034) );
  OAI2BB2X1 U1224 ( .B0(n1498), .B1(n60), .A0N(memory[931]), .A1N(n60), .Y(
        n1035) );
  OAI2BB2X1 U1225 ( .B0(n1496), .B1(n60), .A0N(memory[932]), .A1N(n60), .Y(
        n1036) );
  OAI2BB2X1 U1226 ( .B0(n1494), .B1(n60), .A0N(memory[933]), .A1N(n60), .Y(
        n1037) );
  OAI2BB2X1 U1227 ( .B0(n1492), .B1(n60), .A0N(memory[934]), .A1N(n60), .Y(
        n1038) );
  OAI2BB2X1 U1228 ( .B0(n1490), .B1(n60), .A0N(memory[935]), .A1N(n60), .Y(
        n1039) );
  OAI2BB2X1 U1229 ( .B0(n1480), .B1(n60), .A0N(memory[940]), .A1N(n60), .Y(
        n1044) );
  OAI2BB2X1 U1230 ( .B0(n1478), .B1(n60), .A0N(memory[941]), .A1N(n60), .Y(
        n1045) );
  OAI2BB2X1 U1231 ( .B0(n1476), .B1(n60), .A0N(memory[942]), .A1N(n60), .Y(
        n1046) );
  OAI2BB2X1 U1232 ( .B0(n1474), .B1(n60), .A0N(memory[943]), .A1N(n60), .Y(
        n1047) );
  OAI2BB2X1 U1233 ( .B0(n1504), .B1(n61), .A0N(memory[944]), .A1N(n61), .Y(
        n1048) );
  OAI2BB2X1 U1234 ( .B0(n1502), .B1(n61), .A0N(memory[945]), .A1N(n61), .Y(
        n1049) );
  OAI2BB2X1 U1235 ( .B0(n1500), .B1(n61), .A0N(memory[946]), .A1N(n61), .Y(
        n1050) );
  OAI2BB2X1 U1236 ( .B0(n1498), .B1(n61), .A0N(memory[947]), .A1N(n61), .Y(
        n1051) );
  OAI2BB2X1 U1237 ( .B0(n1496), .B1(n61), .A0N(memory[948]), .A1N(n61), .Y(
        n1052) );
  OAI2BB2X1 U1238 ( .B0(n1494), .B1(n61), .A0N(memory[949]), .A1N(n61), .Y(
        n1053) );
  OAI2BB2X1 U1239 ( .B0(n1492), .B1(n61), .A0N(memory[950]), .A1N(n61), .Y(
        n1054) );
  OAI2BB2X1 U1240 ( .B0(n1490), .B1(n61), .A0N(memory[951]), .A1N(n61), .Y(
        n1055) );
  OAI2BB2X1 U1241 ( .B0(n1480), .B1(n61), .A0N(memory[956]), .A1N(n61), .Y(
        n1060) );
  OAI2BB2X1 U1242 ( .B0(n1478), .B1(n61), .A0N(memory[957]), .A1N(n61), .Y(
        n1061) );
  OAI2BB2X1 U1243 ( .B0(n1476), .B1(n61), .A0N(memory[958]), .A1N(n61), .Y(
        n1062) );
  OAI2BB2X1 U1244 ( .B0(n1474), .B1(n61), .A0N(memory[959]), .A1N(n61), .Y(
        n1063) );
  OAI2BB2X1 U1245 ( .B0(n1504), .B1(n62), .A0N(memory[960]), .A1N(n62), .Y(
        n1064) );
  OAI2BB2X1 U1246 ( .B0(n1502), .B1(n62), .A0N(memory[961]), .A1N(n62), .Y(
        n1065) );
  OAI2BB2X1 U1247 ( .B0(n1500), .B1(n62), .A0N(memory[962]), .A1N(n62), .Y(
        n1066) );
  OAI2BB2X1 U1248 ( .B0(n1498), .B1(n62), .A0N(memory[963]), .A1N(n62), .Y(
        n1067) );
  OAI2BB2X1 U1249 ( .B0(n1496), .B1(n62), .A0N(memory[964]), .A1N(n62), .Y(
        n1068) );
  OAI2BB2X1 U1250 ( .B0(n1494), .B1(n62), .A0N(memory[965]), .A1N(n62), .Y(
        n1069) );
  OAI2BB2X1 U1251 ( .B0(n1492), .B1(n62), .A0N(memory[966]), .A1N(n62), .Y(
        n1070) );
  OAI2BB2X1 U1252 ( .B0(n1490), .B1(n62), .A0N(memory[967]), .A1N(n62), .Y(
        n1071) );
  OAI2BB2X1 U1253 ( .B0(n1480), .B1(n62), .A0N(memory[972]), .A1N(n62), .Y(
        n1076) );
  OAI2BB2X1 U1254 ( .B0(n1478), .B1(n62), .A0N(memory[973]), .A1N(n62), .Y(
        n1077) );
  OAI2BB2X1 U1255 ( .B0(n1476), .B1(n62), .A0N(memory[974]), .A1N(n62), .Y(
        n1078) );
  OAI2BB2X1 U1256 ( .B0(n1474), .B1(n62), .A0N(memory[975]), .A1N(n62), .Y(
        n1079) );
  OAI2BB2X1 U1257 ( .B0(n1504), .B1(n63), .A0N(memory[976]), .A1N(n63), .Y(
        n1080) );
  OAI2BB2X1 U1258 ( .B0(n1502), .B1(n63), .A0N(memory[977]), .A1N(n63), .Y(
        n1081) );
  OAI2BB2X1 U1259 ( .B0(n1500), .B1(n63), .A0N(memory[978]), .A1N(n63), .Y(
        n1082) );
  OAI2BB2X1 U1260 ( .B0(n1498), .B1(n63), .A0N(memory[979]), .A1N(n63), .Y(
        n1083) );
  OAI2BB2X1 U1261 ( .B0(n1496), .B1(n63), .A0N(memory[980]), .A1N(n63), .Y(
        n1084) );
  OAI2BB2X1 U1262 ( .B0(n1494), .B1(n63), .A0N(memory[981]), .A1N(n63), .Y(
        n1085) );
  OAI2BB2X1 U1263 ( .B0(n1492), .B1(n63), .A0N(memory[982]), .A1N(n63), .Y(
        n1086) );
  OAI2BB2X1 U1264 ( .B0(n1490), .B1(n63), .A0N(memory[983]), .A1N(n63), .Y(
        n1087) );
  OAI2BB2X1 U1265 ( .B0(n1480), .B1(n63), .A0N(memory[988]), .A1N(n63), .Y(
        n1092) );
  OAI2BB2X1 U1266 ( .B0(n1478), .B1(n63), .A0N(memory[989]), .A1N(n63), .Y(
        n1093) );
  OAI2BB2X1 U1267 ( .B0(n1476), .B1(n63), .A0N(memory[990]), .A1N(n63), .Y(
        n1094) );
  OAI2BB2X1 U1268 ( .B0(n1474), .B1(n63), .A0N(memory[991]), .A1N(n63), .Y(
        n1095) );
  OAI2BB2X1 U1269 ( .B0(n1504), .B1(n64), .A0N(memory[992]), .A1N(n64), .Y(
        n1096) );
  OAI2BB2X1 U1270 ( .B0(n1502), .B1(n64), .A0N(memory[993]), .A1N(n64), .Y(
        n1097) );
  OAI2BB2X1 U1271 ( .B0(n1500), .B1(n64), .A0N(memory[994]), .A1N(n64), .Y(
        n1098) );
  OAI2BB2X1 U1272 ( .B0(n1498), .B1(n64), .A0N(memory[995]), .A1N(n64), .Y(
        n1099) );
  OAI2BB2X1 U1273 ( .B0(n1496), .B1(n64), .A0N(memory[996]), .A1N(n64), .Y(
        n1100) );
  OAI2BB2X1 U1274 ( .B0(n1494), .B1(n64), .A0N(memory[997]), .A1N(n64), .Y(
        n1101) );
  OAI2BB2X1 U1275 ( .B0(n1492), .B1(n64), .A0N(memory[998]), .A1N(n64), .Y(
        n1102) );
  OAI2BB2X1 U1276 ( .B0(n1490), .B1(n64), .A0N(memory[999]), .A1N(n64), .Y(
        n1103) );
  OAI2BB2X1 U1277 ( .B0(n1480), .B1(n64), .A0N(memory[1004]), .A1N(n64), .Y(
        n1108) );
  OAI2BB2X1 U1278 ( .B0(n1478), .B1(n64), .A0N(memory[1005]), .A1N(n64), .Y(
        n1109) );
  OAI2BB2X1 U1279 ( .B0(n1476), .B1(n64), .A0N(memory[1006]), .A1N(n64), .Y(
        n1110) );
  OAI2BB2X1 U1280 ( .B0(n1474), .B1(n64), .A0N(memory[1007]), .A1N(n64), .Y(
        n1111) );
  OAI2BB2X1 U1281 ( .B0(n1504), .B1(n65), .A0N(memory[1008]), .A1N(n65), .Y(
        n1112) );
  OAI2BB2X1 U1282 ( .B0(n1502), .B1(n65), .A0N(memory[1009]), .A1N(n65), .Y(
        n1113) );
  OAI2BB2X1 U1283 ( .B0(n1500), .B1(n65), .A0N(memory[1010]), .A1N(n65), .Y(
        n1114) );
  OAI2BB2X1 U1284 ( .B0(n1498), .B1(n65), .A0N(memory[1011]), .A1N(n65), .Y(
        n1115) );
  OAI2BB2X1 U1285 ( .B0(n1496), .B1(n65), .A0N(memory[1012]), .A1N(n65), .Y(
        n1116) );
  OAI2BB2X1 U1286 ( .B0(n1494), .B1(n65), .A0N(memory[1013]), .A1N(n65), .Y(
        n1117) );
  OAI2BB2X1 U1287 ( .B0(n1492), .B1(n65), .A0N(memory[1014]), .A1N(n65), .Y(
        n1118) );
  OAI2BB2X1 U1288 ( .B0(n1490), .B1(n65), .A0N(memory[1015]), .A1N(n65), .Y(
        n1119) );
  OAI2BB2X1 U1289 ( .B0(n1480), .B1(n65), .A0N(memory[1020]), .A1N(n65), .Y(
        n1124) );
  OAI2BB2X1 U1290 ( .B0(n1478), .B1(n65), .A0N(memory[1021]), .A1N(n65), .Y(
        n1125) );
  OAI2BB2X1 U1291 ( .B0(n1476), .B1(n65), .A0N(memory[1022]), .A1N(n65), .Y(
        n1126) );
  OAI2BB2X1 U1292 ( .B0(n1474), .B1(n65), .A0N(memory[1023]), .A1N(n65), .Y(
        n1127) );
  OAI2BB2X1 U1293 ( .B0(n1489), .B1(n2), .A0N(memory[24]), .A1N(n2), .Y(n128)
         );
  OAI2BB2X1 U1294 ( .B0(n1487), .B1(n2), .A0N(memory[25]), .A1N(n2), .Y(n129)
         );
  OAI2BB2X1 U1295 ( .B0(n1485), .B1(n2), .A0N(memory[26]), .A1N(n2), .Y(n130)
         );
  OAI2BB2X1 U1296 ( .B0(n1483), .B1(n2), .A0N(memory[27]), .A1N(n2), .Y(n131)
         );
  OAI2BB2X1 U1297 ( .B0(n1488), .B1(n66), .A0N(memory[40]), .A1N(n66), .Y(n144) );
  OAI2BB2X1 U1298 ( .B0(n1486), .B1(n66), .A0N(memory[41]), .A1N(n66), .Y(n145) );
  OAI2BB2X1 U1299 ( .B0(n1484), .B1(n66), .A0N(memory[42]), .A1N(n66), .Y(n146) );
  OAI2BB2X1 U1300 ( .B0(n1482), .B1(n66), .A0N(memory[43]), .A1N(n66), .Y(n147) );
  OAI2BB2X1 U1301 ( .B0(n1489), .B1(n3), .A0N(memory[56]), .A1N(n3), .Y(n160)
         );
  OAI2BB2X1 U1302 ( .B0(n1487), .B1(n3), .A0N(memory[57]), .A1N(n3), .Y(n161)
         );
  OAI2BB2X1 U1303 ( .B0(n1485), .B1(n3), .A0N(memory[58]), .A1N(n3), .Y(n162)
         );
  OAI2BB2X1 U1304 ( .B0(n1483), .B1(n3), .A0N(memory[59]), .A1N(n3), .Y(n163)
         );
  OAI2BB2X1 U1305 ( .B0(n1489), .B1(n67), .A0N(memory[72]), .A1N(n67), .Y(n176) );
  OAI2BB2X1 U1306 ( .B0(n1487), .B1(n67), .A0N(memory[73]), .A1N(n67), .Y(n177) );
  OAI2BB2X1 U1307 ( .B0(n1485), .B1(n67), .A0N(memory[74]), .A1N(n67), .Y(n178) );
  OAI2BB2X1 U1308 ( .B0(n1483), .B1(n67), .A0N(memory[75]), .A1N(n67), .Y(n179) );
  OAI2BB2X1 U1309 ( .B0(n1488), .B1(n4), .A0N(memory[88]), .A1N(n4), .Y(n192)
         );
  OAI2BB2X1 U1310 ( .B0(n1486), .B1(n4), .A0N(memory[89]), .A1N(n4), .Y(n193)
         );
  OAI2BB2X1 U1311 ( .B0(n1484), .B1(n4), .A0N(memory[90]), .A1N(n4), .Y(n194)
         );
  OAI2BB2X1 U1312 ( .B0(n1482), .B1(n4), .A0N(memory[91]), .A1N(n4), .Y(n195)
         );
  OAI2BB2X1 U1313 ( .B0(n1488), .B1(n69), .A0N(memory[104]), .A1N(n69), .Y(
        n208) );
  OAI2BB2X1 U1314 ( .B0(n1486), .B1(n69), .A0N(memory[105]), .A1N(n69), .Y(
        n209) );
  OAI2BB2X1 U1315 ( .B0(n1484), .B1(n69), .A0N(memory[106]), .A1N(n69), .Y(
        n210) );
  OAI2BB2X1 U1316 ( .B0(n1482), .B1(n69), .A0N(memory[107]), .A1N(n69), .Y(
        n211) );
  OAI2BB2X1 U1317 ( .B0(n1489), .B1(n5), .A0N(memory[120]), .A1N(n5), .Y(n224)
         );
  OAI2BB2X1 U1318 ( .B0(n1487), .B1(n5), .A0N(memory[121]), .A1N(n5), .Y(n225)
         );
  OAI2BB2X1 U1319 ( .B0(n1485), .B1(n5), .A0N(memory[122]), .A1N(n5), .Y(n226)
         );
  OAI2BB2X1 U1320 ( .B0(n1483), .B1(n5), .A0N(memory[123]), .A1N(n5), .Y(n227)
         );
  OAI2BB2X1 U1321 ( .B0(n1488), .B1(n6), .A0N(memory[136]), .A1N(n6), .Y(n240)
         );
  OAI2BB2X1 U1322 ( .B0(n1486), .B1(n6), .A0N(memory[137]), .A1N(n6), .Y(n241)
         );
  OAI2BB2X1 U1323 ( .B0(n1484), .B1(n6), .A0N(memory[138]), .A1N(n6), .Y(n242)
         );
  OAI2BB2X1 U1324 ( .B0(n1482), .B1(n6), .A0N(memory[139]), .A1N(n6), .Y(n243)
         );
  OAI2BB2X1 U1325 ( .B0(n1489), .B1(n7), .A0N(memory[152]), .A1N(n7), .Y(n256)
         );
  OAI2BB2X1 U1326 ( .B0(n1487), .B1(n7), .A0N(memory[153]), .A1N(n7), .Y(n257)
         );
  OAI2BB2X1 U1327 ( .B0(n1485), .B1(n7), .A0N(memory[154]), .A1N(n7), .Y(n258)
         );
  OAI2BB2X1 U1328 ( .B0(n1483), .B1(n7), .A0N(memory[155]), .A1N(n7), .Y(n259)
         );
  OAI2BB2X1 U1329 ( .B0(n1488), .B1(n70), .A0N(memory[168]), .A1N(n70), .Y(
        n272) );
  OAI2BB2X1 U1330 ( .B0(n1486), .B1(n70), .A0N(memory[169]), .A1N(n70), .Y(
        n273) );
  OAI2BB2X1 U1331 ( .B0(n1484), .B1(n70), .A0N(memory[170]), .A1N(n70), .Y(
        n274) );
  OAI2BB2X1 U1332 ( .B0(n1482), .B1(n70), .A0N(memory[171]), .A1N(n70), .Y(
        n275) );
  OAI2BB2X1 U1333 ( .B0(n1489), .B1(n8), .A0N(memory[184]), .A1N(n8), .Y(n288)
         );
  OAI2BB2X1 U1334 ( .B0(n1487), .B1(n8), .A0N(memory[185]), .A1N(n8), .Y(n289)
         );
  OAI2BB2X1 U1335 ( .B0(n1485), .B1(n8), .A0N(memory[186]), .A1N(n8), .Y(n290)
         );
  OAI2BB2X1 U1336 ( .B0(n1483), .B1(n8), .A0N(memory[187]), .A1N(n8), .Y(n291)
         );
  OAI2BB2X1 U1337 ( .B0(n1489), .B1(n71), .A0N(memory[200]), .A1N(n71), .Y(
        n304) );
  OAI2BB2X1 U1338 ( .B0(n1487), .B1(n71), .A0N(memory[201]), .A1N(n71), .Y(
        n305) );
  OAI2BB2X1 U1339 ( .B0(n1485), .B1(n71), .A0N(memory[202]), .A1N(n71), .Y(
        n306) );
  OAI2BB2X1 U1340 ( .B0(n1483), .B1(n71), .A0N(memory[203]), .A1N(n71), .Y(
        n307) );
  OAI2BB2X1 U1341 ( .B0(n1489), .B1(n9), .A0N(memory[216]), .A1N(n9), .Y(n320)
         );
  OAI2BB2X1 U1342 ( .B0(n1487), .B1(n9), .A0N(memory[217]), .A1N(n9), .Y(n321)
         );
  OAI2BB2X1 U1343 ( .B0(n1485), .B1(n9), .A0N(memory[218]), .A1N(n9), .Y(n322)
         );
  OAI2BB2X1 U1344 ( .B0(n1483), .B1(n9), .A0N(memory[219]), .A1N(n9), .Y(n323)
         );
  OAI2BB2X1 U1345 ( .B0(n1489), .B1(n72), .A0N(memory[232]), .A1N(n72), .Y(
        n336) );
  OAI2BB2X1 U1346 ( .B0(n1487), .B1(n72), .A0N(memory[233]), .A1N(n72), .Y(
        n337) );
  OAI2BB2X1 U1347 ( .B0(n1485), .B1(n72), .A0N(memory[234]), .A1N(n72), .Y(
        n338) );
  OAI2BB2X1 U1348 ( .B0(n1483), .B1(n72), .A0N(memory[235]), .A1N(n72), .Y(
        n339) );
  OAI2BB2X1 U1349 ( .B0(n1489), .B1(n10), .A0N(memory[248]), .A1N(n10), .Y(
        n352) );
  OAI2BB2X1 U1350 ( .B0(n1487), .B1(n10), .A0N(memory[249]), .A1N(n10), .Y(
        n353) );
  OAI2BB2X1 U1351 ( .B0(n1485), .B1(n10), .A0N(memory[250]), .A1N(n10), .Y(
        n354) );
  OAI2BB2X1 U1352 ( .B0(n1483), .B1(n10), .A0N(memory[251]), .A1N(n10), .Y(
        n355) );
  OAI2BB2X1 U1353 ( .B0(n1489), .B1(n11), .A0N(memory[264]), .A1N(n11), .Y(
        n368) );
  OAI2BB2X1 U1354 ( .B0(n1487), .B1(n11), .A0N(memory[265]), .A1N(n11), .Y(
        n369) );
  OAI2BB2X1 U1355 ( .B0(n1485), .B1(n11), .A0N(memory[266]), .A1N(n11), .Y(
        n370) );
  OAI2BB2X1 U1356 ( .B0(n1483), .B1(n11), .A0N(memory[267]), .A1N(n11), .Y(
        n371) );
  OAI2BB2X1 U1357 ( .B0(n1489), .B1(n12), .A0N(memory[280]), .A1N(n12), .Y(
        n384) );
  OAI2BB2X1 U1358 ( .B0(n1487), .B1(n12), .A0N(memory[281]), .A1N(n12), .Y(
        n385) );
  OAI2BB2X1 U1359 ( .B0(n1485), .B1(n12), .A0N(memory[282]), .A1N(n12), .Y(
        n386) );
  OAI2BB2X1 U1360 ( .B0(n1483), .B1(n12), .A0N(memory[283]), .A1N(n12), .Y(
        n387) );
  OAI2BB2X1 U1361 ( .B0(n1489), .B1(n73), .A0N(memory[296]), .A1N(n73), .Y(
        n400) );
  OAI2BB2X1 U1362 ( .B0(n1487), .B1(n73), .A0N(memory[297]), .A1N(n73), .Y(
        n401) );
  OAI2BB2X1 U1363 ( .B0(n1485), .B1(n73), .A0N(memory[298]), .A1N(n73), .Y(
        n402) );
  OAI2BB2X1 U1364 ( .B0(n1483), .B1(n73), .A0N(memory[299]), .A1N(n73), .Y(
        n403) );
  OAI2BB2X1 U1365 ( .B0(n1489), .B1(n13), .A0N(memory[312]), .A1N(n13), .Y(
        n416) );
  OAI2BB2X1 U1366 ( .B0(n1487), .B1(n13), .A0N(memory[313]), .A1N(n13), .Y(
        n417) );
  OAI2BB2X1 U1367 ( .B0(n1485), .B1(n13), .A0N(memory[314]), .A1N(n13), .Y(
        n418) );
  OAI2BB2X1 U1368 ( .B0(n1483), .B1(n13), .A0N(memory[315]), .A1N(n13), .Y(
        n419) );
  OAI2BB2X1 U1369 ( .B0(n1489), .B1(n74), .A0N(memory[328]), .A1N(n74), .Y(
        n432) );
  OAI2BB2X1 U1370 ( .B0(n1487), .B1(n74), .A0N(memory[329]), .A1N(n74), .Y(
        n433) );
  OAI2BB2X1 U1371 ( .B0(n1485), .B1(n74), .A0N(memory[330]), .A1N(n74), .Y(
        n434) );
  OAI2BB2X1 U1372 ( .B0(n1483), .B1(n74), .A0N(memory[331]), .A1N(n74), .Y(
        n435) );
  OAI2BB2X1 U1373 ( .B0(n1489), .B1(n14), .A0N(memory[344]), .A1N(n14), .Y(
        n448) );
  OAI2BB2X1 U1374 ( .B0(n1487), .B1(n14), .A0N(memory[345]), .A1N(n14), .Y(
        n449) );
  OAI2BB2X1 U1375 ( .B0(n1485), .B1(n14), .A0N(memory[346]), .A1N(n14), .Y(
        n450) );
  OAI2BB2X1 U1376 ( .B0(n1483), .B1(n14), .A0N(memory[347]), .A1N(n14), .Y(
        n451) );
  OAI2BB2X1 U1377 ( .B0(n1489), .B1(n75), .A0N(memory[360]), .A1N(n75), .Y(
        n464) );
  OAI2BB2X1 U1378 ( .B0(n1487), .B1(n75), .A0N(memory[361]), .A1N(n75), .Y(
        n465) );
  OAI2BB2X1 U1379 ( .B0(n1485), .B1(n75), .A0N(memory[362]), .A1N(n75), .Y(
        n466) );
  OAI2BB2X1 U1380 ( .B0(n1483), .B1(n75), .A0N(memory[363]), .A1N(n75), .Y(
        n467) );
  OAI2BB2X1 U1381 ( .B0(n1489), .B1(n15), .A0N(memory[376]), .A1N(n15), .Y(
        n480) );
  OAI2BB2X1 U1382 ( .B0(n1487), .B1(n15), .A0N(memory[377]), .A1N(n15), .Y(
        n481) );
  OAI2BB2X1 U1383 ( .B0(n1485), .B1(n15), .A0N(memory[378]), .A1N(n15), .Y(
        n482) );
  OAI2BB2X1 U1384 ( .B0(n1483), .B1(n15), .A0N(memory[379]), .A1N(n15), .Y(
        n483) );
  OAI2BB2X1 U1385 ( .B0(n1489), .B1(n16), .A0N(memory[392]), .A1N(n16), .Y(
        n496) );
  OAI2BB2X1 U1386 ( .B0(n1487), .B1(n16), .A0N(memory[393]), .A1N(n16), .Y(
        n497) );
  OAI2BB2X1 U1387 ( .B0(n1485), .B1(n16), .A0N(memory[394]), .A1N(n16), .Y(
        n498) );
  OAI2BB2X1 U1388 ( .B0(n1483), .B1(n16), .A0N(memory[395]), .A1N(n16), .Y(
        n499) );
  OAI2BB2X1 U1389 ( .B0(n1488), .B1(n17), .A0N(memory[408]), .A1N(n17), .Y(
        n512) );
  OAI2BB2X1 U1390 ( .B0(n1486), .B1(n17), .A0N(memory[409]), .A1N(n17), .Y(
        n513) );
  OAI2BB2X1 U1391 ( .B0(n1484), .B1(n17), .A0N(memory[410]), .A1N(n17), .Y(
        n514) );
  OAI2BB2X1 U1392 ( .B0(n1482), .B1(n17), .A0N(memory[411]), .A1N(n17), .Y(
        n515) );
  OAI2BB2X1 U1393 ( .B0(n1489), .B1(n76), .A0N(memory[424]), .A1N(n76), .Y(
        n528) );
  OAI2BB2X1 U1394 ( .B0(n1487), .B1(n76), .A0N(memory[425]), .A1N(n76), .Y(
        n529) );
  OAI2BB2X1 U1395 ( .B0(n1485), .B1(n76), .A0N(memory[426]), .A1N(n76), .Y(
        n530) );
  OAI2BB2X1 U1396 ( .B0(n1483), .B1(n76), .A0N(memory[427]), .A1N(n76), .Y(
        n531) );
  OAI2BB2X1 U1397 ( .B0(n1489), .B1(n18), .A0N(memory[440]), .A1N(n18), .Y(
        n544) );
  OAI2BB2X1 U1398 ( .B0(n1487), .B1(n18), .A0N(memory[441]), .A1N(n18), .Y(
        n545) );
  OAI2BB2X1 U1399 ( .B0(n1485), .B1(n18), .A0N(memory[442]), .A1N(n18), .Y(
        n546) );
  OAI2BB2X1 U1400 ( .B0(n1483), .B1(n18), .A0N(memory[443]), .A1N(n18), .Y(
        n547) );
  OAI2BB2X1 U1401 ( .B0(n1489), .B1(n78), .A0N(memory[456]), .A1N(n78), .Y(
        n560) );
  OAI2BB2X1 U1402 ( .B0(n1487), .B1(n78), .A0N(memory[457]), .A1N(n78), .Y(
        n561) );
  OAI2BB2X1 U1403 ( .B0(n1485), .B1(n78), .A0N(memory[458]), .A1N(n78), .Y(
        n562) );
  OAI2BB2X1 U1404 ( .B0(n1483), .B1(n78), .A0N(memory[459]), .A1N(n78), .Y(
        n563) );
  OAI2BB2X1 U1405 ( .B0(n1488), .B1(n19), .A0N(memory[472]), .A1N(n19), .Y(
        n576) );
  OAI2BB2X1 U1406 ( .B0(n1486), .B1(n19), .A0N(memory[473]), .A1N(n19), .Y(
        n577) );
  OAI2BB2X1 U1407 ( .B0(n1484), .B1(n19), .A0N(memory[474]), .A1N(n19), .Y(
        n578) );
  OAI2BB2X1 U1408 ( .B0(n1482), .B1(n19), .A0N(memory[475]), .A1N(n19), .Y(
        n579) );
  OAI2BB2X1 U1409 ( .B0(n1489), .B1(n79), .A0N(memory[488]), .A1N(n79), .Y(
        n592) );
  OAI2BB2X1 U1410 ( .B0(n1487), .B1(n79), .A0N(memory[489]), .A1N(n79), .Y(
        n593) );
  OAI2BB2X1 U1411 ( .B0(n1485), .B1(n79), .A0N(memory[490]), .A1N(n79), .Y(
        n594) );
  OAI2BB2X1 U1412 ( .B0(n1483), .B1(n79), .A0N(memory[491]), .A1N(n79), .Y(
        n595) );
  OAI2BB2X1 U1413 ( .B0(n1488), .B1(n20), .A0N(memory[504]), .A1N(n20), .Y(
        n608) );
  OAI2BB2X1 U1414 ( .B0(n1486), .B1(n20), .A0N(memory[505]), .A1N(n20), .Y(
        n609) );
  OAI2BB2X1 U1415 ( .B0(n1484), .B1(n20), .A0N(memory[506]), .A1N(n20), .Y(
        n610) );
  OAI2BB2X1 U1416 ( .B0(n1482), .B1(n20), .A0N(memory[507]), .A1N(n20), .Y(
        n611) );
  OAI2BB2X1 U1417 ( .B0(n1488), .B1(n21), .A0N(memory[520]), .A1N(n21), .Y(
        n624) );
  OAI2BB2X1 U1418 ( .B0(n1486), .B1(n21), .A0N(memory[521]), .A1N(n21), .Y(
        n625) );
  OAI2BB2X1 U1419 ( .B0(n1484), .B1(n21), .A0N(memory[522]), .A1N(n21), .Y(
        n626) );
  OAI2BB2X1 U1420 ( .B0(n1482), .B1(n21), .A0N(memory[523]), .A1N(n21), .Y(
        n627) );
  OAI2BB2X1 U1421 ( .B0(n1489), .B1(n22), .A0N(memory[536]), .A1N(n22), .Y(
        n640) );
  OAI2BB2X1 U1422 ( .B0(n1487), .B1(n22), .A0N(memory[537]), .A1N(n22), .Y(
        n641) );
  OAI2BB2X1 U1423 ( .B0(n1485), .B1(n22), .A0N(memory[538]), .A1N(n22), .Y(
        n642) );
  OAI2BB2X1 U1424 ( .B0(n1483), .B1(n22), .A0N(memory[539]), .A1N(n22), .Y(
        n643) );
  OAI2BB2X1 U1425 ( .B0(n1488), .B1(n25), .A0N(memory[552]), .A1N(n25), .Y(
        n656) );
  OAI2BB2X1 U1426 ( .B0(n1486), .B1(n25), .A0N(memory[553]), .A1N(n25), .Y(
        n657) );
  OAI2BB2X1 U1427 ( .B0(n1484), .B1(n25), .A0N(memory[554]), .A1N(n25), .Y(
        n658) );
  OAI2BB2X1 U1428 ( .B0(n1482), .B1(n25), .A0N(memory[555]), .A1N(n25), .Y(
        n659) );
  OAI2BB2X1 U1429 ( .B0(n1489), .B1(n27), .A0N(memory[568]), .A1N(n27), .Y(
        n672) );
  OAI2BB2X1 U1430 ( .B0(n1487), .B1(n27), .A0N(memory[569]), .A1N(n27), .Y(
        n673) );
  OAI2BB2X1 U1431 ( .B0(n1485), .B1(n27), .A0N(memory[570]), .A1N(n27), .Y(
        n674) );
  OAI2BB2X1 U1432 ( .B0(n1483), .B1(n27), .A0N(memory[571]), .A1N(n27), .Y(
        n675) );
  OAI2BB2X1 U1433 ( .B0(n1488), .B1(n29), .A0N(memory[584]), .A1N(n29), .Y(
        n688) );
  OAI2BB2X1 U1434 ( .B0(n1486), .B1(n29), .A0N(memory[585]), .A1N(n29), .Y(
        n689) );
  OAI2BB2X1 U1435 ( .B0(n1484), .B1(n29), .A0N(memory[586]), .A1N(n29), .Y(
        n690) );
  OAI2BB2X1 U1436 ( .B0(n1482), .B1(n29), .A0N(memory[587]), .A1N(n29), .Y(
        n691) );
  OAI2BB2X1 U1437 ( .B0(n1489), .B1(n31), .A0N(memory[600]), .A1N(n31), .Y(
        n704) );
  OAI2BB2X1 U1438 ( .B0(n1487), .B1(n31), .A0N(memory[601]), .A1N(n31), .Y(
        n705) );
  OAI2BB2X1 U1439 ( .B0(n1485), .B1(n31), .A0N(memory[602]), .A1N(n31), .Y(
        n706) );
  OAI2BB2X1 U1440 ( .B0(n1483), .B1(n31), .A0N(memory[603]), .A1N(n31), .Y(
        n707) );
  OAI2BB2X1 U1441 ( .B0(n1488), .B1(n33), .A0N(memory[616]), .A1N(n33), .Y(
        n720) );
  OAI2BB2X1 U1442 ( .B0(n1486), .B1(n33), .A0N(memory[617]), .A1N(n33), .Y(
        n721) );
  OAI2BB2X1 U1443 ( .B0(n1484), .B1(n33), .A0N(memory[618]), .A1N(n33), .Y(
        n722) );
  OAI2BB2X1 U1444 ( .B0(n1482), .B1(n33), .A0N(memory[619]), .A1N(n33), .Y(
        n723) );
  OAI2BB2X1 U1445 ( .B0(n1489), .B1(n35), .A0N(memory[632]), .A1N(n35), .Y(
        n736) );
  OAI2BB2X1 U1446 ( .B0(n1487), .B1(n35), .A0N(memory[633]), .A1N(n35), .Y(
        n737) );
  OAI2BB2X1 U1447 ( .B0(n1485), .B1(n35), .A0N(memory[634]), .A1N(n35), .Y(
        n738) );
  OAI2BB2X1 U1448 ( .B0(n1483), .B1(n35), .A0N(memory[635]), .A1N(n35), .Y(
        n739) );
  OAI2BB2X1 U1449 ( .B0(n1488), .B1(n37), .A0N(memory[648]), .A1N(n37), .Y(
        n752) );
  OAI2BB2X1 U1450 ( .B0(n1486), .B1(n37), .A0N(memory[649]), .A1N(n37), .Y(
        n753) );
  OAI2BB2X1 U1451 ( .B0(n1484), .B1(n37), .A0N(memory[650]), .A1N(n37), .Y(
        n754) );
  OAI2BB2X1 U1452 ( .B0(n1482), .B1(n37), .A0N(memory[651]), .A1N(n37), .Y(
        n755) );
  OAI2BB2X1 U1453 ( .B0(n1489), .B1(n40), .A0N(memory[664]), .A1N(n40), .Y(
        n768) );
  OAI2BB2X1 U1454 ( .B0(n1487), .B1(n40), .A0N(memory[665]), .A1N(n40), .Y(
        n769) );
  OAI2BB2X1 U1455 ( .B0(n1485), .B1(n40), .A0N(memory[666]), .A1N(n40), .Y(
        n770) );
  OAI2BB2X1 U1456 ( .B0(n1483), .B1(n40), .A0N(memory[667]), .A1N(n40), .Y(
        n771) );
  OAI2BB2X1 U1457 ( .B0(n1488), .B1(n42), .A0N(memory[680]), .A1N(n42), .Y(
        n784) );
  OAI2BB2X1 U1458 ( .B0(n1486), .B1(n42), .A0N(memory[681]), .A1N(n42), .Y(
        n785) );
  OAI2BB2X1 U1459 ( .B0(n1484), .B1(n42), .A0N(memory[682]), .A1N(n42), .Y(
        n786) );
  OAI2BB2X1 U1460 ( .B0(n1482), .B1(n42), .A0N(memory[683]), .A1N(n42), .Y(
        n787) );
  OAI2BB2X1 U1461 ( .B0(n1488), .B1(n43), .A0N(memory[696]), .A1N(n43), .Y(
        n800) );
  OAI2BB2X1 U1462 ( .B0(n1486), .B1(n43), .A0N(memory[697]), .A1N(n43), .Y(
        n801) );
  OAI2BB2X1 U1463 ( .B0(n1484), .B1(n43), .A0N(memory[698]), .A1N(n43), .Y(
        n802) );
  OAI2BB2X1 U1464 ( .B0(n1482), .B1(n43), .A0N(memory[699]), .A1N(n43), .Y(
        n803) );
  OAI2BB2X1 U1465 ( .B0(n1488), .B1(n44), .A0N(memory[712]), .A1N(n44), .Y(
        n816) );
  OAI2BB2X1 U1466 ( .B0(n1486), .B1(n44), .A0N(memory[713]), .A1N(n44), .Y(
        n817) );
  OAI2BB2X1 U1467 ( .B0(n1484), .B1(n44), .A0N(memory[714]), .A1N(n44), .Y(
        n818) );
  OAI2BB2X1 U1468 ( .B0(n1482), .B1(n44), .A0N(memory[715]), .A1N(n44), .Y(
        n819) );
  OAI2BB2X1 U1469 ( .B0(n1488), .B1(n45), .A0N(memory[728]), .A1N(n45), .Y(
        n832) );
  OAI2BB2X1 U1470 ( .B0(n1486), .B1(n45), .A0N(memory[729]), .A1N(n45), .Y(
        n833) );
  OAI2BB2X1 U1471 ( .B0(n1484), .B1(n45), .A0N(memory[730]), .A1N(n45), .Y(
        n834) );
  OAI2BB2X1 U1472 ( .B0(n1482), .B1(n45), .A0N(memory[731]), .A1N(n45), .Y(
        n835) );
  OAI2BB2X1 U1473 ( .B0(n1489), .B1(n46), .A0N(memory[744]), .A1N(n46), .Y(
        n848) );
  OAI2BB2X1 U1474 ( .B0(n1487), .B1(n46), .A0N(memory[745]), .A1N(n46), .Y(
        n849) );
  OAI2BB2X1 U1475 ( .B0(n1485), .B1(n46), .A0N(memory[746]), .A1N(n46), .Y(
        n850) );
  OAI2BB2X1 U1476 ( .B0(n1483), .B1(n46), .A0N(memory[747]), .A1N(n46), .Y(
        n851) );
  OAI2BB2X1 U1477 ( .B0(n1488), .B1(n47), .A0N(memory[760]), .A1N(n47), .Y(
        n864) );
  OAI2BB2X1 U1478 ( .B0(n1486), .B1(n47), .A0N(memory[761]), .A1N(n47), .Y(
        n865) );
  OAI2BB2X1 U1479 ( .B0(n1484), .B1(n47), .A0N(memory[762]), .A1N(n47), .Y(
        n866) );
  OAI2BB2X1 U1480 ( .B0(n1482), .B1(n47), .A0N(memory[763]), .A1N(n47), .Y(
        n867) );
  OAI2BB2X1 U1481 ( .B0(n1489), .B1(n48), .A0N(memory[776]), .A1N(n48), .Y(
        n880) );
  OAI2BB2X1 U1482 ( .B0(n1487), .B1(n48), .A0N(memory[777]), .A1N(n48), .Y(
        n881) );
  OAI2BB2X1 U1483 ( .B0(n1485), .B1(n48), .A0N(memory[778]), .A1N(n48), .Y(
        n882) );
  OAI2BB2X1 U1484 ( .B0(n1483), .B1(n48), .A0N(memory[779]), .A1N(n48), .Y(
        n883) );
  OAI2BB2X1 U1485 ( .B0(n1488), .B1(n49), .A0N(memory[792]), .A1N(n49), .Y(
        n896) );
  OAI2BB2X1 U1486 ( .B0(n1486), .B1(n49), .A0N(memory[793]), .A1N(n49), .Y(
        n897) );
  OAI2BB2X1 U1487 ( .B0(n1484), .B1(n49), .A0N(memory[794]), .A1N(n49), .Y(
        n898) );
  OAI2BB2X1 U1488 ( .B0(n1482), .B1(n49), .A0N(memory[795]), .A1N(n49), .Y(
        n899) );
  OAI2BB2X1 U1489 ( .B0(n1489), .B1(n51), .A0N(memory[808]), .A1N(n51), .Y(
        n912) );
  OAI2BB2X1 U1490 ( .B0(n1487), .B1(n51), .A0N(memory[809]), .A1N(n51), .Y(
        n913) );
  OAI2BB2X1 U1491 ( .B0(n1485), .B1(n51), .A0N(memory[810]), .A1N(n51), .Y(
        n914) );
  OAI2BB2X1 U1492 ( .B0(n1483), .B1(n51), .A0N(memory[811]), .A1N(n51), .Y(
        n915) );
  OAI2BB2X1 U1493 ( .B0(n1488), .B1(n52), .A0N(memory[824]), .A1N(n52), .Y(
        n928) );
  OAI2BB2X1 U1494 ( .B0(n1486), .B1(n52), .A0N(memory[825]), .A1N(n52), .Y(
        n929) );
  OAI2BB2X1 U1495 ( .B0(n1484), .B1(n52), .A0N(memory[826]), .A1N(n52), .Y(
        n930) );
  OAI2BB2X1 U1496 ( .B0(n1482), .B1(n52), .A0N(memory[827]), .A1N(n52), .Y(
        n931) );
  OAI2BB2X1 U1497 ( .B0(n1488), .B1(n53), .A0N(memory[840]), .A1N(n53), .Y(
        n944) );
  OAI2BB2X1 U1498 ( .B0(n1486), .B1(n53), .A0N(memory[841]), .A1N(n53), .Y(
        n945) );
  OAI2BB2X1 U1499 ( .B0(n1484), .B1(n53), .A0N(memory[842]), .A1N(n53), .Y(
        n946) );
  OAI2BB2X1 U1500 ( .B0(n1482), .B1(n53), .A0N(memory[843]), .A1N(n53), .Y(
        n947) );
  OAI2BB2X1 U1501 ( .B0(n1488), .B1(n54), .A0N(memory[856]), .A1N(n54), .Y(
        n960) );
  OAI2BB2X1 U1502 ( .B0(n1486), .B1(n54), .A0N(memory[857]), .A1N(n54), .Y(
        n961) );
  OAI2BB2X1 U1503 ( .B0(n1484), .B1(n54), .A0N(memory[858]), .A1N(n54), .Y(
        n962) );
  OAI2BB2X1 U1504 ( .B0(n1482), .B1(n54), .A0N(memory[859]), .A1N(n54), .Y(
        n963) );
  OAI2BB2X1 U1505 ( .B0(n1488), .B1(n55), .A0N(memory[872]), .A1N(n55), .Y(
        n976) );
  OAI2BB2X1 U1506 ( .B0(n1486), .B1(n55), .A0N(memory[873]), .A1N(n55), .Y(
        n977) );
  OAI2BB2X1 U1507 ( .B0(n1484), .B1(n55), .A0N(memory[874]), .A1N(n55), .Y(
        n978) );
  OAI2BB2X1 U1508 ( .B0(n1482), .B1(n55), .A0N(memory[875]), .A1N(n55), .Y(
        n979) );
  OAI2BB2X1 U1509 ( .B0(n1488), .B1(n56), .A0N(memory[888]), .A1N(n56), .Y(
        n992) );
  OAI2BB2X1 U1510 ( .B0(n1486), .B1(n56), .A0N(memory[889]), .A1N(n56), .Y(
        n993) );
  OAI2BB2X1 U1511 ( .B0(n1484), .B1(n56), .A0N(memory[890]), .A1N(n56), .Y(
        n994) );
  OAI2BB2X1 U1512 ( .B0(n1482), .B1(n56), .A0N(memory[891]), .A1N(n56), .Y(
        n995) );
  OAI2BB2X1 U1513 ( .B0(n1488), .B1(n57), .A0N(memory[904]), .A1N(n57), .Y(
        n1008) );
  OAI2BB2X1 U1514 ( .B0(n1486), .B1(n57), .A0N(memory[905]), .A1N(n57), .Y(
        n1009) );
  OAI2BB2X1 U1515 ( .B0(n1484), .B1(n57), .A0N(memory[906]), .A1N(n57), .Y(
        n1010) );
  OAI2BB2X1 U1516 ( .B0(n1482), .B1(n57), .A0N(memory[907]), .A1N(n57), .Y(
        n1011) );
  OAI2BB2X1 U1517 ( .B0(n1488), .B1(n58), .A0N(memory[920]), .A1N(n58), .Y(
        n1024) );
  OAI2BB2X1 U1518 ( .B0(n1486), .B1(n58), .A0N(memory[921]), .A1N(n58), .Y(
        n1025) );
  OAI2BB2X1 U1519 ( .B0(n1484), .B1(n58), .A0N(memory[922]), .A1N(n58), .Y(
        n1026) );
  OAI2BB2X1 U1520 ( .B0(n1482), .B1(n58), .A0N(memory[923]), .A1N(n58), .Y(
        n1027) );
  OAI2BB2X1 U1521 ( .B0(n1488), .B1(n60), .A0N(memory[936]), .A1N(n60), .Y(
        n1040) );
  OAI2BB2X1 U1522 ( .B0(n1486), .B1(n60), .A0N(memory[937]), .A1N(n60), .Y(
        n1041) );
  OAI2BB2X1 U1523 ( .B0(n1484), .B1(n60), .A0N(memory[938]), .A1N(n60), .Y(
        n1042) );
  OAI2BB2X1 U1524 ( .B0(n1482), .B1(n60), .A0N(memory[939]), .A1N(n60), .Y(
        n1043) );
  OAI2BB2X1 U1525 ( .B0(n1488), .B1(n61), .A0N(memory[952]), .A1N(n61), .Y(
        n1056) );
  OAI2BB2X1 U1526 ( .B0(n1486), .B1(n61), .A0N(memory[953]), .A1N(n61), .Y(
        n1057) );
  OAI2BB2X1 U1527 ( .B0(n1484), .B1(n61), .A0N(memory[954]), .A1N(n61), .Y(
        n1058) );
  OAI2BB2X1 U1528 ( .B0(n1482), .B1(n61), .A0N(memory[955]), .A1N(n61), .Y(
        n1059) );
  OAI2BB2X1 U1529 ( .B0(n1488), .B1(n62), .A0N(memory[968]), .A1N(n62), .Y(
        n1072) );
  OAI2BB2X1 U1530 ( .B0(n1486), .B1(n62), .A0N(memory[969]), .A1N(n62), .Y(
        n1073) );
  OAI2BB2X1 U1531 ( .B0(n1484), .B1(n62), .A0N(memory[970]), .A1N(n62), .Y(
        n1074) );
  OAI2BB2X1 U1532 ( .B0(n1482), .B1(n62), .A0N(memory[971]), .A1N(n62), .Y(
        n1075) );
  OAI2BB2X1 U1533 ( .B0(n1488), .B1(n63), .A0N(memory[984]), .A1N(n63), .Y(
        n1088) );
  OAI2BB2X1 U1534 ( .B0(n1486), .B1(n63), .A0N(memory[985]), .A1N(n63), .Y(
        n1089) );
  OAI2BB2X1 U1535 ( .B0(n1484), .B1(n63), .A0N(memory[986]), .A1N(n63), .Y(
        n1090) );
  OAI2BB2X1 U1536 ( .B0(n1482), .B1(n63), .A0N(memory[987]), .A1N(n63), .Y(
        n1091) );
  OAI2BB2X1 U1537 ( .B0(n1488), .B1(n64), .A0N(memory[1000]), .A1N(n64), .Y(
        n1104) );
  OAI2BB2X1 U1538 ( .B0(n1486), .B1(n64), .A0N(memory[1001]), .A1N(n64), .Y(
        n1105) );
  OAI2BB2X1 U1539 ( .B0(n1484), .B1(n64), .A0N(memory[1002]), .A1N(n64), .Y(
        n1106) );
  OAI2BB2X1 U1540 ( .B0(n1482), .B1(n64), .A0N(memory[1003]), .A1N(n64), .Y(
        n1107) );
  OAI2BB2X1 U1541 ( .B0(n1488), .B1(n65), .A0N(memory[1016]), .A1N(n65), .Y(
        n1120) );
  OAI2BB2X1 U1542 ( .B0(n1486), .B1(n65), .A0N(memory[1017]), .A1N(n65), .Y(
        n1121) );
  OAI2BB2X1 U1543 ( .B0(n1484), .B1(n65), .A0N(memory[1018]), .A1N(n65), .Y(
        n1122) );
  OAI2BB2X1 U1544 ( .B0(n1482), .B1(n65), .A0N(memory[1019]), .A1N(n65), .Y(
        n1123) );
  BUFX3 U1545 ( .A(addr[5]), .Y(n1511) );
endmodule


module mem8x8_1 ( clk, rstn, en, wr_rd, addr, din, dout );
  input [5:0] addr;
  input [15:0] din;
  output [15:0] dout;
  input clk, rstn, en, wr_rd;
  wire   N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98,
         N99, N100, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n25, n27, n29, n31, n33,
         n35, n37, n40, n42, n43, n44, n45, n46, n47, n48, n49, n51, n52, n53,
         n54, n55, n56, n57, n58, n60, n61, n62, n63, n64, n65, n66, n67, n69,
         n70, n71, n72, n73, n74, n75, n76, n78, n79, n80, n81, n82, n83, n84,
         n85, n87, n88, n89, n90, n91, n92, n93, n94, n96, n97, n98, n99, n100,
         n101, n102, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
         n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
         n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
         n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
         n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
         n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
         n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
         n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
         n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
         n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
         n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
         n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
         n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
         n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
         n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
         n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
         n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
         n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
         n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
         n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
         n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
         n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
         n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
         n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
         n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
         n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
         n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
         n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
         n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
         n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
         n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
         n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
         n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
         n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
         n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495,
         n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
         n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
         n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
         n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
         n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545,
         n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555,
         n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565,
         n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575,
         n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585,
         n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595,
         n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605,
         n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615,
         n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
         n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
         n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
         n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
         n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
         n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
         n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
         n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695,
         n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
         n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715,
         n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725,
         n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735,
         n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745,
         n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755,
         n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765,
         n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775,
         n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785,
         n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795,
         n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805,
         n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815,
         n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825,
         n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835,
         n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845,
         n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855,
         n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865,
         n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875,
         n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885,
         n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895,
         n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905,
         n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915,
         n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925,
         n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935,
         n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945,
         n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955,
         n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965,
         n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975,
         n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985,
         n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995,
         n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005,
         n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015,
         n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025,
         n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035,
         n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045,
         n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055,
         n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065,
         n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075,
         n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085,
         n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095,
         n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105,
         n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115,
         n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125,
         n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135,
         n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145,
         n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155,
         n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165,
         n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175,
         n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185,
         n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195,
         n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205,
         n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215,
         n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225,
         n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
         n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
         n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
         n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265,
         n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275,
         n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285,
         n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295,
         n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305,
         n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315,
         n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325,
         n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335,
         n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345,
         n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355,
         n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365,
         n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375,
         n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385,
         n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395,
         n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405,
         n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415,
         n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425,
         n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435,
         n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445,
         n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455,
         n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465,
         n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475,
         n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485,
         n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495,
         n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505,
         n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515,
         n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525,
         n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535,
         n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545,
         n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553;
  wire   [1023:0] memory;

  DFFRHQX1 memory_reg_1__15_ ( .D(n1528), .CK(clk), .RN(rstn), .Q(memory[1007]) );
  DFFRHQX1 memory_reg_1__14_ ( .D(n1529), .CK(clk), .RN(rstn), .Q(memory[1006]) );
  DFFRHQX1 memory_reg_1__13_ ( .D(n1530), .CK(clk), .RN(rstn), .Q(memory[1005]) );
  DFFRHQX1 memory_reg_1__12_ ( .D(n1531), .CK(clk), .RN(rstn), .Q(memory[1004]) );
  DFFRHQX1 memory_reg_1__11_ ( .D(n1532), .CK(clk), .RN(rstn), .Q(memory[1003]) );
  DFFRHQX1 memory_reg_1__10_ ( .D(n1533), .CK(clk), .RN(rstn), .Q(memory[1002]) );
  DFFRHQX1 memory_reg_1__9_ ( .D(n1534), .CK(clk), .RN(rstn), .Q(memory[1001])
         );
  DFFRHQX1 memory_reg_1__8_ ( .D(n1535), .CK(clk), .RN(rstn), .Q(memory[1000])
         );
  DFFRHQX1 memory_reg_1__7_ ( .D(n1536), .CK(clk), .RN(rstn), .Q(memory[999])
         );
  DFFRHQX1 memory_reg_1__6_ ( .D(n1537), .CK(clk), .RN(rstn), .Q(memory[998])
         );
  DFFRHQX1 memory_reg_1__5_ ( .D(n1538), .CK(clk), .RN(rstn), .Q(memory[997])
         );
  DFFRHQX1 memory_reg_1__4_ ( .D(n1539), .CK(clk), .RN(rstn), .Q(memory[996])
         );
  DFFRHQX1 memory_reg_1__3_ ( .D(n1540), .CK(clk), .RN(rstn), .Q(memory[995])
         );
  DFFRHQX1 memory_reg_1__2_ ( .D(n1541), .CK(clk), .RN(rstn), .Q(memory[994])
         );
  DFFRHQX1 memory_reg_1__1_ ( .D(n1542), .CK(clk), .RN(rstn), .Q(memory[993])
         );
  DFFRHQX1 memory_reg_1__0_ ( .D(n1543), .CK(clk), .RN(rstn), .Q(memory[992])
         );
  DFFRHQX1 memory_reg_5__15_ ( .D(n1592), .CK(clk), .RN(rstn), .Q(memory[943])
         );
  DFFRHQX1 memory_reg_5__14_ ( .D(n1593), .CK(clk), .RN(rstn), .Q(memory[942])
         );
  DFFRHQX1 memory_reg_5__13_ ( .D(n1594), .CK(clk), .RN(rstn), .Q(memory[941])
         );
  DFFRHQX1 memory_reg_5__12_ ( .D(n1595), .CK(clk), .RN(rstn), .Q(memory[940])
         );
  DFFRHQX1 memory_reg_5__11_ ( .D(n1596), .CK(clk), .RN(rstn), .Q(memory[939])
         );
  DFFRHQX1 memory_reg_5__10_ ( .D(n1597), .CK(clk), .RN(rstn), .Q(memory[938])
         );
  DFFRHQX1 memory_reg_5__9_ ( .D(n1598), .CK(clk), .RN(rstn), .Q(memory[937])
         );
  DFFRHQX1 memory_reg_5__8_ ( .D(n1599), .CK(clk), .RN(rstn), .Q(memory[936])
         );
  DFFRHQX1 memory_reg_5__7_ ( .D(n1600), .CK(clk), .RN(rstn), .Q(memory[935])
         );
  DFFRHQX1 memory_reg_5__6_ ( .D(n1601), .CK(clk), .RN(rstn), .Q(memory[934])
         );
  DFFRHQX1 memory_reg_5__5_ ( .D(n1602), .CK(clk), .RN(rstn), .Q(memory[933])
         );
  DFFRHQX1 memory_reg_5__4_ ( .D(n1603), .CK(clk), .RN(rstn), .Q(memory[932])
         );
  DFFRHQX1 memory_reg_5__3_ ( .D(n1604), .CK(clk), .RN(rstn), .Q(memory[931])
         );
  DFFRHQX1 memory_reg_5__2_ ( .D(n1605), .CK(clk), .RN(rstn), .Q(memory[930])
         );
  DFFRHQX1 memory_reg_5__1_ ( .D(n1606), .CK(clk), .RN(rstn), .Q(memory[929])
         );
  DFFRHQX1 memory_reg_5__0_ ( .D(n1607), .CK(clk), .RN(rstn), .Q(memory[928])
         );
  DFFRHQX1 memory_reg_9__15_ ( .D(n1656), .CK(clk), .RN(rstn), .Q(memory[879])
         );
  DFFRHQX1 memory_reg_9__14_ ( .D(n1657), .CK(clk), .RN(rstn), .Q(memory[878])
         );
  DFFRHQX1 memory_reg_9__13_ ( .D(n1658), .CK(clk), .RN(rstn), .Q(memory[877])
         );
  DFFRHQX1 memory_reg_9__12_ ( .D(n1659), .CK(clk), .RN(rstn), .Q(memory[876])
         );
  DFFRHQX1 memory_reg_9__11_ ( .D(n1660), .CK(clk), .RN(rstn), .Q(memory[875])
         );
  DFFRHQX1 memory_reg_9__10_ ( .D(n1661), .CK(clk), .RN(rstn), .Q(memory[874])
         );
  DFFRHQX1 memory_reg_9__9_ ( .D(n1662), .CK(clk), .RN(rstn), .Q(memory[873])
         );
  DFFRHQX1 memory_reg_9__8_ ( .D(n1663), .CK(clk), .RN(rstn), .Q(memory[872])
         );
  DFFRHQX1 memory_reg_9__7_ ( .D(n1664), .CK(clk), .RN(rstn), .Q(memory[871])
         );
  DFFRHQX1 memory_reg_9__6_ ( .D(n1665), .CK(clk), .RN(rstn), .Q(memory[870])
         );
  DFFRHQX1 memory_reg_9__5_ ( .D(n1666), .CK(clk), .RN(rstn), .Q(memory[869])
         );
  DFFRHQX1 memory_reg_9__4_ ( .D(n1667), .CK(clk), .RN(rstn), .Q(memory[868])
         );
  DFFRHQX1 memory_reg_9__3_ ( .D(n1668), .CK(clk), .RN(rstn), .Q(memory[867])
         );
  DFFRHQX1 memory_reg_9__2_ ( .D(n1669), .CK(clk), .RN(rstn), .Q(memory[866])
         );
  DFFRHQX1 memory_reg_9__1_ ( .D(n1670), .CK(clk), .RN(rstn), .Q(memory[865])
         );
  DFFRHQX1 memory_reg_9__0_ ( .D(n1671), .CK(clk), .RN(rstn), .Q(memory[864])
         );
  DFFRHQX1 memory_reg_13__15_ ( .D(n1720), .CK(clk), .RN(rstn), .Q(memory[815]) );
  DFFRHQX1 memory_reg_13__14_ ( .D(n1721), .CK(clk), .RN(rstn), .Q(memory[814]) );
  DFFRHQX1 memory_reg_13__13_ ( .D(n1722), .CK(clk), .RN(rstn), .Q(memory[813]) );
  DFFRHQX1 memory_reg_13__12_ ( .D(n1723), .CK(clk), .RN(rstn), .Q(memory[812]) );
  DFFRHQX1 memory_reg_13__11_ ( .D(n1724), .CK(clk), .RN(rstn), .Q(memory[811]) );
  DFFRHQX1 memory_reg_13__10_ ( .D(n1725), .CK(clk), .RN(rstn), .Q(memory[810]) );
  DFFRHQX1 memory_reg_13__9_ ( .D(n1726), .CK(clk), .RN(rstn), .Q(memory[809])
         );
  DFFRHQX1 memory_reg_13__8_ ( .D(n1727), .CK(clk), .RN(rstn), .Q(memory[808])
         );
  DFFRHQX1 memory_reg_13__7_ ( .D(n1728), .CK(clk), .RN(rstn), .Q(memory[807])
         );
  DFFRHQX1 memory_reg_13__6_ ( .D(n1729), .CK(clk), .RN(rstn), .Q(memory[806])
         );
  DFFRHQX1 memory_reg_13__5_ ( .D(n1730), .CK(clk), .RN(rstn), .Q(memory[805])
         );
  DFFRHQX1 memory_reg_13__4_ ( .D(n1731), .CK(clk), .RN(rstn), .Q(memory[804])
         );
  DFFRHQX1 memory_reg_13__3_ ( .D(n1732), .CK(clk), .RN(rstn), .Q(memory[803])
         );
  DFFRHQX1 memory_reg_13__2_ ( .D(n1733), .CK(clk), .RN(rstn), .Q(memory[802])
         );
  DFFRHQX1 memory_reg_13__1_ ( .D(n1734), .CK(clk), .RN(rstn), .Q(memory[801])
         );
  DFFRHQX1 memory_reg_13__0_ ( .D(n1735), .CK(clk), .RN(rstn), .Q(memory[800])
         );
  DFFRHQX1 memory_reg_17__15_ ( .D(n1784), .CK(clk), .RN(rstn), .Q(memory[751]) );
  DFFRHQX1 memory_reg_17__14_ ( .D(n1785), .CK(clk), .RN(rstn), .Q(memory[750]) );
  DFFRHQX1 memory_reg_17__13_ ( .D(n1786), .CK(clk), .RN(rstn), .Q(memory[749]) );
  DFFRHQX1 memory_reg_17__12_ ( .D(n1787), .CK(clk), .RN(rstn), .Q(memory[748]) );
  DFFRHQX1 memory_reg_17__11_ ( .D(n1788), .CK(clk), .RN(rstn), .Q(memory[747]) );
  DFFRHQX1 memory_reg_17__10_ ( .D(n1789), .CK(clk), .RN(rstn), .Q(memory[746]) );
  DFFRHQX1 memory_reg_17__9_ ( .D(n1790), .CK(clk), .RN(rstn), .Q(memory[745])
         );
  DFFRHQX1 memory_reg_17__8_ ( .D(n1791), .CK(clk), .RN(rstn), .Q(memory[744])
         );
  DFFRHQX1 memory_reg_17__7_ ( .D(n1792), .CK(clk), .RN(rstn), .Q(memory[743])
         );
  DFFRHQX1 memory_reg_17__6_ ( .D(n1793), .CK(clk), .RN(rstn), .Q(memory[742])
         );
  DFFRHQX1 memory_reg_17__5_ ( .D(n1794), .CK(clk), .RN(rstn), .Q(memory[741])
         );
  DFFRHQX1 memory_reg_17__4_ ( .D(n1795), .CK(clk), .RN(rstn), .Q(memory[740])
         );
  DFFRHQX1 memory_reg_17__3_ ( .D(n1796), .CK(clk), .RN(rstn), .Q(memory[739])
         );
  DFFRHQX1 memory_reg_17__2_ ( .D(n1797), .CK(clk), .RN(rstn), .Q(memory[738])
         );
  DFFRHQX1 memory_reg_17__1_ ( .D(n1798), .CK(clk), .RN(rstn), .Q(memory[737])
         );
  DFFRHQX1 memory_reg_17__0_ ( .D(n1799), .CK(clk), .RN(rstn), .Q(memory[736])
         );
  DFFRHQX1 memory_reg_21__15_ ( .D(n1848), .CK(clk), .RN(rstn), .Q(memory[687]) );
  DFFRHQX1 memory_reg_21__14_ ( .D(n1849), .CK(clk), .RN(rstn), .Q(memory[686]) );
  DFFRHQX1 memory_reg_21__13_ ( .D(n1850), .CK(clk), .RN(rstn), .Q(memory[685]) );
  DFFRHQX1 memory_reg_21__12_ ( .D(n1851), .CK(clk), .RN(rstn), .Q(memory[684]) );
  DFFRHQX1 memory_reg_21__11_ ( .D(n1852), .CK(clk), .RN(rstn), .Q(memory[683]) );
  DFFRHQX1 memory_reg_21__10_ ( .D(n1853), .CK(clk), .RN(rstn), .Q(memory[682]) );
  DFFRHQX1 memory_reg_21__9_ ( .D(n1854), .CK(clk), .RN(rstn), .Q(memory[681])
         );
  DFFRHQX1 memory_reg_21__8_ ( .D(n1855), .CK(clk), .RN(rstn), .Q(memory[680])
         );
  DFFRHQX1 memory_reg_21__7_ ( .D(n1856), .CK(clk), .RN(rstn), .Q(memory[679])
         );
  DFFRHQX1 memory_reg_21__6_ ( .D(n1857), .CK(clk), .RN(rstn), .Q(memory[678])
         );
  DFFRHQX1 memory_reg_21__5_ ( .D(n1858), .CK(clk), .RN(rstn), .Q(memory[677])
         );
  DFFRHQX1 memory_reg_21__4_ ( .D(n1859), .CK(clk), .RN(rstn), .Q(memory[676])
         );
  DFFRHQX1 memory_reg_21__3_ ( .D(n1860), .CK(clk), .RN(rstn), .Q(memory[675])
         );
  DFFRHQX1 memory_reg_21__2_ ( .D(n1861), .CK(clk), .RN(rstn), .Q(memory[674])
         );
  DFFRHQX1 memory_reg_21__1_ ( .D(n1862), .CK(clk), .RN(rstn), .Q(memory[673])
         );
  DFFRHQX1 memory_reg_21__0_ ( .D(n1863), .CK(clk), .RN(rstn), .Q(memory[672])
         );
  DFFRHQX1 memory_reg_25__15_ ( .D(n1912), .CK(clk), .RN(rstn), .Q(memory[623]) );
  DFFRHQX1 memory_reg_25__14_ ( .D(n1913), .CK(clk), .RN(rstn), .Q(memory[622]) );
  DFFRHQX1 memory_reg_25__13_ ( .D(n1914), .CK(clk), .RN(rstn), .Q(memory[621]) );
  DFFRHQX1 memory_reg_25__12_ ( .D(n1915), .CK(clk), .RN(rstn), .Q(memory[620]) );
  DFFRHQX1 memory_reg_25__11_ ( .D(n1916), .CK(clk), .RN(rstn), .Q(memory[619]) );
  DFFRHQX1 memory_reg_25__10_ ( .D(n1917), .CK(clk), .RN(rstn), .Q(memory[618]) );
  DFFRHQX1 memory_reg_25__9_ ( .D(n1918), .CK(clk), .RN(rstn), .Q(memory[617])
         );
  DFFRHQX1 memory_reg_25__8_ ( .D(n1919), .CK(clk), .RN(rstn), .Q(memory[616])
         );
  DFFRHQX1 memory_reg_25__7_ ( .D(n1920), .CK(clk), .RN(rstn), .Q(memory[615])
         );
  DFFRHQX1 memory_reg_25__6_ ( .D(n1921), .CK(clk), .RN(rstn), .Q(memory[614])
         );
  DFFRHQX1 memory_reg_25__5_ ( .D(n1922), .CK(clk), .RN(rstn), .Q(memory[613])
         );
  DFFRHQX1 memory_reg_25__4_ ( .D(n1923), .CK(clk), .RN(rstn), .Q(memory[612])
         );
  DFFRHQX1 memory_reg_25__3_ ( .D(n1924), .CK(clk), .RN(rstn), .Q(memory[611])
         );
  DFFRHQX1 memory_reg_25__2_ ( .D(n1925), .CK(clk), .RN(rstn), .Q(memory[610])
         );
  DFFRHQX1 memory_reg_25__1_ ( .D(n1926), .CK(clk), .RN(rstn), .Q(memory[609])
         );
  DFFRHQX1 memory_reg_25__0_ ( .D(n1927), .CK(clk), .RN(rstn), .Q(memory[608])
         );
  DFFRHQX1 memory_reg_29__15_ ( .D(n1976), .CK(clk), .RN(rstn), .Q(memory[559]) );
  DFFRHQX1 memory_reg_29__14_ ( .D(n1977), .CK(clk), .RN(rstn), .Q(memory[558]) );
  DFFRHQX1 memory_reg_29__13_ ( .D(n1978), .CK(clk), .RN(rstn), .Q(memory[557]) );
  DFFRHQX1 memory_reg_29__12_ ( .D(n1979), .CK(clk), .RN(rstn), .Q(memory[556]) );
  DFFRHQX1 memory_reg_29__11_ ( .D(n1980), .CK(clk), .RN(rstn), .Q(memory[555]) );
  DFFRHQX1 memory_reg_29__10_ ( .D(n1981), .CK(clk), .RN(rstn), .Q(memory[554]) );
  DFFRHQX1 memory_reg_29__9_ ( .D(n1982), .CK(clk), .RN(rstn), .Q(memory[553])
         );
  DFFRHQX1 memory_reg_29__8_ ( .D(n1983), .CK(clk), .RN(rstn), .Q(memory[552])
         );
  DFFRHQX1 memory_reg_29__7_ ( .D(n1984), .CK(clk), .RN(rstn), .Q(memory[551])
         );
  DFFRHQX1 memory_reg_29__6_ ( .D(n1985), .CK(clk), .RN(rstn), .Q(memory[550])
         );
  DFFRHQX1 memory_reg_29__5_ ( .D(n1986), .CK(clk), .RN(rstn), .Q(memory[549])
         );
  DFFRHQX1 memory_reg_29__4_ ( .D(n1987), .CK(clk), .RN(rstn), .Q(memory[548])
         );
  DFFRHQX1 memory_reg_29__3_ ( .D(n1988), .CK(clk), .RN(rstn), .Q(memory[547])
         );
  DFFRHQX1 memory_reg_29__2_ ( .D(n1989), .CK(clk), .RN(rstn), .Q(memory[546])
         );
  DFFRHQX1 memory_reg_29__1_ ( .D(n1990), .CK(clk), .RN(rstn), .Q(memory[545])
         );
  DFFRHQX1 memory_reg_29__0_ ( .D(n1991), .CK(clk), .RN(rstn), .Q(memory[544])
         );
  DFFRHQX1 memory_reg_33__15_ ( .D(n2040), .CK(clk), .RN(rstn), .Q(memory[495]) );
  DFFRHQX1 memory_reg_33__14_ ( .D(n2041), .CK(clk), .RN(rstn), .Q(memory[494]) );
  DFFRHQX1 memory_reg_33__13_ ( .D(n2042), .CK(clk), .RN(rstn), .Q(memory[493]) );
  DFFRHQX1 memory_reg_33__12_ ( .D(n2043), .CK(clk), .RN(rstn), .Q(memory[492]) );
  DFFRHQX1 memory_reg_33__11_ ( .D(n2044), .CK(clk), .RN(rstn), .Q(memory[491]) );
  DFFRHQX1 memory_reg_33__10_ ( .D(n2045), .CK(clk), .RN(rstn), .Q(memory[490]) );
  DFFRHQX1 memory_reg_33__9_ ( .D(n2046), .CK(clk), .RN(rstn), .Q(memory[489])
         );
  DFFRHQX1 memory_reg_33__8_ ( .D(n2047), .CK(clk), .RN(rstn), .Q(memory[488])
         );
  DFFRHQX1 memory_reg_33__7_ ( .D(n2048), .CK(clk), .RN(rstn), .Q(memory[487])
         );
  DFFRHQX1 memory_reg_33__6_ ( .D(n2049), .CK(clk), .RN(rstn), .Q(memory[486])
         );
  DFFRHQX1 memory_reg_33__5_ ( .D(n2050), .CK(clk), .RN(rstn), .Q(memory[485])
         );
  DFFRHQX1 memory_reg_33__4_ ( .D(n2051), .CK(clk), .RN(rstn), .Q(memory[484])
         );
  DFFRHQX1 memory_reg_33__3_ ( .D(n2052), .CK(clk), .RN(rstn), .Q(memory[483])
         );
  DFFRHQX1 memory_reg_33__2_ ( .D(n2053), .CK(clk), .RN(rstn), .Q(memory[482])
         );
  DFFRHQX1 memory_reg_33__1_ ( .D(n2054), .CK(clk), .RN(rstn), .Q(memory[481])
         );
  DFFRHQX1 memory_reg_33__0_ ( .D(n2055), .CK(clk), .RN(rstn), .Q(memory[480])
         );
  DFFRHQX1 memory_reg_37__15_ ( .D(n2104), .CK(clk), .RN(rstn), .Q(memory[431]) );
  DFFRHQX1 memory_reg_37__14_ ( .D(n2105), .CK(clk), .RN(rstn), .Q(memory[430]) );
  DFFRHQX1 memory_reg_37__13_ ( .D(n2106), .CK(clk), .RN(rstn), .Q(memory[429]) );
  DFFRHQX1 memory_reg_37__12_ ( .D(n2107), .CK(clk), .RN(rstn), .Q(memory[428]) );
  DFFRHQX1 memory_reg_37__11_ ( .D(n2108), .CK(clk), .RN(rstn), .Q(memory[427]) );
  DFFRHQX1 memory_reg_37__10_ ( .D(n2109), .CK(clk), .RN(rstn), .Q(memory[426]) );
  DFFRHQX1 memory_reg_37__9_ ( .D(n2110), .CK(clk), .RN(rstn), .Q(memory[425])
         );
  DFFRHQX1 memory_reg_37__8_ ( .D(n2111), .CK(clk), .RN(rstn), .Q(memory[424])
         );
  DFFRHQX1 memory_reg_37__7_ ( .D(n2112), .CK(clk), .RN(rstn), .Q(memory[423])
         );
  DFFRHQX1 memory_reg_37__6_ ( .D(n2113), .CK(clk), .RN(rstn), .Q(memory[422])
         );
  DFFRHQX1 memory_reg_37__5_ ( .D(n2114), .CK(clk), .RN(rstn), .Q(memory[421])
         );
  DFFRHQX1 memory_reg_37__4_ ( .D(n2115), .CK(clk), .RN(rstn), .Q(memory[420])
         );
  DFFRHQX1 memory_reg_37__3_ ( .D(n2116), .CK(clk), .RN(rstn), .Q(memory[419])
         );
  DFFRHQX1 memory_reg_37__2_ ( .D(n2117), .CK(clk), .RN(rstn), .Q(memory[418])
         );
  DFFRHQX1 memory_reg_37__1_ ( .D(n2118), .CK(clk), .RN(rstn), .Q(memory[417])
         );
  DFFRHQX1 memory_reg_37__0_ ( .D(n2119), .CK(clk), .RN(rstn), .Q(memory[416])
         );
  DFFRHQX1 memory_reg_41__15_ ( .D(n2168), .CK(clk), .RN(rstn), .Q(memory[367]) );
  DFFRHQX1 memory_reg_41__14_ ( .D(n2169), .CK(clk), .RN(rstn), .Q(memory[366]) );
  DFFRHQX1 memory_reg_41__13_ ( .D(n2170), .CK(clk), .RN(rstn), .Q(memory[365]) );
  DFFRHQX1 memory_reg_41__12_ ( .D(n2171), .CK(clk), .RN(rstn), .Q(memory[364]) );
  DFFRHQX1 memory_reg_41__11_ ( .D(n2172), .CK(clk), .RN(rstn), .Q(memory[363]) );
  DFFRHQX1 memory_reg_41__10_ ( .D(n2173), .CK(clk), .RN(rstn), .Q(memory[362]) );
  DFFRHQX1 memory_reg_41__9_ ( .D(n2174), .CK(clk), .RN(rstn), .Q(memory[361])
         );
  DFFRHQX1 memory_reg_41__8_ ( .D(n2175), .CK(clk), .RN(rstn), .Q(memory[360])
         );
  DFFRHQX1 memory_reg_41__7_ ( .D(n2176), .CK(clk), .RN(rstn), .Q(memory[359])
         );
  DFFRHQX1 memory_reg_41__6_ ( .D(n2177), .CK(clk), .RN(rstn), .Q(memory[358])
         );
  DFFRHQX1 memory_reg_41__5_ ( .D(n2178), .CK(clk), .RN(rstn), .Q(memory[357])
         );
  DFFRHQX1 memory_reg_41__4_ ( .D(n2179), .CK(clk), .RN(rstn), .Q(memory[356])
         );
  DFFRHQX1 memory_reg_41__3_ ( .D(n2180), .CK(clk), .RN(rstn), .Q(memory[355])
         );
  DFFRHQX1 memory_reg_41__2_ ( .D(n2181), .CK(clk), .RN(rstn), .Q(memory[354])
         );
  DFFRHQX1 memory_reg_41__1_ ( .D(n2182), .CK(clk), .RN(rstn), .Q(memory[353])
         );
  DFFRHQX1 memory_reg_41__0_ ( .D(n2183), .CK(clk), .RN(rstn), .Q(memory[352])
         );
  DFFRHQX1 memory_reg_45__15_ ( .D(n2232), .CK(clk), .RN(rstn), .Q(memory[303]) );
  DFFRHQX1 memory_reg_45__14_ ( .D(n2233), .CK(clk), .RN(rstn), .Q(memory[302]) );
  DFFRHQX1 memory_reg_45__13_ ( .D(n2234), .CK(clk), .RN(rstn), .Q(memory[301]) );
  DFFRHQX1 memory_reg_45__12_ ( .D(n2235), .CK(clk), .RN(rstn), .Q(memory[300]) );
  DFFRHQX1 memory_reg_45__11_ ( .D(n2236), .CK(clk), .RN(rstn), .Q(memory[299]) );
  DFFRHQX1 memory_reg_45__10_ ( .D(n2237), .CK(clk), .RN(rstn), .Q(memory[298]) );
  DFFRHQX1 memory_reg_45__9_ ( .D(n2238), .CK(clk), .RN(rstn), .Q(memory[297])
         );
  DFFRHQX1 memory_reg_45__8_ ( .D(n2239), .CK(clk), .RN(rstn), .Q(memory[296])
         );
  DFFRHQX1 memory_reg_45__7_ ( .D(n2240), .CK(clk), .RN(rstn), .Q(memory[295])
         );
  DFFRHQX1 memory_reg_45__6_ ( .D(n2241), .CK(clk), .RN(rstn), .Q(memory[294])
         );
  DFFRHQX1 memory_reg_45__5_ ( .D(n2242), .CK(clk), .RN(rstn), .Q(memory[293])
         );
  DFFRHQX1 memory_reg_45__4_ ( .D(n2243), .CK(clk), .RN(rstn), .Q(memory[292])
         );
  DFFRHQX1 memory_reg_45__3_ ( .D(n2244), .CK(clk), .RN(rstn), .Q(memory[291])
         );
  DFFRHQX1 memory_reg_45__2_ ( .D(n2245), .CK(clk), .RN(rstn), .Q(memory[290])
         );
  DFFRHQX1 memory_reg_45__1_ ( .D(n2246), .CK(clk), .RN(rstn), .Q(memory[289])
         );
  DFFRHQX1 memory_reg_45__0_ ( .D(n2247), .CK(clk), .RN(rstn), .Q(memory[288])
         );
  DFFRHQX1 memory_reg_49__15_ ( .D(n2296), .CK(clk), .RN(rstn), .Q(memory[239]) );
  DFFRHQX1 memory_reg_49__14_ ( .D(n2297), .CK(clk), .RN(rstn), .Q(memory[238]) );
  DFFRHQX1 memory_reg_49__13_ ( .D(n2298), .CK(clk), .RN(rstn), .Q(memory[237]) );
  DFFRHQX1 memory_reg_49__12_ ( .D(n2299), .CK(clk), .RN(rstn), .Q(memory[236]) );
  DFFRHQX1 memory_reg_49__11_ ( .D(n2300), .CK(clk), .RN(rstn), .Q(memory[235]) );
  DFFRHQX1 memory_reg_49__10_ ( .D(n2301), .CK(clk), .RN(rstn), .Q(memory[234]) );
  DFFRHQX1 memory_reg_49__9_ ( .D(n2302), .CK(clk), .RN(rstn), .Q(memory[233])
         );
  DFFRHQX1 memory_reg_49__8_ ( .D(n2303), .CK(clk), .RN(rstn), .Q(memory[232])
         );
  DFFRHQX1 memory_reg_49__7_ ( .D(n2304), .CK(clk), .RN(rstn), .Q(memory[231])
         );
  DFFRHQX1 memory_reg_49__6_ ( .D(n2305), .CK(clk), .RN(rstn), .Q(memory[230])
         );
  DFFRHQX1 memory_reg_49__5_ ( .D(n2306), .CK(clk), .RN(rstn), .Q(memory[229])
         );
  DFFRHQX1 memory_reg_49__4_ ( .D(n2307), .CK(clk), .RN(rstn), .Q(memory[228])
         );
  DFFRHQX1 memory_reg_49__3_ ( .D(n2308), .CK(clk), .RN(rstn), .Q(memory[227])
         );
  DFFRHQX1 memory_reg_49__2_ ( .D(n2309), .CK(clk), .RN(rstn), .Q(memory[226])
         );
  DFFRHQX1 memory_reg_49__1_ ( .D(n2310), .CK(clk), .RN(rstn), .Q(memory[225])
         );
  DFFRHQX1 memory_reg_49__0_ ( .D(n2311), .CK(clk), .RN(rstn), .Q(memory[224])
         );
  DFFRHQX1 memory_reg_53__15_ ( .D(n2360), .CK(clk), .RN(rstn), .Q(memory[175]) );
  DFFRHQX1 memory_reg_53__14_ ( .D(n2361), .CK(clk), .RN(rstn), .Q(memory[174]) );
  DFFRHQX1 memory_reg_53__13_ ( .D(n2362), .CK(clk), .RN(rstn), .Q(memory[173]) );
  DFFRHQX1 memory_reg_53__12_ ( .D(n2363), .CK(clk), .RN(rstn), .Q(memory[172]) );
  DFFRHQX1 memory_reg_53__11_ ( .D(n2364), .CK(clk), .RN(rstn), .Q(memory[171]) );
  DFFRHQX1 memory_reg_53__10_ ( .D(n2365), .CK(clk), .RN(rstn), .Q(memory[170]) );
  DFFRHQX1 memory_reg_53__9_ ( .D(n2366), .CK(clk), .RN(rstn), .Q(memory[169])
         );
  DFFRHQX1 memory_reg_53__8_ ( .D(n2367), .CK(clk), .RN(rstn), .Q(memory[168])
         );
  DFFRHQX1 memory_reg_53__7_ ( .D(n2368), .CK(clk), .RN(rstn), .Q(memory[167])
         );
  DFFRHQX1 memory_reg_53__6_ ( .D(n2369), .CK(clk), .RN(rstn), .Q(memory[166])
         );
  DFFRHQX1 memory_reg_53__5_ ( .D(n2370), .CK(clk), .RN(rstn), .Q(memory[165])
         );
  DFFRHQX1 memory_reg_53__4_ ( .D(n2371), .CK(clk), .RN(rstn), .Q(memory[164])
         );
  DFFRHQX1 memory_reg_53__3_ ( .D(n2372), .CK(clk), .RN(rstn), .Q(memory[163])
         );
  DFFRHQX1 memory_reg_53__2_ ( .D(n2373), .CK(clk), .RN(rstn), .Q(memory[162])
         );
  DFFRHQX1 memory_reg_53__1_ ( .D(n2374), .CK(clk), .RN(rstn), .Q(memory[161])
         );
  DFFRHQX1 memory_reg_53__0_ ( .D(n2375), .CK(clk), .RN(rstn), .Q(memory[160])
         );
  DFFRHQX1 memory_reg_57__15_ ( .D(n2424), .CK(clk), .RN(rstn), .Q(memory[111]) );
  DFFRHQX1 memory_reg_57__14_ ( .D(n2425), .CK(clk), .RN(rstn), .Q(memory[110]) );
  DFFRHQX1 memory_reg_57__13_ ( .D(n2426), .CK(clk), .RN(rstn), .Q(memory[109]) );
  DFFRHQX1 memory_reg_57__12_ ( .D(n2427), .CK(clk), .RN(rstn), .Q(memory[108]) );
  DFFRHQX1 memory_reg_57__11_ ( .D(n2428), .CK(clk), .RN(rstn), .Q(memory[107]) );
  DFFRHQX1 memory_reg_57__10_ ( .D(n2429), .CK(clk), .RN(rstn), .Q(memory[106]) );
  DFFRHQX1 memory_reg_57__9_ ( .D(n2430), .CK(clk), .RN(rstn), .Q(memory[105])
         );
  DFFRHQX1 memory_reg_57__8_ ( .D(n2431), .CK(clk), .RN(rstn), .Q(memory[104])
         );
  DFFRHQX1 memory_reg_57__7_ ( .D(n2432), .CK(clk), .RN(rstn), .Q(memory[103])
         );
  DFFRHQX1 memory_reg_57__6_ ( .D(n2433), .CK(clk), .RN(rstn), .Q(memory[102])
         );
  DFFRHQX1 memory_reg_57__5_ ( .D(n2434), .CK(clk), .RN(rstn), .Q(memory[101])
         );
  DFFRHQX1 memory_reg_57__4_ ( .D(n2435), .CK(clk), .RN(rstn), .Q(memory[100])
         );
  DFFRHQX1 memory_reg_57__3_ ( .D(n2436), .CK(clk), .RN(rstn), .Q(memory[99])
         );
  DFFRHQX1 memory_reg_57__2_ ( .D(n2437), .CK(clk), .RN(rstn), .Q(memory[98])
         );
  DFFRHQX1 memory_reg_57__1_ ( .D(n2438), .CK(clk), .RN(rstn), .Q(memory[97])
         );
  DFFRHQX1 memory_reg_57__0_ ( .D(n2439), .CK(clk), .RN(rstn), .Q(memory[96])
         );
  DFFRHQX1 memory_reg_61__15_ ( .D(n2488), .CK(clk), .RN(rstn), .Q(memory[47])
         );
  DFFRHQX1 memory_reg_61__14_ ( .D(n2489), .CK(clk), .RN(rstn), .Q(memory[46])
         );
  DFFRHQX1 memory_reg_61__13_ ( .D(n2490), .CK(clk), .RN(rstn), .Q(memory[45])
         );
  DFFRHQX1 memory_reg_61__12_ ( .D(n2491), .CK(clk), .RN(rstn), .Q(memory[44])
         );
  DFFRHQX1 memory_reg_61__11_ ( .D(n2492), .CK(clk), .RN(rstn), .Q(memory[43])
         );
  DFFRHQX1 memory_reg_61__10_ ( .D(n2493), .CK(clk), .RN(rstn), .Q(memory[42])
         );
  DFFRHQX1 memory_reg_61__9_ ( .D(n2494), .CK(clk), .RN(rstn), .Q(memory[41])
         );
  DFFRHQX1 memory_reg_61__8_ ( .D(n2495), .CK(clk), .RN(rstn), .Q(memory[40])
         );
  DFFRHQX1 memory_reg_61__7_ ( .D(n2496), .CK(clk), .RN(rstn), .Q(memory[39])
         );
  DFFRHQX1 memory_reg_61__6_ ( .D(n2497), .CK(clk), .RN(rstn), .Q(memory[38])
         );
  DFFRHQX1 memory_reg_61__5_ ( .D(n2498), .CK(clk), .RN(rstn), .Q(memory[37])
         );
  DFFRHQX1 memory_reg_61__4_ ( .D(n2499), .CK(clk), .RN(rstn), .Q(memory[36])
         );
  DFFRHQX1 memory_reg_61__3_ ( .D(n2500), .CK(clk), .RN(rstn), .Q(memory[35])
         );
  DFFRHQX1 memory_reg_61__2_ ( .D(n2501), .CK(clk), .RN(rstn), .Q(memory[34])
         );
  DFFRHQX1 memory_reg_61__1_ ( .D(n2502), .CK(clk), .RN(rstn), .Q(memory[33])
         );
  DFFRHQX1 memory_reg_61__0_ ( .D(n2503), .CK(clk), .RN(rstn), .Q(memory[32])
         );
  DFFRHQX1 memory_reg_3__15_ ( .D(n1560), .CK(clk), .RN(rstn), .Q(memory[975])
         );
  DFFRHQX1 memory_reg_3__14_ ( .D(n1561), .CK(clk), .RN(rstn), .Q(memory[974])
         );
  DFFRHQX1 memory_reg_3__13_ ( .D(n1562), .CK(clk), .RN(rstn), .Q(memory[973])
         );
  DFFRHQX1 memory_reg_3__12_ ( .D(n1563), .CK(clk), .RN(rstn), .Q(memory[972])
         );
  DFFRHQX1 memory_reg_3__11_ ( .D(n1564), .CK(clk), .RN(rstn), .Q(memory[971])
         );
  DFFRHQX1 memory_reg_3__10_ ( .D(n1565), .CK(clk), .RN(rstn), .Q(memory[970])
         );
  DFFRHQX1 memory_reg_3__9_ ( .D(n1566), .CK(clk), .RN(rstn), .Q(memory[969])
         );
  DFFRHQX1 memory_reg_3__8_ ( .D(n1567), .CK(clk), .RN(rstn), .Q(memory[968])
         );
  DFFRHQX1 memory_reg_3__7_ ( .D(n1568), .CK(clk), .RN(rstn), .Q(memory[967])
         );
  DFFRHQX1 memory_reg_3__6_ ( .D(n1569), .CK(clk), .RN(rstn), .Q(memory[966])
         );
  DFFRHQX1 memory_reg_3__5_ ( .D(n1570), .CK(clk), .RN(rstn), .Q(memory[965])
         );
  DFFRHQX1 memory_reg_3__4_ ( .D(n1571), .CK(clk), .RN(rstn), .Q(memory[964])
         );
  DFFRHQX1 memory_reg_3__3_ ( .D(n1572), .CK(clk), .RN(rstn), .Q(memory[963])
         );
  DFFRHQX1 memory_reg_3__2_ ( .D(n1573), .CK(clk), .RN(rstn), .Q(memory[962])
         );
  DFFRHQX1 memory_reg_3__1_ ( .D(n1574), .CK(clk), .RN(rstn), .Q(memory[961])
         );
  DFFRHQX1 memory_reg_3__0_ ( .D(n1575), .CK(clk), .RN(rstn), .Q(memory[960])
         );
  DFFRHQX1 memory_reg_7__15_ ( .D(n1624), .CK(clk), .RN(rstn), .Q(memory[911])
         );
  DFFRHQX1 memory_reg_7__14_ ( .D(n1625), .CK(clk), .RN(rstn), .Q(memory[910])
         );
  DFFRHQX1 memory_reg_7__13_ ( .D(n1626), .CK(clk), .RN(rstn), .Q(memory[909])
         );
  DFFRHQX1 memory_reg_7__12_ ( .D(n1627), .CK(clk), .RN(rstn), .Q(memory[908])
         );
  DFFRHQX1 memory_reg_7__11_ ( .D(n1628), .CK(clk), .RN(rstn), .Q(memory[907])
         );
  DFFRHQX1 memory_reg_7__10_ ( .D(n1629), .CK(clk), .RN(rstn), .Q(memory[906])
         );
  DFFRHQX1 memory_reg_7__9_ ( .D(n1630), .CK(clk), .RN(rstn), .Q(memory[905])
         );
  DFFRHQX1 memory_reg_7__8_ ( .D(n1631), .CK(clk), .RN(rstn), .Q(memory[904])
         );
  DFFRHQX1 memory_reg_7__7_ ( .D(n1632), .CK(clk), .RN(rstn), .Q(memory[903])
         );
  DFFRHQX1 memory_reg_7__6_ ( .D(n1633), .CK(clk), .RN(rstn), .Q(memory[902])
         );
  DFFRHQX1 memory_reg_7__5_ ( .D(n1634), .CK(clk), .RN(rstn), .Q(memory[901])
         );
  DFFRHQX1 memory_reg_7__4_ ( .D(n1635), .CK(clk), .RN(rstn), .Q(memory[900])
         );
  DFFRHQX1 memory_reg_7__3_ ( .D(n1636), .CK(clk), .RN(rstn), .Q(memory[899])
         );
  DFFRHQX1 memory_reg_7__2_ ( .D(n1637), .CK(clk), .RN(rstn), .Q(memory[898])
         );
  DFFRHQX1 memory_reg_7__1_ ( .D(n1638), .CK(clk), .RN(rstn), .Q(memory[897])
         );
  DFFRHQX1 memory_reg_7__0_ ( .D(n1639), .CK(clk), .RN(rstn), .Q(memory[896])
         );
  DFFRHQX1 memory_reg_11__15_ ( .D(n1688), .CK(clk), .RN(rstn), .Q(memory[847]) );
  DFFRHQX1 memory_reg_11__14_ ( .D(n1689), .CK(clk), .RN(rstn), .Q(memory[846]) );
  DFFRHQX1 memory_reg_11__13_ ( .D(n1690), .CK(clk), .RN(rstn), .Q(memory[845]) );
  DFFRHQX1 memory_reg_11__12_ ( .D(n1691), .CK(clk), .RN(rstn), .Q(memory[844]) );
  DFFRHQX1 memory_reg_11__11_ ( .D(n1692), .CK(clk), .RN(rstn), .Q(memory[843]) );
  DFFRHQX1 memory_reg_11__10_ ( .D(n1693), .CK(clk), .RN(rstn), .Q(memory[842]) );
  DFFRHQX1 memory_reg_11__9_ ( .D(n1694), .CK(clk), .RN(rstn), .Q(memory[841])
         );
  DFFRHQX1 memory_reg_11__8_ ( .D(n1695), .CK(clk), .RN(rstn), .Q(memory[840])
         );
  DFFRHQX1 memory_reg_11__7_ ( .D(n1696), .CK(clk), .RN(rstn), .Q(memory[839])
         );
  DFFRHQX1 memory_reg_11__6_ ( .D(n1697), .CK(clk), .RN(rstn), .Q(memory[838])
         );
  DFFRHQX1 memory_reg_11__5_ ( .D(n1698), .CK(clk), .RN(rstn), .Q(memory[837])
         );
  DFFRHQX1 memory_reg_11__4_ ( .D(n1699), .CK(clk), .RN(rstn), .Q(memory[836])
         );
  DFFRHQX1 memory_reg_11__3_ ( .D(n1700), .CK(clk), .RN(rstn), .Q(memory[835])
         );
  DFFRHQX1 memory_reg_11__2_ ( .D(n1701), .CK(clk), .RN(rstn), .Q(memory[834])
         );
  DFFRHQX1 memory_reg_11__1_ ( .D(n1702), .CK(clk), .RN(rstn), .Q(memory[833])
         );
  DFFRHQX1 memory_reg_11__0_ ( .D(n1703), .CK(clk), .RN(rstn), .Q(memory[832])
         );
  DFFRHQX1 memory_reg_15__15_ ( .D(n1752), .CK(clk), .RN(rstn), .Q(memory[783]) );
  DFFRHQX1 memory_reg_15__14_ ( .D(n1753), .CK(clk), .RN(rstn), .Q(memory[782]) );
  DFFRHQX1 memory_reg_15__13_ ( .D(n1754), .CK(clk), .RN(rstn), .Q(memory[781]) );
  DFFRHQX1 memory_reg_15__12_ ( .D(n1755), .CK(clk), .RN(rstn), .Q(memory[780]) );
  DFFRHQX1 memory_reg_15__11_ ( .D(n1756), .CK(clk), .RN(rstn), .Q(memory[779]) );
  DFFRHQX1 memory_reg_15__10_ ( .D(n1757), .CK(clk), .RN(rstn), .Q(memory[778]) );
  DFFRHQX1 memory_reg_15__9_ ( .D(n1758), .CK(clk), .RN(rstn), .Q(memory[777])
         );
  DFFRHQX1 memory_reg_15__8_ ( .D(n1759), .CK(clk), .RN(rstn), .Q(memory[776])
         );
  DFFRHQX1 memory_reg_15__7_ ( .D(n1760), .CK(clk), .RN(rstn), .Q(memory[775])
         );
  DFFRHQX1 memory_reg_15__6_ ( .D(n1761), .CK(clk), .RN(rstn), .Q(memory[774])
         );
  DFFRHQX1 memory_reg_15__5_ ( .D(n1762), .CK(clk), .RN(rstn), .Q(memory[773])
         );
  DFFRHQX1 memory_reg_15__4_ ( .D(n1763), .CK(clk), .RN(rstn), .Q(memory[772])
         );
  DFFRHQX1 memory_reg_15__3_ ( .D(n1764), .CK(clk), .RN(rstn), .Q(memory[771])
         );
  DFFRHQX1 memory_reg_15__2_ ( .D(n1765), .CK(clk), .RN(rstn), .Q(memory[770])
         );
  DFFRHQX1 memory_reg_15__1_ ( .D(n1766), .CK(clk), .RN(rstn), .Q(memory[769])
         );
  DFFRHQX1 memory_reg_15__0_ ( .D(n1767), .CK(clk), .RN(rstn), .Q(memory[768])
         );
  DFFRHQX1 memory_reg_19__15_ ( .D(n1816), .CK(clk), .RN(rstn), .Q(memory[719]) );
  DFFRHQX1 memory_reg_19__14_ ( .D(n1817), .CK(clk), .RN(rstn), .Q(memory[718]) );
  DFFRHQX1 memory_reg_19__13_ ( .D(n1818), .CK(clk), .RN(rstn), .Q(memory[717]) );
  DFFRHQX1 memory_reg_19__12_ ( .D(n1819), .CK(clk), .RN(rstn), .Q(memory[716]) );
  DFFRHQX1 memory_reg_19__11_ ( .D(n1820), .CK(clk), .RN(rstn), .Q(memory[715]) );
  DFFRHQX1 memory_reg_19__10_ ( .D(n1821), .CK(clk), .RN(rstn), .Q(memory[714]) );
  DFFRHQX1 memory_reg_19__9_ ( .D(n1822), .CK(clk), .RN(rstn), .Q(memory[713])
         );
  DFFRHQX1 memory_reg_19__8_ ( .D(n1823), .CK(clk), .RN(rstn), .Q(memory[712])
         );
  DFFRHQX1 memory_reg_19__7_ ( .D(n1824), .CK(clk), .RN(rstn), .Q(memory[711])
         );
  DFFRHQX1 memory_reg_19__6_ ( .D(n1825), .CK(clk), .RN(rstn), .Q(memory[710])
         );
  DFFRHQX1 memory_reg_19__5_ ( .D(n1826), .CK(clk), .RN(rstn), .Q(memory[709])
         );
  DFFRHQX1 memory_reg_19__4_ ( .D(n1827), .CK(clk), .RN(rstn), .Q(memory[708])
         );
  DFFRHQX1 memory_reg_19__3_ ( .D(n1828), .CK(clk), .RN(rstn), .Q(memory[707])
         );
  DFFRHQX1 memory_reg_19__2_ ( .D(n1829), .CK(clk), .RN(rstn), .Q(memory[706])
         );
  DFFRHQX1 memory_reg_19__1_ ( .D(n1830), .CK(clk), .RN(rstn), .Q(memory[705])
         );
  DFFRHQX1 memory_reg_19__0_ ( .D(n1831), .CK(clk), .RN(rstn), .Q(memory[704])
         );
  DFFRHQX1 memory_reg_23__15_ ( .D(n1880), .CK(clk), .RN(rstn), .Q(memory[655]) );
  DFFRHQX1 memory_reg_23__14_ ( .D(n1881), .CK(clk), .RN(rstn), .Q(memory[654]) );
  DFFRHQX1 memory_reg_23__13_ ( .D(n1882), .CK(clk), .RN(rstn), .Q(memory[653]) );
  DFFRHQX1 memory_reg_23__12_ ( .D(n1883), .CK(clk), .RN(rstn), .Q(memory[652]) );
  DFFRHQX1 memory_reg_23__11_ ( .D(n1884), .CK(clk), .RN(rstn), .Q(memory[651]) );
  DFFRHQX1 memory_reg_23__10_ ( .D(n1885), .CK(clk), .RN(rstn), .Q(memory[650]) );
  DFFRHQX1 memory_reg_23__9_ ( .D(n1886), .CK(clk), .RN(rstn), .Q(memory[649])
         );
  DFFRHQX1 memory_reg_23__8_ ( .D(n1887), .CK(clk), .RN(rstn), .Q(memory[648])
         );
  DFFRHQX1 memory_reg_23__7_ ( .D(n1888), .CK(clk), .RN(rstn), .Q(memory[647])
         );
  DFFRHQX1 memory_reg_23__6_ ( .D(n1889), .CK(clk), .RN(rstn), .Q(memory[646])
         );
  DFFRHQX1 memory_reg_23__5_ ( .D(n1890), .CK(clk), .RN(rstn), .Q(memory[645])
         );
  DFFRHQX1 memory_reg_23__4_ ( .D(n1891), .CK(clk), .RN(rstn), .Q(memory[644])
         );
  DFFRHQX1 memory_reg_23__3_ ( .D(n1892), .CK(clk), .RN(rstn), .Q(memory[643])
         );
  DFFRHQX1 memory_reg_23__2_ ( .D(n1893), .CK(clk), .RN(rstn), .Q(memory[642])
         );
  DFFRHQX1 memory_reg_23__1_ ( .D(n1894), .CK(clk), .RN(rstn), .Q(memory[641])
         );
  DFFRHQX1 memory_reg_23__0_ ( .D(n1895), .CK(clk), .RN(rstn), .Q(memory[640])
         );
  DFFRHQX1 memory_reg_27__15_ ( .D(n1944), .CK(clk), .RN(rstn), .Q(memory[591]) );
  DFFRHQX1 memory_reg_27__14_ ( .D(n1945), .CK(clk), .RN(rstn), .Q(memory[590]) );
  DFFRHQX1 memory_reg_27__13_ ( .D(n1946), .CK(clk), .RN(rstn), .Q(memory[589]) );
  DFFRHQX1 memory_reg_27__12_ ( .D(n1947), .CK(clk), .RN(rstn), .Q(memory[588]) );
  DFFRHQX1 memory_reg_27__11_ ( .D(n1948), .CK(clk), .RN(rstn), .Q(memory[587]) );
  DFFRHQX1 memory_reg_27__10_ ( .D(n1949), .CK(clk), .RN(rstn), .Q(memory[586]) );
  DFFRHQX1 memory_reg_27__9_ ( .D(n1950), .CK(clk), .RN(rstn), .Q(memory[585])
         );
  DFFRHQX1 memory_reg_27__8_ ( .D(n1951), .CK(clk), .RN(rstn), .Q(memory[584])
         );
  DFFRHQX1 memory_reg_27__7_ ( .D(n1952), .CK(clk), .RN(rstn), .Q(memory[583])
         );
  DFFRHQX1 memory_reg_27__6_ ( .D(n1953), .CK(clk), .RN(rstn), .Q(memory[582])
         );
  DFFRHQX1 memory_reg_27__5_ ( .D(n1954), .CK(clk), .RN(rstn), .Q(memory[581])
         );
  DFFRHQX1 memory_reg_27__4_ ( .D(n1955), .CK(clk), .RN(rstn), .Q(memory[580])
         );
  DFFRHQX1 memory_reg_27__3_ ( .D(n1956), .CK(clk), .RN(rstn), .Q(memory[579])
         );
  DFFRHQX1 memory_reg_27__2_ ( .D(n1957), .CK(clk), .RN(rstn), .Q(memory[578])
         );
  DFFRHQX1 memory_reg_27__1_ ( .D(n1958), .CK(clk), .RN(rstn), .Q(memory[577])
         );
  DFFRHQX1 memory_reg_27__0_ ( .D(n1959), .CK(clk), .RN(rstn), .Q(memory[576])
         );
  DFFRHQX1 memory_reg_31__15_ ( .D(n2008), .CK(clk), .RN(rstn), .Q(memory[527]) );
  DFFRHQX1 memory_reg_31__14_ ( .D(n2009), .CK(clk), .RN(rstn), .Q(memory[526]) );
  DFFRHQX1 memory_reg_31__13_ ( .D(n2010), .CK(clk), .RN(rstn), .Q(memory[525]) );
  DFFRHQX1 memory_reg_31__12_ ( .D(n2011), .CK(clk), .RN(rstn), .Q(memory[524]) );
  DFFRHQX1 memory_reg_31__11_ ( .D(n2012), .CK(clk), .RN(rstn), .Q(memory[523]) );
  DFFRHQX1 memory_reg_31__10_ ( .D(n2013), .CK(clk), .RN(rstn), .Q(memory[522]) );
  DFFRHQX1 memory_reg_31__9_ ( .D(n2014), .CK(clk), .RN(rstn), .Q(memory[521])
         );
  DFFRHQX1 memory_reg_31__8_ ( .D(n2015), .CK(clk), .RN(rstn), .Q(memory[520])
         );
  DFFRHQX1 memory_reg_31__7_ ( .D(n2016), .CK(clk), .RN(rstn), .Q(memory[519])
         );
  DFFRHQX1 memory_reg_31__6_ ( .D(n2017), .CK(clk), .RN(rstn), .Q(memory[518])
         );
  DFFRHQX1 memory_reg_31__5_ ( .D(n2018), .CK(clk), .RN(rstn), .Q(memory[517])
         );
  DFFRHQX1 memory_reg_31__4_ ( .D(n2019), .CK(clk), .RN(rstn), .Q(memory[516])
         );
  DFFRHQX1 memory_reg_31__3_ ( .D(n2020), .CK(clk), .RN(rstn), .Q(memory[515])
         );
  DFFRHQX1 memory_reg_31__2_ ( .D(n2021), .CK(clk), .RN(rstn), .Q(memory[514])
         );
  DFFRHQX1 memory_reg_31__1_ ( .D(n2022), .CK(clk), .RN(rstn), .Q(memory[513])
         );
  DFFRHQX1 memory_reg_31__0_ ( .D(n2023), .CK(clk), .RN(rstn), .Q(memory[512])
         );
  DFFRHQX1 memory_reg_35__15_ ( .D(n2072), .CK(clk), .RN(rstn), .Q(memory[463]) );
  DFFRHQX1 memory_reg_35__14_ ( .D(n2073), .CK(clk), .RN(rstn), .Q(memory[462]) );
  DFFRHQX1 memory_reg_35__13_ ( .D(n2074), .CK(clk), .RN(rstn), .Q(memory[461]) );
  DFFRHQX1 memory_reg_35__12_ ( .D(n2075), .CK(clk), .RN(rstn), .Q(memory[460]) );
  DFFRHQX1 memory_reg_35__11_ ( .D(n2076), .CK(clk), .RN(rstn), .Q(memory[459]) );
  DFFRHQX1 memory_reg_35__10_ ( .D(n2077), .CK(clk), .RN(rstn), .Q(memory[458]) );
  DFFRHQX1 memory_reg_35__9_ ( .D(n2078), .CK(clk), .RN(rstn), .Q(memory[457])
         );
  DFFRHQX1 memory_reg_35__8_ ( .D(n2079), .CK(clk), .RN(rstn), .Q(memory[456])
         );
  DFFRHQX1 memory_reg_35__7_ ( .D(n2080), .CK(clk), .RN(rstn), .Q(memory[455])
         );
  DFFRHQX1 memory_reg_35__6_ ( .D(n2081), .CK(clk), .RN(rstn), .Q(memory[454])
         );
  DFFRHQX1 memory_reg_35__5_ ( .D(n2082), .CK(clk), .RN(rstn), .Q(memory[453])
         );
  DFFRHQX1 memory_reg_35__4_ ( .D(n2083), .CK(clk), .RN(rstn), .Q(memory[452])
         );
  DFFRHQX1 memory_reg_35__3_ ( .D(n2084), .CK(clk), .RN(rstn), .Q(memory[451])
         );
  DFFRHQX1 memory_reg_35__2_ ( .D(n2085), .CK(clk), .RN(rstn), .Q(memory[450])
         );
  DFFRHQX1 memory_reg_35__1_ ( .D(n2086), .CK(clk), .RN(rstn), .Q(memory[449])
         );
  DFFRHQX1 memory_reg_35__0_ ( .D(n2087), .CK(clk), .RN(rstn), .Q(memory[448])
         );
  DFFRHQX1 memory_reg_39__15_ ( .D(n2136), .CK(clk), .RN(rstn), .Q(memory[399]) );
  DFFRHQX1 memory_reg_39__14_ ( .D(n2137), .CK(clk), .RN(rstn), .Q(memory[398]) );
  DFFRHQX1 memory_reg_39__13_ ( .D(n2138), .CK(clk), .RN(rstn), .Q(memory[397]) );
  DFFRHQX1 memory_reg_39__12_ ( .D(n2139), .CK(clk), .RN(rstn), .Q(memory[396]) );
  DFFRHQX1 memory_reg_39__11_ ( .D(n2140), .CK(clk), .RN(rstn), .Q(memory[395]) );
  DFFRHQX1 memory_reg_39__10_ ( .D(n2141), .CK(clk), .RN(rstn), .Q(memory[394]) );
  DFFRHQX1 memory_reg_39__9_ ( .D(n2142), .CK(clk), .RN(rstn), .Q(memory[393])
         );
  DFFRHQX1 memory_reg_39__8_ ( .D(n2143), .CK(clk), .RN(rstn), .Q(memory[392])
         );
  DFFRHQX1 memory_reg_39__7_ ( .D(n2144), .CK(clk), .RN(rstn), .Q(memory[391])
         );
  DFFRHQX1 memory_reg_39__6_ ( .D(n2145), .CK(clk), .RN(rstn), .Q(memory[390])
         );
  DFFRHQX1 memory_reg_39__5_ ( .D(n2146), .CK(clk), .RN(rstn), .Q(memory[389])
         );
  DFFRHQX1 memory_reg_39__4_ ( .D(n2147), .CK(clk), .RN(rstn), .Q(memory[388])
         );
  DFFRHQX1 memory_reg_39__3_ ( .D(n2148), .CK(clk), .RN(rstn), .Q(memory[387])
         );
  DFFRHQX1 memory_reg_39__2_ ( .D(n2149), .CK(clk), .RN(rstn), .Q(memory[386])
         );
  DFFRHQX1 memory_reg_39__1_ ( .D(n2150), .CK(clk), .RN(rstn), .Q(memory[385])
         );
  DFFRHQX1 memory_reg_39__0_ ( .D(n2151), .CK(clk), .RN(rstn), .Q(memory[384])
         );
  DFFRHQX1 memory_reg_43__15_ ( .D(n2200), .CK(clk), .RN(rstn), .Q(memory[335]) );
  DFFRHQX1 memory_reg_43__14_ ( .D(n2201), .CK(clk), .RN(rstn), .Q(memory[334]) );
  DFFRHQX1 memory_reg_43__13_ ( .D(n2202), .CK(clk), .RN(rstn), .Q(memory[333]) );
  DFFRHQX1 memory_reg_43__12_ ( .D(n2203), .CK(clk), .RN(rstn), .Q(memory[332]) );
  DFFRHQX1 memory_reg_43__11_ ( .D(n2204), .CK(clk), .RN(rstn), .Q(memory[331]) );
  DFFRHQX1 memory_reg_43__10_ ( .D(n2205), .CK(clk), .RN(rstn), .Q(memory[330]) );
  DFFRHQX1 memory_reg_43__9_ ( .D(n2206), .CK(clk), .RN(rstn), .Q(memory[329])
         );
  DFFRHQX1 memory_reg_43__8_ ( .D(n2207), .CK(clk), .RN(rstn), .Q(memory[328])
         );
  DFFRHQX1 memory_reg_43__7_ ( .D(n2208), .CK(clk), .RN(rstn), .Q(memory[327])
         );
  DFFRHQX1 memory_reg_43__6_ ( .D(n2209), .CK(clk), .RN(rstn), .Q(memory[326])
         );
  DFFRHQX1 memory_reg_43__5_ ( .D(n2210), .CK(clk), .RN(rstn), .Q(memory[325])
         );
  DFFRHQX1 memory_reg_43__4_ ( .D(n2211), .CK(clk), .RN(rstn), .Q(memory[324])
         );
  DFFRHQX1 memory_reg_43__3_ ( .D(n2212), .CK(clk), .RN(rstn), .Q(memory[323])
         );
  DFFRHQX1 memory_reg_43__2_ ( .D(n2213), .CK(clk), .RN(rstn), .Q(memory[322])
         );
  DFFRHQX1 memory_reg_43__1_ ( .D(n2214), .CK(clk), .RN(rstn), .Q(memory[321])
         );
  DFFRHQX1 memory_reg_43__0_ ( .D(n2215), .CK(clk), .RN(rstn), .Q(memory[320])
         );
  DFFRHQX1 memory_reg_47__15_ ( .D(n2264), .CK(clk), .RN(rstn), .Q(memory[271]) );
  DFFRHQX1 memory_reg_47__14_ ( .D(n2265), .CK(clk), .RN(rstn), .Q(memory[270]) );
  DFFRHQX1 memory_reg_47__13_ ( .D(n2266), .CK(clk), .RN(rstn), .Q(memory[269]) );
  DFFRHQX1 memory_reg_47__12_ ( .D(n2267), .CK(clk), .RN(rstn), .Q(memory[268]) );
  DFFRHQX1 memory_reg_47__11_ ( .D(n2268), .CK(clk), .RN(rstn), .Q(memory[267]) );
  DFFRHQX1 memory_reg_47__10_ ( .D(n2269), .CK(clk), .RN(rstn), .Q(memory[266]) );
  DFFRHQX1 memory_reg_47__9_ ( .D(n2270), .CK(clk), .RN(rstn), .Q(memory[265])
         );
  DFFRHQX1 memory_reg_47__8_ ( .D(n2271), .CK(clk), .RN(rstn), .Q(memory[264])
         );
  DFFRHQX1 memory_reg_47__7_ ( .D(n2272), .CK(clk), .RN(rstn), .Q(memory[263])
         );
  DFFRHQX1 memory_reg_47__6_ ( .D(n2273), .CK(clk), .RN(rstn), .Q(memory[262])
         );
  DFFRHQX1 memory_reg_47__5_ ( .D(n2274), .CK(clk), .RN(rstn), .Q(memory[261])
         );
  DFFRHQX1 memory_reg_47__4_ ( .D(n2275), .CK(clk), .RN(rstn), .Q(memory[260])
         );
  DFFRHQX1 memory_reg_47__3_ ( .D(n2276), .CK(clk), .RN(rstn), .Q(memory[259])
         );
  DFFRHQX1 memory_reg_47__2_ ( .D(n2277), .CK(clk), .RN(rstn), .Q(memory[258])
         );
  DFFRHQX1 memory_reg_47__1_ ( .D(n2278), .CK(clk), .RN(rstn), .Q(memory[257])
         );
  DFFRHQX1 memory_reg_47__0_ ( .D(n2279), .CK(clk), .RN(rstn), .Q(memory[256])
         );
  DFFRHQX1 memory_reg_51__15_ ( .D(n2328), .CK(clk), .RN(rstn), .Q(memory[207]) );
  DFFRHQX1 memory_reg_51__14_ ( .D(n2329), .CK(clk), .RN(rstn), .Q(memory[206]) );
  DFFRHQX1 memory_reg_51__13_ ( .D(n2330), .CK(clk), .RN(rstn), .Q(memory[205]) );
  DFFRHQX1 memory_reg_51__12_ ( .D(n2331), .CK(clk), .RN(rstn), .Q(memory[204]) );
  DFFRHQX1 memory_reg_51__11_ ( .D(n2332), .CK(clk), .RN(rstn), .Q(memory[203]) );
  DFFRHQX1 memory_reg_51__10_ ( .D(n2333), .CK(clk), .RN(rstn), .Q(memory[202]) );
  DFFRHQX1 memory_reg_51__9_ ( .D(n2334), .CK(clk), .RN(rstn), .Q(memory[201])
         );
  DFFRHQX1 memory_reg_51__8_ ( .D(n2335), .CK(clk), .RN(rstn), .Q(memory[200])
         );
  DFFRHQX1 memory_reg_51__7_ ( .D(n2336), .CK(clk), .RN(rstn), .Q(memory[199])
         );
  DFFRHQX1 memory_reg_51__6_ ( .D(n2337), .CK(clk), .RN(rstn), .Q(memory[198])
         );
  DFFRHQX1 memory_reg_51__5_ ( .D(n2338), .CK(clk), .RN(rstn), .Q(memory[197])
         );
  DFFRHQX1 memory_reg_51__4_ ( .D(n2339), .CK(clk), .RN(rstn), .Q(memory[196])
         );
  DFFRHQX1 memory_reg_51__3_ ( .D(n2340), .CK(clk), .RN(rstn), .Q(memory[195])
         );
  DFFRHQX1 memory_reg_51__2_ ( .D(n2341), .CK(clk), .RN(rstn), .Q(memory[194])
         );
  DFFRHQX1 memory_reg_51__1_ ( .D(n2342), .CK(clk), .RN(rstn), .Q(memory[193])
         );
  DFFRHQX1 memory_reg_51__0_ ( .D(n2343), .CK(clk), .RN(rstn), .Q(memory[192])
         );
  DFFRHQX1 memory_reg_55__15_ ( .D(n2392), .CK(clk), .RN(rstn), .Q(memory[143]) );
  DFFRHQX1 memory_reg_55__14_ ( .D(n2393), .CK(clk), .RN(rstn), .Q(memory[142]) );
  DFFRHQX1 memory_reg_55__13_ ( .D(n2394), .CK(clk), .RN(rstn), .Q(memory[141]) );
  DFFRHQX1 memory_reg_55__12_ ( .D(n2395), .CK(clk), .RN(rstn), .Q(memory[140]) );
  DFFRHQX1 memory_reg_55__11_ ( .D(n2396), .CK(clk), .RN(rstn), .Q(memory[139]) );
  DFFRHQX1 memory_reg_55__10_ ( .D(n2397), .CK(clk), .RN(rstn), .Q(memory[138]) );
  DFFRHQX1 memory_reg_55__9_ ( .D(n2398), .CK(clk), .RN(rstn), .Q(memory[137])
         );
  DFFRHQX1 memory_reg_55__8_ ( .D(n2399), .CK(clk), .RN(rstn), .Q(memory[136])
         );
  DFFRHQX1 memory_reg_55__7_ ( .D(n2400), .CK(clk), .RN(rstn), .Q(memory[135])
         );
  DFFRHQX1 memory_reg_55__6_ ( .D(n2401), .CK(clk), .RN(rstn), .Q(memory[134])
         );
  DFFRHQX1 memory_reg_55__5_ ( .D(n2402), .CK(clk), .RN(rstn), .Q(memory[133])
         );
  DFFRHQX1 memory_reg_55__4_ ( .D(n2403), .CK(clk), .RN(rstn), .Q(memory[132])
         );
  DFFRHQX1 memory_reg_55__3_ ( .D(n2404), .CK(clk), .RN(rstn), .Q(memory[131])
         );
  DFFRHQX1 memory_reg_55__2_ ( .D(n2405), .CK(clk), .RN(rstn), .Q(memory[130])
         );
  DFFRHQX1 memory_reg_55__1_ ( .D(n2406), .CK(clk), .RN(rstn), .Q(memory[129])
         );
  DFFRHQX1 memory_reg_55__0_ ( .D(n2407), .CK(clk), .RN(rstn), .Q(memory[128])
         );
  DFFRHQX1 memory_reg_59__15_ ( .D(n2456), .CK(clk), .RN(rstn), .Q(memory[79])
         );
  DFFRHQX1 memory_reg_59__14_ ( .D(n2457), .CK(clk), .RN(rstn), .Q(memory[78])
         );
  DFFRHQX1 memory_reg_59__13_ ( .D(n2458), .CK(clk), .RN(rstn), .Q(memory[77])
         );
  DFFRHQX1 memory_reg_59__12_ ( .D(n2459), .CK(clk), .RN(rstn), .Q(memory[76])
         );
  DFFRHQX1 memory_reg_59__11_ ( .D(n2460), .CK(clk), .RN(rstn), .Q(memory[75])
         );
  DFFRHQX1 memory_reg_59__10_ ( .D(n2461), .CK(clk), .RN(rstn), .Q(memory[74])
         );
  DFFRHQX1 memory_reg_59__9_ ( .D(n2462), .CK(clk), .RN(rstn), .Q(memory[73])
         );
  DFFRHQX1 memory_reg_59__8_ ( .D(n2463), .CK(clk), .RN(rstn), .Q(memory[72])
         );
  DFFRHQX1 memory_reg_59__7_ ( .D(n2464), .CK(clk), .RN(rstn), .Q(memory[71])
         );
  DFFRHQX1 memory_reg_59__6_ ( .D(n2465), .CK(clk), .RN(rstn), .Q(memory[70])
         );
  DFFRHQX1 memory_reg_59__5_ ( .D(n2466), .CK(clk), .RN(rstn), .Q(memory[69])
         );
  DFFRHQX1 memory_reg_59__4_ ( .D(n2467), .CK(clk), .RN(rstn), .Q(memory[68])
         );
  DFFRHQX1 memory_reg_59__3_ ( .D(n2468), .CK(clk), .RN(rstn), .Q(memory[67])
         );
  DFFRHQX1 memory_reg_59__2_ ( .D(n2469), .CK(clk), .RN(rstn), .Q(memory[66])
         );
  DFFRHQX1 memory_reg_59__1_ ( .D(n2470), .CK(clk), .RN(rstn), .Q(memory[65])
         );
  DFFRHQX1 memory_reg_59__0_ ( .D(n2471), .CK(clk), .RN(rstn), .Q(memory[64])
         );
  DFFRHQX1 memory_reg_63__15_ ( .D(n2520), .CK(clk), .RN(rstn), .Q(memory[15])
         );
  DFFRHQX1 memory_reg_63__14_ ( .D(n2521), .CK(clk), .RN(rstn), .Q(memory[14])
         );
  DFFRHQX1 memory_reg_63__13_ ( .D(n2522), .CK(clk), .RN(rstn), .Q(memory[13])
         );
  DFFRHQX1 memory_reg_63__12_ ( .D(n2523), .CK(clk), .RN(rstn), .Q(memory[12])
         );
  DFFRHQX1 memory_reg_63__11_ ( .D(n2524), .CK(clk), .RN(rstn), .Q(memory[11])
         );
  DFFRHQX1 memory_reg_63__10_ ( .D(n2525), .CK(clk), .RN(rstn), .Q(memory[10])
         );
  DFFRHQX1 memory_reg_63__9_ ( .D(n2526), .CK(clk), .RN(rstn), .Q(memory[9])
         );
  DFFRHQX1 memory_reg_63__8_ ( .D(n2527), .CK(clk), .RN(rstn), .Q(memory[8])
         );
  DFFRHQX1 memory_reg_63__7_ ( .D(n2528), .CK(clk), .RN(rstn), .Q(memory[7])
         );
  DFFRHQX1 memory_reg_63__6_ ( .D(n2529), .CK(clk), .RN(rstn), .Q(memory[6])
         );
  DFFRHQX1 memory_reg_63__5_ ( .D(n2530), .CK(clk), .RN(rstn), .Q(memory[5])
         );
  DFFRHQX1 memory_reg_63__4_ ( .D(n2531), .CK(clk), .RN(rstn), .Q(memory[4])
         );
  DFFRHQX1 memory_reg_63__3_ ( .D(n2532), .CK(clk), .RN(rstn), .Q(memory[3])
         );
  DFFRHQX1 memory_reg_63__2_ ( .D(n2533), .CK(clk), .RN(rstn), .Q(memory[2])
         );
  DFFRHQX1 memory_reg_63__1_ ( .D(n2534), .CK(clk), .RN(rstn), .Q(memory[1])
         );
  DFFRHQX1 memory_reg_63__0_ ( .D(n2535), .CK(clk), .RN(rstn), .Q(memory[0])
         );
  DFFRHQX1 memory_reg_0__15_ ( .D(n1512), .CK(clk), .RN(rstn), .Q(memory[1023]) );
  DFFRHQX1 memory_reg_0__14_ ( .D(n1513), .CK(clk), .RN(rstn), .Q(memory[1022]) );
  DFFRHQX1 memory_reg_0__13_ ( .D(n1514), .CK(clk), .RN(rstn), .Q(memory[1021]) );
  DFFRHQX1 memory_reg_0__12_ ( .D(n1515), .CK(clk), .RN(rstn), .Q(memory[1020]) );
  DFFRHQX1 memory_reg_0__11_ ( .D(n1516), .CK(clk), .RN(rstn), .Q(memory[1019]) );
  DFFRHQX1 memory_reg_0__10_ ( .D(n1517), .CK(clk), .RN(rstn), .Q(memory[1018]) );
  DFFRHQX1 memory_reg_0__9_ ( .D(n1518), .CK(clk), .RN(rstn), .Q(memory[1017])
         );
  DFFRHQX1 memory_reg_0__8_ ( .D(n1519), .CK(clk), .RN(rstn), .Q(memory[1016])
         );
  DFFRHQX1 memory_reg_0__7_ ( .D(n1520), .CK(clk), .RN(rstn), .Q(memory[1015])
         );
  DFFRHQX1 memory_reg_0__6_ ( .D(n1521), .CK(clk), .RN(rstn), .Q(memory[1014])
         );
  DFFRHQX1 memory_reg_0__5_ ( .D(n1522), .CK(clk), .RN(rstn), .Q(memory[1013])
         );
  DFFRHQX1 memory_reg_0__4_ ( .D(n1523), .CK(clk), .RN(rstn), .Q(memory[1012])
         );
  DFFRHQX1 memory_reg_0__3_ ( .D(n1524), .CK(clk), .RN(rstn), .Q(memory[1011])
         );
  DFFRHQX1 memory_reg_0__2_ ( .D(n1525), .CK(clk), .RN(rstn), .Q(memory[1010])
         );
  DFFRHQX1 memory_reg_0__1_ ( .D(n1526), .CK(clk), .RN(rstn), .Q(memory[1009])
         );
  DFFRHQX1 memory_reg_0__0_ ( .D(n1527), .CK(clk), .RN(rstn), .Q(memory[1008])
         );
  DFFRHQX1 memory_reg_4__15_ ( .D(n1576), .CK(clk), .RN(rstn), .Q(memory[959])
         );
  DFFRHQX1 memory_reg_4__14_ ( .D(n1577), .CK(clk), .RN(rstn), .Q(memory[958])
         );
  DFFRHQX1 memory_reg_4__13_ ( .D(n1578), .CK(clk), .RN(rstn), .Q(memory[957])
         );
  DFFRHQX1 memory_reg_4__12_ ( .D(n1579), .CK(clk), .RN(rstn), .Q(memory[956])
         );
  DFFRHQX1 memory_reg_4__11_ ( .D(n1580), .CK(clk), .RN(rstn), .Q(memory[955])
         );
  DFFRHQX1 memory_reg_4__10_ ( .D(n1581), .CK(clk), .RN(rstn), .Q(memory[954])
         );
  DFFRHQX1 memory_reg_4__9_ ( .D(n1582), .CK(clk), .RN(rstn), .Q(memory[953])
         );
  DFFRHQX1 memory_reg_4__8_ ( .D(n1583), .CK(clk), .RN(rstn), .Q(memory[952])
         );
  DFFRHQX1 memory_reg_4__7_ ( .D(n1584), .CK(clk), .RN(rstn), .Q(memory[951])
         );
  DFFRHQX1 memory_reg_4__6_ ( .D(n1585), .CK(clk), .RN(rstn), .Q(memory[950])
         );
  DFFRHQX1 memory_reg_4__5_ ( .D(n1586), .CK(clk), .RN(rstn), .Q(memory[949])
         );
  DFFRHQX1 memory_reg_4__4_ ( .D(n1587), .CK(clk), .RN(rstn), .Q(memory[948])
         );
  DFFRHQX1 memory_reg_4__3_ ( .D(n1588), .CK(clk), .RN(rstn), .Q(memory[947])
         );
  DFFRHQX1 memory_reg_4__2_ ( .D(n1589), .CK(clk), .RN(rstn), .Q(memory[946])
         );
  DFFRHQX1 memory_reg_4__1_ ( .D(n1590), .CK(clk), .RN(rstn), .Q(memory[945])
         );
  DFFRHQX1 memory_reg_4__0_ ( .D(n1591), .CK(clk), .RN(rstn), .Q(memory[944])
         );
  DFFRHQX1 memory_reg_8__15_ ( .D(n1640), .CK(clk), .RN(rstn), .Q(memory[895])
         );
  DFFRHQX1 memory_reg_8__14_ ( .D(n1641), .CK(clk), .RN(rstn), .Q(memory[894])
         );
  DFFRHQX1 memory_reg_8__13_ ( .D(n1642), .CK(clk), .RN(rstn), .Q(memory[893])
         );
  DFFRHQX1 memory_reg_8__12_ ( .D(n1643), .CK(clk), .RN(rstn), .Q(memory[892])
         );
  DFFRHQX1 memory_reg_8__11_ ( .D(n1644), .CK(clk), .RN(rstn), .Q(memory[891])
         );
  DFFRHQX1 memory_reg_8__10_ ( .D(n1645), .CK(clk), .RN(rstn), .Q(memory[890])
         );
  DFFRHQX1 memory_reg_8__9_ ( .D(n1646), .CK(clk), .RN(rstn), .Q(memory[889])
         );
  DFFRHQX1 memory_reg_8__8_ ( .D(n1647), .CK(clk), .RN(rstn), .Q(memory[888])
         );
  DFFRHQX1 memory_reg_8__7_ ( .D(n1648), .CK(clk), .RN(rstn), .Q(memory[887])
         );
  DFFRHQX1 memory_reg_8__6_ ( .D(n1649), .CK(clk), .RN(rstn), .Q(memory[886])
         );
  DFFRHQX1 memory_reg_8__5_ ( .D(n1650), .CK(clk), .RN(rstn), .Q(memory[885])
         );
  DFFRHQX1 memory_reg_8__4_ ( .D(n1651), .CK(clk), .RN(rstn), .Q(memory[884])
         );
  DFFRHQX1 memory_reg_8__3_ ( .D(n1652), .CK(clk), .RN(rstn), .Q(memory[883])
         );
  DFFRHQX1 memory_reg_8__2_ ( .D(n1653), .CK(clk), .RN(rstn), .Q(memory[882])
         );
  DFFRHQX1 memory_reg_8__1_ ( .D(n1654), .CK(clk), .RN(rstn), .Q(memory[881])
         );
  DFFRHQX1 memory_reg_8__0_ ( .D(n1655), .CK(clk), .RN(rstn), .Q(memory[880])
         );
  DFFRHQX1 memory_reg_12__15_ ( .D(n1704), .CK(clk), .RN(rstn), .Q(memory[831]) );
  DFFRHQX1 memory_reg_12__14_ ( .D(n1705), .CK(clk), .RN(rstn), .Q(memory[830]) );
  DFFRHQX1 memory_reg_12__13_ ( .D(n1706), .CK(clk), .RN(rstn), .Q(memory[829]) );
  DFFRHQX1 memory_reg_12__12_ ( .D(n1707), .CK(clk), .RN(rstn), .Q(memory[828]) );
  DFFRHQX1 memory_reg_12__11_ ( .D(n1708), .CK(clk), .RN(rstn), .Q(memory[827]) );
  DFFRHQX1 memory_reg_12__10_ ( .D(n1709), .CK(clk), .RN(rstn), .Q(memory[826]) );
  DFFRHQX1 memory_reg_12__9_ ( .D(n1710), .CK(clk), .RN(rstn), .Q(memory[825])
         );
  DFFRHQX1 memory_reg_12__8_ ( .D(n1711), .CK(clk), .RN(rstn), .Q(memory[824])
         );
  DFFRHQX1 memory_reg_12__7_ ( .D(n1712), .CK(clk), .RN(rstn), .Q(memory[823])
         );
  DFFRHQX1 memory_reg_12__6_ ( .D(n1713), .CK(clk), .RN(rstn), .Q(memory[822])
         );
  DFFRHQX1 memory_reg_12__5_ ( .D(n1714), .CK(clk), .RN(rstn), .Q(memory[821])
         );
  DFFRHQX1 memory_reg_12__4_ ( .D(n1715), .CK(clk), .RN(rstn), .Q(memory[820])
         );
  DFFRHQX1 memory_reg_12__3_ ( .D(n1716), .CK(clk), .RN(rstn), .Q(memory[819])
         );
  DFFRHQX1 memory_reg_12__2_ ( .D(n1717), .CK(clk), .RN(rstn), .Q(memory[818])
         );
  DFFRHQX1 memory_reg_12__1_ ( .D(n1718), .CK(clk), .RN(rstn), .Q(memory[817])
         );
  DFFRHQX1 memory_reg_12__0_ ( .D(n1719), .CK(clk), .RN(rstn), .Q(memory[816])
         );
  DFFRHQX1 memory_reg_16__15_ ( .D(n1768), .CK(clk), .RN(rstn), .Q(memory[767]) );
  DFFRHQX1 memory_reg_16__14_ ( .D(n1769), .CK(clk), .RN(rstn), .Q(memory[766]) );
  DFFRHQX1 memory_reg_16__13_ ( .D(n1770), .CK(clk), .RN(rstn), .Q(memory[765]) );
  DFFRHQX1 memory_reg_16__12_ ( .D(n1771), .CK(clk), .RN(rstn), .Q(memory[764]) );
  DFFRHQX1 memory_reg_16__11_ ( .D(n1772), .CK(clk), .RN(rstn), .Q(memory[763]) );
  DFFRHQX1 memory_reg_16__10_ ( .D(n1773), .CK(clk), .RN(rstn), .Q(memory[762]) );
  DFFRHQX1 memory_reg_16__9_ ( .D(n1774), .CK(clk), .RN(rstn), .Q(memory[761])
         );
  DFFRHQX1 memory_reg_16__8_ ( .D(n1775), .CK(clk), .RN(rstn), .Q(memory[760])
         );
  DFFRHQX1 memory_reg_16__7_ ( .D(n1776), .CK(clk), .RN(rstn), .Q(memory[759])
         );
  DFFRHQX1 memory_reg_16__6_ ( .D(n1777), .CK(clk), .RN(rstn), .Q(memory[758])
         );
  DFFRHQX1 memory_reg_16__5_ ( .D(n1778), .CK(clk), .RN(rstn), .Q(memory[757])
         );
  DFFRHQX1 memory_reg_16__4_ ( .D(n1779), .CK(clk), .RN(rstn), .Q(memory[756])
         );
  DFFRHQX1 memory_reg_16__3_ ( .D(n1780), .CK(clk), .RN(rstn), .Q(memory[755])
         );
  DFFRHQX1 memory_reg_16__2_ ( .D(n1781), .CK(clk), .RN(rstn), .Q(memory[754])
         );
  DFFRHQX1 memory_reg_16__1_ ( .D(n1782), .CK(clk), .RN(rstn), .Q(memory[753])
         );
  DFFRHQX1 memory_reg_16__0_ ( .D(n1783), .CK(clk), .RN(rstn), .Q(memory[752])
         );
  DFFRHQX1 memory_reg_20__15_ ( .D(n1832), .CK(clk), .RN(rstn), .Q(memory[703]) );
  DFFRHQX1 memory_reg_20__14_ ( .D(n1833), .CK(clk), .RN(rstn), .Q(memory[702]) );
  DFFRHQX1 memory_reg_20__13_ ( .D(n1834), .CK(clk), .RN(rstn), .Q(memory[701]) );
  DFFRHQX1 memory_reg_20__12_ ( .D(n1835), .CK(clk), .RN(rstn), .Q(memory[700]) );
  DFFRHQX1 memory_reg_20__11_ ( .D(n1836), .CK(clk), .RN(rstn), .Q(memory[699]) );
  DFFRHQX1 memory_reg_20__10_ ( .D(n1837), .CK(clk), .RN(rstn), .Q(memory[698]) );
  DFFRHQX1 memory_reg_20__9_ ( .D(n1838), .CK(clk), .RN(rstn), .Q(memory[697])
         );
  DFFRHQX1 memory_reg_20__8_ ( .D(n1839), .CK(clk), .RN(rstn), .Q(memory[696])
         );
  DFFRHQX1 memory_reg_20__7_ ( .D(n1840), .CK(clk), .RN(rstn), .Q(memory[695])
         );
  DFFRHQX1 memory_reg_20__6_ ( .D(n1841), .CK(clk), .RN(rstn), .Q(memory[694])
         );
  DFFRHQX1 memory_reg_20__5_ ( .D(n1842), .CK(clk), .RN(rstn), .Q(memory[693])
         );
  DFFRHQX1 memory_reg_20__4_ ( .D(n1843), .CK(clk), .RN(rstn), .Q(memory[692])
         );
  DFFRHQX1 memory_reg_20__3_ ( .D(n1844), .CK(clk), .RN(rstn), .Q(memory[691])
         );
  DFFRHQX1 memory_reg_20__2_ ( .D(n1845), .CK(clk), .RN(rstn), .Q(memory[690])
         );
  DFFRHQX1 memory_reg_20__1_ ( .D(n1846), .CK(clk), .RN(rstn), .Q(memory[689])
         );
  DFFRHQX1 memory_reg_20__0_ ( .D(n1847), .CK(clk), .RN(rstn), .Q(memory[688])
         );
  DFFRHQX1 memory_reg_24__15_ ( .D(n1896), .CK(clk), .RN(rstn), .Q(memory[639]) );
  DFFRHQX1 memory_reg_24__14_ ( .D(n1897), .CK(clk), .RN(rstn), .Q(memory[638]) );
  DFFRHQX1 memory_reg_24__13_ ( .D(n1898), .CK(clk), .RN(rstn), .Q(memory[637]) );
  DFFRHQX1 memory_reg_24__12_ ( .D(n1899), .CK(clk), .RN(rstn), .Q(memory[636]) );
  DFFRHQX1 memory_reg_24__11_ ( .D(n1900), .CK(clk), .RN(rstn), .Q(memory[635]) );
  DFFRHQX1 memory_reg_24__10_ ( .D(n1901), .CK(clk), .RN(rstn), .Q(memory[634]) );
  DFFRHQX1 memory_reg_24__9_ ( .D(n1902), .CK(clk), .RN(rstn), .Q(memory[633])
         );
  DFFRHQX1 memory_reg_24__8_ ( .D(n1903), .CK(clk), .RN(rstn), .Q(memory[632])
         );
  DFFRHQX1 memory_reg_24__7_ ( .D(n1904), .CK(clk), .RN(rstn), .Q(memory[631])
         );
  DFFRHQX1 memory_reg_24__6_ ( .D(n1905), .CK(clk), .RN(rstn), .Q(memory[630])
         );
  DFFRHQX1 memory_reg_24__5_ ( .D(n1906), .CK(clk), .RN(rstn), .Q(memory[629])
         );
  DFFRHQX1 memory_reg_24__4_ ( .D(n1907), .CK(clk), .RN(rstn), .Q(memory[628])
         );
  DFFRHQX1 memory_reg_24__3_ ( .D(n1908), .CK(clk), .RN(rstn), .Q(memory[627])
         );
  DFFRHQX1 memory_reg_24__2_ ( .D(n1909), .CK(clk), .RN(rstn), .Q(memory[626])
         );
  DFFRHQX1 memory_reg_24__1_ ( .D(n1910), .CK(clk), .RN(rstn), .Q(memory[625])
         );
  DFFRHQX1 memory_reg_24__0_ ( .D(n1911), .CK(clk), .RN(rstn), .Q(memory[624])
         );
  DFFRHQX1 memory_reg_28__15_ ( .D(n1960), .CK(clk), .RN(rstn), .Q(memory[575]) );
  DFFRHQX1 memory_reg_28__14_ ( .D(n1961), .CK(clk), .RN(rstn), .Q(memory[574]) );
  DFFRHQX1 memory_reg_28__13_ ( .D(n1962), .CK(clk), .RN(rstn), .Q(memory[573]) );
  DFFRHQX1 memory_reg_28__12_ ( .D(n1963), .CK(clk), .RN(rstn), .Q(memory[572]) );
  DFFRHQX1 memory_reg_28__11_ ( .D(n1964), .CK(clk), .RN(rstn), .Q(memory[571]) );
  DFFRHQX1 memory_reg_28__10_ ( .D(n1965), .CK(clk), .RN(rstn), .Q(memory[570]) );
  DFFRHQX1 memory_reg_28__9_ ( .D(n1966), .CK(clk), .RN(rstn), .Q(memory[569])
         );
  DFFRHQX1 memory_reg_28__8_ ( .D(n1967), .CK(clk), .RN(rstn), .Q(memory[568])
         );
  DFFRHQX1 memory_reg_28__7_ ( .D(n1968), .CK(clk), .RN(rstn), .Q(memory[567])
         );
  DFFRHQX1 memory_reg_28__6_ ( .D(n1969), .CK(clk), .RN(rstn), .Q(memory[566])
         );
  DFFRHQX1 memory_reg_28__5_ ( .D(n1970), .CK(clk), .RN(rstn), .Q(memory[565])
         );
  DFFRHQX1 memory_reg_28__4_ ( .D(n1971), .CK(clk), .RN(rstn), .Q(memory[564])
         );
  DFFRHQX1 memory_reg_28__3_ ( .D(n1972), .CK(clk), .RN(rstn), .Q(memory[563])
         );
  DFFRHQX1 memory_reg_28__2_ ( .D(n1973), .CK(clk), .RN(rstn), .Q(memory[562])
         );
  DFFRHQX1 memory_reg_28__1_ ( .D(n1974), .CK(clk), .RN(rstn), .Q(memory[561])
         );
  DFFRHQX1 memory_reg_28__0_ ( .D(n1975), .CK(clk), .RN(rstn), .Q(memory[560])
         );
  DFFRHQX1 memory_reg_32__15_ ( .D(n2024), .CK(clk), .RN(rstn), .Q(memory[511]) );
  DFFRHQX1 memory_reg_32__14_ ( .D(n2025), .CK(clk), .RN(rstn), .Q(memory[510]) );
  DFFRHQX1 memory_reg_32__13_ ( .D(n2026), .CK(clk), .RN(rstn), .Q(memory[509]) );
  DFFRHQX1 memory_reg_32__12_ ( .D(n2027), .CK(clk), .RN(rstn), .Q(memory[508]) );
  DFFRHQX1 memory_reg_32__11_ ( .D(n2028), .CK(clk), .RN(rstn), .Q(memory[507]) );
  DFFRHQX1 memory_reg_32__10_ ( .D(n2029), .CK(clk), .RN(rstn), .Q(memory[506]) );
  DFFRHQX1 memory_reg_32__9_ ( .D(n2030), .CK(clk), .RN(rstn), .Q(memory[505])
         );
  DFFRHQX1 memory_reg_32__8_ ( .D(n2031), .CK(clk), .RN(rstn), .Q(memory[504])
         );
  DFFRHQX1 memory_reg_32__7_ ( .D(n2032), .CK(clk), .RN(rstn), .Q(memory[503])
         );
  DFFRHQX1 memory_reg_32__6_ ( .D(n2033), .CK(clk), .RN(rstn), .Q(memory[502])
         );
  DFFRHQX1 memory_reg_32__5_ ( .D(n2034), .CK(clk), .RN(rstn), .Q(memory[501])
         );
  DFFRHQX1 memory_reg_32__4_ ( .D(n2035), .CK(clk), .RN(rstn), .Q(memory[500])
         );
  DFFRHQX1 memory_reg_32__3_ ( .D(n2036), .CK(clk), .RN(rstn), .Q(memory[499])
         );
  DFFRHQX1 memory_reg_32__2_ ( .D(n2037), .CK(clk), .RN(rstn), .Q(memory[498])
         );
  DFFRHQX1 memory_reg_32__1_ ( .D(n2038), .CK(clk), .RN(rstn), .Q(memory[497])
         );
  DFFRHQX1 memory_reg_32__0_ ( .D(n2039), .CK(clk), .RN(rstn), .Q(memory[496])
         );
  DFFRHQX1 memory_reg_36__15_ ( .D(n2088), .CK(clk), .RN(rstn), .Q(memory[447]) );
  DFFRHQX1 memory_reg_36__14_ ( .D(n2089), .CK(clk), .RN(rstn), .Q(memory[446]) );
  DFFRHQX1 memory_reg_36__13_ ( .D(n2090), .CK(clk), .RN(rstn), .Q(memory[445]) );
  DFFRHQX1 memory_reg_36__12_ ( .D(n2091), .CK(clk), .RN(rstn), .Q(memory[444]) );
  DFFRHQX1 memory_reg_36__11_ ( .D(n2092), .CK(clk), .RN(rstn), .Q(memory[443]) );
  DFFRHQX1 memory_reg_36__10_ ( .D(n2093), .CK(clk), .RN(rstn), .Q(memory[442]) );
  DFFRHQX1 memory_reg_36__9_ ( .D(n2094), .CK(clk), .RN(rstn), .Q(memory[441])
         );
  DFFRHQX1 memory_reg_36__8_ ( .D(n2095), .CK(clk), .RN(rstn), .Q(memory[440])
         );
  DFFRHQX1 memory_reg_36__7_ ( .D(n2096), .CK(clk), .RN(rstn), .Q(memory[439])
         );
  DFFRHQX1 memory_reg_36__6_ ( .D(n2097), .CK(clk), .RN(rstn), .Q(memory[438])
         );
  DFFRHQX1 memory_reg_36__5_ ( .D(n2098), .CK(clk), .RN(rstn), .Q(memory[437])
         );
  DFFRHQX1 memory_reg_36__4_ ( .D(n2099), .CK(clk), .RN(rstn), .Q(memory[436])
         );
  DFFRHQX1 memory_reg_36__3_ ( .D(n2100), .CK(clk), .RN(rstn), .Q(memory[435])
         );
  DFFRHQX1 memory_reg_36__2_ ( .D(n2101), .CK(clk), .RN(rstn), .Q(memory[434])
         );
  DFFRHQX1 memory_reg_36__1_ ( .D(n2102), .CK(clk), .RN(rstn), .Q(memory[433])
         );
  DFFRHQX1 memory_reg_36__0_ ( .D(n2103), .CK(clk), .RN(rstn), .Q(memory[432])
         );
  DFFRHQX1 memory_reg_40__15_ ( .D(n2152), .CK(clk), .RN(rstn), .Q(memory[383]) );
  DFFRHQX1 memory_reg_40__14_ ( .D(n2153), .CK(clk), .RN(rstn), .Q(memory[382]) );
  DFFRHQX1 memory_reg_40__13_ ( .D(n2154), .CK(clk), .RN(rstn), .Q(memory[381]) );
  DFFRHQX1 memory_reg_40__12_ ( .D(n2155), .CK(clk), .RN(rstn), .Q(memory[380]) );
  DFFRHQX1 memory_reg_40__11_ ( .D(n2156), .CK(clk), .RN(rstn), .Q(memory[379]) );
  DFFRHQX1 memory_reg_40__10_ ( .D(n2157), .CK(clk), .RN(rstn), .Q(memory[378]) );
  DFFRHQX1 memory_reg_40__9_ ( .D(n2158), .CK(clk), .RN(rstn), .Q(memory[377])
         );
  DFFRHQX1 memory_reg_40__8_ ( .D(n2159), .CK(clk), .RN(rstn), .Q(memory[376])
         );
  DFFRHQX1 memory_reg_40__7_ ( .D(n2160), .CK(clk), .RN(rstn), .Q(memory[375])
         );
  DFFRHQX1 memory_reg_40__6_ ( .D(n2161), .CK(clk), .RN(rstn), .Q(memory[374])
         );
  DFFRHQX1 memory_reg_40__5_ ( .D(n2162), .CK(clk), .RN(rstn), .Q(memory[373])
         );
  DFFRHQX1 memory_reg_40__4_ ( .D(n2163), .CK(clk), .RN(rstn), .Q(memory[372])
         );
  DFFRHQX1 memory_reg_40__3_ ( .D(n2164), .CK(clk), .RN(rstn), .Q(memory[371])
         );
  DFFRHQX1 memory_reg_40__2_ ( .D(n2165), .CK(clk), .RN(rstn), .Q(memory[370])
         );
  DFFRHQX1 memory_reg_40__1_ ( .D(n2166), .CK(clk), .RN(rstn), .Q(memory[369])
         );
  DFFRHQX1 memory_reg_40__0_ ( .D(n2167), .CK(clk), .RN(rstn), .Q(memory[368])
         );
  DFFRHQX1 memory_reg_44__15_ ( .D(n2216), .CK(clk), .RN(rstn), .Q(memory[319]) );
  DFFRHQX1 memory_reg_44__14_ ( .D(n2217), .CK(clk), .RN(rstn), .Q(memory[318]) );
  DFFRHQX1 memory_reg_44__13_ ( .D(n2218), .CK(clk), .RN(rstn), .Q(memory[317]) );
  DFFRHQX1 memory_reg_44__12_ ( .D(n2219), .CK(clk), .RN(rstn), .Q(memory[316]) );
  DFFRHQX1 memory_reg_44__11_ ( .D(n2220), .CK(clk), .RN(rstn), .Q(memory[315]) );
  DFFRHQX1 memory_reg_44__10_ ( .D(n2221), .CK(clk), .RN(rstn), .Q(memory[314]) );
  DFFRHQX1 memory_reg_44__9_ ( .D(n2222), .CK(clk), .RN(rstn), .Q(memory[313])
         );
  DFFRHQX1 memory_reg_44__8_ ( .D(n2223), .CK(clk), .RN(rstn), .Q(memory[312])
         );
  DFFRHQX1 memory_reg_44__7_ ( .D(n2224), .CK(clk), .RN(rstn), .Q(memory[311])
         );
  DFFRHQX1 memory_reg_44__6_ ( .D(n2225), .CK(clk), .RN(rstn), .Q(memory[310])
         );
  DFFRHQX1 memory_reg_44__5_ ( .D(n2226), .CK(clk), .RN(rstn), .Q(memory[309])
         );
  DFFRHQX1 memory_reg_44__4_ ( .D(n2227), .CK(clk), .RN(rstn), .Q(memory[308])
         );
  DFFRHQX1 memory_reg_44__3_ ( .D(n2228), .CK(clk), .RN(rstn), .Q(memory[307])
         );
  DFFRHQX1 memory_reg_44__2_ ( .D(n2229), .CK(clk), .RN(rstn), .Q(memory[306])
         );
  DFFRHQX1 memory_reg_44__1_ ( .D(n2230), .CK(clk), .RN(rstn), .Q(memory[305])
         );
  DFFRHQX1 memory_reg_44__0_ ( .D(n2231), .CK(clk), .RN(rstn), .Q(memory[304])
         );
  DFFRHQX1 memory_reg_48__15_ ( .D(n2280), .CK(clk), .RN(rstn), .Q(memory[255]) );
  DFFRHQX1 memory_reg_48__14_ ( .D(n2281), .CK(clk), .RN(rstn), .Q(memory[254]) );
  DFFRHQX1 memory_reg_48__13_ ( .D(n2282), .CK(clk), .RN(rstn), .Q(memory[253]) );
  DFFRHQX1 memory_reg_48__12_ ( .D(n2283), .CK(clk), .RN(rstn), .Q(memory[252]) );
  DFFRHQX1 memory_reg_48__11_ ( .D(n2284), .CK(clk), .RN(rstn), .Q(memory[251]) );
  DFFRHQX1 memory_reg_48__10_ ( .D(n2285), .CK(clk), .RN(rstn), .Q(memory[250]) );
  DFFRHQX1 memory_reg_48__9_ ( .D(n2286), .CK(clk), .RN(rstn), .Q(memory[249])
         );
  DFFRHQX1 memory_reg_48__8_ ( .D(n2287), .CK(clk), .RN(rstn), .Q(memory[248])
         );
  DFFRHQX1 memory_reg_48__7_ ( .D(n2288), .CK(clk), .RN(rstn), .Q(memory[247])
         );
  DFFRHQX1 memory_reg_48__6_ ( .D(n2289), .CK(clk), .RN(rstn), .Q(memory[246])
         );
  DFFRHQX1 memory_reg_48__5_ ( .D(n2290), .CK(clk), .RN(rstn), .Q(memory[245])
         );
  DFFRHQX1 memory_reg_48__4_ ( .D(n2291), .CK(clk), .RN(rstn), .Q(memory[244])
         );
  DFFRHQX1 memory_reg_48__3_ ( .D(n2292), .CK(clk), .RN(rstn), .Q(memory[243])
         );
  DFFRHQX1 memory_reg_48__2_ ( .D(n2293), .CK(clk), .RN(rstn), .Q(memory[242])
         );
  DFFRHQX1 memory_reg_48__1_ ( .D(n2294), .CK(clk), .RN(rstn), .Q(memory[241])
         );
  DFFRHQX1 memory_reg_48__0_ ( .D(n2295), .CK(clk), .RN(rstn), .Q(memory[240])
         );
  DFFRHQX1 memory_reg_52__15_ ( .D(n2344), .CK(clk), .RN(rstn), .Q(memory[191]) );
  DFFRHQX1 memory_reg_52__14_ ( .D(n2345), .CK(clk), .RN(rstn), .Q(memory[190]) );
  DFFRHQX1 memory_reg_52__13_ ( .D(n2346), .CK(clk), .RN(rstn), .Q(memory[189]) );
  DFFRHQX1 memory_reg_52__12_ ( .D(n2347), .CK(clk), .RN(rstn), .Q(memory[188]) );
  DFFRHQX1 memory_reg_52__11_ ( .D(n2348), .CK(clk), .RN(rstn), .Q(memory[187]) );
  DFFRHQX1 memory_reg_52__10_ ( .D(n2349), .CK(clk), .RN(rstn), .Q(memory[186]) );
  DFFRHQX1 memory_reg_52__9_ ( .D(n2350), .CK(clk), .RN(rstn), .Q(memory[185])
         );
  DFFRHQX1 memory_reg_52__8_ ( .D(n2351), .CK(clk), .RN(rstn), .Q(memory[184])
         );
  DFFRHQX1 memory_reg_52__7_ ( .D(n2352), .CK(clk), .RN(rstn), .Q(memory[183])
         );
  DFFRHQX1 memory_reg_52__6_ ( .D(n2353), .CK(clk), .RN(rstn), .Q(memory[182])
         );
  DFFRHQX1 memory_reg_52__5_ ( .D(n2354), .CK(clk), .RN(rstn), .Q(memory[181])
         );
  DFFRHQX1 memory_reg_52__4_ ( .D(n2355), .CK(clk), .RN(rstn), .Q(memory[180])
         );
  DFFRHQX1 memory_reg_52__3_ ( .D(n2356), .CK(clk), .RN(rstn), .Q(memory[179])
         );
  DFFRHQX1 memory_reg_52__2_ ( .D(n2357), .CK(clk), .RN(rstn), .Q(memory[178])
         );
  DFFRHQX1 memory_reg_52__1_ ( .D(n2358), .CK(clk), .RN(rstn), .Q(memory[177])
         );
  DFFRHQX1 memory_reg_52__0_ ( .D(n2359), .CK(clk), .RN(rstn), .Q(memory[176])
         );
  DFFRHQX1 memory_reg_56__15_ ( .D(n2408), .CK(clk), .RN(rstn), .Q(memory[127]) );
  DFFRHQX1 memory_reg_56__14_ ( .D(n2409), .CK(clk), .RN(rstn), .Q(memory[126]) );
  DFFRHQX1 memory_reg_56__13_ ( .D(n2410), .CK(clk), .RN(rstn), .Q(memory[125]) );
  DFFRHQX1 memory_reg_56__12_ ( .D(n2411), .CK(clk), .RN(rstn), .Q(memory[124]) );
  DFFRHQX1 memory_reg_56__11_ ( .D(n2412), .CK(clk), .RN(rstn), .Q(memory[123]) );
  DFFRHQX1 memory_reg_56__10_ ( .D(n2413), .CK(clk), .RN(rstn), .Q(memory[122]) );
  DFFRHQX1 memory_reg_56__9_ ( .D(n2414), .CK(clk), .RN(rstn), .Q(memory[121])
         );
  DFFRHQX1 memory_reg_56__8_ ( .D(n2415), .CK(clk), .RN(rstn), .Q(memory[120])
         );
  DFFRHQX1 memory_reg_56__7_ ( .D(n2416), .CK(clk), .RN(rstn), .Q(memory[119])
         );
  DFFRHQX1 memory_reg_56__6_ ( .D(n2417), .CK(clk), .RN(rstn), .Q(memory[118])
         );
  DFFRHQX1 memory_reg_56__5_ ( .D(n2418), .CK(clk), .RN(rstn), .Q(memory[117])
         );
  DFFRHQX1 memory_reg_56__4_ ( .D(n2419), .CK(clk), .RN(rstn), .Q(memory[116])
         );
  DFFRHQX1 memory_reg_56__3_ ( .D(n2420), .CK(clk), .RN(rstn), .Q(memory[115])
         );
  DFFRHQX1 memory_reg_56__2_ ( .D(n2421), .CK(clk), .RN(rstn), .Q(memory[114])
         );
  DFFRHQX1 memory_reg_56__1_ ( .D(n2422), .CK(clk), .RN(rstn), .Q(memory[113])
         );
  DFFRHQX1 memory_reg_56__0_ ( .D(n2423), .CK(clk), .RN(rstn), .Q(memory[112])
         );
  DFFRHQX1 memory_reg_60__15_ ( .D(n2472), .CK(clk), .RN(rstn), .Q(memory[63])
         );
  DFFRHQX1 memory_reg_60__14_ ( .D(n2473), .CK(clk), .RN(rstn), .Q(memory[62])
         );
  DFFRHQX1 memory_reg_60__13_ ( .D(n2474), .CK(clk), .RN(rstn), .Q(memory[61])
         );
  DFFRHQX1 memory_reg_60__12_ ( .D(n2475), .CK(clk), .RN(rstn), .Q(memory[60])
         );
  DFFRHQX1 memory_reg_60__11_ ( .D(n2476), .CK(clk), .RN(rstn), .Q(memory[59])
         );
  DFFRHQX1 memory_reg_60__10_ ( .D(n2477), .CK(clk), .RN(rstn), .Q(memory[58])
         );
  DFFRHQX1 memory_reg_60__9_ ( .D(n2478), .CK(clk), .RN(rstn), .Q(memory[57])
         );
  DFFRHQX1 memory_reg_60__8_ ( .D(n2479), .CK(clk), .RN(rstn), .Q(memory[56])
         );
  DFFRHQX1 memory_reg_60__7_ ( .D(n2480), .CK(clk), .RN(rstn), .Q(memory[55])
         );
  DFFRHQX1 memory_reg_60__6_ ( .D(n2481), .CK(clk), .RN(rstn), .Q(memory[54])
         );
  DFFRHQX1 memory_reg_60__5_ ( .D(n2482), .CK(clk), .RN(rstn), .Q(memory[53])
         );
  DFFRHQX1 memory_reg_60__4_ ( .D(n2483), .CK(clk), .RN(rstn), .Q(memory[52])
         );
  DFFRHQX1 memory_reg_60__3_ ( .D(n2484), .CK(clk), .RN(rstn), .Q(memory[51])
         );
  DFFRHQX1 memory_reg_60__2_ ( .D(n2485), .CK(clk), .RN(rstn), .Q(memory[50])
         );
  DFFRHQX1 memory_reg_60__1_ ( .D(n2486), .CK(clk), .RN(rstn), .Q(memory[49])
         );
  DFFRHQX1 memory_reg_60__0_ ( .D(n2487), .CK(clk), .RN(rstn), .Q(memory[48])
         );
  DFFRHQX1 memory_reg_2__15_ ( .D(n1544), .CK(clk), .RN(rstn), .Q(memory[991])
         );
  DFFRHQX1 memory_reg_2__14_ ( .D(n1545), .CK(clk), .RN(rstn), .Q(memory[990])
         );
  DFFRHQX1 memory_reg_2__13_ ( .D(n1546), .CK(clk), .RN(rstn), .Q(memory[989])
         );
  DFFRHQX1 memory_reg_2__12_ ( .D(n1547), .CK(clk), .RN(rstn), .Q(memory[988])
         );
  DFFRHQX1 memory_reg_2__11_ ( .D(n1548), .CK(clk), .RN(rstn), .Q(memory[987])
         );
  DFFRHQX1 memory_reg_2__10_ ( .D(n1549), .CK(clk), .RN(rstn), .Q(memory[986])
         );
  DFFRHQX1 memory_reg_2__9_ ( .D(n1550), .CK(clk), .RN(rstn), .Q(memory[985])
         );
  DFFRHQX1 memory_reg_2__8_ ( .D(n1551), .CK(clk), .RN(rstn), .Q(memory[984])
         );
  DFFRHQX1 memory_reg_2__7_ ( .D(n1552), .CK(clk), .RN(rstn), .Q(memory[983])
         );
  DFFRHQX1 memory_reg_2__6_ ( .D(n1553), .CK(clk), .RN(rstn), .Q(memory[982])
         );
  DFFRHQX1 memory_reg_2__5_ ( .D(n1554), .CK(clk), .RN(rstn), .Q(memory[981])
         );
  DFFRHQX1 memory_reg_2__4_ ( .D(n1555), .CK(clk), .RN(rstn), .Q(memory[980])
         );
  DFFRHQX1 memory_reg_2__3_ ( .D(n1556), .CK(clk), .RN(rstn), .Q(memory[979])
         );
  DFFRHQX1 memory_reg_2__2_ ( .D(n1557), .CK(clk), .RN(rstn), .Q(memory[978])
         );
  DFFRHQX1 memory_reg_2__1_ ( .D(n1558), .CK(clk), .RN(rstn), .Q(memory[977])
         );
  DFFRHQX1 memory_reg_2__0_ ( .D(n1559), .CK(clk), .RN(rstn), .Q(memory[976])
         );
  DFFRHQX1 memory_reg_6__15_ ( .D(n1608), .CK(clk), .RN(rstn), .Q(memory[927])
         );
  DFFRHQX1 memory_reg_6__14_ ( .D(n1609), .CK(clk), .RN(rstn), .Q(memory[926])
         );
  DFFRHQX1 memory_reg_6__13_ ( .D(n1610), .CK(clk), .RN(rstn), .Q(memory[925])
         );
  DFFRHQX1 memory_reg_6__12_ ( .D(n1611), .CK(clk), .RN(rstn), .Q(memory[924])
         );
  DFFRHQX1 memory_reg_6__11_ ( .D(n1612), .CK(clk), .RN(rstn), .Q(memory[923])
         );
  DFFRHQX1 memory_reg_6__10_ ( .D(n1613), .CK(clk), .RN(rstn), .Q(memory[922])
         );
  DFFRHQX1 memory_reg_6__9_ ( .D(n1614), .CK(clk), .RN(rstn), .Q(memory[921])
         );
  DFFRHQX1 memory_reg_6__8_ ( .D(n1615), .CK(clk), .RN(rstn), .Q(memory[920])
         );
  DFFRHQX1 memory_reg_6__7_ ( .D(n1616), .CK(clk), .RN(rstn), .Q(memory[919])
         );
  DFFRHQX1 memory_reg_6__6_ ( .D(n1617), .CK(clk), .RN(rstn), .Q(memory[918])
         );
  DFFRHQX1 memory_reg_6__5_ ( .D(n1618), .CK(clk), .RN(rstn), .Q(memory[917])
         );
  DFFRHQX1 memory_reg_6__4_ ( .D(n1619), .CK(clk), .RN(rstn), .Q(memory[916])
         );
  DFFRHQX1 memory_reg_6__3_ ( .D(n1620), .CK(clk), .RN(rstn), .Q(memory[915])
         );
  DFFRHQX1 memory_reg_6__2_ ( .D(n1621), .CK(clk), .RN(rstn), .Q(memory[914])
         );
  DFFRHQX1 memory_reg_6__1_ ( .D(n1622), .CK(clk), .RN(rstn), .Q(memory[913])
         );
  DFFRHQX1 memory_reg_6__0_ ( .D(n1623), .CK(clk), .RN(rstn), .Q(memory[912])
         );
  DFFRHQX1 memory_reg_10__15_ ( .D(n1672), .CK(clk), .RN(rstn), .Q(memory[863]) );
  DFFRHQX1 memory_reg_10__14_ ( .D(n1673), .CK(clk), .RN(rstn), .Q(memory[862]) );
  DFFRHQX1 memory_reg_10__13_ ( .D(n1674), .CK(clk), .RN(rstn), .Q(memory[861]) );
  DFFRHQX1 memory_reg_10__12_ ( .D(n1675), .CK(clk), .RN(rstn), .Q(memory[860]) );
  DFFRHQX1 memory_reg_10__11_ ( .D(n1676), .CK(clk), .RN(rstn), .Q(memory[859]) );
  DFFRHQX1 memory_reg_10__10_ ( .D(n1677), .CK(clk), .RN(rstn), .Q(memory[858]) );
  DFFRHQX1 memory_reg_10__9_ ( .D(n1678), .CK(clk), .RN(rstn), .Q(memory[857])
         );
  DFFRHQX1 memory_reg_10__8_ ( .D(n1679), .CK(clk), .RN(rstn), .Q(memory[856])
         );
  DFFRHQX1 memory_reg_10__7_ ( .D(n1680), .CK(clk), .RN(rstn), .Q(memory[855])
         );
  DFFRHQX1 memory_reg_10__6_ ( .D(n1681), .CK(clk), .RN(rstn), .Q(memory[854])
         );
  DFFRHQX1 memory_reg_10__5_ ( .D(n1682), .CK(clk), .RN(rstn), .Q(memory[853])
         );
  DFFRHQX1 memory_reg_10__4_ ( .D(n1683), .CK(clk), .RN(rstn), .Q(memory[852])
         );
  DFFRHQX1 memory_reg_10__3_ ( .D(n1684), .CK(clk), .RN(rstn), .Q(memory[851])
         );
  DFFRHQX1 memory_reg_10__2_ ( .D(n1685), .CK(clk), .RN(rstn), .Q(memory[850])
         );
  DFFRHQX1 memory_reg_10__1_ ( .D(n1686), .CK(clk), .RN(rstn), .Q(memory[849])
         );
  DFFRHQX1 memory_reg_10__0_ ( .D(n1687), .CK(clk), .RN(rstn), .Q(memory[848])
         );
  DFFRHQX1 memory_reg_14__15_ ( .D(n1736), .CK(clk), .RN(rstn), .Q(memory[799]) );
  DFFRHQX1 memory_reg_14__14_ ( .D(n1737), .CK(clk), .RN(rstn), .Q(memory[798]) );
  DFFRHQX1 memory_reg_14__13_ ( .D(n1738), .CK(clk), .RN(rstn), .Q(memory[797]) );
  DFFRHQX1 memory_reg_14__12_ ( .D(n1739), .CK(clk), .RN(rstn), .Q(memory[796]) );
  DFFRHQX1 memory_reg_14__11_ ( .D(n1740), .CK(clk), .RN(rstn), .Q(memory[795]) );
  DFFRHQX1 memory_reg_14__10_ ( .D(n1741), .CK(clk), .RN(rstn), .Q(memory[794]) );
  DFFRHQX1 memory_reg_14__9_ ( .D(n1742), .CK(clk), .RN(rstn), .Q(memory[793])
         );
  DFFRHQX1 memory_reg_14__8_ ( .D(n1743), .CK(clk), .RN(rstn), .Q(memory[792])
         );
  DFFRHQX1 memory_reg_14__7_ ( .D(n1744), .CK(clk), .RN(rstn), .Q(memory[791])
         );
  DFFRHQX1 memory_reg_14__6_ ( .D(n1745), .CK(clk), .RN(rstn), .Q(memory[790])
         );
  DFFRHQX1 memory_reg_14__5_ ( .D(n1746), .CK(clk), .RN(rstn), .Q(memory[789])
         );
  DFFRHQX1 memory_reg_14__4_ ( .D(n1747), .CK(clk), .RN(rstn), .Q(memory[788])
         );
  DFFRHQX1 memory_reg_14__3_ ( .D(n1748), .CK(clk), .RN(rstn), .Q(memory[787])
         );
  DFFRHQX1 memory_reg_14__2_ ( .D(n1749), .CK(clk), .RN(rstn), .Q(memory[786])
         );
  DFFRHQX1 memory_reg_14__1_ ( .D(n1750), .CK(clk), .RN(rstn), .Q(memory[785])
         );
  DFFRHQX1 memory_reg_14__0_ ( .D(n1751), .CK(clk), .RN(rstn), .Q(memory[784])
         );
  DFFRHQX1 memory_reg_18__15_ ( .D(n1800), .CK(clk), .RN(rstn), .Q(memory[735]) );
  DFFRHQX1 memory_reg_18__14_ ( .D(n1801), .CK(clk), .RN(rstn), .Q(memory[734]) );
  DFFRHQX1 memory_reg_18__13_ ( .D(n1802), .CK(clk), .RN(rstn), .Q(memory[733]) );
  DFFRHQX1 memory_reg_18__12_ ( .D(n1803), .CK(clk), .RN(rstn), .Q(memory[732]) );
  DFFRHQX1 memory_reg_18__11_ ( .D(n1804), .CK(clk), .RN(rstn), .Q(memory[731]) );
  DFFRHQX1 memory_reg_18__10_ ( .D(n1805), .CK(clk), .RN(rstn), .Q(memory[730]) );
  DFFRHQX1 memory_reg_18__9_ ( .D(n1806), .CK(clk), .RN(rstn), .Q(memory[729])
         );
  DFFRHQX1 memory_reg_18__8_ ( .D(n1807), .CK(clk), .RN(rstn), .Q(memory[728])
         );
  DFFRHQX1 memory_reg_18__7_ ( .D(n1808), .CK(clk), .RN(rstn), .Q(memory[727])
         );
  DFFRHQX1 memory_reg_18__6_ ( .D(n1809), .CK(clk), .RN(rstn), .Q(memory[726])
         );
  DFFRHQX1 memory_reg_18__5_ ( .D(n1810), .CK(clk), .RN(rstn), .Q(memory[725])
         );
  DFFRHQX1 memory_reg_18__4_ ( .D(n1811), .CK(clk), .RN(rstn), .Q(memory[724])
         );
  DFFRHQX1 memory_reg_18__3_ ( .D(n1812), .CK(clk), .RN(rstn), .Q(memory[723])
         );
  DFFRHQX1 memory_reg_18__2_ ( .D(n1813), .CK(clk), .RN(rstn), .Q(memory[722])
         );
  DFFRHQX1 memory_reg_18__1_ ( .D(n1814), .CK(clk), .RN(rstn), .Q(memory[721])
         );
  DFFRHQX1 memory_reg_18__0_ ( .D(n1815), .CK(clk), .RN(rstn), .Q(memory[720])
         );
  DFFRHQX1 memory_reg_22__15_ ( .D(n1864), .CK(clk), .RN(rstn), .Q(memory[671]) );
  DFFRHQX1 memory_reg_22__14_ ( .D(n1865), .CK(clk), .RN(rstn), .Q(memory[670]) );
  DFFRHQX1 memory_reg_22__13_ ( .D(n1866), .CK(clk), .RN(rstn), .Q(memory[669]) );
  DFFRHQX1 memory_reg_22__12_ ( .D(n1867), .CK(clk), .RN(rstn), .Q(memory[668]) );
  DFFRHQX1 memory_reg_22__11_ ( .D(n1868), .CK(clk), .RN(rstn), .Q(memory[667]) );
  DFFRHQX1 memory_reg_22__10_ ( .D(n1869), .CK(clk), .RN(rstn), .Q(memory[666]) );
  DFFRHQX1 memory_reg_22__9_ ( .D(n1870), .CK(clk), .RN(rstn), .Q(memory[665])
         );
  DFFRHQX1 memory_reg_22__8_ ( .D(n1871), .CK(clk), .RN(rstn), .Q(memory[664])
         );
  DFFRHQX1 memory_reg_22__7_ ( .D(n1872), .CK(clk), .RN(rstn), .Q(memory[663])
         );
  DFFRHQX1 memory_reg_22__6_ ( .D(n1873), .CK(clk), .RN(rstn), .Q(memory[662])
         );
  DFFRHQX1 memory_reg_22__5_ ( .D(n1874), .CK(clk), .RN(rstn), .Q(memory[661])
         );
  DFFRHQX1 memory_reg_22__4_ ( .D(n1875), .CK(clk), .RN(rstn), .Q(memory[660])
         );
  DFFRHQX1 memory_reg_22__3_ ( .D(n1876), .CK(clk), .RN(rstn), .Q(memory[659])
         );
  DFFRHQX1 memory_reg_22__2_ ( .D(n1877), .CK(clk), .RN(rstn), .Q(memory[658])
         );
  DFFRHQX1 memory_reg_22__1_ ( .D(n1878), .CK(clk), .RN(rstn), .Q(memory[657])
         );
  DFFRHQX1 memory_reg_22__0_ ( .D(n1879), .CK(clk), .RN(rstn), .Q(memory[656])
         );
  DFFRHQX1 memory_reg_26__15_ ( .D(n1928), .CK(clk), .RN(rstn), .Q(memory[607]) );
  DFFRHQX1 memory_reg_26__14_ ( .D(n1929), .CK(clk), .RN(rstn), .Q(memory[606]) );
  DFFRHQX1 memory_reg_26__13_ ( .D(n1930), .CK(clk), .RN(rstn), .Q(memory[605]) );
  DFFRHQX1 memory_reg_26__12_ ( .D(n1931), .CK(clk), .RN(rstn), .Q(memory[604]) );
  DFFRHQX1 memory_reg_26__11_ ( .D(n1932), .CK(clk), .RN(rstn), .Q(memory[603]) );
  DFFRHQX1 memory_reg_26__10_ ( .D(n1933), .CK(clk), .RN(rstn), .Q(memory[602]) );
  DFFRHQX1 memory_reg_26__9_ ( .D(n1934), .CK(clk), .RN(rstn), .Q(memory[601])
         );
  DFFRHQX1 memory_reg_26__8_ ( .D(n1935), .CK(clk), .RN(rstn), .Q(memory[600])
         );
  DFFRHQX1 memory_reg_26__7_ ( .D(n1936), .CK(clk), .RN(rstn), .Q(memory[599])
         );
  DFFRHQX1 memory_reg_26__6_ ( .D(n1937), .CK(clk), .RN(rstn), .Q(memory[598])
         );
  DFFRHQX1 memory_reg_26__5_ ( .D(n1938), .CK(clk), .RN(rstn), .Q(memory[597])
         );
  DFFRHQX1 memory_reg_26__4_ ( .D(n1939), .CK(clk), .RN(rstn), .Q(memory[596])
         );
  DFFRHQX1 memory_reg_26__3_ ( .D(n1940), .CK(clk), .RN(rstn), .Q(memory[595])
         );
  DFFRHQX1 memory_reg_26__2_ ( .D(n1941), .CK(clk), .RN(rstn), .Q(memory[594])
         );
  DFFRHQX1 memory_reg_26__1_ ( .D(n1942), .CK(clk), .RN(rstn), .Q(memory[593])
         );
  DFFRHQX1 memory_reg_26__0_ ( .D(n1943), .CK(clk), .RN(rstn), .Q(memory[592])
         );
  DFFRHQX1 memory_reg_30__15_ ( .D(n1992), .CK(clk), .RN(rstn), .Q(memory[543]) );
  DFFRHQX1 memory_reg_30__14_ ( .D(n1993), .CK(clk), .RN(rstn), .Q(memory[542]) );
  DFFRHQX1 memory_reg_30__13_ ( .D(n1994), .CK(clk), .RN(rstn), .Q(memory[541]) );
  DFFRHQX1 memory_reg_30__12_ ( .D(n1995), .CK(clk), .RN(rstn), .Q(memory[540]) );
  DFFRHQX1 memory_reg_30__11_ ( .D(n1996), .CK(clk), .RN(rstn), .Q(memory[539]) );
  DFFRHQX1 memory_reg_30__10_ ( .D(n1997), .CK(clk), .RN(rstn), .Q(memory[538]) );
  DFFRHQX1 memory_reg_30__9_ ( .D(n1998), .CK(clk), .RN(rstn), .Q(memory[537])
         );
  DFFRHQX1 memory_reg_30__8_ ( .D(n1999), .CK(clk), .RN(rstn), .Q(memory[536])
         );
  DFFRHQX1 memory_reg_30__7_ ( .D(n2000), .CK(clk), .RN(rstn), .Q(memory[535])
         );
  DFFRHQX1 memory_reg_30__6_ ( .D(n2001), .CK(clk), .RN(rstn), .Q(memory[534])
         );
  DFFRHQX1 memory_reg_30__5_ ( .D(n2002), .CK(clk), .RN(rstn), .Q(memory[533])
         );
  DFFRHQX1 memory_reg_30__4_ ( .D(n2003), .CK(clk), .RN(rstn), .Q(memory[532])
         );
  DFFRHQX1 memory_reg_30__3_ ( .D(n2004), .CK(clk), .RN(rstn), .Q(memory[531])
         );
  DFFRHQX1 memory_reg_30__2_ ( .D(n2005), .CK(clk), .RN(rstn), .Q(memory[530])
         );
  DFFRHQX1 memory_reg_30__1_ ( .D(n2006), .CK(clk), .RN(rstn), .Q(memory[529])
         );
  DFFRHQX1 memory_reg_30__0_ ( .D(n2007), .CK(clk), .RN(rstn), .Q(memory[528])
         );
  DFFRHQX1 memory_reg_34__15_ ( .D(n2056), .CK(clk), .RN(rstn), .Q(memory[479]) );
  DFFRHQX1 memory_reg_34__14_ ( .D(n2057), .CK(clk), .RN(rstn), .Q(memory[478]) );
  DFFRHQX1 memory_reg_34__13_ ( .D(n2058), .CK(clk), .RN(rstn), .Q(memory[477]) );
  DFFRHQX1 memory_reg_34__12_ ( .D(n2059), .CK(clk), .RN(rstn), .Q(memory[476]) );
  DFFRHQX1 memory_reg_34__11_ ( .D(n2060), .CK(clk), .RN(rstn), .Q(memory[475]) );
  DFFRHQX1 memory_reg_34__10_ ( .D(n2061), .CK(clk), .RN(rstn), .Q(memory[474]) );
  DFFRHQX1 memory_reg_34__9_ ( .D(n2062), .CK(clk), .RN(rstn), .Q(memory[473])
         );
  DFFRHQX1 memory_reg_34__8_ ( .D(n2063), .CK(clk), .RN(rstn), .Q(memory[472])
         );
  DFFRHQX1 memory_reg_34__7_ ( .D(n2064), .CK(clk), .RN(rstn), .Q(memory[471])
         );
  DFFRHQX1 memory_reg_34__6_ ( .D(n2065), .CK(clk), .RN(rstn), .Q(memory[470])
         );
  DFFRHQX1 memory_reg_34__5_ ( .D(n2066), .CK(clk), .RN(rstn), .Q(memory[469])
         );
  DFFRHQX1 memory_reg_34__4_ ( .D(n2067), .CK(clk), .RN(rstn), .Q(memory[468])
         );
  DFFRHQX1 memory_reg_34__3_ ( .D(n2068), .CK(clk), .RN(rstn), .Q(memory[467])
         );
  DFFRHQX1 memory_reg_34__2_ ( .D(n2069), .CK(clk), .RN(rstn), .Q(memory[466])
         );
  DFFRHQX1 memory_reg_34__1_ ( .D(n2070), .CK(clk), .RN(rstn), .Q(memory[465])
         );
  DFFRHQX1 memory_reg_34__0_ ( .D(n2071), .CK(clk), .RN(rstn), .Q(memory[464])
         );
  DFFRHQX1 memory_reg_38__15_ ( .D(n2120), .CK(clk), .RN(rstn), .Q(memory[415]) );
  DFFRHQX1 memory_reg_38__14_ ( .D(n2121), .CK(clk), .RN(rstn), .Q(memory[414]) );
  DFFRHQX1 memory_reg_38__13_ ( .D(n2122), .CK(clk), .RN(rstn), .Q(memory[413]) );
  DFFRHQX1 memory_reg_38__12_ ( .D(n2123), .CK(clk), .RN(rstn), .Q(memory[412]) );
  DFFRHQX1 memory_reg_38__11_ ( .D(n2124), .CK(clk), .RN(rstn), .Q(memory[411]) );
  DFFRHQX1 memory_reg_38__10_ ( .D(n2125), .CK(clk), .RN(rstn), .Q(memory[410]) );
  DFFRHQX1 memory_reg_38__9_ ( .D(n2126), .CK(clk), .RN(rstn), .Q(memory[409])
         );
  DFFRHQX1 memory_reg_38__8_ ( .D(n2127), .CK(clk), .RN(rstn), .Q(memory[408])
         );
  DFFRHQX1 memory_reg_38__7_ ( .D(n2128), .CK(clk), .RN(rstn), .Q(memory[407])
         );
  DFFRHQX1 memory_reg_38__6_ ( .D(n2129), .CK(clk), .RN(rstn), .Q(memory[406])
         );
  DFFRHQX1 memory_reg_38__5_ ( .D(n2130), .CK(clk), .RN(rstn), .Q(memory[405])
         );
  DFFRHQX1 memory_reg_38__4_ ( .D(n2131), .CK(clk), .RN(rstn), .Q(memory[404])
         );
  DFFRHQX1 memory_reg_38__3_ ( .D(n2132), .CK(clk), .RN(rstn), .Q(memory[403])
         );
  DFFRHQX1 memory_reg_38__2_ ( .D(n2133), .CK(clk), .RN(rstn), .Q(memory[402])
         );
  DFFRHQX1 memory_reg_38__1_ ( .D(n2134), .CK(clk), .RN(rstn), .Q(memory[401])
         );
  DFFRHQX1 memory_reg_38__0_ ( .D(n2135), .CK(clk), .RN(rstn), .Q(memory[400])
         );
  DFFRHQX1 memory_reg_42__15_ ( .D(n2184), .CK(clk), .RN(rstn), .Q(memory[351]) );
  DFFRHQX1 memory_reg_42__14_ ( .D(n2185), .CK(clk), .RN(rstn), .Q(memory[350]) );
  DFFRHQX1 memory_reg_42__13_ ( .D(n2186), .CK(clk), .RN(rstn), .Q(memory[349]) );
  DFFRHQX1 memory_reg_42__12_ ( .D(n2187), .CK(clk), .RN(rstn), .Q(memory[348]) );
  DFFRHQX1 memory_reg_42__11_ ( .D(n2188), .CK(clk), .RN(rstn), .Q(memory[347]) );
  DFFRHQX1 memory_reg_42__10_ ( .D(n2189), .CK(clk), .RN(rstn), .Q(memory[346]) );
  DFFRHQX1 memory_reg_42__9_ ( .D(n2190), .CK(clk), .RN(rstn), .Q(memory[345])
         );
  DFFRHQX1 memory_reg_42__8_ ( .D(n2191), .CK(clk), .RN(rstn), .Q(memory[344])
         );
  DFFRHQX1 memory_reg_42__7_ ( .D(n2192), .CK(clk), .RN(rstn), .Q(memory[343])
         );
  DFFRHQX1 memory_reg_42__6_ ( .D(n2193), .CK(clk), .RN(rstn), .Q(memory[342])
         );
  DFFRHQX1 memory_reg_42__5_ ( .D(n2194), .CK(clk), .RN(rstn), .Q(memory[341])
         );
  DFFRHQX1 memory_reg_42__4_ ( .D(n2195), .CK(clk), .RN(rstn), .Q(memory[340])
         );
  DFFRHQX1 memory_reg_42__3_ ( .D(n2196), .CK(clk), .RN(rstn), .Q(memory[339])
         );
  DFFRHQX1 memory_reg_42__2_ ( .D(n2197), .CK(clk), .RN(rstn), .Q(memory[338])
         );
  DFFRHQX1 memory_reg_42__1_ ( .D(n2198), .CK(clk), .RN(rstn), .Q(memory[337])
         );
  DFFRHQX1 memory_reg_42__0_ ( .D(n2199), .CK(clk), .RN(rstn), .Q(memory[336])
         );
  DFFRHQX1 memory_reg_46__15_ ( .D(n2248), .CK(clk), .RN(rstn), .Q(memory[287]) );
  DFFRHQX1 memory_reg_46__14_ ( .D(n2249), .CK(clk), .RN(rstn), .Q(memory[286]) );
  DFFRHQX1 memory_reg_46__13_ ( .D(n2250), .CK(clk), .RN(rstn), .Q(memory[285]) );
  DFFRHQX1 memory_reg_46__12_ ( .D(n2251), .CK(clk), .RN(rstn), .Q(memory[284]) );
  DFFRHQX1 memory_reg_46__11_ ( .D(n2252), .CK(clk), .RN(rstn), .Q(memory[283]) );
  DFFRHQX1 memory_reg_46__10_ ( .D(n2253), .CK(clk), .RN(rstn), .Q(memory[282]) );
  DFFRHQX1 memory_reg_46__9_ ( .D(n2254), .CK(clk), .RN(rstn), .Q(memory[281])
         );
  DFFRHQX1 memory_reg_46__8_ ( .D(n2255), .CK(clk), .RN(rstn), .Q(memory[280])
         );
  DFFRHQX1 memory_reg_46__7_ ( .D(n2256), .CK(clk), .RN(rstn), .Q(memory[279])
         );
  DFFRHQX1 memory_reg_46__6_ ( .D(n2257), .CK(clk), .RN(rstn), .Q(memory[278])
         );
  DFFRHQX1 memory_reg_46__5_ ( .D(n2258), .CK(clk), .RN(rstn), .Q(memory[277])
         );
  DFFRHQX1 memory_reg_46__4_ ( .D(n2259), .CK(clk), .RN(rstn), .Q(memory[276])
         );
  DFFRHQX1 memory_reg_46__3_ ( .D(n2260), .CK(clk), .RN(rstn), .Q(memory[275])
         );
  DFFRHQX1 memory_reg_46__2_ ( .D(n2261), .CK(clk), .RN(rstn), .Q(memory[274])
         );
  DFFRHQX1 memory_reg_46__1_ ( .D(n2262), .CK(clk), .RN(rstn), .Q(memory[273])
         );
  DFFRHQX1 memory_reg_46__0_ ( .D(n2263), .CK(clk), .RN(rstn), .Q(memory[272])
         );
  DFFRHQX1 memory_reg_50__15_ ( .D(n2312), .CK(clk), .RN(rstn), .Q(memory[223]) );
  DFFRHQX1 memory_reg_50__14_ ( .D(n2313), .CK(clk), .RN(rstn), .Q(memory[222]) );
  DFFRHQX1 memory_reg_50__13_ ( .D(n2314), .CK(clk), .RN(rstn), .Q(memory[221]) );
  DFFRHQX1 memory_reg_50__12_ ( .D(n2315), .CK(clk), .RN(rstn), .Q(memory[220]) );
  DFFRHQX1 memory_reg_50__11_ ( .D(n2316), .CK(clk), .RN(rstn), .Q(memory[219]) );
  DFFRHQX1 memory_reg_50__10_ ( .D(n2317), .CK(clk), .RN(rstn), .Q(memory[218]) );
  DFFRHQX1 memory_reg_50__9_ ( .D(n2318), .CK(clk), .RN(rstn), .Q(memory[217])
         );
  DFFRHQX1 memory_reg_50__8_ ( .D(n2319), .CK(clk), .RN(rstn), .Q(memory[216])
         );
  DFFRHQX1 memory_reg_50__7_ ( .D(n2320), .CK(clk), .RN(rstn), .Q(memory[215])
         );
  DFFRHQX1 memory_reg_50__6_ ( .D(n2321), .CK(clk), .RN(rstn), .Q(memory[214])
         );
  DFFRHQX1 memory_reg_50__5_ ( .D(n2322), .CK(clk), .RN(rstn), .Q(memory[213])
         );
  DFFRHQX1 memory_reg_50__4_ ( .D(n2323), .CK(clk), .RN(rstn), .Q(memory[212])
         );
  DFFRHQX1 memory_reg_50__3_ ( .D(n2324), .CK(clk), .RN(rstn), .Q(memory[211])
         );
  DFFRHQX1 memory_reg_50__2_ ( .D(n2325), .CK(clk), .RN(rstn), .Q(memory[210])
         );
  DFFRHQX1 memory_reg_50__1_ ( .D(n2326), .CK(clk), .RN(rstn), .Q(memory[209])
         );
  DFFRHQX1 memory_reg_50__0_ ( .D(n2327), .CK(clk), .RN(rstn), .Q(memory[208])
         );
  DFFRHQX1 memory_reg_54__15_ ( .D(n2376), .CK(clk), .RN(rstn), .Q(memory[159]) );
  DFFRHQX1 memory_reg_54__14_ ( .D(n2377), .CK(clk), .RN(rstn), .Q(memory[158]) );
  DFFRHQX1 memory_reg_54__13_ ( .D(n2378), .CK(clk), .RN(rstn), .Q(memory[157]) );
  DFFRHQX1 memory_reg_54__12_ ( .D(n2379), .CK(clk), .RN(rstn), .Q(memory[156]) );
  DFFRHQX1 memory_reg_54__11_ ( .D(n2380), .CK(clk), .RN(rstn), .Q(memory[155]) );
  DFFRHQX1 memory_reg_54__10_ ( .D(n2381), .CK(clk), .RN(rstn), .Q(memory[154]) );
  DFFRHQX1 memory_reg_54__9_ ( .D(n2382), .CK(clk), .RN(rstn), .Q(memory[153])
         );
  DFFRHQX1 memory_reg_54__8_ ( .D(n2383), .CK(clk), .RN(rstn), .Q(memory[152])
         );
  DFFRHQX1 memory_reg_54__7_ ( .D(n2384), .CK(clk), .RN(rstn), .Q(memory[151])
         );
  DFFRHQX1 memory_reg_54__6_ ( .D(n2385), .CK(clk), .RN(rstn), .Q(memory[150])
         );
  DFFRHQX1 memory_reg_54__5_ ( .D(n2386), .CK(clk), .RN(rstn), .Q(memory[149])
         );
  DFFRHQX1 memory_reg_54__4_ ( .D(n2387), .CK(clk), .RN(rstn), .Q(memory[148])
         );
  DFFRHQX1 memory_reg_54__3_ ( .D(n2388), .CK(clk), .RN(rstn), .Q(memory[147])
         );
  DFFRHQX1 memory_reg_54__2_ ( .D(n2389), .CK(clk), .RN(rstn), .Q(memory[146])
         );
  DFFRHQX1 memory_reg_54__1_ ( .D(n2390), .CK(clk), .RN(rstn), .Q(memory[145])
         );
  DFFRHQX1 memory_reg_54__0_ ( .D(n2391), .CK(clk), .RN(rstn), .Q(memory[144])
         );
  DFFRHQX1 memory_reg_58__15_ ( .D(n2440), .CK(clk), .RN(rstn), .Q(memory[95])
         );
  DFFRHQX1 memory_reg_58__14_ ( .D(n2441), .CK(clk), .RN(rstn), .Q(memory[94])
         );
  DFFRHQX1 memory_reg_58__13_ ( .D(n2442), .CK(clk), .RN(rstn), .Q(memory[93])
         );
  DFFRHQX1 memory_reg_58__12_ ( .D(n2443), .CK(clk), .RN(rstn), .Q(memory[92])
         );
  DFFRHQX1 memory_reg_58__11_ ( .D(n2444), .CK(clk), .RN(rstn), .Q(memory[91])
         );
  DFFRHQX1 memory_reg_58__10_ ( .D(n2445), .CK(clk), .RN(rstn), .Q(memory[90])
         );
  DFFRHQX1 memory_reg_58__9_ ( .D(n2446), .CK(clk), .RN(rstn), .Q(memory[89])
         );
  DFFRHQX1 memory_reg_58__8_ ( .D(n2447), .CK(clk), .RN(rstn), .Q(memory[88])
         );
  DFFRHQX1 memory_reg_58__7_ ( .D(n2448), .CK(clk), .RN(rstn), .Q(memory[87])
         );
  DFFRHQX1 memory_reg_58__6_ ( .D(n2449), .CK(clk), .RN(rstn), .Q(memory[86])
         );
  DFFRHQX1 memory_reg_58__5_ ( .D(n2450), .CK(clk), .RN(rstn), .Q(memory[85])
         );
  DFFRHQX1 memory_reg_58__4_ ( .D(n2451), .CK(clk), .RN(rstn), .Q(memory[84])
         );
  DFFRHQX1 memory_reg_58__3_ ( .D(n2452), .CK(clk), .RN(rstn), .Q(memory[83])
         );
  DFFRHQX1 memory_reg_58__2_ ( .D(n2453), .CK(clk), .RN(rstn), .Q(memory[82])
         );
  DFFRHQX1 memory_reg_58__1_ ( .D(n2454), .CK(clk), .RN(rstn), .Q(memory[81])
         );
  DFFRHQX1 memory_reg_58__0_ ( .D(n2455), .CK(clk), .RN(rstn), .Q(memory[80])
         );
  DFFRHQX1 memory_reg_62__15_ ( .D(n2504), .CK(clk), .RN(rstn), .Q(memory[31])
         );
  DFFRHQX1 memory_reg_62__14_ ( .D(n2505), .CK(clk), .RN(rstn), .Q(memory[30])
         );
  DFFRHQX1 memory_reg_62__13_ ( .D(n2506), .CK(clk), .RN(rstn), .Q(memory[29])
         );
  DFFRHQX1 memory_reg_62__12_ ( .D(n2507), .CK(clk), .RN(rstn), .Q(memory[28])
         );
  DFFRHQX1 memory_reg_62__11_ ( .D(n2508), .CK(clk), .RN(rstn), .Q(memory[27])
         );
  DFFRHQX1 memory_reg_62__10_ ( .D(n2509), .CK(clk), .RN(rstn), .Q(memory[26])
         );
  DFFRHQX1 memory_reg_62__9_ ( .D(n2510), .CK(clk), .RN(rstn), .Q(memory[25])
         );
  DFFRHQX1 memory_reg_62__8_ ( .D(n2511), .CK(clk), .RN(rstn), .Q(memory[24])
         );
  DFFRHQX1 memory_reg_62__7_ ( .D(n2512), .CK(clk), .RN(rstn), .Q(memory[23])
         );
  DFFRHQX1 memory_reg_62__6_ ( .D(n2513), .CK(clk), .RN(rstn), .Q(memory[22])
         );
  DFFRHQX1 memory_reg_62__5_ ( .D(n2514), .CK(clk), .RN(rstn), .Q(memory[21])
         );
  DFFRHQX1 memory_reg_62__4_ ( .D(n2515), .CK(clk), .RN(rstn), .Q(memory[20])
         );
  DFFRHQX1 memory_reg_62__3_ ( .D(n2516), .CK(clk), .RN(rstn), .Q(memory[19])
         );
  DFFRHQX1 memory_reg_62__2_ ( .D(n2517), .CK(clk), .RN(rstn), .Q(memory[18])
         );
  DFFRHQX1 memory_reg_62__1_ ( .D(n2518), .CK(clk), .RN(rstn), .Q(memory[17])
         );
  DFFRHQX1 memory_reg_62__0_ ( .D(n2519), .CK(clk), .RN(rstn), .Q(memory[16])
         );
  INVXL U2 ( .A(addr[2]), .Y(n1508) );
  NAND2X1 U3 ( .A(n2553), .B(n2552), .Y(n1) );
  NAND2X1 U4 ( .A(n2551), .B(n2552), .Y(n2) );
  NAND2X1 U5 ( .A(n2545), .B(n2552), .Y(n3) );
  NAND2X1 U6 ( .A(n2543), .B(n2553), .Y(n4) );
  NAND2X1 U7 ( .A(n2543), .B(n2551), .Y(n5) );
  NAND2X1 U8 ( .A(n2543), .B(n2545), .Y(n6) );
  NAND2X1 U9 ( .A(n2542), .B(n2553), .Y(n7) );
  NAND2X1 U10 ( .A(n2542), .B(n2551), .Y(n8) );
  NAND2X1 U11 ( .A(n2542), .B(n2545), .Y(n9) );
  NAND2X1 U12 ( .A(n2541), .B(n2553), .Y(n10) );
  NAND2X1 U13 ( .A(n2541), .B(n2551), .Y(n11) );
  NAND2X1 U14 ( .A(n2541), .B(n2545), .Y(n12) );
  NAND2X1 U15 ( .A(n2540), .B(n2553), .Y(n13) );
  NAND2X1 U16 ( .A(n2540), .B(n2551), .Y(n14) );
  NAND2X1 U17 ( .A(n2540), .B(n2550), .Y(n15) );
  NAND2X1 U18 ( .A(n2540), .B(n2549), .Y(n16) );
  NAND2X1 U19 ( .A(n2540), .B(n2548), .Y(n17) );
  NAND2X1 U20 ( .A(n2540), .B(n2547), .Y(n18) );
  NAND2X1 U21 ( .A(n2540), .B(n2546), .Y(n19) );
  NAND2X1 U22 ( .A(n2540), .B(n2545), .Y(n20) );
  NAND2X1 U23 ( .A(n2539), .B(n2553), .Y(n21) );
  NAND2X1 U24 ( .A(n2539), .B(n2551), .Y(n22) );
  NAND2X1 U25 ( .A(n2539), .B(n2550), .Y(n25) );
  NAND2X1 U26 ( .A(n2539), .B(n2549), .Y(n27) );
  NAND2X1 U27 ( .A(n2539), .B(n2548), .Y(n29) );
  NAND2X1 U28 ( .A(n2539), .B(n2547), .Y(n31) );
  NAND2X1 U29 ( .A(n2539), .B(n2546), .Y(n33) );
  NAND2X1 U30 ( .A(n2539), .B(n2545), .Y(n35) );
  NAND2X1 U31 ( .A(n2538), .B(n2553), .Y(n37) );
  NAND2X1 U32 ( .A(n2538), .B(n2551), .Y(n40) );
  NAND2X1 U33 ( .A(n2538), .B(n2550), .Y(n42) );
  NAND2X1 U34 ( .A(n2538), .B(n2549), .Y(n43) );
  NAND2X1 U35 ( .A(n2538), .B(n2548), .Y(n44) );
  NAND2X1 U36 ( .A(n2538), .B(n2547), .Y(n45) );
  NAND2X1 U37 ( .A(n2538), .B(n2546), .Y(n46) );
  NAND2X1 U38 ( .A(n2538), .B(n2545), .Y(n47) );
  NAND2X1 U39 ( .A(n2537), .B(n2553), .Y(n48) );
  NAND2X1 U40 ( .A(n2537), .B(n2551), .Y(n49) );
  NAND2X1 U41 ( .A(n2537), .B(n2550), .Y(n51) );
  NAND2X1 U42 ( .A(n2537), .B(n2549), .Y(n52) );
  NAND2X1 U43 ( .A(n2537), .B(n2548), .Y(n53) );
  NAND2X1 U44 ( .A(n2537), .B(n2547), .Y(n54) );
  NAND2X1 U45 ( .A(n2537), .B(n2546), .Y(n55) );
  NAND2X1 U46 ( .A(n2537), .B(n2545), .Y(n56) );
  NAND2X1 U47 ( .A(n2550), .B(n2552), .Y(n57) );
  NAND2X1 U48 ( .A(n2549), .B(n2552), .Y(n58) );
  NAND2X1 U49 ( .A(n2548), .B(n2552), .Y(n60) );
  NAND2X1 U50 ( .A(n2547), .B(n2552), .Y(n61) );
  NAND2X1 U51 ( .A(n2546), .B(n2552), .Y(n62) );
  NAND2X1 U52 ( .A(n2543), .B(n2550), .Y(n63) );
  NAND2X1 U53 ( .A(n2543), .B(n2549), .Y(n64) );
  NAND2X1 U54 ( .A(n2543), .B(n2548), .Y(n65) );
  NAND2X1 U55 ( .A(n2543), .B(n2547), .Y(n66) );
  NAND2X1 U56 ( .A(n2543), .B(n2546), .Y(n67) );
  NAND2X1 U57 ( .A(n2542), .B(n2550), .Y(n69) );
  NAND2X1 U58 ( .A(n2542), .B(n2549), .Y(n70) );
  NAND2X1 U59 ( .A(n2542), .B(n2548), .Y(n71) );
  NAND2X1 U60 ( .A(n2542), .B(n2547), .Y(n72) );
  NAND2X1 U61 ( .A(n2542), .B(n2546), .Y(n73) );
  NAND2X1 U62 ( .A(n2541), .B(n2550), .Y(n74) );
  NAND2X1 U63 ( .A(n2541), .B(n2549), .Y(n75) );
  NAND2X1 U64 ( .A(n2541), .B(n2548), .Y(n76) );
  NAND2X1 U65 ( .A(n2541), .B(n2547), .Y(n78) );
  NAND2X1 U66 ( .A(n2541), .B(n2546), .Y(n79) );
  NOR4BX1 U67 ( .AN(n2544), .B(n1509), .C(addr[4]), .D(n1510), .Y(n2538) );
  NOR4BX1 U68 ( .AN(n2544), .B(addr[3]), .C(addr[4]), .D(n1510), .Y(n2537) );
  NOR4BX1 U69 ( .AN(n2544), .B(n1511), .C(n1509), .D(n1510), .Y(n2540) );
  NOR4BX1 U70 ( .AN(n2544), .B(n1511), .C(addr[3]), .D(n1510), .Y(n2539) );
  INVX1 U71 ( .A(n1506), .Y(n1454) );
  INVX1 U72 ( .A(n1506), .Y(n1455) );
  INVX1 U73 ( .A(n1506), .Y(n1456) );
  INVX1 U74 ( .A(n1506), .Y(n1457) );
  INVX1 U75 ( .A(n1506), .Y(n1458) );
  INVX1 U76 ( .A(n1506), .Y(n1459) );
  INVX1 U77 ( .A(n1506), .Y(n1460) );
  INVX1 U78 ( .A(n1506), .Y(n1461) );
  INVX1 U79 ( .A(n1453), .Y(n1462) );
  INVX1 U80 ( .A(n1453), .Y(n1463) );
  INVX1 U81 ( .A(n1453), .Y(n1464) );
  INVX1 U82 ( .A(n1453), .Y(n1465) );
  INVX1 U83 ( .A(n1453), .Y(n1466) );
  INVX1 U84 ( .A(n1453), .Y(n1467) );
  INVX1 U85 ( .A(n1506), .Y(n1468) );
  INVX1 U86 ( .A(n1506), .Y(n1469) );
  INVX1 U87 ( .A(n1506), .Y(n1470) );
  INVX1 U88 ( .A(n1433), .Y(n1434) );
  INVX1 U89 ( .A(n1433), .Y(n1435) );
  INVX1 U90 ( .A(n1507), .Y(n1436) );
  INVX1 U91 ( .A(n1433), .Y(n1437) );
  INVX1 U92 ( .A(n1433), .Y(n1438) );
  INVX1 U93 ( .A(n1507), .Y(n1439) );
  INVX1 U94 ( .A(n1507), .Y(n1440) );
  INVX1 U95 ( .A(n1433), .Y(n1441) );
  INVX1 U96 ( .A(n1433), .Y(n1442) );
  INVX1 U97 ( .A(n1433), .Y(n1443) );
  INVX1 U98 ( .A(n1507), .Y(n1444) );
  INVX1 U99 ( .A(n1433), .Y(n1445) );
  INVX1 U100 ( .A(n1433), .Y(n1446) );
  INVX1 U101 ( .A(n1433), .Y(n1447) );
  INVX1 U102 ( .A(n1433), .Y(n1448) );
  INVX1 U103 ( .A(n1433), .Y(n1449) );
  INVX1 U104 ( .A(n1507), .Y(n1450) );
  INVX1 U105 ( .A(n1507), .Y(n1451) );
  INVX1 U106 ( .A(n1471), .Y(n1453) );
  INVX1 U107 ( .A(addr[1]), .Y(n1433) );
  INVX1 U108 ( .A(n1507), .Y(n1452) );
  INVX1 U109 ( .A(n1509), .Y(n1427) );
  INVX1 U110 ( .A(n1509), .Y(n1428) );
  INVX1 U111 ( .A(n1509), .Y(n1429) );
  INVX1 U112 ( .A(n1509), .Y(n1430) );
  INVX1 U113 ( .A(n1506), .Y(n1471) );
  INVX1 U114 ( .A(n1508), .Y(n1431) );
  INVX1 U115 ( .A(n1508), .Y(n1432) );
  NOR3X1 U116 ( .A(n1507), .B(n1506), .C(n1508), .Y(n2553) );
  NOR3X1 U117 ( .A(n1507), .B(n1463), .C(n1508), .Y(n2551) );
  NOR3X1 U118 ( .A(n1506), .B(n1439), .C(n1508), .Y(n2550) );
  NOR3X1 U119 ( .A(n1467), .B(n1436), .C(n1508), .Y(n2549) );
  NOR3X1 U120 ( .A(n1506), .B(addr[2]), .C(n1507), .Y(n2548) );
  NOR3X1 U121 ( .A(n1464), .B(addr[2]), .C(n1507), .Y(n2547) );
  NOR3X1 U122 ( .A(n1440), .B(addr[2]), .C(n1506), .Y(n2546) );
  NOR3X1 U123 ( .A(n1452), .B(addr[2]), .C(n1462), .Y(n2545) );
  AND2X2 U124 ( .A(wr_rd), .B(en), .Y(n2544) );
  BUFX3 U125 ( .A(n2536), .Y(n1473) );
  NAND2BX1 U126 ( .AN(wr_rd), .B(en), .Y(n2536) );
  INVX1 U127 ( .A(din[0]), .Y(n1505) );
  INVX1 U128 ( .A(din[1]), .Y(n1503) );
  INVX1 U129 ( .A(din[2]), .Y(n1501) );
  INVX1 U130 ( .A(din[3]), .Y(n1499) );
  INVX1 U131 ( .A(din[4]), .Y(n1497) );
  INVX1 U132 ( .A(din[5]), .Y(n1495) );
  INVX1 U133 ( .A(din[6]), .Y(n1493) );
  INVX1 U134 ( .A(din[7]), .Y(n1491) );
  INVX1 U135 ( .A(din[8]), .Y(n1489) );
  INVX1 U136 ( .A(din[9]), .Y(n1487) );
  INVX1 U137 ( .A(din[10]), .Y(n1485) );
  INVX1 U138 ( .A(din[11]), .Y(n1483) );
  INVX1 U139 ( .A(din[12]), .Y(n1481) );
  INVX1 U140 ( .A(din[13]), .Y(n1479) );
  INVX1 U141 ( .A(din[14]), .Y(n1477) );
  INVX1 U142 ( .A(din[15]), .Y(n1475) );
  INVX1 U143 ( .A(din[0]), .Y(n1504) );
  INVX1 U144 ( .A(din[1]), .Y(n1502) );
  INVX1 U145 ( .A(din[2]), .Y(n1500) );
  INVX1 U146 ( .A(din[3]), .Y(n1498) );
  INVX1 U147 ( .A(din[4]), .Y(n1496) );
  INVX1 U148 ( .A(din[5]), .Y(n1494) );
  INVX1 U149 ( .A(din[6]), .Y(n1492) );
  INVX1 U150 ( .A(din[7]), .Y(n1490) );
  INVX1 U151 ( .A(din[8]), .Y(n1488) );
  INVX1 U152 ( .A(din[9]), .Y(n1486) );
  INVX1 U153 ( .A(din[10]), .Y(n1484) );
  INVX1 U154 ( .A(din[11]), .Y(n1482) );
  INVX1 U155 ( .A(din[12]), .Y(n1480) );
  INVX1 U156 ( .A(din[13]), .Y(n1478) );
  INVX1 U157 ( .A(din[14]), .Y(n1476) );
  INVX1 U158 ( .A(din[15]), .Y(n1474) );
  NOR2BX1 U159 ( .AN(N100), .B(n1473), .Y(dout[0]) );
  MX4X1 U160 ( .A(n101), .B(n90), .C(n96), .D(n84), .S0(n1510), .S1(n1472), 
        .Y(N100) );
  MX4X1 U161 ( .A(n83), .B(n81), .C(n82), .D(n80), .S0(n1427), .S1(n1431), .Y(
        n84) );
  MX4X1 U162 ( .A(n100), .B(n98), .C(n99), .D(n97), .S0(n1430), .S1(n1432), 
        .Y(n101) );
  NOR2BX1 U163 ( .AN(N99), .B(n1473), .Y(dout[1]) );
  MX4X1 U164 ( .A(n1146), .B(n1136), .C(n1141), .D(n1131), .S0(n1510), .S1(
        n1472), .Y(N99) );
  MX4X1 U165 ( .A(n1145), .B(n1143), .C(n1144), .D(n1142), .S0(n1427), .S1(
        n1431), .Y(n1146) );
  MX4X1 U166 ( .A(n1135), .B(n1133), .C(n1134), .D(n1132), .S0(n1427), .S1(
        n1431), .Y(n1136) );
  NOR2BX1 U167 ( .AN(N98), .B(n1473), .Y(dout[2]) );
  MX4X1 U168 ( .A(n1166), .B(n1156), .C(n1161), .D(n1151), .S0(n1510), .S1(
        n1472), .Y(N98) );
  MX4X1 U169 ( .A(n1165), .B(n1163), .C(n1164), .D(n1162), .S0(n1427), .S1(
        n1431), .Y(n1166) );
  MX4X1 U170 ( .A(n1155), .B(n1153), .C(n1154), .D(n1152), .S0(n1427), .S1(
        n1431), .Y(n1156) );
  NOR2BX1 U171 ( .AN(N97), .B(n1473), .Y(dout[3]) );
  MX4X1 U172 ( .A(n1186), .B(n1176), .C(n1181), .D(n1171), .S0(n1510), .S1(
        n1472), .Y(N97) );
  MX4X1 U173 ( .A(n1185), .B(n1183), .C(n1184), .D(n1182), .S0(n1427), .S1(
        n1431), .Y(n1186) );
  MX4X1 U174 ( .A(n1175), .B(n1173), .C(n1174), .D(n1172), .S0(n1427), .S1(
        n1431), .Y(n1176) );
  NOR2BX1 U175 ( .AN(N96), .B(n1473), .Y(dout[4]) );
  MX4X1 U176 ( .A(n1206), .B(n1196), .C(n1201), .D(n1191), .S0(addr[5]), .S1(
        n1472), .Y(N96) );
  MX4X1 U177 ( .A(n1205), .B(n1203), .C(n1204), .D(n1202), .S0(n1428), .S1(
        n1432), .Y(n1206) );
  MX4X1 U178 ( .A(n1195), .B(n1193), .C(n1194), .D(n1192), .S0(n1428), .S1(
        n1432), .Y(n1196) );
  NOR2BX1 U179 ( .AN(N95), .B(n1473), .Y(dout[5]) );
  MX4X1 U180 ( .A(n1226), .B(n1216), .C(n1221), .D(n1211), .S0(n1510), .S1(
        n1472), .Y(N95) );
  MX4X1 U181 ( .A(n1225), .B(n1223), .C(n1224), .D(n1222), .S0(n1428), .S1(
        n1432), .Y(n1226) );
  MX4X1 U182 ( .A(n1215), .B(n1213), .C(n1214), .D(n1212), .S0(n1428), .S1(
        n1432), .Y(n1216) );
  NOR2BX1 U183 ( .AN(N94), .B(n1473), .Y(dout[6]) );
  MX4X1 U184 ( .A(n1246), .B(n1236), .C(n1241), .D(n1231), .S0(n1510), .S1(
        n1472), .Y(N94) );
  MX4X1 U185 ( .A(n1245), .B(n1243), .C(n1244), .D(n1242), .S0(n1428), .S1(
        n1432), .Y(n1246) );
  MX4X1 U186 ( .A(n1235), .B(n1233), .C(n1234), .D(n1232), .S0(n1428), .S1(
        n1432), .Y(n1236) );
  NOR2BX1 U187 ( .AN(N93), .B(n1473), .Y(dout[7]) );
  MX4X1 U188 ( .A(n1266), .B(n1256), .C(n1261), .D(n1251), .S0(n1510), .S1(
        n1472), .Y(N93) );
  MX4X1 U189 ( .A(n1265), .B(n1263), .C(n1264), .D(n1262), .S0(n1429), .S1(
        n1431), .Y(n1266) );
  MX4X1 U190 ( .A(n1255), .B(n1253), .C(n1254), .D(n1252), .S0(n1429), .S1(
        n1431), .Y(n1256) );
  NOR2BX1 U191 ( .AN(N92), .B(n1473), .Y(dout[8]) );
  MX4X1 U192 ( .A(n1286), .B(n1276), .C(n1281), .D(n1271), .S0(n1510), .S1(
        n1472), .Y(N92) );
  MX4X1 U193 ( .A(n1285), .B(n1283), .C(n1284), .D(n1282), .S0(n1429), .S1(
        n1432), .Y(n1286) );
  MX4X1 U194 ( .A(n1275), .B(n1273), .C(n1274), .D(n1272), .S0(n1429), .S1(
        n1432), .Y(n1276) );
  NOR2BX1 U195 ( .AN(N91), .B(n1473), .Y(dout[9]) );
  MX4X1 U196 ( .A(n1306), .B(n1296), .C(n1301), .D(n1291), .S0(addr[5]), .S1(
        n1472), .Y(N91) );
  MX4X1 U197 ( .A(n1305), .B(n1303), .C(n1304), .D(n1302), .S0(n1429), .S1(
        n1432), .Y(n1306) );
  MX4X1 U198 ( .A(n1295), .B(n1293), .C(n1294), .D(n1292), .S0(n1429), .S1(
        n1431), .Y(n1296) );
  NOR2BX1 U199 ( .AN(N90), .B(n1473), .Y(dout[10]) );
  MX4X1 U200 ( .A(n1326), .B(n1316), .C(n1321), .D(n1311), .S0(addr[5]), .S1(
        n1472), .Y(N90) );
  MX4X1 U201 ( .A(n1325), .B(n1323), .C(n1324), .D(n1322), .S0(n1430), .S1(
        addr[2]), .Y(n1326) );
  MX4X1 U202 ( .A(n1315), .B(n1313), .C(n1314), .D(n1312), .S0(n1430), .S1(
        addr[2]), .Y(n1316) );
  NOR2BX1 U203 ( .AN(N89), .B(n1473), .Y(dout[11]) );
  MX4X1 U204 ( .A(n1346), .B(n1336), .C(n1341), .D(n1331), .S0(addr[5]), .S1(
        n1472), .Y(N89) );
  MX4X1 U205 ( .A(n1345), .B(n1343), .C(n1344), .D(n1342), .S0(n1430), .S1(
        addr[2]), .Y(n1346) );
  MX4X1 U206 ( .A(n1335), .B(n1333), .C(n1334), .D(n1332), .S0(n1430), .S1(
        addr[2]), .Y(n1336) );
  NOR2BX1 U207 ( .AN(N88), .B(n1473), .Y(dout[12]) );
  MX4X1 U208 ( .A(n1366), .B(n1356), .C(n1361), .D(n1351), .S0(addr[5]), .S1(
        n1472), .Y(N88) );
  MX4X1 U209 ( .A(n1365), .B(n1363), .C(n1364), .D(n1362), .S0(n1430), .S1(
        addr[2]), .Y(n1366) );
  MX4X1 U210 ( .A(n1355), .B(n1353), .C(n1354), .D(n1352), .S0(n1430), .S1(
        addr[2]), .Y(n1356) );
  NOR2BX1 U211 ( .AN(N87), .B(n1473), .Y(dout[13]) );
  MX4X1 U212 ( .A(n1386), .B(n1376), .C(n1381), .D(n1371), .S0(addr[5]), .S1(
        n1472), .Y(N87) );
  MX4X1 U213 ( .A(n1385), .B(n1383), .C(n1384), .D(n1382), .S0(addr[3]), .S1(
        addr[2]), .Y(n1386) );
  MX4X1 U214 ( .A(n1375), .B(n1373), .C(n1374), .D(n1372), .S0(addr[3]), .S1(
        n1431), .Y(n1376) );
  NOR2BX1 U215 ( .AN(N86), .B(n1473), .Y(dout[14]) );
  MX4X1 U216 ( .A(n1406), .B(n1396), .C(n1401), .D(n1391), .S0(addr[5]), .S1(
        n1472), .Y(N86) );
  MX4X1 U217 ( .A(n1405), .B(n1403), .C(n1404), .D(n1402), .S0(addr[3]), .S1(
        addr[2]), .Y(n1406) );
  MX4X1 U218 ( .A(n1395), .B(n1393), .C(n1394), .D(n1392), .S0(addr[3]), .S1(
        n1432), .Y(n1396) );
  NOR2BX1 U219 ( .AN(N85), .B(n1473), .Y(dout[15]) );
  MX4X1 U220 ( .A(n1426), .B(n1416), .C(n1421), .D(n1411), .S0(addr[5]), .S1(
        n1472), .Y(N85) );
  MX4X1 U221 ( .A(n1425), .B(n1423), .C(n1424), .D(n1422), .S0(addr[3]), .S1(
        addr[2]), .Y(n1426) );
  MX4X1 U222 ( .A(n1415), .B(n1413), .C(n1414), .D(n1412), .S0(addr[3]), .S1(
        addr[2]), .Y(n1416) );
  INVX1 U223 ( .A(addr[0]), .Y(n1506) );
  INVX1 U224 ( .A(addr[1]), .Y(n1507) );
  INVX1 U225 ( .A(addr[3]), .Y(n1509) );
  AND4X2 U226 ( .A(n2544), .B(n1510), .C(addr[4]), .D(n1509), .Y(n2543) );
  AND4X2 U227 ( .A(n2544), .B(n1510), .C(addr[4]), .D(n1427), .Y(n2552) );
  AND4X2 U228 ( .A(n2544), .B(n1510), .C(addr[3]), .D(n1511), .Y(n2542) );
  AND4X2 U229 ( .A(n2544), .B(n1510), .C(n1509), .D(n1511), .Y(n2541) );
  INVX1 U230 ( .A(addr[4]), .Y(n1511) );
  BUFX3 U231 ( .A(addr[4]), .Y(n1472) );
  MX4X1 U232 ( .A(memory[944]), .B(memory[928]), .C(memory[912]), .D(
        memory[896]), .S0(n1454), .S1(n1450), .Y(n99) );
  MX4X1 U233 ( .A(memory[176]), .B(memory[160]), .C(memory[144]), .D(
        memory[128]), .S0(n1454), .S1(n1451), .Y(n82) );
  MX4X1 U234 ( .A(memory[433]), .B(memory[417]), .C(memory[401]), .D(
        memory[385]), .S0(n1455), .S1(n1434), .Y(n1134) );
  MX4X1 U235 ( .A(memory[945]), .B(memory[929]), .C(memory[913]), .D(
        memory[897]), .S0(n1456), .S1(n1435), .Y(n1144) );
  MX4X1 U236 ( .A(memory[434]), .B(memory[418]), .C(memory[402]), .D(
        memory[386]), .S0(n1456), .S1(n1435), .Y(n1154) );
  MX4X1 U237 ( .A(memory[946]), .B(memory[930]), .C(memory[914]), .D(
        memory[898]), .S0(n1457), .S1(n1436), .Y(n1164) );
  MX4X1 U238 ( .A(memory[435]), .B(memory[419]), .C(memory[403]), .D(
        memory[387]), .S0(n1458), .S1(n1437), .Y(n1174) );
  MX4X1 U239 ( .A(memory[947]), .B(memory[931]), .C(memory[915]), .D(
        memory[899]), .S0(n1458), .S1(n1437), .Y(n1184) );
  MX4X1 U240 ( .A(memory[436]), .B(memory[420]), .C(memory[404]), .D(
        memory[388]), .S0(n1459), .S1(n1438), .Y(n1194) );
  MX4X1 U241 ( .A(memory[948]), .B(memory[932]), .C(memory[916]), .D(
        memory[900]), .S0(n1460), .S1(n1439), .Y(n1204) );
  MX4X1 U242 ( .A(memory[437]), .B(memory[421]), .C(memory[405]), .D(
        memory[389]), .S0(n1460), .S1(n1439), .Y(n1214) );
  MX4X1 U243 ( .A(memory[949]), .B(memory[933]), .C(memory[917]), .D(
        memory[901]), .S0(n1461), .S1(n1440), .Y(n1224) );
  MX4X1 U244 ( .A(memory[438]), .B(memory[422]), .C(memory[406]), .D(
        memory[390]), .S0(n1462), .S1(n1441), .Y(n1234) );
  MX4X1 U245 ( .A(memory[950]), .B(memory[934]), .C(memory[918]), .D(
        memory[902]), .S0(n1462), .S1(n1441), .Y(n1244) );
  MX4X1 U246 ( .A(memory[439]), .B(memory[423]), .C(memory[407]), .D(
        memory[391]), .S0(n1463), .S1(n1442), .Y(n1254) );
  MX4X1 U247 ( .A(memory[951]), .B(memory[935]), .C(memory[919]), .D(
        memory[903]), .S0(n1464), .S1(n1443), .Y(n1264) );
  MX4X1 U248 ( .A(memory[440]), .B(memory[424]), .C(memory[408]), .D(
        memory[392]), .S0(n1464), .S1(n1443), .Y(n1274) );
  MX4X1 U249 ( .A(memory[952]), .B(memory[936]), .C(memory[920]), .D(
        memory[904]), .S0(n1469), .S1(n1444), .Y(n1284) );
  MX4X1 U250 ( .A(memory[441]), .B(memory[425]), .C(memory[409]), .D(
        memory[393]), .S0(n1469), .S1(n1445), .Y(n1294) );
  MX4X1 U251 ( .A(memory[953]), .B(memory[937]), .C(memory[921]), .D(
        memory[905]), .S0(n1456), .S1(n1445), .Y(n1304) );
  MX4X1 U252 ( .A(memory[442]), .B(memory[426]), .C(memory[410]), .D(
        memory[394]), .S0(n1465), .S1(n1446), .Y(n1314) );
  MX4X1 U253 ( .A(memory[954]), .B(memory[938]), .C(memory[922]), .D(
        memory[906]), .S0(n1466), .S1(n1447), .Y(n1324) );
  MX4X1 U254 ( .A(memory[443]), .B(memory[427]), .C(memory[411]), .D(
        memory[395]), .S0(n1466), .S1(n1447), .Y(n1334) );
  MX4X1 U255 ( .A(memory[955]), .B(memory[939]), .C(memory[923]), .D(
        memory[907]), .S0(n1467), .S1(n1448), .Y(n1344) );
  MX4X1 U256 ( .A(memory[444]), .B(memory[428]), .C(memory[412]), .D(
        memory[396]), .S0(n1467), .S1(n1449), .Y(n1354) );
  MX4X1 U257 ( .A(memory[956]), .B(memory[940]), .C(memory[924]), .D(
        memory[908]), .S0(n1466), .S1(n1449), .Y(n1364) );
  MX4X1 U258 ( .A(memory[445]), .B(memory[429]), .C(memory[413]), .D(
        memory[397]), .S0(n1468), .S1(n1450), .Y(n1374) );
  MX4X1 U259 ( .A(memory[957]), .B(memory[941]), .C(memory[925]), .D(
        memory[909]), .S0(n1469), .S1(n1450), .Y(n1384) );
  MX4X1 U260 ( .A(memory[446]), .B(memory[430]), .C(memory[414]), .D(
        memory[398]), .S0(n1469), .S1(n1451), .Y(n1394) );
  MX4X1 U261 ( .A(memory[958]), .B(memory[942]), .C(memory[926]), .D(
        memory[910]), .S0(n1470), .S1(n1451), .Y(n1404) );
  MX4X1 U262 ( .A(memory[447]), .B(memory[431]), .C(memory[415]), .D(
        memory[399]), .S0(n1460), .S1(n1452), .Y(n1414) );
  MX4X1 U263 ( .A(memory[959]), .B(memory[943]), .C(memory[927]), .D(
        memory[911]), .S0(n1458), .S1(n1452), .Y(n1424) );
  MX4X1 U264 ( .A(n94), .B(n92), .C(n93), .D(n91), .S0(n1428), .S1(n1432), .Y(
        n96) );
  MX4X1 U265 ( .A(memory[752]), .B(memory[736]), .C(memory[720]), .D(
        memory[704]), .S0(n1454), .S1(addr[1]), .Y(n94) );
  MX4X1 U266 ( .A(memory[624]), .B(memory[608]), .C(memory[592]), .D(
        memory[576]), .S0(n1454), .S1(addr[1]), .Y(n92) );
  MX4X1 U267 ( .A(memory[688]), .B(memory[672]), .C(memory[656]), .D(
        memory[640]), .S0(n1454), .S1(n1451), .Y(n93) );
  MX4X1 U268 ( .A(n1140), .B(n1138), .C(n1139), .D(n1137), .S0(n1427), .S1(
        n1431), .Y(n1141) );
  MX4X1 U269 ( .A(memory[753]), .B(memory[737]), .C(memory[721]), .D(
        memory[705]), .S0(n1455), .S1(n1434), .Y(n1140) );
  MX4X1 U270 ( .A(memory[625]), .B(memory[609]), .C(memory[593]), .D(
        memory[577]), .S0(n1455), .S1(n1434), .Y(n1138) );
  MX4X1 U271 ( .A(memory[689]), .B(memory[673]), .C(memory[657]), .D(
        memory[641]), .S0(n1455), .S1(n1434), .Y(n1139) );
  MX4X1 U272 ( .A(n1160), .B(n1158), .C(n1159), .D(n1157), .S0(n1427), .S1(
        n1431), .Y(n1161) );
  MX4X1 U273 ( .A(memory[754]), .B(memory[738]), .C(memory[722]), .D(
        memory[706]), .S0(n1457), .S1(n1436), .Y(n1160) );
  MX4X1 U274 ( .A(memory[626]), .B(memory[610]), .C(memory[594]), .D(
        memory[578]), .S0(n1457), .S1(n1436), .Y(n1158) );
  MX4X1 U275 ( .A(memory[690]), .B(memory[674]), .C(memory[658]), .D(
        memory[642]), .S0(n1457), .S1(n1436), .Y(n1159) );
  MX4X1 U276 ( .A(n1180), .B(n1178), .C(n1179), .D(n1177), .S0(n1427), .S1(
        n1431), .Y(n1181) );
  MX4X1 U277 ( .A(memory[755]), .B(memory[739]), .C(memory[723]), .D(
        memory[707]), .S0(n1458), .S1(n1437), .Y(n1180) );
  MX4X1 U278 ( .A(memory[627]), .B(memory[611]), .C(memory[595]), .D(
        memory[579]), .S0(n1458), .S1(n1437), .Y(n1178) );
  MX4X1 U279 ( .A(memory[691]), .B(memory[675]), .C(memory[659]), .D(
        memory[643]), .S0(n1458), .S1(n1437), .Y(n1179) );
  MX4X1 U280 ( .A(n1200), .B(n1198), .C(n1199), .D(n1197), .S0(n1428), .S1(
        n1432), .Y(n1201) );
  MX4X1 U281 ( .A(memory[756]), .B(memory[740]), .C(memory[724]), .D(
        memory[708]), .S0(n1459), .S1(n1438), .Y(n1200) );
  MX4X1 U282 ( .A(memory[628]), .B(memory[612]), .C(memory[596]), .D(
        memory[580]), .S0(n1459), .S1(n1438), .Y(n1198) );
  MX4X1 U283 ( .A(memory[692]), .B(memory[676]), .C(memory[660]), .D(
        memory[644]), .S0(n1459), .S1(n1438), .Y(n1199) );
  MX4X1 U284 ( .A(n1220), .B(n1218), .C(n1219), .D(n1217), .S0(n1428), .S1(
        n1432), .Y(n1221) );
  MX4X1 U285 ( .A(memory[757]), .B(memory[741]), .C(memory[725]), .D(
        memory[709]), .S0(n1461), .S1(n1440), .Y(n1220) );
  MX4X1 U286 ( .A(memory[629]), .B(memory[613]), .C(memory[597]), .D(
        memory[581]), .S0(n1461), .S1(n1440), .Y(n1218) );
  MX4X1 U287 ( .A(memory[693]), .B(memory[677]), .C(memory[661]), .D(
        memory[645]), .S0(n1461), .S1(n1440), .Y(n1219) );
  MX4X1 U288 ( .A(n1240), .B(n1238), .C(n1239), .D(n1237), .S0(n1428), .S1(
        n1432), .Y(n1241) );
  MX4X1 U289 ( .A(memory[758]), .B(memory[742]), .C(memory[726]), .D(
        memory[710]), .S0(n1462), .S1(n1441), .Y(n1240) );
  MX4X1 U290 ( .A(memory[630]), .B(memory[614]), .C(memory[598]), .D(
        memory[582]), .S0(n1462), .S1(n1441), .Y(n1238) );
  MX4X1 U291 ( .A(memory[694]), .B(memory[678]), .C(memory[662]), .D(
        memory[646]), .S0(n1462), .S1(n1441), .Y(n1239) );
  MX4X1 U292 ( .A(n1260), .B(n1258), .C(n1259), .D(n1257), .S0(n1429), .S1(
        n1431), .Y(n1261) );
  MX4X1 U293 ( .A(memory[759]), .B(memory[743]), .C(memory[727]), .D(
        memory[711]), .S0(n1463), .S1(n1442), .Y(n1260) );
  MX4X1 U294 ( .A(memory[631]), .B(memory[615]), .C(memory[599]), .D(
        memory[583]), .S0(n1463), .S1(n1442), .Y(n1258) );
  MX4X1 U295 ( .A(memory[695]), .B(memory[679]), .C(memory[663]), .D(
        memory[647]), .S0(n1463), .S1(n1442), .Y(n1259) );
  MX4X1 U296 ( .A(n1280), .B(n1278), .C(n1279), .D(n1277), .S0(n1429), .S1(
        n1432), .Y(n1281) );
  MX4X1 U297 ( .A(memory[760]), .B(memory[744]), .C(memory[728]), .D(
        memory[712]), .S0(n1468), .S1(n1444), .Y(n1280) );
  MX4X1 U298 ( .A(memory[632]), .B(memory[616]), .C(memory[600]), .D(
        memory[584]), .S0(n1459), .S1(n1444), .Y(n1278) );
  MX4X1 U299 ( .A(memory[696]), .B(memory[680]), .C(memory[664]), .D(
        memory[648]), .S0(n1460), .S1(n1444), .Y(n1279) );
  MX4X1 U300 ( .A(n1300), .B(n1298), .C(n1299), .D(n1297), .S0(n1429), .S1(
        n1432), .Y(n1301) );
  MX4X1 U301 ( .A(memory[761]), .B(memory[745]), .C(memory[729]), .D(
        memory[713]), .S0(n1458), .S1(n1445), .Y(n1300) );
  MX4X1 U302 ( .A(memory[633]), .B(memory[617]), .C(memory[601]), .D(
        memory[585]), .S0(n1468), .S1(n1445), .Y(n1298) );
  MX4X1 U303 ( .A(memory[697]), .B(memory[681]), .C(memory[665]), .D(
        memory[649]), .S0(n1464), .S1(n1445), .Y(n1299) );
  MX4X1 U304 ( .A(n1320), .B(n1318), .C(n1319), .D(n1317), .S0(n1430), .S1(
        addr[2]), .Y(n1321) );
  MX4X1 U305 ( .A(memory[762]), .B(memory[746]), .C(memory[730]), .D(
        memory[714]), .S0(n1465), .S1(n1446), .Y(n1320) );
  MX4X1 U306 ( .A(memory[634]), .B(memory[618]), .C(memory[602]), .D(
        memory[586]), .S0(n1465), .S1(n1446), .Y(n1318) );
  MX4X1 U307 ( .A(memory[698]), .B(memory[682]), .C(memory[666]), .D(
        memory[650]), .S0(n1465), .S1(n1446), .Y(n1319) );
  MX4X1 U308 ( .A(n1340), .B(n1338), .C(n1339), .D(n1337), .S0(n1430), .S1(
        addr[2]), .Y(n1341) );
  MX4X1 U309 ( .A(memory[763]), .B(memory[747]), .C(memory[731]), .D(
        memory[715]), .S0(n1467), .S1(n1448), .Y(n1340) );
  MX4X1 U310 ( .A(memory[635]), .B(memory[619]), .C(memory[603]), .D(
        memory[587]), .S0(n1467), .S1(n1448), .Y(n1338) );
  MX4X1 U311 ( .A(memory[699]), .B(memory[683]), .C(memory[667]), .D(
        memory[651]), .S0(n1467), .S1(n1448), .Y(n1339) );
  MX4X1 U312 ( .A(n1360), .B(n1358), .C(n1359), .D(n1357), .S0(n1430), .S1(
        addr[2]), .Y(n1361) );
  MX4X1 U313 ( .A(memory[764]), .B(memory[748]), .C(memory[732]), .D(
        memory[716]), .S0(n1465), .S1(n1449), .Y(n1360) );
  MX4X1 U314 ( .A(memory[636]), .B(memory[620]), .C(memory[604]), .D(
        memory[588]), .S0(n1469), .S1(n1449), .Y(n1358) );
  MX4X1 U315 ( .A(memory[700]), .B(memory[684]), .C(memory[668]), .D(
        memory[652]), .S0(n1459), .S1(n1449), .Y(n1359) );
  MX4X1 U316 ( .A(n1380), .B(n1378), .C(n1379), .D(n1377), .S0(n1427), .S1(
        addr[2]), .Y(n1381) );
  MX4X1 U317 ( .A(memory[765]), .B(memory[749]), .C(memory[733]), .D(
        memory[717]), .S0(n1468), .S1(n1450), .Y(n1380) );
  MX4X1 U318 ( .A(memory[637]), .B(memory[621]), .C(memory[605]), .D(
        memory[589]), .S0(n1468), .S1(n1450), .Y(n1378) );
  MX4X1 U319 ( .A(memory[701]), .B(memory[685]), .C(memory[669]), .D(
        memory[653]), .S0(n1468), .S1(n1450), .Y(n1379) );
  MX4X1 U320 ( .A(n1400), .B(n1398), .C(n1399), .D(n1397), .S0(addr[3]), .S1(
        addr[2]), .Y(n1401) );
  MX4X1 U321 ( .A(memory[766]), .B(memory[750]), .C(memory[734]), .D(
        memory[718]), .S0(n1470), .S1(n1451), .Y(n1400) );
  MX4X1 U322 ( .A(memory[638]), .B(memory[622]), .C(memory[606]), .D(
        memory[590]), .S0(n1470), .S1(n1451), .Y(n1398) );
  MX4X1 U323 ( .A(memory[702]), .B(memory[686]), .C(memory[670]), .D(
        memory[654]), .S0(n1470), .S1(n1451), .Y(n1399) );
  MX4X1 U324 ( .A(n1420), .B(n1418), .C(n1419), .D(n1417), .S0(addr[3]), .S1(
        n1431), .Y(n1421) );
  MX4X1 U325 ( .A(memory[767]), .B(memory[751]), .C(memory[735]), .D(
        memory[719]), .S0(n1461), .S1(n1452), .Y(n1420) );
  MX4X1 U326 ( .A(memory[639]), .B(memory[623]), .C(memory[607]), .D(
        memory[591]), .S0(n1457), .S1(n1452), .Y(n1418) );
  MX4X1 U327 ( .A(memory[703]), .B(memory[687]), .C(memory[671]), .D(
        memory[655]), .S0(n1471), .S1(n1452), .Y(n1419) );
  MX4X1 U328 ( .A(memory[1008]), .B(memory[992]), .C(memory[976]), .D(
        memory[960]), .S0(n1454), .S1(n1451), .Y(n100) );
  MX4X1 U329 ( .A(memory[240]), .B(memory[224]), .C(memory[208]), .D(
        memory[192]), .S0(n1469), .S1(addr[1]), .Y(n83) );
  MX4X1 U330 ( .A(memory[497]), .B(memory[481]), .C(memory[465]), .D(
        memory[449]), .S0(n1455), .S1(n1434), .Y(n1135) );
  MX4X1 U331 ( .A(memory[1009]), .B(memory[993]), .C(memory[977]), .D(
        memory[961]), .S0(n1456), .S1(n1435), .Y(n1145) );
  MX4X1 U332 ( .A(memory[498]), .B(memory[482]), .C(memory[466]), .D(
        memory[450]), .S0(n1456), .S1(n1435), .Y(n1155) );
  MX4X1 U333 ( .A(memory[1010]), .B(memory[994]), .C(memory[978]), .D(
        memory[962]), .S0(n1457), .S1(n1436), .Y(n1165) );
  MX4X1 U334 ( .A(memory[499]), .B(memory[483]), .C(memory[467]), .D(
        memory[451]), .S0(n1458), .S1(n1437), .Y(n1175) );
  MX4X1 U335 ( .A(memory[1011]), .B(memory[995]), .C(memory[979]), .D(
        memory[963]), .S0(n1458), .S1(n1437), .Y(n1185) );
  MX4X1 U336 ( .A(memory[500]), .B(memory[484]), .C(memory[468]), .D(
        memory[452]), .S0(n1459), .S1(n1438), .Y(n1195) );
  MX4X1 U337 ( .A(memory[1012]), .B(memory[996]), .C(memory[980]), .D(
        memory[964]), .S0(n1460), .S1(n1439), .Y(n1205) );
  MX4X1 U338 ( .A(memory[501]), .B(memory[485]), .C(memory[469]), .D(
        memory[453]), .S0(n1460), .S1(n1439), .Y(n1215) );
  MX4X1 U339 ( .A(memory[1013]), .B(memory[997]), .C(memory[981]), .D(
        memory[965]), .S0(n1461), .S1(n1440), .Y(n1225) );
  MX4X1 U340 ( .A(memory[502]), .B(memory[486]), .C(memory[470]), .D(
        memory[454]), .S0(n1462), .S1(n1441), .Y(n1235) );
  MX4X1 U341 ( .A(memory[1014]), .B(memory[998]), .C(memory[982]), .D(
        memory[966]), .S0(n1462), .S1(n1441), .Y(n1245) );
  MX4X1 U342 ( .A(memory[503]), .B(memory[487]), .C(memory[471]), .D(
        memory[455]), .S0(n1463), .S1(n1442), .Y(n1255) );
  MX4X1 U343 ( .A(memory[1015]), .B(memory[999]), .C(memory[983]), .D(
        memory[967]), .S0(n1464), .S1(n1443), .Y(n1265) );
  MX4X1 U344 ( .A(memory[504]), .B(memory[488]), .C(memory[472]), .D(
        memory[456]), .S0(n1464), .S1(n1443), .Y(n1275) );
  MX4X1 U345 ( .A(memory[1016]), .B(memory[1000]), .C(memory[984]), .D(
        memory[968]), .S0(n1460), .S1(n1444), .Y(n1285) );
  MX4X1 U346 ( .A(memory[505]), .B(memory[489]), .C(memory[473]), .D(
        memory[457]), .S0(n1455), .S1(n1445), .Y(n1295) );
  MX4X1 U347 ( .A(memory[1017]), .B(memory[1001]), .C(memory[985]), .D(
        memory[969]), .S0(n1464), .S1(n1445), .Y(n1305) );
  MX4X1 U348 ( .A(memory[506]), .B(memory[490]), .C(memory[474]), .D(
        memory[458]), .S0(n1465), .S1(n1446), .Y(n1315) );
  MX4X1 U349 ( .A(memory[1018]), .B(memory[1002]), .C(memory[986]), .D(
        memory[970]), .S0(n1466), .S1(n1447), .Y(n1325) );
  MX4X1 U350 ( .A(memory[507]), .B(memory[491]), .C(memory[475]), .D(
        memory[459]), .S0(n1466), .S1(n1447), .Y(n1335) );
  MX4X1 U351 ( .A(memory[1019]), .B(memory[1003]), .C(memory[987]), .D(
        memory[971]), .S0(n1467), .S1(n1448), .Y(n1345) );
  MX4X1 U352 ( .A(memory[508]), .B(memory[492]), .C(memory[476]), .D(
        memory[460]), .S0(n1459), .S1(n1449), .Y(n1355) );
  MX4X1 U353 ( .A(memory[1020]), .B(memory[1004]), .C(memory[988]), .D(
        memory[972]), .S0(n1470), .S1(n1449), .Y(n1365) );
  MX4X1 U354 ( .A(memory[509]), .B(memory[493]), .C(memory[477]), .D(
        memory[461]), .S0(n1468), .S1(n1450), .Y(n1375) );
  MX4X1 U355 ( .A(memory[1021]), .B(memory[1005]), .C(memory[989]), .D(
        memory[973]), .S0(n1469), .S1(n1436), .Y(n1385) );
  MX4X1 U356 ( .A(memory[510]), .B(memory[494]), .C(memory[478]), .D(
        memory[462]), .S0(n1469), .S1(n1450), .Y(n1395) );
  MX4X1 U357 ( .A(memory[1022]), .B(memory[1006]), .C(memory[990]), .D(
        memory[974]), .S0(n1470), .S1(n1451), .Y(n1405) );
  MX4X1 U358 ( .A(memory[511]), .B(memory[495]), .C(memory[479]), .D(
        memory[463]), .S0(n1468), .S1(n1452), .Y(n1415) );
  MX4X1 U359 ( .A(memory[1023]), .B(memory[1007]), .C(memory[991]), .D(
        memory[975]), .S0(n1470), .S1(n1452), .Y(n1425) );
  MX4X1 U360 ( .A(memory[560]), .B(memory[544]), .C(memory[528]), .D(
        memory[512]), .S0(n1454), .S1(n1450), .Y(n91) );
  MX4X1 U361 ( .A(memory[304]), .B(memory[288]), .C(memory[272]), .D(
        memory[256]), .S0(n1454), .S1(n1451), .Y(n85) );
  MX4X1 U362 ( .A(memory[816]), .B(memory[800]), .C(memory[784]), .D(
        memory[768]), .S0(n1454), .S1(n1450), .Y(n97) );
  MX4X1 U363 ( .A(memory[48]), .B(memory[32]), .C(memory[16]), .D(memory[0]), 
        .S0(n1455), .S1(n1451), .Y(n80) );
  MX4X1 U364 ( .A(memory[49]), .B(memory[33]), .C(memory[17]), .D(memory[1]), 
        .S0(n1455), .S1(n1434), .Y(n102) );
  MX4X1 U365 ( .A(memory[561]), .B(memory[545]), .C(memory[529]), .D(
        memory[513]), .S0(n1455), .S1(n1434), .Y(n1137) );
  MX4X1 U366 ( .A(memory[305]), .B(memory[289]), .C(memory[273]), .D(
        memory[257]), .S0(n1455), .S1(n1434), .Y(n1132) );
  MX4X1 U367 ( .A(memory[817]), .B(memory[801]), .C(memory[785]), .D(
        memory[769]), .S0(n1456), .S1(n1435), .Y(n1142) );
  MX4X1 U368 ( .A(memory[50]), .B(memory[34]), .C(memory[18]), .D(memory[2]), 
        .S0(n1456), .S1(n1435), .Y(n1147) );
  MX4X1 U369 ( .A(memory[562]), .B(memory[546]), .C(memory[530]), .D(
        memory[514]), .S0(n1457), .S1(n1436), .Y(n1157) );
  MX4X1 U370 ( .A(memory[306]), .B(memory[290]), .C(memory[274]), .D(
        memory[258]), .S0(n1456), .S1(n1435), .Y(n1152) );
  MX4X1 U371 ( .A(memory[818]), .B(memory[802]), .C(memory[786]), .D(
        memory[770]), .S0(n1457), .S1(n1436), .Y(n1162) );
  MX4X1 U372 ( .A(memory[51]), .B(memory[35]), .C(memory[19]), .D(memory[3]), 
        .S0(n1457), .S1(n1436), .Y(n1167) );
  MX4X1 U373 ( .A(memory[563]), .B(memory[547]), .C(memory[531]), .D(
        memory[515]), .S0(n1458), .S1(n1437), .Y(n1177) );
  MX4X1 U374 ( .A(memory[307]), .B(memory[291]), .C(memory[275]), .D(
        memory[259]), .S0(n1458), .S1(n1437), .Y(n1172) );
  MX4X1 U375 ( .A(memory[819]), .B(memory[803]), .C(memory[787]), .D(
        memory[771]), .S0(n1458), .S1(n1437), .Y(n1182) );
  MX4X1 U376 ( .A(memory[52]), .B(memory[36]), .C(memory[20]), .D(memory[4]), 
        .S0(n1459), .S1(n1438), .Y(n1187) );
  MX4X1 U377 ( .A(memory[564]), .B(memory[548]), .C(memory[532]), .D(
        memory[516]), .S0(n1459), .S1(n1438), .Y(n1197) );
  MX4X1 U378 ( .A(memory[308]), .B(memory[292]), .C(memory[276]), .D(
        memory[260]), .S0(n1459), .S1(n1438), .Y(n1192) );
  MX4X1 U379 ( .A(memory[820]), .B(memory[804]), .C(memory[788]), .D(
        memory[772]), .S0(n1460), .S1(n1439), .Y(n1202) );
  MX4X1 U380 ( .A(memory[53]), .B(memory[37]), .C(memory[21]), .D(memory[5]), 
        .S0(n1460), .S1(n1439), .Y(n1207) );
  MX4X1 U381 ( .A(memory[565]), .B(memory[549]), .C(memory[533]), .D(
        memory[517]), .S0(n1461), .S1(n1440), .Y(n1217) );
  MX4X1 U382 ( .A(memory[309]), .B(memory[293]), .C(memory[277]), .D(
        memory[261]), .S0(n1460), .S1(n1439), .Y(n1212) );
  MX4X1 U383 ( .A(memory[821]), .B(memory[805]), .C(memory[789]), .D(
        memory[773]), .S0(n1461), .S1(n1440), .Y(n1222) );
  MX4X1 U384 ( .A(memory[54]), .B(memory[38]), .C(memory[22]), .D(memory[6]), 
        .S0(n1461), .S1(n1440), .Y(n1227) );
  MX4X1 U385 ( .A(memory[566]), .B(memory[550]), .C(memory[534]), .D(
        memory[518]), .S0(n1462), .S1(n1441), .Y(n1237) );
  MX4X1 U386 ( .A(memory[310]), .B(memory[294]), .C(memory[278]), .D(
        memory[262]), .S0(n1462), .S1(n1441), .Y(n1232) );
  MX4X1 U387 ( .A(memory[822]), .B(memory[806]), .C(memory[790]), .D(
        memory[774]), .S0(n1462), .S1(n1441), .Y(n1242) );
  MX4X1 U388 ( .A(memory[55]), .B(memory[39]), .C(memory[23]), .D(memory[7]), 
        .S0(n1463), .S1(n1442), .Y(n1247) );
  MX4X1 U389 ( .A(memory[567]), .B(memory[551]), .C(memory[535]), .D(
        memory[519]), .S0(n1463), .S1(n1442), .Y(n1257) );
  MX4X1 U390 ( .A(memory[311]), .B(memory[295]), .C(memory[279]), .D(
        memory[263]), .S0(n1463), .S1(n1442), .Y(n1252) );
  MX4X1 U391 ( .A(memory[823]), .B(memory[807]), .C(memory[791]), .D(
        memory[775]), .S0(n1464), .S1(n1443), .Y(n1262) );
  MX4X1 U392 ( .A(memory[56]), .B(memory[40]), .C(memory[24]), .D(memory[8]), 
        .S0(n1464), .S1(n1443), .Y(n1267) );
  MX4X1 U393 ( .A(memory[568]), .B(memory[552]), .C(memory[536]), .D(
        memory[520]), .S0(n1461), .S1(n1444), .Y(n1277) );
  MX4X1 U394 ( .A(memory[312]), .B(memory[296]), .C(memory[280]), .D(
        memory[264]), .S0(n1464), .S1(n1443), .Y(n1272) );
  MX4X1 U395 ( .A(memory[824]), .B(memory[808]), .C(memory[792]), .D(
        memory[776]), .S0(n1461), .S1(n1444), .Y(n1282) );
  MX4X1 U396 ( .A(memory[57]), .B(memory[41]), .C(memory[25]), .D(memory[9]), 
        .S0(n1454), .S1(n1444), .Y(n1287) );
  MX4X1 U397 ( .A(memory[569]), .B(memory[553]), .C(memory[537]), .D(
        memory[521]), .S0(n1463), .S1(n1445), .Y(n1297) );
  MX4X1 U398 ( .A(memory[313]), .B(memory[297]), .C(memory[281]), .D(
        memory[265]), .S0(n1460), .S1(n1445), .Y(n1292) );
  MX4X1 U399 ( .A(memory[825]), .B(memory[809]), .C(memory[793]), .D(
        memory[777]), .S0(n1454), .S1(n1445), .Y(n1302) );
  MX4X1 U400 ( .A(memory[58]), .B(memory[42]), .C(memory[26]), .D(memory[10]), 
        .S0(n1465), .S1(n1446), .Y(n1307) );
  MX4X1 U401 ( .A(memory[570]), .B(memory[554]), .C(memory[538]), .D(
        memory[522]), .S0(n1465), .S1(n1446), .Y(n1317) );
  MX4X1 U402 ( .A(memory[314]), .B(memory[298]), .C(memory[282]), .D(
        memory[266]), .S0(n1465), .S1(n1446), .Y(n1312) );
  MX4X1 U403 ( .A(memory[826]), .B(memory[810]), .C(memory[794]), .D(
        memory[778]), .S0(n1466), .S1(n1447), .Y(n1322) );
  MX4X1 U404 ( .A(memory[59]), .B(memory[43]), .C(memory[27]), .D(memory[11]), 
        .S0(n1466), .S1(n1447), .Y(n1327) );
  MX4X1 U405 ( .A(memory[571]), .B(memory[555]), .C(memory[539]), .D(
        memory[523]), .S0(n1467), .S1(n1448), .Y(n1337) );
  MX4X1 U406 ( .A(memory[315]), .B(memory[299]), .C(memory[283]), .D(
        memory[267]), .S0(n1466), .S1(n1447), .Y(n1332) );
  MX4X1 U407 ( .A(memory[827]), .B(memory[811]), .C(memory[795]), .D(
        memory[779]), .S0(n1467), .S1(n1448), .Y(n1342) );
  MX4X1 U408 ( .A(memory[60]), .B(memory[44]), .C(memory[28]), .D(memory[12]), 
        .S0(n1467), .S1(n1448), .Y(n1347) );
  MX4X1 U409 ( .A(memory[572]), .B(memory[556]), .C(memory[540]), .D(
        memory[524]), .S0(n1461), .S1(n1449), .Y(n1357) );
  MX4X1 U410 ( .A(memory[316]), .B(memory[300]), .C(memory[284]), .D(
        memory[268]), .S0(n1470), .S1(n1449), .Y(n1352) );
  MX4X1 U411 ( .A(memory[828]), .B(memory[812]), .C(memory[796]), .D(
        memory[780]), .S0(n1468), .S1(n1449), .Y(n1362) );
  MX4X1 U412 ( .A(memory[61]), .B(memory[45]), .C(memory[29]), .D(memory[13]), 
        .S0(n1468), .S1(n1450), .Y(n1367) );
  MX4X1 U413 ( .A(memory[573]), .B(memory[557]), .C(memory[541]), .D(
        memory[525]), .S0(n1468), .S1(n1450), .Y(n1377) );
  MX4X1 U414 ( .A(memory[317]), .B(memory[301]), .C(memory[285]), .D(
        memory[269]), .S0(n1468), .S1(n1450), .Y(n1372) );
  MX4X1 U415 ( .A(memory[829]), .B(memory[813]), .C(memory[797]), .D(
        memory[781]), .S0(n1469), .S1(n1451), .Y(n1382) );
  MX4X1 U416 ( .A(memory[62]), .B(memory[46]), .C(memory[30]), .D(memory[14]), 
        .S0(n1469), .S1(n1450), .Y(n1387) );
  MX4X1 U417 ( .A(memory[574]), .B(memory[558]), .C(memory[542]), .D(
        memory[526]), .S0(n1470), .S1(n1451), .Y(n1397) );
  MX4X1 U418 ( .A(memory[318]), .B(memory[302]), .C(memory[286]), .D(
        memory[270]), .S0(n1469), .S1(n1451), .Y(n1392) );
  MX4X1 U419 ( .A(memory[830]), .B(memory[814]), .C(memory[798]), .D(
        memory[782]), .S0(n1470), .S1(n1451), .Y(n1402) );
  MX4X1 U420 ( .A(memory[63]), .B(memory[47]), .C(memory[31]), .D(memory[15]), 
        .S0(n1470), .S1(n1451), .Y(n1407) );
  MX4X1 U421 ( .A(memory[575]), .B(memory[559]), .C(memory[543]), .D(
        memory[527]), .S0(n1470), .S1(n1452), .Y(n1417) );
  MX4X1 U422 ( .A(memory[319]), .B(memory[303]), .C(memory[287]), .D(
        memory[271]), .S0(n1459), .S1(n1452), .Y(n1412) );
  MX4X1 U423 ( .A(memory[831]), .B(memory[815]), .C(memory[799]), .D(
        memory[783]), .S0(n1456), .S1(n1452), .Y(n1422) );
  MX4X1 U424 ( .A(n1130), .B(n1128), .C(n1129), .D(n102), .S0(n1427), .S1(
        n1431), .Y(n1131) );
  MX4X1 U425 ( .A(memory[241]), .B(memory[225]), .C(memory[209]), .D(
        memory[193]), .S0(n1455), .S1(n1434), .Y(n1130) );
  MX4X1 U426 ( .A(memory[113]), .B(memory[97]), .C(memory[81]), .D(memory[65]), 
        .S0(n1455), .S1(n1434), .Y(n1128) );
  MX4X1 U427 ( .A(memory[177]), .B(memory[161]), .C(memory[145]), .D(
        memory[129]), .S0(n1455), .S1(n1434), .Y(n1129) );
  MX4X1 U428 ( .A(n1150), .B(n1148), .C(n1149), .D(n1147), .S0(n1427), .S1(
        n1431), .Y(n1151) );
  MX4X1 U429 ( .A(memory[242]), .B(memory[226]), .C(memory[210]), .D(
        memory[194]), .S0(n1456), .S1(n1435), .Y(n1150) );
  MX4X1 U430 ( .A(memory[114]), .B(memory[98]), .C(memory[82]), .D(memory[66]), 
        .S0(n1456), .S1(n1435), .Y(n1148) );
  MX4X1 U431 ( .A(memory[178]), .B(memory[162]), .C(memory[146]), .D(
        memory[130]), .S0(n1456), .S1(n1435), .Y(n1149) );
  MX4X1 U432 ( .A(n1170), .B(n1168), .C(n1169), .D(n1167), .S0(n1427), .S1(
        n1431), .Y(n1171) );
  MX4X1 U433 ( .A(memory[243]), .B(memory[227]), .C(memory[211]), .D(
        memory[195]), .S0(n1457), .S1(n1436), .Y(n1170) );
  MX4X1 U434 ( .A(memory[115]), .B(memory[99]), .C(memory[83]), .D(memory[67]), 
        .S0(n1457), .S1(n1436), .Y(n1168) );
  MX4X1 U435 ( .A(memory[179]), .B(memory[163]), .C(memory[147]), .D(
        memory[131]), .S0(n1457), .S1(n1436), .Y(n1169) );
  MX4X1 U436 ( .A(n1190), .B(n1188), .C(n1189), .D(n1187), .S0(n1428), .S1(
        n1432), .Y(n1191) );
  MX4X1 U437 ( .A(memory[244]), .B(memory[228]), .C(memory[212]), .D(
        memory[196]), .S0(n1459), .S1(n1438), .Y(n1190) );
  MX4X1 U438 ( .A(memory[116]), .B(memory[100]), .C(memory[84]), .D(memory[68]), .S0(n1459), .S1(n1438), .Y(n1188) );
  MX4X1 U439 ( .A(memory[180]), .B(memory[164]), .C(memory[148]), .D(
        memory[132]), .S0(n1459), .S1(n1438), .Y(n1189) );
  MX4X1 U440 ( .A(n1210), .B(n1208), .C(n1209), .D(n1207), .S0(n1428), .S1(
        n1432), .Y(n1211) );
  MX4X1 U441 ( .A(memory[245]), .B(memory[229]), .C(memory[213]), .D(
        memory[197]), .S0(n1460), .S1(n1439), .Y(n1210) );
  MX4X1 U442 ( .A(memory[117]), .B(memory[101]), .C(memory[85]), .D(memory[69]), .S0(n1460), .S1(n1439), .Y(n1208) );
  MX4X1 U443 ( .A(memory[181]), .B(memory[165]), .C(memory[149]), .D(
        memory[133]), .S0(n1460), .S1(n1439), .Y(n1209) );
  MX4X1 U444 ( .A(n1230), .B(n1228), .C(n1229), .D(n1227), .S0(n1428), .S1(
        n1432), .Y(n1231) );
  MX4X1 U445 ( .A(memory[246]), .B(memory[230]), .C(memory[214]), .D(
        memory[198]), .S0(n1461), .S1(n1440), .Y(n1230) );
  MX4X1 U446 ( .A(memory[118]), .B(memory[102]), .C(memory[86]), .D(memory[70]), .S0(n1461), .S1(n1440), .Y(n1228) );
  MX4X1 U447 ( .A(memory[182]), .B(memory[166]), .C(memory[150]), .D(
        memory[134]), .S0(n1461), .S1(n1440), .Y(n1229) );
  MX4X1 U448 ( .A(n1250), .B(n1248), .C(n1249), .D(n1247), .S0(n1429), .S1(
        n1431), .Y(n1251) );
  MX4X1 U449 ( .A(memory[247]), .B(memory[231]), .C(memory[215]), .D(
        memory[199]), .S0(n1463), .S1(n1442), .Y(n1250) );
  MX4X1 U450 ( .A(memory[119]), .B(memory[103]), .C(memory[87]), .D(memory[71]), .S0(n1463), .S1(n1442), .Y(n1248) );
  MX4X1 U451 ( .A(memory[183]), .B(memory[167]), .C(memory[151]), .D(
        memory[135]), .S0(n1463), .S1(n1442), .Y(n1249) );
  MX4X1 U452 ( .A(n1270), .B(n1268), .C(n1269), .D(n1267), .S0(n1429), .S1(
        n1432), .Y(n1271) );
  MX4X1 U453 ( .A(memory[248]), .B(memory[232]), .C(memory[216]), .D(
        memory[200]), .S0(n1464), .S1(n1443), .Y(n1270) );
  MX4X1 U454 ( .A(memory[120]), .B(memory[104]), .C(memory[88]), .D(memory[72]), .S0(n1464), .S1(n1443), .Y(n1268) );
  MX4X1 U455 ( .A(memory[184]), .B(memory[168]), .C(memory[152]), .D(
        memory[136]), .S0(n1464), .S1(n1443), .Y(n1269) );
  MX4X1 U456 ( .A(n1290), .B(n1288), .C(n1289), .D(n1287), .S0(n1429), .S1(
        addr[2]), .Y(n1291) );
  MX4X1 U457 ( .A(memory[249]), .B(memory[233]), .C(memory[217]), .D(
        memory[201]), .S0(n1454), .S1(n1444), .Y(n1290) );
  MX4X1 U458 ( .A(memory[121]), .B(memory[105]), .C(memory[89]), .D(memory[73]), .S0(n1459), .S1(n1444), .Y(n1288) );
  MX4X1 U459 ( .A(memory[185]), .B(memory[169]), .C(memory[153]), .D(
        memory[137]), .S0(n1460), .S1(n1444), .Y(n1289) );
  MX4X1 U460 ( .A(n1310), .B(n1308), .C(n1309), .D(n1307), .S0(n1430), .S1(
        n1431), .Y(n1311) );
  MX4X1 U461 ( .A(memory[250]), .B(memory[234]), .C(memory[218]), .D(
        memory[202]), .S0(n1465), .S1(n1446), .Y(n1310) );
  MX4X1 U462 ( .A(memory[122]), .B(memory[106]), .C(memory[90]), .D(memory[74]), .S0(n1465), .S1(n1446), .Y(n1308) );
  MX4X1 U463 ( .A(memory[186]), .B(memory[170]), .C(memory[154]), .D(
        memory[138]), .S0(n1465), .S1(n1446), .Y(n1309) );
  MX4X1 U464 ( .A(n1330), .B(n1328), .C(n1329), .D(n1327), .S0(n1430), .S1(
        n1432), .Y(n1331) );
  MX4X1 U465 ( .A(memory[251]), .B(memory[235]), .C(memory[219]), .D(
        memory[203]), .S0(n1466), .S1(n1447), .Y(n1330) );
  MX4X1 U466 ( .A(memory[123]), .B(memory[107]), .C(memory[91]), .D(memory[75]), .S0(n1466), .S1(n1447), .Y(n1328) );
  MX4X1 U467 ( .A(memory[187]), .B(memory[171]), .C(memory[155]), .D(
        memory[139]), .S0(n1466), .S1(n1447), .Y(n1329) );
  MX4X1 U468 ( .A(n1350), .B(n1348), .C(n1349), .D(n1347), .S0(n1430), .S1(
        addr[2]), .Y(n1351) );
  MX4X1 U469 ( .A(memory[252]), .B(memory[236]), .C(memory[220]), .D(
        memory[204]), .S0(n1467), .S1(n1448), .Y(n1350) );
  MX4X1 U470 ( .A(memory[124]), .B(memory[108]), .C(memory[92]), .D(memory[76]), .S0(n1467), .S1(n1448), .Y(n1348) );
  MX4X1 U471 ( .A(memory[188]), .B(memory[172]), .C(memory[156]), .D(
        memory[140]), .S0(n1467), .S1(n1448), .Y(n1349) );
  MX4X1 U472 ( .A(n1370), .B(n1368), .C(n1369), .D(n1367), .S0(n1429), .S1(
        n1431), .Y(n1371) );
  MX4X1 U473 ( .A(memory[253]), .B(memory[237]), .C(memory[221]), .D(
        memory[205]), .S0(n1468), .S1(n1450), .Y(n1370) );
  MX4X1 U474 ( .A(memory[125]), .B(memory[109]), .C(memory[93]), .D(memory[77]), .S0(n1468), .S1(n1450), .Y(n1368) );
  MX4X1 U475 ( .A(memory[189]), .B(memory[173]), .C(memory[157]), .D(
        memory[141]), .S0(n1468), .S1(n1450), .Y(n1369) );
  MX4X1 U476 ( .A(n1390), .B(n1388), .C(n1389), .D(n1387), .S0(n1430), .S1(
        n1432), .Y(n1391) );
  MX4X1 U477 ( .A(memory[254]), .B(memory[238]), .C(memory[222]), .D(
        memory[206]), .S0(n1469), .S1(n1450), .Y(n1390) );
  MX4X1 U478 ( .A(memory[126]), .B(memory[110]), .C(memory[94]), .D(memory[78]), .S0(n1469), .S1(n1450), .Y(n1388) );
  MX4X1 U479 ( .A(memory[190]), .B(memory[174]), .C(memory[158]), .D(
        memory[142]), .S0(n1469), .S1(n1450), .Y(n1389) );
  MX4X1 U480 ( .A(n1410), .B(n1408), .C(n1409), .D(n1407), .S0(n1428), .S1(
        addr[2]), .Y(n1411) );
  MX4X1 U481 ( .A(memory[255]), .B(memory[239]), .C(memory[223]), .D(
        memory[207]), .S0(n1470), .S1(n1451), .Y(n1410) );
  MX4X1 U482 ( .A(memory[127]), .B(memory[111]), .C(memory[95]), .D(memory[79]), .S0(n1470), .S1(n1451), .Y(n1408) );
  MX4X1 U483 ( .A(memory[191]), .B(memory[175]), .C(memory[159]), .D(
        memory[143]), .S0(n1470), .S1(n1451), .Y(n1409) );
  MX4X1 U484 ( .A(memory[880]), .B(memory[864]), .C(memory[848]), .D(
        memory[832]), .S0(n1454), .S1(n1450), .Y(n98) );
  MX4X1 U485 ( .A(memory[112]), .B(memory[96]), .C(memory[80]), .D(memory[64]), 
        .S0(n1468), .S1(n1450), .Y(n81) );
  MX4X1 U486 ( .A(memory[369]), .B(memory[353]), .C(memory[337]), .D(
        memory[321]), .S0(n1455), .S1(n1434), .Y(n1133) );
  MX4X1 U487 ( .A(memory[881]), .B(memory[865]), .C(memory[849]), .D(
        memory[833]), .S0(n1456), .S1(n1435), .Y(n1143) );
  MX4X1 U488 ( .A(memory[370]), .B(memory[354]), .C(memory[338]), .D(
        memory[322]), .S0(n1456), .S1(n1435), .Y(n1153) );
  MX4X1 U489 ( .A(memory[882]), .B(memory[866]), .C(memory[850]), .D(
        memory[834]), .S0(n1457), .S1(n1436), .Y(n1163) );
  MX4X1 U490 ( .A(memory[371]), .B(memory[355]), .C(memory[339]), .D(
        memory[323]), .S0(n1458), .S1(n1437), .Y(n1173) );
  MX4X1 U491 ( .A(memory[883]), .B(memory[867]), .C(memory[851]), .D(
        memory[835]), .S0(n1458), .S1(n1437), .Y(n1183) );
  MX4X1 U492 ( .A(memory[372]), .B(memory[356]), .C(memory[340]), .D(
        memory[324]), .S0(n1459), .S1(n1438), .Y(n1193) );
  MX4X1 U493 ( .A(memory[884]), .B(memory[868]), .C(memory[852]), .D(
        memory[836]), .S0(n1460), .S1(n1439), .Y(n1203) );
  MX4X1 U494 ( .A(memory[373]), .B(memory[357]), .C(memory[341]), .D(
        memory[325]), .S0(n1460), .S1(n1439), .Y(n1213) );
  MX4X1 U495 ( .A(memory[885]), .B(memory[869]), .C(memory[853]), .D(
        memory[837]), .S0(n1461), .S1(n1440), .Y(n1223) );
  MX4X1 U496 ( .A(memory[374]), .B(memory[358]), .C(memory[342]), .D(
        memory[326]), .S0(n1462), .S1(n1441), .Y(n1233) );
  MX4X1 U497 ( .A(memory[886]), .B(memory[870]), .C(memory[854]), .D(
        memory[838]), .S0(n1462), .S1(n1441), .Y(n1243) );
  MX4X1 U498 ( .A(memory[375]), .B(memory[359]), .C(memory[343]), .D(
        memory[327]), .S0(n1463), .S1(n1442), .Y(n1253) );
  MX4X1 U499 ( .A(memory[887]), .B(memory[871]), .C(memory[855]), .D(
        memory[839]), .S0(n1464), .S1(n1443), .Y(n1263) );
  MX4X1 U500 ( .A(memory[376]), .B(memory[360]), .C(memory[344]), .D(
        memory[328]), .S0(n1464), .S1(n1443), .Y(n1273) );
  MX4X1 U501 ( .A(memory[888]), .B(memory[872]), .C(memory[856]), .D(
        memory[840]), .S0(n1454), .S1(n1444), .Y(n1283) );
  MX4X1 U502 ( .A(memory[377]), .B(memory[361]), .C(memory[345]), .D(
        memory[329]), .S0(n1457), .S1(n1445), .Y(n1293) );
  MX4X1 U503 ( .A(memory[889]), .B(memory[873]), .C(memory[857]), .D(
        memory[841]), .S0(n1463), .S1(n1445), .Y(n1303) );
  MX4X1 U504 ( .A(memory[378]), .B(memory[362]), .C(memory[346]), .D(
        memory[330]), .S0(n1465), .S1(n1446), .Y(n1313) );
  MX4X1 U505 ( .A(memory[890]), .B(memory[874]), .C(memory[858]), .D(
        memory[842]), .S0(n1466), .S1(n1447), .Y(n1323) );
  MX4X1 U506 ( .A(memory[379]), .B(memory[363]), .C(memory[347]), .D(
        memory[331]), .S0(n1466), .S1(n1447), .Y(n1333) );
  MX4X1 U507 ( .A(memory[891]), .B(memory[875]), .C(memory[859]), .D(
        memory[843]), .S0(n1467), .S1(n1448), .Y(n1343) );
  MX4X1 U508 ( .A(memory[380]), .B(memory[364]), .C(memory[348]), .D(
        memory[332]), .S0(n1461), .S1(n1449), .Y(n1353) );
  MX4X1 U509 ( .A(memory[892]), .B(memory[876]), .C(memory[860]), .D(
        memory[844]), .S0(n1462), .S1(n1449), .Y(n1363) );
  MX4X1 U510 ( .A(memory[381]), .B(memory[365]), .C(memory[349]), .D(
        memory[333]), .S0(n1468), .S1(n1450), .Y(n1373) );
  MX4X1 U511 ( .A(memory[893]), .B(memory[877]), .C(memory[861]), .D(
        memory[845]), .S0(n1469), .S1(n1444), .Y(n1383) );
  MX4X1 U512 ( .A(memory[382]), .B(memory[366]), .C(memory[350]), .D(
        memory[334]), .S0(n1469), .S1(n1451), .Y(n1393) );
  MX4X1 U513 ( .A(memory[894]), .B(memory[878]), .C(memory[862]), .D(
        memory[846]), .S0(n1470), .S1(n1451), .Y(n1403) );
  MX4X1 U514 ( .A(memory[383]), .B(memory[367]), .C(memory[351]), .D(
        memory[335]), .S0(n1470), .S1(n1452), .Y(n1413) );
  MX4X1 U515 ( .A(memory[895]), .B(memory[879]), .C(memory[863]), .D(
        memory[847]), .S0(n1469), .S1(n1452), .Y(n1423) );
  MX4X1 U516 ( .A(n89), .B(n87), .C(n88), .D(n85), .S0(n1429), .S1(n1431), .Y(
        n90) );
  MX4X1 U517 ( .A(memory[496]), .B(memory[480]), .C(memory[464]), .D(
        memory[448]), .S0(n1454), .S1(addr[1]), .Y(n89) );
  MX4X1 U518 ( .A(memory[368]), .B(memory[352]), .C(memory[336]), .D(
        memory[320]), .S0(n1454), .S1(n1451), .Y(n87) );
  MX4X1 U519 ( .A(memory[432]), .B(memory[416]), .C(memory[400]), .D(
        memory[384]), .S0(n1454), .S1(n1451), .Y(n88) );
  OAI2BB2X1 U520 ( .B0(n1), .B1(n1505), .A0N(memory[0]), .A1N(n1), .Y(n2535)
         );
  OAI2BB2X1 U521 ( .B0(n1), .B1(n1503), .A0N(memory[1]), .A1N(n1), .Y(n2534)
         );
  OAI2BB2X1 U522 ( .B0(n1), .B1(n1501), .A0N(memory[2]), .A1N(n1), .Y(n2533)
         );
  OAI2BB2X1 U523 ( .B0(n1), .B1(n1499), .A0N(memory[3]), .A1N(n1), .Y(n2532)
         );
  OAI2BB2X1 U524 ( .B0(n1), .B1(n1497), .A0N(memory[4]), .A1N(n1), .Y(n2531)
         );
  OAI2BB2X1 U525 ( .B0(n1), .B1(n1495), .A0N(memory[5]), .A1N(n1), .Y(n2530)
         );
  OAI2BB2X1 U526 ( .B0(n1), .B1(n1493), .A0N(memory[6]), .A1N(n1), .Y(n2529)
         );
  OAI2BB2X1 U527 ( .B0(n1), .B1(n1491), .A0N(memory[7]), .A1N(n1), .Y(n2528)
         );
  OAI2BB2X1 U528 ( .B0(n1), .B1(n1489), .A0N(memory[8]), .A1N(n1), .Y(n2527)
         );
  OAI2BB2X1 U529 ( .B0(n1), .B1(n1487), .A0N(memory[9]), .A1N(n1), .Y(n2526)
         );
  OAI2BB2X1 U530 ( .B0(n1), .B1(n1485), .A0N(memory[10]), .A1N(n1), .Y(n2525)
         );
  OAI2BB2X1 U531 ( .B0(n1), .B1(n1483), .A0N(memory[11]), .A1N(n1), .Y(n2524)
         );
  OAI2BB2X1 U532 ( .B0(n1), .B1(n1481), .A0N(memory[12]), .A1N(n1), .Y(n2523)
         );
  OAI2BB2X1 U533 ( .B0(n1), .B1(n1479), .A0N(memory[13]), .A1N(n1), .Y(n2522)
         );
  OAI2BB2X1 U534 ( .B0(n1), .B1(n1477), .A0N(memory[14]), .A1N(n1), .Y(n2521)
         );
  OAI2BB2X1 U535 ( .B0(n1), .B1(n1475), .A0N(memory[15]), .A1N(n1), .Y(n2520)
         );
  OAI2BB2X1 U536 ( .B0(n1504), .B1(n2), .A0N(memory[16]), .A1N(n2), .Y(n2519)
         );
  OAI2BB2X1 U537 ( .B0(n1502), .B1(n2), .A0N(memory[17]), .A1N(n2), .Y(n2518)
         );
  OAI2BB2X1 U538 ( .B0(n1500), .B1(n2), .A0N(memory[18]), .A1N(n2), .Y(n2517)
         );
  OAI2BB2X1 U539 ( .B0(n1498), .B1(n2), .A0N(memory[19]), .A1N(n2), .Y(n2516)
         );
  OAI2BB2X1 U540 ( .B0(n1496), .B1(n2), .A0N(memory[20]), .A1N(n2), .Y(n2515)
         );
  OAI2BB2X1 U541 ( .B0(n1494), .B1(n2), .A0N(memory[21]), .A1N(n2), .Y(n2514)
         );
  OAI2BB2X1 U542 ( .B0(n1492), .B1(n2), .A0N(memory[22]), .A1N(n2), .Y(n2513)
         );
  OAI2BB2X1 U543 ( .B0(n1490), .B1(n2), .A0N(memory[23]), .A1N(n2), .Y(n2512)
         );
  OAI2BB2X1 U544 ( .B0(n1480), .B1(n2), .A0N(memory[28]), .A1N(n2), .Y(n2507)
         );
  OAI2BB2X1 U545 ( .B0(n1478), .B1(n2), .A0N(memory[29]), .A1N(n2), .Y(n2506)
         );
  OAI2BB2X1 U546 ( .B0(n1476), .B1(n2), .A0N(memory[30]), .A1N(n2), .Y(n2505)
         );
  OAI2BB2X1 U547 ( .B0(n1474), .B1(n2), .A0N(memory[31]), .A1N(n2), .Y(n2504)
         );
  OAI2BB2X1 U548 ( .B0(n1504), .B1(n57), .A0N(memory[32]), .A1N(n57), .Y(n2503) );
  OAI2BB2X1 U549 ( .B0(n1502), .B1(n57), .A0N(memory[33]), .A1N(n57), .Y(n2502) );
  OAI2BB2X1 U550 ( .B0(n1500), .B1(n57), .A0N(memory[34]), .A1N(n57), .Y(n2501) );
  OAI2BB2X1 U551 ( .B0(n1498), .B1(n57), .A0N(memory[35]), .A1N(n57), .Y(n2500) );
  OAI2BB2X1 U552 ( .B0(n1496), .B1(n57), .A0N(memory[36]), .A1N(n57), .Y(n2499) );
  OAI2BB2X1 U553 ( .B0(n1494), .B1(n57), .A0N(memory[37]), .A1N(n57), .Y(n2498) );
  OAI2BB2X1 U554 ( .B0(n1492), .B1(n57), .A0N(memory[38]), .A1N(n57), .Y(n2497) );
  OAI2BB2X1 U555 ( .B0(n1490), .B1(n57), .A0N(memory[39]), .A1N(n57), .Y(n2496) );
  OAI2BB2X1 U556 ( .B0(n1480), .B1(n57), .A0N(memory[44]), .A1N(n57), .Y(n2491) );
  OAI2BB2X1 U557 ( .B0(n1478), .B1(n57), .A0N(memory[45]), .A1N(n57), .Y(n2490) );
  OAI2BB2X1 U558 ( .B0(n1476), .B1(n57), .A0N(memory[46]), .A1N(n57), .Y(n2489) );
  OAI2BB2X1 U559 ( .B0(n1474), .B1(n57), .A0N(memory[47]), .A1N(n57), .Y(n2488) );
  OAI2BB2X1 U560 ( .B0(n1505), .B1(n58), .A0N(memory[48]), .A1N(n58), .Y(n2487) );
  OAI2BB2X1 U561 ( .B0(n1503), .B1(n58), .A0N(memory[49]), .A1N(n58), .Y(n2486) );
  OAI2BB2X1 U562 ( .B0(n1501), .B1(n58), .A0N(memory[50]), .A1N(n58), .Y(n2485) );
  OAI2BB2X1 U563 ( .B0(n1499), .B1(n58), .A0N(memory[51]), .A1N(n58), .Y(n2484) );
  OAI2BB2X1 U564 ( .B0(n1497), .B1(n58), .A0N(memory[52]), .A1N(n58), .Y(n2483) );
  OAI2BB2X1 U565 ( .B0(n1495), .B1(n58), .A0N(memory[53]), .A1N(n58), .Y(n2482) );
  OAI2BB2X1 U566 ( .B0(n1493), .B1(n58), .A0N(memory[54]), .A1N(n58), .Y(n2481) );
  OAI2BB2X1 U567 ( .B0(n1491), .B1(n58), .A0N(memory[55]), .A1N(n58), .Y(n2480) );
  OAI2BB2X1 U568 ( .B0(n1481), .B1(n58), .A0N(memory[60]), .A1N(n58), .Y(n2475) );
  OAI2BB2X1 U569 ( .B0(n1479), .B1(n58), .A0N(memory[61]), .A1N(n58), .Y(n2474) );
  OAI2BB2X1 U570 ( .B0(n1477), .B1(n58), .A0N(memory[62]), .A1N(n58), .Y(n2473) );
  OAI2BB2X1 U571 ( .B0(n1475), .B1(n58), .A0N(memory[63]), .A1N(n58), .Y(n2472) );
  OAI2BB2X1 U572 ( .B0(n1504), .B1(n60), .A0N(memory[64]), .A1N(n60), .Y(n2471) );
  OAI2BB2X1 U573 ( .B0(n1502), .B1(n60), .A0N(memory[65]), .A1N(n60), .Y(n2470) );
  OAI2BB2X1 U574 ( .B0(n1500), .B1(n60), .A0N(memory[66]), .A1N(n60), .Y(n2469) );
  OAI2BB2X1 U575 ( .B0(n1498), .B1(n60), .A0N(memory[67]), .A1N(n60), .Y(n2468) );
  OAI2BB2X1 U576 ( .B0(n1496), .B1(n60), .A0N(memory[68]), .A1N(n60), .Y(n2467) );
  OAI2BB2X1 U577 ( .B0(n1494), .B1(n60), .A0N(memory[69]), .A1N(n60), .Y(n2466) );
  OAI2BB2X1 U578 ( .B0(n1492), .B1(n60), .A0N(memory[70]), .A1N(n60), .Y(n2465) );
  OAI2BB2X1 U579 ( .B0(n1490), .B1(n60), .A0N(memory[71]), .A1N(n60), .Y(n2464) );
  OAI2BB2X1 U580 ( .B0(n1480), .B1(n60), .A0N(memory[76]), .A1N(n60), .Y(n2459) );
  OAI2BB2X1 U581 ( .B0(n1478), .B1(n60), .A0N(memory[77]), .A1N(n60), .Y(n2458) );
  OAI2BB2X1 U582 ( .B0(n1476), .B1(n60), .A0N(memory[78]), .A1N(n60), .Y(n2457) );
  OAI2BB2X1 U583 ( .B0(n1474), .B1(n60), .A0N(memory[79]), .A1N(n60), .Y(n2456) );
  OAI2BB2X1 U584 ( .B0(n1505), .B1(n61), .A0N(memory[80]), .A1N(n61), .Y(n2455) );
  OAI2BB2X1 U585 ( .B0(n1503), .B1(n61), .A0N(memory[81]), .A1N(n61), .Y(n2454) );
  OAI2BB2X1 U586 ( .B0(n1501), .B1(n61), .A0N(memory[82]), .A1N(n61), .Y(n2453) );
  OAI2BB2X1 U587 ( .B0(n1499), .B1(n61), .A0N(memory[83]), .A1N(n61), .Y(n2452) );
  OAI2BB2X1 U588 ( .B0(n1497), .B1(n61), .A0N(memory[84]), .A1N(n61), .Y(n2451) );
  OAI2BB2X1 U589 ( .B0(n1495), .B1(n61), .A0N(memory[85]), .A1N(n61), .Y(n2450) );
  OAI2BB2X1 U590 ( .B0(n1493), .B1(n61), .A0N(memory[86]), .A1N(n61), .Y(n2449) );
  OAI2BB2X1 U591 ( .B0(n1491), .B1(n61), .A0N(memory[87]), .A1N(n61), .Y(n2448) );
  OAI2BB2X1 U592 ( .B0(n1481), .B1(n61), .A0N(memory[92]), .A1N(n61), .Y(n2443) );
  OAI2BB2X1 U593 ( .B0(n1479), .B1(n61), .A0N(memory[93]), .A1N(n61), .Y(n2442) );
  OAI2BB2X1 U594 ( .B0(n1477), .B1(n61), .A0N(memory[94]), .A1N(n61), .Y(n2441) );
  OAI2BB2X1 U595 ( .B0(n1475), .B1(n61), .A0N(memory[95]), .A1N(n61), .Y(n2440) );
  OAI2BB2X1 U596 ( .B0(n1504), .B1(n62), .A0N(memory[96]), .A1N(n62), .Y(n2439) );
  OAI2BB2X1 U597 ( .B0(n1502), .B1(n62), .A0N(memory[97]), .A1N(n62), .Y(n2438) );
  OAI2BB2X1 U598 ( .B0(n1500), .B1(n62), .A0N(memory[98]), .A1N(n62), .Y(n2437) );
  OAI2BB2X1 U599 ( .B0(n1498), .B1(n62), .A0N(memory[99]), .A1N(n62), .Y(n2436) );
  OAI2BB2X1 U600 ( .B0(n1496), .B1(n62), .A0N(memory[100]), .A1N(n62), .Y(
        n2435) );
  OAI2BB2X1 U601 ( .B0(n1494), .B1(n62), .A0N(memory[101]), .A1N(n62), .Y(
        n2434) );
  OAI2BB2X1 U602 ( .B0(n1492), .B1(n62), .A0N(memory[102]), .A1N(n62), .Y(
        n2433) );
  OAI2BB2X1 U603 ( .B0(n1490), .B1(n62), .A0N(memory[103]), .A1N(n62), .Y(
        n2432) );
  OAI2BB2X1 U604 ( .B0(n1480), .B1(n62), .A0N(memory[108]), .A1N(n62), .Y(
        n2427) );
  OAI2BB2X1 U605 ( .B0(n1478), .B1(n62), .A0N(memory[109]), .A1N(n62), .Y(
        n2426) );
  OAI2BB2X1 U606 ( .B0(n1476), .B1(n62), .A0N(memory[110]), .A1N(n62), .Y(
        n2425) );
  OAI2BB2X1 U607 ( .B0(n1474), .B1(n62), .A0N(memory[111]), .A1N(n62), .Y(
        n2424) );
  OAI2BB2X1 U608 ( .B0(n1505), .B1(n3), .A0N(memory[112]), .A1N(n3), .Y(n2423)
         );
  OAI2BB2X1 U609 ( .B0(n1503), .B1(n3), .A0N(memory[113]), .A1N(n3), .Y(n2422)
         );
  OAI2BB2X1 U610 ( .B0(n1501), .B1(n3), .A0N(memory[114]), .A1N(n3), .Y(n2421)
         );
  OAI2BB2X1 U611 ( .B0(n1499), .B1(n3), .A0N(memory[115]), .A1N(n3), .Y(n2420)
         );
  OAI2BB2X1 U612 ( .B0(n1497), .B1(n3), .A0N(memory[116]), .A1N(n3), .Y(n2419)
         );
  OAI2BB2X1 U613 ( .B0(n1495), .B1(n3), .A0N(memory[117]), .A1N(n3), .Y(n2418)
         );
  OAI2BB2X1 U614 ( .B0(n1493), .B1(n3), .A0N(memory[118]), .A1N(n3), .Y(n2417)
         );
  OAI2BB2X1 U615 ( .B0(n1491), .B1(n3), .A0N(memory[119]), .A1N(n3), .Y(n2416)
         );
  OAI2BB2X1 U616 ( .B0(n1481), .B1(n3), .A0N(memory[124]), .A1N(n3), .Y(n2411)
         );
  OAI2BB2X1 U617 ( .B0(n1479), .B1(n3), .A0N(memory[125]), .A1N(n3), .Y(n2410)
         );
  OAI2BB2X1 U618 ( .B0(n1477), .B1(n3), .A0N(memory[126]), .A1N(n3), .Y(n2409)
         );
  OAI2BB2X1 U619 ( .B0(n1475), .B1(n3), .A0N(memory[127]), .A1N(n3), .Y(n2408)
         );
  OAI2BB2X1 U620 ( .B0(n1505), .B1(n4), .A0N(memory[128]), .A1N(n4), .Y(n2407)
         );
  OAI2BB2X1 U621 ( .B0(n1503), .B1(n4), .A0N(memory[129]), .A1N(n4), .Y(n2406)
         );
  OAI2BB2X1 U622 ( .B0(n1501), .B1(n4), .A0N(memory[130]), .A1N(n4), .Y(n2405)
         );
  OAI2BB2X1 U623 ( .B0(n1499), .B1(n4), .A0N(memory[131]), .A1N(n4), .Y(n2404)
         );
  OAI2BB2X1 U624 ( .B0(n1497), .B1(n4), .A0N(memory[132]), .A1N(n4), .Y(n2403)
         );
  OAI2BB2X1 U625 ( .B0(n1495), .B1(n4), .A0N(memory[133]), .A1N(n4), .Y(n2402)
         );
  OAI2BB2X1 U626 ( .B0(n1493), .B1(n4), .A0N(memory[134]), .A1N(n4), .Y(n2401)
         );
  OAI2BB2X1 U627 ( .B0(n1491), .B1(n4), .A0N(memory[135]), .A1N(n4), .Y(n2400)
         );
  OAI2BB2X1 U628 ( .B0(n1481), .B1(n4), .A0N(memory[140]), .A1N(n4), .Y(n2395)
         );
  OAI2BB2X1 U629 ( .B0(n1479), .B1(n4), .A0N(memory[141]), .A1N(n4), .Y(n2394)
         );
  OAI2BB2X1 U630 ( .B0(n1477), .B1(n4), .A0N(memory[142]), .A1N(n4), .Y(n2393)
         );
  OAI2BB2X1 U631 ( .B0(n1475), .B1(n4), .A0N(memory[143]), .A1N(n4), .Y(n2392)
         );
  OAI2BB2X1 U632 ( .B0(n1505), .B1(n5), .A0N(memory[144]), .A1N(n5), .Y(n2391)
         );
  OAI2BB2X1 U633 ( .B0(n1503), .B1(n5), .A0N(memory[145]), .A1N(n5), .Y(n2390)
         );
  OAI2BB2X1 U634 ( .B0(n1501), .B1(n5), .A0N(memory[146]), .A1N(n5), .Y(n2389)
         );
  OAI2BB2X1 U635 ( .B0(n1499), .B1(n5), .A0N(memory[147]), .A1N(n5), .Y(n2388)
         );
  OAI2BB2X1 U636 ( .B0(n1497), .B1(n5), .A0N(memory[148]), .A1N(n5), .Y(n2387)
         );
  OAI2BB2X1 U637 ( .B0(n1495), .B1(n5), .A0N(memory[149]), .A1N(n5), .Y(n2386)
         );
  OAI2BB2X1 U638 ( .B0(n1493), .B1(n5), .A0N(memory[150]), .A1N(n5), .Y(n2385)
         );
  OAI2BB2X1 U639 ( .B0(n1491), .B1(n5), .A0N(memory[151]), .A1N(n5), .Y(n2384)
         );
  OAI2BB2X1 U640 ( .B0(n1481), .B1(n5), .A0N(memory[156]), .A1N(n5), .Y(n2379)
         );
  OAI2BB2X1 U641 ( .B0(n1479), .B1(n5), .A0N(memory[157]), .A1N(n5), .Y(n2378)
         );
  OAI2BB2X1 U642 ( .B0(n1477), .B1(n5), .A0N(memory[158]), .A1N(n5), .Y(n2377)
         );
  OAI2BB2X1 U643 ( .B0(n1475), .B1(n5), .A0N(memory[159]), .A1N(n5), .Y(n2376)
         );
  OAI2BB2X1 U644 ( .B0(n1504), .B1(n63), .A0N(memory[160]), .A1N(n63), .Y(
        n2375) );
  OAI2BB2X1 U645 ( .B0(n1502), .B1(n63), .A0N(memory[161]), .A1N(n63), .Y(
        n2374) );
  OAI2BB2X1 U646 ( .B0(n1500), .B1(n63), .A0N(memory[162]), .A1N(n63), .Y(
        n2373) );
  OAI2BB2X1 U647 ( .B0(n1498), .B1(n63), .A0N(memory[163]), .A1N(n63), .Y(
        n2372) );
  OAI2BB2X1 U648 ( .B0(n1496), .B1(n63), .A0N(memory[164]), .A1N(n63), .Y(
        n2371) );
  OAI2BB2X1 U649 ( .B0(n1494), .B1(n63), .A0N(memory[165]), .A1N(n63), .Y(
        n2370) );
  OAI2BB2X1 U650 ( .B0(n1492), .B1(n63), .A0N(memory[166]), .A1N(n63), .Y(
        n2369) );
  OAI2BB2X1 U651 ( .B0(n1490), .B1(n63), .A0N(memory[167]), .A1N(n63), .Y(
        n2368) );
  OAI2BB2X1 U652 ( .B0(n1480), .B1(n63), .A0N(memory[172]), .A1N(n63), .Y(
        n2363) );
  OAI2BB2X1 U653 ( .B0(n1478), .B1(n63), .A0N(memory[173]), .A1N(n63), .Y(
        n2362) );
  OAI2BB2X1 U654 ( .B0(n1476), .B1(n63), .A0N(memory[174]), .A1N(n63), .Y(
        n2361) );
  OAI2BB2X1 U655 ( .B0(n1474), .B1(n63), .A0N(memory[175]), .A1N(n63), .Y(
        n2360) );
  OAI2BB2X1 U656 ( .B0(n1505), .B1(n64), .A0N(memory[176]), .A1N(n64), .Y(
        n2359) );
  OAI2BB2X1 U657 ( .B0(n1503), .B1(n64), .A0N(memory[177]), .A1N(n64), .Y(
        n2358) );
  OAI2BB2X1 U658 ( .B0(n1501), .B1(n64), .A0N(memory[178]), .A1N(n64), .Y(
        n2357) );
  OAI2BB2X1 U659 ( .B0(n1499), .B1(n64), .A0N(memory[179]), .A1N(n64), .Y(
        n2356) );
  OAI2BB2X1 U660 ( .B0(n1497), .B1(n64), .A0N(memory[180]), .A1N(n64), .Y(
        n2355) );
  OAI2BB2X1 U661 ( .B0(n1495), .B1(n64), .A0N(memory[181]), .A1N(n64), .Y(
        n2354) );
  OAI2BB2X1 U662 ( .B0(n1493), .B1(n64), .A0N(memory[182]), .A1N(n64), .Y(
        n2353) );
  OAI2BB2X1 U663 ( .B0(n1491), .B1(n64), .A0N(memory[183]), .A1N(n64), .Y(
        n2352) );
  OAI2BB2X1 U664 ( .B0(n1481), .B1(n64), .A0N(memory[188]), .A1N(n64), .Y(
        n2347) );
  OAI2BB2X1 U665 ( .B0(n1479), .B1(n64), .A0N(memory[189]), .A1N(n64), .Y(
        n2346) );
  OAI2BB2X1 U666 ( .B0(n1477), .B1(n64), .A0N(memory[190]), .A1N(n64), .Y(
        n2345) );
  OAI2BB2X1 U667 ( .B0(n1475), .B1(n64), .A0N(memory[191]), .A1N(n64), .Y(
        n2344) );
  OAI2BB2X1 U668 ( .B0(n1505), .B1(n65), .A0N(memory[192]), .A1N(n65), .Y(
        n2343) );
  OAI2BB2X1 U669 ( .B0(n1503), .B1(n65), .A0N(memory[193]), .A1N(n65), .Y(
        n2342) );
  OAI2BB2X1 U670 ( .B0(n1501), .B1(n65), .A0N(memory[194]), .A1N(n65), .Y(
        n2341) );
  OAI2BB2X1 U671 ( .B0(n1499), .B1(n65), .A0N(memory[195]), .A1N(n65), .Y(
        n2340) );
  OAI2BB2X1 U672 ( .B0(n1497), .B1(n65), .A0N(memory[196]), .A1N(n65), .Y(
        n2339) );
  OAI2BB2X1 U673 ( .B0(n1495), .B1(n65), .A0N(memory[197]), .A1N(n65), .Y(
        n2338) );
  OAI2BB2X1 U674 ( .B0(n1493), .B1(n65), .A0N(memory[198]), .A1N(n65), .Y(
        n2337) );
  OAI2BB2X1 U675 ( .B0(n1491), .B1(n65), .A0N(memory[199]), .A1N(n65), .Y(
        n2336) );
  OAI2BB2X1 U676 ( .B0(n1481), .B1(n65), .A0N(memory[204]), .A1N(n65), .Y(
        n2331) );
  OAI2BB2X1 U677 ( .B0(n1479), .B1(n65), .A0N(memory[205]), .A1N(n65), .Y(
        n2330) );
  OAI2BB2X1 U678 ( .B0(n1477), .B1(n65), .A0N(memory[206]), .A1N(n65), .Y(
        n2329) );
  OAI2BB2X1 U679 ( .B0(n1475), .B1(n65), .A0N(memory[207]), .A1N(n65), .Y(
        n2328) );
  OAI2BB2X1 U680 ( .B0(n1505), .B1(n66), .A0N(memory[208]), .A1N(n66), .Y(
        n2327) );
  OAI2BB2X1 U681 ( .B0(n1503), .B1(n66), .A0N(memory[209]), .A1N(n66), .Y(
        n2326) );
  OAI2BB2X1 U682 ( .B0(n1501), .B1(n66), .A0N(memory[210]), .A1N(n66), .Y(
        n2325) );
  OAI2BB2X1 U683 ( .B0(n1499), .B1(n66), .A0N(memory[211]), .A1N(n66), .Y(
        n2324) );
  OAI2BB2X1 U684 ( .B0(n1497), .B1(n66), .A0N(memory[212]), .A1N(n66), .Y(
        n2323) );
  OAI2BB2X1 U685 ( .B0(n1495), .B1(n66), .A0N(memory[213]), .A1N(n66), .Y(
        n2322) );
  OAI2BB2X1 U686 ( .B0(n1493), .B1(n66), .A0N(memory[214]), .A1N(n66), .Y(
        n2321) );
  OAI2BB2X1 U687 ( .B0(n1491), .B1(n66), .A0N(memory[215]), .A1N(n66), .Y(
        n2320) );
  OAI2BB2X1 U688 ( .B0(n1481), .B1(n66), .A0N(memory[220]), .A1N(n66), .Y(
        n2315) );
  OAI2BB2X1 U689 ( .B0(n1479), .B1(n66), .A0N(memory[221]), .A1N(n66), .Y(
        n2314) );
  OAI2BB2X1 U690 ( .B0(n1477), .B1(n66), .A0N(memory[222]), .A1N(n66), .Y(
        n2313) );
  OAI2BB2X1 U691 ( .B0(n1475), .B1(n66), .A0N(memory[223]), .A1N(n66), .Y(
        n2312) );
  OAI2BB2X1 U692 ( .B0(n1505), .B1(n67), .A0N(memory[224]), .A1N(n67), .Y(
        n2311) );
  OAI2BB2X1 U693 ( .B0(n1503), .B1(n67), .A0N(memory[225]), .A1N(n67), .Y(
        n2310) );
  OAI2BB2X1 U694 ( .B0(n1501), .B1(n67), .A0N(memory[226]), .A1N(n67), .Y(
        n2309) );
  OAI2BB2X1 U695 ( .B0(n1499), .B1(n67), .A0N(memory[227]), .A1N(n67), .Y(
        n2308) );
  OAI2BB2X1 U696 ( .B0(n1497), .B1(n67), .A0N(memory[228]), .A1N(n67), .Y(
        n2307) );
  OAI2BB2X1 U697 ( .B0(n1495), .B1(n67), .A0N(memory[229]), .A1N(n67), .Y(
        n2306) );
  OAI2BB2X1 U698 ( .B0(n1493), .B1(n67), .A0N(memory[230]), .A1N(n67), .Y(
        n2305) );
  OAI2BB2X1 U699 ( .B0(n1491), .B1(n67), .A0N(memory[231]), .A1N(n67), .Y(
        n2304) );
  OAI2BB2X1 U700 ( .B0(n1481), .B1(n67), .A0N(memory[236]), .A1N(n67), .Y(
        n2299) );
  OAI2BB2X1 U701 ( .B0(n1479), .B1(n67), .A0N(memory[237]), .A1N(n67), .Y(
        n2298) );
  OAI2BB2X1 U702 ( .B0(n1477), .B1(n67), .A0N(memory[238]), .A1N(n67), .Y(
        n2297) );
  OAI2BB2X1 U703 ( .B0(n1475), .B1(n67), .A0N(memory[239]), .A1N(n67), .Y(
        n2296) );
  OAI2BB2X1 U704 ( .B0(n1505), .B1(n6), .A0N(memory[240]), .A1N(n6), .Y(n2295)
         );
  OAI2BB2X1 U705 ( .B0(n1503), .B1(n6), .A0N(memory[241]), .A1N(n6), .Y(n2294)
         );
  OAI2BB2X1 U706 ( .B0(n1501), .B1(n6), .A0N(memory[242]), .A1N(n6), .Y(n2293)
         );
  OAI2BB2X1 U707 ( .B0(n1499), .B1(n6), .A0N(memory[243]), .A1N(n6), .Y(n2292)
         );
  OAI2BB2X1 U708 ( .B0(n1497), .B1(n6), .A0N(memory[244]), .A1N(n6), .Y(n2291)
         );
  OAI2BB2X1 U709 ( .B0(n1495), .B1(n6), .A0N(memory[245]), .A1N(n6), .Y(n2290)
         );
  OAI2BB2X1 U710 ( .B0(n1493), .B1(n6), .A0N(memory[246]), .A1N(n6), .Y(n2289)
         );
  OAI2BB2X1 U711 ( .B0(n1491), .B1(n6), .A0N(memory[247]), .A1N(n6), .Y(n2288)
         );
  OAI2BB2X1 U712 ( .B0(n1481), .B1(n6), .A0N(memory[252]), .A1N(n6), .Y(n2283)
         );
  OAI2BB2X1 U713 ( .B0(n1479), .B1(n6), .A0N(memory[253]), .A1N(n6), .Y(n2282)
         );
  OAI2BB2X1 U714 ( .B0(n1477), .B1(n6), .A0N(memory[254]), .A1N(n6), .Y(n2281)
         );
  OAI2BB2X1 U715 ( .B0(n1475), .B1(n6), .A0N(memory[255]), .A1N(n6), .Y(n2280)
         );
  OAI2BB2X1 U716 ( .B0(n1505), .B1(n7), .A0N(memory[256]), .A1N(n7), .Y(n2279)
         );
  OAI2BB2X1 U717 ( .B0(n1503), .B1(n7), .A0N(memory[257]), .A1N(n7), .Y(n2278)
         );
  OAI2BB2X1 U718 ( .B0(n1501), .B1(n7), .A0N(memory[258]), .A1N(n7), .Y(n2277)
         );
  OAI2BB2X1 U719 ( .B0(n1499), .B1(n7), .A0N(memory[259]), .A1N(n7), .Y(n2276)
         );
  OAI2BB2X1 U720 ( .B0(n1497), .B1(n7), .A0N(memory[260]), .A1N(n7), .Y(n2275)
         );
  OAI2BB2X1 U721 ( .B0(n1495), .B1(n7), .A0N(memory[261]), .A1N(n7), .Y(n2274)
         );
  OAI2BB2X1 U722 ( .B0(n1493), .B1(n7), .A0N(memory[262]), .A1N(n7), .Y(n2273)
         );
  OAI2BB2X1 U723 ( .B0(n1491), .B1(n7), .A0N(memory[263]), .A1N(n7), .Y(n2272)
         );
  OAI2BB2X1 U724 ( .B0(n1481), .B1(n7), .A0N(memory[268]), .A1N(n7), .Y(n2267)
         );
  OAI2BB2X1 U725 ( .B0(n1479), .B1(n7), .A0N(memory[269]), .A1N(n7), .Y(n2266)
         );
  OAI2BB2X1 U726 ( .B0(n1477), .B1(n7), .A0N(memory[270]), .A1N(n7), .Y(n2265)
         );
  OAI2BB2X1 U727 ( .B0(n1475), .B1(n7), .A0N(memory[271]), .A1N(n7), .Y(n2264)
         );
  OAI2BB2X1 U728 ( .B0(n1505), .B1(n8), .A0N(memory[272]), .A1N(n8), .Y(n2263)
         );
  OAI2BB2X1 U729 ( .B0(n1503), .B1(n8), .A0N(memory[273]), .A1N(n8), .Y(n2262)
         );
  OAI2BB2X1 U730 ( .B0(n1501), .B1(n8), .A0N(memory[274]), .A1N(n8), .Y(n2261)
         );
  OAI2BB2X1 U731 ( .B0(n1499), .B1(n8), .A0N(memory[275]), .A1N(n8), .Y(n2260)
         );
  OAI2BB2X1 U732 ( .B0(n1497), .B1(n8), .A0N(memory[276]), .A1N(n8), .Y(n2259)
         );
  OAI2BB2X1 U733 ( .B0(n1495), .B1(n8), .A0N(memory[277]), .A1N(n8), .Y(n2258)
         );
  OAI2BB2X1 U734 ( .B0(n1493), .B1(n8), .A0N(memory[278]), .A1N(n8), .Y(n2257)
         );
  OAI2BB2X1 U735 ( .B0(n1491), .B1(n8), .A0N(memory[279]), .A1N(n8), .Y(n2256)
         );
  OAI2BB2X1 U736 ( .B0(n1481), .B1(n8), .A0N(memory[284]), .A1N(n8), .Y(n2251)
         );
  OAI2BB2X1 U737 ( .B0(n1479), .B1(n8), .A0N(memory[285]), .A1N(n8), .Y(n2250)
         );
  OAI2BB2X1 U738 ( .B0(n1477), .B1(n8), .A0N(memory[286]), .A1N(n8), .Y(n2249)
         );
  OAI2BB2X1 U739 ( .B0(n1475), .B1(n8), .A0N(memory[287]), .A1N(n8), .Y(n2248)
         );
  OAI2BB2X1 U740 ( .B0(n1505), .B1(n69), .A0N(memory[288]), .A1N(n69), .Y(
        n2247) );
  OAI2BB2X1 U741 ( .B0(n1503), .B1(n69), .A0N(memory[289]), .A1N(n69), .Y(
        n2246) );
  OAI2BB2X1 U742 ( .B0(n1501), .B1(n69), .A0N(memory[290]), .A1N(n69), .Y(
        n2245) );
  OAI2BB2X1 U743 ( .B0(n1499), .B1(n69), .A0N(memory[291]), .A1N(n69), .Y(
        n2244) );
  OAI2BB2X1 U744 ( .B0(n1497), .B1(n69), .A0N(memory[292]), .A1N(n69), .Y(
        n2243) );
  OAI2BB2X1 U745 ( .B0(n1495), .B1(n69), .A0N(memory[293]), .A1N(n69), .Y(
        n2242) );
  OAI2BB2X1 U746 ( .B0(n1493), .B1(n69), .A0N(memory[294]), .A1N(n69), .Y(
        n2241) );
  OAI2BB2X1 U747 ( .B0(n1491), .B1(n69), .A0N(memory[295]), .A1N(n69), .Y(
        n2240) );
  OAI2BB2X1 U748 ( .B0(n1481), .B1(n69), .A0N(memory[300]), .A1N(n69), .Y(
        n2235) );
  OAI2BB2X1 U749 ( .B0(n1479), .B1(n69), .A0N(memory[301]), .A1N(n69), .Y(
        n2234) );
  OAI2BB2X1 U750 ( .B0(n1477), .B1(n69), .A0N(memory[302]), .A1N(n69), .Y(
        n2233) );
  OAI2BB2X1 U751 ( .B0(n1475), .B1(n69), .A0N(memory[303]), .A1N(n69), .Y(
        n2232) );
  OAI2BB2X1 U752 ( .B0(n1505), .B1(n70), .A0N(memory[304]), .A1N(n70), .Y(
        n2231) );
  OAI2BB2X1 U753 ( .B0(n1503), .B1(n70), .A0N(memory[305]), .A1N(n70), .Y(
        n2230) );
  OAI2BB2X1 U754 ( .B0(n1501), .B1(n70), .A0N(memory[306]), .A1N(n70), .Y(
        n2229) );
  OAI2BB2X1 U755 ( .B0(n1499), .B1(n70), .A0N(memory[307]), .A1N(n70), .Y(
        n2228) );
  OAI2BB2X1 U756 ( .B0(n1497), .B1(n70), .A0N(memory[308]), .A1N(n70), .Y(
        n2227) );
  OAI2BB2X1 U757 ( .B0(n1495), .B1(n70), .A0N(memory[309]), .A1N(n70), .Y(
        n2226) );
  OAI2BB2X1 U758 ( .B0(n1493), .B1(n70), .A0N(memory[310]), .A1N(n70), .Y(
        n2225) );
  OAI2BB2X1 U759 ( .B0(n1491), .B1(n70), .A0N(memory[311]), .A1N(n70), .Y(
        n2224) );
  OAI2BB2X1 U760 ( .B0(n1481), .B1(n70), .A0N(memory[316]), .A1N(n70), .Y(
        n2219) );
  OAI2BB2X1 U761 ( .B0(n1479), .B1(n70), .A0N(memory[317]), .A1N(n70), .Y(
        n2218) );
  OAI2BB2X1 U762 ( .B0(n1477), .B1(n70), .A0N(memory[318]), .A1N(n70), .Y(
        n2217) );
  OAI2BB2X1 U763 ( .B0(n1475), .B1(n70), .A0N(memory[319]), .A1N(n70), .Y(
        n2216) );
  OAI2BB2X1 U764 ( .B0(n1505), .B1(n71), .A0N(memory[320]), .A1N(n71), .Y(
        n2215) );
  OAI2BB2X1 U765 ( .B0(n1503), .B1(n71), .A0N(memory[321]), .A1N(n71), .Y(
        n2214) );
  OAI2BB2X1 U766 ( .B0(n1501), .B1(n71), .A0N(memory[322]), .A1N(n71), .Y(
        n2213) );
  OAI2BB2X1 U767 ( .B0(n1499), .B1(n71), .A0N(memory[323]), .A1N(n71), .Y(
        n2212) );
  OAI2BB2X1 U768 ( .B0(n1497), .B1(n71), .A0N(memory[324]), .A1N(n71), .Y(
        n2211) );
  OAI2BB2X1 U769 ( .B0(n1495), .B1(n71), .A0N(memory[325]), .A1N(n71), .Y(
        n2210) );
  OAI2BB2X1 U770 ( .B0(n1493), .B1(n71), .A0N(memory[326]), .A1N(n71), .Y(
        n2209) );
  OAI2BB2X1 U771 ( .B0(n1491), .B1(n71), .A0N(memory[327]), .A1N(n71), .Y(
        n2208) );
  OAI2BB2X1 U772 ( .B0(n1481), .B1(n71), .A0N(memory[332]), .A1N(n71), .Y(
        n2203) );
  OAI2BB2X1 U773 ( .B0(n1479), .B1(n71), .A0N(memory[333]), .A1N(n71), .Y(
        n2202) );
  OAI2BB2X1 U774 ( .B0(n1477), .B1(n71), .A0N(memory[334]), .A1N(n71), .Y(
        n2201) );
  OAI2BB2X1 U775 ( .B0(n1475), .B1(n71), .A0N(memory[335]), .A1N(n71), .Y(
        n2200) );
  OAI2BB2X1 U776 ( .B0(n1505), .B1(n72), .A0N(memory[336]), .A1N(n72), .Y(
        n2199) );
  OAI2BB2X1 U777 ( .B0(n1503), .B1(n72), .A0N(memory[337]), .A1N(n72), .Y(
        n2198) );
  OAI2BB2X1 U778 ( .B0(n1501), .B1(n72), .A0N(memory[338]), .A1N(n72), .Y(
        n2197) );
  OAI2BB2X1 U779 ( .B0(n1499), .B1(n72), .A0N(memory[339]), .A1N(n72), .Y(
        n2196) );
  OAI2BB2X1 U780 ( .B0(n1497), .B1(n72), .A0N(memory[340]), .A1N(n72), .Y(
        n2195) );
  OAI2BB2X1 U781 ( .B0(n1495), .B1(n72), .A0N(memory[341]), .A1N(n72), .Y(
        n2194) );
  OAI2BB2X1 U782 ( .B0(n1493), .B1(n72), .A0N(memory[342]), .A1N(n72), .Y(
        n2193) );
  OAI2BB2X1 U783 ( .B0(n1491), .B1(n72), .A0N(memory[343]), .A1N(n72), .Y(
        n2192) );
  OAI2BB2X1 U784 ( .B0(n1481), .B1(n72), .A0N(memory[348]), .A1N(n72), .Y(
        n2187) );
  OAI2BB2X1 U785 ( .B0(n1479), .B1(n72), .A0N(memory[349]), .A1N(n72), .Y(
        n2186) );
  OAI2BB2X1 U786 ( .B0(n1477), .B1(n72), .A0N(memory[350]), .A1N(n72), .Y(
        n2185) );
  OAI2BB2X1 U787 ( .B0(n1475), .B1(n72), .A0N(memory[351]), .A1N(n72), .Y(
        n2184) );
  OAI2BB2X1 U788 ( .B0(n1505), .B1(n73), .A0N(memory[352]), .A1N(n73), .Y(
        n2183) );
  OAI2BB2X1 U789 ( .B0(n1503), .B1(n73), .A0N(memory[353]), .A1N(n73), .Y(
        n2182) );
  OAI2BB2X1 U790 ( .B0(n1501), .B1(n73), .A0N(memory[354]), .A1N(n73), .Y(
        n2181) );
  OAI2BB2X1 U791 ( .B0(n1499), .B1(n73), .A0N(memory[355]), .A1N(n73), .Y(
        n2180) );
  OAI2BB2X1 U792 ( .B0(n1497), .B1(n73), .A0N(memory[356]), .A1N(n73), .Y(
        n2179) );
  OAI2BB2X1 U793 ( .B0(n1495), .B1(n73), .A0N(memory[357]), .A1N(n73), .Y(
        n2178) );
  OAI2BB2X1 U794 ( .B0(n1493), .B1(n73), .A0N(memory[358]), .A1N(n73), .Y(
        n2177) );
  OAI2BB2X1 U795 ( .B0(n1491), .B1(n73), .A0N(memory[359]), .A1N(n73), .Y(
        n2176) );
  OAI2BB2X1 U796 ( .B0(n1481), .B1(n73), .A0N(memory[364]), .A1N(n73), .Y(
        n2171) );
  OAI2BB2X1 U797 ( .B0(n1479), .B1(n73), .A0N(memory[365]), .A1N(n73), .Y(
        n2170) );
  OAI2BB2X1 U798 ( .B0(n1477), .B1(n73), .A0N(memory[366]), .A1N(n73), .Y(
        n2169) );
  OAI2BB2X1 U799 ( .B0(n1475), .B1(n73), .A0N(memory[367]), .A1N(n73), .Y(
        n2168) );
  OAI2BB2X1 U800 ( .B0(n1505), .B1(n9), .A0N(memory[368]), .A1N(n9), .Y(n2167)
         );
  OAI2BB2X1 U801 ( .B0(n1503), .B1(n9), .A0N(memory[369]), .A1N(n9), .Y(n2166)
         );
  OAI2BB2X1 U802 ( .B0(n1501), .B1(n9), .A0N(memory[370]), .A1N(n9), .Y(n2165)
         );
  OAI2BB2X1 U803 ( .B0(n1499), .B1(n9), .A0N(memory[371]), .A1N(n9), .Y(n2164)
         );
  OAI2BB2X1 U804 ( .B0(n1497), .B1(n9), .A0N(memory[372]), .A1N(n9), .Y(n2163)
         );
  OAI2BB2X1 U805 ( .B0(n1495), .B1(n9), .A0N(memory[373]), .A1N(n9), .Y(n2162)
         );
  OAI2BB2X1 U806 ( .B0(n1493), .B1(n9), .A0N(memory[374]), .A1N(n9), .Y(n2161)
         );
  OAI2BB2X1 U807 ( .B0(n1491), .B1(n9), .A0N(memory[375]), .A1N(n9), .Y(n2160)
         );
  OAI2BB2X1 U808 ( .B0(n1481), .B1(n9), .A0N(memory[380]), .A1N(n9), .Y(n2155)
         );
  OAI2BB2X1 U809 ( .B0(n1479), .B1(n9), .A0N(memory[381]), .A1N(n9), .Y(n2154)
         );
  OAI2BB2X1 U810 ( .B0(n1477), .B1(n9), .A0N(memory[382]), .A1N(n9), .Y(n2153)
         );
  OAI2BB2X1 U811 ( .B0(n1475), .B1(n9), .A0N(memory[383]), .A1N(n9), .Y(n2152)
         );
  OAI2BB2X1 U812 ( .B0(n1505), .B1(n10), .A0N(memory[384]), .A1N(n10), .Y(
        n2151) );
  OAI2BB2X1 U813 ( .B0(n1503), .B1(n10), .A0N(memory[385]), .A1N(n10), .Y(
        n2150) );
  OAI2BB2X1 U814 ( .B0(n1501), .B1(n10), .A0N(memory[386]), .A1N(n10), .Y(
        n2149) );
  OAI2BB2X1 U815 ( .B0(n1499), .B1(n10), .A0N(memory[387]), .A1N(n10), .Y(
        n2148) );
  OAI2BB2X1 U816 ( .B0(n1497), .B1(n10), .A0N(memory[388]), .A1N(n10), .Y(
        n2147) );
  OAI2BB2X1 U817 ( .B0(n1495), .B1(n10), .A0N(memory[389]), .A1N(n10), .Y(
        n2146) );
  OAI2BB2X1 U818 ( .B0(n1493), .B1(n10), .A0N(memory[390]), .A1N(n10), .Y(
        n2145) );
  OAI2BB2X1 U819 ( .B0(n1491), .B1(n10), .A0N(memory[391]), .A1N(n10), .Y(
        n2144) );
  OAI2BB2X1 U820 ( .B0(n1481), .B1(n10), .A0N(memory[396]), .A1N(n10), .Y(
        n2139) );
  OAI2BB2X1 U821 ( .B0(n1479), .B1(n10), .A0N(memory[397]), .A1N(n10), .Y(
        n2138) );
  OAI2BB2X1 U822 ( .B0(n1477), .B1(n10), .A0N(memory[398]), .A1N(n10), .Y(
        n2137) );
  OAI2BB2X1 U823 ( .B0(n1475), .B1(n10), .A0N(memory[399]), .A1N(n10), .Y(
        n2136) );
  OAI2BB2X1 U824 ( .B0(n1504), .B1(n11), .A0N(memory[400]), .A1N(n11), .Y(
        n2135) );
  OAI2BB2X1 U825 ( .B0(n1502), .B1(n11), .A0N(memory[401]), .A1N(n11), .Y(
        n2134) );
  OAI2BB2X1 U826 ( .B0(n1500), .B1(n11), .A0N(memory[402]), .A1N(n11), .Y(
        n2133) );
  OAI2BB2X1 U827 ( .B0(n1498), .B1(n11), .A0N(memory[403]), .A1N(n11), .Y(
        n2132) );
  OAI2BB2X1 U828 ( .B0(n1496), .B1(n11), .A0N(memory[404]), .A1N(n11), .Y(
        n2131) );
  OAI2BB2X1 U829 ( .B0(n1494), .B1(n11), .A0N(memory[405]), .A1N(n11), .Y(
        n2130) );
  OAI2BB2X1 U830 ( .B0(n1492), .B1(n11), .A0N(memory[406]), .A1N(n11), .Y(
        n2129) );
  OAI2BB2X1 U831 ( .B0(n1490), .B1(n11), .A0N(memory[407]), .A1N(n11), .Y(
        n2128) );
  OAI2BB2X1 U832 ( .B0(n1480), .B1(n11), .A0N(memory[412]), .A1N(n11), .Y(
        n2123) );
  OAI2BB2X1 U833 ( .B0(n1478), .B1(n11), .A0N(memory[413]), .A1N(n11), .Y(
        n2122) );
  OAI2BB2X1 U834 ( .B0(n1476), .B1(n11), .A0N(memory[414]), .A1N(n11), .Y(
        n2121) );
  OAI2BB2X1 U835 ( .B0(n1474), .B1(n11), .A0N(memory[415]), .A1N(n11), .Y(
        n2120) );
  OAI2BB2X1 U836 ( .B0(n1505), .B1(n74), .A0N(memory[416]), .A1N(n74), .Y(
        n2119) );
  OAI2BB2X1 U837 ( .B0(n1503), .B1(n74), .A0N(memory[417]), .A1N(n74), .Y(
        n2118) );
  OAI2BB2X1 U838 ( .B0(n1501), .B1(n74), .A0N(memory[418]), .A1N(n74), .Y(
        n2117) );
  OAI2BB2X1 U839 ( .B0(n1499), .B1(n74), .A0N(memory[419]), .A1N(n74), .Y(
        n2116) );
  OAI2BB2X1 U840 ( .B0(n1497), .B1(n74), .A0N(memory[420]), .A1N(n74), .Y(
        n2115) );
  OAI2BB2X1 U841 ( .B0(n1495), .B1(n74), .A0N(memory[421]), .A1N(n74), .Y(
        n2114) );
  OAI2BB2X1 U842 ( .B0(n1493), .B1(n74), .A0N(memory[422]), .A1N(n74), .Y(
        n2113) );
  OAI2BB2X1 U843 ( .B0(n1491), .B1(n74), .A0N(memory[423]), .A1N(n74), .Y(
        n2112) );
  OAI2BB2X1 U844 ( .B0(n1481), .B1(n74), .A0N(memory[428]), .A1N(n74), .Y(
        n2107) );
  OAI2BB2X1 U845 ( .B0(n1479), .B1(n74), .A0N(memory[429]), .A1N(n74), .Y(
        n2106) );
  OAI2BB2X1 U846 ( .B0(n1477), .B1(n74), .A0N(memory[430]), .A1N(n74), .Y(
        n2105) );
  OAI2BB2X1 U847 ( .B0(n1475), .B1(n74), .A0N(memory[431]), .A1N(n74), .Y(
        n2104) );
  OAI2BB2X1 U848 ( .B0(n1505), .B1(n75), .A0N(memory[432]), .A1N(n75), .Y(
        n2103) );
  OAI2BB2X1 U849 ( .B0(n1503), .B1(n75), .A0N(memory[433]), .A1N(n75), .Y(
        n2102) );
  OAI2BB2X1 U850 ( .B0(n1501), .B1(n75), .A0N(memory[434]), .A1N(n75), .Y(
        n2101) );
  OAI2BB2X1 U851 ( .B0(n1499), .B1(n75), .A0N(memory[435]), .A1N(n75), .Y(
        n2100) );
  OAI2BB2X1 U852 ( .B0(n1497), .B1(n75), .A0N(memory[436]), .A1N(n75), .Y(
        n2099) );
  OAI2BB2X1 U853 ( .B0(n1495), .B1(n75), .A0N(memory[437]), .A1N(n75), .Y(
        n2098) );
  OAI2BB2X1 U854 ( .B0(n1493), .B1(n75), .A0N(memory[438]), .A1N(n75), .Y(
        n2097) );
  OAI2BB2X1 U855 ( .B0(n1491), .B1(n75), .A0N(memory[439]), .A1N(n75), .Y(
        n2096) );
  OAI2BB2X1 U856 ( .B0(n1481), .B1(n75), .A0N(memory[444]), .A1N(n75), .Y(
        n2091) );
  OAI2BB2X1 U857 ( .B0(n1479), .B1(n75), .A0N(memory[445]), .A1N(n75), .Y(
        n2090) );
  OAI2BB2X1 U858 ( .B0(n1477), .B1(n75), .A0N(memory[446]), .A1N(n75), .Y(
        n2089) );
  OAI2BB2X1 U859 ( .B0(n1475), .B1(n75), .A0N(memory[447]), .A1N(n75), .Y(
        n2088) );
  OAI2BB2X1 U860 ( .B0(n1505), .B1(n76), .A0N(memory[448]), .A1N(n76), .Y(
        n2087) );
  OAI2BB2X1 U861 ( .B0(n1503), .B1(n76), .A0N(memory[449]), .A1N(n76), .Y(
        n2086) );
  OAI2BB2X1 U862 ( .B0(n1501), .B1(n76), .A0N(memory[450]), .A1N(n76), .Y(
        n2085) );
  OAI2BB2X1 U863 ( .B0(n1499), .B1(n76), .A0N(memory[451]), .A1N(n76), .Y(
        n2084) );
  OAI2BB2X1 U864 ( .B0(n1497), .B1(n76), .A0N(memory[452]), .A1N(n76), .Y(
        n2083) );
  OAI2BB2X1 U865 ( .B0(n1495), .B1(n76), .A0N(memory[453]), .A1N(n76), .Y(
        n2082) );
  OAI2BB2X1 U866 ( .B0(n1493), .B1(n76), .A0N(memory[454]), .A1N(n76), .Y(
        n2081) );
  OAI2BB2X1 U867 ( .B0(n1491), .B1(n76), .A0N(memory[455]), .A1N(n76), .Y(
        n2080) );
  OAI2BB2X1 U868 ( .B0(n1481), .B1(n76), .A0N(memory[460]), .A1N(n76), .Y(
        n2075) );
  OAI2BB2X1 U869 ( .B0(n1479), .B1(n76), .A0N(memory[461]), .A1N(n76), .Y(
        n2074) );
  OAI2BB2X1 U870 ( .B0(n1477), .B1(n76), .A0N(memory[462]), .A1N(n76), .Y(
        n2073) );
  OAI2BB2X1 U871 ( .B0(n1475), .B1(n76), .A0N(memory[463]), .A1N(n76), .Y(
        n2072) );
  OAI2BB2X1 U872 ( .B0(n1504), .B1(n78), .A0N(memory[464]), .A1N(n78), .Y(
        n2071) );
  OAI2BB2X1 U873 ( .B0(n1502), .B1(n78), .A0N(memory[465]), .A1N(n78), .Y(
        n2070) );
  OAI2BB2X1 U874 ( .B0(n1500), .B1(n78), .A0N(memory[466]), .A1N(n78), .Y(
        n2069) );
  OAI2BB2X1 U875 ( .B0(n1498), .B1(n78), .A0N(memory[467]), .A1N(n78), .Y(
        n2068) );
  OAI2BB2X1 U876 ( .B0(n1496), .B1(n78), .A0N(memory[468]), .A1N(n78), .Y(
        n2067) );
  OAI2BB2X1 U877 ( .B0(n1494), .B1(n78), .A0N(memory[469]), .A1N(n78), .Y(
        n2066) );
  OAI2BB2X1 U878 ( .B0(n1492), .B1(n78), .A0N(memory[470]), .A1N(n78), .Y(
        n2065) );
  OAI2BB2X1 U879 ( .B0(n1490), .B1(n78), .A0N(memory[471]), .A1N(n78), .Y(
        n2064) );
  OAI2BB2X1 U880 ( .B0(n1480), .B1(n78), .A0N(memory[476]), .A1N(n78), .Y(
        n2059) );
  OAI2BB2X1 U881 ( .B0(n1478), .B1(n78), .A0N(memory[477]), .A1N(n78), .Y(
        n2058) );
  OAI2BB2X1 U882 ( .B0(n1476), .B1(n78), .A0N(memory[478]), .A1N(n78), .Y(
        n2057) );
  OAI2BB2X1 U883 ( .B0(n1474), .B1(n78), .A0N(memory[479]), .A1N(n78), .Y(
        n2056) );
  OAI2BB2X1 U884 ( .B0(n1505), .B1(n79), .A0N(memory[480]), .A1N(n79), .Y(
        n2055) );
  OAI2BB2X1 U885 ( .B0(n1503), .B1(n79), .A0N(memory[481]), .A1N(n79), .Y(
        n2054) );
  OAI2BB2X1 U886 ( .B0(n1501), .B1(n79), .A0N(memory[482]), .A1N(n79), .Y(
        n2053) );
  OAI2BB2X1 U887 ( .B0(n1499), .B1(n79), .A0N(memory[483]), .A1N(n79), .Y(
        n2052) );
  OAI2BB2X1 U888 ( .B0(n1497), .B1(n79), .A0N(memory[484]), .A1N(n79), .Y(
        n2051) );
  OAI2BB2X1 U889 ( .B0(n1495), .B1(n79), .A0N(memory[485]), .A1N(n79), .Y(
        n2050) );
  OAI2BB2X1 U890 ( .B0(n1493), .B1(n79), .A0N(memory[486]), .A1N(n79), .Y(
        n2049) );
  OAI2BB2X1 U891 ( .B0(n1491), .B1(n79), .A0N(memory[487]), .A1N(n79), .Y(
        n2048) );
  OAI2BB2X1 U892 ( .B0(n1481), .B1(n79), .A0N(memory[492]), .A1N(n79), .Y(
        n2043) );
  OAI2BB2X1 U893 ( .B0(n1479), .B1(n79), .A0N(memory[493]), .A1N(n79), .Y(
        n2042) );
  OAI2BB2X1 U894 ( .B0(n1477), .B1(n79), .A0N(memory[494]), .A1N(n79), .Y(
        n2041) );
  OAI2BB2X1 U895 ( .B0(n1475), .B1(n79), .A0N(memory[495]), .A1N(n79), .Y(
        n2040) );
  OAI2BB2X1 U896 ( .B0(n1504), .B1(n12), .A0N(memory[496]), .A1N(n12), .Y(
        n2039) );
  OAI2BB2X1 U897 ( .B0(n1502), .B1(n12), .A0N(memory[497]), .A1N(n12), .Y(
        n2038) );
  OAI2BB2X1 U898 ( .B0(n1500), .B1(n12), .A0N(memory[498]), .A1N(n12), .Y(
        n2037) );
  OAI2BB2X1 U899 ( .B0(n1498), .B1(n12), .A0N(memory[499]), .A1N(n12), .Y(
        n2036) );
  OAI2BB2X1 U900 ( .B0(n1496), .B1(n12), .A0N(memory[500]), .A1N(n12), .Y(
        n2035) );
  OAI2BB2X1 U901 ( .B0(n1494), .B1(n12), .A0N(memory[501]), .A1N(n12), .Y(
        n2034) );
  OAI2BB2X1 U902 ( .B0(n1492), .B1(n12), .A0N(memory[502]), .A1N(n12), .Y(
        n2033) );
  OAI2BB2X1 U903 ( .B0(n1490), .B1(n12), .A0N(memory[503]), .A1N(n12), .Y(
        n2032) );
  OAI2BB2X1 U904 ( .B0(n1480), .B1(n12), .A0N(memory[508]), .A1N(n12), .Y(
        n2027) );
  OAI2BB2X1 U905 ( .B0(n1478), .B1(n12), .A0N(memory[509]), .A1N(n12), .Y(
        n2026) );
  OAI2BB2X1 U906 ( .B0(n1476), .B1(n12), .A0N(memory[510]), .A1N(n12), .Y(
        n2025) );
  OAI2BB2X1 U907 ( .B0(n1474), .B1(n12), .A0N(memory[511]), .A1N(n12), .Y(
        n2024) );
  OAI2BB2X1 U908 ( .B0(n1505), .B1(n13), .A0N(memory[512]), .A1N(n13), .Y(
        n2023) );
  OAI2BB2X1 U909 ( .B0(n1503), .B1(n13), .A0N(memory[513]), .A1N(n13), .Y(
        n2022) );
  OAI2BB2X1 U910 ( .B0(n1501), .B1(n13), .A0N(memory[514]), .A1N(n13), .Y(
        n2021) );
  OAI2BB2X1 U911 ( .B0(n1499), .B1(n13), .A0N(memory[515]), .A1N(n13), .Y(
        n2020) );
  OAI2BB2X1 U912 ( .B0(n1497), .B1(n13), .A0N(memory[516]), .A1N(n13), .Y(
        n2019) );
  OAI2BB2X1 U913 ( .B0(n1495), .B1(n13), .A0N(memory[517]), .A1N(n13), .Y(
        n2018) );
  OAI2BB2X1 U914 ( .B0(n1493), .B1(n13), .A0N(memory[518]), .A1N(n13), .Y(
        n2017) );
  OAI2BB2X1 U915 ( .B0(n1491), .B1(n13), .A0N(memory[519]), .A1N(n13), .Y(
        n2016) );
  OAI2BB2X1 U916 ( .B0(n1481), .B1(n13), .A0N(memory[524]), .A1N(n13), .Y(
        n2011) );
  OAI2BB2X1 U917 ( .B0(n1479), .B1(n13), .A0N(memory[525]), .A1N(n13), .Y(
        n2010) );
  OAI2BB2X1 U918 ( .B0(n1477), .B1(n13), .A0N(memory[526]), .A1N(n13), .Y(
        n2009) );
  OAI2BB2X1 U919 ( .B0(n1475), .B1(n13), .A0N(memory[527]), .A1N(n13), .Y(
        n2008) );
  OAI2BB2X1 U920 ( .B0(n1504), .B1(n14), .A0N(memory[528]), .A1N(n14), .Y(
        n2007) );
  OAI2BB2X1 U921 ( .B0(n1502), .B1(n14), .A0N(memory[529]), .A1N(n14), .Y(
        n2006) );
  OAI2BB2X1 U922 ( .B0(n1500), .B1(n14), .A0N(memory[530]), .A1N(n14), .Y(
        n2005) );
  OAI2BB2X1 U923 ( .B0(n1498), .B1(n14), .A0N(memory[531]), .A1N(n14), .Y(
        n2004) );
  OAI2BB2X1 U924 ( .B0(n1496), .B1(n14), .A0N(memory[532]), .A1N(n14), .Y(
        n2003) );
  OAI2BB2X1 U925 ( .B0(n1494), .B1(n14), .A0N(memory[533]), .A1N(n14), .Y(
        n2002) );
  OAI2BB2X1 U926 ( .B0(n1492), .B1(n14), .A0N(memory[534]), .A1N(n14), .Y(
        n2001) );
  OAI2BB2X1 U927 ( .B0(n1490), .B1(n14), .A0N(memory[535]), .A1N(n14), .Y(
        n2000) );
  OAI2BB2X1 U928 ( .B0(n1480), .B1(n14), .A0N(memory[540]), .A1N(n14), .Y(
        n1995) );
  OAI2BB2X1 U929 ( .B0(n1478), .B1(n14), .A0N(memory[541]), .A1N(n14), .Y(
        n1994) );
  OAI2BB2X1 U930 ( .B0(n1476), .B1(n14), .A0N(memory[542]), .A1N(n14), .Y(
        n1993) );
  OAI2BB2X1 U931 ( .B0(n1474), .B1(n14), .A0N(memory[543]), .A1N(n14), .Y(
        n1992) );
  OAI2BB2X1 U932 ( .B0(n1505), .B1(n15), .A0N(memory[544]), .A1N(n15), .Y(
        n1991) );
  OAI2BB2X1 U933 ( .B0(n1503), .B1(n15), .A0N(memory[545]), .A1N(n15), .Y(
        n1990) );
  OAI2BB2X1 U934 ( .B0(n1501), .B1(n15), .A0N(memory[546]), .A1N(n15), .Y(
        n1989) );
  OAI2BB2X1 U935 ( .B0(n1499), .B1(n15), .A0N(memory[547]), .A1N(n15), .Y(
        n1988) );
  OAI2BB2X1 U936 ( .B0(n1497), .B1(n15), .A0N(memory[548]), .A1N(n15), .Y(
        n1987) );
  OAI2BB2X1 U937 ( .B0(n1495), .B1(n15), .A0N(memory[549]), .A1N(n15), .Y(
        n1986) );
  OAI2BB2X1 U938 ( .B0(n1493), .B1(n15), .A0N(memory[550]), .A1N(n15), .Y(
        n1985) );
  OAI2BB2X1 U939 ( .B0(n1491), .B1(n15), .A0N(memory[551]), .A1N(n15), .Y(
        n1984) );
  OAI2BB2X1 U940 ( .B0(n1481), .B1(n15), .A0N(memory[556]), .A1N(n15), .Y(
        n1979) );
  OAI2BB2X1 U941 ( .B0(n1479), .B1(n15), .A0N(memory[557]), .A1N(n15), .Y(
        n1978) );
  OAI2BB2X1 U942 ( .B0(n1477), .B1(n15), .A0N(memory[558]), .A1N(n15), .Y(
        n1977) );
  OAI2BB2X1 U943 ( .B0(n1475), .B1(n15), .A0N(memory[559]), .A1N(n15), .Y(
        n1976) );
  OAI2BB2X1 U944 ( .B0(n1504), .B1(n16), .A0N(memory[560]), .A1N(n16), .Y(
        n1975) );
  OAI2BB2X1 U945 ( .B0(n1502), .B1(n16), .A0N(memory[561]), .A1N(n16), .Y(
        n1974) );
  OAI2BB2X1 U946 ( .B0(n1500), .B1(n16), .A0N(memory[562]), .A1N(n16), .Y(
        n1973) );
  OAI2BB2X1 U947 ( .B0(n1498), .B1(n16), .A0N(memory[563]), .A1N(n16), .Y(
        n1972) );
  OAI2BB2X1 U948 ( .B0(n1496), .B1(n16), .A0N(memory[564]), .A1N(n16), .Y(
        n1971) );
  OAI2BB2X1 U949 ( .B0(n1494), .B1(n16), .A0N(memory[565]), .A1N(n16), .Y(
        n1970) );
  OAI2BB2X1 U950 ( .B0(n1492), .B1(n16), .A0N(memory[566]), .A1N(n16), .Y(
        n1969) );
  OAI2BB2X1 U951 ( .B0(n1490), .B1(n16), .A0N(memory[567]), .A1N(n16), .Y(
        n1968) );
  OAI2BB2X1 U952 ( .B0(n1480), .B1(n16), .A0N(memory[572]), .A1N(n16), .Y(
        n1963) );
  OAI2BB2X1 U953 ( .B0(n1478), .B1(n16), .A0N(memory[573]), .A1N(n16), .Y(
        n1962) );
  OAI2BB2X1 U954 ( .B0(n1476), .B1(n16), .A0N(memory[574]), .A1N(n16), .Y(
        n1961) );
  OAI2BB2X1 U955 ( .B0(n1474), .B1(n16), .A0N(memory[575]), .A1N(n16), .Y(
        n1960) );
  OAI2BB2X1 U956 ( .B0(n1505), .B1(n17), .A0N(memory[576]), .A1N(n17), .Y(
        n1959) );
  OAI2BB2X1 U957 ( .B0(n1503), .B1(n17), .A0N(memory[577]), .A1N(n17), .Y(
        n1958) );
  OAI2BB2X1 U958 ( .B0(n1501), .B1(n17), .A0N(memory[578]), .A1N(n17), .Y(
        n1957) );
  OAI2BB2X1 U959 ( .B0(n1499), .B1(n17), .A0N(memory[579]), .A1N(n17), .Y(
        n1956) );
  OAI2BB2X1 U960 ( .B0(n1497), .B1(n17), .A0N(memory[580]), .A1N(n17), .Y(
        n1955) );
  OAI2BB2X1 U961 ( .B0(n1495), .B1(n17), .A0N(memory[581]), .A1N(n17), .Y(
        n1954) );
  OAI2BB2X1 U962 ( .B0(n1493), .B1(n17), .A0N(memory[582]), .A1N(n17), .Y(
        n1953) );
  OAI2BB2X1 U963 ( .B0(n1491), .B1(n17), .A0N(memory[583]), .A1N(n17), .Y(
        n1952) );
  OAI2BB2X1 U964 ( .B0(n1481), .B1(n17), .A0N(memory[588]), .A1N(n17), .Y(
        n1947) );
  OAI2BB2X1 U965 ( .B0(n1479), .B1(n17), .A0N(memory[589]), .A1N(n17), .Y(
        n1946) );
  OAI2BB2X1 U966 ( .B0(n1477), .B1(n17), .A0N(memory[590]), .A1N(n17), .Y(
        n1945) );
  OAI2BB2X1 U967 ( .B0(n1475), .B1(n17), .A0N(memory[591]), .A1N(n17), .Y(
        n1944) );
  OAI2BB2X1 U968 ( .B0(n1504), .B1(n18), .A0N(memory[592]), .A1N(n18), .Y(
        n1943) );
  OAI2BB2X1 U969 ( .B0(n1502), .B1(n18), .A0N(memory[593]), .A1N(n18), .Y(
        n1942) );
  OAI2BB2X1 U970 ( .B0(n1500), .B1(n18), .A0N(memory[594]), .A1N(n18), .Y(
        n1941) );
  OAI2BB2X1 U971 ( .B0(n1498), .B1(n18), .A0N(memory[595]), .A1N(n18), .Y(
        n1940) );
  OAI2BB2X1 U972 ( .B0(n1496), .B1(n18), .A0N(memory[596]), .A1N(n18), .Y(
        n1939) );
  OAI2BB2X1 U973 ( .B0(n1494), .B1(n18), .A0N(memory[597]), .A1N(n18), .Y(
        n1938) );
  OAI2BB2X1 U974 ( .B0(n1492), .B1(n18), .A0N(memory[598]), .A1N(n18), .Y(
        n1937) );
  OAI2BB2X1 U975 ( .B0(n1490), .B1(n18), .A0N(memory[599]), .A1N(n18), .Y(
        n1936) );
  OAI2BB2X1 U976 ( .B0(n1480), .B1(n18), .A0N(memory[604]), .A1N(n18), .Y(
        n1931) );
  OAI2BB2X1 U977 ( .B0(n1478), .B1(n18), .A0N(memory[605]), .A1N(n18), .Y(
        n1930) );
  OAI2BB2X1 U978 ( .B0(n1476), .B1(n18), .A0N(memory[606]), .A1N(n18), .Y(
        n1929) );
  OAI2BB2X1 U979 ( .B0(n1474), .B1(n18), .A0N(memory[607]), .A1N(n18), .Y(
        n1928) );
  OAI2BB2X1 U980 ( .B0(n1504), .B1(n19), .A0N(memory[608]), .A1N(n19), .Y(
        n1927) );
  OAI2BB2X1 U981 ( .B0(n1502), .B1(n19), .A0N(memory[609]), .A1N(n19), .Y(
        n1926) );
  OAI2BB2X1 U982 ( .B0(n1500), .B1(n19), .A0N(memory[610]), .A1N(n19), .Y(
        n1925) );
  OAI2BB2X1 U983 ( .B0(n1498), .B1(n19), .A0N(memory[611]), .A1N(n19), .Y(
        n1924) );
  OAI2BB2X1 U984 ( .B0(n1496), .B1(n19), .A0N(memory[612]), .A1N(n19), .Y(
        n1923) );
  OAI2BB2X1 U985 ( .B0(n1494), .B1(n19), .A0N(memory[613]), .A1N(n19), .Y(
        n1922) );
  OAI2BB2X1 U986 ( .B0(n1492), .B1(n19), .A0N(memory[614]), .A1N(n19), .Y(
        n1921) );
  OAI2BB2X1 U987 ( .B0(n1490), .B1(n19), .A0N(memory[615]), .A1N(n19), .Y(
        n1920) );
  OAI2BB2X1 U988 ( .B0(n1480), .B1(n19), .A0N(memory[620]), .A1N(n19), .Y(
        n1915) );
  OAI2BB2X1 U989 ( .B0(n1478), .B1(n19), .A0N(memory[621]), .A1N(n19), .Y(
        n1914) );
  OAI2BB2X1 U990 ( .B0(n1476), .B1(n19), .A0N(memory[622]), .A1N(n19), .Y(
        n1913) );
  OAI2BB2X1 U991 ( .B0(n1474), .B1(n19), .A0N(memory[623]), .A1N(n19), .Y(
        n1912) );
  OAI2BB2X1 U992 ( .B0(n1505), .B1(n20), .A0N(memory[624]), .A1N(n20), .Y(
        n1911) );
  OAI2BB2X1 U993 ( .B0(n1503), .B1(n20), .A0N(memory[625]), .A1N(n20), .Y(
        n1910) );
  OAI2BB2X1 U994 ( .B0(n1501), .B1(n20), .A0N(memory[626]), .A1N(n20), .Y(
        n1909) );
  OAI2BB2X1 U995 ( .B0(n1499), .B1(n20), .A0N(memory[627]), .A1N(n20), .Y(
        n1908) );
  OAI2BB2X1 U996 ( .B0(n1497), .B1(n20), .A0N(memory[628]), .A1N(n20), .Y(
        n1907) );
  OAI2BB2X1 U997 ( .B0(n1495), .B1(n20), .A0N(memory[629]), .A1N(n20), .Y(
        n1906) );
  OAI2BB2X1 U998 ( .B0(n1493), .B1(n20), .A0N(memory[630]), .A1N(n20), .Y(
        n1905) );
  OAI2BB2X1 U999 ( .B0(n1491), .B1(n20), .A0N(memory[631]), .A1N(n20), .Y(
        n1904) );
  OAI2BB2X1 U1000 ( .B0(n1481), .B1(n20), .A0N(memory[636]), .A1N(n20), .Y(
        n1899) );
  OAI2BB2X1 U1001 ( .B0(n1479), .B1(n20), .A0N(memory[637]), .A1N(n20), .Y(
        n1898) );
  OAI2BB2X1 U1002 ( .B0(n1477), .B1(n20), .A0N(memory[638]), .A1N(n20), .Y(
        n1897) );
  OAI2BB2X1 U1003 ( .B0(n1475), .B1(n20), .A0N(memory[639]), .A1N(n20), .Y(
        n1896) );
  OAI2BB2X1 U1004 ( .B0(n1504), .B1(n21), .A0N(memory[640]), .A1N(n21), .Y(
        n1895) );
  OAI2BB2X1 U1005 ( .B0(n1502), .B1(n21), .A0N(memory[641]), .A1N(n21), .Y(
        n1894) );
  OAI2BB2X1 U1006 ( .B0(n1500), .B1(n21), .A0N(memory[642]), .A1N(n21), .Y(
        n1893) );
  OAI2BB2X1 U1007 ( .B0(n1498), .B1(n21), .A0N(memory[643]), .A1N(n21), .Y(
        n1892) );
  OAI2BB2X1 U1008 ( .B0(n1496), .B1(n21), .A0N(memory[644]), .A1N(n21), .Y(
        n1891) );
  OAI2BB2X1 U1009 ( .B0(n1494), .B1(n21), .A0N(memory[645]), .A1N(n21), .Y(
        n1890) );
  OAI2BB2X1 U1010 ( .B0(n1492), .B1(n21), .A0N(memory[646]), .A1N(n21), .Y(
        n1889) );
  OAI2BB2X1 U1011 ( .B0(n1490), .B1(n21), .A0N(memory[647]), .A1N(n21), .Y(
        n1888) );
  OAI2BB2X1 U1012 ( .B0(n1480), .B1(n21), .A0N(memory[652]), .A1N(n21), .Y(
        n1883) );
  OAI2BB2X1 U1013 ( .B0(n1478), .B1(n21), .A0N(memory[653]), .A1N(n21), .Y(
        n1882) );
  OAI2BB2X1 U1014 ( .B0(n1476), .B1(n21), .A0N(memory[654]), .A1N(n21), .Y(
        n1881) );
  OAI2BB2X1 U1015 ( .B0(n1474), .B1(n21), .A0N(memory[655]), .A1N(n21), .Y(
        n1880) );
  OAI2BB2X1 U1016 ( .B0(n1504), .B1(n22), .A0N(memory[656]), .A1N(n22), .Y(
        n1879) );
  OAI2BB2X1 U1017 ( .B0(n1502), .B1(n22), .A0N(memory[657]), .A1N(n22), .Y(
        n1878) );
  OAI2BB2X1 U1018 ( .B0(n1500), .B1(n22), .A0N(memory[658]), .A1N(n22), .Y(
        n1877) );
  OAI2BB2X1 U1019 ( .B0(n1498), .B1(n22), .A0N(memory[659]), .A1N(n22), .Y(
        n1876) );
  OAI2BB2X1 U1020 ( .B0(n1496), .B1(n22), .A0N(memory[660]), .A1N(n22), .Y(
        n1875) );
  OAI2BB2X1 U1021 ( .B0(n1494), .B1(n22), .A0N(memory[661]), .A1N(n22), .Y(
        n1874) );
  OAI2BB2X1 U1022 ( .B0(n1492), .B1(n22), .A0N(memory[662]), .A1N(n22), .Y(
        n1873) );
  OAI2BB2X1 U1023 ( .B0(n1490), .B1(n22), .A0N(memory[663]), .A1N(n22), .Y(
        n1872) );
  OAI2BB2X1 U1024 ( .B0(n1480), .B1(n22), .A0N(memory[668]), .A1N(n22), .Y(
        n1867) );
  OAI2BB2X1 U1025 ( .B0(n1478), .B1(n22), .A0N(memory[669]), .A1N(n22), .Y(
        n1866) );
  OAI2BB2X1 U1026 ( .B0(n1476), .B1(n22), .A0N(memory[670]), .A1N(n22), .Y(
        n1865) );
  OAI2BB2X1 U1027 ( .B0(n1474), .B1(n22), .A0N(memory[671]), .A1N(n22), .Y(
        n1864) );
  OAI2BB2X1 U1028 ( .B0(n1505), .B1(n25), .A0N(memory[672]), .A1N(n25), .Y(
        n1863) );
  OAI2BB2X1 U1029 ( .B0(n1503), .B1(n25), .A0N(memory[673]), .A1N(n25), .Y(
        n1862) );
  OAI2BB2X1 U1030 ( .B0(n1501), .B1(n25), .A0N(memory[674]), .A1N(n25), .Y(
        n1861) );
  OAI2BB2X1 U1031 ( .B0(n1499), .B1(n25), .A0N(memory[675]), .A1N(n25), .Y(
        n1860) );
  OAI2BB2X1 U1032 ( .B0(n1497), .B1(n25), .A0N(memory[676]), .A1N(n25), .Y(
        n1859) );
  OAI2BB2X1 U1033 ( .B0(n1495), .B1(n25), .A0N(memory[677]), .A1N(n25), .Y(
        n1858) );
  OAI2BB2X1 U1034 ( .B0(n1493), .B1(n25), .A0N(memory[678]), .A1N(n25), .Y(
        n1857) );
  OAI2BB2X1 U1035 ( .B0(n1491), .B1(n25), .A0N(memory[679]), .A1N(n25), .Y(
        n1856) );
  OAI2BB2X1 U1036 ( .B0(n1481), .B1(n25), .A0N(memory[684]), .A1N(n25), .Y(
        n1851) );
  OAI2BB2X1 U1037 ( .B0(n1479), .B1(n25), .A0N(memory[685]), .A1N(n25), .Y(
        n1850) );
  OAI2BB2X1 U1038 ( .B0(n1477), .B1(n25), .A0N(memory[686]), .A1N(n25), .Y(
        n1849) );
  OAI2BB2X1 U1039 ( .B0(n1475), .B1(n25), .A0N(memory[687]), .A1N(n25), .Y(
        n1848) );
  OAI2BB2X1 U1040 ( .B0(n1504), .B1(n27), .A0N(memory[688]), .A1N(n27), .Y(
        n1847) );
  OAI2BB2X1 U1041 ( .B0(n1502), .B1(n27), .A0N(memory[689]), .A1N(n27), .Y(
        n1846) );
  OAI2BB2X1 U1042 ( .B0(n1500), .B1(n27), .A0N(memory[690]), .A1N(n27), .Y(
        n1845) );
  OAI2BB2X1 U1043 ( .B0(n1498), .B1(n27), .A0N(memory[691]), .A1N(n27), .Y(
        n1844) );
  OAI2BB2X1 U1044 ( .B0(n1496), .B1(n27), .A0N(memory[692]), .A1N(n27), .Y(
        n1843) );
  OAI2BB2X1 U1045 ( .B0(n1494), .B1(n27), .A0N(memory[693]), .A1N(n27), .Y(
        n1842) );
  OAI2BB2X1 U1046 ( .B0(n1492), .B1(n27), .A0N(memory[694]), .A1N(n27), .Y(
        n1841) );
  OAI2BB2X1 U1047 ( .B0(n1490), .B1(n27), .A0N(memory[695]), .A1N(n27), .Y(
        n1840) );
  OAI2BB2X1 U1048 ( .B0(n1480), .B1(n27), .A0N(memory[700]), .A1N(n27), .Y(
        n1835) );
  OAI2BB2X1 U1049 ( .B0(n1478), .B1(n27), .A0N(memory[701]), .A1N(n27), .Y(
        n1834) );
  OAI2BB2X1 U1050 ( .B0(n1476), .B1(n27), .A0N(memory[702]), .A1N(n27), .Y(
        n1833) );
  OAI2BB2X1 U1051 ( .B0(n1474), .B1(n27), .A0N(memory[703]), .A1N(n27), .Y(
        n1832) );
  OAI2BB2X1 U1052 ( .B0(n1505), .B1(n29), .A0N(memory[704]), .A1N(n29), .Y(
        n1831) );
  OAI2BB2X1 U1053 ( .B0(n1503), .B1(n29), .A0N(memory[705]), .A1N(n29), .Y(
        n1830) );
  OAI2BB2X1 U1054 ( .B0(n1501), .B1(n29), .A0N(memory[706]), .A1N(n29), .Y(
        n1829) );
  OAI2BB2X1 U1055 ( .B0(n1499), .B1(n29), .A0N(memory[707]), .A1N(n29), .Y(
        n1828) );
  OAI2BB2X1 U1056 ( .B0(n1497), .B1(n29), .A0N(memory[708]), .A1N(n29), .Y(
        n1827) );
  OAI2BB2X1 U1057 ( .B0(n1495), .B1(n29), .A0N(memory[709]), .A1N(n29), .Y(
        n1826) );
  OAI2BB2X1 U1058 ( .B0(n1493), .B1(n29), .A0N(memory[710]), .A1N(n29), .Y(
        n1825) );
  OAI2BB2X1 U1059 ( .B0(n1491), .B1(n29), .A0N(memory[711]), .A1N(n29), .Y(
        n1824) );
  OAI2BB2X1 U1060 ( .B0(n1481), .B1(n29), .A0N(memory[716]), .A1N(n29), .Y(
        n1819) );
  OAI2BB2X1 U1061 ( .B0(n1479), .B1(n29), .A0N(memory[717]), .A1N(n29), .Y(
        n1818) );
  OAI2BB2X1 U1062 ( .B0(n1477), .B1(n29), .A0N(memory[718]), .A1N(n29), .Y(
        n1817) );
  OAI2BB2X1 U1063 ( .B0(n1475), .B1(n29), .A0N(memory[719]), .A1N(n29), .Y(
        n1816) );
  OAI2BB2X1 U1064 ( .B0(n1504), .B1(n31), .A0N(memory[720]), .A1N(n31), .Y(
        n1815) );
  OAI2BB2X1 U1065 ( .B0(n1502), .B1(n31), .A0N(memory[721]), .A1N(n31), .Y(
        n1814) );
  OAI2BB2X1 U1066 ( .B0(n1500), .B1(n31), .A0N(memory[722]), .A1N(n31), .Y(
        n1813) );
  OAI2BB2X1 U1067 ( .B0(n1498), .B1(n31), .A0N(memory[723]), .A1N(n31), .Y(
        n1812) );
  OAI2BB2X1 U1068 ( .B0(n1496), .B1(n31), .A0N(memory[724]), .A1N(n31), .Y(
        n1811) );
  OAI2BB2X1 U1069 ( .B0(n1494), .B1(n31), .A0N(memory[725]), .A1N(n31), .Y(
        n1810) );
  OAI2BB2X1 U1070 ( .B0(n1492), .B1(n31), .A0N(memory[726]), .A1N(n31), .Y(
        n1809) );
  OAI2BB2X1 U1071 ( .B0(n1490), .B1(n31), .A0N(memory[727]), .A1N(n31), .Y(
        n1808) );
  OAI2BB2X1 U1072 ( .B0(n1480), .B1(n31), .A0N(memory[732]), .A1N(n31), .Y(
        n1803) );
  OAI2BB2X1 U1073 ( .B0(n1478), .B1(n31), .A0N(memory[733]), .A1N(n31), .Y(
        n1802) );
  OAI2BB2X1 U1074 ( .B0(n1476), .B1(n31), .A0N(memory[734]), .A1N(n31), .Y(
        n1801) );
  OAI2BB2X1 U1075 ( .B0(n1474), .B1(n31), .A0N(memory[735]), .A1N(n31), .Y(
        n1800) );
  OAI2BB2X1 U1076 ( .B0(n1505), .B1(n33), .A0N(memory[736]), .A1N(n33), .Y(
        n1799) );
  OAI2BB2X1 U1077 ( .B0(n1503), .B1(n33), .A0N(memory[737]), .A1N(n33), .Y(
        n1798) );
  OAI2BB2X1 U1078 ( .B0(n1501), .B1(n33), .A0N(memory[738]), .A1N(n33), .Y(
        n1797) );
  OAI2BB2X1 U1079 ( .B0(n1499), .B1(n33), .A0N(memory[739]), .A1N(n33), .Y(
        n1796) );
  OAI2BB2X1 U1080 ( .B0(n1497), .B1(n33), .A0N(memory[740]), .A1N(n33), .Y(
        n1795) );
  OAI2BB2X1 U1081 ( .B0(n1495), .B1(n33), .A0N(memory[741]), .A1N(n33), .Y(
        n1794) );
  OAI2BB2X1 U1082 ( .B0(n1493), .B1(n33), .A0N(memory[742]), .A1N(n33), .Y(
        n1793) );
  OAI2BB2X1 U1083 ( .B0(n1491), .B1(n33), .A0N(memory[743]), .A1N(n33), .Y(
        n1792) );
  OAI2BB2X1 U1084 ( .B0(n1481), .B1(n33), .A0N(memory[748]), .A1N(n33), .Y(
        n1787) );
  OAI2BB2X1 U1085 ( .B0(n1479), .B1(n33), .A0N(memory[749]), .A1N(n33), .Y(
        n1786) );
  OAI2BB2X1 U1086 ( .B0(n1477), .B1(n33), .A0N(memory[750]), .A1N(n33), .Y(
        n1785) );
  OAI2BB2X1 U1087 ( .B0(n1475), .B1(n33), .A0N(memory[751]), .A1N(n33), .Y(
        n1784) );
  OAI2BB2X1 U1088 ( .B0(n1504), .B1(n35), .A0N(memory[752]), .A1N(n35), .Y(
        n1783) );
  OAI2BB2X1 U1089 ( .B0(n1502), .B1(n35), .A0N(memory[753]), .A1N(n35), .Y(
        n1782) );
  OAI2BB2X1 U1090 ( .B0(n1500), .B1(n35), .A0N(memory[754]), .A1N(n35), .Y(
        n1781) );
  OAI2BB2X1 U1091 ( .B0(n1498), .B1(n35), .A0N(memory[755]), .A1N(n35), .Y(
        n1780) );
  OAI2BB2X1 U1092 ( .B0(n1496), .B1(n35), .A0N(memory[756]), .A1N(n35), .Y(
        n1779) );
  OAI2BB2X1 U1093 ( .B0(n1494), .B1(n35), .A0N(memory[757]), .A1N(n35), .Y(
        n1778) );
  OAI2BB2X1 U1094 ( .B0(n1492), .B1(n35), .A0N(memory[758]), .A1N(n35), .Y(
        n1777) );
  OAI2BB2X1 U1095 ( .B0(n1490), .B1(n35), .A0N(memory[759]), .A1N(n35), .Y(
        n1776) );
  OAI2BB2X1 U1096 ( .B0(n1480), .B1(n35), .A0N(memory[764]), .A1N(n35), .Y(
        n1771) );
  OAI2BB2X1 U1097 ( .B0(n1478), .B1(n35), .A0N(memory[765]), .A1N(n35), .Y(
        n1770) );
  OAI2BB2X1 U1098 ( .B0(n1476), .B1(n35), .A0N(memory[766]), .A1N(n35), .Y(
        n1769) );
  OAI2BB2X1 U1099 ( .B0(n1474), .B1(n35), .A0N(memory[767]), .A1N(n35), .Y(
        n1768) );
  OAI2BB2X1 U1100 ( .B0(n1504), .B1(n37), .A0N(memory[768]), .A1N(n37), .Y(
        n1767) );
  OAI2BB2X1 U1101 ( .B0(n1502), .B1(n37), .A0N(memory[769]), .A1N(n37), .Y(
        n1766) );
  OAI2BB2X1 U1102 ( .B0(n1500), .B1(n37), .A0N(memory[770]), .A1N(n37), .Y(
        n1765) );
  OAI2BB2X1 U1103 ( .B0(n1498), .B1(n37), .A0N(memory[771]), .A1N(n37), .Y(
        n1764) );
  OAI2BB2X1 U1104 ( .B0(n1496), .B1(n37), .A0N(memory[772]), .A1N(n37), .Y(
        n1763) );
  OAI2BB2X1 U1105 ( .B0(n1494), .B1(n37), .A0N(memory[773]), .A1N(n37), .Y(
        n1762) );
  OAI2BB2X1 U1106 ( .B0(n1492), .B1(n37), .A0N(memory[774]), .A1N(n37), .Y(
        n1761) );
  OAI2BB2X1 U1107 ( .B0(n1490), .B1(n37), .A0N(memory[775]), .A1N(n37), .Y(
        n1760) );
  OAI2BB2X1 U1108 ( .B0(n1480), .B1(n37), .A0N(memory[780]), .A1N(n37), .Y(
        n1755) );
  OAI2BB2X1 U1109 ( .B0(n1478), .B1(n37), .A0N(memory[781]), .A1N(n37), .Y(
        n1754) );
  OAI2BB2X1 U1110 ( .B0(n1476), .B1(n37), .A0N(memory[782]), .A1N(n37), .Y(
        n1753) );
  OAI2BB2X1 U1111 ( .B0(n1474), .B1(n37), .A0N(memory[783]), .A1N(n37), .Y(
        n1752) );
  OAI2BB2X1 U1112 ( .B0(n1505), .B1(n40), .A0N(memory[784]), .A1N(n40), .Y(
        n1751) );
  OAI2BB2X1 U1113 ( .B0(n1503), .B1(n40), .A0N(memory[785]), .A1N(n40), .Y(
        n1750) );
  OAI2BB2X1 U1114 ( .B0(n1501), .B1(n40), .A0N(memory[786]), .A1N(n40), .Y(
        n1749) );
  OAI2BB2X1 U1115 ( .B0(n1499), .B1(n40), .A0N(memory[787]), .A1N(n40), .Y(
        n1748) );
  OAI2BB2X1 U1116 ( .B0(n1497), .B1(n40), .A0N(memory[788]), .A1N(n40), .Y(
        n1747) );
  OAI2BB2X1 U1117 ( .B0(n1495), .B1(n40), .A0N(memory[789]), .A1N(n40), .Y(
        n1746) );
  OAI2BB2X1 U1118 ( .B0(n1493), .B1(n40), .A0N(memory[790]), .A1N(n40), .Y(
        n1745) );
  OAI2BB2X1 U1119 ( .B0(n1491), .B1(n40), .A0N(memory[791]), .A1N(n40), .Y(
        n1744) );
  OAI2BB2X1 U1120 ( .B0(n1481), .B1(n40), .A0N(memory[796]), .A1N(n40), .Y(
        n1739) );
  OAI2BB2X1 U1121 ( .B0(n1479), .B1(n40), .A0N(memory[797]), .A1N(n40), .Y(
        n1738) );
  OAI2BB2X1 U1122 ( .B0(n1477), .B1(n40), .A0N(memory[798]), .A1N(n40), .Y(
        n1737) );
  OAI2BB2X1 U1123 ( .B0(n1475), .B1(n40), .A0N(memory[799]), .A1N(n40), .Y(
        n1736) );
  OAI2BB2X1 U1124 ( .B0(n1504), .B1(n42), .A0N(memory[800]), .A1N(n42), .Y(
        n1735) );
  OAI2BB2X1 U1125 ( .B0(n1502), .B1(n42), .A0N(memory[801]), .A1N(n42), .Y(
        n1734) );
  OAI2BB2X1 U1126 ( .B0(n1500), .B1(n42), .A0N(memory[802]), .A1N(n42), .Y(
        n1733) );
  OAI2BB2X1 U1127 ( .B0(n1498), .B1(n42), .A0N(memory[803]), .A1N(n42), .Y(
        n1732) );
  OAI2BB2X1 U1128 ( .B0(n1496), .B1(n42), .A0N(memory[804]), .A1N(n42), .Y(
        n1731) );
  OAI2BB2X1 U1129 ( .B0(n1494), .B1(n42), .A0N(memory[805]), .A1N(n42), .Y(
        n1730) );
  OAI2BB2X1 U1130 ( .B0(n1492), .B1(n42), .A0N(memory[806]), .A1N(n42), .Y(
        n1729) );
  OAI2BB2X1 U1131 ( .B0(n1490), .B1(n42), .A0N(memory[807]), .A1N(n42), .Y(
        n1728) );
  OAI2BB2X1 U1132 ( .B0(n1480), .B1(n42), .A0N(memory[812]), .A1N(n42), .Y(
        n1723) );
  OAI2BB2X1 U1133 ( .B0(n1478), .B1(n42), .A0N(memory[813]), .A1N(n42), .Y(
        n1722) );
  OAI2BB2X1 U1134 ( .B0(n1476), .B1(n42), .A0N(memory[814]), .A1N(n42), .Y(
        n1721) );
  OAI2BB2X1 U1135 ( .B0(n1474), .B1(n42), .A0N(memory[815]), .A1N(n42), .Y(
        n1720) );
  OAI2BB2X1 U1136 ( .B0(n1504), .B1(n43), .A0N(memory[816]), .A1N(n43), .Y(
        n1719) );
  OAI2BB2X1 U1137 ( .B0(n1502), .B1(n43), .A0N(memory[817]), .A1N(n43), .Y(
        n1718) );
  OAI2BB2X1 U1138 ( .B0(n1500), .B1(n43), .A0N(memory[818]), .A1N(n43), .Y(
        n1717) );
  OAI2BB2X1 U1139 ( .B0(n1498), .B1(n43), .A0N(memory[819]), .A1N(n43), .Y(
        n1716) );
  OAI2BB2X1 U1140 ( .B0(n1496), .B1(n43), .A0N(memory[820]), .A1N(n43), .Y(
        n1715) );
  OAI2BB2X1 U1141 ( .B0(n1494), .B1(n43), .A0N(memory[821]), .A1N(n43), .Y(
        n1714) );
  OAI2BB2X1 U1142 ( .B0(n1492), .B1(n43), .A0N(memory[822]), .A1N(n43), .Y(
        n1713) );
  OAI2BB2X1 U1143 ( .B0(n1490), .B1(n43), .A0N(memory[823]), .A1N(n43), .Y(
        n1712) );
  OAI2BB2X1 U1144 ( .B0(n1480), .B1(n43), .A0N(memory[828]), .A1N(n43), .Y(
        n1707) );
  OAI2BB2X1 U1145 ( .B0(n1478), .B1(n43), .A0N(memory[829]), .A1N(n43), .Y(
        n1706) );
  OAI2BB2X1 U1146 ( .B0(n1476), .B1(n43), .A0N(memory[830]), .A1N(n43), .Y(
        n1705) );
  OAI2BB2X1 U1147 ( .B0(n1474), .B1(n43), .A0N(memory[831]), .A1N(n43), .Y(
        n1704) );
  OAI2BB2X1 U1148 ( .B0(n1504), .B1(n44), .A0N(memory[832]), .A1N(n44), .Y(
        n1703) );
  OAI2BB2X1 U1149 ( .B0(n1502), .B1(n44), .A0N(memory[833]), .A1N(n44), .Y(
        n1702) );
  OAI2BB2X1 U1150 ( .B0(n1500), .B1(n44), .A0N(memory[834]), .A1N(n44), .Y(
        n1701) );
  OAI2BB2X1 U1151 ( .B0(n1498), .B1(n44), .A0N(memory[835]), .A1N(n44), .Y(
        n1700) );
  OAI2BB2X1 U1152 ( .B0(n1496), .B1(n44), .A0N(memory[836]), .A1N(n44), .Y(
        n1699) );
  OAI2BB2X1 U1153 ( .B0(n1494), .B1(n44), .A0N(memory[837]), .A1N(n44), .Y(
        n1698) );
  OAI2BB2X1 U1154 ( .B0(n1492), .B1(n44), .A0N(memory[838]), .A1N(n44), .Y(
        n1697) );
  OAI2BB2X1 U1155 ( .B0(n1490), .B1(n44), .A0N(memory[839]), .A1N(n44), .Y(
        n1696) );
  OAI2BB2X1 U1156 ( .B0(n1480), .B1(n44), .A0N(memory[844]), .A1N(n44), .Y(
        n1691) );
  OAI2BB2X1 U1157 ( .B0(n1478), .B1(n44), .A0N(memory[845]), .A1N(n44), .Y(
        n1690) );
  OAI2BB2X1 U1158 ( .B0(n1476), .B1(n44), .A0N(memory[846]), .A1N(n44), .Y(
        n1689) );
  OAI2BB2X1 U1159 ( .B0(n1474), .B1(n44), .A0N(memory[847]), .A1N(n44), .Y(
        n1688) );
  OAI2BB2X1 U1160 ( .B0(n1504), .B1(n45), .A0N(memory[848]), .A1N(n45), .Y(
        n1687) );
  OAI2BB2X1 U1161 ( .B0(n1502), .B1(n45), .A0N(memory[849]), .A1N(n45), .Y(
        n1686) );
  OAI2BB2X1 U1162 ( .B0(n1500), .B1(n45), .A0N(memory[850]), .A1N(n45), .Y(
        n1685) );
  OAI2BB2X1 U1163 ( .B0(n1498), .B1(n45), .A0N(memory[851]), .A1N(n45), .Y(
        n1684) );
  OAI2BB2X1 U1164 ( .B0(n1496), .B1(n45), .A0N(memory[852]), .A1N(n45), .Y(
        n1683) );
  OAI2BB2X1 U1165 ( .B0(n1494), .B1(n45), .A0N(memory[853]), .A1N(n45), .Y(
        n1682) );
  OAI2BB2X1 U1166 ( .B0(n1492), .B1(n45), .A0N(memory[854]), .A1N(n45), .Y(
        n1681) );
  OAI2BB2X1 U1167 ( .B0(n1490), .B1(n45), .A0N(memory[855]), .A1N(n45), .Y(
        n1680) );
  OAI2BB2X1 U1168 ( .B0(n1480), .B1(n45), .A0N(memory[860]), .A1N(n45), .Y(
        n1675) );
  OAI2BB2X1 U1169 ( .B0(n1478), .B1(n45), .A0N(memory[861]), .A1N(n45), .Y(
        n1674) );
  OAI2BB2X1 U1170 ( .B0(n1476), .B1(n45), .A0N(memory[862]), .A1N(n45), .Y(
        n1673) );
  OAI2BB2X1 U1171 ( .B0(n1474), .B1(n45), .A0N(memory[863]), .A1N(n45), .Y(
        n1672) );
  OAI2BB2X1 U1172 ( .B0(n1504), .B1(n46), .A0N(memory[864]), .A1N(n46), .Y(
        n1671) );
  OAI2BB2X1 U1173 ( .B0(n1502), .B1(n46), .A0N(memory[865]), .A1N(n46), .Y(
        n1670) );
  OAI2BB2X1 U1174 ( .B0(n1500), .B1(n46), .A0N(memory[866]), .A1N(n46), .Y(
        n1669) );
  OAI2BB2X1 U1175 ( .B0(n1498), .B1(n46), .A0N(memory[867]), .A1N(n46), .Y(
        n1668) );
  OAI2BB2X1 U1176 ( .B0(n1496), .B1(n46), .A0N(memory[868]), .A1N(n46), .Y(
        n1667) );
  OAI2BB2X1 U1177 ( .B0(n1494), .B1(n46), .A0N(memory[869]), .A1N(n46), .Y(
        n1666) );
  OAI2BB2X1 U1178 ( .B0(n1492), .B1(n46), .A0N(memory[870]), .A1N(n46), .Y(
        n1665) );
  OAI2BB2X1 U1179 ( .B0(n1490), .B1(n46), .A0N(memory[871]), .A1N(n46), .Y(
        n1664) );
  OAI2BB2X1 U1180 ( .B0(n1480), .B1(n46), .A0N(memory[876]), .A1N(n46), .Y(
        n1659) );
  OAI2BB2X1 U1181 ( .B0(n1478), .B1(n46), .A0N(memory[877]), .A1N(n46), .Y(
        n1658) );
  OAI2BB2X1 U1182 ( .B0(n1476), .B1(n46), .A0N(memory[878]), .A1N(n46), .Y(
        n1657) );
  OAI2BB2X1 U1183 ( .B0(n1474), .B1(n46), .A0N(memory[879]), .A1N(n46), .Y(
        n1656) );
  OAI2BB2X1 U1184 ( .B0(n1504), .B1(n47), .A0N(memory[880]), .A1N(n47), .Y(
        n1655) );
  OAI2BB2X1 U1185 ( .B0(n1502), .B1(n47), .A0N(memory[881]), .A1N(n47), .Y(
        n1654) );
  OAI2BB2X1 U1186 ( .B0(n1500), .B1(n47), .A0N(memory[882]), .A1N(n47), .Y(
        n1653) );
  OAI2BB2X1 U1187 ( .B0(n1498), .B1(n47), .A0N(memory[883]), .A1N(n47), .Y(
        n1652) );
  OAI2BB2X1 U1188 ( .B0(n1496), .B1(n47), .A0N(memory[884]), .A1N(n47), .Y(
        n1651) );
  OAI2BB2X1 U1189 ( .B0(n1494), .B1(n47), .A0N(memory[885]), .A1N(n47), .Y(
        n1650) );
  OAI2BB2X1 U1190 ( .B0(n1492), .B1(n47), .A0N(memory[886]), .A1N(n47), .Y(
        n1649) );
  OAI2BB2X1 U1191 ( .B0(n1490), .B1(n47), .A0N(memory[887]), .A1N(n47), .Y(
        n1648) );
  OAI2BB2X1 U1192 ( .B0(n1480), .B1(n47), .A0N(memory[892]), .A1N(n47), .Y(
        n1643) );
  OAI2BB2X1 U1193 ( .B0(n1478), .B1(n47), .A0N(memory[893]), .A1N(n47), .Y(
        n1642) );
  OAI2BB2X1 U1194 ( .B0(n1476), .B1(n47), .A0N(memory[894]), .A1N(n47), .Y(
        n1641) );
  OAI2BB2X1 U1195 ( .B0(n1474), .B1(n47), .A0N(memory[895]), .A1N(n47), .Y(
        n1640) );
  OAI2BB2X1 U1196 ( .B0(n1504), .B1(n48), .A0N(memory[896]), .A1N(n48), .Y(
        n1639) );
  OAI2BB2X1 U1197 ( .B0(n1502), .B1(n48), .A0N(memory[897]), .A1N(n48), .Y(
        n1638) );
  OAI2BB2X1 U1198 ( .B0(n1500), .B1(n48), .A0N(memory[898]), .A1N(n48), .Y(
        n1637) );
  OAI2BB2X1 U1199 ( .B0(n1498), .B1(n48), .A0N(memory[899]), .A1N(n48), .Y(
        n1636) );
  OAI2BB2X1 U1200 ( .B0(n1496), .B1(n48), .A0N(memory[900]), .A1N(n48), .Y(
        n1635) );
  OAI2BB2X1 U1201 ( .B0(n1494), .B1(n48), .A0N(memory[901]), .A1N(n48), .Y(
        n1634) );
  OAI2BB2X1 U1202 ( .B0(n1492), .B1(n48), .A0N(memory[902]), .A1N(n48), .Y(
        n1633) );
  OAI2BB2X1 U1203 ( .B0(n1490), .B1(n48), .A0N(memory[903]), .A1N(n48), .Y(
        n1632) );
  OAI2BB2X1 U1204 ( .B0(n1480), .B1(n48), .A0N(memory[908]), .A1N(n48), .Y(
        n1627) );
  OAI2BB2X1 U1205 ( .B0(n1478), .B1(n48), .A0N(memory[909]), .A1N(n48), .Y(
        n1626) );
  OAI2BB2X1 U1206 ( .B0(n1476), .B1(n48), .A0N(memory[910]), .A1N(n48), .Y(
        n1625) );
  OAI2BB2X1 U1207 ( .B0(n1474), .B1(n48), .A0N(memory[911]), .A1N(n48), .Y(
        n1624) );
  OAI2BB2X1 U1208 ( .B0(n1504), .B1(n49), .A0N(memory[912]), .A1N(n49), .Y(
        n1623) );
  OAI2BB2X1 U1209 ( .B0(n1502), .B1(n49), .A0N(memory[913]), .A1N(n49), .Y(
        n1622) );
  OAI2BB2X1 U1210 ( .B0(n1500), .B1(n49), .A0N(memory[914]), .A1N(n49), .Y(
        n1621) );
  OAI2BB2X1 U1211 ( .B0(n1498), .B1(n49), .A0N(memory[915]), .A1N(n49), .Y(
        n1620) );
  OAI2BB2X1 U1212 ( .B0(n1496), .B1(n49), .A0N(memory[916]), .A1N(n49), .Y(
        n1619) );
  OAI2BB2X1 U1213 ( .B0(n1494), .B1(n49), .A0N(memory[917]), .A1N(n49), .Y(
        n1618) );
  OAI2BB2X1 U1214 ( .B0(n1492), .B1(n49), .A0N(memory[918]), .A1N(n49), .Y(
        n1617) );
  OAI2BB2X1 U1215 ( .B0(n1490), .B1(n49), .A0N(memory[919]), .A1N(n49), .Y(
        n1616) );
  OAI2BB2X1 U1216 ( .B0(n1480), .B1(n49), .A0N(memory[924]), .A1N(n49), .Y(
        n1611) );
  OAI2BB2X1 U1217 ( .B0(n1478), .B1(n49), .A0N(memory[925]), .A1N(n49), .Y(
        n1610) );
  OAI2BB2X1 U1218 ( .B0(n1476), .B1(n49), .A0N(memory[926]), .A1N(n49), .Y(
        n1609) );
  OAI2BB2X1 U1219 ( .B0(n1474), .B1(n49), .A0N(memory[927]), .A1N(n49), .Y(
        n1608) );
  OAI2BB2X1 U1220 ( .B0(n1504), .B1(n51), .A0N(memory[928]), .A1N(n51), .Y(
        n1607) );
  OAI2BB2X1 U1221 ( .B0(n1502), .B1(n51), .A0N(memory[929]), .A1N(n51), .Y(
        n1606) );
  OAI2BB2X1 U1222 ( .B0(n1500), .B1(n51), .A0N(memory[930]), .A1N(n51), .Y(
        n1605) );
  OAI2BB2X1 U1223 ( .B0(n1498), .B1(n51), .A0N(memory[931]), .A1N(n51), .Y(
        n1604) );
  OAI2BB2X1 U1224 ( .B0(n1496), .B1(n51), .A0N(memory[932]), .A1N(n51), .Y(
        n1603) );
  OAI2BB2X1 U1225 ( .B0(n1494), .B1(n51), .A0N(memory[933]), .A1N(n51), .Y(
        n1602) );
  OAI2BB2X1 U1226 ( .B0(n1492), .B1(n51), .A0N(memory[934]), .A1N(n51), .Y(
        n1601) );
  OAI2BB2X1 U1227 ( .B0(n1490), .B1(n51), .A0N(memory[935]), .A1N(n51), .Y(
        n1600) );
  OAI2BB2X1 U1228 ( .B0(n1480), .B1(n51), .A0N(memory[940]), .A1N(n51), .Y(
        n1595) );
  OAI2BB2X1 U1229 ( .B0(n1478), .B1(n51), .A0N(memory[941]), .A1N(n51), .Y(
        n1594) );
  OAI2BB2X1 U1230 ( .B0(n1476), .B1(n51), .A0N(memory[942]), .A1N(n51), .Y(
        n1593) );
  OAI2BB2X1 U1231 ( .B0(n1474), .B1(n51), .A0N(memory[943]), .A1N(n51), .Y(
        n1592) );
  OAI2BB2X1 U1232 ( .B0(n1504), .B1(n52), .A0N(memory[944]), .A1N(n52), .Y(
        n1591) );
  OAI2BB2X1 U1233 ( .B0(n1502), .B1(n52), .A0N(memory[945]), .A1N(n52), .Y(
        n1590) );
  OAI2BB2X1 U1234 ( .B0(n1500), .B1(n52), .A0N(memory[946]), .A1N(n52), .Y(
        n1589) );
  OAI2BB2X1 U1235 ( .B0(n1498), .B1(n52), .A0N(memory[947]), .A1N(n52), .Y(
        n1588) );
  OAI2BB2X1 U1236 ( .B0(n1496), .B1(n52), .A0N(memory[948]), .A1N(n52), .Y(
        n1587) );
  OAI2BB2X1 U1237 ( .B0(n1494), .B1(n52), .A0N(memory[949]), .A1N(n52), .Y(
        n1586) );
  OAI2BB2X1 U1238 ( .B0(n1492), .B1(n52), .A0N(memory[950]), .A1N(n52), .Y(
        n1585) );
  OAI2BB2X1 U1239 ( .B0(n1490), .B1(n52), .A0N(memory[951]), .A1N(n52), .Y(
        n1584) );
  OAI2BB2X1 U1240 ( .B0(n1480), .B1(n52), .A0N(memory[956]), .A1N(n52), .Y(
        n1579) );
  OAI2BB2X1 U1241 ( .B0(n1478), .B1(n52), .A0N(memory[957]), .A1N(n52), .Y(
        n1578) );
  OAI2BB2X1 U1242 ( .B0(n1476), .B1(n52), .A0N(memory[958]), .A1N(n52), .Y(
        n1577) );
  OAI2BB2X1 U1243 ( .B0(n1474), .B1(n52), .A0N(memory[959]), .A1N(n52), .Y(
        n1576) );
  OAI2BB2X1 U1244 ( .B0(n1504), .B1(n53), .A0N(memory[960]), .A1N(n53), .Y(
        n1575) );
  OAI2BB2X1 U1245 ( .B0(n1502), .B1(n53), .A0N(memory[961]), .A1N(n53), .Y(
        n1574) );
  OAI2BB2X1 U1246 ( .B0(n1500), .B1(n53), .A0N(memory[962]), .A1N(n53), .Y(
        n1573) );
  OAI2BB2X1 U1247 ( .B0(n1498), .B1(n53), .A0N(memory[963]), .A1N(n53), .Y(
        n1572) );
  OAI2BB2X1 U1248 ( .B0(n1496), .B1(n53), .A0N(memory[964]), .A1N(n53), .Y(
        n1571) );
  OAI2BB2X1 U1249 ( .B0(n1494), .B1(n53), .A0N(memory[965]), .A1N(n53), .Y(
        n1570) );
  OAI2BB2X1 U1250 ( .B0(n1492), .B1(n53), .A0N(memory[966]), .A1N(n53), .Y(
        n1569) );
  OAI2BB2X1 U1251 ( .B0(n1490), .B1(n53), .A0N(memory[967]), .A1N(n53), .Y(
        n1568) );
  OAI2BB2X1 U1252 ( .B0(n1480), .B1(n53), .A0N(memory[972]), .A1N(n53), .Y(
        n1563) );
  OAI2BB2X1 U1253 ( .B0(n1478), .B1(n53), .A0N(memory[973]), .A1N(n53), .Y(
        n1562) );
  OAI2BB2X1 U1254 ( .B0(n1476), .B1(n53), .A0N(memory[974]), .A1N(n53), .Y(
        n1561) );
  OAI2BB2X1 U1255 ( .B0(n1474), .B1(n53), .A0N(memory[975]), .A1N(n53), .Y(
        n1560) );
  OAI2BB2X1 U1256 ( .B0(n1504), .B1(n54), .A0N(memory[976]), .A1N(n54), .Y(
        n1559) );
  OAI2BB2X1 U1257 ( .B0(n1502), .B1(n54), .A0N(memory[977]), .A1N(n54), .Y(
        n1558) );
  OAI2BB2X1 U1258 ( .B0(n1500), .B1(n54), .A0N(memory[978]), .A1N(n54), .Y(
        n1557) );
  OAI2BB2X1 U1259 ( .B0(n1498), .B1(n54), .A0N(memory[979]), .A1N(n54), .Y(
        n1556) );
  OAI2BB2X1 U1260 ( .B0(n1496), .B1(n54), .A0N(memory[980]), .A1N(n54), .Y(
        n1555) );
  OAI2BB2X1 U1261 ( .B0(n1494), .B1(n54), .A0N(memory[981]), .A1N(n54), .Y(
        n1554) );
  OAI2BB2X1 U1262 ( .B0(n1492), .B1(n54), .A0N(memory[982]), .A1N(n54), .Y(
        n1553) );
  OAI2BB2X1 U1263 ( .B0(n1490), .B1(n54), .A0N(memory[983]), .A1N(n54), .Y(
        n1552) );
  OAI2BB2X1 U1264 ( .B0(n1480), .B1(n54), .A0N(memory[988]), .A1N(n54), .Y(
        n1547) );
  OAI2BB2X1 U1265 ( .B0(n1478), .B1(n54), .A0N(memory[989]), .A1N(n54), .Y(
        n1546) );
  OAI2BB2X1 U1266 ( .B0(n1476), .B1(n54), .A0N(memory[990]), .A1N(n54), .Y(
        n1545) );
  OAI2BB2X1 U1267 ( .B0(n1474), .B1(n54), .A0N(memory[991]), .A1N(n54), .Y(
        n1544) );
  OAI2BB2X1 U1268 ( .B0(n1504), .B1(n55), .A0N(memory[992]), .A1N(n55), .Y(
        n1543) );
  OAI2BB2X1 U1269 ( .B0(n1502), .B1(n55), .A0N(memory[993]), .A1N(n55), .Y(
        n1542) );
  OAI2BB2X1 U1270 ( .B0(n1500), .B1(n55), .A0N(memory[994]), .A1N(n55), .Y(
        n1541) );
  OAI2BB2X1 U1271 ( .B0(n1498), .B1(n55), .A0N(memory[995]), .A1N(n55), .Y(
        n1540) );
  OAI2BB2X1 U1272 ( .B0(n1496), .B1(n55), .A0N(memory[996]), .A1N(n55), .Y(
        n1539) );
  OAI2BB2X1 U1273 ( .B0(n1494), .B1(n55), .A0N(memory[997]), .A1N(n55), .Y(
        n1538) );
  OAI2BB2X1 U1274 ( .B0(n1492), .B1(n55), .A0N(memory[998]), .A1N(n55), .Y(
        n1537) );
  OAI2BB2X1 U1275 ( .B0(n1490), .B1(n55), .A0N(memory[999]), .A1N(n55), .Y(
        n1536) );
  OAI2BB2X1 U1276 ( .B0(n1480), .B1(n55), .A0N(memory[1004]), .A1N(n55), .Y(
        n1531) );
  OAI2BB2X1 U1277 ( .B0(n1478), .B1(n55), .A0N(memory[1005]), .A1N(n55), .Y(
        n1530) );
  OAI2BB2X1 U1278 ( .B0(n1476), .B1(n55), .A0N(memory[1006]), .A1N(n55), .Y(
        n1529) );
  OAI2BB2X1 U1279 ( .B0(n1474), .B1(n55), .A0N(memory[1007]), .A1N(n55), .Y(
        n1528) );
  OAI2BB2X1 U1280 ( .B0(n1504), .B1(n56), .A0N(memory[1008]), .A1N(n56), .Y(
        n1527) );
  OAI2BB2X1 U1281 ( .B0(n1502), .B1(n56), .A0N(memory[1009]), .A1N(n56), .Y(
        n1526) );
  OAI2BB2X1 U1282 ( .B0(n1500), .B1(n56), .A0N(memory[1010]), .A1N(n56), .Y(
        n1525) );
  OAI2BB2X1 U1283 ( .B0(n1498), .B1(n56), .A0N(memory[1011]), .A1N(n56), .Y(
        n1524) );
  OAI2BB2X1 U1284 ( .B0(n1496), .B1(n56), .A0N(memory[1012]), .A1N(n56), .Y(
        n1523) );
  OAI2BB2X1 U1285 ( .B0(n1494), .B1(n56), .A0N(memory[1013]), .A1N(n56), .Y(
        n1522) );
  OAI2BB2X1 U1286 ( .B0(n1492), .B1(n56), .A0N(memory[1014]), .A1N(n56), .Y(
        n1521) );
  OAI2BB2X1 U1287 ( .B0(n1490), .B1(n56), .A0N(memory[1015]), .A1N(n56), .Y(
        n1520) );
  OAI2BB2X1 U1288 ( .B0(n1480), .B1(n56), .A0N(memory[1020]), .A1N(n56), .Y(
        n1515) );
  OAI2BB2X1 U1289 ( .B0(n1478), .B1(n56), .A0N(memory[1021]), .A1N(n56), .Y(
        n1514) );
  OAI2BB2X1 U1290 ( .B0(n1476), .B1(n56), .A0N(memory[1022]), .A1N(n56), .Y(
        n1513) );
  OAI2BB2X1 U1291 ( .B0(n1474), .B1(n56), .A0N(memory[1023]), .A1N(n56), .Y(
        n1512) );
  OAI2BB2X1 U1292 ( .B0(n1488), .B1(n2), .A0N(memory[24]), .A1N(n2), .Y(n2511)
         );
  OAI2BB2X1 U1293 ( .B0(n1486), .B1(n2), .A0N(memory[25]), .A1N(n2), .Y(n2510)
         );
  OAI2BB2X1 U1294 ( .B0(n1484), .B1(n2), .A0N(memory[26]), .A1N(n2), .Y(n2509)
         );
  OAI2BB2X1 U1295 ( .B0(n1482), .B1(n2), .A0N(memory[27]), .A1N(n2), .Y(n2508)
         );
  OAI2BB2X1 U1296 ( .B0(n1488), .B1(n57), .A0N(memory[40]), .A1N(n57), .Y(
        n2495) );
  OAI2BB2X1 U1297 ( .B0(n1486), .B1(n57), .A0N(memory[41]), .A1N(n57), .Y(
        n2494) );
  OAI2BB2X1 U1298 ( .B0(n1484), .B1(n57), .A0N(memory[42]), .A1N(n57), .Y(
        n2493) );
  OAI2BB2X1 U1299 ( .B0(n1482), .B1(n57), .A0N(memory[43]), .A1N(n57), .Y(
        n2492) );
  OAI2BB2X1 U1300 ( .B0(n1489), .B1(n58), .A0N(memory[56]), .A1N(n58), .Y(
        n2479) );
  OAI2BB2X1 U1301 ( .B0(n1487), .B1(n58), .A0N(memory[57]), .A1N(n58), .Y(
        n2478) );
  OAI2BB2X1 U1302 ( .B0(n1485), .B1(n58), .A0N(memory[58]), .A1N(n58), .Y(
        n2477) );
  OAI2BB2X1 U1303 ( .B0(n1483), .B1(n58), .A0N(memory[59]), .A1N(n58), .Y(
        n2476) );
  OAI2BB2X1 U1304 ( .B0(n1488), .B1(n60), .A0N(memory[72]), .A1N(n60), .Y(
        n2463) );
  OAI2BB2X1 U1305 ( .B0(n1486), .B1(n60), .A0N(memory[73]), .A1N(n60), .Y(
        n2462) );
  OAI2BB2X1 U1306 ( .B0(n1484), .B1(n60), .A0N(memory[74]), .A1N(n60), .Y(
        n2461) );
  OAI2BB2X1 U1307 ( .B0(n1482), .B1(n60), .A0N(memory[75]), .A1N(n60), .Y(
        n2460) );
  OAI2BB2X1 U1308 ( .B0(n1489), .B1(n61), .A0N(memory[88]), .A1N(n61), .Y(
        n2447) );
  OAI2BB2X1 U1309 ( .B0(n1487), .B1(n61), .A0N(memory[89]), .A1N(n61), .Y(
        n2446) );
  OAI2BB2X1 U1310 ( .B0(n1485), .B1(n61), .A0N(memory[90]), .A1N(n61), .Y(
        n2445) );
  OAI2BB2X1 U1311 ( .B0(n1483), .B1(n61), .A0N(memory[91]), .A1N(n61), .Y(
        n2444) );
  OAI2BB2X1 U1312 ( .B0(n1488), .B1(n62), .A0N(memory[104]), .A1N(n62), .Y(
        n2431) );
  OAI2BB2X1 U1313 ( .B0(n1486), .B1(n62), .A0N(memory[105]), .A1N(n62), .Y(
        n2430) );
  OAI2BB2X1 U1314 ( .B0(n1484), .B1(n62), .A0N(memory[106]), .A1N(n62), .Y(
        n2429) );
  OAI2BB2X1 U1315 ( .B0(n1482), .B1(n62), .A0N(memory[107]), .A1N(n62), .Y(
        n2428) );
  OAI2BB2X1 U1316 ( .B0(n1489), .B1(n3), .A0N(memory[120]), .A1N(n3), .Y(n2415) );
  OAI2BB2X1 U1317 ( .B0(n1487), .B1(n3), .A0N(memory[121]), .A1N(n3), .Y(n2414) );
  OAI2BB2X1 U1318 ( .B0(n1485), .B1(n3), .A0N(memory[122]), .A1N(n3), .Y(n2413) );
  OAI2BB2X1 U1319 ( .B0(n1483), .B1(n3), .A0N(memory[123]), .A1N(n3), .Y(n2412) );
  OAI2BB2X1 U1320 ( .B0(n1489), .B1(n4), .A0N(memory[136]), .A1N(n4), .Y(n2399) );
  OAI2BB2X1 U1321 ( .B0(n1487), .B1(n4), .A0N(memory[137]), .A1N(n4), .Y(n2398) );
  OAI2BB2X1 U1322 ( .B0(n1485), .B1(n4), .A0N(memory[138]), .A1N(n4), .Y(n2397) );
  OAI2BB2X1 U1323 ( .B0(n1483), .B1(n4), .A0N(memory[139]), .A1N(n4), .Y(n2396) );
  OAI2BB2X1 U1324 ( .B0(n1489), .B1(n5), .A0N(memory[152]), .A1N(n5), .Y(n2383) );
  OAI2BB2X1 U1325 ( .B0(n1487), .B1(n5), .A0N(memory[153]), .A1N(n5), .Y(n2382) );
  OAI2BB2X1 U1326 ( .B0(n1485), .B1(n5), .A0N(memory[154]), .A1N(n5), .Y(n2381) );
  OAI2BB2X1 U1327 ( .B0(n1483), .B1(n5), .A0N(memory[155]), .A1N(n5), .Y(n2380) );
  OAI2BB2X1 U1328 ( .B0(n1488), .B1(n63), .A0N(memory[168]), .A1N(n63), .Y(
        n2367) );
  OAI2BB2X1 U1329 ( .B0(n1486), .B1(n63), .A0N(memory[169]), .A1N(n63), .Y(
        n2366) );
  OAI2BB2X1 U1330 ( .B0(n1484), .B1(n63), .A0N(memory[170]), .A1N(n63), .Y(
        n2365) );
  OAI2BB2X1 U1331 ( .B0(n1482), .B1(n63), .A0N(memory[171]), .A1N(n63), .Y(
        n2364) );
  OAI2BB2X1 U1332 ( .B0(n1489), .B1(n64), .A0N(memory[184]), .A1N(n64), .Y(
        n2351) );
  OAI2BB2X1 U1333 ( .B0(n1487), .B1(n64), .A0N(memory[185]), .A1N(n64), .Y(
        n2350) );
  OAI2BB2X1 U1334 ( .B0(n1485), .B1(n64), .A0N(memory[186]), .A1N(n64), .Y(
        n2349) );
  OAI2BB2X1 U1335 ( .B0(n1483), .B1(n64), .A0N(memory[187]), .A1N(n64), .Y(
        n2348) );
  OAI2BB2X1 U1336 ( .B0(n1489), .B1(n65), .A0N(memory[200]), .A1N(n65), .Y(
        n2335) );
  OAI2BB2X1 U1337 ( .B0(n1487), .B1(n65), .A0N(memory[201]), .A1N(n65), .Y(
        n2334) );
  OAI2BB2X1 U1338 ( .B0(n1485), .B1(n65), .A0N(memory[202]), .A1N(n65), .Y(
        n2333) );
  OAI2BB2X1 U1339 ( .B0(n1483), .B1(n65), .A0N(memory[203]), .A1N(n65), .Y(
        n2332) );
  OAI2BB2X1 U1340 ( .B0(n1489), .B1(n66), .A0N(memory[216]), .A1N(n66), .Y(
        n2319) );
  OAI2BB2X1 U1341 ( .B0(n1487), .B1(n66), .A0N(memory[217]), .A1N(n66), .Y(
        n2318) );
  OAI2BB2X1 U1342 ( .B0(n1485), .B1(n66), .A0N(memory[218]), .A1N(n66), .Y(
        n2317) );
  OAI2BB2X1 U1343 ( .B0(n1483), .B1(n66), .A0N(memory[219]), .A1N(n66), .Y(
        n2316) );
  OAI2BB2X1 U1344 ( .B0(n1489), .B1(n67), .A0N(memory[232]), .A1N(n67), .Y(
        n2303) );
  OAI2BB2X1 U1345 ( .B0(n1487), .B1(n67), .A0N(memory[233]), .A1N(n67), .Y(
        n2302) );
  OAI2BB2X1 U1346 ( .B0(n1485), .B1(n67), .A0N(memory[234]), .A1N(n67), .Y(
        n2301) );
  OAI2BB2X1 U1347 ( .B0(n1483), .B1(n67), .A0N(memory[235]), .A1N(n67), .Y(
        n2300) );
  OAI2BB2X1 U1348 ( .B0(n1489), .B1(n6), .A0N(memory[248]), .A1N(n6), .Y(n2287) );
  OAI2BB2X1 U1349 ( .B0(n1487), .B1(n6), .A0N(memory[249]), .A1N(n6), .Y(n2286) );
  OAI2BB2X1 U1350 ( .B0(n1485), .B1(n6), .A0N(memory[250]), .A1N(n6), .Y(n2285) );
  OAI2BB2X1 U1351 ( .B0(n1483), .B1(n6), .A0N(memory[251]), .A1N(n6), .Y(n2284) );
  OAI2BB2X1 U1352 ( .B0(n1489), .B1(n7), .A0N(memory[264]), .A1N(n7), .Y(n2271) );
  OAI2BB2X1 U1353 ( .B0(n1487), .B1(n7), .A0N(memory[265]), .A1N(n7), .Y(n2270) );
  OAI2BB2X1 U1354 ( .B0(n1485), .B1(n7), .A0N(memory[266]), .A1N(n7), .Y(n2269) );
  OAI2BB2X1 U1355 ( .B0(n1483), .B1(n7), .A0N(memory[267]), .A1N(n7), .Y(n2268) );
  OAI2BB2X1 U1356 ( .B0(n1489), .B1(n8), .A0N(memory[280]), .A1N(n8), .Y(n2255) );
  OAI2BB2X1 U1357 ( .B0(n1487), .B1(n8), .A0N(memory[281]), .A1N(n8), .Y(n2254) );
  OAI2BB2X1 U1358 ( .B0(n1485), .B1(n8), .A0N(memory[282]), .A1N(n8), .Y(n2253) );
  OAI2BB2X1 U1359 ( .B0(n1483), .B1(n8), .A0N(memory[283]), .A1N(n8), .Y(n2252) );
  OAI2BB2X1 U1360 ( .B0(n1489), .B1(n69), .A0N(memory[296]), .A1N(n69), .Y(
        n2239) );
  OAI2BB2X1 U1361 ( .B0(n1487), .B1(n69), .A0N(memory[297]), .A1N(n69), .Y(
        n2238) );
  OAI2BB2X1 U1362 ( .B0(n1485), .B1(n69), .A0N(memory[298]), .A1N(n69), .Y(
        n2237) );
  OAI2BB2X1 U1363 ( .B0(n1483), .B1(n69), .A0N(memory[299]), .A1N(n69), .Y(
        n2236) );
  OAI2BB2X1 U1364 ( .B0(n1489), .B1(n70), .A0N(memory[312]), .A1N(n70), .Y(
        n2223) );
  OAI2BB2X1 U1365 ( .B0(n1487), .B1(n70), .A0N(memory[313]), .A1N(n70), .Y(
        n2222) );
  OAI2BB2X1 U1366 ( .B0(n1485), .B1(n70), .A0N(memory[314]), .A1N(n70), .Y(
        n2221) );
  OAI2BB2X1 U1367 ( .B0(n1483), .B1(n70), .A0N(memory[315]), .A1N(n70), .Y(
        n2220) );
  OAI2BB2X1 U1368 ( .B0(n1489), .B1(n71), .A0N(memory[328]), .A1N(n71), .Y(
        n2207) );
  OAI2BB2X1 U1369 ( .B0(n1487), .B1(n71), .A0N(memory[329]), .A1N(n71), .Y(
        n2206) );
  OAI2BB2X1 U1370 ( .B0(n1485), .B1(n71), .A0N(memory[330]), .A1N(n71), .Y(
        n2205) );
  OAI2BB2X1 U1371 ( .B0(n1483), .B1(n71), .A0N(memory[331]), .A1N(n71), .Y(
        n2204) );
  OAI2BB2X1 U1372 ( .B0(n1489), .B1(n72), .A0N(memory[344]), .A1N(n72), .Y(
        n2191) );
  OAI2BB2X1 U1373 ( .B0(n1487), .B1(n72), .A0N(memory[345]), .A1N(n72), .Y(
        n2190) );
  OAI2BB2X1 U1374 ( .B0(n1485), .B1(n72), .A0N(memory[346]), .A1N(n72), .Y(
        n2189) );
  OAI2BB2X1 U1375 ( .B0(n1483), .B1(n72), .A0N(memory[347]), .A1N(n72), .Y(
        n2188) );
  OAI2BB2X1 U1376 ( .B0(n1489), .B1(n73), .A0N(memory[360]), .A1N(n73), .Y(
        n2175) );
  OAI2BB2X1 U1377 ( .B0(n1487), .B1(n73), .A0N(memory[361]), .A1N(n73), .Y(
        n2174) );
  OAI2BB2X1 U1378 ( .B0(n1485), .B1(n73), .A0N(memory[362]), .A1N(n73), .Y(
        n2173) );
  OAI2BB2X1 U1379 ( .B0(n1483), .B1(n73), .A0N(memory[363]), .A1N(n73), .Y(
        n2172) );
  OAI2BB2X1 U1380 ( .B0(n1489), .B1(n9), .A0N(memory[376]), .A1N(n9), .Y(n2159) );
  OAI2BB2X1 U1381 ( .B0(n1487), .B1(n9), .A0N(memory[377]), .A1N(n9), .Y(n2158) );
  OAI2BB2X1 U1382 ( .B0(n1485), .B1(n9), .A0N(memory[378]), .A1N(n9), .Y(n2157) );
  OAI2BB2X1 U1383 ( .B0(n1483), .B1(n9), .A0N(memory[379]), .A1N(n9), .Y(n2156) );
  OAI2BB2X1 U1384 ( .B0(n1489), .B1(n10), .A0N(memory[392]), .A1N(n10), .Y(
        n2143) );
  OAI2BB2X1 U1385 ( .B0(n1487), .B1(n10), .A0N(memory[393]), .A1N(n10), .Y(
        n2142) );
  OAI2BB2X1 U1386 ( .B0(n1485), .B1(n10), .A0N(memory[394]), .A1N(n10), .Y(
        n2141) );
  OAI2BB2X1 U1387 ( .B0(n1483), .B1(n10), .A0N(memory[395]), .A1N(n10), .Y(
        n2140) );
  OAI2BB2X1 U1388 ( .B0(n1488), .B1(n11), .A0N(memory[408]), .A1N(n11), .Y(
        n2127) );
  OAI2BB2X1 U1389 ( .B0(n1486), .B1(n11), .A0N(memory[409]), .A1N(n11), .Y(
        n2126) );
  OAI2BB2X1 U1390 ( .B0(n1484), .B1(n11), .A0N(memory[410]), .A1N(n11), .Y(
        n2125) );
  OAI2BB2X1 U1391 ( .B0(n1482), .B1(n11), .A0N(memory[411]), .A1N(n11), .Y(
        n2124) );
  OAI2BB2X1 U1392 ( .B0(n1489), .B1(n74), .A0N(memory[424]), .A1N(n74), .Y(
        n2111) );
  OAI2BB2X1 U1393 ( .B0(n1487), .B1(n74), .A0N(memory[425]), .A1N(n74), .Y(
        n2110) );
  OAI2BB2X1 U1394 ( .B0(n1485), .B1(n74), .A0N(memory[426]), .A1N(n74), .Y(
        n2109) );
  OAI2BB2X1 U1395 ( .B0(n1483), .B1(n74), .A0N(memory[427]), .A1N(n74), .Y(
        n2108) );
  OAI2BB2X1 U1396 ( .B0(n1489), .B1(n75), .A0N(memory[440]), .A1N(n75), .Y(
        n2095) );
  OAI2BB2X1 U1397 ( .B0(n1487), .B1(n75), .A0N(memory[441]), .A1N(n75), .Y(
        n2094) );
  OAI2BB2X1 U1398 ( .B0(n1485), .B1(n75), .A0N(memory[442]), .A1N(n75), .Y(
        n2093) );
  OAI2BB2X1 U1399 ( .B0(n1483), .B1(n75), .A0N(memory[443]), .A1N(n75), .Y(
        n2092) );
  OAI2BB2X1 U1400 ( .B0(n1489), .B1(n76), .A0N(memory[456]), .A1N(n76), .Y(
        n2079) );
  OAI2BB2X1 U1401 ( .B0(n1487), .B1(n76), .A0N(memory[457]), .A1N(n76), .Y(
        n2078) );
  OAI2BB2X1 U1402 ( .B0(n1485), .B1(n76), .A0N(memory[458]), .A1N(n76), .Y(
        n2077) );
  OAI2BB2X1 U1403 ( .B0(n1483), .B1(n76), .A0N(memory[459]), .A1N(n76), .Y(
        n2076) );
  OAI2BB2X1 U1404 ( .B0(n1488), .B1(n78), .A0N(memory[472]), .A1N(n78), .Y(
        n2063) );
  OAI2BB2X1 U1405 ( .B0(n1486), .B1(n78), .A0N(memory[473]), .A1N(n78), .Y(
        n2062) );
  OAI2BB2X1 U1406 ( .B0(n1484), .B1(n78), .A0N(memory[474]), .A1N(n78), .Y(
        n2061) );
  OAI2BB2X1 U1407 ( .B0(n1482), .B1(n78), .A0N(memory[475]), .A1N(n78), .Y(
        n2060) );
  OAI2BB2X1 U1408 ( .B0(n1489), .B1(n79), .A0N(memory[488]), .A1N(n79), .Y(
        n2047) );
  OAI2BB2X1 U1409 ( .B0(n1487), .B1(n79), .A0N(memory[489]), .A1N(n79), .Y(
        n2046) );
  OAI2BB2X1 U1410 ( .B0(n1485), .B1(n79), .A0N(memory[490]), .A1N(n79), .Y(
        n2045) );
  OAI2BB2X1 U1411 ( .B0(n1483), .B1(n79), .A0N(memory[491]), .A1N(n79), .Y(
        n2044) );
  OAI2BB2X1 U1412 ( .B0(n1488), .B1(n12), .A0N(memory[504]), .A1N(n12), .Y(
        n2031) );
  OAI2BB2X1 U1413 ( .B0(n1486), .B1(n12), .A0N(memory[505]), .A1N(n12), .Y(
        n2030) );
  OAI2BB2X1 U1414 ( .B0(n1484), .B1(n12), .A0N(memory[506]), .A1N(n12), .Y(
        n2029) );
  OAI2BB2X1 U1415 ( .B0(n1482), .B1(n12), .A0N(memory[507]), .A1N(n12), .Y(
        n2028) );
  OAI2BB2X1 U1416 ( .B0(n1489), .B1(n13), .A0N(memory[520]), .A1N(n13), .Y(
        n2015) );
  OAI2BB2X1 U1417 ( .B0(n1487), .B1(n13), .A0N(memory[521]), .A1N(n13), .Y(
        n2014) );
  OAI2BB2X1 U1418 ( .B0(n1485), .B1(n13), .A0N(memory[522]), .A1N(n13), .Y(
        n2013) );
  OAI2BB2X1 U1419 ( .B0(n1483), .B1(n13), .A0N(memory[523]), .A1N(n13), .Y(
        n2012) );
  OAI2BB2X1 U1420 ( .B0(n1488), .B1(n14), .A0N(memory[536]), .A1N(n14), .Y(
        n1999) );
  OAI2BB2X1 U1421 ( .B0(n1486), .B1(n14), .A0N(memory[537]), .A1N(n14), .Y(
        n1998) );
  OAI2BB2X1 U1422 ( .B0(n1484), .B1(n14), .A0N(memory[538]), .A1N(n14), .Y(
        n1997) );
  OAI2BB2X1 U1423 ( .B0(n1482), .B1(n14), .A0N(memory[539]), .A1N(n14), .Y(
        n1996) );
  OAI2BB2X1 U1424 ( .B0(n1489), .B1(n15), .A0N(memory[552]), .A1N(n15), .Y(
        n1983) );
  OAI2BB2X1 U1425 ( .B0(n1487), .B1(n15), .A0N(memory[553]), .A1N(n15), .Y(
        n1982) );
  OAI2BB2X1 U1426 ( .B0(n1485), .B1(n15), .A0N(memory[554]), .A1N(n15), .Y(
        n1981) );
  OAI2BB2X1 U1427 ( .B0(n1483), .B1(n15), .A0N(memory[555]), .A1N(n15), .Y(
        n1980) );
  OAI2BB2X1 U1428 ( .B0(n1488), .B1(n16), .A0N(memory[568]), .A1N(n16), .Y(
        n1967) );
  OAI2BB2X1 U1429 ( .B0(n1486), .B1(n16), .A0N(memory[569]), .A1N(n16), .Y(
        n1966) );
  OAI2BB2X1 U1430 ( .B0(n1484), .B1(n16), .A0N(memory[570]), .A1N(n16), .Y(
        n1965) );
  OAI2BB2X1 U1431 ( .B0(n1482), .B1(n16), .A0N(memory[571]), .A1N(n16), .Y(
        n1964) );
  OAI2BB2X1 U1432 ( .B0(n1489), .B1(n17), .A0N(memory[584]), .A1N(n17), .Y(
        n1951) );
  OAI2BB2X1 U1433 ( .B0(n1487), .B1(n17), .A0N(memory[585]), .A1N(n17), .Y(
        n1950) );
  OAI2BB2X1 U1434 ( .B0(n1485), .B1(n17), .A0N(memory[586]), .A1N(n17), .Y(
        n1949) );
  OAI2BB2X1 U1435 ( .B0(n1483), .B1(n17), .A0N(memory[587]), .A1N(n17), .Y(
        n1948) );
  OAI2BB2X1 U1436 ( .B0(n1488), .B1(n18), .A0N(memory[600]), .A1N(n18), .Y(
        n1935) );
  OAI2BB2X1 U1437 ( .B0(n1486), .B1(n18), .A0N(memory[601]), .A1N(n18), .Y(
        n1934) );
  OAI2BB2X1 U1438 ( .B0(n1484), .B1(n18), .A0N(memory[602]), .A1N(n18), .Y(
        n1933) );
  OAI2BB2X1 U1439 ( .B0(n1482), .B1(n18), .A0N(memory[603]), .A1N(n18), .Y(
        n1932) );
  OAI2BB2X1 U1440 ( .B0(n1488), .B1(n19), .A0N(memory[616]), .A1N(n19), .Y(
        n1919) );
  OAI2BB2X1 U1441 ( .B0(n1486), .B1(n19), .A0N(memory[617]), .A1N(n19), .Y(
        n1918) );
  OAI2BB2X1 U1442 ( .B0(n1484), .B1(n19), .A0N(memory[618]), .A1N(n19), .Y(
        n1917) );
  OAI2BB2X1 U1443 ( .B0(n1482), .B1(n19), .A0N(memory[619]), .A1N(n19), .Y(
        n1916) );
  OAI2BB2X1 U1444 ( .B0(n1489), .B1(n20), .A0N(memory[632]), .A1N(n20), .Y(
        n1903) );
  OAI2BB2X1 U1445 ( .B0(n1487), .B1(n20), .A0N(memory[633]), .A1N(n20), .Y(
        n1902) );
  OAI2BB2X1 U1446 ( .B0(n1485), .B1(n20), .A0N(memory[634]), .A1N(n20), .Y(
        n1901) );
  OAI2BB2X1 U1447 ( .B0(n1483), .B1(n20), .A0N(memory[635]), .A1N(n20), .Y(
        n1900) );
  OAI2BB2X1 U1448 ( .B0(n1488), .B1(n21), .A0N(memory[648]), .A1N(n21), .Y(
        n1887) );
  OAI2BB2X1 U1449 ( .B0(n1486), .B1(n21), .A0N(memory[649]), .A1N(n21), .Y(
        n1886) );
  OAI2BB2X1 U1450 ( .B0(n1484), .B1(n21), .A0N(memory[650]), .A1N(n21), .Y(
        n1885) );
  OAI2BB2X1 U1451 ( .B0(n1482), .B1(n21), .A0N(memory[651]), .A1N(n21), .Y(
        n1884) );
  OAI2BB2X1 U1452 ( .B0(n1488), .B1(n22), .A0N(memory[664]), .A1N(n22), .Y(
        n1871) );
  OAI2BB2X1 U1453 ( .B0(n1486), .B1(n22), .A0N(memory[665]), .A1N(n22), .Y(
        n1870) );
  OAI2BB2X1 U1454 ( .B0(n1484), .B1(n22), .A0N(memory[666]), .A1N(n22), .Y(
        n1869) );
  OAI2BB2X1 U1455 ( .B0(n1482), .B1(n22), .A0N(memory[667]), .A1N(n22), .Y(
        n1868) );
  OAI2BB2X1 U1456 ( .B0(n1489), .B1(n25), .A0N(memory[680]), .A1N(n25), .Y(
        n1855) );
  OAI2BB2X1 U1457 ( .B0(n1487), .B1(n25), .A0N(memory[681]), .A1N(n25), .Y(
        n1854) );
  OAI2BB2X1 U1458 ( .B0(n1485), .B1(n25), .A0N(memory[682]), .A1N(n25), .Y(
        n1853) );
  OAI2BB2X1 U1459 ( .B0(n1483), .B1(n25), .A0N(memory[683]), .A1N(n25), .Y(
        n1852) );
  OAI2BB2X1 U1460 ( .B0(n1488), .B1(n27), .A0N(memory[696]), .A1N(n27), .Y(
        n1839) );
  OAI2BB2X1 U1461 ( .B0(n1486), .B1(n27), .A0N(memory[697]), .A1N(n27), .Y(
        n1838) );
  OAI2BB2X1 U1462 ( .B0(n1484), .B1(n27), .A0N(memory[698]), .A1N(n27), .Y(
        n1837) );
  OAI2BB2X1 U1463 ( .B0(n1482), .B1(n27), .A0N(memory[699]), .A1N(n27), .Y(
        n1836) );
  OAI2BB2X1 U1464 ( .B0(n1489), .B1(n29), .A0N(memory[712]), .A1N(n29), .Y(
        n1823) );
  OAI2BB2X1 U1465 ( .B0(n1487), .B1(n29), .A0N(memory[713]), .A1N(n29), .Y(
        n1822) );
  OAI2BB2X1 U1466 ( .B0(n1485), .B1(n29), .A0N(memory[714]), .A1N(n29), .Y(
        n1821) );
  OAI2BB2X1 U1467 ( .B0(n1483), .B1(n29), .A0N(memory[715]), .A1N(n29), .Y(
        n1820) );
  OAI2BB2X1 U1468 ( .B0(n1488), .B1(n31), .A0N(memory[728]), .A1N(n31), .Y(
        n1807) );
  OAI2BB2X1 U1469 ( .B0(n1486), .B1(n31), .A0N(memory[729]), .A1N(n31), .Y(
        n1806) );
  OAI2BB2X1 U1470 ( .B0(n1484), .B1(n31), .A0N(memory[730]), .A1N(n31), .Y(
        n1805) );
  OAI2BB2X1 U1471 ( .B0(n1482), .B1(n31), .A0N(memory[731]), .A1N(n31), .Y(
        n1804) );
  OAI2BB2X1 U1472 ( .B0(n1489), .B1(n33), .A0N(memory[744]), .A1N(n33), .Y(
        n1791) );
  OAI2BB2X1 U1473 ( .B0(n1487), .B1(n33), .A0N(memory[745]), .A1N(n33), .Y(
        n1790) );
  OAI2BB2X1 U1474 ( .B0(n1485), .B1(n33), .A0N(memory[746]), .A1N(n33), .Y(
        n1789) );
  OAI2BB2X1 U1475 ( .B0(n1483), .B1(n33), .A0N(memory[747]), .A1N(n33), .Y(
        n1788) );
  OAI2BB2X1 U1476 ( .B0(n1488), .B1(n35), .A0N(memory[760]), .A1N(n35), .Y(
        n1775) );
  OAI2BB2X1 U1477 ( .B0(n1486), .B1(n35), .A0N(memory[761]), .A1N(n35), .Y(
        n1774) );
  OAI2BB2X1 U1478 ( .B0(n1484), .B1(n35), .A0N(memory[762]), .A1N(n35), .Y(
        n1773) );
  OAI2BB2X1 U1479 ( .B0(n1482), .B1(n35), .A0N(memory[763]), .A1N(n35), .Y(
        n1772) );
  OAI2BB2X1 U1480 ( .B0(n1488), .B1(n37), .A0N(memory[776]), .A1N(n37), .Y(
        n1759) );
  OAI2BB2X1 U1481 ( .B0(n1486), .B1(n37), .A0N(memory[777]), .A1N(n37), .Y(
        n1758) );
  OAI2BB2X1 U1482 ( .B0(n1484), .B1(n37), .A0N(memory[778]), .A1N(n37), .Y(
        n1757) );
  OAI2BB2X1 U1483 ( .B0(n1482), .B1(n37), .A0N(memory[779]), .A1N(n37), .Y(
        n1756) );
  OAI2BB2X1 U1484 ( .B0(n1489), .B1(n40), .A0N(memory[792]), .A1N(n40), .Y(
        n1743) );
  OAI2BB2X1 U1485 ( .B0(n1487), .B1(n40), .A0N(memory[793]), .A1N(n40), .Y(
        n1742) );
  OAI2BB2X1 U1486 ( .B0(n1485), .B1(n40), .A0N(memory[794]), .A1N(n40), .Y(
        n1741) );
  OAI2BB2X1 U1487 ( .B0(n1483), .B1(n40), .A0N(memory[795]), .A1N(n40), .Y(
        n1740) );
  OAI2BB2X1 U1488 ( .B0(n1488), .B1(n42), .A0N(memory[808]), .A1N(n42), .Y(
        n1727) );
  OAI2BB2X1 U1489 ( .B0(n1486), .B1(n42), .A0N(memory[809]), .A1N(n42), .Y(
        n1726) );
  OAI2BB2X1 U1490 ( .B0(n1484), .B1(n42), .A0N(memory[810]), .A1N(n42), .Y(
        n1725) );
  OAI2BB2X1 U1491 ( .B0(n1482), .B1(n42), .A0N(memory[811]), .A1N(n42), .Y(
        n1724) );
  OAI2BB2X1 U1492 ( .B0(n1488), .B1(n43), .A0N(memory[824]), .A1N(n43), .Y(
        n1711) );
  OAI2BB2X1 U1493 ( .B0(n1486), .B1(n43), .A0N(memory[825]), .A1N(n43), .Y(
        n1710) );
  OAI2BB2X1 U1494 ( .B0(n1484), .B1(n43), .A0N(memory[826]), .A1N(n43), .Y(
        n1709) );
  OAI2BB2X1 U1495 ( .B0(n1482), .B1(n43), .A0N(memory[827]), .A1N(n43), .Y(
        n1708) );
  OAI2BB2X1 U1496 ( .B0(n1488), .B1(n44), .A0N(memory[840]), .A1N(n44), .Y(
        n1695) );
  OAI2BB2X1 U1497 ( .B0(n1486), .B1(n44), .A0N(memory[841]), .A1N(n44), .Y(
        n1694) );
  OAI2BB2X1 U1498 ( .B0(n1484), .B1(n44), .A0N(memory[842]), .A1N(n44), .Y(
        n1693) );
  OAI2BB2X1 U1499 ( .B0(n1482), .B1(n44), .A0N(memory[843]), .A1N(n44), .Y(
        n1692) );
  OAI2BB2X1 U1500 ( .B0(n1488), .B1(n45), .A0N(memory[856]), .A1N(n45), .Y(
        n1679) );
  OAI2BB2X1 U1501 ( .B0(n1486), .B1(n45), .A0N(memory[857]), .A1N(n45), .Y(
        n1678) );
  OAI2BB2X1 U1502 ( .B0(n1484), .B1(n45), .A0N(memory[858]), .A1N(n45), .Y(
        n1677) );
  OAI2BB2X1 U1503 ( .B0(n1482), .B1(n45), .A0N(memory[859]), .A1N(n45), .Y(
        n1676) );
  OAI2BB2X1 U1504 ( .B0(n1488), .B1(n46), .A0N(memory[872]), .A1N(n46), .Y(
        n1663) );
  OAI2BB2X1 U1505 ( .B0(n1486), .B1(n46), .A0N(memory[873]), .A1N(n46), .Y(
        n1662) );
  OAI2BB2X1 U1506 ( .B0(n1484), .B1(n46), .A0N(memory[874]), .A1N(n46), .Y(
        n1661) );
  OAI2BB2X1 U1507 ( .B0(n1482), .B1(n46), .A0N(memory[875]), .A1N(n46), .Y(
        n1660) );
  OAI2BB2X1 U1508 ( .B0(n1488), .B1(n47), .A0N(memory[888]), .A1N(n47), .Y(
        n1647) );
  OAI2BB2X1 U1509 ( .B0(n1486), .B1(n47), .A0N(memory[889]), .A1N(n47), .Y(
        n1646) );
  OAI2BB2X1 U1510 ( .B0(n1484), .B1(n47), .A0N(memory[890]), .A1N(n47), .Y(
        n1645) );
  OAI2BB2X1 U1511 ( .B0(n1482), .B1(n47), .A0N(memory[891]), .A1N(n47), .Y(
        n1644) );
  OAI2BB2X1 U1512 ( .B0(n1488), .B1(n48), .A0N(memory[904]), .A1N(n48), .Y(
        n1631) );
  OAI2BB2X1 U1513 ( .B0(n1486), .B1(n48), .A0N(memory[905]), .A1N(n48), .Y(
        n1630) );
  OAI2BB2X1 U1514 ( .B0(n1484), .B1(n48), .A0N(memory[906]), .A1N(n48), .Y(
        n1629) );
  OAI2BB2X1 U1515 ( .B0(n1482), .B1(n48), .A0N(memory[907]), .A1N(n48), .Y(
        n1628) );
  OAI2BB2X1 U1516 ( .B0(n1488), .B1(n49), .A0N(memory[920]), .A1N(n49), .Y(
        n1615) );
  OAI2BB2X1 U1517 ( .B0(n1486), .B1(n49), .A0N(memory[921]), .A1N(n49), .Y(
        n1614) );
  OAI2BB2X1 U1518 ( .B0(n1484), .B1(n49), .A0N(memory[922]), .A1N(n49), .Y(
        n1613) );
  OAI2BB2X1 U1519 ( .B0(n1482), .B1(n49), .A0N(memory[923]), .A1N(n49), .Y(
        n1612) );
  OAI2BB2X1 U1520 ( .B0(n1488), .B1(n51), .A0N(memory[936]), .A1N(n51), .Y(
        n1599) );
  OAI2BB2X1 U1521 ( .B0(n1486), .B1(n51), .A0N(memory[937]), .A1N(n51), .Y(
        n1598) );
  OAI2BB2X1 U1522 ( .B0(n1484), .B1(n51), .A0N(memory[938]), .A1N(n51), .Y(
        n1597) );
  OAI2BB2X1 U1523 ( .B0(n1482), .B1(n51), .A0N(memory[939]), .A1N(n51), .Y(
        n1596) );
  OAI2BB2X1 U1524 ( .B0(n1488), .B1(n52), .A0N(memory[952]), .A1N(n52), .Y(
        n1583) );
  OAI2BB2X1 U1525 ( .B0(n1486), .B1(n52), .A0N(memory[953]), .A1N(n52), .Y(
        n1582) );
  OAI2BB2X1 U1526 ( .B0(n1484), .B1(n52), .A0N(memory[954]), .A1N(n52), .Y(
        n1581) );
  OAI2BB2X1 U1527 ( .B0(n1482), .B1(n52), .A0N(memory[955]), .A1N(n52), .Y(
        n1580) );
  OAI2BB2X1 U1528 ( .B0(n1488), .B1(n53), .A0N(memory[968]), .A1N(n53), .Y(
        n1567) );
  OAI2BB2X1 U1529 ( .B0(n1486), .B1(n53), .A0N(memory[969]), .A1N(n53), .Y(
        n1566) );
  OAI2BB2X1 U1530 ( .B0(n1484), .B1(n53), .A0N(memory[970]), .A1N(n53), .Y(
        n1565) );
  OAI2BB2X1 U1531 ( .B0(n1482), .B1(n53), .A0N(memory[971]), .A1N(n53), .Y(
        n1564) );
  OAI2BB2X1 U1532 ( .B0(n1488), .B1(n54), .A0N(memory[984]), .A1N(n54), .Y(
        n1551) );
  OAI2BB2X1 U1533 ( .B0(n1486), .B1(n54), .A0N(memory[985]), .A1N(n54), .Y(
        n1550) );
  OAI2BB2X1 U1534 ( .B0(n1484), .B1(n54), .A0N(memory[986]), .A1N(n54), .Y(
        n1549) );
  OAI2BB2X1 U1535 ( .B0(n1482), .B1(n54), .A0N(memory[987]), .A1N(n54), .Y(
        n1548) );
  OAI2BB2X1 U1536 ( .B0(n1488), .B1(n55), .A0N(memory[1000]), .A1N(n55), .Y(
        n1535) );
  OAI2BB2X1 U1537 ( .B0(n1486), .B1(n55), .A0N(memory[1001]), .A1N(n55), .Y(
        n1534) );
  OAI2BB2X1 U1538 ( .B0(n1484), .B1(n55), .A0N(memory[1002]), .A1N(n55), .Y(
        n1533) );
  OAI2BB2X1 U1539 ( .B0(n1482), .B1(n55), .A0N(memory[1003]), .A1N(n55), .Y(
        n1532) );
  OAI2BB2X1 U1540 ( .B0(n1488), .B1(n56), .A0N(memory[1016]), .A1N(n56), .Y(
        n1519) );
  OAI2BB2X1 U1541 ( .B0(n1486), .B1(n56), .A0N(memory[1017]), .A1N(n56), .Y(
        n1518) );
  OAI2BB2X1 U1542 ( .B0(n1484), .B1(n56), .A0N(memory[1018]), .A1N(n56), .Y(
        n1517) );
  OAI2BB2X1 U1543 ( .B0(n1482), .B1(n56), .A0N(memory[1019]), .A1N(n56), .Y(
        n1516) );
  BUFX3 U1544 ( .A(addr[5]), .Y(n1510) );
endmodule


module mem4x4_0 ( clk, rstn, en, wr_rd, addr, din, dout );
  input [3:0] addr;
  input [15:0] din;
  output [15:0] dout;
  input clk, rstn, en, wr_rd;
  wire   N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48,
         N49, N50, n21, n22, n24, n26, n29, n32, n33, n35, n37, n39, n45, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n23, n25, n27, n28, n30, n31,
         n34, n36, n38, n40, n41, n42, n43, n44, n46, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375;
  wire   [255:0] memory;

  DFFRHQX1 memory_reg_1__15_ ( .D(n287), .CK(clk), .RN(rstn), .Q(memory[239])
         );
  DFFRHQX1 memory_reg_1__14_ ( .D(n286), .CK(clk), .RN(rstn), .Q(memory[238])
         );
  DFFRHQX1 memory_reg_1__13_ ( .D(n285), .CK(clk), .RN(rstn), .Q(memory[237])
         );
  DFFRHQX1 memory_reg_1__12_ ( .D(n284), .CK(clk), .RN(rstn), .Q(memory[236])
         );
  DFFRHQX1 memory_reg_1__11_ ( .D(n283), .CK(clk), .RN(rstn), .Q(memory[235])
         );
  DFFRHQX1 memory_reg_1__10_ ( .D(n282), .CK(clk), .RN(rstn), .Q(memory[234])
         );
  DFFRHQX1 memory_reg_1__9_ ( .D(n281), .CK(clk), .RN(rstn), .Q(memory[233])
         );
  DFFRHQX1 memory_reg_1__8_ ( .D(n280), .CK(clk), .RN(rstn), .Q(memory[232])
         );
  DFFRHQX1 memory_reg_1__7_ ( .D(n279), .CK(clk), .RN(rstn), .Q(memory[231])
         );
  DFFRHQX1 memory_reg_1__6_ ( .D(n278), .CK(clk), .RN(rstn), .Q(memory[230])
         );
  DFFRHQX1 memory_reg_1__5_ ( .D(n277), .CK(clk), .RN(rstn), .Q(memory[229])
         );
  DFFRHQX1 memory_reg_1__4_ ( .D(n276), .CK(clk), .RN(rstn), .Q(memory[228])
         );
  DFFRHQX1 memory_reg_1__3_ ( .D(n275), .CK(clk), .RN(rstn), .Q(memory[227])
         );
  DFFRHQX1 memory_reg_1__2_ ( .D(n274), .CK(clk), .RN(rstn), .Q(memory[226])
         );
  DFFRHQX1 memory_reg_1__1_ ( .D(n273), .CK(clk), .RN(rstn), .Q(memory[225])
         );
  DFFRHQX1 memory_reg_1__0_ ( .D(n272), .CK(clk), .RN(rstn), .Q(memory[224])
         );
  DFFRHQX1 memory_reg_5__15_ ( .D(n223), .CK(clk), .RN(rstn), .Q(memory[175])
         );
  DFFRHQX1 memory_reg_5__14_ ( .D(n222), .CK(clk), .RN(rstn), .Q(memory[174])
         );
  DFFRHQX1 memory_reg_5__13_ ( .D(n221), .CK(clk), .RN(rstn), .Q(memory[173])
         );
  DFFRHQX1 memory_reg_5__12_ ( .D(n220), .CK(clk), .RN(rstn), .Q(memory[172])
         );
  DFFRHQX1 memory_reg_5__11_ ( .D(n219), .CK(clk), .RN(rstn), .Q(memory[171])
         );
  DFFRHQX1 memory_reg_5__10_ ( .D(n218), .CK(clk), .RN(rstn), .Q(memory[170])
         );
  DFFRHQX1 memory_reg_5__9_ ( .D(n217), .CK(clk), .RN(rstn), .Q(memory[169])
         );
  DFFRHQX1 memory_reg_5__8_ ( .D(n216), .CK(clk), .RN(rstn), .Q(memory[168])
         );
  DFFRHQX1 memory_reg_5__7_ ( .D(n215), .CK(clk), .RN(rstn), .Q(memory[167])
         );
  DFFRHQX1 memory_reg_5__6_ ( .D(n214), .CK(clk), .RN(rstn), .Q(memory[166])
         );
  DFFRHQX1 memory_reg_5__5_ ( .D(n213), .CK(clk), .RN(rstn), .Q(memory[165])
         );
  DFFRHQX1 memory_reg_5__4_ ( .D(n212), .CK(clk), .RN(rstn), .Q(memory[164])
         );
  DFFRHQX1 memory_reg_5__3_ ( .D(n211), .CK(clk), .RN(rstn), .Q(memory[163])
         );
  DFFRHQX1 memory_reg_5__2_ ( .D(n210), .CK(clk), .RN(rstn), .Q(memory[162])
         );
  DFFRHQX1 memory_reg_5__1_ ( .D(n209), .CK(clk), .RN(rstn), .Q(memory[161])
         );
  DFFRHQX1 memory_reg_5__0_ ( .D(n208), .CK(clk), .RN(rstn), .Q(memory[160])
         );
  DFFRHQX1 memory_reg_9__15_ ( .D(n159), .CK(clk), .RN(rstn), .Q(memory[111])
         );
  DFFRHQX1 memory_reg_9__14_ ( .D(n158), .CK(clk), .RN(rstn), .Q(memory[110])
         );
  DFFRHQX1 memory_reg_9__13_ ( .D(n157), .CK(clk), .RN(rstn), .Q(memory[109])
         );
  DFFRHQX1 memory_reg_9__12_ ( .D(n156), .CK(clk), .RN(rstn), .Q(memory[108])
         );
  DFFRHQX1 memory_reg_9__11_ ( .D(n155), .CK(clk), .RN(rstn), .Q(memory[107])
         );
  DFFRHQX1 memory_reg_9__10_ ( .D(n154), .CK(clk), .RN(rstn), .Q(memory[106])
         );
  DFFRHQX1 memory_reg_9__9_ ( .D(n153), .CK(clk), .RN(rstn), .Q(memory[105])
         );
  DFFRHQX1 memory_reg_9__8_ ( .D(n152), .CK(clk), .RN(rstn), .Q(memory[104])
         );
  DFFRHQX1 memory_reg_9__7_ ( .D(n151), .CK(clk), .RN(rstn), .Q(memory[103])
         );
  DFFRHQX1 memory_reg_9__6_ ( .D(n150), .CK(clk), .RN(rstn), .Q(memory[102])
         );
  DFFRHQX1 memory_reg_9__5_ ( .D(n149), .CK(clk), .RN(rstn), .Q(memory[101])
         );
  DFFRHQX1 memory_reg_9__4_ ( .D(n148), .CK(clk), .RN(rstn), .Q(memory[100])
         );
  DFFRHQX1 memory_reg_9__3_ ( .D(n147), .CK(clk), .RN(rstn), .Q(memory[99]) );
  DFFRHQX1 memory_reg_9__2_ ( .D(n146), .CK(clk), .RN(rstn), .Q(memory[98]) );
  DFFRHQX1 memory_reg_9__1_ ( .D(n145), .CK(clk), .RN(rstn), .Q(memory[97]) );
  DFFRHQX1 memory_reg_9__0_ ( .D(n144), .CK(clk), .RN(rstn), .Q(memory[96]) );
  DFFRHQX1 memory_reg_13__15_ ( .D(n95), .CK(clk), .RN(rstn), .Q(memory[47])
         );
  DFFRHQX1 memory_reg_13__14_ ( .D(n94), .CK(clk), .RN(rstn), .Q(memory[46])
         );
  DFFRHQX1 memory_reg_13__13_ ( .D(n93), .CK(clk), .RN(rstn), .Q(memory[45])
         );
  DFFRHQX1 memory_reg_13__12_ ( .D(n92), .CK(clk), .RN(rstn), .Q(memory[44])
         );
  DFFRHQX1 memory_reg_13__11_ ( .D(n91), .CK(clk), .RN(rstn), .Q(memory[43])
         );
  DFFRHQX1 memory_reg_13__10_ ( .D(n90), .CK(clk), .RN(rstn), .Q(memory[42])
         );
  DFFRHQX1 memory_reg_13__9_ ( .D(n89), .CK(clk), .RN(rstn), .Q(memory[41]) );
  DFFRHQX1 memory_reg_13__8_ ( .D(n88), .CK(clk), .RN(rstn), .Q(memory[40]) );
  DFFRHQX1 memory_reg_13__7_ ( .D(n87), .CK(clk), .RN(rstn), .Q(memory[39]) );
  DFFRHQX1 memory_reg_13__6_ ( .D(n86), .CK(clk), .RN(rstn), .Q(memory[38]) );
  DFFRHQX1 memory_reg_13__5_ ( .D(n85), .CK(clk), .RN(rstn), .Q(memory[37]) );
  DFFRHQX1 memory_reg_13__4_ ( .D(n84), .CK(clk), .RN(rstn), .Q(memory[36]) );
  DFFRHQX1 memory_reg_13__3_ ( .D(n83), .CK(clk), .RN(rstn), .Q(memory[35]) );
  DFFRHQX1 memory_reg_13__2_ ( .D(n82), .CK(clk), .RN(rstn), .Q(memory[34]) );
  DFFRHQX1 memory_reg_13__1_ ( .D(n81), .CK(clk), .RN(rstn), .Q(memory[33]) );
  DFFRHQX1 memory_reg_13__0_ ( .D(n80), .CK(clk), .RN(rstn), .Q(memory[32]) );
  DFFRHQX1 memory_reg_3__15_ ( .D(n255), .CK(clk), .RN(rstn), .Q(memory[207])
         );
  DFFRHQX1 memory_reg_3__14_ ( .D(n254), .CK(clk), .RN(rstn), .Q(memory[206])
         );
  DFFRHQX1 memory_reg_3__13_ ( .D(n253), .CK(clk), .RN(rstn), .Q(memory[205])
         );
  DFFRHQX1 memory_reg_3__12_ ( .D(n252), .CK(clk), .RN(rstn), .Q(memory[204])
         );
  DFFRHQX1 memory_reg_3__11_ ( .D(n251), .CK(clk), .RN(rstn), .Q(memory[203])
         );
  DFFRHQX1 memory_reg_3__10_ ( .D(n250), .CK(clk), .RN(rstn), .Q(memory[202])
         );
  DFFRHQX1 memory_reg_3__9_ ( .D(n249), .CK(clk), .RN(rstn), .Q(memory[201])
         );
  DFFRHQX1 memory_reg_3__8_ ( .D(n248), .CK(clk), .RN(rstn), .Q(memory[200])
         );
  DFFRHQX1 memory_reg_3__7_ ( .D(n247), .CK(clk), .RN(rstn), .Q(memory[199])
         );
  DFFRHQX1 memory_reg_3__6_ ( .D(n246), .CK(clk), .RN(rstn), .Q(memory[198])
         );
  DFFRHQX1 memory_reg_3__5_ ( .D(n245), .CK(clk), .RN(rstn), .Q(memory[197])
         );
  DFFRHQX1 memory_reg_3__4_ ( .D(n244), .CK(clk), .RN(rstn), .Q(memory[196])
         );
  DFFRHQX1 memory_reg_3__3_ ( .D(n243), .CK(clk), .RN(rstn), .Q(memory[195])
         );
  DFFRHQX1 memory_reg_3__2_ ( .D(n242), .CK(clk), .RN(rstn), .Q(memory[194])
         );
  DFFRHQX1 memory_reg_3__1_ ( .D(n241), .CK(clk), .RN(rstn), .Q(memory[193])
         );
  DFFRHQX1 memory_reg_3__0_ ( .D(n240), .CK(clk), .RN(rstn), .Q(memory[192])
         );
  DFFRHQX1 memory_reg_7__15_ ( .D(n191), .CK(clk), .RN(rstn), .Q(memory[143])
         );
  DFFRHQX1 memory_reg_7__14_ ( .D(n190), .CK(clk), .RN(rstn), .Q(memory[142])
         );
  DFFRHQX1 memory_reg_7__13_ ( .D(n189), .CK(clk), .RN(rstn), .Q(memory[141])
         );
  DFFRHQX1 memory_reg_7__12_ ( .D(n188), .CK(clk), .RN(rstn), .Q(memory[140])
         );
  DFFRHQX1 memory_reg_7__11_ ( .D(n187), .CK(clk), .RN(rstn), .Q(memory[139])
         );
  DFFRHQX1 memory_reg_7__10_ ( .D(n186), .CK(clk), .RN(rstn), .Q(memory[138])
         );
  DFFRHQX1 memory_reg_7__9_ ( .D(n185), .CK(clk), .RN(rstn), .Q(memory[137])
         );
  DFFRHQX1 memory_reg_7__8_ ( .D(n184), .CK(clk), .RN(rstn), .Q(memory[136])
         );
  DFFRHQX1 memory_reg_7__7_ ( .D(n183), .CK(clk), .RN(rstn), .Q(memory[135])
         );
  DFFRHQX1 memory_reg_7__6_ ( .D(n182), .CK(clk), .RN(rstn), .Q(memory[134])
         );
  DFFRHQX1 memory_reg_7__5_ ( .D(n181), .CK(clk), .RN(rstn), .Q(memory[133])
         );
  DFFRHQX1 memory_reg_7__4_ ( .D(n180), .CK(clk), .RN(rstn), .Q(memory[132])
         );
  DFFRHQX1 memory_reg_7__3_ ( .D(n179), .CK(clk), .RN(rstn), .Q(memory[131])
         );
  DFFRHQX1 memory_reg_7__2_ ( .D(n178), .CK(clk), .RN(rstn), .Q(memory[130])
         );
  DFFRHQX1 memory_reg_7__1_ ( .D(n177), .CK(clk), .RN(rstn), .Q(memory[129])
         );
  DFFRHQX1 memory_reg_7__0_ ( .D(n176), .CK(clk), .RN(rstn), .Q(memory[128])
         );
  DFFRHQX1 memory_reg_11__15_ ( .D(n127), .CK(clk), .RN(rstn), .Q(memory[79])
         );
  DFFRHQX1 memory_reg_11__14_ ( .D(n126), .CK(clk), .RN(rstn), .Q(memory[78])
         );
  DFFRHQX1 memory_reg_11__13_ ( .D(n125), .CK(clk), .RN(rstn), .Q(memory[77])
         );
  DFFRHQX1 memory_reg_11__12_ ( .D(n124), .CK(clk), .RN(rstn), .Q(memory[76])
         );
  DFFRHQX1 memory_reg_11__11_ ( .D(n123), .CK(clk), .RN(rstn), .Q(memory[75])
         );
  DFFRHQX1 memory_reg_11__10_ ( .D(n122), .CK(clk), .RN(rstn), .Q(memory[74])
         );
  DFFRHQX1 memory_reg_11__9_ ( .D(n121), .CK(clk), .RN(rstn), .Q(memory[73])
         );
  DFFRHQX1 memory_reg_11__8_ ( .D(n120), .CK(clk), .RN(rstn), .Q(memory[72])
         );
  DFFRHQX1 memory_reg_11__7_ ( .D(n119), .CK(clk), .RN(rstn), .Q(memory[71])
         );
  DFFRHQX1 memory_reg_11__6_ ( .D(n118), .CK(clk), .RN(rstn), .Q(memory[70])
         );
  DFFRHQX1 memory_reg_11__5_ ( .D(n117), .CK(clk), .RN(rstn), .Q(memory[69])
         );
  DFFRHQX1 memory_reg_11__4_ ( .D(n116), .CK(clk), .RN(rstn), .Q(memory[68])
         );
  DFFRHQX1 memory_reg_11__3_ ( .D(n115), .CK(clk), .RN(rstn), .Q(memory[67])
         );
  DFFRHQX1 memory_reg_11__2_ ( .D(n114), .CK(clk), .RN(rstn), .Q(memory[66])
         );
  DFFRHQX1 memory_reg_11__1_ ( .D(n113), .CK(clk), .RN(rstn), .Q(memory[65])
         );
  DFFRHQX1 memory_reg_11__0_ ( .D(n112), .CK(clk), .RN(rstn), .Q(memory[64])
         );
  DFFRHQX1 memory_reg_15__15_ ( .D(n63), .CK(clk), .RN(rstn), .Q(memory[15])
         );
  DFFRHQX1 memory_reg_15__14_ ( .D(n62), .CK(clk), .RN(rstn), .Q(memory[14])
         );
  DFFRHQX1 memory_reg_15__13_ ( .D(n61), .CK(clk), .RN(rstn), .Q(memory[13])
         );
  DFFRHQX1 memory_reg_15__12_ ( .D(n60), .CK(clk), .RN(rstn), .Q(memory[12])
         );
  DFFRHQX1 memory_reg_15__11_ ( .D(n59), .CK(clk), .RN(rstn), .Q(memory[11])
         );
  DFFRHQX1 memory_reg_15__10_ ( .D(n58), .CK(clk), .RN(rstn), .Q(memory[10])
         );
  DFFRHQX1 memory_reg_15__9_ ( .D(n57), .CK(clk), .RN(rstn), .Q(memory[9]) );
  DFFRHQX1 memory_reg_15__8_ ( .D(n56), .CK(clk), .RN(rstn), .Q(memory[8]) );
  DFFRHQX1 memory_reg_15__7_ ( .D(n55), .CK(clk), .RN(rstn), .Q(memory[7]) );
  DFFRHQX1 memory_reg_15__6_ ( .D(n54), .CK(clk), .RN(rstn), .Q(memory[6]) );
  DFFRHQX1 memory_reg_15__5_ ( .D(n53), .CK(clk), .RN(rstn), .Q(memory[5]) );
  DFFRHQX1 memory_reg_15__4_ ( .D(n52), .CK(clk), .RN(rstn), .Q(memory[4]) );
  DFFRHQX1 memory_reg_15__3_ ( .D(n51), .CK(clk), .RN(rstn), .Q(memory[3]) );
  DFFRHQX1 memory_reg_15__2_ ( .D(n50), .CK(clk), .RN(rstn), .Q(memory[2]) );
  DFFRHQX1 memory_reg_15__1_ ( .D(n49), .CK(clk), .RN(rstn), .Q(memory[1]) );
  DFFRHQX1 memory_reg_15__0_ ( .D(n48), .CK(clk), .RN(rstn), .Q(memory[0]) );
  DFFRHQX1 memory_reg_0__15_ ( .D(n303), .CK(clk), .RN(rstn), .Q(memory[255])
         );
  DFFRHQX1 memory_reg_0__14_ ( .D(n302), .CK(clk), .RN(rstn), .Q(memory[254])
         );
  DFFRHQX1 memory_reg_0__13_ ( .D(n301), .CK(clk), .RN(rstn), .Q(memory[253])
         );
  DFFRHQX1 memory_reg_0__12_ ( .D(n300), .CK(clk), .RN(rstn), .Q(memory[252])
         );
  DFFRHQX1 memory_reg_0__11_ ( .D(n299), .CK(clk), .RN(rstn), .Q(memory[251])
         );
  DFFRHQX1 memory_reg_0__10_ ( .D(n298), .CK(clk), .RN(rstn), .Q(memory[250])
         );
  DFFRHQX1 memory_reg_0__9_ ( .D(n297), .CK(clk), .RN(rstn), .Q(memory[249])
         );
  DFFRHQX1 memory_reg_0__8_ ( .D(n296), .CK(clk), .RN(rstn), .Q(memory[248])
         );
  DFFRHQX1 memory_reg_0__7_ ( .D(n295), .CK(clk), .RN(rstn), .Q(memory[247])
         );
  DFFRHQX1 memory_reg_0__6_ ( .D(n294), .CK(clk), .RN(rstn), .Q(memory[246])
         );
  DFFRHQX1 memory_reg_0__5_ ( .D(n293), .CK(clk), .RN(rstn), .Q(memory[245])
         );
  DFFRHQX1 memory_reg_0__4_ ( .D(n292), .CK(clk), .RN(rstn), .Q(memory[244])
         );
  DFFRHQX1 memory_reg_0__3_ ( .D(n291), .CK(clk), .RN(rstn), .Q(memory[243])
         );
  DFFRHQX1 memory_reg_0__2_ ( .D(n290), .CK(clk), .RN(rstn), .Q(memory[242])
         );
  DFFRHQX1 memory_reg_0__1_ ( .D(n289), .CK(clk), .RN(rstn), .Q(memory[241])
         );
  DFFRHQX1 memory_reg_0__0_ ( .D(n288), .CK(clk), .RN(rstn), .Q(memory[240])
         );
  DFFRHQX1 memory_reg_4__15_ ( .D(n239), .CK(clk), .RN(rstn), .Q(memory[191])
         );
  DFFRHQX1 memory_reg_4__14_ ( .D(n238), .CK(clk), .RN(rstn), .Q(memory[190])
         );
  DFFRHQX1 memory_reg_4__13_ ( .D(n237), .CK(clk), .RN(rstn), .Q(memory[189])
         );
  DFFRHQX1 memory_reg_4__12_ ( .D(n236), .CK(clk), .RN(rstn), .Q(memory[188])
         );
  DFFRHQX1 memory_reg_4__11_ ( .D(n235), .CK(clk), .RN(rstn), .Q(memory[187])
         );
  DFFRHQX1 memory_reg_4__10_ ( .D(n234), .CK(clk), .RN(rstn), .Q(memory[186])
         );
  DFFRHQX1 memory_reg_4__9_ ( .D(n233), .CK(clk), .RN(rstn), .Q(memory[185])
         );
  DFFRHQX1 memory_reg_4__8_ ( .D(n232), .CK(clk), .RN(rstn), .Q(memory[184])
         );
  DFFRHQX1 memory_reg_4__7_ ( .D(n231), .CK(clk), .RN(rstn), .Q(memory[183])
         );
  DFFRHQX1 memory_reg_4__6_ ( .D(n230), .CK(clk), .RN(rstn), .Q(memory[182])
         );
  DFFRHQX1 memory_reg_4__5_ ( .D(n229), .CK(clk), .RN(rstn), .Q(memory[181])
         );
  DFFRHQX1 memory_reg_4__4_ ( .D(n228), .CK(clk), .RN(rstn), .Q(memory[180])
         );
  DFFRHQX1 memory_reg_4__3_ ( .D(n227), .CK(clk), .RN(rstn), .Q(memory[179])
         );
  DFFRHQX1 memory_reg_4__2_ ( .D(n226), .CK(clk), .RN(rstn), .Q(memory[178])
         );
  DFFRHQX1 memory_reg_4__1_ ( .D(n225), .CK(clk), .RN(rstn), .Q(memory[177])
         );
  DFFRHQX1 memory_reg_4__0_ ( .D(n224), .CK(clk), .RN(rstn), .Q(memory[176])
         );
  DFFRHQX1 memory_reg_8__15_ ( .D(n175), .CK(clk), .RN(rstn), .Q(memory[127])
         );
  DFFRHQX1 memory_reg_8__14_ ( .D(n174), .CK(clk), .RN(rstn), .Q(memory[126])
         );
  DFFRHQX1 memory_reg_8__13_ ( .D(n173), .CK(clk), .RN(rstn), .Q(memory[125])
         );
  DFFRHQX1 memory_reg_8__12_ ( .D(n172), .CK(clk), .RN(rstn), .Q(memory[124])
         );
  DFFRHQX1 memory_reg_8__11_ ( .D(n171), .CK(clk), .RN(rstn), .Q(memory[123])
         );
  DFFRHQX1 memory_reg_8__10_ ( .D(n170), .CK(clk), .RN(rstn), .Q(memory[122])
         );
  DFFRHQX1 memory_reg_8__9_ ( .D(n169), .CK(clk), .RN(rstn), .Q(memory[121])
         );
  DFFRHQX1 memory_reg_8__8_ ( .D(n168), .CK(clk), .RN(rstn), .Q(memory[120])
         );
  DFFRHQX1 memory_reg_8__7_ ( .D(n167), .CK(clk), .RN(rstn), .Q(memory[119])
         );
  DFFRHQX1 memory_reg_8__6_ ( .D(n166), .CK(clk), .RN(rstn), .Q(memory[118])
         );
  DFFRHQX1 memory_reg_8__5_ ( .D(n165), .CK(clk), .RN(rstn), .Q(memory[117])
         );
  DFFRHQX1 memory_reg_8__4_ ( .D(n164), .CK(clk), .RN(rstn), .Q(memory[116])
         );
  DFFRHQX1 memory_reg_8__3_ ( .D(n163), .CK(clk), .RN(rstn), .Q(memory[115])
         );
  DFFRHQX1 memory_reg_8__2_ ( .D(n162), .CK(clk), .RN(rstn), .Q(memory[114])
         );
  DFFRHQX1 memory_reg_8__1_ ( .D(n161), .CK(clk), .RN(rstn), .Q(memory[113])
         );
  DFFRHQX1 memory_reg_8__0_ ( .D(n160), .CK(clk), .RN(rstn), .Q(memory[112])
         );
  DFFRHQX1 memory_reg_12__15_ ( .D(n111), .CK(clk), .RN(rstn), .Q(memory[63])
         );
  DFFRHQX1 memory_reg_12__14_ ( .D(n110), .CK(clk), .RN(rstn), .Q(memory[62])
         );
  DFFRHQX1 memory_reg_12__13_ ( .D(n109), .CK(clk), .RN(rstn), .Q(memory[61])
         );
  DFFRHQX1 memory_reg_12__12_ ( .D(n108), .CK(clk), .RN(rstn), .Q(memory[60])
         );
  DFFRHQX1 memory_reg_12__11_ ( .D(n107), .CK(clk), .RN(rstn), .Q(memory[59])
         );
  DFFRHQX1 memory_reg_12__10_ ( .D(n106), .CK(clk), .RN(rstn), .Q(memory[58])
         );
  DFFRHQX1 memory_reg_12__9_ ( .D(n105), .CK(clk), .RN(rstn), .Q(memory[57])
         );
  DFFRHQX1 memory_reg_12__8_ ( .D(n104), .CK(clk), .RN(rstn), .Q(memory[56])
         );
  DFFRHQX1 memory_reg_12__7_ ( .D(n103), .CK(clk), .RN(rstn), .Q(memory[55])
         );
  DFFRHQX1 memory_reg_12__6_ ( .D(n102), .CK(clk), .RN(rstn), .Q(memory[54])
         );
  DFFRHQX1 memory_reg_12__5_ ( .D(n101), .CK(clk), .RN(rstn), .Q(memory[53])
         );
  DFFRHQX1 memory_reg_12__4_ ( .D(n100), .CK(clk), .RN(rstn), .Q(memory[52])
         );
  DFFRHQX1 memory_reg_12__3_ ( .D(n99), .CK(clk), .RN(rstn), .Q(memory[51]) );
  DFFRHQX1 memory_reg_12__2_ ( .D(n98), .CK(clk), .RN(rstn), .Q(memory[50]) );
  DFFRHQX1 memory_reg_12__1_ ( .D(n97), .CK(clk), .RN(rstn), .Q(memory[49]) );
  DFFRHQX1 memory_reg_12__0_ ( .D(n96), .CK(clk), .RN(rstn), .Q(memory[48]) );
  DFFRHQX1 memory_reg_2__15_ ( .D(n271), .CK(clk), .RN(rstn), .Q(memory[223])
         );
  DFFRHQX1 memory_reg_2__14_ ( .D(n270), .CK(clk), .RN(rstn), .Q(memory[222])
         );
  DFFRHQX1 memory_reg_2__13_ ( .D(n269), .CK(clk), .RN(rstn), .Q(memory[221])
         );
  DFFRHQX1 memory_reg_2__12_ ( .D(n268), .CK(clk), .RN(rstn), .Q(memory[220])
         );
  DFFRHQX1 memory_reg_2__11_ ( .D(n267), .CK(clk), .RN(rstn), .Q(memory[219])
         );
  DFFRHQX1 memory_reg_2__10_ ( .D(n266), .CK(clk), .RN(rstn), .Q(memory[218])
         );
  DFFRHQX1 memory_reg_2__9_ ( .D(n265), .CK(clk), .RN(rstn), .Q(memory[217])
         );
  DFFRHQX1 memory_reg_2__8_ ( .D(n264), .CK(clk), .RN(rstn), .Q(memory[216])
         );
  DFFRHQX1 memory_reg_2__7_ ( .D(n263), .CK(clk), .RN(rstn), .Q(memory[215])
         );
  DFFRHQX1 memory_reg_2__6_ ( .D(n262), .CK(clk), .RN(rstn), .Q(memory[214])
         );
  DFFRHQX1 memory_reg_2__5_ ( .D(n261), .CK(clk), .RN(rstn), .Q(memory[213])
         );
  DFFRHQX1 memory_reg_2__4_ ( .D(n260), .CK(clk), .RN(rstn), .Q(memory[212])
         );
  DFFRHQX1 memory_reg_2__3_ ( .D(n259), .CK(clk), .RN(rstn), .Q(memory[211])
         );
  DFFRHQX1 memory_reg_2__2_ ( .D(n258), .CK(clk), .RN(rstn), .Q(memory[210])
         );
  DFFRHQX1 memory_reg_2__1_ ( .D(n257), .CK(clk), .RN(rstn), .Q(memory[209])
         );
  DFFRHQX1 memory_reg_2__0_ ( .D(n256), .CK(clk), .RN(rstn), .Q(memory[208])
         );
  DFFRHQX1 memory_reg_6__15_ ( .D(n207), .CK(clk), .RN(rstn), .Q(memory[159])
         );
  DFFRHQX1 memory_reg_6__14_ ( .D(n206), .CK(clk), .RN(rstn), .Q(memory[158])
         );
  DFFRHQX1 memory_reg_6__13_ ( .D(n205), .CK(clk), .RN(rstn), .Q(memory[157])
         );
  DFFRHQX1 memory_reg_6__12_ ( .D(n204), .CK(clk), .RN(rstn), .Q(memory[156])
         );
  DFFRHQX1 memory_reg_6__11_ ( .D(n203), .CK(clk), .RN(rstn), .Q(memory[155])
         );
  DFFRHQX1 memory_reg_6__10_ ( .D(n202), .CK(clk), .RN(rstn), .Q(memory[154])
         );
  DFFRHQX1 memory_reg_6__9_ ( .D(n201), .CK(clk), .RN(rstn), .Q(memory[153])
         );
  DFFRHQX1 memory_reg_6__8_ ( .D(n200), .CK(clk), .RN(rstn), .Q(memory[152])
         );
  DFFRHQX1 memory_reg_6__7_ ( .D(n199), .CK(clk), .RN(rstn), .Q(memory[151])
         );
  DFFRHQX1 memory_reg_6__6_ ( .D(n198), .CK(clk), .RN(rstn), .Q(memory[150])
         );
  DFFRHQX1 memory_reg_6__5_ ( .D(n197), .CK(clk), .RN(rstn), .Q(memory[149])
         );
  DFFRHQX1 memory_reg_6__4_ ( .D(n196), .CK(clk), .RN(rstn), .Q(memory[148])
         );
  DFFRHQX1 memory_reg_6__3_ ( .D(n195), .CK(clk), .RN(rstn), .Q(memory[147])
         );
  DFFRHQX1 memory_reg_6__2_ ( .D(n194), .CK(clk), .RN(rstn), .Q(memory[146])
         );
  DFFRHQX1 memory_reg_6__1_ ( .D(n193), .CK(clk), .RN(rstn), .Q(memory[145])
         );
  DFFRHQX1 memory_reg_6__0_ ( .D(n192), .CK(clk), .RN(rstn), .Q(memory[144])
         );
  DFFRHQX1 memory_reg_10__15_ ( .D(n143), .CK(clk), .RN(rstn), .Q(memory[95])
         );
  DFFRHQX1 memory_reg_10__14_ ( .D(n142), .CK(clk), .RN(rstn), .Q(memory[94])
         );
  DFFRHQX1 memory_reg_10__13_ ( .D(n141), .CK(clk), .RN(rstn), .Q(memory[93])
         );
  DFFRHQX1 memory_reg_10__12_ ( .D(n140), .CK(clk), .RN(rstn), .Q(memory[92])
         );
  DFFRHQX1 memory_reg_10__11_ ( .D(n139), .CK(clk), .RN(rstn), .Q(memory[91])
         );
  DFFRHQX1 memory_reg_10__10_ ( .D(n138), .CK(clk), .RN(rstn), .Q(memory[90])
         );
  DFFRHQX1 memory_reg_10__9_ ( .D(n137), .CK(clk), .RN(rstn), .Q(memory[89])
         );
  DFFRHQX1 memory_reg_10__8_ ( .D(n136), .CK(clk), .RN(rstn), .Q(memory[88])
         );
  DFFRHQX1 memory_reg_10__7_ ( .D(n135), .CK(clk), .RN(rstn), .Q(memory[87])
         );
  DFFRHQX1 memory_reg_10__6_ ( .D(n134), .CK(clk), .RN(rstn), .Q(memory[86])
         );
  DFFRHQX1 memory_reg_10__5_ ( .D(n133), .CK(clk), .RN(rstn), .Q(memory[85])
         );
  DFFRHQX1 memory_reg_10__4_ ( .D(n132), .CK(clk), .RN(rstn), .Q(memory[84])
         );
  DFFRHQX1 memory_reg_10__3_ ( .D(n131), .CK(clk), .RN(rstn), .Q(memory[83])
         );
  DFFRHQX1 memory_reg_10__2_ ( .D(n130), .CK(clk), .RN(rstn), .Q(memory[82])
         );
  DFFRHQX1 memory_reg_10__1_ ( .D(n129), .CK(clk), .RN(rstn), .Q(memory[81])
         );
  DFFRHQX1 memory_reg_10__0_ ( .D(n128), .CK(clk), .RN(rstn), .Q(memory[80])
         );
  DFFRHQX1 memory_reg_14__15_ ( .D(n79), .CK(clk), .RN(rstn), .Q(memory[31])
         );
  DFFRHQX1 memory_reg_14__14_ ( .D(n78), .CK(clk), .RN(rstn), .Q(memory[30])
         );
  DFFRHQX1 memory_reg_14__13_ ( .D(n77), .CK(clk), .RN(rstn), .Q(memory[29])
         );
  DFFRHQX1 memory_reg_14__12_ ( .D(n76), .CK(clk), .RN(rstn), .Q(memory[28])
         );
  DFFRHQX1 memory_reg_14__11_ ( .D(n75), .CK(clk), .RN(rstn), .Q(memory[27])
         );
  DFFRHQX1 memory_reg_14__10_ ( .D(n74), .CK(clk), .RN(rstn), .Q(memory[26])
         );
  DFFRHQX1 memory_reg_14__9_ ( .D(n73), .CK(clk), .RN(rstn), .Q(memory[25]) );
  DFFRHQX1 memory_reg_14__8_ ( .D(n72), .CK(clk), .RN(rstn), .Q(memory[24]) );
  DFFRHQX1 memory_reg_14__7_ ( .D(n71), .CK(clk), .RN(rstn), .Q(memory[23]) );
  DFFRHQX1 memory_reg_14__6_ ( .D(n70), .CK(clk), .RN(rstn), .Q(memory[22]) );
  DFFRHQX1 memory_reg_14__5_ ( .D(n69), .CK(clk), .RN(rstn), .Q(memory[21]) );
  DFFRHQX1 memory_reg_14__4_ ( .D(n68), .CK(clk), .RN(rstn), .Q(memory[20]) );
  DFFRHQX1 memory_reg_14__3_ ( .D(n67), .CK(clk), .RN(rstn), .Q(memory[19]) );
  DFFRHQX1 memory_reg_14__2_ ( .D(n66), .CK(clk), .RN(rstn), .Q(memory[18]) );
  DFFRHQX1 memory_reg_14__1_ ( .D(n65), .CK(clk), .RN(rstn), .Q(memory[17]) );
  DFFRHQX1 memory_reg_14__0_ ( .D(n64), .CK(clk), .RN(rstn), .Q(memory[16]) );
  INVXL U2 ( .A(addr[0]), .Y(n351) );
  NAND2X1 U3 ( .A(n21), .B(n22), .Y(n1) );
  NAND2X1 U4 ( .A(n24), .B(n21), .Y(n2) );
  NAND2X1 U5 ( .A(n26), .B(n22), .Y(n3) );
  NAND2X1 U6 ( .A(n26), .B(n24), .Y(n4) );
  NAND2X1 U7 ( .A(n29), .B(n22), .Y(n5) );
  NAND2X1 U8 ( .A(n29), .B(n24), .Y(n6) );
  NAND2X1 U9 ( .A(n32), .B(n22), .Y(n7) );
  NAND2X1 U10 ( .A(n32), .B(n24), .Y(n8) );
  NAND2X1 U11 ( .A(n37), .B(n21), .Y(n9) );
  NAND2X1 U12 ( .A(n39), .B(n21), .Y(n10) );
  NAND2X1 U13 ( .A(n37), .B(n26), .Y(n11) );
  NAND2X1 U14 ( .A(n39), .B(n26), .Y(n12) );
  NAND2X1 U15 ( .A(n37), .B(n29), .Y(n13) );
  NAND2X1 U16 ( .A(n39), .B(n29), .Y(n14) );
  NAND2X1 U17 ( .A(n37), .B(n32), .Y(n15) );
  NAND2X1 U18 ( .A(n39), .B(n32), .Y(n16) );
  INVX1 U19 ( .A(n351), .Y(n352) );
  INVX1 U20 ( .A(n351), .Y(n353) );
  INVX1 U21 ( .A(n351), .Y(n354) );
  INVX1 U22 ( .A(n358), .Y(n349) );
  INVX1 U23 ( .A(n358), .Y(n350) );
  NOR2X1 U24 ( .A(n359), .B(addr[1]), .Y(n26) );
  NOR2X1 U25 ( .A(n359), .B(n358), .Y(n21) );
  AND2X2 U26 ( .A(n45), .B(addr[0]), .Y(n37) );
  AND2X2 U27 ( .A(n45), .B(n351), .Y(n39) );
  AND2X2 U28 ( .A(n33), .B(n351), .Y(n24) );
  AND2X2 U29 ( .A(n33), .B(n353), .Y(n22) );
  MX4X1 U30 ( .A(memory[176]), .B(memory[160]), .C(memory[144]), .D(
        memory[128]), .S0(n353), .S1(n349), .Y(n19) );
  MX4X1 U31 ( .A(memory[177]), .B(memory[161]), .C(memory[145]), .D(
        memory[129]), .S0(n352), .S1(n349), .Y(n27) );
  MX4X1 U32 ( .A(memory[178]), .B(memory[162]), .C(memory[146]), .D(
        memory[130]), .S0(n352), .S1(n349), .Y(n34) );
  MX4X1 U33 ( .A(memory[179]), .B(memory[163]), .C(memory[147]), .D(
        memory[131]), .S0(n352), .S1(n349), .Y(n41) );
  MX4X1 U34 ( .A(memory[180]), .B(memory[164]), .C(memory[148]), .D(
        memory[132]), .S0(n353), .S1(n350), .Y(n46) );
  MX4X1 U35 ( .A(memory[181]), .B(memory[165]), .C(memory[149]), .D(
        memory[133]), .S0(n353), .S1(n350), .Y(n307) );
  MX4X1 U36 ( .A(memory[182]), .B(memory[166]), .C(memory[150]), .D(
        memory[134]), .S0(n353), .S1(n350), .Y(n311) );
  MX4X1 U37 ( .A(memory[183]), .B(memory[167]), .C(memory[151]), .D(
        memory[135]), .S0(n352), .S1(n350), .Y(n315) );
  MX4X1 U38 ( .A(memory[184]), .B(memory[168]), .C(memory[152]), .D(
        memory[136]), .S0(n354), .S1(n349), .Y(n319) );
  MX4X1 U39 ( .A(memory[185]), .B(memory[169]), .C(memory[153]), .D(
        memory[137]), .S0(n353), .S1(n350), .Y(n323) );
  MX4X1 U40 ( .A(memory[186]), .B(memory[170]), .C(memory[154]), .D(
        memory[138]), .S0(n354), .S1(n350), .Y(n327) );
  MX4X1 U41 ( .A(memory[187]), .B(memory[171]), .C(memory[155]), .D(
        memory[139]), .S0(n354), .S1(addr[1]), .Y(n331) );
  MX4X1 U42 ( .A(memory[188]), .B(memory[172]), .C(memory[156]), .D(
        memory[140]), .S0(n354), .S1(addr[1]), .Y(n335) );
  MX4X1 U43 ( .A(memory[189]), .B(memory[173]), .C(memory[157]), .D(
        memory[141]), .S0(n354), .S1(addr[1]), .Y(n339) );
  MX4X1 U44 ( .A(memory[190]), .B(memory[174]), .C(memory[158]), .D(
        memory[142]), .S0(n353), .S1(addr[1]), .Y(n343) );
  MX4X1 U45 ( .A(memory[191]), .B(memory[175]), .C(memory[159]), .D(
        memory[143]), .S0(addr[0]), .S1(addr[1]), .Y(n347) );
  MX4X1 U46 ( .A(memory[48]), .B(memory[32]), .C(memory[16]), .D(memory[0]), 
        .S0(n352), .S1(n350), .Y(n17) );
  MX4X1 U47 ( .A(memory[49]), .B(memory[33]), .C(memory[17]), .D(memory[1]), 
        .S0(n352), .S1(n349), .Y(n23) );
  MX4X1 U48 ( .A(memory[50]), .B(memory[34]), .C(memory[18]), .D(memory[2]), 
        .S0(n352), .S1(n349), .Y(n30) );
  MX4X1 U49 ( .A(memory[51]), .B(memory[35]), .C(memory[19]), .D(memory[3]), 
        .S0(n352), .S1(n349), .Y(n38) );
  MX4X1 U50 ( .A(memory[52]), .B(memory[36]), .C(memory[20]), .D(memory[4]), 
        .S0(n353), .S1(n350), .Y(n43) );
  MX4X1 U51 ( .A(memory[53]), .B(memory[37]), .C(memory[21]), .D(memory[5]), 
        .S0(n353), .S1(n350), .Y(n305) );
  MX4X1 U52 ( .A(memory[54]), .B(memory[38]), .C(memory[22]), .D(memory[6]), 
        .S0(n353), .S1(n350), .Y(n309) );
  MX4X1 U53 ( .A(memory[55]), .B(memory[39]), .C(memory[23]), .D(memory[7]), 
        .S0(n354), .S1(n349), .Y(n313) );
  MX4X1 U54 ( .A(memory[56]), .B(memory[40]), .C(memory[24]), .D(memory[8]), 
        .S0(n353), .S1(n349), .Y(n317) );
  MX4X1 U55 ( .A(memory[57]), .B(memory[41]), .C(memory[25]), .D(memory[9]), 
        .S0(addr[0]), .S1(n350), .Y(n321) );
  MX4X1 U56 ( .A(memory[58]), .B(memory[42]), .C(memory[26]), .D(memory[10]), 
        .S0(n354), .S1(n350), .Y(n325) );
  MX4X1 U57 ( .A(memory[59]), .B(memory[43]), .C(memory[27]), .D(memory[11]), 
        .S0(n354), .S1(n349), .Y(n329) );
  MX4X1 U58 ( .A(memory[60]), .B(memory[44]), .C(memory[28]), .D(memory[12]), 
        .S0(n354), .S1(n349), .Y(n333) );
  MX4X1 U59 ( .A(memory[61]), .B(memory[45]), .C(memory[29]), .D(memory[13]), 
        .S0(n352), .S1(n349), .Y(n337) );
  MX4X1 U60 ( .A(memory[62]), .B(memory[46]), .C(memory[30]), .D(memory[14]), 
        .S0(n352), .S1(n350), .Y(n341) );
  MX4X1 U61 ( .A(memory[63]), .B(memory[47]), .C(memory[31]), .D(memory[15]), 
        .S0(addr[0]), .S1(addr[1]), .Y(n345) );
  NOR2BX1 U62 ( .AN(N50), .B(n357), .Y(dout[0]) );
  MX4X1 U63 ( .A(n20), .B(n18), .C(n19), .D(n17), .S0(n356), .S1(n355), .Y(N50) );
  MX4X1 U64 ( .A(memory[240]), .B(memory[224]), .C(memory[208]), .D(
        memory[192]), .S0(n354), .S1(addr[1]), .Y(n20) );
  MX4X1 U65 ( .A(memory[112]), .B(memory[96]), .C(memory[80]), .D(memory[64]), 
        .S0(n352), .S1(n349), .Y(n18) );
  NOR2BX1 U66 ( .AN(N49), .B(n357), .Y(dout[1]) );
  MX4X1 U67 ( .A(n28), .B(n25), .C(n27), .D(n23), .S0(n356), .S1(n355), .Y(N49) );
  MX4X1 U68 ( .A(memory[241]), .B(memory[225]), .C(memory[209]), .D(
        memory[193]), .S0(n352), .S1(n349), .Y(n28) );
  MX4X1 U69 ( .A(memory[113]), .B(memory[97]), .C(memory[81]), .D(memory[65]), 
        .S0(n352), .S1(n349), .Y(n25) );
  NOR2BX1 U70 ( .AN(N48), .B(n357), .Y(dout[2]) );
  MX4X1 U71 ( .A(n36), .B(n31), .C(n34), .D(n30), .S0(n356), .S1(n355), .Y(N48) );
  MX4X1 U72 ( .A(memory[242]), .B(memory[226]), .C(memory[210]), .D(
        memory[194]), .S0(n352), .S1(n349), .Y(n36) );
  MX4X1 U73 ( .A(memory[114]), .B(memory[98]), .C(memory[82]), .D(memory[66]), 
        .S0(n352), .S1(n349), .Y(n31) );
  NOR2BX1 U74 ( .AN(N47), .B(n357), .Y(dout[3]) );
  MX4X1 U75 ( .A(n42), .B(n40), .C(n41), .D(n38), .S0(n356), .S1(n355), .Y(N47) );
  MX4X1 U76 ( .A(memory[243]), .B(memory[227]), .C(memory[211]), .D(
        memory[195]), .S0(n352), .S1(n349), .Y(n42) );
  MX4X1 U77 ( .A(memory[115]), .B(memory[99]), .C(memory[83]), .D(memory[67]), 
        .S0(n352), .S1(n349), .Y(n40) );
  NOR2BX1 U78 ( .AN(N46), .B(n357), .Y(dout[4]) );
  MX4X1 U79 ( .A(n304), .B(n44), .C(n46), .D(n43), .S0(n356), .S1(n355), .Y(
        N46) );
  MX4X1 U80 ( .A(memory[244]), .B(memory[228]), .C(memory[212]), .D(
        memory[196]), .S0(n353), .S1(n350), .Y(n304) );
  MX4X1 U81 ( .A(memory[116]), .B(memory[100]), .C(memory[84]), .D(memory[68]), 
        .S0(n353), .S1(n350), .Y(n44) );
  NOR2BX1 U82 ( .AN(N45), .B(n357), .Y(dout[5]) );
  MX4X1 U83 ( .A(n308), .B(n306), .C(n307), .D(n305), .S0(n356), .S1(n355), 
        .Y(N45) );
  MX4X1 U84 ( .A(memory[245]), .B(memory[229]), .C(memory[213]), .D(
        memory[197]), .S0(n353), .S1(n350), .Y(n308) );
  MX4X1 U85 ( .A(memory[117]), .B(memory[101]), .C(memory[85]), .D(memory[69]), 
        .S0(n353), .S1(n350), .Y(n306) );
  NOR2BX1 U86 ( .AN(N44), .B(n357), .Y(dout[6]) );
  MX4X1 U87 ( .A(n312), .B(n310), .C(n311), .D(n309), .S0(n356), .S1(n355), 
        .Y(N44) );
  MX4X1 U88 ( .A(memory[246]), .B(memory[230]), .C(memory[214]), .D(
        memory[198]), .S0(n353), .S1(n350), .Y(n312) );
  MX4X1 U89 ( .A(memory[118]), .B(memory[102]), .C(memory[86]), .D(memory[70]), 
        .S0(n353), .S1(n350), .Y(n310) );
  NOR2BX1 U90 ( .AN(N43), .B(n357), .Y(dout[7]) );
  MX4X1 U91 ( .A(n316), .B(n314), .C(n315), .D(n313), .S0(n356), .S1(n355), 
        .Y(N43) );
  MX4X1 U92 ( .A(memory[247]), .B(memory[231]), .C(memory[215]), .D(
        memory[199]), .S0(n354), .S1(n349), .Y(n316) );
  MX4X1 U93 ( .A(memory[119]), .B(memory[103]), .C(memory[87]), .D(memory[71]), 
        .S0(n354), .S1(n350), .Y(n314) );
  NOR2BX1 U94 ( .AN(N42), .B(n357), .Y(dout[8]) );
  MX4X1 U95 ( .A(n320), .B(n318), .C(n319), .D(n317), .S0(n356), .S1(n355), 
        .Y(N42) );
  MX4X1 U96 ( .A(memory[248]), .B(memory[232]), .C(memory[216]), .D(
        memory[200]), .S0(addr[0]), .S1(n350), .Y(n320) );
  MX4X1 U97 ( .A(memory[120]), .B(memory[104]), .C(memory[88]), .D(memory[72]), 
        .S0(n353), .S1(n350), .Y(n318) );
  NOR2BX1 U98 ( .AN(N41), .B(n357), .Y(dout[9]) );
  MX4X1 U99 ( .A(n324), .B(n322), .C(n323), .D(n321), .S0(n356), .S1(n355), 
        .Y(N41) );
  MX4X1 U100 ( .A(memory[249]), .B(memory[233]), .C(memory[217]), .D(
        memory[201]), .S0(addr[0]), .S1(n349), .Y(n324) );
  MX4X1 U101 ( .A(memory[121]), .B(memory[105]), .C(memory[89]), .D(memory[73]), .S0(n352), .S1(n349), .Y(n322) );
  NOR2BX1 U102 ( .AN(N40), .B(n357), .Y(dout[10]) );
  MX4X1 U103 ( .A(n328), .B(n326), .C(n327), .D(n325), .S0(n356), .S1(n355), 
        .Y(N40) );
  MX4X1 U104 ( .A(memory[250]), .B(memory[234]), .C(memory[218]), .D(
        memory[202]), .S0(n354), .S1(addr[1]), .Y(n328) );
  MX4X1 U105 ( .A(memory[122]), .B(memory[106]), .C(memory[90]), .D(memory[74]), .S0(n354), .S1(addr[1]), .Y(n326) );
  NOR2BX1 U106 ( .AN(N39), .B(n357), .Y(dout[11]) );
  MX4X1 U107 ( .A(n332), .B(n330), .C(n331), .D(n329), .S0(n356), .S1(n355), 
        .Y(N39) );
  MX4X1 U108 ( .A(memory[251]), .B(memory[235]), .C(memory[219]), .D(
        memory[203]), .S0(n354), .S1(addr[1]), .Y(n332) );
  MX4X1 U109 ( .A(memory[123]), .B(memory[107]), .C(memory[91]), .D(memory[75]), .S0(n354), .S1(addr[1]), .Y(n330) );
  NOR2BX1 U110 ( .AN(N38), .B(n357), .Y(dout[12]) );
  MX4X1 U111 ( .A(n336), .B(n334), .C(n335), .D(n333), .S0(n356), .S1(n355), 
        .Y(N38) );
  MX4X1 U112 ( .A(memory[252]), .B(memory[236]), .C(memory[220]), .D(
        memory[204]), .S0(n354), .S1(addr[1]), .Y(n336) );
  MX4X1 U113 ( .A(memory[124]), .B(memory[108]), .C(memory[92]), .D(memory[76]), .S0(n354), .S1(addr[1]), .Y(n334) );
  NOR2BX1 U114 ( .AN(N37), .B(n357), .Y(dout[13]) );
  MX4X1 U115 ( .A(n340), .B(n338), .C(n339), .D(n337), .S0(n356), .S1(n355), 
        .Y(N37) );
  MX4X1 U116 ( .A(memory[253]), .B(memory[237]), .C(memory[221]), .D(
        memory[205]), .S0(addr[0]), .S1(addr[1]), .Y(n340) );
  MX4X1 U117 ( .A(memory[125]), .B(memory[109]), .C(memory[93]), .D(memory[77]), .S0(addr[0]), .S1(addr[1]), .Y(n338) );
  NOR2BX1 U118 ( .AN(N36), .B(n357), .Y(dout[14]) );
  MX4X1 U119 ( .A(n344), .B(n342), .C(n343), .D(n341), .S0(n356), .S1(n355), 
        .Y(N36) );
  MX4X1 U120 ( .A(memory[254]), .B(memory[238]), .C(memory[222]), .D(
        memory[206]), .S0(addr[0]), .S1(addr[1]), .Y(n344) );
  MX4X1 U121 ( .A(memory[126]), .B(memory[110]), .C(memory[94]), .D(memory[78]), .S0(addr[0]), .S1(addr[1]), .Y(n342) );
  NOR2BX1 U122 ( .AN(N35), .B(n357), .Y(dout[15]) );
  MX4X1 U123 ( .A(n348), .B(n346), .C(n347), .D(n345), .S0(n356), .S1(n355), 
        .Y(N35) );
  MX4X1 U124 ( .A(memory[255]), .B(memory[239]), .C(memory[223]), .D(
        memory[207]), .S0(addr[0]), .S1(addr[1]), .Y(n348) );
  MX4X1 U125 ( .A(memory[127]), .B(memory[111]), .C(memory[95]), .D(memory[79]), .S0(addr[0]), .S1(addr[1]), .Y(n346) );
  INVX1 U126 ( .A(addr[1]), .Y(n358) );
  NOR2X1 U127 ( .A(n358), .B(addr[2]), .Y(n29) );
  NOR2X1 U128 ( .A(addr[1]), .B(addr[2]), .Y(n32) );
  BUFX3 U129 ( .A(addr[3]), .Y(n356) );
  OAI2BB2X1 U130 ( .B0(n1), .B1(n375), .A0N(memory[0]), .A1N(n1), .Y(n48) );
  OAI2BB2X1 U131 ( .B0(n1), .B1(n374), .A0N(memory[1]), .A1N(n1), .Y(n49) );
  OAI2BB2X1 U132 ( .B0(n1), .B1(n373), .A0N(memory[2]), .A1N(n1), .Y(n50) );
  OAI2BB2X1 U133 ( .B0(n1), .B1(n372), .A0N(memory[3]), .A1N(n1), .Y(n51) );
  OAI2BB2X1 U134 ( .B0(n1), .B1(n371), .A0N(memory[4]), .A1N(n1), .Y(n52) );
  OAI2BB2X1 U135 ( .B0(n1), .B1(n370), .A0N(memory[5]), .A1N(n1), .Y(n53) );
  OAI2BB2X1 U136 ( .B0(n1), .B1(n369), .A0N(memory[6]), .A1N(n1), .Y(n54) );
  OAI2BB2X1 U137 ( .B0(n1), .B1(n368), .A0N(memory[7]), .A1N(n1), .Y(n55) );
  OAI2BB2X1 U138 ( .B0(n1), .B1(n367), .A0N(memory[8]), .A1N(n1), .Y(n56) );
  OAI2BB2X1 U139 ( .B0(n1), .B1(n366), .A0N(memory[9]), .A1N(n1), .Y(n57) );
  OAI2BB2X1 U140 ( .B0(n1), .B1(n365), .A0N(memory[10]), .A1N(n1), .Y(n58) );
  OAI2BB2X1 U141 ( .B0(n1), .B1(n364), .A0N(memory[11]), .A1N(n1), .Y(n59) );
  OAI2BB2X1 U142 ( .B0(n1), .B1(n363), .A0N(memory[12]), .A1N(n1), .Y(n60) );
  OAI2BB2X1 U143 ( .B0(n1), .B1(n362), .A0N(memory[13]), .A1N(n1), .Y(n61) );
  OAI2BB2X1 U144 ( .B0(n1), .B1(n361), .A0N(memory[14]), .A1N(n1), .Y(n62) );
  OAI2BB2X1 U145 ( .B0(n1), .B1(n360), .A0N(memory[15]), .A1N(n1), .Y(n63) );
  OAI2BB2X1 U146 ( .B0(n375), .B1(n2), .A0N(memory[16]), .A1N(n2), .Y(n64) );
  OAI2BB2X1 U147 ( .B0(n374), .B1(n2), .A0N(memory[17]), .A1N(n2), .Y(n65) );
  OAI2BB2X1 U148 ( .B0(n373), .B1(n2), .A0N(memory[18]), .A1N(n2), .Y(n66) );
  OAI2BB2X1 U149 ( .B0(n372), .B1(n2), .A0N(memory[19]), .A1N(n2), .Y(n67) );
  OAI2BB2X1 U150 ( .B0(n371), .B1(n2), .A0N(memory[20]), .A1N(n2), .Y(n68) );
  OAI2BB2X1 U151 ( .B0(n370), .B1(n2), .A0N(memory[21]), .A1N(n2), .Y(n69) );
  OAI2BB2X1 U152 ( .B0(n369), .B1(n2), .A0N(memory[22]), .A1N(n2), .Y(n70) );
  OAI2BB2X1 U153 ( .B0(n368), .B1(n2), .A0N(memory[23]), .A1N(n2), .Y(n71) );
  OAI2BB2X1 U154 ( .B0(n363), .B1(n2), .A0N(memory[28]), .A1N(n2), .Y(n76) );
  OAI2BB2X1 U155 ( .B0(n362), .B1(n2), .A0N(memory[29]), .A1N(n2), .Y(n77) );
  OAI2BB2X1 U156 ( .B0(n361), .B1(n2), .A0N(memory[30]), .A1N(n2), .Y(n78) );
  OAI2BB2X1 U157 ( .B0(n360), .B1(n2), .A0N(memory[31]), .A1N(n2), .Y(n79) );
  OAI2BB2X1 U158 ( .B0(n375), .B1(n3), .A0N(memory[32]), .A1N(n3), .Y(n80) );
  OAI2BB2X1 U159 ( .B0(n374), .B1(n3), .A0N(memory[33]), .A1N(n3), .Y(n81) );
  OAI2BB2X1 U160 ( .B0(n373), .B1(n3), .A0N(memory[34]), .A1N(n3), .Y(n82) );
  OAI2BB2X1 U161 ( .B0(n372), .B1(n3), .A0N(memory[35]), .A1N(n3), .Y(n83) );
  OAI2BB2X1 U162 ( .B0(n371), .B1(n3), .A0N(memory[36]), .A1N(n3), .Y(n84) );
  OAI2BB2X1 U163 ( .B0(n370), .B1(n3), .A0N(memory[37]), .A1N(n3), .Y(n85) );
  OAI2BB2X1 U164 ( .B0(n369), .B1(n3), .A0N(memory[38]), .A1N(n3), .Y(n86) );
  OAI2BB2X1 U165 ( .B0(n368), .B1(n3), .A0N(memory[39]), .A1N(n3), .Y(n87) );
  OAI2BB2X1 U166 ( .B0(n363), .B1(n3), .A0N(memory[44]), .A1N(n3), .Y(n92) );
  OAI2BB2X1 U167 ( .B0(n362), .B1(n3), .A0N(memory[45]), .A1N(n3), .Y(n93) );
  OAI2BB2X1 U168 ( .B0(n361), .B1(n3), .A0N(memory[46]), .A1N(n3), .Y(n94) );
  OAI2BB2X1 U169 ( .B0(n360), .B1(n3), .A0N(memory[47]), .A1N(n3), .Y(n95) );
  OAI2BB2X1 U170 ( .B0(n375), .B1(n4), .A0N(memory[48]), .A1N(n4), .Y(n96) );
  OAI2BB2X1 U171 ( .B0(n374), .B1(n4), .A0N(memory[49]), .A1N(n4), .Y(n97) );
  OAI2BB2X1 U172 ( .B0(n373), .B1(n4), .A0N(memory[50]), .A1N(n4), .Y(n98) );
  OAI2BB2X1 U173 ( .B0(n372), .B1(n4), .A0N(memory[51]), .A1N(n4), .Y(n99) );
  OAI2BB2X1 U174 ( .B0(n371), .B1(n4), .A0N(memory[52]), .A1N(n4), .Y(n100) );
  OAI2BB2X1 U175 ( .B0(n370), .B1(n4), .A0N(memory[53]), .A1N(n4), .Y(n101) );
  OAI2BB2X1 U176 ( .B0(n369), .B1(n4), .A0N(memory[54]), .A1N(n4), .Y(n102) );
  OAI2BB2X1 U177 ( .B0(n368), .B1(n4), .A0N(memory[55]), .A1N(n4), .Y(n103) );
  OAI2BB2X1 U178 ( .B0(n363), .B1(n4), .A0N(memory[60]), .A1N(n4), .Y(n108) );
  OAI2BB2X1 U179 ( .B0(n362), .B1(n4), .A0N(memory[61]), .A1N(n4), .Y(n109) );
  OAI2BB2X1 U180 ( .B0(n361), .B1(n4), .A0N(memory[62]), .A1N(n4), .Y(n110) );
  OAI2BB2X1 U181 ( .B0(n360), .B1(n4), .A0N(memory[63]), .A1N(n4), .Y(n111) );
  OAI2BB2X1 U182 ( .B0(n375), .B1(n5), .A0N(memory[64]), .A1N(n5), .Y(n112) );
  OAI2BB2X1 U183 ( .B0(n374), .B1(n5), .A0N(memory[65]), .A1N(n5), .Y(n113) );
  OAI2BB2X1 U184 ( .B0(n373), .B1(n5), .A0N(memory[66]), .A1N(n5), .Y(n114) );
  OAI2BB2X1 U185 ( .B0(n372), .B1(n5), .A0N(memory[67]), .A1N(n5), .Y(n115) );
  OAI2BB2X1 U186 ( .B0(n371), .B1(n5), .A0N(memory[68]), .A1N(n5), .Y(n116) );
  OAI2BB2X1 U187 ( .B0(n370), .B1(n5), .A0N(memory[69]), .A1N(n5), .Y(n117) );
  OAI2BB2X1 U188 ( .B0(n369), .B1(n5), .A0N(memory[70]), .A1N(n5), .Y(n118) );
  OAI2BB2X1 U189 ( .B0(n368), .B1(n5), .A0N(memory[71]), .A1N(n5), .Y(n119) );
  OAI2BB2X1 U190 ( .B0(n363), .B1(n5), .A0N(memory[76]), .A1N(n5), .Y(n124) );
  OAI2BB2X1 U191 ( .B0(n362), .B1(n5), .A0N(memory[77]), .A1N(n5), .Y(n125) );
  OAI2BB2X1 U192 ( .B0(n361), .B1(n5), .A0N(memory[78]), .A1N(n5), .Y(n126) );
  OAI2BB2X1 U193 ( .B0(n360), .B1(n5), .A0N(memory[79]), .A1N(n5), .Y(n127) );
  OAI2BB2X1 U194 ( .B0(n375), .B1(n6), .A0N(memory[80]), .A1N(n6), .Y(n128) );
  OAI2BB2X1 U195 ( .B0(n374), .B1(n6), .A0N(memory[81]), .A1N(n6), .Y(n129) );
  OAI2BB2X1 U196 ( .B0(n373), .B1(n6), .A0N(memory[82]), .A1N(n6), .Y(n130) );
  OAI2BB2X1 U197 ( .B0(n372), .B1(n6), .A0N(memory[83]), .A1N(n6), .Y(n131) );
  OAI2BB2X1 U198 ( .B0(n371), .B1(n6), .A0N(memory[84]), .A1N(n6), .Y(n132) );
  OAI2BB2X1 U199 ( .B0(n370), .B1(n6), .A0N(memory[85]), .A1N(n6), .Y(n133) );
  OAI2BB2X1 U200 ( .B0(n369), .B1(n6), .A0N(memory[86]), .A1N(n6), .Y(n134) );
  OAI2BB2X1 U201 ( .B0(n368), .B1(n6), .A0N(memory[87]), .A1N(n6), .Y(n135) );
  OAI2BB2X1 U202 ( .B0(n363), .B1(n6), .A0N(memory[92]), .A1N(n6), .Y(n140) );
  OAI2BB2X1 U203 ( .B0(n362), .B1(n6), .A0N(memory[93]), .A1N(n6), .Y(n141) );
  OAI2BB2X1 U204 ( .B0(n361), .B1(n6), .A0N(memory[94]), .A1N(n6), .Y(n142) );
  OAI2BB2X1 U205 ( .B0(n360), .B1(n6), .A0N(memory[95]), .A1N(n6), .Y(n143) );
  OAI2BB2X1 U206 ( .B0(n375), .B1(n7), .A0N(memory[96]), .A1N(n7), .Y(n144) );
  OAI2BB2X1 U207 ( .B0(n374), .B1(n7), .A0N(memory[97]), .A1N(n7), .Y(n145) );
  OAI2BB2X1 U208 ( .B0(n373), .B1(n7), .A0N(memory[98]), .A1N(n7), .Y(n146) );
  OAI2BB2X1 U209 ( .B0(n372), .B1(n7), .A0N(memory[99]), .A1N(n7), .Y(n147) );
  OAI2BB2X1 U210 ( .B0(n371), .B1(n7), .A0N(memory[100]), .A1N(n7), .Y(n148)
         );
  OAI2BB2X1 U211 ( .B0(n370), .B1(n7), .A0N(memory[101]), .A1N(n7), .Y(n149)
         );
  OAI2BB2X1 U212 ( .B0(n369), .B1(n7), .A0N(memory[102]), .A1N(n7), .Y(n150)
         );
  OAI2BB2X1 U213 ( .B0(n368), .B1(n7), .A0N(memory[103]), .A1N(n7), .Y(n151)
         );
  OAI2BB2X1 U214 ( .B0(n363), .B1(n7), .A0N(memory[108]), .A1N(n7), .Y(n156)
         );
  OAI2BB2X1 U215 ( .B0(n362), .B1(n7), .A0N(memory[109]), .A1N(n7), .Y(n157)
         );
  OAI2BB2X1 U216 ( .B0(n361), .B1(n7), .A0N(memory[110]), .A1N(n7), .Y(n158)
         );
  OAI2BB2X1 U217 ( .B0(n360), .B1(n7), .A0N(memory[111]), .A1N(n7), .Y(n159)
         );
  OAI2BB2X1 U218 ( .B0(n375), .B1(n8), .A0N(memory[112]), .A1N(n8), .Y(n160)
         );
  OAI2BB2X1 U219 ( .B0(n374), .B1(n8), .A0N(memory[113]), .A1N(n8), .Y(n161)
         );
  OAI2BB2X1 U220 ( .B0(n373), .B1(n8), .A0N(memory[114]), .A1N(n8), .Y(n162)
         );
  OAI2BB2X1 U221 ( .B0(n372), .B1(n8), .A0N(memory[115]), .A1N(n8), .Y(n163)
         );
  OAI2BB2X1 U222 ( .B0(n371), .B1(n8), .A0N(memory[116]), .A1N(n8), .Y(n164)
         );
  OAI2BB2X1 U223 ( .B0(n370), .B1(n8), .A0N(memory[117]), .A1N(n8), .Y(n165)
         );
  OAI2BB2X1 U224 ( .B0(n369), .B1(n8), .A0N(memory[118]), .A1N(n8), .Y(n166)
         );
  OAI2BB2X1 U225 ( .B0(n368), .B1(n8), .A0N(memory[119]), .A1N(n8), .Y(n167)
         );
  OAI2BB2X1 U226 ( .B0(n363), .B1(n8), .A0N(memory[124]), .A1N(n8), .Y(n172)
         );
  OAI2BB2X1 U227 ( .B0(n362), .B1(n8), .A0N(memory[125]), .A1N(n8), .Y(n173)
         );
  OAI2BB2X1 U228 ( .B0(n361), .B1(n8), .A0N(memory[126]), .A1N(n8), .Y(n174)
         );
  OAI2BB2X1 U229 ( .B0(n360), .B1(n8), .A0N(memory[127]), .A1N(n8), .Y(n175)
         );
  OAI2BB2X1 U230 ( .B0(n375), .B1(n9), .A0N(memory[128]), .A1N(n9), .Y(n176)
         );
  OAI2BB2X1 U231 ( .B0(n374), .B1(n9), .A0N(memory[129]), .A1N(n9), .Y(n177)
         );
  OAI2BB2X1 U232 ( .B0(n373), .B1(n9), .A0N(memory[130]), .A1N(n9), .Y(n178)
         );
  OAI2BB2X1 U233 ( .B0(n372), .B1(n9), .A0N(memory[131]), .A1N(n9), .Y(n179)
         );
  OAI2BB2X1 U234 ( .B0(n371), .B1(n9), .A0N(memory[132]), .A1N(n9), .Y(n180)
         );
  OAI2BB2X1 U235 ( .B0(n370), .B1(n9), .A0N(memory[133]), .A1N(n9), .Y(n181)
         );
  OAI2BB2X1 U236 ( .B0(n369), .B1(n9), .A0N(memory[134]), .A1N(n9), .Y(n182)
         );
  OAI2BB2X1 U237 ( .B0(n368), .B1(n9), .A0N(memory[135]), .A1N(n9), .Y(n183)
         );
  OAI2BB2X1 U238 ( .B0(n363), .B1(n9), .A0N(memory[140]), .A1N(n9), .Y(n188)
         );
  OAI2BB2X1 U239 ( .B0(n362), .B1(n9), .A0N(memory[141]), .A1N(n9), .Y(n189)
         );
  OAI2BB2X1 U240 ( .B0(n361), .B1(n9), .A0N(memory[142]), .A1N(n9), .Y(n190)
         );
  OAI2BB2X1 U241 ( .B0(n360), .B1(n9), .A0N(memory[143]), .A1N(n9), .Y(n191)
         );
  OAI2BB2X1 U242 ( .B0(n375), .B1(n10), .A0N(memory[144]), .A1N(n10), .Y(n192)
         );
  OAI2BB2X1 U243 ( .B0(n374), .B1(n10), .A0N(memory[145]), .A1N(n10), .Y(n193)
         );
  OAI2BB2X1 U244 ( .B0(n373), .B1(n10), .A0N(memory[146]), .A1N(n10), .Y(n194)
         );
  OAI2BB2X1 U245 ( .B0(n372), .B1(n10), .A0N(memory[147]), .A1N(n10), .Y(n195)
         );
  OAI2BB2X1 U246 ( .B0(n371), .B1(n10), .A0N(memory[148]), .A1N(n10), .Y(n196)
         );
  OAI2BB2X1 U247 ( .B0(n370), .B1(n10), .A0N(memory[149]), .A1N(n10), .Y(n197)
         );
  OAI2BB2X1 U248 ( .B0(n369), .B1(n10), .A0N(memory[150]), .A1N(n10), .Y(n198)
         );
  OAI2BB2X1 U249 ( .B0(n368), .B1(n10), .A0N(memory[151]), .A1N(n10), .Y(n199)
         );
  OAI2BB2X1 U250 ( .B0(n363), .B1(n10), .A0N(memory[156]), .A1N(n10), .Y(n204)
         );
  OAI2BB2X1 U251 ( .B0(n362), .B1(n10), .A0N(memory[157]), .A1N(n10), .Y(n205)
         );
  OAI2BB2X1 U252 ( .B0(n361), .B1(n10), .A0N(memory[158]), .A1N(n10), .Y(n206)
         );
  OAI2BB2X1 U253 ( .B0(n360), .B1(n10), .A0N(memory[159]), .A1N(n10), .Y(n207)
         );
  OAI2BB2X1 U254 ( .B0(n375), .B1(n11), .A0N(memory[160]), .A1N(n11), .Y(n208)
         );
  OAI2BB2X1 U255 ( .B0(n374), .B1(n11), .A0N(memory[161]), .A1N(n11), .Y(n209)
         );
  OAI2BB2X1 U256 ( .B0(n373), .B1(n11), .A0N(memory[162]), .A1N(n11), .Y(n210)
         );
  OAI2BB2X1 U257 ( .B0(n372), .B1(n11), .A0N(memory[163]), .A1N(n11), .Y(n211)
         );
  OAI2BB2X1 U258 ( .B0(n371), .B1(n11), .A0N(memory[164]), .A1N(n11), .Y(n212)
         );
  OAI2BB2X1 U259 ( .B0(n370), .B1(n11), .A0N(memory[165]), .A1N(n11), .Y(n213)
         );
  OAI2BB2X1 U260 ( .B0(n369), .B1(n11), .A0N(memory[166]), .A1N(n11), .Y(n214)
         );
  OAI2BB2X1 U261 ( .B0(n368), .B1(n11), .A0N(memory[167]), .A1N(n11), .Y(n215)
         );
  OAI2BB2X1 U262 ( .B0(n363), .B1(n11), .A0N(memory[172]), .A1N(n11), .Y(n220)
         );
  OAI2BB2X1 U263 ( .B0(n362), .B1(n11), .A0N(memory[173]), .A1N(n11), .Y(n221)
         );
  OAI2BB2X1 U264 ( .B0(n361), .B1(n11), .A0N(memory[174]), .A1N(n11), .Y(n222)
         );
  OAI2BB2X1 U265 ( .B0(n360), .B1(n11), .A0N(memory[175]), .A1N(n11), .Y(n223)
         );
  OAI2BB2X1 U266 ( .B0(n375), .B1(n12), .A0N(memory[176]), .A1N(n12), .Y(n224)
         );
  OAI2BB2X1 U267 ( .B0(n374), .B1(n12), .A0N(memory[177]), .A1N(n12), .Y(n225)
         );
  OAI2BB2X1 U268 ( .B0(n373), .B1(n12), .A0N(memory[178]), .A1N(n12), .Y(n226)
         );
  OAI2BB2X1 U269 ( .B0(n372), .B1(n12), .A0N(memory[179]), .A1N(n12), .Y(n227)
         );
  OAI2BB2X1 U270 ( .B0(n371), .B1(n12), .A0N(memory[180]), .A1N(n12), .Y(n228)
         );
  OAI2BB2X1 U271 ( .B0(n370), .B1(n12), .A0N(memory[181]), .A1N(n12), .Y(n229)
         );
  OAI2BB2X1 U272 ( .B0(n369), .B1(n12), .A0N(memory[182]), .A1N(n12), .Y(n230)
         );
  OAI2BB2X1 U273 ( .B0(n368), .B1(n12), .A0N(memory[183]), .A1N(n12), .Y(n231)
         );
  OAI2BB2X1 U274 ( .B0(n363), .B1(n12), .A0N(memory[188]), .A1N(n12), .Y(n236)
         );
  OAI2BB2X1 U275 ( .B0(n362), .B1(n12), .A0N(memory[189]), .A1N(n12), .Y(n237)
         );
  OAI2BB2X1 U276 ( .B0(n361), .B1(n12), .A0N(memory[190]), .A1N(n12), .Y(n238)
         );
  OAI2BB2X1 U277 ( .B0(n360), .B1(n12), .A0N(memory[191]), .A1N(n12), .Y(n239)
         );
  OAI2BB2X1 U278 ( .B0(n375), .B1(n13), .A0N(memory[192]), .A1N(n13), .Y(n240)
         );
  OAI2BB2X1 U279 ( .B0(n374), .B1(n13), .A0N(memory[193]), .A1N(n13), .Y(n241)
         );
  OAI2BB2X1 U280 ( .B0(n373), .B1(n13), .A0N(memory[194]), .A1N(n13), .Y(n242)
         );
  OAI2BB2X1 U281 ( .B0(n372), .B1(n13), .A0N(memory[195]), .A1N(n13), .Y(n243)
         );
  OAI2BB2X1 U282 ( .B0(n371), .B1(n13), .A0N(memory[196]), .A1N(n13), .Y(n244)
         );
  OAI2BB2X1 U283 ( .B0(n370), .B1(n13), .A0N(memory[197]), .A1N(n13), .Y(n245)
         );
  OAI2BB2X1 U284 ( .B0(n369), .B1(n13), .A0N(memory[198]), .A1N(n13), .Y(n246)
         );
  OAI2BB2X1 U285 ( .B0(n368), .B1(n13), .A0N(memory[199]), .A1N(n13), .Y(n247)
         );
  OAI2BB2X1 U286 ( .B0(n363), .B1(n13), .A0N(memory[204]), .A1N(n13), .Y(n252)
         );
  OAI2BB2X1 U287 ( .B0(n362), .B1(n13), .A0N(memory[205]), .A1N(n13), .Y(n253)
         );
  OAI2BB2X1 U288 ( .B0(n361), .B1(n13), .A0N(memory[206]), .A1N(n13), .Y(n254)
         );
  OAI2BB2X1 U289 ( .B0(n360), .B1(n13), .A0N(memory[207]), .A1N(n13), .Y(n255)
         );
  OAI2BB2X1 U290 ( .B0(n375), .B1(n14), .A0N(memory[208]), .A1N(n14), .Y(n256)
         );
  OAI2BB2X1 U291 ( .B0(n374), .B1(n14), .A0N(memory[209]), .A1N(n14), .Y(n257)
         );
  OAI2BB2X1 U292 ( .B0(n373), .B1(n14), .A0N(memory[210]), .A1N(n14), .Y(n258)
         );
  OAI2BB2X1 U293 ( .B0(n372), .B1(n14), .A0N(memory[211]), .A1N(n14), .Y(n259)
         );
  OAI2BB2X1 U294 ( .B0(n371), .B1(n14), .A0N(memory[212]), .A1N(n14), .Y(n260)
         );
  OAI2BB2X1 U295 ( .B0(n370), .B1(n14), .A0N(memory[213]), .A1N(n14), .Y(n261)
         );
  OAI2BB2X1 U296 ( .B0(n369), .B1(n14), .A0N(memory[214]), .A1N(n14), .Y(n262)
         );
  OAI2BB2X1 U297 ( .B0(n368), .B1(n14), .A0N(memory[215]), .A1N(n14), .Y(n263)
         );
  OAI2BB2X1 U298 ( .B0(n363), .B1(n14), .A0N(memory[220]), .A1N(n14), .Y(n268)
         );
  OAI2BB2X1 U299 ( .B0(n362), .B1(n14), .A0N(memory[221]), .A1N(n14), .Y(n269)
         );
  OAI2BB2X1 U300 ( .B0(n361), .B1(n14), .A0N(memory[222]), .A1N(n14), .Y(n270)
         );
  OAI2BB2X1 U301 ( .B0(n360), .B1(n14), .A0N(memory[223]), .A1N(n14), .Y(n271)
         );
  OAI2BB2X1 U302 ( .B0(n375), .B1(n15), .A0N(memory[224]), .A1N(n15), .Y(n272)
         );
  OAI2BB2X1 U303 ( .B0(n374), .B1(n15), .A0N(memory[225]), .A1N(n15), .Y(n273)
         );
  OAI2BB2X1 U304 ( .B0(n373), .B1(n15), .A0N(memory[226]), .A1N(n15), .Y(n274)
         );
  OAI2BB2X1 U305 ( .B0(n372), .B1(n15), .A0N(memory[227]), .A1N(n15), .Y(n275)
         );
  OAI2BB2X1 U306 ( .B0(n371), .B1(n15), .A0N(memory[228]), .A1N(n15), .Y(n276)
         );
  OAI2BB2X1 U307 ( .B0(n370), .B1(n15), .A0N(memory[229]), .A1N(n15), .Y(n277)
         );
  OAI2BB2X1 U308 ( .B0(n369), .B1(n15), .A0N(memory[230]), .A1N(n15), .Y(n278)
         );
  OAI2BB2X1 U309 ( .B0(n368), .B1(n15), .A0N(memory[231]), .A1N(n15), .Y(n279)
         );
  OAI2BB2X1 U310 ( .B0(n363), .B1(n15), .A0N(memory[236]), .A1N(n15), .Y(n284)
         );
  OAI2BB2X1 U311 ( .B0(n362), .B1(n15), .A0N(memory[237]), .A1N(n15), .Y(n285)
         );
  OAI2BB2X1 U312 ( .B0(n361), .B1(n15), .A0N(memory[238]), .A1N(n15), .Y(n286)
         );
  OAI2BB2X1 U313 ( .B0(n360), .B1(n15), .A0N(memory[239]), .A1N(n15), .Y(n287)
         );
  OAI2BB2X1 U314 ( .B0(n375), .B1(n16), .A0N(memory[240]), .A1N(n16), .Y(n288)
         );
  OAI2BB2X1 U315 ( .B0(n374), .B1(n16), .A0N(memory[241]), .A1N(n16), .Y(n289)
         );
  OAI2BB2X1 U316 ( .B0(n373), .B1(n16), .A0N(memory[242]), .A1N(n16), .Y(n290)
         );
  OAI2BB2X1 U317 ( .B0(n372), .B1(n16), .A0N(memory[243]), .A1N(n16), .Y(n291)
         );
  OAI2BB2X1 U318 ( .B0(n371), .B1(n16), .A0N(memory[244]), .A1N(n16), .Y(n292)
         );
  OAI2BB2X1 U319 ( .B0(n370), .B1(n16), .A0N(memory[245]), .A1N(n16), .Y(n293)
         );
  OAI2BB2X1 U320 ( .B0(n369), .B1(n16), .A0N(memory[246]), .A1N(n16), .Y(n294)
         );
  OAI2BB2X1 U321 ( .B0(n368), .B1(n16), .A0N(memory[247]), .A1N(n16), .Y(n295)
         );
  OAI2BB2X1 U322 ( .B0(n363), .B1(n16), .A0N(memory[252]), .A1N(n16), .Y(n300)
         );
  OAI2BB2X1 U323 ( .B0(n362), .B1(n16), .A0N(memory[253]), .A1N(n16), .Y(n301)
         );
  OAI2BB2X1 U324 ( .B0(n361), .B1(n16), .A0N(memory[254]), .A1N(n16), .Y(n302)
         );
  OAI2BB2X1 U325 ( .B0(n360), .B1(n16), .A0N(memory[255]), .A1N(n16), .Y(n303)
         );
  OAI2BB2X1 U326 ( .B0(n367), .B1(n2), .A0N(memory[24]), .A1N(n2), .Y(n72) );
  OAI2BB2X1 U327 ( .B0(n366), .B1(n2), .A0N(memory[25]), .A1N(n2), .Y(n73) );
  OAI2BB2X1 U328 ( .B0(n365), .B1(n2), .A0N(memory[26]), .A1N(n2), .Y(n74) );
  OAI2BB2X1 U329 ( .B0(n364), .B1(n2), .A0N(memory[27]), .A1N(n2), .Y(n75) );
  OAI2BB2X1 U330 ( .B0(n367), .B1(n3), .A0N(memory[40]), .A1N(n3), .Y(n88) );
  OAI2BB2X1 U331 ( .B0(n366), .B1(n3), .A0N(memory[41]), .A1N(n3), .Y(n89) );
  OAI2BB2X1 U332 ( .B0(n365), .B1(n3), .A0N(memory[42]), .A1N(n3), .Y(n90) );
  OAI2BB2X1 U333 ( .B0(n364), .B1(n3), .A0N(memory[43]), .A1N(n3), .Y(n91) );
  OAI2BB2X1 U334 ( .B0(n367), .B1(n4), .A0N(memory[56]), .A1N(n4), .Y(n104) );
  OAI2BB2X1 U335 ( .B0(n366), .B1(n4), .A0N(memory[57]), .A1N(n4), .Y(n105) );
  OAI2BB2X1 U336 ( .B0(n365), .B1(n4), .A0N(memory[58]), .A1N(n4), .Y(n106) );
  OAI2BB2X1 U337 ( .B0(n364), .B1(n4), .A0N(memory[59]), .A1N(n4), .Y(n107) );
  OAI2BB2X1 U338 ( .B0(n367), .B1(n5), .A0N(memory[72]), .A1N(n5), .Y(n120) );
  OAI2BB2X1 U339 ( .B0(n366), .B1(n5), .A0N(memory[73]), .A1N(n5), .Y(n121) );
  OAI2BB2X1 U340 ( .B0(n365), .B1(n5), .A0N(memory[74]), .A1N(n5), .Y(n122) );
  OAI2BB2X1 U341 ( .B0(n364), .B1(n5), .A0N(memory[75]), .A1N(n5), .Y(n123) );
  OAI2BB2X1 U342 ( .B0(n367), .B1(n6), .A0N(memory[88]), .A1N(n6), .Y(n136) );
  OAI2BB2X1 U343 ( .B0(n366), .B1(n6), .A0N(memory[89]), .A1N(n6), .Y(n137) );
  OAI2BB2X1 U344 ( .B0(n365), .B1(n6), .A0N(memory[90]), .A1N(n6), .Y(n138) );
  OAI2BB2X1 U345 ( .B0(n364), .B1(n6), .A0N(memory[91]), .A1N(n6), .Y(n139) );
  OAI2BB2X1 U346 ( .B0(n367), .B1(n7), .A0N(memory[104]), .A1N(n7), .Y(n152)
         );
  OAI2BB2X1 U347 ( .B0(n366), .B1(n7), .A0N(memory[105]), .A1N(n7), .Y(n153)
         );
  OAI2BB2X1 U348 ( .B0(n365), .B1(n7), .A0N(memory[106]), .A1N(n7), .Y(n154)
         );
  OAI2BB2X1 U349 ( .B0(n364), .B1(n7), .A0N(memory[107]), .A1N(n7), .Y(n155)
         );
  OAI2BB2X1 U350 ( .B0(n367), .B1(n8), .A0N(memory[120]), .A1N(n8), .Y(n168)
         );
  OAI2BB2X1 U351 ( .B0(n366), .B1(n8), .A0N(memory[121]), .A1N(n8), .Y(n169)
         );
  OAI2BB2X1 U352 ( .B0(n365), .B1(n8), .A0N(memory[122]), .A1N(n8), .Y(n170)
         );
  OAI2BB2X1 U353 ( .B0(n364), .B1(n8), .A0N(memory[123]), .A1N(n8), .Y(n171)
         );
  OAI2BB2X1 U354 ( .B0(n367), .B1(n9), .A0N(memory[136]), .A1N(n9), .Y(n184)
         );
  OAI2BB2X1 U355 ( .B0(n366), .B1(n9), .A0N(memory[137]), .A1N(n9), .Y(n185)
         );
  OAI2BB2X1 U356 ( .B0(n365), .B1(n9), .A0N(memory[138]), .A1N(n9), .Y(n186)
         );
  OAI2BB2X1 U357 ( .B0(n364), .B1(n9), .A0N(memory[139]), .A1N(n9), .Y(n187)
         );
  OAI2BB2X1 U358 ( .B0(n367), .B1(n10), .A0N(memory[152]), .A1N(n10), .Y(n200)
         );
  OAI2BB2X1 U359 ( .B0(n366), .B1(n10), .A0N(memory[153]), .A1N(n10), .Y(n201)
         );
  OAI2BB2X1 U360 ( .B0(n365), .B1(n10), .A0N(memory[154]), .A1N(n10), .Y(n202)
         );
  OAI2BB2X1 U361 ( .B0(n364), .B1(n10), .A0N(memory[155]), .A1N(n10), .Y(n203)
         );
  OAI2BB2X1 U362 ( .B0(n367), .B1(n11), .A0N(memory[168]), .A1N(n11), .Y(n216)
         );
  OAI2BB2X1 U363 ( .B0(n366), .B1(n11), .A0N(memory[169]), .A1N(n11), .Y(n217)
         );
  OAI2BB2X1 U364 ( .B0(n365), .B1(n11), .A0N(memory[170]), .A1N(n11), .Y(n218)
         );
  OAI2BB2X1 U365 ( .B0(n364), .B1(n11), .A0N(memory[171]), .A1N(n11), .Y(n219)
         );
  OAI2BB2X1 U366 ( .B0(n367), .B1(n12), .A0N(memory[184]), .A1N(n12), .Y(n232)
         );
  OAI2BB2X1 U367 ( .B0(n366), .B1(n12), .A0N(memory[185]), .A1N(n12), .Y(n233)
         );
  OAI2BB2X1 U368 ( .B0(n365), .B1(n12), .A0N(memory[186]), .A1N(n12), .Y(n234)
         );
  OAI2BB2X1 U369 ( .B0(n364), .B1(n12), .A0N(memory[187]), .A1N(n12), .Y(n235)
         );
  OAI2BB2X1 U370 ( .B0(n367), .B1(n13), .A0N(memory[200]), .A1N(n13), .Y(n248)
         );
  OAI2BB2X1 U371 ( .B0(n366), .B1(n13), .A0N(memory[201]), .A1N(n13), .Y(n249)
         );
  OAI2BB2X1 U372 ( .B0(n365), .B1(n13), .A0N(memory[202]), .A1N(n13), .Y(n250)
         );
  OAI2BB2X1 U373 ( .B0(n364), .B1(n13), .A0N(memory[203]), .A1N(n13), .Y(n251)
         );
  OAI2BB2X1 U374 ( .B0(n367), .B1(n14), .A0N(memory[216]), .A1N(n14), .Y(n264)
         );
  OAI2BB2X1 U375 ( .B0(n366), .B1(n14), .A0N(memory[217]), .A1N(n14), .Y(n265)
         );
  OAI2BB2X1 U376 ( .B0(n365), .B1(n14), .A0N(memory[218]), .A1N(n14), .Y(n266)
         );
  OAI2BB2X1 U377 ( .B0(n364), .B1(n14), .A0N(memory[219]), .A1N(n14), .Y(n267)
         );
  OAI2BB2X1 U378 ( .B0(n367), .B1(n15), .A0N(memory[232]), .A1N(n15), .Y(n280)
         );
  OAI2BB2X1 U379 ( .B0(n366), .B1(n15), .A0N(memory[233]), .A1N(n15), .Y(n281)
         );
  OAI2BB2X1 U380 ( .B0(n365), .B1(n15), .A0N(memory[234]), .A1N(n15), .Y(n282)
         );
  OAI2BB2X1 U381 ( .B0(n364), .B1(n15), .A0N(memory[235]), .A1N(n15), .Y(n283)
         );
  OAI2BB2X1 U382 ( .B0(n367), .B1(n16), .A0N(memory[248]), .A1N(n16), .Y(n296)
         );
  OAI2BB2X1 U383 ( .B0(n366), .B1(n16), .A0N(memory[249]), .A1N(n16), .Y(n297)
         );
  OAI2BB2X1 U384 ( .B0(n365), .B1(n16), .A0N(memory[250]), .A1N(n16), .Y(n298)
         );
  OAI2BB2X1 U385 ( .B0(n364), .B1(n16), .A0N(memory[251]), .A1N(n16), .Y(n299)
         );
  BUFX3 U386 ( .A(n47), .Y(n357) );
  NAND2BX1 U387 ( .AN(wr_rd), .B(en), .Y(n47) );
  NOR2BX1 U388 ( .AN(n35), .B(addr[3]), .Y(n45) );
  BUFX3 U389 ( .A(addr[2]), .Y(n355) );
  INVX1 U390 ( .A(addr[2]), .Y(n359) );
  AND2X2 U391 ( .A(wr_rd), .B(en), .Y(n35) );
  AND2X2 U392 ( .A(addr[3]), .B(n35), .Y(n33) );
  INVX1 U393 ( .A(din[0]), .Y(n375) );
  INVX1 U394 ( .A(din[1]), .Y(n374) );
  INVX1 U395 ( .A(din[2]), .Y(n373) );
  INVX1 U396 ( .A(din[3]), .Y(n372) );
  INVX1 U397 ( .A(din[4]), .Y(n371) );
  INVX1 U398 ( .A(din[5]), .Y(n370) );
  INVX1 U399 ( .A(din[6]), .Y(n369) );
  INVX1 U400 ( .A(din[7]), .Y(n368) );
  INVX1 U401 ( .A(din[8]), .Y(n367) );
  INVX1 U402 ( .A(din[9]), .Y(n366) );
  INVX1 U403 ( .A(din[10]), .Y(n365) );
  INVX1 U404 ( .A(din[11]), .Y(n364) );
  INVX1 U405 ( .A(din[12]), .Y(n363) );
  INVX1 U406 ( .A(din[13]), .Y(n362) );
  INVX1 U407 ( .A(din[14]), .Y(n361) );
  INVX1 U408 ( .A(din[15]), .Y(n360) );
endmodule


module mem4x4_3 ( clk, rstn, en, wr_rd, addr, din, dout );
  input [3:0] addr;
  input [15:0] din;
  output [15:0] dout;
  input clk, rstn, en, wr_rd;
  wire   N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48,
         N49, N50, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n23, n25, n27, n28, n30, n31, n34, n36,
         n38, n40, n41, n42, n43, n44, n46, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643;
  wire   [255:0] memory;

  DFFRHQX1 memory_reg_1__15_ ( .D(n392), .CK(clk), .RN(rstn), .Q(memory[239])
         );
  DFFRHQX1 memory_reg_1__14_ ( .D(n393), .CK(clk), .RN(rstn), .Q(memory[238])
         );
  DFFRHQX1 memory_reg_1__13_ ( .D(n394), .CK(clk), .RN(rstn), .Q(memory[237])
         );
  DFFRHQX1 memory_reg_1__12_ ( .D(n395), .CK(clk), .RN(rstn), .Q(memory[236])
         );
  DFFRHQX1 memory_reg_1__11_ ( .D(n396), .CK(clk), .RN(rstn), .Q(memory[235])
         );
  DFFRHQX1 memory_reg_1__10_ ( .D(n397), .CK(clk), .RN(rstn), .Q(memory[234])
         );
  DFFRHQX1 memory_reg_1__9_ ( .D(n398), .CK(clk), .RN(rstn), .Q(memory[233])
         );
  DFFRHQX1 memory_reg_1__8_ ( .D(n399), .CK(clk), .RN(rstn), .Q(memory[232])
         );
  DFFRHQX1 memory_reg_1__7_ ( .D(n400), .CK(clk), .RN(rstn), .Q(memory[231])
         );
  DFFRHQX1 memory_reg_1__6_ ( .D(n401), .CK(clk), .RN(rstn), .Q(memory[230])
         );
  DFFRHQX1 memory_reg_1__5_ ( .D(n402), .CK(clk), .RN(rstn), .Q(memory[229])
         );
  DFFRHQX1 memory_reg_1__4_ ( .D(n403), .CK(clk), .RN(rstn), .Q(memory[228])
         );
  DFFRHQX1 memory_reg_1__3_ ( .D(n404), .CK(clk), .RN(rstn), .Q(memory[227])
         );
  DFFRHQX1 memory_reg_1__2_ ( .D(n405), .CK(clk), .RN(rstn), .Q(memory[226])
         );
  DFFRHQX1 memory_reg_1__1_ ( .D(n406), .CK(clk), .RN(rstn), .Q(memory[225])
         );
  DFFRHQX1 memory_reg_1__0_ ( .D(n407), .CK(clk), .RN(rstn), .Q(memory[224])
         );
  DFFRHQX1 memory_reg_5__15_ ( .D(n456), .CK(clk), .RN(rstn), .Q(memory[175])
         );
  DFFRHQX1 memory_reg_5__14_ ( .D(n457), .CK(clk), .RN(rstn), .Q(memory[174])
         );
  DFFRHQX1 memory_reg_5__13_ ( .D(n458), .CK(clk), .RN(rstn), .Q(memory[173])
         );
  DFFRHQX1 memory_reg_5__12_ ( .D(n459), .CK(clk), .RN(rstn), .Q(memory[172])
         );
  DFFRHQX1 memory_reg_5__11_ ( .D(n460), .CK(clk), .RN(rstn), .Q(memory[171])
         );
  DFFRHQX1 memory_reg_5__10_ ( .D(n461), .CK(clk), .RN(rstn), .Q(memory[170])
         );
  DFFRHQX1 memory_reg_5__9_ ( .D(n462), .CK(clk), .RN(rstn), .Q(memory[169])
         );
  DFFRHQX1 memory_reg_5__8_ ( .D(n463), .CK(clk), .RN(rstn), .Q(memory[168])
         );
  DFFRHQX1 memory_reg_5__7_ ( .D(n464), .CK(clk), .RN(rstn), .Q(memory[167])
         );
  DFFRHQX1 memory_reg_5__6_ ( .D(n465), .CK(clk), .RN(rstn), .Q(memory[166])
         );
  DFFRHQX1 memory_reg_5__5_ ( .D(n466), .CK(clk), .RN(rstn), .Q(memory[165])
         );
  DFFRHQX1 memory_reg_5__4_ ( .D(n467), .CK(clk), .RN(rstn), .Q(memory[164])
         );
  DFFRHQX1 memory_reg_5__3_ ( .D(n468), .CK(clk), .RN(rstn), .Q(memory[163])
         );
  DFFRHQX1 memory_reg_5__2_ ( .D(n469), .CK(clk), .RN(rstn), .Q(memory[162])
         );
  DFFRHQX1 memory_reg_5__1_ ( .D(n470), .CK(clk), .RN(rstn), .Q(memory[161])
         );
  DFFRHQX1 memory_reg_5__0_ ( .D(n471), .CK(clk), .RN(rstn), .Q(memory[160])
         );
  DFFRHQX1 memory_reg_9__15_ ( .D(n520), .CK(clk), .RN(rstn), .Q(memory[111])
         );
  DFFRHQX1 memory_reg_9__14_ ( .D(n521), .CK(clk), .RN(rstn), .Q(memory[110])
         );
  DFFRHQX1 memory_reg_9__13_ ( .D(n522), .CK(clk), .RN(rstn), .Q(memory[109])
         );
  DFFRHQX1 memory_reg_9__12_ ( .D(n523), .CK(clk), .RN(rstn), .Q(memory[108])
         );
  DFFRHQX1 memory_reg_9__11_ ( .D(n524), .CK(clk), .RN(rstn), .Q(memory[107])
         );
  DFFRHQX1 memory_reg_9__10_ ( .D(n525), .CK(clk), .RN(rstn), .Q(memory[106])
         );
  DFFRHQX1 memory_reg_9__9_ ( .D(n526), .CK(clk), .RN(rstn), .Q(memory[105])
         );
  DFFRHQX1 memory_reg_9__8_ ( .D(n527), .CK(clk), .RN(rstn), .Q(memory[104])
         );
  DFFRHQX1 memory_reg_9__7_ ( .D(n528), .CK(clk), .RN(rstn), .Q(memory[103])
         );
  DFFRHQX1 memory_reg_9__6_ ( .D(n529), .CK(clk), .RN(rstn), .Q(memory[102])
         );
  DFFRHQX1 memory_reg_9__5_ ( .D(n530), .CK(clk), .RN(rstn), .Q(memory[101])
         );
  DFFRHQX1 memory_reg_9__4_ ( .D(n531), .CK(clk), .RN(rstn), .Q(memory[100])
         );
  DFFRHQX1 memory_reg_9__3_ ( .D(n532), .CK(clk), .RN(rstn), .Q(memory[99]) );
  DFFRHQX1 memory_reg_9__2_ ( .D(n533), .CK(clk), .RN(rstn), .Q(memory[98]) );
  DFFRHQX1 memory_reg_9__1_ ( .D(n534), .CK(clk), .RN(rstn), .Q(memory[97]) );
  DFFRHQX1 memory_reg_9__0_ ( .D(n535), .CK(clk), .RN(rstn), .Q(memory[96]) );
  DFFRHQX1 memory_reg_13__15_ ( .D(n584), .CK(clk), .RN(rstn), .Q(memory[47])
         );
  DFFRHQX1 memory_reg_13__14_ ( .D(n585), .CK(clk), .RN(rstn), .Q(memory[46])
         );
  DFFRHQX1 memory_reg_13__13_ ( .D(n586), .CK(clk), .RN(rstn), .Q(memory[45])
         );
  DFFRHQX1 memory_reg_13__12_ ( .D(n587), .CK(clk), .RN(rstn), .Q(memory[44])
         );
  DFFRHQX1 memory_reg_13__11_ ( .D(n588), .CK(clk), .RN(rstn), .Q(memory[43])
         );
  DFFRHQX1 memory_reg_13__10_ ( .D(n589), .CK(clk), .RN(rstn), .Q(memory[42])
         );
  DFFRHQX1 memory_reg_13__9_ ( .D(n590), .CK(clk), .RN(rstn), .Q(memory[41])
         );
  DFFRHQX1 memory_reg_13__8_ ( .D(n591), .CK(clk), .RN(rstn), .Q(memory[40])
         );
  DFFRHQX1 memory_reg_13__7_ ( .D(n592), .CK(clk), .RN(rstn), .Q(memory[39])
         );
  DFFRHQX1 memory_reg_13__6_ ( .D(n593), .CK(clk), .RN(rstn), .Q(memory[38])
         );
  DFFRHQX1 memory_reg_13__5_ ( .D(n594), .CK(clk), .RN(rstn), .Q(memory[37])
         );
  DFFRHQX1 memory_reg_13__4_ ( .D(n595), .CK(clk), .RN(rstn), .Q(memory[36])
         );
  DFFRHQX1 memory_reg_13__3_ ( .D(n596), .CK(clk), .RN(rstn), .Q(memory[35])
         );
  DFFRHQX1 memory_reg_13__2_ ( .D(n597), .CK(clk), .RN(rstn), .Q(memory[34])
         );
  DFFRHQX1 memory_reg_13__1_ ( .D(n598), .CK(clk), .RN(rstn), .Q(memory[33])
         );
  DFFRHQX1 memory_reg_13__0_ ( .D(n599), .CK(clk), .RN(rstn), .Q(memory[32])
         );
  DFFRHQX1 memory_reg_3__15_ ( .D(n424), .CK(clk), .RN(rstn), .Q(memory[207])
         );
  DFFRHQX1 memory_reg_3__14_ ( .D(n425), .CK(clk), .RN(rstn), .Q(memory[206])
         );
  DFFRHQX1 memory_reg_3__13_ ( .D(n426), .CK(clk), .RN(rstn), .Q(memory[205])
         );
  DFFRHQX1 memory_reg_3__12_ ( .D(n427), .CK(clk), .RN(rstn), .Q(memory[204])
         );
  DFFRHQX1 memory_reg_3__11_ ( .D(n428), .CK(clk), .RN(rstn), .Q(memory[203])
         );
  DFFRHQX1 memory_reg_3__10_ ( .D(n429), .CK(clk), .RN(rstn), .Q(memory[202])
         );
  DFFRHQX1 memory_reg_3__9_ ( .D(n430), .CK(clk), .RN(rstn), .Q(memory[201])
         );
  DFFRHQX1 memory_reg_3__8_ ( .D(n431), .CK(clk), .RN(rstn), .Q(memory[200])
         );
  DFFRHQX1 memory_reg_3__7_ ( .D(n432), .CK(clk), .RN(rstn), .Q(memory[199])
         );
  DFFRHQX1 memory_reg_3__6_ ( .D(n433), .CK(clk), .RN(rstn), .Q(memory[198])
         );
  DFFRHQX1 memory_reg_3__5_ ( .D(n434), .CK(clk), .RN(rstn), .Q(memory[197])
         );
  DFFRHQX1 memory_reg_3__4_ ( .D(n435), .CK(clk), .RN(rstn), .Q(memory[196])
         );
  DFFRHQX1 memory_reg_3__3_ ( .D(n436), .CK(clk), .RN(rstn), .Q(memory[195])
         );
  DFFRHQX1 memory_reg_3__2_ ( .D(n437), .CK(clk), .RN(rstn), .Q(memory[194])
         );
  DFFRHQX1 memory_reg_3__1_ ( .D(n438), .CK(clk), .RN(rstn), .Q(memory[193])
         );
  DFFRHQX1 memory_reg_3__0_ ( .D(n439), .CK(clk), .RN(rstn), .Q(memory[192])
         );
  DFFRHQX1 memory_reg_7__15_ ( .D(n488), .CK(clk), .RN(rstn), .Q(memory[143])
         );
  DFFRHQX1 memory_reg_7__14_ ( .D(n489), .CK(clk), .RN(rstn), .Q(memory[142])
         );
  DFFRHQX1 memory_reg_7__13_ ( .D(n490), .CK(clk), .RN(rstn), .Q(memory[141])
         );
  DFFRHQX1 memory_reg_7__12_ ( .D(n491), .CK(clk), .RN(rstn), .Q(memory[140])
         );
  DFFRHQX1 memory_reg_7__11_ ( .D(n492), .CK(clk), .RN(rstn), .Q(memory[139])
         );
  DFFRHQX1 memory_reg_7__10_ ( .D(n493), .CK(clk), .RN(rstn), .Q(memory[138])
         );
  DFFRHQX1 memory_reg_7__9_ ( .D(n494), .CK(clk), .RN(rstn), .Q(memory[137])
         );
  DFFRHQX1 memory_reg_7__8_ ( .D(n495), .CK(clk), .RN(rstn), .Q(memory[136])
         );
  DFFRHQX1 memory_reg_7__7_ ( .D(n496), .CK(clk), .RN(rstn), .Q(memory[135])
         );
  DFFRHQX1 memory_reg_7__6_ ( .D(n497), .CK(clk), .RN(rstn), .Q(memory[134])
         );
  DFFRHQX1 memory_reg_7__5_ ( .D(n498), .CK(clk), .RN(rstn), .Q(memory[133])
         );
  DFFRHQX1 memory_reg_7__4_ ( .D(n499), .CK(clk), .RN(rstn), .Q(memory[132])
         );
  DFFRHQX1 memory_reg_7__3_ ( .D(n500), .CK(clk), .RN(rstn), .Q(memory[131])
         );
  DFFRHQX1 memory_reg_7__2_ ( .D(n501), .CK(clk), .RN(rstn), .Q(memory[130])
         );
  DFFRHQX1 memory_reg_7__1_ ( .D(n502), .CK(clk), .RN(rstn), .Q(memory[129])
         );
  DFFRHQX1 memory_reg_7__0_ ( .D(n503), .CK(clk), .RN(rstn), .Q(memory[128])
         );
  DFFRHQX1 memory_reg_11__15_ ( .D(n552), .CK(clk), .RN(rstn), .Q(memory[79])
         );
  DFFRHQX1 memory_reg_11__14_ ( .D(n553), .CK(clk), .RN(rstn), .Q(memory[78])
         );
  DFFRHQX1 memory_reg_11__13_ ( .D(n554), .CK(clk), .RN(rstn), .Q(memory[77])
         );
  DFFRHQX1 memory_reg_11__12_ ( .D(n555), .CK(clk), .RN(rstn), .Q(memory[76])
         );
  DFFRHQX1 memory_reg_11__11_ ( .D(n556), .CK(clk), .RN(rstn), .Q(memory[75])
         );
  DFFRHQX1 memory_reg_11__10_ ( .D(n557), .CK(clk), .RN(rstn), .Q(memory[74])
         );
  DFFRHQX1 memory_reg_11__9_ ( .D(n558), .CK(clk), .RN(rstn), .Q(memory[73])
         );
  DFFRHQX1 memory_reg_11__8_ ( .D(n559), .CK(clk), .RN(rstn), .Q(memory[72])
         );
  DFFRHQX1 memory_reg_11__7_ ( .D(n560), .CK(clk), .RN(rstn), .Q(memory[71])
         );
  DFFRHQX1 memory_reg_11__6_ ( .D(n561), .CK(clk), .RN(rstn), .Q(memory[70])
         );
  DFFRHQX1 memory_reg_11__5_ ( .D(n562), .CK(clk), .RN(rstn), .Q(memory[69])
         );
  DFFRHQX1 memory_reg_11__4_ ( .D(n563), .CK(clk), .RN(rstn), .Q(memory[68])
         );
  DFFRHQX1 memory_reg_11__3_ ( .D(n564), .CK(clk), .RN(rstn), .Q(memory[67])
         );
  DFFRHQX1 memory_reg_11__2_ ( .D(n565), .CK(clk), .RN(rstn), .Q(memory[66])
         );
  DFFRHQX1 memory_reg_11__1_ ( .D(n566), .CK(clk), .RN(rstn), .Q(memory[65])
         );
  DFFRHQX1 memory_reg_11__0_ ( .D(n567), .CK(clk), .RN(rstn), .Q(memory[64])
         );
  DFFRHQX1 memory_reg_15__15_ ( .D(n616), .CK(clk), .RN(rstn), .Q(memory[15])
         );
  DFFRHQX1 memory_reg_15__14_ ( .D(n617), .CK(clk), .RN(rstn), .Q(memory[14])
         );
  DFFRHQX1 memory_reg_15__13_ ( .D(n618), .CK(clk), .RN(rstn), .Q(memory[13])
         );
  DFFRHQX1 memory_reg_15__12_ ( .D(n619), .CK(clk), .RN(rstn), .Q(memory[12])
         );
  DFFRHQX1 memory_reg_15__11_ ( .D(n620), .CK(clk), .RN(rstn), .Q(memory[11])
         );
  DFFRHQX1 memory_reg_15__10_ ( .D(n621), .CK(clk), .RN(rstn), .Q(memory[10])
         );
  DFFRHQX1 memory_reg_15__9_ ( .D(n622), .CK(clk), .RN(rstn), .Q(memory[9]) );
  DFFRHQX1 memory_reg_15__8_ ( .D(n623), .CK(clk), .RN(rstn), .Q(memory[8]) );
  DFFRHQX1 memory_reg_15__7_ ( .D(n624), .CK(clk), .RN(rstn), .Q(memory[7]) );
  DFFRHQX1 memory_reg_15__6_ ( .D(n625), .CK(clk), .RN(rstn), .Q(memory[6]) );
  DFFRHQX1 memory_reg_15__5_ ( .D(n626), .CK(clk), .RN(rstn), .Q(memory[5]) );
  DFFRHQX1 memory_reg_15__4_ ( .D(n627), .CK(clk), .RN(rstn), .Q(memory[4]) );
  DFFRHQX1 memory_reg_15__3_ ( .D(n628), .CK(clk), .RN(rstn), .Q(memory[3]) );
  DFFRHQX1 memory_reg_15__2_ ( .D(n629), .CK(clk), .RN(rstn), .Q(memory[2]) );
  DFFRHQX1 memory_reg_15__1_ ( .D(n630), .CK(clk), .RN(rstn), .Q(memory[1]) );
  DFFRHQX1 memory_reg_15__0_ ( .D(n631), .CK(clk), .RN(rstn), .Q(memory[0]) );
  DFFRHQX1 memory_reg_0__15_ ( .D(n376), .CK(clk), .RN(rstn), .Q(memory[255])
         );
  DFFRHQX1 memory_reg_0__14_ ( .D(n377), .CK(clk), .RN(rstn), .Q(memory[254])
         );
  DFFRHQX1 memory_reg_0__13_ ( .D(n378), .CK(clk), .RN(rstn), .Q(memory[253])
         );
  DFFRHQX1 memory_reg_0__12_ ( .D(n379), .CK(clk), .RN(rstn), .Q(memory[252])
         );
  DFFRHQX1 memory_reg_0__11_ ( .D(n380), .CK(clk), .RN(rstn), .Q(memory[251])
         );
  DFFRHQX1 memory_reg_0__10_ ( .D(n381), .CK(clk), .RN(rstn), .Q(memory[250])
         );
  DFFRHQX1 memory_reg_0__9_ ( .D(n382), .CK(clk), .RN(rstn), .Q(memory[249])
         );
  DFFRHQX1 memory_reg_0__8_ ( .D(n383), .CK(clk), .RN(rstn), .Q(memory[248])
         );
  DFFRHQX1 memory_reg_0__7_ ( .D(n384), .CK(clk), .RN(rstn), .Q(memory[247])
         );
  DFFRHQX1 memory_reg_0__6_ ( .D(n385), .CK(clk), .RN(rstn), .Q(memory[246])
         );
  DFFRHQX1 memory_reg_0__5_ ( .D(n386), .CK(clk), .RN(rstn), .Q(memory[245])
         );
  DFFRHQX1 memory_reg_0__4_ ( .D(n387), .CK(clk), .RN(rstn), .Q(memory[244])
         );
  DFFRHQX1 memory_reg_0__3_ ( .D(n388), .CK(clk), .RN(rstn), .Q(memory[243])
         );
  DFFRHQX1 memory_reg_0__2_ ( .D(n389), .CK(clk), .RN(rstn), .Q(memory[242])
         );
  DFFRHQX1 memory_reg_0__1_ ( .D(n390), .CK(clk), .RN(rstn), .Q(memory[241])
         );
  DFFRHQX1 memory_reg_0__0_ ( .D(n391), .CK(clk), .RN(rstn), .Q(memory[240])
         );
  DFFRHQX1 memory_reg_4__15_ ( .D(n440), .CK(clk), .RN(rstn), .Q(memory[191])
         );
  DFFRHQX1 memory_reg_4__14_ ( .D(n441), .CK(clk), .RN(rstn), .Q(memory[190])
         );
  DFFRHQX1 memory_reg_4__13_ ( .D(n442), .CK(clk), .RN(rstn), .Q(memory[189])
         );
  DFFRHQX1 memory_reg_4__12_ ( .D(n443), .CK(clk), .RN(rstn), .Q(memory[188])
         );
  DFFRHQX1 memory_reg_4__11_ ( .D(n444), .CK(clk), .RN(rstn), .Q(memory[187])
         );
  DFFRHQX1 memory_reg_4__10_ ( .D(n445), .CK(clk), .RN(rstn), .Q(memory[186])
         );
  DFFRHQX1 memory_reg_4__9_ ( .D(n446), .CK(clk), .RN(rstn), .Q(memory[185])
         );
  DFFRHQX1 memory_reg_4__8_ ( .D(n447), .CK(clk), .RN(rstn), .Q(memory[184])
         );
  DFFRHQX1 memory_reg_4__7_ ( .D(n448), .CK(clk), .RN(rstn), .Q(memory[183])
         );
  DFFRHQX1 memory_reg_4__6_ ( .D(n449), .CK(clk), .RN(rstn), .Q(memory[182])
         );
  DFFRHQX1 memory_reg_4__5_ ( .D(n450), .CK(clk), .RN(rstn), .Q(memory[181])
         );
  DFFRHQX1 memory_reg_4__4_ ( .D(n451), .CK(clk), .RN(rstn), .Q(memory[180])
         );
  DFFRHQX1 memory_reg_4__3_ ( .D(n452), .CK(clk), .RN(rstn), .Q(memory[179])
         );
  DFFRHQX1 memory_reg_4__2_ ( .D(n453), .CK(clk), .RN(rstn), .Q(memory[178])
         );
  DFFRHQX1 memory_reg_4__1_ ( .D(n454), .CK(clk), .RN(rstn), .Q(memory[177])
         );
  DFFRHQX1 memory_reg_4__0_ ( .D(n455), .CK(clk), .RN(rstn), .Q(memory[176])
         );
  DFFRHQX1 memory_reg_8__15_ ( .D(n504), .CK(clk), .RN(rstn), .Q(memory[127])
         );
  DFFRHQX1 memory_reg_8__14_ ( .D(n505), .CK(clk), .RN(rstn), .Q(memory[126])
         );
  DFFRHQX1 memory_reg_8__13_ ( .D(n506), .CK(clk), .RN(rstn), .Q(memory[125])
         );
  DFFRHQX1 memory_reg_8__12_ ( .D(n507), .CK(clk), .RN(rstn), .Q(memory[124])
         );
  DFFRHQX1 memory_reg_8__11_ ( .D(n508), .CK(clk), .RN(rstn), .Q(memory[123])
         );
  DFFRHQX1 memory_reg_8__10_ ( .D(n509), .CK(clk), .RN(rstn), .Q(memory[122])
         );
  DFFRHQX1 memory_reg_8__9_ ( .D(n510), .CK(clk), .RN(rstn), .Q(memory[121])
         );
  DFFRHQX1 memory_reg_8__8_ ( .D(n511), .CK(clk), .RN(rstn), .Q(memory[120])
         );
  DFFRHQX1 memory_reg_8__7_ ( .D(n512), .CK(clk), .RN(rstn), .Q(memory[119])
         );
  DFFRHQX1 memory_reg_8__6_ ( .D(n513), .CK(clk), .RN(rstn), .Q(memory[118])
         );
  DFFRHQX1 memory_reg_8__5_ ( .D(n514), .CK(clk), .RN(rstn), .Q(memory[117])
         );
  DFFRHQX1 memory_reg_8__4_ ( .D(n515), .CK(clk), .RN(rstn), .Q(memory[116])
         );
  DFFRHQX1 memory_reg_8__3_ ( .D(n516), .CK(clk), .RN(rstn), .Q(memory[115])
         );
  DFFRHQX1 memory_reg_8__2_ ( .D(n517), .CK(clk), .RN(rstn), .Q(memory[114])
         );
  DFFRHQX1 memory_reg_8__1_ ( .D(n518), .CK(clk), .RN(rstn), .Q(memory[113])
         );
  DFFRHQX1 memory_reg_8__0_ ( .D(n519), .CK(clk), .RN(rstn), .Q(memory[112])
         );
  DFFRHQX1 memory_reg_12__15_ ( .D(n568), .CK(clk), .RN(rstn), .Q(memory[63])
         );
  DFFRHQX1 memory_reg_12__14_ ( .D(n569), .CK(clk), .RN(rstn), .Q(memory[62])
         );
  DFFRHQX1 memory_reg_12__13_ ( .D(n570), .CK(clk), .RN(rstn), .Q(memory[61])
         );
  DFFRHQX1 memory_reg_12__12_ ( .D(n571), .CK(clk), .RN(rstn), .Q(memory[60])
         );
  DFFRHQX1 memory_reg_12__11_ ( .D(n572), .CK(clk), .RN(rstn), .Q(memory[59])
         );
  DFFRHQX1 memory_reg_12__10_ ( .D(n573), .CK(clk), .RN(rstn), .Q(memory[58])
         );
  DFFRHQX1 memory_reg_12__9_ ( .D(n574), .CK(clk), .RN(rstn), .Q(memory[57])
         );
  DFFRHQX1 memory_reg_12__8_ ( .D(n575), .CK(clk), .RN(rstn), .Q(memory[56])
         );
  DFFRHQX1 memory_reg_12__7_ ( .D(n576), .CK(clk), .RN(rstn), .Q(memory[55])
         );
  DFFRHQX1 memory_reg_12__6_ ( .D(n577), .CK(clk), .RN(rstn), .Q(memory[54])
         );
  DFFRHQX1 memory_reg_12__5_ ( .D(n578), .CK(clk), .RN(rstn), .Q(memory[53])
         );
  DFFRHQX1 memory_reg_12__4_ ( .D(n579), .CK(clk), .RN(rstn), .Q(memory[52])
         );
  DFFRHQX1 memory_reg_12__3_ ( .D(n580), .CK(clk), .RN(rstn), .Q(memory[51])
         );
  DFFRHQX1 memory_reg_12__2_ ( .D(n581), .CK(clk), .RN(rstn), .Q(memory[50])
         );
  DFFRHQX1 memory_reg_12__1_ ( .D(n582), .CK(clk), .RN(rstn), .Q(memory[49])
         );
  DFFRHQX1 memory_reg_12__0_ ( .D(n583), .CK(clk), .RN(rstn), .Q(memory[48])
         );
  DFFRHQX1 memory_reg_2__15_ ( .D(n408), .CK(clk), .RN(rstn), .Q(memory[223])
         );
  DFFRHQX1 memory_reg_2__14_ ( .D(n409), .CK(clk), .RN(rstn), .Q(memory[222])
         );
  DFFRHQX1 memory_reg_2__13_ ( .D(n410), .CK(clk), .RN(rstn), .Q(memory[221])
         );
  DFFRHQX1 memory_reg_2__12_ ( .D(n411), .CK(clk), .RN(rstn), .Q(memory[220])
         );
  DFFRHQX1 memory_reg_2__11_ ( .D(n412), .CK(clk), .RN(rstn), .Q(memory[219])
         );
  DFFRHQX1 memory_reg_2__10_ ( .D(n413), .CK(clk), .RN(rstn), .Q(memory[218])
         );
  DFFRHQX1 memory_reg_2__9_ ( .D(n414), .CK(clk), .RN(rstn), .Q(memory[217])
         );
  DFFRHQX1 memory_reg_2__8_ ( .D(n415), .CK(clk), .RN(rstn), .Q(memory[216])
         );
  DFFRHQX1 memory_reg_2__7_ ( .D(n416), .CK(clk), .RN(rstn), .Q(memory[215])
         );
  DFFRHQX1 memory_reg_2__6_ ( .D(n417), .CK(clk), .RN(rstn), .Q(memory[214])
         );
  DFFRHQX1 memory_reg_2__5_ ( .D(n418), .CK(clk), .RN(rstn), .Q(memory[213])
         );
  DFFRHQX1 memory_reg_2__4_ ( .D(n419), .CK(clk), .RN(rstn), .Q(memory[212])
         );
  DFFRHQX1 memory_reg_2__3_ ( .D(n420), .CK(clk), .RN(rstn), .Q(memory[211])
         );
  DFFRHQX1 memory_reg_2__2_ ( .D(n421), .CK(clk), .RN(rstn), .Q(memory[210])
         );
  DFFRHQX1 memory_reg_2__1_ ( .D(n422), .CK(clk), .RN(rstn), .Q(memory[209])
         );
  DFFRHQX1 memory_reg_2__0_ ( .D(n423), .CK(clk), .RN(rstn), .Q(memory[208])
         );
  DFFRHQX1 memory_reg_6__15_ ( .D(n472), .CK(clk), .RN(rstn), .Q(memory[159])
         );
  DFFRHQX1 memory_reg_6__14_ ( .D(n473), .CK(clk), .RN(rstn), .Q(memory[158])
         );
  DFFRHQX1 memory_reg_6__13_ ( .D(n474), .CK(clk), .RN(rstn), .Q(memory[157])
         );
  DFFRHQX1 memory_reg_6__12_ ( .D(n475), .CK(clk), .RN(rstn), .Q(memory[156])
         );
  DFFRHQX1 memory_reg_6__11_ ( .D(n476), .CK(clk), .RN(rstn), .Q(memory[155])
         );
  DFFRHQX1 memory_reg_6__10_ ( .D(n477), .CK(clk), .RN(rstn), .Q(memory[154])
         );
  DFFRHQX1 memory_reg_6__9_ ( .D(n478), .CK(clk), .RN(rstn), .Q(memory[153])
         );
  DFFRHQX1 memory_reg_6__8_ ( .D(n479), .CK(clk), .RN(rstn), .Q(memory[152])
         );
  DFFRHQX1 memory_reg_6__7_ ( .D(n480), .CK(clk), .RN(rstn), .Q(memory[151])
         );
  DFFRHQX1 memory_reg_6__6_ ( .D(n481), .CK(clk), .RN(rstn), .Q(memory[150])
         );
  DFFRHQX1 memory_reg_6__5_ ( .D(n482), .CK(clk), .RN(rstn), .Q(memory[149])
         );
  DFFRHQX1 memory_reg_6__4_ ( .D(n483), .CK(clk), .RN(rstn), .Q(memory[148])
         );
  DFFRHQX1 memory_reg_6__3_ ( .D(n484), .CK(clk), .RN(rstn), .Q(memory[147])
         );
  DFFRHQX1 memory_reg_6__2_ ( .D(n485), .CK(clk), .RN(rstn), .Q(memory[146])
         );
  DFFRHQX1 memory_reg_6__1_ ( .D(n486), .CK(clk), .RN(rstn), .Q(memory[145])
         );
  DFFRHQX1 memory_reg_6__0_ ( .D(n487), .CK(clk), .RN(rstn), .Q(memory[144])
         );
  DFFRHQX1 memory_reg_10__15_ ( .D(n536), .CK(clk), .RN(rstn), .Q(memory[95])
         );
  DFFRHQX1 memory_reg_10__14_ ( .D(n537), .CK(clk), .RN(rstn), .Q(memory[94])
         );
  DFFRHQX1 memory_reg_10__13_ ( .D(n538), .CK(clk), .RN(rstn), .Q(memory[93])
         );
  DFFRHQX1 memory_reg_10__12_ ( .D(n539), .CK(clk), .RN(rstn), .Q(memory[92])
         );
  DFFRHQX1 memory_reg_10__11_ ( .D(n540), .CK(clk), .RN(rstn), .Q(memory[91])
         );
  DFFRHQX1 memory_reg_10__10_ ( .D(n541), .CK(clk), .RN(rstn), .Q(memory[90])
         );
  DFFRHQX1 memory_reg_10__9_ ( .D(n542), .CK(clk), .RN(rstn), .Q(memory[89])
         );
  DFFRHQX1 memory_reg_10__8_ ( .D(n543), .CK(clk), .RN(rstn), .Q(memory[88])
         );
  DFFRHQX1 memory_reg_10__7_ ( .D(n544), .CK(clk), .RN(rstn), .Q(memory[87])
         );
  DFFRHQX1 memory_reg_10__6_ ( .D(n545), .CK(clk), .RN(rstn), .Q(memory[86])
         );
  DFFRHQX1 memory_reg_10__5_ ( .D(n546), .CK(clk), .RN(rstn), .Q(memory[85])
         );
  DFFRHQX1 memory_reg_10__4_ ( .D(n547), .CK(clk), .RN(rstn), .Q(memory[84])
         );
  DFFRHQX1 memory_reg_10__3_ ( .D(n548), .CK(clk), .RN(rstn), .Q(memory[83])
         );
  DFFRHQX1 memory_reg_10__2_ ( .D(n549), .CK(clk), .RN(rstn), .Q(memory[82])
         );
  DFFRHQX1 memory_reg_10__1_ ( .D(n550), .CK(clk), .RN(rstn), .Q(memory[81])
         );
  DFFRHQX1 memory_reg_10__0_ ( .D(n551), .CK(clk), .RN(rstn), .Q(memory[80])
         );
  DFFRHQX1 memory_reg_14__15_ ( .D(n600), .CK(clk), .RN(rstn), .Q(memory[31])
         );
  DFFRHQX1 memory_reg_14__14_ ( .D(n601), .CK(clk), .RN(rstn), .Q(memory[30])
         );
  DFFRHQX1 memory_reg_14__13_ ( .D(n602), .CK(clk), .RN(rstn), .Q(memory[29])
         );
  DFFRHQX1 memory_reg_14__12_ ( .D(n603), .CK(clk), .RN(rstn), .Q(memory[28])
         );
  DFFRHQX1 memory_reg_14__11_ ( .D(n604), .CK(clk), .RN(rstn), .Q(memory[27])
         );
  DFFRHQX1 memory_reg_14__10_ ( .D(n605), .CK(clk), .RN(rstn), .Q(memory[26])
         );
  DFFRHQX1 memory_reg_14__9_ ( .D(n606), .CK(clk), .RN(rstn), .Q(memory[25])
         );
  DFFRHQX1 memory_reg_14__8_ ( .D(n607), .CK(clk), .RN(rstn), .Q(memory[24])
         );
  DFFRHQX1 memory_reg_14__7_ ( .D(n608), .CK(clk), .RN(rstn), .Q(memory[23])
         );
  DFFRHQX1 memory_reg_14__6_ ( .D(n609), .CK(clk), .RN(rstn), .Q(memory[22])
         );
  DFFRHQX1 memory_reg_14__5_ ( .D(n610), .CK(clk), .RN(rstn), .Q(memory[21])
         );
  DFFRHQX1 memory_reg_14__4_ ( .D(n611), .CK(clk), .RN(rstn), .Q(memory[20])
         );
  DFFRHQX1 memory_reg_14__3_ ( .D(n612), .CK(clk), .RN(rstn), .Q(memory[19])
         );
  DFFRHQX1 memory_reg_14__2_ ( .D(n613), .CK(clk), .RN(rstn), .Q(memory[18])
         );
  DFFRHQX1 memory_reg_14__1_ ( .D(n614), .CK(clk), .RN(rstn), .Q(memory[17])
         );
  DFFRHQX1 memory_reg_14__0_ ( .D(n615), .CK(clk), .RN(rstn), .Q(memory[16])
         );
  NAND2X1 U2 ( .A(n643), .B(n642), .Y(n1) );
  NAND2X1 U3 ( .A(n641), .B(n643), .Y(n2) );
  NAND2X1 U4 ( .A(n640), .B(n642), .Y(n3) );
  NAND2X1 U5 ( .A(n640), .B(n641), .Y(n4) );
  NAND2X1 U6 ( .A(n639), .B(n642), .Y(n5) );
  NAND2X1 U7 ( .A(n639), .B(n641), .Y(n6) );
  NAND2X1 U8 ( .A(n638), .B(n642), .Y(n7) );
  NAND2X1 U9 ( .A(n638), .B(n641), .Y(n8) );
  NAND2X1 U10 ( .A(n635), .B(n643), .Y(n9) );
  NAND2X1 U11 ( .A(n634), .B(n643), .Y(n10) );
  NAND2X1 U12 ( .A(n635), .B(n640), .Y(n11) );
  NAND2X1 U13 ( .A(n634), .B(n640), .Y(n12) );
  NAND2X1 U14 ( .A(n635), .B(n639), .Y(n13) );
  NAND2X1 U15 ( .A(n634), .B(n639), .Y(n14) );
  NAND2X1 U16 ( .A(n635), .B(n638), .Y(n15) );
  NAND2X1 U17 ( .A(n634), .B(n638), .Y(n16) );
  INVX1 U18 ( .A(n351), .Y(n352) );
  INVX1 U19 ( .A(n351), .Y(n353) );
  INVX1 U20 ( .A(n351), .Y(n354) );
  INVX1 U21 ( .A(n358), .Y(n349) );
  INVX1 U22 ( .A(n358), .Y(n350) );
  INVX1 U23 ( .A(addr[0]), .Y(n351) );
  NOR2X1 U24 ( .A(n359), .B(addr[1]), .Y(n640) );
  NOR2X1 U25 ( .A(n359), .B(n358), .Y(n643) );
  AND2X2 U26 ( .A(n633), .B(addr[0]), .Y(n635) );
  AND2X2 U27 ( .A(n633), .B(n351), .Y(n634) );
  AND2X2 U28 ( .A(n637), .B(n351), .Y(n641) );
  AND2X2 U29 ( .A(n637), .B(n353), .Y(n642) );
  MX4X1 U30 ( .A(memory[176]), .B(memory[160]), .C(memory[144]), .D(
        memory[128]), .S0(n353), .S1(n349), .Y(n19) );
  MX4X1 U31 ( .A(memory[177]), .B(memory[161]), .C(memory[145]), .D(
        memory[129]), .S0(n352), .S1(n349), .Y(n27) );
  MX4X1 U32 ( .A(memory[178]), .B(memory[162]), .C(memory[146]), .D(
        memory[130]), .S0(n352), .S1(n349), .Y(n34) );
  MX4X1 U33 ( .A(memory[179]), .B(memory[163]), .C(memory[147]), .D(
        memory[131]), .S0(n352), .S1(n349), .Y(n41) );
  MX4X1 U34 ( .A(memory[180]), .B(memory[164]), .C(memory[148]), .D(
        memory[132]), .S0(n353), .S1(n350), .Y(n46) );
  MX4X1 U35 ( .A(memory[181]), .B(memory[165]), .C(memory[149]), .D(
        memory[133]), .S0(n353), .S1(n350), .Y(n307) );
  MX4X1 U36 ( .A(memory[182]), .B(memory[166]), .C(memory[150]), .D(
        memory[134]), .S0(n353), .S1(n350), .Y(n311) );
  MX4X1 U37 ( .A(memory[183]), .B(memory[167]), .C(memory[151]), .D(
        memory[135]), .S0(n352), .S1(n350), .Y(n315) );
  MX4X1 U38 ( .A(memory[184]), .B(memory[168]), .C(memory[152]), .D(
        memory[136]), .S0(n354), .S1(n349), .Y(n319) );
  MX4X1 U39 ( .A(memory[185]), .B(memory[169]), .C(memory[153]), .D(
        memory[137]), .S0(n353), .S1(n350), .Y(n323) );
  MX4X1 U40 ( .A(memory[186]), .B(memory[170]), .C(memory[154]), .D(
        memory[138]), .S0(n354), .S1(n350), .Y(n327) );
  MX4X1 U41 ( .A(memory[187]), .B(memory[171]), .C(memory[155]), .D(
        memory[139]), .S0(n354), .S1(addr[1]), .Y(n331) );
  MX4X1 U42 ( .A(memory[188]), .B(memory[172]), .C(memory[156]), .D(
        memory[140]), .S0(n354), .S1(addr[1]), .Y(n335) );
  MX4X1 U43 ( .A(memory[189]), .B(memory[173]), .C(memory[157]), .D(
        memory[141]), .S0(n354), .S1(addr[1]), .Y(n339) );
  MX4X1 U44 ( .A(memory[190]), .B(memory[174]), .C(memory[158]), .D(
        memory[142]), .S0(n353), .S1(addr[1]), .Y(n343) );
  MX4X1 U45 ( .A(memory[191]), .B(memory[175]), .C(memory[159]), .D(
        memory[143]), .S0(addr[0]), .S1(addr[1]), .Y(n347) );
  MX4X1 U46 ( .A(memory[48]), .B(memory[32]), .C(memory[16]), .D(memory[0]), 
        .S0(n352), .S1(n350), .Y(n17) );
  MX4X1 U47 ( .A(memory[49]), .B(memory[33]), .C(memory[17]), .D(memory[1]), 
        .S0(n352), .S1(n349), .Y(n23) );
  MX4X1 U48 ( .A(memory[50]), .B(memory[34]), .C(memory[18]), .D(memory[2]), 
        .S0(n352), .S1(n349), .Y(n30) );
  MX4X1 U49 ( .A(memory[51]), .B(memory[35]), .C(memory[19]), .D(memory[3]), 
        .S0(n352), .S1(n349), .Y(n38) );
  MX4X1 U50 ( .A(memory[52]), .B(memory[36]), .C(memory[20]), .D(memory[4]), 
        .S0(n353), .S1(n350), .Y(n43) );
  MX4X1 U51 ( .A(memory[53]), .B(memory[37]), .C(memory[21]), .D(memory[5]), 
        .S0(n353), .S1(n350), .Y(n305) );
  MX4X1 U52 ( .A(memory[54]), .B(memory[38]), .C(memory[22]), .D(memory[6]), 
        .S0(n353), .S1(n350), .Y(n309) );
  MX4X1 U53 ( .A(memory[55]), .B(memory[39]), .C(memory[23]), .D(memory[7]), 
        .S0(n354), .S1(n349), .Y(n313) );
  MX4X1 U54 ( .A(memory[56]), .B(memory[40]), .C(memory[24]), .D(memory[8]), 
        .S0(n353), .S1(n350), .Y(n317) );
  MX4X1 U55 ( .A(memory[57]), .B(memory[41]), .C(memory[25]), .D(memory[9]), 
        .S0(addr[0]), .S1(n349), .Y(n321) );
  MX4X1 U56 ( .A(memory[58]), .B(memory[42]), .C(memory[26]), .D(memory[10]), 
        .S0(n354), .S1(n350), .Y(n325) );
  MX4X1 U57 ( .A(memory[59]), .B(memory[43]), .C(memory[27]), .D(memory[11]), 
        .S0(n354), .S1(n349), .Y(n329) );
  MX4X1 U58 ( .A(memory[60]), .B(memory[44]), .C(memory[28]), .D(memory[12]), 
        .S0(n354), .S1(n349), .Y(n333) );
  MX4X1 U59 ( .A(memory[61]), .B(memory[45]), .C(memory[29]), .D(memory[13]), 
        .S0(n352), .S1(n349), .Y(n337) );
  MX4X1 U60 ( .A(memory[62]), .B(memory[46]), .C(memory[30]), .D(memory[14]), 
        .S0(n352), .S1(n350), .Y(n341) );
  MX4X1 U61 ( .A(memory[63]), .B(memory[47]), .C(memory[31]), .D(memory[15]), 
        .S0(addr[0]), .S1(addr[1]), .Y(n345) );
  NOR2BX1 U62 ( .AN(N50), .B(n357), .Y(dout[0]) );
  MX4X1 U63 ( .A(n20), .B(n18), .C(n19), .D(n17), .S0(n356), .S1(n355), .Y(N50) );
  MX4X1 U64 ( .A(memory[240]), .B(memory[224]), .C(memory[208]), .D(
        memory[192]), .S0(n354), .S1(addr[1]), .Y(n20) );
  MX4X1 U65 ( .A(memory[112]), .B(memory[96]), .C(memory[80]), .D(memory[64]), 
        .S0(n352), .S1(n349), .Y(n18) );
  NOR2BX1 U66 ( .AN(N49), .B(n357), .Y(dout[1]) );
  MX4X1 U67 ( .A(n28), .B(n25), .C(n27), .D(n23), .S0(n356), .S1(n355), .Y(N49) );
  MX4X1 U68 ( .A(memory[241]), .B(memory[225]), .C(memory[209]), .D(
        memory[193]), .S0(n352), .S1(n349), .Y(n28) );
  MX4X1 U69 ( .A(memory[113]), .B(memory[97]), .C(memory[81]), .D(memory[65]), 
        .S0(n352), .S1(n349), .Y(n25) );
  NOR2BX1 U70 ( .AN(N48), .B(n357), .Y(dout[2]) );
  MX4X1 U71 ( .A(n36), .B(n31), .C(n34), .D(n30), .S0(n356), .S1(n355), .Y(N48) );
  MX4X1 U72 ( .A(memory[242]), .B(memory[226]), .C(memory[210]), .D(
        memory[194]), .S0(n352), .S1(n349), .Y(n36) );
  MX4X1 U73 ( .A(memory[114]), .B(memory[98]), .C(memory[82]), .D(memory[66]), 
        .S0(n352), .S1(n349), .Y(n31) );
  NOR2BX1 U74 ( .AN(N47), .B(n357), .Y(dout[3]) );
  MX4X1 U75 ( .A(n42), .B(n40), .C(n41), .D(n38), .S0(n356), .S1(n355), .Y(N47) );
  MX4X1 U76 ( .A(memory[243]), .B(memory[227]), .C(memory[211]), .D(
        memory[195]), .S0(n352), .S1(n349), .Y(n42) );
  MX4X1 U77 ( .A(memory[115]), .B(memory[99]), .C(memory[83]), .D(memory[67]), 
        .S0(n352), .S1(n349), .Y(n40) );
  NOR2BX1 U78 ( .AN(N46), .B(n357), .Y(dout[4]) );
  MX4X1 U79 ( .A(n304), .B(n44), .C(n46), .D(n43), .S0(n356), .S1(n355), .Y(
        N46) );
  MX4X1 U80 ( .A(memory[244]), .B(memory[228]), .C(memory[212]), .D(
        memory[196]), .S0(n353), .S1(n350), .Y(n304) );
  MX4X1 U81 ( .A(memory[116]), .B(memory[100]), .C(memory[84]), .D(memory[68]), 
        .S0(n353), .S1(n350), .Y(n44) );
  NOR2BX1 U82 ( .AN(N45), .B(n357), .Y(dout[5]) );
  MX4X1 U83 ( .A(n308), .B(n306), .C(n307), .D(n305), .S0(n356), .S1(n355), 
        .Y(N45) );
  MX4X1 U84 ( .A(memory[245]), .B(memory[229]), .C(memory[213]), .D(
        memory[197]), .S0(n353), .S1(n350), .Y(n308) );
  MX4X1 U85 ( .A(memory[117]), .B(memory[101]), .C(memory[85]), .D(memory[69]), 
        .S0(n353), .S1(n350), .Y(n306) );
  NOR2BX1 U86 ( .AN(N44), .B(n357), .Y(dout[6]) );
  MX4X1 U87 ( .A(n312), .B(n310), .C(n311), .D(n309), .S0(n356), .S1(n355), 
        .Y(N44) );
  MX4X1 U88 ( .A(memory[246]), .B(memory[230]), .C(memory[214]), .D(
        memory[198]), .S0(n353), .S1(n350), .Y(n312) );
  MX4X1 U89 ( .A(memory[118]), .B(memory[102]), .C(memory[86]), .D(memory[70]), 
        .S0(n353), .S1(n350), .Y(n310) );
  NOR2BX1 U90 ( .AN(N43), .B(n357), .Y(dout[7]) );
  MX4X1 U91 ( .A(n316), .B(n314), .C(n315), .D(n313), .S0(n356), .S1(n355), 
        .Y(N43) );
  MX4X1 U92 ( .A(memory[247]), .B(memory[231]), .C(memory[215]), .D(
        memory[199]), .S0(n354), .S1(n349), .Y(n316) );
  MX4X1 U93 ( .A(memory[119]), .B(memory[103]), .C(memory[87]), .D(memory[71]), 
        .S0(n354), .S1(n350), .Y(n314) );
  NOR2BX1 U94 ( .AN(N42), .B(n357), .Y(dout[8]) );
  MX4X1 U95 ( .A(n320), .B(n318), .C(n319), .D(n317), .S0(n356), .S1(n355), 
        .Y(N42) );
  MX4X1 U96 ( .A(memory[248]), .B(memory[232]), .C(memory[216]), .D(
        memory[200]), .S0(addr[0]), .S1(n350), .Y(n320) );
  MX4X1 U97 ( .A(memory[120]), .B(memory[104]), .C(memory[88]), .D(memory[72]), 
        .S0(n353), .S1(n350), .Y(n318) );
  NOR2BX1 U98 ( .AN(N41), .B(n357), .Y(dout[9]) );
  MX4X1 U99 ( .A(n324), .B(n322), .C(n323), .D(n321), .S0(n356), .S1(n355), 
        .Y(N41) );
  MX4X1 U100 ( .A(memory[249]), .B(memory[233]), .C(memory[217]), .D(
        memory[201]), .S0(addr[0]), .S1(n349), .Y(n324) );
  MX4X1 U101 ( .A(memory[121]), .B(memory[105]), .C(memory[89]), .D(memory[73]), .S0(n352), .S1(n349), .Y(n322) );
  NOR2BX1 U102 ( .AN(N40), .B(n357), .Y(dout[10]) );
  MX4X1 U103 ( .A(n328), .B(n326), .C(n327), .D(n325), .S0(n356), .S1(n355), 
        .Y(N40) );
  MX4X1 U104 ( .A(memory[250]), .B(memory[234]), .C(memory[218]), .D(
        memory[202]), .S0(n354), .S1(addr[1]), .Y(n328) );
  MX4X1 U105 ( .A(memory[122]), .B(memory[106]), .C(memory[90]), .D(memory[74]), .S0(n354), .S1(addr[1]), .Y(n326) );
  NOR2BX1 U106 ( .AN(N39), .B(n357), .Y(dout[11]) );
  MX4X1 U107 ( .A(n332), .B(n330), .C(n331), .D(n329), .S0(n356), .S1(n355), 
        .Y(N39) );
  MX4X1 U108 ( .A(memory[251]), .B(memory[235]), .C(memory[219]), .D(
        memory[203]), .S0(n354), .S1(addr[1]), .Y(n332) );
  MX4X1 U109 ( .A(memory[123]), .B(memory[107]), .C(memory[91]), .D(memory[75]), .S0(n354), .S1(addr[1]), .Y(n330) );
  NOR2BX1 U110 ( .AN(N38), .B(n357), .Y(dout[12]) );
  MX4X1 U111 ( .A(n336), .B(n334), .C(n335), .D(n333), .S0(n356), .S1(n355), 
        .Y(N38) );
  MX4X1 U112 ( .A(memory[252]), .B(memory[236]), .C(memory[220]), .D(
        memory[204]), .S0(n354), .S1(addr[1]), .Y(n336) );
  MX4X1 U113 ( .A(memory[124]), .B(memory[108]), .C(memory[92]), .D(memory[76]), .S0(n354), .S1(addr[1]), .Y(n334) );
  NOR2BX1 U114 ( .AN(N37), .B(n357), .Y(dout[13]) );
  MX4X1 U115 ( .A(n340), .B(n338), .C(n339), .D(n337), .S0(n356), .S1(n355), 
        .Y(N37) );
  MX4X1 U116 ( .A(memory[253]), .B(memory[237]), .C(memory[221]), .D(
        memory[205]), .S0(addr[0]), .S1(addr[1]), .Y(n340) );
  MX4X1 U117 ( .A(memory[125]), .B(memory[109]), .C(memory[93]), .D(memory[77]), .S0(addr[0]), .S1(addr[1]), .Y(n338) );
  NOR2BX1 U118 ( .AN(N36), .B(n357), .Y(dout[14]) );
  MX4X1 U119 ( .A(n344), .B(n342), .C(n343), .D(n341), .S0(n356), .S1(n355), 
        .Y(N36) );
  MX4X1 U120 ( .A(memory[254]), .B(memory[238]), .C(memory[222]), .D(
        memory[206]), .S0(addr[0]), .S1(addr[1]), .Y(n344) );
  MX4X1 U121 ( .A(memory[126]), .B(memory[110]), .C(memory[94]), .D(memory[78]), .S0(addr[0]), .S1(addr[1]), .Y(n342) );
  NOR2BX1 U122 ( .AN(N35), .B(n357), .Y(dout[15]) );
  MX4X1 U123 ( .A(n348), .B(n346), .C(n347), .D(n345), .S0(n356), .S1(n355), 
        .Y(N35) );
  MX4X1 U124 ( .A(memory[255]), .B(memory[239]), .C(memory[223]), .D(
        memory[207]), .S0(addr[0]), .S1(addr[1]), .Y(n348) );
  MX4X1 U125 ( .A(memory[127]), .B(memory[111]), .C(memory[95]), .D(memory[79]), .S0(addr[0]), .S1(addr[1]), .Y(n346) );
  INVX1 U126 ( .A(addr[1]), .Y(n358) );
  NOR2X1 U127 ( .A(n358), .B(addr[2]), .Y(n639) );
  NOR2X1 U128 ( .A(addr[1]), .B(addr[2]), .Y(n638) );
  BUFX3 U129 ( .A(addr[3]), .Y(n356) );
  OAI2BB2X1 U130 ( .B0(n1), .B1(n375), .A0N(memory[0]), .A1N(n1), .Y(n631) );
  OAI2BB2X1 U131 ( .B0(n1), .B1(n374), .A0N(memory[1]), .A1N(n1), .Y(n630) );
  OAI2BB2X1 U132 ( .B0(n1), .B1(n373), .A0N(memory[2]), .A1N(n1), .Y(n629) );
  OAI2BB2X1 U133 ( .B0(n1), .B1(n372), .A0N(memory[3]), .A1N(n1), .Y(n628) );
  OAI2BB2X1 U134 ( .B0(n1), .B1(n371), .A0N(memory[4]), .A1N(n1), .Y(n627) );
  OAI2BB2X1 U135 ( .B0(n1), .B1(n370), .A0N(memory[5]), .A1N(n1), .Y(n626) );
  OAI2BB2X1 U136 ( .B0(n1), .B1(n369), .A0N(memory[6]), .A1N(n1), .Y(n625) );
  OAI2BB2X1 U137 ( .B0(n1), .B1(n368), .A0N(memory[7]), .A1N(n1), .Y(n624) );
  OAI2BB2X1 U138 ( .B0(n1), .B1(n367), .A0N(memory[8]), .A1N(n1), .Y(n623) );
  OAI2BB2X1 U139 ( .B0(n1), .B1(n366), .A0N(memory[9]), .A1N(n1), .Y(n622) );
  OAI2BB2X1 U140 ( .B0(n1), .B1(n365), .A0N(memory[10]), .A1N(n1), .Y(n621) );
  OAI2BB2X1 U141 ( .B0(n1), .B1(n364), .A0N(memory[11]), .A1N(n1), .Y(n620) );
  OAI2BB2X1 U142 ( .B0(n1), .B1(n363), .A0N(memory[12]), .A1N(n1), .Y(n619) );
  OAI2BB2X1 U143 ( .B0(n1), .B1(n362), .A0N(memory[13]), .A1N(n1), .Y(n618) );
  OAI2BB2X1 U144 ( .B0(n1), .B1(n361), .A0N(memory[14]), .A1N(n1), .Y(n617) );
  OAI2BB2X1 U145 ( .B0(n1), .B1(n360), .A0N(memory[15]), .A1N(n1), .Y(n616) );
  OAI2BB2X1 U146 ( .B0(n375), .B1(n2), .A0N(memory[16]), .A1N(n2), .Y(n615) );
  OAI2BB2X1 U147 ( .B0(n374), .B1(n2), .A0N(memory[17]), .A1N(n2), .Y(n614) );
  OAI2BB2X1 U148 ( .B0(n373), .B1(n2), .A0N(memory[18]), .A1N(n2), .Y(n613) );
  OAI2BB2X1 U149 ( .B0(n372), .B1(n2), .A0N(memory[19]), .A1N(n2), .Y(n612) );
  OAI2BB2X1 U150 ( .B0(n371), .B1(n2), .A0N(memory[20]), .A1N(n2), .Y(n611) );
  OAI2BB2X1 U151 ( .B0(n370), .B1(n2), .A0N(memory[21]), .A1N(n2), .Y(n610) );
  OAI2BB2X1 U152 ( .B0(n369), .B1(n2), .A0N(memory[22]), .A1N(n2), .Y(n609) );
  OAI2BB2X1 U153 ( .B0(n368), .B1(n2), .A0N(memory[23]), .A1N(n2), .Y(n608) );
  OAI2BB2X1 U154 ( .B0(n363), .B1(n2), .A0N(memory[28]), .A1N(n2), .Y(n603) );
  OAI2BB2X1 U155 ( .B0(n362), .B1(n2), .A0N(memory[29]), .A1N(n2), .Y(n602) );
  OAI2BB2X1 U156 ( .B0(n361), .B1(n2), .A0N(memory[30]), .A1N(n2), .Y(n601) );
  OAI2BB2X1 U157 ( .B0(n360), .B1(n2), .A0N(memory[31]), .A1N(n2), .Y(n600) );
  OAI2BB2X1 U158 ( .B0(n375), .B1(n3), .A0N(memory[32]), .A1N(n3), .Y(n599) );
  OAI2BB2X1 U159 ( .B0(n374), .B1(n3), .A0N(memory[33]), .A1N(n3), .Y(n598) );
  OAI2BB2X1 U160 ( .B0(n373), .B1(n3), .A0N(memory[34]), .A1N(n3), .Y(n597) );
  OAI2BB2X1 U161 ( .B0(n372), .B1(n3), .A0N(memory[35]), .A1N(n3), .Y(n596) );
  OAI2BB2X1 U162 ( .B0(n371), .B1(n3), .A0N(memory[36]), .A1N(n3), .Y(n595) );
  OAI2BB2X1 U163 ( .B0(n370), .B1(n3), .A0N(memory[37]), .A1N(n3), .Y(n594) );
  OAI2BB2X1 U164 ( .B0(n369), .B1(n3), .A0N(memory[38]), .A1N(n3), .Y(n593) );
  OAI2BB2X1 U165 ( .B0(n368), .B1(n3), .A0N(memory[39]), .A1N(n3), .Y(n592) );
  OAI2BB2X1 U166 ( .B0(n363), .B1(n3), .A0N(memory[44]), .A1N(n3), .Y(n587) );
  OAI2BB2X1 U167 ( .B0(n362), .B1(n3), .A0N(memory[45]), .A1N(n3), .Y(n586) );
  OAI2BB2X1 U168 ( .B0(n361), .B1(n3), .A0N(memory[46]), .A1N(n3), .Y(n585) );
  OAI2BB2X1 U169 ( .B0(n360), .B1(n3), .A0N(memory[47]), .A1N(n3), .Y(n584) );
  OAI2BB2X1 U170 ( .B0(n375), .B1(n4), .A0N(memory[48]), .A1N(n4), .Y(n583) );
  OAI2BB2X1 U171 ( .B0(n374), .B1(n4), .A0N(memory[49]), .A1N(n4), .Y(n582) );
  OAI2BB2X1 U172 ( .B0(n373), .B1(n4), .A0N(memory[50]), .A1N(n4), .Y(n581) );
  OAI2BB2X1 U173 ( .B0(n372), .B1(n4), .A0N(memory[51]), .A1N(n4), .Y(n580) );
  OAI2BB2X1 U174 ( .B0(n371), .B1(n4), .A0N(memory[52]), .A1N(n4), .Y(n579) );
  OAI2BB2X1 U175 ( .B0(n370), .B1(n4), .A0N(memory[53]), .A1N(n4), .Y(n578) );
  OAI2BB2X1 U176 ( .B0(n369), .B1(n4), .A0N(memory[54]), .A1N(n4), .Y(n577) );
  OAI2BB2X1 U177 ( .B0(n368), .B1(n4), .A0N(memory[55]), .A1N(n4), .Y(n576) );
  OAI2BB2X1 U178 ( .B0(n363), .B1(n4), .A0N(memory[60]), .A1N(n4), .Y(n571) );
  OAI2BB2X1 U179 ( .B0(n362), .B1(n4), .A0N(memory[61]), .A1N(n4), .Y(n570) );
  OAI2BB2X1 U180 ( .B0(n361), .B1(n4), .A0N(memory[62]), .A1N(n4), .Y(n569) );
  OAI2BB2X1 U181 ( .B0(n360), .B1(n4), .A0N(memory[63]), .A1N(n4), .Y(n568) );
  OAI2BB2X1 U182 ( .B0(n375), .B1(n5), .A0N(memory[64]), .A1N(n5), .Y(n567) );
  OAI2BB2X1 U183 ( .B0(n374), .B1(n5), .A0N(memory[65]), .A1N(n5), .Y(n566) );
  OAI2BB2X1 U184 ( .B0(n373), .B1(n5), .A0N(memory[66]), .A1N(n5), .Y(n565) );
  OAI2BB2X1 U185 ( .B0(n372), .B1(n5), .A0N(memory[67]), .A1N(n5), .Y(n564) );
  OAI2BB2X1 U186 ( .B0(n371), .B1(n5), .A0N(memory[68]), .A1N(n5), .Y(n563) );
  OAI2BB2X1 U187 ( .B0(n370), .B1(n5), .A0N(memory[69]), .A1N(n5), .Y(n562) );
  OAI2BB2X1 U188 ( .B0(n369), .B1(n5), .A0N(memory[70]), .A1N(n5), .Y(n561) );
  OAI2BB2X1 U189 ( .B0(n368), .B1(n5), .A0N(memory[71]), .A1N(n5), .Y(n560) );
  OAI2BB2X1 U190 ( .B0(n363), .B1(n5), .A0N(memory[76]), .A1N(n5), .Y(n555) );
  OAI2BB2X1 U191 ( .B0(n362), .B1(n5), .A0N(memory[77]), .A1N(n5), .Y(n554) );
  OAI2BB2X1 U192 ( .B0(n361), .B1(n5), .A0N(memory[78]), .A1N(n5), .Y(n553) );
  OAI2BB2X1 U193 ( .B0(n360), .B1(n5), .A0N(memory[79]), .A1N(n5), .Y(n552) );
  OAI2BB2X1 U194 ( .B0(n375), .B1(n6), .A0N(memory[80]), .A1N(n6), .Y(n551) );
  OAI2BB2X1 U195 ( .B0(n374), .B1(n6), .A0N(memory[81]), .A1N(n6), .Y(n550) );
  OAI2BB2X1 U196 ( .B0(n373), .B1(n6), .A0N(memory[82]), .A1N(n6), .Y(n549) );
  OAI2BB2X1 U197 ( .B0(n372), .B1(n6), .A0N(memory[83]), .A1N(n6), .Y(n548) );
  OAI2BB2X1 U198 ( .B0(n371), .B1(n6), .A0N(memory[84]), .A1N(n6), .Y(n547) );
  OAI2BB2X1 U199 ( .B0(n370), .B1(n6), .A0N(memory[85]), .A1N(n6), .Y(n546) );
  OAI2BB2X1 U200 ( .B0(n369), .B1(n6), .A0N(memory[86]), .A1N(n6), .Y(n545) );
  OAI2BB2X1 U201 ( .B0(n368), .B1(n6), .A0N(memory[87]), .A1N(n6), .Y(n544) );
  OAI2BB2X1 U202 ( .B0(n363), .B1(n6), .A0N(memory[92]), .A1N(n6), .Y(n539) );
  OAI2BB2X1 U203 ( .B0(n362), .B1(n6), .A0N(memory[93]), .A1N(n6), .Y(n538) );
  OAI2BB2X1 U204 ( .B0(n361), .B1(n6), .A0N(memory[94]), .A1N(n6), .Y(n537) );
  OAI2BB2X1 U205 ( .B0(n360), .B1(n6), .A0N(memory[95]), .A1N(n6), .Y(n536) );
  OAI2BB2X1 U206 ( .B0(n375), .B1(n7), .A0N(memory[96]), .A1N(n7), .Y(n535) );
  OAI2BB2X1 U207 ( .B0(n374), .B1(n7), .A0N(memory[97]), .A1N(n7), .Y(n534) );
  OAI2BB2X1 U208 ( .B0(n373), .B1(n7), .A0N(memory[98]), .A1N(n7), .Y(n533) );
  OAI2BB2X1 U209 ( .B0(n372), .B1(n7), .A0N(memory[99]), .A1N(n7), .Y(n532) );
  OAI2BB2X1 U210 ( .B0(n371), .B1(n7), .A0N(memory[100]), .A1N(n7), .Y(n531)
         );
  OAI2BB2X1 U211 ( .B0(n370), .B1(n7), .A0N(memory[101]), .A1N(n7), .Y(n530)
         );
  OAI2BB2X1 U212 ( .B0(n369), .B1(n7), .A0N(memory[102]), .A1N(n7), .Y(n529)
         );
  OAI2BB2X1 U213 ( .B0(n368), .B1(n7), .A0N(memory[103]), .A1N(n7), .Y(n528)
         );
  OAI2BB2X1 U214 ( .B0(n363), .B1(n7), .A0N(memory[108]), .A1N(n7), .Y(n523)
         );
  OAI2BB2X1 U215 ( .B0(n362), .B1(n7), .A0N(memory[109]), .A1N(n7), .Y(n522)
         );
  OAI2BB2X1 U216 ( .B0(n361), .B1(n7), .A0N(memory[110]), .A1N(n7), .Y(n521)
         );
  OAI2BB2X1 U217 ( .B0(n360), .B1(n7), .A0N(memory[111]), .A1N(n7), .Y(n520)
         );
  OAI2BB2X1 U218 ( .B0(n375), .B1(n8), .A0N(memory[112]), .A1N(n8), .Y(n519)
         );
  OAI2BB2X1 U219 ( .B0(n374), .B1(n8), .A0N(memory[113]), .A1N(n8), .Y(n518)
         );
  OAI2BB2X1 U220 ( .B0(n373), .B1(n8), .A0N(memory[114]), .A1N(n8), .Y(n517)
         );
  OAI2BB2X1 U221 ( .B0(n372), .B1(n8), .A0N(memory[115]), .A1N(n8), .Y(n516)
         );
  OAI2BB2X1 U222 ( .B0(n371), .B1(n8), .A0N(memory[116]), .A1N(n8), .Y(n515)
         );
  OAI2BB2X1 U223 ( .B0(n370), .B1(n8), .A0N(memory[117]), .A1N(n8), .Y(n514)
         );
  OAI2BB2X1 U224 ( .B0(n369), .B1(n8), .A0N(memory[118]), .A1N(n8), .Y(n513)
         );
  OAI2BB2X1 U225 ( .B0(n368), .B1(n8), .A0N(memory[119]), .A1N(n8), .Y(n512)
         );
  OAI2BB2X1 U226 ( .B0(n363), .B1(n8), .A0N(memory[124]), .A1N(n8), .Y(n507)
         );
  OAI2BB2X1 U227 ( .B0(n362), .B1(n8), .A0N(memory[125]), .A1N(n8), .Y(n506)
         );
  OAI2BB2X1 U228 ( .B0(n361), .B1(n8), .A0N(memory[126]), .A1N(n8), .Y(n505)
         );
  OAI2BB2X1 U229 ( .B0(n360), .B1(n8), .A0N(memory[127]), .A1N(n8), .Y(n504)
         );
  OAI2BB2X1 U230 ( .B0(n375), .B1(n9), .A0N(memory[128]), .A1N(n9), .Y(n503)
         );
  OAI2BB2X1 U231 ( .B0(n374), .B1(n9), .A0N(memory[129]), .A1N(n9), .Y(n502)
         );
  OAI2BB2X1 U232 ( .B0(n373), .B1(n9), .A0N(memory[130]), .A1N(n9), .Y(n501)
         );
  OAI2BB2X1 U233 ( .B0(n372), .B1(n9), .A0N(memory[131]), .A1N(n9), .Y(n500)
         );
  OAI2BB2X1 U234 ( .B0(n371), .B1(n9), .A0N(memory[132]), .A1N(n9), .Y(n499)
         );
  OAI2BB2X1 U235 ( .B0(n370), .B1(n9), .A0N(memory[133]), .A1N(n9), .Y(n498)
         );
  OAI2BB2X1 U236 ( .B0(n369), .B1(n9), .A0N(memory[134]), .A1N(n9), .Y(n497)
         );
  OAI2BB2X1 U237 ( .B0(n368), .B1(n9), .A0N(memory[135]), .A1N(n9), .Y(n496)
         );
  OAI2BB2X1 U238 ( .B0(n363), .B1(n9), .A0N(memory[140]), .A1N(n9), .Y(n491)
         );
  OAI2BB2X1 U239 ( .B0(n362), .B1(n9), .A0N(memory[141]), .A1N(n9), .Y(n490)
         );
  OAI2BB2X1 U240 ( .B0(n361), .B1(n9), .A0N(memory[142]), .A1N(n9), .Y(n489)
         );
  OAI2BB2X1 U241 ( .B0(n360), .B1(n9), .A0N(memory[143]), .A1N(n9), .Y(n488)
         );
  OAI2BB2X1 U242 ( .B0(n375), .B1(n10), .A0N(memory[144]), .A1N(n10), .Y(n487)
         );
  OAI2BB2X1 U243 ( .B0(n374), .B1(n10), .A0N(memory[145]), .A1N(n10), .Y(n486)
         );
  OAI2BB2X1 U244 ( .B0(n373), .B1(n10), .A0N(memory[146]), .A1N(n10), .Y(n485)
         );
  OAI2BB2X1 U245 ( .B0(n372), .B1(n10), .A0N(memory[147]), .A1N(n10), .Y(n484)
         );
  OAI2BB2X1 U246 ( .B0(n371), .B1(n10), .A0N(memory[148]), .A1N(n10), .Y(n483)
         );
  OAI2BB2X1 U247 ( .B0(n370), .B1(n10), .A0N(memory[149]), .A1N(n10), .Y(n482)
         );
  OAI2BB2X1 U248 ( .B0(n369), .B1(n10), .A0N(memory[150]), .A1N(n10), .Y(n481)
         );
  OAI2BB2X1 U249 ( .B0(n368), .B1(n10), .A0N(memory[151]), .A1N(n10), .Y(n480)
         );
  OAI2BB2X1 U250 ( .B0(n363), .B1(n10), .A0N(memory[156]), .A1N(n10), .Y(n475)
         );
  OAI2BB2X1 U251 ( .B0(n362), .B1(n10), .A0N(memory[157]), .A1N(n10), .Y(n474)
         );
  OAI2BB2X1 U252 ( .B0(n361), .B1(n10), .A0N(memory[158]), .A1N(n10), .Y(n473)
         );
  OAI2BB2X1 U253 ( .B0(n360), .B1(n10), .A0N(memory[159]), .A1N(n10), .Y(n472)
         );
  OAI2BB2X1 U254 ( .B0(n375), .B1(n11), .A0N(memory[160]), .A1N(n11), .Y(n471)
         );
  OAI2BB2X1 U255 ( .B0(n374), .B1(n11), .A0N(memory[161]), .A1N(n11), .Y(n470)
         );
  OAI2BB2X1 U256 ( .B0(n373), .B1(n11), .A0N(memory[162]), .A1N(n11), .Y(n469)
         );
  OAI2BB2X1 U257 ( .B0(n372), .B1(n11), .A0N(memory[163]), .A1N(n11), .Y(n468)
         );
  OAI2BB2X1 U258 ( .B0(n371), .B1(n11), .A0N(memory[164]), .A1N(n11), .Y(n467)
         );
  OAI2BB2X1 U259 ( .B0(n370), .B1(n11), .A0N(memory[165]), .A1N(n11), .Y(n466)
         );
  OAI2BB2X1 U260 ( .B0(n369), .B1(n11), .A0N(memory[166]), .A1N(n11), .Y(n465)
         );
  OAI2BB2X1 U261 ( .B0(n368), .B1(n11), .A0N(memory[167]), .A1N(n11), .Y(n464)
         );
  OAI2BB2X1 U262 ( .B0(n363), .B1(n11), .A0N(memory[172]), .A1N(n11), .Y(n459)
         );
  OAI2BB2X1 U263 ( .B0(n362), .B1(n11), .A0N(memory[173]), .A1N(n11), .Y(n458)
         );
  OAI2BB2X1 U264 ( .B0(n361), .B1(n11), .A0N(memory[174]), .A1N(n11), .Y(n457)
         );
  OAI2BB2X1 U265 ( .B0(n360), .B1(n11), .A0N(memory[175]), .A1N(n11), .Y(n456)
         );
  OAI2BB2X1 U266 ( .B0(n375), .B1(n12), .A0N(memory[176]), .A1N(n12), .Y(n455)
         );
  OAI2BB2X1 U267 ( .B0(n374), .B1(n12), .A0N(memory[177]), .A1N(n12), .Y(n454)
         );
  OAI2BB2X1 U268 ( .B0(n373), .B1(n12), .A0N(memory[178]), .A1N(n12), .Y(n453)
         );
  OAI2BB2X1 U269 ( .B0(n372), .B1(n12), .A0N(memory[179]), .A1N(n12), .Y(n452)
         );
  OAI2BB2X1 U270 ( .B0(n371), .B1(n12), .A0N(memory[180]), .A1N(n12), .Y(n451)
         );
  OAI2BB2X1 U271 ( .B0(n370), .B1(n12), .A0N(memory[181]), .A1N(n12), .Y(n450)
         );
  OAI2BB2X1 U272 ( .B0(n369), .B1(n12), .A0N(memory[182]), .A1N(n12), .Y(n449)
         );
  OAI2BB2X1 U273 ( .B0(n368), .B1(n12), .A0N(memory[183]), .A1N(n12), .Y(n448)
         );
  OAI2BB2X1 U274 ( .B0(n363), .B1(n12), .A0N(memory[188]), .A1N(n12), .Y(n443)
         );
  OAI2BB2X1 U275 ( .B0(n362), .B1(n12), .A0N(memory[189]), .A1N(n12), .Y(n442)
         );
  OAI2BB2X1 U276 ( .B0(n361), .B1(n12), .A0N(memory[190]), .A1N(n12), .Y(n441)
         );
  OAI2BB2X1 U277 ( .B0(n360), .B1(n12), .A0N(memory[191]), .A1N(n12), .Y(n440)
         );
  OAI2BB2X1 U278 ( .B0(n375), .B1(n13), .A0N(memory[192]), .A1N(n13), .Y(n439)
         );
  OAI2BB2X1 U279 ( .B0(n374), .B1(n13), .A0N(memory[193]), .A1N(n13), .Y(n438)
         );
  OAI2BB2X1 U280 ( .B0(n373), .B1(n13), .A0N(memory[194]), .A1N(n13), .Y(n437)
         );
  OAI2BB2X1 U281 ( .B0(n372), .B1(n13), .A0N(memory[195]), .A1N(n13), .Y(n436)
         );
  OAI2BB2X1 U282 ( .B0(n371), .B1(n13), .A0N(memory[196]), .A1N(n13), .Y(n435)
         );
  OAI2BB2X1 U283 ( .B0(n370), .B1(n13), .A0N(memory[197]), .A1N(n13), .Y(n434)
         );
  OAI2BB2X1 U284 ( .B0(n369), .B1(n13), .A0N(memory[198]), .A1N(n13), .Y(n433)
         );
  OAI2BB2X1 U285 ( .B0(n368), .B1(n13), .A0N(memory[199]), .A1N(n13), .Y(n432)
         );
  OAI2BB2X1 U286 ( .B0(n363), .B1(n13), .A0N(memory[204]), .A1N(n13), .Y(n427)
         );
  OAI2BB2X1 U287 ( .B0(n362), .B1(n13), .A0N(memory[205]), .A1N(n13), .Y(n426)
         );
  OAI2BB2X1 U288 ( .B0(n361), .B1(n13), .A0N(memory[206]), .A1N(n13), .Y(n425)
         );
  OAI2BB2X1 U289 ( .B0(n360), .B1(n13), .A0N(memory[207]), .A1N(n13), .Y(n424)
         );
  OAI2BB2X1 U290 ( .B0(n375), .B1(n14), .A0N(memory[208]), .A1N(n14), .Y(n423)
         );
  OAI2BB2X1 U291 ( .B0(n374), .B1(n14), .A0N(memory[209]), .A1N(n14), .Y(n422)
         );
  OAI2BB2X1 U292 ( .B0(n373), .B1(n14), .A0N(memory[210]), .A1N(n14), .Y(n421)
         );
  OAI2BB2X1 U293 ( .B0(n372), .B1(n14), .A0N(memory[211]), .A1N(n14), .Y(n420)
         );
  OAI2BB2X1 U294 ( .B0(n371), .B1(n14), .A0N(memory[212]), .A1N(n14), .Y(n419)
         );
  OAI2BB2X1 U295 ( .B0(n370), .B1(n14), .A0N(memory[213]), .A1N(n14), .Y(n418)
         );
  OAI2BB2X1 U296 ( .B0(n369), .B1(n14), .A0N(memory[214]), .A1N(n14), .Y(n417)
         );
  OAI2BB2X1 U297 ( .B0(n368), .B1(n14), .A0N(memory[215]), .A1N(n14), .Y(n416)
         );
  OAI2BB2X1 U298 ( .B0(n363), .B1(n14), .A0N(memory[220]), .A1N(n14), .Y(n411)
         );
  OAI2BB2X1 U299 ( .B0(n362), .B1(n14), .A0N(memory[221]), .A1N(n14), .Y(n410)
         );
  OAI2BB2X1 U300 ( .B0(n361), .B1(n14), .A0N(memory[222]), .A1N(n14), .Y(n409)
         );
  OAI2BB2X1 U301 ( .B0(n360), .B1(n14), .A0N(memory[223]), .A1N(n14), .Y(n408)
         );
  OAI2BB2X1 U302 ( .B0(n375), .B1(n15), .A0N(memory[224]), .A1N(n15), .Y(n407)
         );
  OAI2BB2X1 U303 ( .B0(n374), .B1(n15), .A0N(memory[225]), .A1N(n15), .Y(n406)
         );
  OAI2BB2X1 U304 ( .B0(n373), .B1(n15), .A0N(memory[226]), .A1N(n15), .Y(n405)
         );
  OAI2BB2X1 U305 ( .B0(n372), .B1(n15), .A0N(memory[227]), .A1N(n15), .Y(n404)
         );
  OAI2BB2X1 U306 ( .B0(n371), .B1(n15), .A0N(memory[228]), .A1N(n15), .Y(n403)
         );
  OAI2BB2X1 U307 ( .B0(n370), .B1(n15), .A0N(memory[229]), .A1N(n15), .Y(n402)
         );
  OAI2BB2X1 U308 ( .B0(n369), .B1(n15), .A0N(memory[230]), .A1N(n15), .Y(n401)
         );
  OAI2BB2X1 U309 ( .B0(n368), .B1(n15), .A0N(memory[231]), .A1N(n15), .Y(n400)
         );
  OAI2BB2X1 U310 ( .B0(n363), .B1(n15), .A0N(memory[236]), .A1N(n15), .Y(n395)
         );
  OAI2BB2X1 U311 ( .B0(n362), .B1(n15), .A0N(memory[237]), .A1N(n15), .Y(n394)
         );
  OAI2BB2X1 U312 ( .B0(n361), .B1(n15), .A0N(memory[238]), .A1N(n15), .Y(n393)
         );
  OAI2BB2X1 U313 ( .B0(n360), .B1(n15), .A0N(memory[239]), .A1N(n15), .Y(n392)
         );
  OAI2BB2X1 U314 ( .B0(n375), .B1(n16), .A0N(memory[240]), .A1N(n16), .Y(n391)
         );
  OAI2BB2X1 U315 ( .B0(n374), .B1(n16), .A0N(memory[241]), .A1N(n16), .Y(n390)
         );
  OAI2BB2X1 U316 ( .B0(n373), .B1(n16), .A0N(memory[242]), .A1N(n16), .Y(n389)
         );
  OAI2BB2X1 U317 ( .B0(n372), .B1(n16), .A0N(memory[243]), .A1N(n16), .Y(n388)
         );
  OAI2BB2X1 U318 ( .B0(n371), .B1(n16), .A0N(memory[244]), .A1N(n16), .Y(n387)
         );
  OAI2BB2X1 U319 ( .B0(n370), .B1(n16), .A0N(memory[245]), .A1N(n16), .Y(n386)
         );
  OAI2BB2X1 U320 ( .B0(n369), .B1(n16), .A0N(memory[246]), .A1N(n16), .Y(n385)
         );
  OAI2BB2X1 U321 ( .B0(n368), .B1(n16), .A0N(memory[247]), .A1N(n16), .Y(n384)
         );
  OAI2BB2X1 U322 ( .B0(n363), .B1(n16), .A0N(memory[252]), .A1N(n16), .Y(n379)
         );
  OAI2BB2X1 U323 ( .B0(n362), .B1(n16), .A0N(memory[253]), .A1N(n16), .Y(n378)
         );
  OAI2BB2X1 U324 ( .B0(n361), .B1(n16), .A0N(memory[254]), .A1N(n16), .Y(n377)
         );
  OAI2BB2X1 U325 ( .B0(n360), .B1(n16), .A0N(memory[255]), .A1N(n16), .Y(n376)
         );
  OAI2BB2X1 U326 ( .B0(n367), .B1(n2), .A0N(memory[24]), .A1N(n2), .Y(n607) );
  OAI2BB2X1 U327 ( .B0(n366), .B1(n2), .A0N(memory[25]), .A1N(n2), .Y(n606) );
  OAI2BB2X1 U328 ( .B0(n365), .B1(n2), .A0N(memory[26]), .A1N(n2), .Y(n605) );
  OAI2BB2X1 U329 ( .B0(n364), .B1(n2), .A0N(memory[27]), .A1N(n2), .Y(n604) );
  OAI2BB2X1 U330 ( .B0(n367), .B1(n3), .A0N(memory[40]), .A1N(n3), .Y(n591) );
  OAI2BB2X1 U331 ( .B0(n366), .B1(n3), .A0N(memory[41]), .A1N(n3), .Y(n590) );
  OAI2BB2X1 U332 ( .B0(n365), .B1(n3), .A0N(memory[42]), .A1N(n3), .Y(n589) );
  OAI2BB2X1 U333 ( .B0(n364), .B1(n3), .A0N(memory[43]), .A1N(n3), .Y(n588) );
  OAI2BB2X1 U334 ( .B0(n367), .B1(n4), .A0N(memory[56]), .A1N(n4), .Y(n575) );
  OAI2BB2X1 U335 ( .B0(n366), .B1(n4), .A0N(memory[57]), .A1N(n4), .Y(n574) );
  OAI2BB2X1 U336 ( .B0(n365), .B1(n4), .A0N(memory[58]), .A1N(n4), .Y(n573) );
  OAI2BB2X1 U337 ( .B0(n364), .B1(n4), .A0N(memory[59]), .A1N(n4), .Y(n572) );
  OAI2BB2X1 U338 ( .B0(n367), .B1(n5), .A0N(memory[72]), .A1N(n5), .Y(n559) );
  OAI2BB2X1 U339 ( .B0(n366), .B1(n5), .A0N(memory[73]), .A1N(n5), .Y(n558) );
  OAI2BB2X1 U340 ( .B0(n365), .B1(n5), .A0N(memory[74]), .A1N(n5), .Y(n557) );
  OAI2BB2X1 U341 ( .B0(n364), .B1(n5), .A0N(memory[75]), .A1N(n5), .Y(n556) );
  OAI2BB2X1 U342 ( .B0(n367), .B1(n6), .A0N(memory[88]), .A1N(n6), .Y(n543) );
  OAI2BB2X1 U343 ( .B0(n366), .B1(n6), .A0N(memory[89]), .A1N(n6), .Y(n542) );
  OAI2BB2X1 U344 ( .B0(n365), .B1(n6), .A0N(memory[90]), .A1N(n6), .Y(n541) );
  OAI2BB2X1 U345 ( .B0(n364), .B1(n6), .A0N(memory[91]), .A1N(n6), .Y(n540) );
  OAI2BB2X1 U346 ( .B0(n367), .B1(n7), .A0N(memory[104]), .A1N(n7), .Y(n527)
         );
  OAI2BB2X1 U347 ( .B0(n366), .B1(n7), .A0N(memory[105]), .A1N(n7), .Y(n526)
         );
  OAI2BB2X1 U348 ( .B0(n365), .B1(n7), .A0N(memory[106]), .A1N(n7), .Y(n525)
         );
  OAI2BB2X1 U349 ( .B0(n364), .B1(n7), .A0N(memory[107]), .A1N(n7), .Y(n524)
         );
  OAI2BB2X1 U350 ( .B0(n367), .B1(n8), .A0N(memory[120]), .A1N(n8), .Y(n511)
         );
  OAI2BB2X1 U351 ( .B0(n366), .B1(n8), .A0N(memory[121]), .A1N(n8), .Y(n510)
         );
  OAI2BB2X1 U352 ( .B0(n365), .B1(n8), .A0N(memory[122]), .A1N(n8), .Y(n509)
         );
  OAI2BB2X1 U353 ( .B0(n364), .B1(n8), .A0N(memory[123]), .A1N(n8), .Y(n508)
         );
  OAI2BB2X1 U354 ( .B0(n367), .B1(n9), .A0N(memory[136]), .A1N(n9), .Y(n495)
         );
  OAI2BB2X1 U355 ( .B0(n366), .B1(n9), .A0N(memory[137]), .A1N(n9), .Y(n494)
         );
  OAI2BB2X1 U356 ( .B0(n365), .B1(n9), .A0N(memory[138]), .A1N(n9), .Y(n493)
         );
  OAI2BB2X1 U357 ( .B0(n364), .B1(n9), .A0N(memory[139]), .A1N(n9), .Y(n492)
         );
  OAI2BB2X1 U358 ( .B0(n367), .B1(n10), .A0N(memory[152]), .A1N(n10), .Y(n479)
         );
  OAI2BB2X1 U359 ( .B0(n366), .B1(n10), .A0N(memory[153]), .A1N(n10), .Y(n478)
         );
  OAI2BB2X1 U360 ( .B0(n365), .B1(n10), .A0N(memory[154]), .A1N(n10), .Y(n477)
         );
  OAI2BB2X1 U361 ( .B0(n364), .B1(n10), .A0N(memory[155]), .A1N(n10), .Y(n476)
         );
  OAI2BB2X1 U362 ( .B0(n367), .B1(n11), .A0N(memory[168]), .A1N(n11), .Y(n463)
         );
  OAI2BB2X1 U363 ( .B0(n366), .B1(n11), .A0N(memory[169]), .A1N(n11), .Y(n462)
         );
  OAI2BB2X1 U364 ( .B0(n365), .B1(n11), .A0N(memory[170]), .A1N(n11), .Y(n461)
         );
  OAI2BB2X1 U365 ( .B0(n364), .B1(n11), .A0N(memory[171]), .A1N(n11), .Y(n460)
         );
  OAI2BB2X1 U366 ( .B0(n367), .B1(n12), .A0N(memory[184]), .A1N(n12), .Y(n447)
         );
  OAI2BB2X1 U367 ( .B0(n366), .B1(n12), .A0N(memory[185]), .A1N(n12), .Y(n446)
         );
  OAI2BB2X1 U368 ( .B0(n365), .B1(n12), .A0N(memory[186]), .A1N(n12), .Y(n445)
         );
  OAI2BB2X1 U369 ( .B0(n364), .B1(n12), .A0N(memory[187]), .A1N(n12), .Y(n444)
         );
  OAI2BB2X1 U370 ( .B0(n367), .B1(n13), .A0N(memory[200]), .A1N(n13), .Y(n431)
         );
  OAI2BB2X1 U371 ( .B0(n366), .B1(n13), .A0N(memory[201]), .A1N(n13), .Y(n430)
         );
  OAI2BB2X1 U372 ( .B0(n365), .B1(n13), .A0N(memory[202]), .A1N(n13), .Y(n429)
         );
  OAI2BB2X1 U373 ( .B0(n364), .B1(n13), .A0N(memory[203]), .A1N(n13), .Y(n428)
         );
  OAI2BB2X1 U374 ( .B0(n367), .B1(n14), .A0N(memory[216]), .A1N(n14), .Y(n415)
         );
  OAI2BB2X1 U375 ( .B0(n366), .B1(n14), .A0N(memory[217]), .A1N(n14), .Y(n414)
         );
  OAI2BB2X1 U376 ( .B0(n365), .B1(n14), .A0N(memory[218]), .A1N(n14), .Y(n413)
         );
  OAI2BB2X1 U377 ( .B0(n364), .B1(n14), .A0N(memory[219]), .A1N(n14), .Y(n412)
         );
  OAI2BB2X1 U378 ( .B0(n367), .B1(n15), .A0N(memory[232]), .A1N(n15), .Y(n399)
         );
  OAI2BB2X1 U379 ( .B0(n366), .B1(n15), .A0N(memory[233]), .A1N(n15), .Y(n398)
         );
  OAI2BB2X1 U380 ( .B0(n365), .B1(n15), .A0N(memory[234]), .A1N(n15), .Y(n397)
         );
  OAI2BB2X1 U381 ( .B0(n364), .B1(n15), .A0N(memory[235]), .A1N(n15), .Y(n396)
         );
  OAI2BB2X1 U382 ( .B0(n367), .B1(n16), .A0N(memory[248]), .A1N(n16), .Y(n383)
         );
  OAI2BB2X1 U383 ( .B0(n366), .B1(n16), .A0N(memory[249]), .A1N(n16), .Y(n382)
         );
  OAI2BB2X1 U384 ( .B0(n365), .B1(n16), .A0N(memory[250]), .A1N(n16), .Y(n381)
         );
  OAI2BB2X1 U385 ( .B0(n364), .B1(n16), .A0N(memory[251]), .A1N(n16), .Y(n380)
         );
  BUFX3 U386 ( .A(n632), .Y(n357) );
  NAND2BX1 U387 ( .AN(wr_rd), .B(en), .Y(n632) );
  NOR2BX1 U388 ( .AN(n636), .B(addr[3]), .Y(n633) );
  BUFX3 U389 ( .A(addr[2]), .Y(n355) );
  INVX1 U390 ( .A(addr[2]), .Y(n359) );
  AND2X2 U391 ( .A(wr_rd), .B(en), .Y(n636) );
  AND2X2 U392 ( .A(addr[3]), .B(n636), .Y(n637) );
  INVX1 U393 ( .A(din[0]), .Y(n375) );
  INVX1 U394 ( .A(din[1]), .Y(n374) );
  INVX1 U395 ( .A(din[2]), .Y(n373) );
  INVX1 U396 ( .A(din[3]), .Y(n372) );
  INVX1 U397 ( .A(din[4]), .Y(n371) );
  INVX1 U398 ( .A(din[5]), .Y(n370) );
  INVX1 U399 ( .A(din[6]), .Y(n369) );
  INVX1 U400 ( .A(din[7]), .Y(n368) );
  INVX1 U401 ( .A(din[8]), .Y(n367) );
  INVX1 U402 ( .A(din[9]), .Y(n366) );
  INVX1 U403 ( .A(din[10]), .Y(n365) );
  INVX1 U404 ( .A(din[11]), .Y(n364) );
  INVX1 U405 ( .A(din[12]), .Y(n363) );
  INVX1 U406 ( .A(din[13]), .Y(n362) );
  INVX1 U407 ( .A(din[14]), .Y(n361) );
  INVX1 U408 ( .A(din[15]), .Y(n360) );
endmodule


module mem4x4_2 ( clk, rstn, en, wr_rd, addr, din, dout );
  input [3:0] addr;
  input [15:0] din;
  output [15:0] dout;
  input clk, rstn, en, wr_rd;
  wire   N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48,
         N49, N50, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n23, n25, n27, n28, n30, n31, n34, n36,
         n38, n40, n41, n42, n43, n44, n46, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643;
  wire   [255:0] memory;

  DFFRHQX1 memory_reg_1__15_ ( .D(n392), .CK(clk), .RN(rstn), .Q(memory[239])
         );
  DFFRHQX1 memory_reg_1__14_ ( .D(n393), .CK(clk), .RN(rstn), .Q(memory[238])
         );
  DFFRHQX1 memory_reg_1__13_ ( .D(n394), .CK(clk), .RN(rstn), .Q(memory[237])
         );
  DFFRHQX1 memory_reg_1__12_ ( .D(n395), .CK(clk), .RN(rstn), .Q(memory[236])
         );
  DFFRHQX1 memory_reg_1__11_ ( .D(n396), .CK(clk), .RN(rstn), .Q(memory[235])
         );
  DFFRHQX1 memory_reg_1__10_ ( .D(n397), .CK(clk), .RN(rstn), .Q(memory[234])
         );
  DFFRHQX1 memory_reg_1__9_ ( .D(n398), .CK(clk), .RN(rstn), .Q(memory[233])
         );
  DFFRHQX1 memory_reg_1__8_ ( .D(n399), .CK(clk), .RN(rstn), .Q(memory[232])
         );
  DFFRHQX1 memory_reg_1__7_ ( .D(n400), .CK(clk), .RN(rstn), .Q(memory[231])
         );
  DFFRHQX1 memory_reg_1__6_ ( .D(n401), .CK(clk), .RN(rstn), .Q(memory[230])
         );
  DFFRHQX1 memory_reg_1__5_ ( .D(n402), .CK(clk), .RN(rstn), .Q(memory[229])
         );
  DFFRHQX1 memory_reg_1__4_ ( .D(n403), .CK(clk), .RN(rstn), .Q(memory[228])
         );
  DFFRHQX1 memory_reg_1__3_ ( .D(n404), .CK(clk), .RN(rstn), .Q(memory[227])
         );
  DFFRHQX1 memory_reg_1__2_ ( .D(n405), .CK(clk), .RN(rstn), .Q(memory[226])
         );
  DFFRHQX1 memory_reg_1__1_ ( .D(n406), .CK(clk), .RN(rstn), .Q(memory[225])
         );
  DFFRHQX1 memory_reg_1__0_ ( .D(n407), .CK(clk), .RN(rstn), .Q(memory[224])
         );
  DFFRHQX1 memory_reg_5__15_ ( .D(n456), .CK(clk), .RN(rstn), .Q(memory[175])
         );
  DFFRHQX1 memory_reg_5__14_ ( .D(n457), .CK(clk), .RN(rstn), .Q(memory[174])
         );
  DFFRHQX1 memory_reg_5__13_ ( .D(n458), .CK(clk), .RN(rstn), .Q(memory[173])
         );
  DFFRHQX1 memory_reg_5__12_ ( .D(n459), .CK(clk), .RN(rstn), .Q(memory[172])
         );
  DFFRHQX1 memory_reg_5__11_ ( .D(n460), .CK(clk), .RN(rstn), .Q(memory[171])
         );
  DFFRHQX1 memory_reg_5__10_ ( .D(n461), .CK(clk), .RN(rstn), .Q(memory[170])
         );
  DFFRHQX1 memory_reg_5__9_ ( .D(n462), .CK(clk), .RN(rstn), .Q(memory[169])
         );
  DFFRHQX1 memory_reg_5__8_ ( .D(n463), .CK(clk), .RN(rstn), .Q(memory[168])
         );
  DFFRHQX1 memory_reg_5__7_ ( .D(n464), .CK(clk), .RN(rstn), .Q(memory[167])
         );
  DFFRHQX1 memory_reg_5__6_ ( .D(n465), .CK(clk), .RN(rstn), .Q(memory[166])
         );
  DFFRHQX1 memory_reg_5__5_ ( .D(n466), .CK(clk), .RN(rstn), .Q(memory[165])
         );
  DFFRHQX1 memory_reg_5__4_ ( .D(n467), .CK(clk), .RN(rstn), .Q(memory[164])
         );
  DFFRHQX1 memory_reg_5__3_ ( .D(n468), .CK(clk), .RN(rstn), .Q(memory[163])
         );
  DFFRHQX1 memory_reg_5__2_ ( .D(n469), .CK(clk), .RN(rstn), .Q(memory[162])
         );
  DFFRHQX1 memory_reg_5__1_ ( .D(n470), .CK(clk), .RN(rstn), .Q(memory[161])
         );
  DFFRHQX1 memory_reg_5__0_ ( .D(n471), .CK(clk), .RN(rstn), .Q(memory[160])
         );
  DFFRHQX1 memory_reg_9__15_ ( .D(n520), .CK(clk), .RN(rstn), .Q(memory[111])
         );
  DFFRHQX1 memory_reg_9__14_ ( .D(n521), .CK(clk), .RN(rstn), .Q(memory[110])
         );
  DFFRHQX1 memory_reg_9__13_ ( .D(n522), .CK(clk), .RN(rstn), .Q(memory[109])
         );
  DFFRHQX1 memory_reg_9__12_ ( .D(n523), .CK(clk), .RN(rstn), .Q(memory[108])
         );
  DFFRHQX1 memory_reg_9__11_ ( .D(n524), .CK(clk), .RN(rstn), .Q(memory[107])
         );
  DFFRHQX1 memory_reg_9__10_ ( .D(n525), .CK(clk), .RN(rstn), .Q(memory[106])
         );
  DFFRHQX1 memory_reg_9__9_ ( .D(n526), .CK(clk), .RN(rstn), .Q(memory[105])
         );
  DFFRHQX1 memory_reg_9__8_ ( .D(n527), .CK(clk), .RN(rstn), .Q(memory[104])
         );
  DFFRHQX1 memory_reg_9__7_ ( .D(n528), .CK(clk), .RN(rstn), .Q(memory[103])
         );
  DFFRHQX1 memory_reg_9__6_ ( .D(n529), .CK(clk), .RN(rstn), .Q(memory[102])
         );
  DFFRHQX1 memory_reg_9__5_ ( .D(n530), .CK(clk), .RN(rstn), .Q(memory[101])
         );
  DFFRHQX1 memory_reg_9__4_ ( .D(n531), .CK(clk), .RN(rstn), .Q(memory[100])
         );
  DFFRHQX1 memory_reg_9__3_ ( .D(n532), .CK(clk), .RN(rstn), .Q(memory[99]) );
  DFFRHQX1 memory_reg_9__2_ ( .D(n533), .CK(clk), .RN(rstn), .Q(memory[98]) );
  DFFRHQX1 memory_reg_9__1_ ( .D(n534), .CK(clk), .RN(rstn), .Q(memory[97]) );
  DFFRHQX1 memory_reg_9__0_ ( .D(n535), .CK(clk), .RN(rstn), .Q(memory[96]) );
  DFFRHQX1 memory_reg_13__15_ ( .D(n584), .CK(clk), .RN(rstn), .Q(memory[47])
         );
  DFFRHQX1 memory_reg_13__14_ ( .D(n585), .CK(clk), .RN(rstn), .Q(memory[46])
         );
  DFFRHQX1 memory_reg_13__13_ ( .D(n586), .CK(clk), .RN(rstn), .Q(memory[45])
         );
  DFFRHQX1 memory_reg_13__12_ ( .D(n587), .CK(clk), .RN(rstn), .Q(memory[44])
         );
  DFFRHQX1 memory_reg_13__11_ ( .D(n588), .CK(clk), .RN(rstn), .Q(memory[43])
         );
  DFFRHQX1 memory_reg_13__10_ ( .D(n589), .CK(clk), .RN(rstn), .Q(memory[42])
         );
  DFFRHQX1 memory_reg_13__9_ ( .D(n590), .CK(clk), .RN(rstn), .Q(memory[41])
         );
  DFFRHQX1 memory_reg_13__8_ ( .D(n591), .CK(clk), .RN(rstn), .Q(memory[40])
         );
  DFFRHQX1 memory_reg_13__7_ ( .D(n592), .CK(clk), .RN(rstn), .Q(memory[39])
         );
  DFFRHQX1 memory_reg_13__6_ ( .D(n593), .CK(clk), .RN(rstn), .Q(memory[38])
         );
  DFFRHQX1 memory_reg_13__5_ ( .D(n594), .CK(clk), .RN(rstn), .Q(memory[37])
         );
  DFFRHQX1 memory_reg_13__4_ ( .D(n595), .CK(clk), .RN(rstn), .Q(memory[36])
         );
  DFFRHQX1 memory_reg_13__3_ ( .D(n596), .CK(clk), .RN(rstn), .Q(memory[35])
         );
  DFFRHQX1 memory_reg_13__2_ ( .D(n597), .CK(clk), .RN(rstn), .Q(memory[34])
         );
  DFFRHQX1 memory_reg_13__1_ ( .D(n598), .CK(clk), .RN(rstn), .Q(memory[33])
         );
  DFFRHQX1 memory_reg_13__0_ ( .D(n599), .CK(clk), .RN(rstn), .Q(memory[32])
         );
  DFFRHQX1 memory_reg_3__15_ ( .D(n424), .CK(clk), .RN(rstn), .Q(memory[207])
         );
  DFFRHQX1 memory_reg_3__14_ ( .D(n425), .CK(clk), .RN(rstn), .Q(memory[206])
         );
  DFFRHQX1 memory_reg_3__13_ ( .D(n426), .CK(clk), .RN(rstn), .Q(memory[205])
         );
  DFFRHQX1 memory_reg_3__12_ ( .D(n427), .CK(clk), .RN(rstn), .Q(memory[204])
         );
  DFFRHQX1 memory_reg_3__11_ ( .D(n428), .CK(clk), .RN(rstn), .Q(memory[203])
         );
  DFFRHQX1 memory_reg_3__10_ ( .D(n429), .CK(clk), .RN(rstn), .Q(memory[202])
         );
  DFFRHQX1 memory_reg_3__9_ ( .D(n430), .CK(clk), .RN(rstn), .Q(memory[201])
         );
  DFFRHQX1 memory_reg_3__8_ ( .D(n431), .CK(clk), .RN(rstn), .Q(memory[200])
         );
  DFFRHQX1 memory_reg_3__7_ ( .D(n432), .CK(clk), .RN(rstn), .Q(memory[199])
         );
  DFFRHQX1 memory_reg_3__6_ ( .D(n433), .CK(clk), .RN(rstn), .Q(memory[198])
         );
  DFFRHQX1 memory_reg_3__5_ ( .D(n434), .CK(clk), .RN(rstn), .Q(memory[197])
         );
  DFFRHQX1 memory_reg_3__4_ ( .D(n435), .CK(clk), .RN(rstn), .Q(memory[196])
         );
  DFFRHQX1 memory_reg_3__3_ ( .D(n436), .CK(clk), .RN(rstn), .Q(memory[195])
         );
  DFFRHQX1 memory_reg_3__2_ ( .D(n437), .CK(clk), .RN(rstn), .Q(memory[194])
         );
  DFFRHQX1 memory_reg_3__1_ ( .D(n438), .CK(clk), .RN(rstn), .Q(memory[193])
         );
  DFFRHQX1 memory_reg_3__0_ ( .D(n439), .CK(clk), .RN(rstn), .Q(memory[192])
         );
  DFFRHQX1 memory_reg_7__15_ ( .D(n488), .CK(clk), .RN(rstn), .Q(memory[143])
         );
  DFFRHQX1 memory_reg_7__14_ ( .D(n489), .CK(clk), .RN(rstn), .Q(memory[142])
         );
  DFFRHQX1 memory_reg_7__13_ ( .D(n490), .CK(clk), .RN(rstn), .Q(memory[141])
         );
  DFFRHQX1 memory_reg_7__12_ ( .D(n491), .CK(clk), .RN(rstn), .Q(memory[140])
         );
  DFFRHQX1 memory_reg_7__11_ ( .D(n492), .CK(clk), .RN(rstn), .Q(memory[139])
         );
  DFFRHQX1 memory_reg_7__10_ ( .D(n493), .CK(clk), .RN(rstn), .Q(memory[138])
         );
  DFFRHQX1 memory_reg_7__9_ ( .D(n494), .CK(clk), .RN(rstn), .Q(memory[137])
         );
  DFFRHQX1 memory_reg_7__8_ ( .D(n495), .CK(clk), .RN(rstn), .Q(memory[136])
         );
  DFFRHQX1 memory_reg_7__7_ ( .D(n496), .CK(clk), .RN(rstn), .Q(memory[135])
         );
  DFFRHQX1 memory_reg_7__6_ ( .D(n497), .CK(clk), .RN(rstn), .Q(memory[134])
         );
  DFFRHQX1 memory_reg_7__5_ ( .D(n498), .CK(clk), .RN(rstn), .Q(memory[133])
         );
  DFFRHQX1 memory_reg_7__4_ ( .D(n499), .CK(clk), .RN(rstn), .Q(memory[132])
         );
  DFFRHQX1 memory_reg_7__3_ ( .D(n500), .CK(clk), .RN(rstn), .Q(memory[131])
         );
  DFFRHQX1 memory_reg_7__2_ ( .D(n501), .CK(clk), .RN(rstn), .Q(memory[130])
         );
  DFFRHQX1 memory_reg_7__1_ ( .D(n502), .CK(clk), .RN(rstn), .Q(memory[129])
         );
  DFFRHQX1 memory_reg_7__0_ ( .D(n503), .CK(clk), .RN(rstn), .Q(memory[128])
         );
  DFFRHQX1 memory_reg_11__15_ ( .D(n552), .CK(clk), .RN(rstn), .Q(memory[79])
         );
  DFFRHQX1 memory_reg_11__14_ ( .D(n553), .CK(clk), .RN(rstn), .Q(memory[78])
         );
  DFFRHQX1 memory_reg_11__13_ ( .D(n554), .CK(clk), .RN(rstn), .Q(memory[77])
         );
  DFFRHQX1 memory_reg_11__12_ ( .D(n555), .CK(clk), .RN(rstn), .Q(memory[76])
         );
  DFFRHQX1 memory_reg_11__11_ ( .D(n556), .CK(clk), .RN(rstn), .Q(memory[75])
         );
  DFFRHQX1 memory_reg_11__10_ ( .D(n557), .CK(clk), .RN(rstn), .Q(memory[74])
         );
  DFFRHQX1 memory_reg_11__9_ ( .D(n558), .CK(clk), .RN(rstn), .Q(memory[73])
         );
  DFFRHQX1 memory_reg_11__8_ ( .D(n559), .CK(clk), .RN(rstn), .Q(memory[72])
         );
  DFFRHQX1 memory_reg_11__7_ ( .D(n560), .CK(clk), .RN(rstn), .Q(memory[71])
         );
  DFFRHQX1 memory_reg_11__6_ ( .D(n561), .CK(clk), .RN(rstn), .Q(memory[70])
         );
  DFFRHQX1 memory_reg_11__5_ ( .D(n562), .CK(clk), .RN(rstn), .Q(memory[69])
         );
  DFFRHQX1 memory_reg_11__4_ ( .D(n563), .CK(clk), .RN(rstn), .Q(memory[68])
         );
  DFFRHQX1 memory_reg_11__3_ ( .D(n564), .CK(clk), .RN(rstn), .Q(memory[67])
         );
  DFFRHQX1 memory_reg_11__2_ ( .D(n565), .CK(clk), .RN(rstn), .Q(memory[66])
         );
  DFFRHQX1 memory_reg_11__1_ ( .D(n566), .CK(clk), .RN(rstn), .Q(memory[65])
         );
  DFFRHQX1 memory_reg_11__0_ ( .D(n567), .CK(clk), .RN(rstn), .Q(memory[64])
         );
  DFFRHQX1 memory_reg_15__15_ ( .D(n616), .CK(clk), .RN(rstn), .Q(memory[15])
         );
  DFFRHQX1 memory_reg_15__14_ ( .D(n617), .CK(clk), .RN(rstn), .Q(memory[14])
         );
  DFFRHQX1 memory_reg_15__13_ ( .D(n618), .CK(clk), .RN(rstn), .Q(memory[13])
         );
  DFFRHQX1 memory_reg_15__12_ ( .D(n619), .CK(clk), .RN(rstn), .Q(memory[12])
         );
  DFFRHQX1 memory_reg_15__11_ ( .D(n620), .CK(clk), .RN(rstn), .Q(memory[11])
         );
  DFFRHQX1 memory_reg_15__10_ ( .D(n621), .CK(clk), .RN(rstn), .Q(memory[10])
         );
  DFFRHQX1 memory_reg_15__9_ ( .D(n622), .CK(clk), .RN(rstn), .Q(memory[9]) );
  DFFRHQX1 memory_reg_15__8_ ( .D(n623), .CK(clk), .RN(rstn), .Q(memory[8]) );
  DFFRHQX1 memory_reg_15__7_ ( .D(n624), .CK(clk), .RN(rstn), .Q(memory[7]) );
  DFFRHQX1 memory_reg_15__6_ ( .D(n625), .CK(clk), .RN(rstn), .Q(memory[6]) );
  DFFRHQX1 memory_reg_15__5_ ( .D(n626), .CK(clk), .RN(rstn), .Q(memory[5]) );
  DFFRHQX1 memory_reg_15__4_ ( .D(n627), .CK(clk), .RN(rstn), .Q(memory[4]) );
  DFFRHQX1 memory_reg_15__3_ ( .D(n628), .CK(clk), .RN(rstn), .Q(memory[3]) );
  DFFRHQX1 memory_reg_15__2_ ( .D(n629), .CK(clk), .RN(rstn), .Q(memory[2]) );
  DFFRHQX1 memory_reg_15__1_ ( .D(n630), .CK(clk), .RN(rstn), .Q(memory[1]) );
  DFFRHQX1 memory_reg_15__0_ ( .D(n631), .CK(clk), .RN(rstn), .Q(memory[0]) );
  DFFRHQX1 memory_reg_0__15_ ( .D(n376), .CK(clk), .RN(rstn), .Q(memory[255])
         );
  DFFRHQX1 memory_reg_0__14_ ( .D(n377), .CK(clk), .RN(rstn), .Q(memory[254])
         );
  DFFRHQX1 memory_reg_0__13_ ( .D(n378), .CK(clk), .RN(rstn), .Q(memory[253])
         );
  DFFRHQX1 memory_reg_0__12_ ( .D(n379), .CK(clk), .RN(rstn), .Q(memory[252])
         );
  DFFRHQX1 memory_reg_0__11_ ( .D(n380), .CK(clk), .RN(rstn), .Q(memory[251])
         );
  DFFRHQX1 memory_reg_0__10_ ( .D(n381), .CK(clk), .RN(rstn), .Q(memory[250])
         );
  DFFRHQX1 memory_reg_0__9_ ( .D(n382), .CK(clk), .RN(rstn), .Q(memory[249])
         );
  DFFRHQX1 memory_reg_0__8_ ( .D(n383), .CK(clk), .RN(rstn), .Q(memory[248])
         );
  DFFRHQX1 memory_reg_0__7_ ( .D(n384), .CK(clk), .RN(rstn), .Q(memory[247])
         );
  DFFRHQX1 memory_reg_0__6_ ( .D(n385), .CK(clk), .RN(rstn), .Q(memory[246])
         );
  DFFRHQX1 memory_reg_0__5_ ( .D(n386), .CK(clk), .RN(rstn), .Q(memory[245])
         );
  DFFRHQX1 memory_reg_0__4_ ( .D(n387), .CK(clk), .RN(rstn), .Q(memory[244])
         );
  DFFRHQX1 memory_reg_0__3_ ( .D(n388), .CK(clk), .RN(rstn), .Q(memory[243])
         );
  DFFRHQX1 memory_reg_0__2_ ( .D(n389), .CK(clk), .RN(rstn), .Q(memory[242])
         );
  DFFRHQX1 memory_reg_0__1_ ( .D(n390), .CK(clk), .RN(rstn), .Q(memory[241])
         );
  DFFRHQX1 memory_reg_0__0_ ( .D(n391), .CK(clk), .RN(rstn), .Q(memory[240])
         );
  DFFRHQX1 memory_reg_4__15_ ( .D(n440), .CK(clk), .RN(rstn), .Q(memory[191])
         );
  DFFRHQX1 memory_reg_4__14_ ( .D(n441), .CK(clk), .RN(rstn), .Q(memory[190])
         );
  DFFRHQX1 memory_reg_4__13_ ( .D(n442), .CK(clk), .RN(rstn), .Q(memory[189])
         );
  DFFRHQX1 memory_reg_4__12_ ( .D(n443), .CK(clk), .RN(rstn), .Q(memory[188])
         );
  DFFRHQX1 memory_reg_4__11_ ( .D(n444), .CK(clk), .RN(rstn), .Q(memory[187])
         );
  DFFRHQX1 memory_reg_4__10_ ( .D(n445), .CK(clk), .RN(rstn), .Q(memory[186])
         );
  DFFRHQX1 memory_reg_4__9_ ( .D(n446), .CK(clk), .RN(rstn), .Q(memory[185])
         );
  DFFRHQX1 memory_reg_4__8_ ( .D(n447), .CK(clk), .RN(rstn), .Q(memory[184])
         );
  DFFRHQX1 memory_reg_4__7_ ( .D(n448), .CK(clk), .RN(rstn), .Q(memory[183])
         );
  DFFRHQX1 memory_reg_4__6_ ( .D(n449), .CK(clk), .RN(rstn), .Q(memory[182])
         );
  DFFRHQX1 memory_reg_4__5_ ( .D(n450), .CK(clk), .RN(rstn), .Q(memory[181])
         );
  DFFRHQX1 memory_reg_4__4_ ( .D(n451), .CK(clk), .RN(rstn), .Q(memory[180])
         );
  DFFRHQX1 memory_reg_4__3_ ( .D(n452), .CK(clk), .RN(rstn), .Q(memory[179])
         );
  DFFRHQX1 memory_reg_4__2_ ( .D(n453), .CK(clk), .RN(rstn), .Q(memory[178])
         );
  DFFRHQX1 memory_reg_4__1_ ( .D(n454), .CK(clk), .RN(rstn), .Q(memory[177])
         );
  DFFRHQX1 memory_reg_4__0_ ( .D(n455), .CK(clk), .RN(rstn), .Q(memory[176])
         );
  DFFRHQX1 memory_reg_8__15_ ( .D(n504), .CK(clk), .RN(rstn), .Q(memory[127])
         );
  DFFRHQX1 memory_reg_8__14_ ( .D(n505), .CK(clk), .RN(rstn), .Q(memory[126])
         );
  DFFRHQX1 memory_reg_8__13_ ( .D(n506), .CK(clk), .RN(rstn), .Q(memory[125])
         );
  DFFRHQX1 memory_reg_8__12_ ( .D(n507), .CK(clk), .RN(rstn), .Q(memory[124])
         );
  DFFRHQX1 memory_reg_8__11_ ( .D(n508), .CK(clk), .RN(rstn), .Q(memory[123])
         );
  DFFRHQX1 memory_reg_8__10_ ( .D(n509), .CK(clk), .RN(rstn), .Q(memory[122])
         );
  DFFRHQX1 memory_reg_8__9_ ( .D(n510), .CK(clk), .RN(rstn), .Q(memory[121])
         );
  DFFRHQX1 memory_reg_8__8_ ( .D(n511), .CK(clk), .RN(rstn), .Q(memory[120])
         );
  DFFRHQX1 memory_reg_8__7_ ( .D(n512), .CK(clk), .RN(rstn), .Q(memory[119])
         );
  DFFRHQX1 memory_reg_8__6_ ( .D(n513), .CK(clk), .RN(rstn), .Q(memory[118])
         );
  DFFRHQX1 memory_reg_8__5_ ( .D(n514), .CK(clk), .RN(rstn), .Q(memory[117])
         );
  DFFRHQX1 memory_reg_8__4_ ( .D(n515), .CK(clk), .RN(rstn), .Q(memory[116])
         );
  DFFRHQX1 memory_reg_8__3_ ( .D(n516), .CK(clk), .RN(rstn), .Q(memory[115])
         );
  DFFRHQX1 memory_reg_8__2_ ( .D(n517), .CK(clk), .RN(rstn), .Q(memory[114])
         );
  DFFRHQX1 memory_reg_8__1_ ( .D(n518), .CK(clk), .RN(rstn), .Q(memory[113])
         );
  DFFRHQX1 memory_reg_8__0_ ( .D(n519), .CK(clk), .RN(rstn), .Q(memory[112])
         );
  DFFRHQX1 memory_reg_12__15_ ( .D(n568), .CK(clk), .RN(rstn), .Q(memory[63])
         );
  DFFRHQX1 memory_reg_12__14_ ( .D(n569), .CK(clk), .RN(rstn), .Q(memory[62])
         );
  DFFRHQX1 memory_reg_12__13_ ( .D(n570), .CK(clk), .RN(rstn), .Q(memory[61])
         );
  DFFRHQX1 memory_reg_12__12_ ( .D(n571), .CK(clk), .RN(rstn), .Q(memory[60])
         );
  DFFRHQX1 memory_reg_12__11_ ( .D(n572), .CK(clk), .RN(rstn), .Q(memory[59])
         );
  DFFRHQX1 memory_reg_12__10_ ( .D(n573), .CK(clk), .RN(rstn), .Q(memory[58])
         );
  DFFRHQX1 memory_reg_12__9_ ( .D(n574), .CK(clk), .RN(rstn), .Q(memory[57])
         );
  DFFRHQX1 memory_reg_12__8_ ( .D(n575), .CK(clk), .RN(rstn), .Q(memory[56])
         );
  DFFRHQX1 memory_reg_12__7_ ( .D(n576), .CK(clk), .RN(rstn), .Q(memory[55])
         );
  DFFRHQX1 memory_reg_12__6_ ( .D(n577), .CK(clk), .RN(rstn), .Q(memory[54])
         );
  DFFRHQX1 memory_reg_12__5_ ( .D(n578), .CK(clk), .RN(rstn), .Q(memory[53])
         );
  DFFRHQX1 memory_reg_12__4_ ( .D(n579), .CK(clk), .RN(rstn), .Q(memory[52])
         );
  DFFRHQX1 memory_reg_12__3_ ( .D(n580), .CK(clk), .RN(rstn), .Q(memory[51])
         );
  DFFRHQX1 memory_reg_12__2_ ( .D(n581), .CK(clk), .RN(rstn), .Q(memory[50])
         );
  DFFRHQX1 memory_reg_12__1_ ( .D(n582), .CK(clk), .RN(rstn), .Q(memory[49])
         );
  DFFRHQX1 memory_reg_12__0_ ( .D(n583), .CK(clk), .RN(rstn), .Q(memory[48])
         );
  DFFRHQX1 memory_reg_2__15_ ( .D(n408), .CK(clk), .RN(rstn), .Q(memory[223])
         );
  DFFRHQX1 memory_reg_2__14_ ( .D(n409), .CK(clk), .RN(rstn), .Q(memory[222])
         );
  DFFRHQX1 memory_reg_2__13_ ( .D(n410), .CK(clk), .RN(rstn), .Q(memory[221])
         );
  DFFRHQX1 memory_reg_2__12_ ( .D(n411), .CK(clk), .RN(rstn), .Q(memory[220])
         );
  DFFRHQX1 memory_reg_2__11_ ( .D(n412), .CK(clk), .RN(rstn), .Q(memory[219])
         );
  DFFRHQX1 memory_reg_2__10_ ( .D(n413), .CK(clk), .RN(rstn), .Q(memory[218])
         );
  DFFRHQX1 memory_reg_2__9_ ( .D(n414), .CK(clk), .RN(rstn), .Q(memory[217])
         );
  DFFRHQX1 memory_reg_2__8_ ( .D(n415), .CK(clk), .RN(rstn), .Q(memory[216])
         );
  DFFRHQX1 memory_reg_2__7_ ( .D(n416), .CK(clk), .RN(rstn), .Q(memory[215])
         );
  DFFRHQX1 memory_reg_2__6_ ( .D(n417), .CK(clk), .RN(rstn), .Q(memory[214])
         );
  DFFRHQX1 memory_reg_2__5_ ( .D(n418), .CK(clk), .RN(rstn), .Q(memory[213])
         );
  DFFRHQX1 memory_reg_2__4_ ( .D(n419), .CK(clk), .RN(rstn), .Q(memory[212])
         );
  DFFRHQX1 memory_reg_2__3_ ( .D(n420), .CK(clk), .RN(rstn), .Q(memory[211])
         );
  DFFRHQX1 memory_reg_2__2_ ( .D(n421), .CK(clk), .RN(rstn), .Q(memory[210])
         );
  DFFRHQX1 memory_reg_2__1_ ( .D(n422), .CK(clk), .RN(rstn), .Q(memory[209])
         );
  DFFRHQX1 memory_reg_2__0_ ( .D(n423), .CK(clk), .RN(rstn), .Q(memory[208])
         );
  DFFRHQX1 memory_reg_6__15_ ( .D(n472), .CK(clk), .RN(rstn), .Q(memory[159])
         );
  DFFRHQX1 memory_reg_6__14_ ( .D(n473), .CK(clk), .RN(rstn), .Q(memory[158])
         );
  DFFRHQX1 memory_reg_6__13_ ( .D(n474), .CK(clk), .RN(rstn), .Q(memory[157])
         );
  DFFRHQX1 memory_reg_6__12_ ( .D(n475), .CK(clk), .RN(rstn), .Q(memory[156])
         );
  DFFRHQX1 memory_reg_6__11_ ( .D(n476), .CK(clk), .RN(rstn), .Q(memory[155])
         );
  DFFRHQX1 memory_reg_6__10_ ( .D(n477), .CK(clk), .RN(rstn), .Q(memory[154])
         );
  DFFRHQX1 memory_reg_6__9_ ( .D(n478), .CK(clk), .RN(rstn), .Q(memory[153])
         );
  DFFRHQX1 memory_reg_6__8_ ( .D(n479), .CK(clk), .RN(rstn), .Q(memory[152])
         );
  DFFRHQX1 memory_reg_6__7_ ( .D(n480), .CK(clk), .RN(rstn), .Q(memory[151])
         );
  DFFRHQX1 memory_reg_6__6_ ( .D(n481), .CK(clk), .RN(rstn), .Q(memory[150])
         );
  DFFRHQX1 memory_reg_6__5_ ( .D(n482), .CK(clk), .RN(rstn), .Q(memory[149])
         );
  DFFRHQX1 memory_reg_6__4_ ( .D(n483), .CK(clk), .RN(rstn), .Q(memory[148])
         );
  DFFRHQX1 memory_reg_6__3_ ( .D(n484), .CK(clk), .RN(rstn), .Q(memory[147])
         );
  DFFRHQX1 memory_reg_6__2_ ( .D(n485), .CK(clk), .RN(rstn), .Q(memory[146])
         );
  DFFRHQX1 memory_reg_6__1_ ( .D(n486), .CK(clk), .RN(rstn), .Q(memory[145])
         );
  DFFRHQX1 memory_reg_6__0_ ( .D(n487), .CK(clk), .RN(rstn), .Q(memory[144])
         );
  DFFRHQX1 memory_reg_10__15_ ( .D(n536), .CK(clk), .RN(rstn), .Q(memory[95])
         );
  DFFRHQX1 memory_reg_10__14_ ( .D(n537), .CK(clk), .RN(rstn), .Q(memory[94])
         );
  DFFRHQX1 memory_reg_10__13_ ( .D(n538), .CK(clk), .RN(rstn), .Q(memory[93])
         );
  DFFRHQX1 memory_reg_10__12_ ( .D(n539), .CK(clk), .RN(rstn), .Q(memory[92])
         );
  DFFRHQX1 memory_reg_10__11_ ( .D(n540), .CK(clk), .RN(rstn), .Q(memory[91])
         );
  DFFRHQX1 memory_reg_10__10_ ( .D(n541), .CK(clk), .RN(rstn), .Q(memory[90])
         );
  DFFRHQX1 memory_reg_10__9_ ( .D(n542), .CK(clk), .RN(rstn), .Q(memory[89])
         );
  DFFRHQX1 memory_reg_10__8_ ( .D(n543), .CK(clk), .RN(rstn), .Q(memory[88])
         );
  DFFRHQX1 memory_reg_10__7_ ( .D(n544), .CK(clk), .RN(rstn), .Q(memory[87])
         );
  DFFRHQX1 memory_reg_10__6_ ( .D(n545), .CK(clk), .RN(rstn), .Q(memory[86])
         );
  DFFRHQX1 memory_reg_10__5_ ( .D(n546), .CK(clk), .RN(rstn), .Q(memory[85])
         );
  DFFRHQX1 memory_reg_10__4_ ( .D(n547), .CK(clk), .RN(rstn), .Q(memory[84])
         );
  DFFRHQX1 memory_reg_10__3_ ( .D(n548), .CK(clk), .RN(rstn), .Q(memory[83])
         );
  DFFRHQX1 memory_reg_10__2_ ( .D(n549), .CK(clk), .RN(rstn), .Q(memory[82])
         );
  DFFRHQX1 memory_reg_10__1_ ( .D(n550), .CK(clk), .RN(rstn), .Q(memory[81])
         );
  DFFRHQX1 memory_reg_10__0_ ( .D(n551), .CK(clk), .RN(rstn), .Q(memory[80])
         );
  DFFRHQX1 memory_reg_14__15_ ( .D(n600), .CK(clk), .RN(rstn), .Q(memory[31])
         );
  DFFRHQX1 memory_reg_14__14_ ( .D(n601), .CK(clk), .RN(rstn), .Q(memory[30])
         );
  DFFRHQX1 memory_reg_14__13_ ( .D(n602), .CK(clk), .RN(rstn), .Q(memory[29])
         );
  DFFRHQX1 memory_reg_14__12_ ( .D(n603), .CK(clk), .RN(rstn), .Q(memory[28])
         );
  DFFRHQX1 memory_reg_14__11_ ( .D(n604), .CK(clk), .RN(rstn), .Q(memory[27])
         );
  DFFRHQX1 memory_reg_14__10_ ( .D(n605), .CK(clk), .RN(rstn), .Q(memory[26])
         );
  DFFRHQX1 memory_reg_14__9_ ( .D(n606), .CK(clk), .RN(rstn), .Q(memory[25])
         );
  DFFRHQX1 memory_reg_14__8_ ( .D(n607), .CK(clk), .RN(rstn), .Q(memory[24])
         );
  DFFRHQX1 memory_reg_14__7_ ( .D(n608), .CK(clk), .RN(rstn), .Q(memory[23])
         );
  DFFRHQX1 memory_reg_14__6_ ( .D(n609), .CK(clk), .RN(rstn), .Q(memory[22])
         );
  DFFRHQX1 memory_reg_14__5_ ( .D(n610), .CK(clk), .RN(rstn), .Q(memory[21])
         );
  DFFRHQX1 memory_reg_14__4_ ( .D(n611), .CK(clk), .RN(rstn), .Q(memory[20])
         );
  DFFRHQX1 memory_reg_14__3_ ( .D(n612), .CK(clk), .RN(rstn), .Q(memory[19])
         );
  DFFRHQX1 memory_reg_14__2_ ( .D(n613), .CK(clk), .RN(rstn), .Q(memory[18])
         );
  DFFRHQX1 memory_reg_14__1_ ( .D(n614), .CK(clk), .RN(rstn), .Q(memory[17])
         );
  DFFRHQX1 memory_reg_14__0_ ( .D(n615), .CK(clk), .RN(rstn), .Q(memory[16])
         );
  NAND2X1 U2 ( .A(n643), .B(n642), .Y(n1) );
  NAND2X1 U3 ( .A(n641), .B(n643), .Y(n2) );
  NAND2X1 U4 ( .A(n640), .B(n642), .Y(n3) );
  NAND2X1 U5 ( .A(n640), .B(n641), .Y(n4) );
  NAND2X1 U6 ( .A(n639), .B(n642), .Y(n5) );
  NAND2X1 U7 ( .A(n639), .B(n641), .Y(n6) );
  NAND2X1 U8 ( .A(n638), .B(n642), .Y(n7) );
  NAND2X1 U9 ( .A(n638), .B(n641), .Y(n8) );
  NAND2X1 U10 ( .A(n635), .B(n643), .Y(n9) );
  NAND2X1 U11 ( .A(n634), .B(n643), .Y(n10) );
  NAND2X1 U12 ( .A(n635), .B(n640), .Y(n11) );
  NAND2X1 U13 ( .A(n634), .B(n640), .Y(n12) );
  NAND2X1 U14 ( .A(n635), .B(n639), .Y(n13) );
  NAND2X1 U15 ( .A(n634), .B(n639), .Y(n14) );
  NAND2X1 U16 ( .A(n635), .B(n638), .Y(n15) );
  NAND2X1 U17 ( .A(n634), .B(n638), .Y(n16) );
  INVX1 U18 ( .A(n357), .Y(n351) );
  INVX1 U19 ( .A(n357), .Y(n352) );
  INVX1 U20 ( .A(n357), .Y(n353) );
  INVX1 U21 ( .A(n358), .Y(n349) );
  INVX1 U22 ( .A(n358), .Y(n350) );
  NOR2X1 U23 ( .A(n359), .B(addr[1]), .Y(n640) );
  NOR2X1 U24 ( .A(n359), .B(n358), .Y(n643) );
  AND2X2 U25 ( .A(n633), .B(addr[0]), .Y(n635) );
  AND2X2 U26 ( .A(n633), .B(n357), .Y(n634) );
  AND2X2 U27 ( .A(n637), .B(n357), .Y(n641) );
  AND2X2 U28 ( .A(n637), .B(addr[0]), .Y(n642) );
  MX4X1 U29 ( .A(memory[176]), .B(memory[160]), .C(memory[144]), .D(
        memory[128]), .S0(n352), .S1(n349), .Y(n19) );
  MX4X1 U30 ( .A(memory[177]), .B(memory[161]), .C(memory[145]), .D(
        memory[129]), .S0(n351), .S1(n349), .Y(n27) );
  MX4X1 U31 ( .A(memory[178]), .B(memory[162]), .C(memory[146]), .D(
        memory[130]), .S0(n351), .S1(n349), .Y(n34) );
  MX4X1 U32 ( .A(memory[179]), .B(memory[163]), .C(memory[147]), .D(
        memory[131]), .S0(n351), .S1(n349), .Y(n41) );
  MX4X1 U33 ( .A(memory[180]), .B(memory[164]), .C(memory[148]), .D(
        memory[132]), .S0(n352), .S1(addr[1]), .Y(n46) );
  MX4X1 U34 ( .A(memory[181]), .B(memory[165]), .C(memory[149]), .D(
        memory[133]), .S0(n352), .S1(addr[1]), .Y(n307) );
  MX4X1 U35 ( .A(memory[182]), .B(memory[166]), .C(memory[150]), .D(
        memory[134]), .S0(n352), .S1(addr[1]), .Y(n311) );
  MX4X1 U36 ( .A(memory[183]), .B(memory[167]), .C(memory[151]), .D(
        memory[135]), .S0(n353), .S1(addr[1]), .Y(n315) );
  MX4X1 U37 ( .A(memory[184]), .B(memory[168]), .C(memory[152]), .D(
        memory[136]), .S0(n353), .S1(n349), .Y(n319) );
  MX4X1 U38 ( .A(memory[185]), .B(memory[169]), .C(memory[153]), .D(
        memory[137]), .S0(n353), .S1(n350), .Y(n323) );
  MX4X1 U39 ( .A(memory[186]), .B(memory[170]), .C(memory[154]), .D(
        memory[138]), .S0(addr[0]), .S1(n350), .Y(n327) );
  MX4X1 U40 ( .A(memory[187]), .B(memory[171]), .C(memory[155]), .D(
        memory[139]), .S0(n353), .S1(n350), .Y(n331) );
  MX4X1 U41 ( .A(memory[188]), .B(memory[172]), .C(memory[156]), .D(
        memory[140]), .S0(n351), .S1(n350), .Y(n335) );
  MX4X1 U42 ( .A(memory[189]), .B(memory[173]), .C(memory[157]), .D(
        memory[141]), .S0(n352), .S1(addr[1]), .Y(n339) );
  MX4X1 U43 ( .A(memory[190]), .B(memory[174]), .C(memory[158]), .D(
        memory[142]), .S0(addr[0]), .S1(addr[1]), .Y(n343) );
  MX4X1 U44 ( .A(memory[191]), .B(memory[175]), .C(memory[159]), .D(
        memory[143]), .S0(addr[0]), .S1(n350), .Y(n347) );
  MX4X1 U45 ( .A(memory[48]), .B(memory[32]), .C(memory[16]), .D(memory[0]), 
        .S0(n351), .S1(n349), .Y(n17) );
  MX4X1 U46 ( .A(memory[49]), .B(memory[33]), .C(memory[17]), .D(memory[1]), 
        .S0(n351), .S1(n349), .Y(n23) );
  MX4X1 U47 ( .A(memory[50]), .B(memory[34]), .C(memory[18]), .D(memory[2]), 
        .S0(n351), .S1(n349), .Y(n30) );
  MX4X1 U48 ( .A(memory[51]), .B(memory[35]), .C(memory[19]), .D(memory[3]), 
        .S0(n351), .S1(n349), .Y(n38) );
  MX4X1 U49 ( .A(memory[52]), .B(memory[36]), .C(memory[20]), .D(memory[4]), 
        .S0(n352), .S1(n349), .Y(n43) );
  MX4X1 U50 ( .A(memory[53]), .B(memory[37]), .C(memory[21]), .D(memory[5]), 
        .S0(n352), .S1(n350), .Y(n305) );
  MX4X1 U51 ( .A(memory[54]), .B(memory[38]), .C(memory[22]), .D(memory[6]), 
        .S0(n352), .S1(addr[1]), .Y(n309) );
  MX4X1 U52 ( .A(memory[55]), .B(memory[39]), .C(memory[23]), .D(memory[7]), 
        .S0(n353), .S1(n349), .Y(n313) );
  MX4X1 U53 ( .A(memory[56]), .B(memory[40]), .C(memory[24]), .D(memory[8]), 
        .S0(n353), .S1(n350), .Y(n317) );
  MX4X1 U54 ( .A(memory[57]), .B(memory[41]), .C(memory[25]), .D(memory[9]), 
        .S0(n353), .S1(n349), .Y(n321) );
  MX4X1 U55 ( .A(memory[58]), .B(memory[42]), .C(memory[26]), .D(memory[10]), 
        .S0(n353), .S1(n350), .Y(n325) );
  MX4X1 U56 ( .A(memory[59]), .B(memory[43]), .C(memory[27]), .D(memory[11]), 
        .S0(n351), .S1(n350), .Y(n329) );
  MX4X1 U57 ( .A(memory[60]), .B(memory[44]), .C(memory[28]), .D(memory[12]), 
        .S0(n352), .S1(n350), .Y(n333) );
  MX4X1 U58 ( .A(memory[61]), .B(memory[45]), .C(memory[29]), .D(memory[13]), 
        .S0(n353), .S1(n349), .Y(n337) );
  MX4X1 U59 ( .A(memory[62]), .B(memory[46]), .C(memory[30]), .D(memory[14]), 
        .S0(n351), .S1(n350), .Y(n341) );
  MX4X1 U60 ( .A(memory[63]), .B(memory[47]), .C(memory[31]), .D(memory[15]), 
        .S0(addr[0]), .S1(n350), .Y(n345) );
  NOR2BX1 U61 ( .AN(N50), .B(n356), .Y(dout[0]) );
  MX4X1 U62 ( .A(n20), .B(n18), .C(n19), .D(n17), .S0(n355), .S1(n354), .Y(N50) );
  MX4X1 U63 ( .A(memory[240]), .B(memory[224]), .C(memory[208]), .D(
        memory[192]), .S0(n352), .S1(addr[1]), .Y(n20) );
  MX4X1 U64 ( .A(memory[112]), .B(memory[96]), .C(memory[80]), .D(memory[64]), 
        .S0(n353), .S1(n350), .Y(n18) );
  NOR2BX1 U65 ( .AN(N49), .B(n356), .Y(dout[1]) );
  MX4X1 U66 ( .A(n28), .B(n25), .C(n27), .D(n23), .S0(n355), .S1(n354), .Y(N49) );
  MX4X1 U67 ( .A(memory[241]), .B(memory[225]), .C(memory[209]), .D(
        memory[193]), .S0(n351), .S1(n349), .Y(n28) );
  MX4X1 U68 ( .A(memory[113]), .B(memory[97]), .C(memory[81]), .D(memory[65]), 
        .S0(n351), .S1(n349), .Y(n25) );
  NOR2BX1 U69 ( .AN(N48), .B(n356), .Y(dout[2]) );
  MX4X1 U70 ( .A(n36), .B(n31), .C(n34), .D(n30), .S0(n355), .S1(n354), .Y(N48) );
  MX4X1 U71 ( .A(memory[242]), .B(memory[226]), .C(memory[210]), .D(
        memory[194]), .S0(n351), .S1(n349), .Y(n36) );
  MX4X1 U72 ( .A(memory[114]), .B(memory[98]), .C(memory[82]), .D(memory[66]), 
        .S0(n351), .S1(n349), .Y(n31) );
  NOR2BX1 U73 ( .AN(N47), .B(n356), .Y(dout[3]) );
  MX4X1 U74 ( .A(n42), .B(n40), .C(n41), .D(n38), .S0(n355), .S1(n354), .Y(N47) );
  MX4X1 U75 ( .A(memory[243]), .B(memory[227]), .C(memory[211]), .D(
        memory[195]), .S0(n351), .S1(n349), .Y(n42) );
  MX4X1 U76 ( .A(memory[115]), .B(memory[99]), .C(memory[83]), .D(memory[67]), 
        .S0(n351), .S1(n349), .Y(n40) );
  NOR2BX1 U77 ( .AN(N46), .B(n356), .Y(dout[4]) );
  MX4X1 U78 ( .A(n304), .B(n44), .C(n46), .D(n43), .S0(n355), .S1(n354), .Y(
        N46) );
  MX4X1 U79 ( .A(memory[244]), .B(memory[228]), .C(memory[212]), .D(
        memory[196]), .S0(n352), .S1(addr[1]), .Y(n304) );
  MX4X1 U80 ( .A(memory[116]), .B(memory[100]), .C(memory[84]), .D(memory[68]), 
        .S0(n352), .S1(addr[1]), .Y(n44) );
  NOR2BX1 U81 ( .AN(N45), .B(n356), .Y(dout[5]) );
  MX4X1 U82 ( .A(n308), .B(n306), .C(n307), .D(n305), .S0(n355), .S1(n354), 
        .Y(N45) );
  MX4X1 U83 ( .A(memory[245]), .B(memory[229]), .C(memory[213]), .D(
        memory[197]), .S0(n352), .S1(addr[1]), .Y(n308) );
  MX4X1 U84 ( .A(memory[117]), .B(memory[101]), .C(memory[85]), .D(memory[69]), 
        .S0(n352), .S1(addr[1]), .Y(n306) );
  NOR2BX1 U85 ( .AN(N44), .B(n356), .Y(dout[6]) );
  MX4X1 U86 ( .A(n312), .B(n310), .C(n311), .D(n309), .S0(n355), .S1(n354), 
        .Y(N44) );
  MX4X1 U87 ( .A(memory[246]), .B(memory[230]), .C(memory[214]), .D(
        memory[198]), .S0(n352), .S1(addr[1]), .Y(n312) );
  MX4X1 U88 ( .A(memory[118]), .B(memory[102]), .C(memory[86]), .D(memory[70]), 
        .S0(n352), .S1(addr[1]), .Y(n310) );
  NOR2BX1 U89 ( .AN(N43), .B(n356), .Y(dout[7]) );
  MX4X1 U90 ( .A(n316), .B(n314), .C(n315), .D(n313), .S0(n355), .S1(n354), 
        .Y(N43) );
  MX4X1 U91 ( .A(memory[247]), .B(memory[231]), .C(memory[215]), .D(
        memory[199]), .S0(n353), .S1(addr[1]), .Y(n316) );
  MX4X1 U92 ( .A(memory[119]), .B(memory[103]), .C(memory[87]), .D(memory[71]), 
        .S0(n353), .S1(n349), .Y(n314) );
  NOR2BX1 U93 ( .AN(N42), .B(n356), .Y(dout[8]) );
  MX4X1 U94 ( .A(n320), .B(n318), .C(n319), .D(n317), .S0(n355), .S1(n354), 
        .Y(N42) );
  MX4X1 U95 ( .A(memory[248]), .B(memory[232]), .C(memory[216]), .D(
        memory[200]), .S0(n353), .S1(addr[1]), .Y(n320) );
  MX4X1 U96 ( .A(memory[120]), .B(memory[104]), .C(memory[88]), .D(memory[72]), 
        .S0(n353), .S1(addr[1]), .Y(n318) );
  NOR2BX1 U97 ( .AN(N41), .B(n356), .Y(dout[9]) );
  MX4X1 U98 ( .A(n324), .B(n322), .C(n323), .D(n321), .S0(n355), .S1(n354), 
        .Y(N41) );
  MX4X1 U99 ( .A(memory[249]), .B(memory[233]), .C(memory[217]), .D(
        memory[201]), .S0(n353), .S1(addr[1]), .Y(n324) );
  MX4X1 U100 ( .A(memory[121]), .B(memory[105]), .C(memory[89]), .D(memory[73]), .S0(n353), .S1(addr[1]), .Y(n322) );
  NOR2BX1 U101 ( .AN(N40), .B(n356), .Y(dout[10]) );
  MX4X1 U102 ( .A(n328), .B(n326), .C(n327), .D(n325), .S0(n355), .S1(n354), 
        .Y(N40) );
  MX4X1 U103 ( .A(memory[250]), .B(memory[234]), .C(memory[218]), .D(
        memory[202]), .S0(n353), .S1(n350), .Y(n328) );
  MX4X1 U104 ( .A(memory[122]), .B(memory[106]), .C(memory[90]), .D(memory[74]), .S0(n352), .S1(n350), .Y(n326) );
  NOR2BX1 U105 ( .AN(N39), .B(n356), .Y(dout[11]) );
  MX4X1 U106 ( .A(n332), .B(n330), .C(n331), .D(n329), .S0(n355), .S1(n354), 
        .Y(N39) );
  MX4X1 U107 ( .A(memory[251]), .B(memory[235]), .C(memory[219]), .D(
        memory[203]), .S0(n351), .S1(n350), .Y(n332) );
  MX4X1 U108 ( .A(memory[123]), .B(memory[107]), .C(memory[91]), .D(memory[75]), .S0(n353), .S1(n350), .Y(n330) );
  NOR2BX1 U109 ( .AN(N38), .B(n356), .Y(dout[12]) );
  MX4X1 U110 ( .A(n336), .B(n334), .C(n335), .D(n333), .S0(n355), .S1(n354), 
        .Y(N38) );
  MX4X1 U111 ( .A(memory[252]), .B(memory[236]), .C(memory[220]), .D(
        memory[204]), .S0(n352), .S1(n350), .Y(n336) );
  MX4X1 U112 ( .A(memory[124]), .B(memory[108]), .C(memory[92]), .D(memory[76]), .S0(n351), .S1(n350), .Y(n334) );
  NOR2BX1 U113 ( .AN(N37), .B(n356), .Y(dout[13]) );
  MX4X1 U114 ( .A(n340), .B(n338), .C(n339), .D(n337), .S0(n355), .S1(n354), 
        .Y(N37) );
  MX4X1 U115 ( .A(memory[253]), .B(memory[237]), .C(memory[221]), .D(
        memory[205]), .S0(addr[0]), .S1(n349), .Y(n340) );
  MX4X1 U116 ( .A(memory[125]), .B(memory[109]), .C(memory[93]), .D(memory[77]), .S0(addr[0]), .S1(n349), .Y(n338) );
  NOR2BX1 U117 ( .AN(N36), .B(n356), .Y(dout[14]) );
  MX4X1 U118 ( .A(n344), .B(n342), .C(n343), .D(n341), .S0(n355), .S1(n354), 
        .Y(N36) );
  MX4X1 U119 ( .A(memory[254]), .B(memory[238]), .C(memory[222]), .D(
        memory[206]), .S0(addr[0]), .S1(n350), .Y(n344) );
  MX4X1 U120 ( .A(memory[126]), .B(memory[110]), .C(memory[94]), .D(memory[78]), .S0(addr[0]), .S1(n350), .Y(n342) );
  NOR2BX1 U121 ( .AN(N35), .B(n356), .Y(dout[15]) );
  MX4X1 U122 ( .A(n348), .B(n346), .C(n347), .D(n345), .S0(n355), .S1(n354), 
        .Y(N35) );
  MX4X1 U123 ( .A(memory[255]), .B(memory[239]), .C(memory[223]), .D(
        memory[207]), .S0(addr[0]), .S1(n349), .Y(n348) );
  MX4X1 U124 ( .A(memory[127]), .B(memory[111]), .C(memory[95]), .D(memory[79]), .S0(addr[0]), .S1(n350), .Y(n346) );
  INVX1 U125 ( .A(addr[1]), .Y(n358) );
  INVX1 U126 ( .A(addr[0]), .Y(n357) );
  NOR2X1 U127 ( .A(n358), .B(addr[2]), .Y(n639) );
  NOR2X1 U128 ( .A(addr[1]), .B(addr[2]), .Y(n638) );
  BUFX3 U129 ( .A(addr[3]), .Y(n355) );
  OAI2BB2X1 U130 ( .B0(n1), .B1(n375), .A0N(memory[0]), .A1N(n1), .Y(n631) );
  OAI2BB2X1 U131 ( .B0(n1), .B1(n374), .A0N(memory[1]), .A1N(n1), .Y(n630) );
  OAI2BB2X1 U132 ( .B0(n1), .B1(n373), .A0N(memory[2]), .A1N(n1), .Y(n629) );
  OAI2BB2X1 U133 ( .B0(n1), .B1(n372), .A0N(memory[3]), .A1N(n1), .Y(n628) );
  OAI2BB2X1 U134 ( .B0(n1), .B1(n371), .A0N(memory[4]), .A1N(n1), .Y(n627) );
  OAI2BB2X1 U135 ( .B0(n1), .B1(n370), .A0N(memory[5]), .A1N(n1), .Y(n626) );
  OAI2BB2X1 U136 ( .B0(n1), .B1(n369), .A0N(memory[6]), .A1N(n1), .Y(n625) );
  OAI2BB2X1 U137 ( .B0(n1), .B1(n368), .A0N(memory[7]), .A1N(n1), .Y(n624) );
  OAI2BB2X1 U138 ( .B0(n1), .B1(n367), .A0N(memory[8]), .A1N(n1), .Y(n623) );
  OAI2BB2X1 U139 ( .B0(n1), .B1(n366), .A0N(memory[9]), .A1N(n1), .Y(n622) );
  OAI2BB2X1 U140 ( .B0(n1), .B1(n365), .A0N(memory[10]), .A1N(n1), .Y(n621) );
  OAI2BB2X1 U141 ( .B0(n1), .B1(n364), .A0N(memory[11]), .A1N(n1), .Y(n620) );
  OAI2BB2X1 U142 ( .B0(n1), .B1(n363), .A0N(memory[12]), .A1N(n1), .Y(n619) );
  OAI2BB2X1 U143 ( .B0(n1), .B1(n362), .A0N(memory[13]), .A1N(n1), .Y(n618) );
  OAI2BB2X1 U144 ( .B0(n1), .B1(n361), .A0N(memory[14]), .A1N(n1), .Y(n617) );
  OAI2BB2X1 U145 ( .B0(n1), .B1(n360), .A0N(memory[15]), .A1N(n1), .Y(n616) );
  OAI2BB2X1 U146 ( .B0(n375), .B1(n2), .A0N(memory[16]), .A1N(n2), .Y(n615) );
  OAI2BB2X1 U147 ( .B0(n374), .B1(n2), .A0N(memory[17]), .A1N(n2), .Y(n614) );
  OAI2BB2X1 U148 ( .B0(n373), .B1(n2), .A0N(memory[18]), .A1N(n2), .Y(n613) );
  OAI2BB2X1 U149 ( .B0(n372), .B1(n2), .A0N(memory[19]), .A1N(n2), .Y(n612) );
  OAI2BB2X1 U150 ( .B0(n371), .B1(n2), .A0N(memory[20]), .A1N(n2), .Y(n611) );
  OAI2BB2X1 U151 ( .B0(n370), .B1(n2), .A0N(memory[21]), .A1N(n2), .Y(n610) );
  OAI2BB2X1 U152 ( .B0(n369), .B1(n2), .A0N(memory[22]), .A1N(n2), .Y(n609) );
  OAI2BB2X1 U153 ( .B0(n368), .B1(n2), .A0N(memory[23]), .A1N(n2), .Y(n608) );
  OAI2BB2X1 U154 ( .B0(n363), .B1(n2), .A0N(memory[28]), .A1N(n2), .Y(n603) );
  OAI2BB2X1 U155 ( .B0(n362), .B1(n2), .A0N(memory[29]), .A1N(n2), .Y(n602) );
  OAI2BB2X1 U156 ( .B0(n361), .B1(n2), .A0N(memory[30]), .A1N(n2), .Y(n601) );
  OAI2BB2X1 U157 ( .B0(n360), .B1(n2), .A0N(memory[31]), .A1N(n2), .Y(n600) );
  OAI2BB2X1 U158 ( .B0(n375), .B1(n3), .A0N(memory[32]), .A1N(n3), .Y(n599) );
  OAI2BB2X1 U159 ( .B0(n374), .B1(n3), .A0N(memory[33]), .A1N(n3), .Y(n598) );
  OAI2BB2X1 U160 ( .B0(n373), .B1(n3), .A0N(memory[34]), .A1N(n3), .Y(n597) );
  OAI2BB2X1 U161 ( .B0(n372), .B1(n3), .A0N(memory[35]), .A1N(n3), .Y(n596) );
  OAI2BB2X1 U162 ( .B0(n371), .B1(n3), .A0N(memory[36]), .A1N(n3), .Y(n595) );
  OAI2BB2X1 U163 ( .B0(n370), .B1(n3), .A0N(memory[37]), .A1N(n3), .Y(n594) );
  OAI2BB2X1 U164 ( .B0(n369), .B1(n3), .A0N(memory[38]), .A1N(n3), .Y(n593) );
  OAI2BB2X1 U165 ( .B0(n368), .B1(n3), .A0N(memory[39]), .A1N(n3), .Y(n592) );
  OAI2BB2X1 U166 ( .B0(n363), .B1(n3), .A0N(memory[44]), .A1N(n3), .Y(n587) );
  OAI2BB2X1 U167 ( .B0(n362), .B1(n3), .A0N(memory[45]), .A1N(n3), .Y(n586) );
  OAI2BB2X1 U168 ( .B0(n361), .B1(n3), .A0N(memory[46]), .A1N(n3), .Y(n585) );
  OAI2BB2X1 U169 ( .B0(n360), .B1(n3), .A0N(memory[47]), .A1N(n3), .Y(n584) );
  OAI2BB2X1 U170 ( .B0(n375), .B1(n4), .A0N(memory[48]), .A1N(n4), .Y(n583) );
  OAI2BB2X1 U171 ( .B0(n374), .B1(n4), .A0N(memory[49]), .A1N(n4), .Y(n582) );
  OAI2BB2X1 U172 ( .B0(n373), .B1(n4), .A0N(memory[50]), .A1N(n4), .Y(n581) );
  OAI2BB2X1 U173 ( .B0(n372), .B1(n4), .A0N(memory[51]), .A1N(n4), .Y(n580) );
  OAI2BB2X1 U174 ( .B0(n371), .B1(n4), .A0N(memory[52]), .A1N(n4), .Y(n579) );
  OAI2BB2X1 U175 ( .B0(n370), .B1(n4), .A0N(memory[53]), .A1N(n4), .Y(n578) );
  OAI2BB2X1 U176 ( .B0(n369), .B1(n4), .A0N(memory[54]), .A1N(n4), .Y(n577) );
  OAI2BB2X1 U177 ( .B0(n368), .B1(n4), .A0N(memory[55]), .A1N(n4), .Y(n576) );
  OAI2BB2X1 U178 ( .B0(n363), .B1(n4), .A0N(memory[60]), .A1N(n4), .Y(n571) );
  OAI2BB2X1 U179 ( .B0(n362), .B1(n4), .A0N(memory[61]), .A1N(n4), .Y(n570) );
  OAI2BB2X1 U180 ( .B0(n361), .B1(n4), .A0N(memory[62]), .A1N(n4), .Y(n569) );
  OAI2BB2X1 U181 ( .B0(n360), .B1(n4), .A0N(memory[63]), .A1N(n4), .Y(n568) );
  OAI2BB2X1 U182 ( .B0(n375), .B1(n5), .A0N(memory[64]), .A1N(n5), .Y(n567) );
  OAI2BB2X1 U183 ( .B0(n374), .B1(n5), .A0N(memory[65]), .A1N(n5), .Y(n566) );
  OAI2BB2X1 U184 ( .B0(n373), .B1(n5), .A0N(memory[66]), .A1N(n5), .Y(n565) );
  OAI2BB2X1 U185 ( .B0(n372), .B1(n5), .A0N(memory[67]), .A1N(n5), .Y(n564) );
  OAI2BB2X1 U186 ( .B0(n371), .B1(n5), .A0N(memory[68]), .A1N(n5), .Y(n563) );
  OAI2BB2X1 U187 ( .B0(n370), .B1(n5), .A0N(memory[69]), .A1N(n5), .Y(n562) );
  OAI2BB2X1 U188 ( .B0(n369), .B1(n5), .A0N(memory[70]), .A1N(n5), .Y(n561) );
  OAI2BB2X1 U189 ( .B0(n368), .B1(n5), .A0N(memory[71]), .A1N(n5), .Y(n560) );
  OAI2BB2X1 U190 ( .B0(n363), .B1(n5), .A0N(memory[76]), .A1N(n5), .Y(n555) );
  OAI2BB2X1 U191 ( .B0(n362), .B1(n5), .A0N(memory[77]), .A1N(n5), .Y(n554) );
  OAI2BB2X1 U192 ( .B0(n361), .B1(n5), .A0N(memory[78]), .A1N(n5), .Y(n553) );
  OAI2BB2X1 U193 ( .B0(n360), .B1(n5), .A0N(memory[79]), .A1N(n5), .Y(n552) );
  OAI2BB2X1 U194 ( .B0(n375), .B1(n6), .A0N(memory[80]), .A1N(n6), .Y(n551) );
  OAI2BB2X1 U195 ( .B0(n374), .B1(n6), .A0N(memory[81]), .A1N(n6), .Y(n550) );
  OAI2BB2X1 U196 ( .B0(n373), .B1(n6), .A0N(memory[82]), .A1N(n6), .Y(n549) );
  OAI2BB2X1 U197 ( .B0(n372), .B1(n6), .A0N(memory[83]), .A1N(n6), .Y(n548) );
  OAI2BB2X1 U198 ( .B0(n371), .B1(n6), .A0N(memory[84]), .A1N(n6), .Y(n547) );
  OAI2BB2X1 U199 ( .B0(n370), .B1(n6), .A0N(memory[85]), .A1N(n6), .Y(n546) );
  OAI2BB2X1 U200 ( .B0(n369), .B1(n6), .A0N(memory[86]), .A1N(n6), .Y(n545) );
  OAI2BB2X1 U201 ( .B0(n368), .B1(n6), .A0N(memory[87]), .A1N(n6), .Y(n544) );
  OAI2BB2X1 U202 ( .B0(n363), .B1(n6), .A0N(memory[92]), .A1N(n6), .Y(n539) );
  OAI2BB2X1 U203 ( .B0(n362), .B1(n6), .A0N(memory[93]), .A1N(n6), .Y(n538) );
  OAI2BB2X1 U204 ( .B0(n361), .B1(n6), .A0N(memory[94]), .A1N(n6), .Y(n537) );
  OAI2BB2X1 U205 ( .B0(n360), .B1(n6), .A0N(memory[95]), .A1N(n6), .Y(n536) );
  OAI2BB2X1 U206 ( .B0(n375), .B1(n7), .A0N(memory[96]), .A1N(n7), .Y(n535) );
  OAI2BB2X1 U207 ( .B0(n374), .B1(n7), .A0N(memory[97]), .A1N(n7), .Y(n534) );
  OAI2BB2X1 U208 ( .B0(n373), .B1(n7), .A0N(memory[98]), .A1N(n7), .Y(n533) );
  OAI2BB2X1 U209 ( .B0(n372), .B1(n7), .A0N(memory[99]), .A1N(n7), .Y(n532) );
  OAI2BB2X1 U210 ( .B0(n371), .B1(n7), .A0N(memory[100]), .A1N(n7), .Y(n531)
         );
  OAI2BB2X1 U211 ( .B0(n370), .B1(n7), .A0N(memory[101]), .A1N(n7), .Y(n530)
         );
  OAI2BB2X1 U212 ( .B0(n369), .B1(n7), .A0N(memory[102]), .A1N(n7), .Y(n529)
         );
  OAI2BB2X1 U213 ( .B0(n368), .B1(n7), .A0N(memory[103]), .A1N(n7), .Y(n528)
         );
  OAI2BB2X1 U214 ( .B0(n363), .B1(n7), .A0N(memory[108]), .A1N(n7), .Y(n523)
         );
  OAI2BB2X1 U215 ( .B0(n362), .B1(n7), .A0N(memory[109]), .A1N(n7), .Y(n522)
         );
  OAI2BB2X1 U216 ( .B0(n361), .B1(n7), .A0N(memory[110]), .A1N(n7), .Y(n521)
         );
  OAI2BB2X1 U217 ( .B0(n360), .B1(n7), .A0N(memory[111]), .A1N(n7), .Y(n520)
         );
  OAI2BB2X1 U218 ( .B0(n375), .B1(n8), .A0N(memory[112]), .A1N(n8), .Y(n519)
         );
  OAI2BB2X1 U219 ( .B0(n374), .B1(n8), .A0N(memory[113]), .A1N(n8), .Y(n518)
         );
  OAI2BB2X1 U220 ( .B0(n373), .B1(n8), .A0N(memory[114]), .A1N(n8), .Y(n517)
         );
  OAI2BB2X1 U221 ( .B0(n372), .B1(n8), .A0N(memory[115]), .A1N(n8), .Y(n516)
         );
  OAI2BB2X1 U222 ( .B0(n371), .B1(n8), .A0N(memory[116]), .A1N(n8), .Y(n515)
         );
  OAI2BB2X1 U223 ( .B0(n370), .B1(n8), .A0N(memory[117]), .A1N(n8), .Y(n514)
         );
  OAI2BB2X1 U224 ( .B0(n369), .B1(n8), .A0N(memory[118]), .A1N(n8), .Y(n513)
         );
  OAI2BB2X1 U225 ( .B0(n368), .B1(n8), .A0N(memory[119]), .A1N(n8), .Y(n512)
         );
  OAI2BB2X1 U226 ( .B0(n363), .B1(n8), .A0N(memory[124]), .A1N(n8), .Y(n507)
         );
  OAI2BB2X1 U227 ( .B0(n362), .B1(n8), .A0N(memory[125]), .A1N(n8), .Y(n506)
         );
  OAI2BB2X1 U228 ( .B0(n361), .B1(n8), .A0N(memory[126]), .A1N(n8), .Y(n505)
         );
  OAI2BB2X1 U229 ( .B0(n360), .B1(n8), .A0N(memory[127]), .A1N(n8), .Y(n504)
         );
  OAI2BB2X1 U230 ( .B0(n375), .B1(n9), .A0N(memory[128]), .A1N(n9), .Y(n503)
         );
  OAI2BB2X1 U231 ( .B0(n374), .B1(n9), .A0N(memory[129]), .A1N(n9), .Y(n502)
         );
  OAI2BB2X1 U232 ( .B0(n373), .B1(n9), .A0N(memory[130]), .A1N(n9), .Y(n501)
         );
  OAI2BB2X1 U233 ( .B0(n372), .B1(n9), .A0N(memory[131]), .A1N(n9), .Y(n500)
         );
  OAI2BB2X1 U234 ( .B0(n371), .B1(n9), .A0N(memory[132]), .A1N(n9), .Y(n499)
         );
  OAI2BB2X1 U235 ( .B0(n370), .B1(n9), .A0N(memory[133]), .A1N(n9), .Y(n498)
         );
  OAI2BB2X1 U236 ( .B0(n369), .B1(n9), .A0N(memory[134]), .A1N(n9), .Y(n497)
         );
  OAI2BB2X1 U237 ( .B0(n368), .B1(n9), .A0N(memory[135]), .A1N(n9), .Y(n496)
         );
  OAI2BB2X1 U238 ( .B0(n363), .B1(n9), .A0N(memory[140]), .A1N(n9), .Y(n491)
         );
  OAI2BB2X1 U239 ( .B0(n362), .B1(n9), .A0N(memory[141]), .A1N(n9), .Y(n490)
         );
  OAI2BB2X1 U240 ( .B0(n361), .B1(n9), .A0N(memory[142]), .A1N(n9), .Y(n489)
         );
  OAI2BB2X1 U241 ( .B0(n360), .B1(n9), .A0N(memory[143]), .A1N(n9), .Y(n488)
         );
  OAI2BB2X1 U242 ( .B0(n375), .B1(n10), .A0N(memory[144]), .A1N(n10), .Y(n487)
         );
  OAI2BB2X1 U243 ( .B0(n374), .B1(n10), .A0N(memory[145]), .A1N(n10), .Y(n486)
         );
  OAI2BB2X1 U244 ( .B0(n373), .B1(n10), .A0N(memory[146]), .A1N(n10), .Y(n485)
         );
  OAI2BB2X1 U245 ( .B0(n372), .B1(n10), .A0N(memory[147]), .A1N(n10), .Y(n484)
         );
  OAI2BB2X1 U246 ( .B0(n371), .B1(n10), .A0N(memory[148]), .A1N(n10), .Y(n483)
         );
  OAI2BB2X1 U247 ( .B0(n370), .B1(n10), .A0N(memory[149]), .A1N(n10), .Y(n482)
         );
  OAI2BB2X1 U248 ( .B0(n369), .B1(n10), .A0N(memory[150]), .A1N(n10), .Y(n481)
         );
  OAI2BB2X1 U249 ( .B0(n368), .B1(n10), .A0N(memory[151]), .A1N(n10), .Y(n480)
         );
  OAI2BB2X1 U250 ( .B0(n363), .B1(n10), .A0N(memory[156]), .A1N(n10), .Y(n475)
         );
  OAI2BB2X1 U251 ( .B0(n362), .B1(n10), .A0N(memory[157]), .A1N(n10), .Y(n474)
         );
  OAI2BB2X1 U252 ( .B0(n361), .B1(n10), .A0N(memory[158]), .A1N(n10), .Y(n473)
         );
  OAI2BB2X1 U253 ( .B0(n360), .B1(n10), .A0N(memory[159]), .A1N(n10), .Y(n472)
         );
  OAI2BB2X1 U254 ( .B0(n375), .B1(n11), .A0N(memory[160]), .A1N(n11), .Y(n471)
         );
  OAI2BB2X1 U255 ( .B0(n374), .B1(n11), .A0N(memory[161]), .A1N(n11), .Y(n470)
         );
  OAI2BB2X1 U256 ( .B0(n373), .B1(n11), .A0N(memory[162]), .A1N(n11), .Y(n469)
         );
  OAI2BB2X1 U257 ( .B0(n372), .B1(n11), .A0N(memory[163]), .A1N(n11), .Y(n468)
         );
  OAI2BB2X1 U258 ( .B0(n371), .B1(n11), .A0N(memory[164]), .A1N(n11), .Y(n467)
         );
  OAI2BB2X1 U259 ( .B0(n370), .B1(n11), .A0N(memory[165]), .A1N(n11), .Y(n466)
         );
  OAI2BB2X1 U260 ( .B0(n369), .B1(n11), .A0N(memory[166]), .A1N(n11), .Y(n465)
         );
  OAI2BB2X1 U261 ( .B0(n368), .B1(n11), .A0N(memory[167]), .A1N(n11), .Y(n464)
         );
  OAI2BB2X1 U262 ( .B0(n363), .B1(n11), .A0N(memory[172]), .A1N(n11), .Y(n459)
         );
  OAI2BB2X1 U263 ( .B0(n362), .B1(n11), .A0N(memory[173]), .A1N(n11), .Y(n458)
         );
  OAI2BB2X1 U264 ( .B0(n361), .B1(n11), .A0N(memory[174]), .A1N(n11), .Y(n457)
         );
  OAI2BB2X1 U265 ( .B0(n360), .B1(n11), .A0N(memory[175]), .A1N(n11), .Y(n456)
         );
  OAI2BB2X1 U266 ( .B0(n375), .B1(n12), .A0N(memory[176]), .A1N(n12), .Y(n455)
         );
  OAI2BB2X1 U267 ( .B0(n374), .B1(n12), .A0N(memory[177]), .A1N(n12), .Y(n454)
         );
  OAI2BB2X1 U268 ( .B0(n373), .B1(n12), .A0N(memory[178]), .A1N(n12), .Y(n453)
         );
  OAI2BB2X1 U269 ( .B0(n372), .B1(n12), .A0N(memory[179]), .A1N(n12), .Y(n452)
         );
  OAI2BB2X1 U270 ( .B0(n371), .B1(n12), .A0N(memory[180]), .A1N(n12), .Y(n451)
         );
  OAI2BB2X1 U271 ( .B0(n370), .B1(n12), .A0N(memory[181]), .A1N(n12), .Y(n450)
         );
  OAI2BB2X1 U272 ( .B0(n369), .B1(n12), .A0N(memory[182]), .A1N(n12), .Y(n449)
         );
  OAI2BB2X1 U273 ( .B0(n368), .B1(n12), .A0N(memory[183]), .A1N(n12), .Y(n448)
         );
  OAI2BB2X1 U274 ( .B0(n363), .B1(n12), .A0N(memory[188]), .A1N(n12), .Y(n443)
         );
  OAI2BB2X1 U275 ( .B0(n362), .B1(n12), .A0N(memory[189]), .A1N(n12), .Y(n442)
         );
  OAI2BB2X1 U276 ( .B0(n361), .B1(n12), .A0N(memory[190]), .A1N(n12), .Y(n441)
         );
  OAI2BB2X1 U277 ( .B0(n360), .B1(n12), .A0N(memory[191]), .A1N(n12), .Y(n440)
         );
  OAI2BB2X1 U278 ( .B0(n375), .B1(n13), .A0N(memory[192]), .A1N(n13), .Y(n439)
         );
  OAI2BB2X1 U279 ( .B0(n374), .B1(n13), .A0N(memory[193]), .A1N(n13), .Y(n438)
         );
  OAI2BB2X1 U280 ( .B0(n373), .B1(n13), .A0N(memory[194]), .A1N(n13), .Y(n437)
         );
  OAI2BB2X1 U281 ( .B0(n372), .B1(n13), .A0N(memory[195]), .A1N(n13), .Y(n436)
         );
  OAI2BB2X1 U282 ( .B0(n371), .B1(n13), .A0N(memory[196]), .A1N(n13), .Y(n435)
         );
  OAI2BB2X1 U283 ( .B0(n370), .B1(n13), .A0N(memory[197]), .A1N(n13), .Y(n434)
         );
  OAI2BB2X1 U284 ( .B0(n369), .B1(n13), .A0N(memory[198]), .A1N(n13), .Y(n433)
         );
  OAI2BB2X1 U285 ( .B0(n368), .B1(n13), .A0N(memory[199]), .A1N(n13), .Y(n432)
         );
  OAI2BB2X1 U286 ( .B0(n363), .B1(n13), .A0N(memory[204]), .A1N(n13), .Y(n427)
         );
  OAI2BB2X1 U287 ( .B0(n362), .B1(n13), .A0N(memory[205]), .A1N(n13), .Y(n426)
         );
  OAI2BB2X1 U288 ( .B0(n361), .B1(n13), .A0N(memory[206]), .A1N(n13), .Y(n425)
         );
  OAI2BB2X1 U289 ( .B0(n360), .B1(n13), .A0N(memory[207]), .A1N(n13), .Y(n424)
         );
  OAI2BB2X1 U290 ( .B0(n375), .B1(n14), .A0N(memory[208]), .A1N(n14), .Y(n423)
         );
  OAI2BB2X1 U291 ( .B0(n374), .B1(n14), .A0N(memory[209]), .A1N(n14), .Y(n422)
         );
  OAI2BB2X1 U292 ( .B0(n373), .B1(n14), .A0N(memory[210]), .A1N(n14), .Y(n421)
         );
  OAI2BB2X1 U293 ( .B0(n372), .B1(n14), .A0N(memory[211]), .A1N(n14), .Y(n420)
         );
  OAI2BB2X1 U294 ( .B0(n371), .B1(n14), .A0N(memory[212]), .A1N(n14), .Y(n419)
         );
  OAI2BB2X1 U295 ( .B0(n370), .B1(n14), .A0N(memory[213]), .A1N(n14), .Y(n418)
         );
  OAI2BB2X1 U296 ( .B0(n369), .B1(n14), .A0N(memory[214]), .A1N(n14), .Y(n417)
         );
  OAI2BB2X1 U297 ( .B0(n368), .B1(n14), .A0N(memory[215]), .A1N(n14), .Y(n416)
         );
  OAI2BB2X1 U298 ( .B0(n363), .B1(n14), .A0N(memory[220]), .A1N(n14), .Y(n411)
         );
  OAI2BB2X1 U299 ( .B0(n362), .B1(n14), .A0N(memory[221]), .A1N(n14), .Y(n410)
         );
  OAI2BB2X1 U300 ( .B0(n361), .B1(n14), .A0N(memory[222]), .A1N(n14), .Y(n409)
         );
  OAI2BB2X1 U301 ( .B0(n360), .B1(n14), .A0N(memory[223]), .A1N(n14), .Y(n408)
         );
  OAI2BB2X1 U302 ( .B0(n375), .B1(n15), .A0N(memory[224]), .A1N(n15), .Y(n407)
         );
  OAI2BB2X1 U303 ( .B0(n374), .B1(n15), .A0N(memory[225]), .A1N(n15), .Y(n406)
         );
  OAI2BB2X1 U304 ( .B0(n373), .B1(n15), .A0N(memory[226]), .A1N(n15), .Y(n405)
         );
  OAI2BB2X1 U305 ( .B0(n372), .B1(n15), .A0N(memory[227]), .A1N(n15), .Y(n404)
         );
  OAI2BB2X1 U306 ( .B0(n371), .B1(n15), .A0N(memory[228]), .A1N(n15), .Y(n403)
         );
  OAI2BB2X1 U307 ( .B0(n370), .B1(n15), .A0N(memory[229]), .A1N(n15), .Y(n402)
         );
  OAI2BB2X1 U308 ( .B0(n369), .B1(n15), .A0N(memory[230]), .A1N(n15), .Y(n401)
         );
  OAI2BB2X1 U309 ( .B0(n368), .B1(n15), .A0N(memory[231]), .A1N(n15), .Y(n400)
         );
  OAI2BB2X1 U310 ( .B0(n363), .B1(n15), .A0N(memory[236]), .A1N(n15), .Y(n395)
         );
  OAI2BB2X1 U311 ( .B0(n362), .B1(n15), .A0N(memory[237]), .A1N(n15), .Y(n394)
         );
  OAI2BB2X1 U312 ( .B0(n361), .B1(n15), .A0N(memory[238]), .A1N(n15), .Y(n393)
         );
  OAI2BB2X1 U313 ( .B0(n360), .B1(n15), .A0N(memory[239]), .A1N(n15), .Y(n392)
         );
  OAI2BB2X1 U314 ( .B0(n375), .B1(n16), .A0N(memory[240]), .A1N(n16), .Y(n391)
         );
  OAI2BB2X1 U315 ( .B0(n374), .B1(n16), .A0N(memory[241]), .A1N(n16), .Y(n390)
         );
  OAI2BB2X1 U316 ( .B0(n373), .B1(n16), .A0N(memory[242]), .A1N(n16), .Y(n389)
         );
  OAI2BB2X1 U317 ( .B0(n372), .B1(n16), .A0N(memory[243]), .A1N(n16), .Y(n388)
         );
  OAI2BB2X1 U318 ( .B0(n371), .B1(n16), .A0N(memory[244]), .A1N(n16), .Y(n387)
         );
  OAI2BB2X1 U319 ( .B0(n370), .B1(n16), .A0N(memory[245]), .A1N(n16), .Y(n386)
         );
  OAI2BB2X1 U320 ( .B0(n369), .B1(n16), .A0N(memory[246]), .A1N(n16), .Y(n385)
         );
  OAI2BB2X1 U321 ( .B0(n368), .B1(n16), .A0N(memory[247]), .A1N(n16), .Y(n384)
         );
  OAI2BB2X1 U322 ( .B0(n363), .B1(n16), .A0N(memory[252]), .A1N(n16), .Y(n379)
         );
  OAI2BB2X1 U323 ( .B0(n362), .B1(n16), .A0N(memory[253]), .A1N(n16), .Y(n378)
         );
  OAI2BB2X1 U324 ( .B0(n361), .B1(n16), .A0N(memory[254]), .A1N(n16), .Y(n377)
         );
  OAI2BB2X1 U325 ( .B0(n360), .B1(n16), .A0N(memory[255]), .A1N(n16), .Y(n376)
         );
  OAI2BB2X1 U326 ( .B0(n367), .B1(n2), .A0N(memory[24]), .A1N(n2), .Y(n607) );
  OAI2BB2X1 U327 ( .B0(n366), .B1(n2), .A0N(memory[25]), .A1N(n2), .Y(n606) );
  OAI2BB2X1 U328 ( .B0(n365), .B1(n2), .A0N(memory[26]), .A1N(n2), .Y(n605) );
  OAI2BB2X1 U329 ( .B0(n364), .B1(n2), .A0N(memory[27]), .A1N(n2), .Y(n604) );
  OAI2BB2X1 U330 ( .B0(n367), .B1(n3), .A0N(memory[40]), .A1N(n3), .Y(n591) );
  OAI2BB2X1 U331 ( .B0(n366), .B1(n3), .A0N(memory[41]), .A1N(n3), .Y(n590) );
  OAI2BB2X1 U332 ( .B0(n365), .B1(n3), .A0N(memory[42]), .A1N(n3), .Y(n589) );
  OAI2BB2X1 U333 ( .B0(n364), .B1(n3), .A0N(memory[43]), .A1N(n3), .Y(n588) );
  OAI2BB2X1 U334 ( .B0(n367), .B1(n4), .A0N(memory[56]), .A1N(n4), .Y(n575) );
  OAI2BB2X1 U335 ( .B0(n366), .B1(n4), .A0N(memory[57]), .A1N(n4), .Y(n574) );
  OAI2BB2X1 U336 ( .B0(n365), .B1(n4), .A0N(memory[58]), .A1N(n4), .Y(n573) );
  OAI2BB2X1 U337 ( .B0(n364), .B1(n4), .A0N(memory[59]), .A1N(n4), .Y(n572) );
  OAI2BB2X1 U338 ( .B0(n367), .B1(n5), .A0N(memory[72]), .A1N(n5), .Y(n559) );
  OAI2BB2X1 U339 ( .B0(n366), .B1(n5), .A0N(memory[73]), .A1N(n5), .Y(n558) );
  OAI2BB2X1 U340 ( .B0(n365), .B1(n5), .A0N(memory[74]), .A1N(n5), .Y(n557) );
  OAI2BB2X1 U341 ( .B0(n364), .B1(n5), .A0N(memory[75]), .A1N(n5), .Y(n556) );
  OAI2BB2X1 U342 ( .B0(n367), .B1(n6), .A0N(memory[88]), .A1N(n6), .Y(n543) );
  OAI2BB2X1 U343 ( .B0(n366), .B1(n6), .A0N(memory[89]), .A1N(n6), .Y(n542) );
  OAI2BB2X1 U344 ( .B0(n365), .B1(n6), .A0N(memory[90]), .A1N(n6), .Y(n541) );
  OAI2BB2X1 U345 ( .B0(n364), .B1(n6), .A0N(memory[91]), .A1N(n6), .Y(n540) );
  OAI2BB2X1 U346 ( .B0(n367), .B1(n7), .A0N(memory[104]), .A1N(n7), .Y(n527)
         );
  OAI2BB2X1 U347 ( .B0(n366), .B1(n7), .A0N(memory[105]), .A1N(n7), .Y(n526)
         );
  OAI2BB2X1 U348 ( .B0(n365), .B1(n7), .A0N(memory[106]), .A1N(n7), .Y(n525)
         );
  OAI2BB2X1 U349 ( .B0(n364), .B1(n7), .A0N(memory[107]), .A1N(n7), .Y(n524)
         );
  OAI2BB2X1 U350 ( .B0(n367), .B1(n8), .A0N(memory[120]), .A1N(n8), .Y(n511)
         );
  OAI2BB2X1 U351 ( .B0(n366), .B1(n8), .A0N(memory[121]), .A1N(n8), .Y(n510)
         );
  OAI2BB2X1 U352 ( .B0(n365), .B1(n8), .A0N(memory[122]), .A1N(n8), .Y(n509)
         );
  OAI2BB2X1 U353 ( .B0(n364), .B1(n8), .A0N(memory[123]), .A1N(n8), .Y(n508)
         );
  OAI2BB2X1 U354 ( .B0(n367), .B1(n9), .A0N(memory[136]), .A1N(n9), .Y(n495)
         );
  OAI2BB2X1 U355 ( .B0(n366), .B1(n9), .A0N(memory[137]), .A1N(n9), .Y(n494)
         );
  OAI2BB2X1 U356 ( .B0(n365), .B1(n9), .A0N(memory[138]), .A1N(n9), .Y(n493)
         );
  OAI2BB2X1 U357 ( .B0(n364), .B1(n9), .A0N(memory[139]), .A1N(n9), .Y(n492)
         );
  OAI2BB2X1 U358 ( .B0(n367), .B1(n10), .A0N(memory[152]), .A1N(n10), .Y(n479)
         );
  OAI2BB2X1 U359 ( .B0(n366), .B1(n10), .A0N(memory[153]), .A1N(n10), .Y(n478)
         );
  OAI2BB2X1 U360 ( .B0(n365), .B1(n10), .A0N(memory[154]), .A1N(n10), .Y(n477)
         );
  OAI2BB2X1 U361 ( .B0(n364), .B1(n10), .A0N(memory[155]), .A1N(n10), .Y(n476)
         );
  OAI2BB2X1 U362 ( .B0(n367), .B1(n11), .A0N(memory[168]), .A1N(n11), .Y(n463)
         );
  OAI2BB2X1 U363 ( .B0(n366), .B1(n11), .A0N(memory[169]), .A1N(n11), .Y(n462)
         );
  OAI2BB2X1 U364 ( .B0(n365), .B1(n11), .A0N(memory[170]), .A1N(n11), .Y(n461)
         );
  OAI2BB2X1 U365 ( .B0(n364), .B1(n11), .A0N(memory[171]), .A1N(n11), .Y(n460)
         );
  OAI2BB2X1 U366 ( .B0(n367), .B1(n12), .A0N(memory[184]), .A1N(n12), .Y(n447)
         );
  OAI2BB2X1 U367 ( .B0(n366), .B1(n12), .A0N(memory[185]), .A1N(n12), .Y(n446)
         );
  OAI2BB2X1 U368 ( .B0(n365), .B1(n12), .A0N(memory[186]), .A1N(n12), .Y(n445)
         );
  OAI2BB2X1 U369 ( .B0(n364), .B1(n12), .A0N(memory[187]), .A1N(n12), .Y(n444)
         );
  OAI2BB2X1 U370 ( .B0(n367), .B1(n13), .A0N(memory[200]), .A1N(n13), .Y(n431)
         );
  OAI2BB2X1 U371 ( .B0(n366), .B1(n13), .A0N(memory[201]), .A1N(n13), .Y(n430)
         );
  OAI2BB2X1 U372 ( .B0(n365), .B1(n13), .A0N(memory[202]), .A1N(n13), .Y(n429)
         );
  OAI2BB2X1 U373 ( .B0(n364), .B1(n13), .A0N(memory[203]), .A1N(n13), .Y(n428)
         );
  OAI2BB2X1 U374 ( .B0(n367), .B1(n14), .A0N(memory[216]), .A1N(n14), .Y(n415)
         );
  OAI2BB2X1 U375 ( .B0(n366), .B1(n14), .A0N(memory[217]), .A1N(n14), .Y(n414)
         );
  OAI2BB2X1 U376 ( .B0(n365), .B1(n14), .A0N(memory[218]), .A1N(n14), .Y(n413)
         );
  OAI2BB2X1 U377 ( .B0(n364), .B1(n14), .A0N(memory[219]), .A1N(n14), .Y(n412)
         );
  OAI2BB2X1 U378 ( .B0(n367), .B1(n15), .A0N(memory[232]), .A1N(n15), .Y(n399)
         );
  OAI2BB2X1 U379 ( .B0(n366), .B1(n15), .A0N(memory[233]), .A1N(n15), .Y(n398)
         );
  OAI2BB2X1 U380 ( .B0(n365), .B1(n15), .A0N(memory[234]), .A1N(n15), .Y(n397)
         );
  OAI2BB2X1 U381 ( .B0(n364), .B1(n15), .A0N(memory[235]), .A1N(n15), .Y(n396)
         );
  OAI2BB2X1 U382 ( .B0(n367), .B1(n16), .A0N(memory[248]), .A1N(n16), .Y(n383)
         );
  OAI2BB2X1 U383 ( .B0(n366), .B1(n16), .A0N(memory[249]), .A1N(n16), .Y(n382)
         );
  OAI2BB2X1 U384 ( .B0(n365), .B1(n16), .A0N(memory[250]), .A1N(n16), .Y(n381)
         );
  OAI2BB2X1 U385 ( .B0(n364), .B1(n16), .A0N(memory[251]), .A1N(n16), .Y(n380)
         );
  NOR2BX1 U386 ( .AN(n636), .B(addr[3]), .Y(n633) );
  BUFX3 U387 ( .A(addr[2]), .Y(n354) );
  INVX1 U388 ( .A(addr[2]), .Y(n359) );
  AND2X2 U389 ( .A(wr_rd), .B(en), .Y(n636) );
  AND2X2 U390 ( .A(addr[3]), .B(n636), .Y(n637) );
  INVX1 U391 ( .A(din[0]), .Y(n375) );
  INVX1 U392 ( .A(din[1]), .Y(n374) );
  INVX1 U393 ( .A(din[2]), .Y(n373) );
  INVX1 U394 ( .A(din[3]), .Y(n372) );
  INVX1 U395 ( .A(din[4]), .Y(n371) );
  INVX1 U396 ( .A(din[5]), .Y(n370) );
  INVX1 U397 ( .A(din[6]), .Y(n369) );
  INVX1 U398 ( .A(din[7]), .Y(n368) );
  INVX1 U399 ( .A(din[8]), .Y(n367) );
  INVX1 U400 ( .A(din[9]), .Y(n366) );
  INVX1 U401 ( .A(din[10]), .Y(n365) );
  INVX1 U402 ( .A(din[11]), .Y(n364) );
  INVX1 U403 ( .A(din[12]), .Y(n363) );
  INVX1 U404 ( .A(din[13]), .Y(n362) );
  INVX1 U405 ( .A(din[14]), .Y(n361) );
  INVX1 U406 ( .A(din[15]), .Y(n360) );
  BUFX3 U407 ( .A(n632), .Y(n356) );
  NAND2BX1 U408 ( .AN(wr_rd), .B(en), .Y(n632) );
endmodule


module mem4x4_1 ( clk, rstn, en, wr_rd, addr, din, dout );
  input [3:0] addr;
  input [15:0] din;
  output [15:0] dout;
  input clk, rstn, en, wr_rd;
  wire   N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48,
         N49, N50, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n23, n25, n27, n28, n30, n31, n34, n36,
         n38, n40, n41, n42, n43, n44, n46, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643;
  wire   [255:0] memory;

  DFFRHQX1 memory_reg_1__15_ ( .D(n392), .CK(clk), .RN(rstn), .Q(memory[239])
         );
  DFFRHQX1 memory_reg_1__14_ ( .D(n393), .CK(clk), .RN(rstn), .Q(memory[238])
         );
  DFFRHQX1 memory_reg_1__13_ ( .D(n394), .CK(clk), .RN(rstn), .Q(memory[237])
         );
  DFFRHQX1 memory_reg_1__12_ ( .D(n395), .CK(clk), .RN(rstn), .Q(memory[236])
         );
  DFFRHQX1 memory_reg_1__11_ ( .D(n396), .CK(clk), .RN(rstn), .Q(memory[235])
         );
  DFFRHQX1 memory_reg_1__10_ ( .D(n397), .CK(clk), .RN(rstn), .Q(memory[234])
         );
  DFFRHQX1 memory_reg_1__9_ ( .D(n398), .CK(clk), .RN(rstn), .Q(memory[233])
         );
  DFFRHQX1 memory_reg_1__8_ ( .D(n399), .CK(clk), .RN(rstn), .Q(memory[232])
         );
  DFFRHQX1 memory_reg_1__7_ ( .D(n400), .CK(clk), .RN(rstn), .Q(memory[231])
         );
  DFFRHQX1 memory_reg_1__6_ ( .D(n401), .CK(clk), .RN(rstn), .Q(memory[230])
         );
  DFFRHQX1 memory_reg_1__5_ ( .D(n402), .CK(clk), .RN(rstn), .Q(memory[229])
         );
  DFFRHQX1 memory_reg_1__4_ ( .D(n403), .CK(clk), .RN(rstn), .Q(memory[228])
         );
  DFFRHQX1 memory_reg_1__3_ ( .D(n404), .CK(clk), .RN(rstn), .Q(memory[227])
         );
  DFFRHQX1 memory_reg_1__2_ ( .D(n405), .CK(clk), .RN(rstn), .Q(memory[226])
         );
  DFFRHQX1 memory_reg_1__1_ ( .D(n406), .CK(clk), .RN(rstn), .Q(memory[225])
         );
  DFFRHQX1 memory_reg_1__0_ ( .D(n407), .CK(clk), .RN(rstn), .Q(memory[224])
         );
  DFFRHQX1 memory_reg_5__15_ ( .D(n456), .CK(clk), .RN(rstn), .Q(memory[175])
         );
  DFFRHQX1 memory_reg_5__14_ ( .D(n457), .CK(clk), .RN(rstn), .Q(memory[174])
         );
  DFFRHQX1 memory_reg_5__13_ ( .D(n458), .CK(clk), .RN(rstn), .Q(memory[173])
         );
  DFFRHQX1 memory_reg_5__12_ ( .D(n459), .CK(clk), .RN(rstn), .Q(memory[172])
         );
  DFFRHQX1 memory_reg_5__11_ ( .D(n460), .CK(clk), .RN(rstn), .Q(memory[171])
         );
  DFFRHQX1 memory_reg_5__10_ ( .D(n461), .CK(clk), .RN(rstn), .Q(memory[170])
         );
  DFFRHQX1 memory_reg_5__9_ ( .D(n462), .CK(clk), .RN(rstn), .Q(memory[169])
         );
  DFFRHQX1 memory_reg_5__8_ ( .D(n463), .CK(clk), .RN(rstn), .Q(memory[168])
         );
  DFFRHQX1 memory_reg_5__7_ ( .D(n464), .CK(clk), .RN(rstn), .Q(memory[167])
         );
  DFFRHQX1 memory_reg_5__6_ ( .D(n465), .CK(clk), .RN(rstn), .Q(memory[166])
         );
  DFFRHQX1 memory_reg_5__5_ ( .D(n466), .CK(clk), .RN(rstn), .Q(memory[165])
         );
  DFFRHQX1 memory_reg_5__4_ ( .D(n467), .CK(clk), .RN(rstn), .Q(memory[164])
         );
  DFFRHQX1 memory_reg_5__3_ ( .D(n468), .CK(clk), .RN(rstn), .Q(memory[163])
         );
  DFFRHQX1 memory_reg_5__2_ ( .D(n469), .CK(clk), .RN(rstn), .Q(memory[162])
         );
  DFFRHQX1 memory_reg_5__1_ ( .D(n470), .CK(clk), .RN(rstn), .Q(memory[161])
         );
  DFFRHQX1 memory_reg_5__0_ ( .D(n471), .CK(clk), .RN(rstn), .Q(memory[160])
         );
  DFFRHQX1 memory_reg_9__15_ ( .D(n520), .CK(clk), .RN(rstn), .Q(memory[111])
         );
  DFFRHQX1 memory_reg_9__14_ ( .D(n521), .CK(clk), .RN(rstn), .Q(memory[110])
         );
  DFFRHQX1 memory_reg_9__13_ ( .D(n522), .CK(clk), .RN(rstn), .Q(memory[109])
         );
  DFFRHQX1 memory_reg_9__12_ ( .D(n523), .CK(clk), .RN(rstn), .Q(memory[108])
         );
  DFFRHQX1 memory_reg_9__11_ ( .D(n524), .CK(clk), .RN(rstn), .Q(memory[107])
         );
  DFFRHQX1 memory_reg_9__10_ ( .D(n525), .CK(clk), .RN(rstn), .Q(memory[106])
         );
  DFFRHQX1 memory_reg_9__9_ ( .D(n526), .CK(clk), .RN(rstn), .Q(memory[105])
         );
  DFFRHQX1 memory_reg_9__8_ ( .D(n527), .CK(clk), .RN(rstn), .Q(memory[104])
         );
  DFFRHQX1 memory_reg_9__7_ ( .D(n528), .CK(clk), .RN(rstn), .Q(memory[103])
         );
  DFFRHQX1 memory_reg_9__6_ ( .D(n529), .CK(clk), .RN(rstn), .Q(memory[102])
         );
  DFFRHQX1 memory_reg_9__5_ ( .D(n530), .CK(clk), .RN(rstn), .Q(memory[101])
         );
  DFFRHQX1 memory_reg_9__4_ ( .D(n531), .CK(clk), .RN(rstn), .Q(memory[100])
         );
  DFFRHQX1 memory_reg_9__3_ ( .D(n532), .CK(clk), .RN(rstn), .Q(memory[99]) );
  DFFRHQX1 memory_reg_9__2_ ( .D(n533), .CK(clk), .RN(rstn), .Q(memory[98]) );
  DFFRHQX1 memory_reg_9__1_ ( .D(n534), .CK(clk), .RN(rstn), .Q(memory[97]) );
  DFFRHQX1 memory_reg_9__0_ ( .D(n535), .CK(clk), .RN(rstn), .Q(memory[96]) );
  DFFRHQX1 memory_reg_13__15_ ( .D(n584), .CK(clk), .RN(rstn), .Q(memory[47])
         );
  DFFRHQX1 memory_reg_13__14_ ( .D(n585), .CK(clk), .RN(rstn), .Q(memory[46])
         );
  DFFRHQX1 memory_reg_13__13_ ( .D(n586), .CK(clk), .RN(rstn), .Q(memory[45])
         );
  DFFRHQX1 memory_reg_13__12_ ( .D(n587), .CK(clk), .RN(rstn), .Q(memory[44])
         );
  DFFRHQX1 memory_reg_13__11_ ( .D(n588), .CK(clk), .RN(rstn), .Q(memory[43])
         );
  DFFRHQX1 memory_reg_13__10_ ( .D(n589), .CK(clk), .RN(rstn), .Q(memory[42])
         );
  DFFRHQX1 memory_reg_13__9_ ( .D(n590), .CK(clk), .RN(rstn), .Q(memory[41])
         );
  DFFRHQX1 memory_reg_13__8_ ( .D(n591), .CK(clk), .RN(rstn), .Q(memory[40])
         );
  DFFRHQX1 memory_reg_13__7_ ( .D(n592), .CK(clk), .RN(rstn), .Q(memory[39])
         );
  DFFRHQX1 memory_reg_13__6_ ( .D(n593), .CK(clk), .RN(rstn), .Q(memory[38])
         );
  DFFRHQX1 memory_reg_13__5_ ( .D(n594), .CK(clk), .RN(rstn), .Q(memory[37])
         );
  DFFRHQX1 memory_reg_13__4_ ( .D(n595), .CK(clk), .RN(rstn), .Q(memory[36])
         );
  DFFRHQX1 memory_reg_13__3_ ( .D(n596), .CK(clk), .RN(rstn), .Q(memory[35])
         );
  DFFRHQX1 memory_reg_13__2_ ( .D(n597), .CK(clk), .RN(rstn), .Q(memory[34])
         );
  DFFRHQX1 memory_reg_13__1_ ( .D(n598), .CK(clk), .RN(rstn), .Q(memory[33])
         );
  DFFRHQX1 memory_reg_13__0_ ( .D(n599), .CK(clk), .RN(rstn), .Q(memory[32])
         );
  DFFRHQX1 memory_reg_3__15_ ( .D(n424), .CK(clk), .RN(rstn), .Q(memory[207])
         );
  DFFRHQX1 memory_reg_3__14_ ( .D(n425), .CK(clk), .RN(rstn), .Q(memory[206])
         );
  DFFRHQX1 memory_reg_3__13_ ( .D(n426), .CK(clk), .RN(rstn), .Q(memory[205])
         );
  DFFRHQX1 memory_reg_3__12_ ( .D(n427), .CK(clk), .RN(rstn), .Q(memory[204])
         );
  DFFRHQX1 memory_reg_3__11_ ( .D(n428), .CK(clk), .RN(rstn), .Q(memory[203])
         );
  DFFRHQX1 memory_reg_3__10_ ( .D(n429), .CK(clk), .RN(rstn), .Q(memory[202])
         );
  DFFRHQX1 memory_reg_3__9_ ( .D(n430), .CK(clk), .RN(rstn), .Q(memory[201])
         );
  DFFRHQX1 memory_reg_3__8_ ( .D(n431), .CK(clk), .RN(rstn), .Q(memory[200])
         );
  DFFRHQX1 memory_reg_3__7_ ( .D(n432), .CK(clk), .RN(rstn), .Q(memory[199])
         );
  DFFRHQX1 memory_reg_3__6_ ( .D(n433), .CK(clk), .RN(rstn), .Q(memory[198])
         );
  DFFRHQX1 memory_reg_3__5_ ( .D(n434), .CK(clk), .RN(rstn), .Q(memory[197])
         );
  DFFRHQX1 memory_reg_3__4_ ( .D(n435), .CK(clk), .RN(rstn), .Q(memory[196])
         );
  DFFRHQX1 memory_reg_3__3_ ( .D(n436), .CK(clk), .RN(rstn), .Q(memory[195])
         );
  DFFRHQX1 memory_reg_3__2_ ( .D(n437), .CK(clk), .RN(rstn), .Q(memory[194])
         );
  DFFRHQX1 memory_reg_3__1_ ( .D(n438), .CK(clk), .RN(rstn), .Q(memory[193])
         );
  DFFRHQX1 memory_reg_3__0_ ( .D(n439), .CK(clk), .RN(rstn), .Q(memory[192])
         );
  DFFRHQX1 memory_reg_7__15_ ( .D(n488), .CK(clk), .RN(rstn), .Q(memory[143])
         );
  DFFRHQX1 memory_reg_7__14_ ( .D(n489), .CK(clk), .RN(rstn), .Q(memory[142])
         );
  DFFRHQX1 memory_reg_7__13_ ( .D(n490), .CK(clk), .RN(rstn), .Q(memory[141])
         );
  DFFRHQX1 memory_reg_7__12_ ( .D(n491), .CK(clk), .RN(rstn), .Q(memory[140])
         );
  DFFRHQX1 memory_reg_7__11_ ( .D(n492), .CK(clk), .RN(rstn), .Q(memory[139])
         );
  DFFRHQX1 memory_reg_7__10_ ( .D(n493), .CK(clk), .RN(rstn), .Q(memory[138])
         );
  DFFRHQX1 memory_reg_7__9_ ( .D(n494), .CK(clk), .RN(rstn), .Q(memory[137])
         );
  DFFRHQX1 memory_reg_7__8_ ( .D(n495), .CK(clk), .RN(rstn), .Q(memory[136])
         );
  DFFRHQX1 memory_reg_7__7_ ( .D(n496), .CK(clk), .RN(rstn), .Q(memory[135])
         );
  DFFRHQX1 memory_reg_7__6_ ( .D(n497), .CK(clk), .RN(rstn), .Q(memory[134])
         );
  DFFRHQX1 memory_reg_7__5_ ( .D(n498), .CK(clk), .RN(rstn), .Q(memory[133])
         );
  DFFRHQX1 memory_reg_7__4_ ( .D(n499), .CK(clk), .RN(rstn), .Q(memory[132])
         );
  DFFRHQX1 memory_reg_7__3_ ( .D(n500), .CK(clk), .RN(rstn), .Q(memory[131])
         );
  DFFRHQX1 memory_reg_7__2_ ( .D(n501), .CK(clk), .RN(rstn), .Q(memory[130])
         );
  DFFRHQX1 memory_reg_7__1_ ( .D(n502), .CK(clk), .RN(rstn), .Q(memory[129])
         );
  DFFRHQX1 memory_reg_7__0_ ( .D(n503), .CK(clk), .RN(rstn), .Q(memory[128])
         );
  DFFRHQX1 memory_reg_11__15_ ( .D(n552), .CK(clk), .RN(rstn), .Q(memory[79])
         );
  DFFRHQX1 memory_reg_11__14_ ( .D(n553), .CK(clk), .RN(rstn), .Q(memory[78])
         );
  DFFRHQX1 memory_reg_11__13_ ( .D(n554), .CK(clk), .RN(rstn), .Q(memory[77])
         );
  DFFRHQX1 memory_reg_11__12_ ( .D(n555), .CK(clk), .RN(rstn), .Q(memory[76])
         );
  DFFRHQX1 memory_reg_11__11_ ( .D(n556), .CK(clk), .RN(rstn), .Q(memory[75])
         );
  DFFRHQX1 memory_reg_11__10_ ( .D(n557), .CK(clk), .RN(rstn), .Q(memory[74])
         );
  DFFRHQX1 memory_reg_11__9_ ( .D(n558), .CK(clk), .RN(rstn), .Q(memory[73])
         );
  DFFRHQX1 memory_reg_11__8_ ( .D(n559), .CK(clk), .RN(rstn), .Q(memory[72])
         );
  DFFRHQX1 memory_reg_11__7_ ( .D(n560), .CK(clk), .RN(rstn), .Q(memory[71])
         );
  DFFRHQX1 memory_reg_11__6_ ( .D(n561), .CK(clk), .RN(rstn), .Q(memory[70])
         );
  DFFRHQX1 memory_reg_11__5_ ( .D(n562), .CK(clk), .RN(rstn), .Q(memory[69])
         );
  DFFRHQX1 memory_reg_11__4_ ( .D(n563), .CK(clk), .RN(rstn), .Q(memory[68])
         );
  DFFRHQX1 memory_reg_11__3_ ( .D(n564), .CK(clk), .RN(rstn), .Q(memory[67])
         );
  DFFRHQX1 memory_reg_11__2_ ( .D(n565), .CK(clk), .RN(rstn), .Q(memory[66])
         );
  DFFRHQX1 memory_reg_11__1_ ( .D(n566), .CK(clk), .RN(rstn), .Q(memory[65])
         );
  DFFRHQX1 memory_reg_11__0_ ( .D(n567), .CK(clk), .RN(rstn), .Q(memory[64])
         );
  DFFRHQX1 memory_reg_15__15_ ( .D(n616), .CK(clk), .RN(rstn), .Q(memory[15])
         );
  DFFRHQX1 memory_reg_15__14_ ( .D(n617), .CK(clk), .RN(rstn), .Q(memory[14])
         );
  DFFRHQX1 memory_reg_15__13_ ( .D(n618), .CK(clk), .RN(rstn), .Q(memory[13])
         );
  DFFRHQX1 memory_reg_15__12_ ( .D(n619), .CK(clk), .RN(rstn), .Q(memory[12])
         );
  DFFRHQX1 memory_reg_15__11_ ( .D(n620), .CK(clk), .RN(rstn), .Q(memory[11])
         );
  DFFRHQX1 memory_reg_15__10_ ( .D(n621), .CK(clk), .RN(rstn), .Q(memory[10])
         );
  DFFRHQX1 memory_reg_15__9_ ( .D(n622), .CK(clk), .RN(rstn), .Q(memory[9]) );
  DFFRHQX1 memory_reg_15__8_ ( .D(n623), .CK(clk), .RN(rstn), .Q(memory[8]) );
  DFFRHQX1 memory_reg_15__7_ ( .D(n624), .CK(clk), .RN(rstn), .Q(memory[7]) );
  DFFRHQX1 memory_reg_15__6_ ( .D(n625), .CK(clk), .RN(rstn), .Q(memory[6]) );
  DFFRHQX1 memory_reg_15__5_ ( .D(n626), .CK(clk), .RN(rstn), .Q(memory[5]) );
  DFFRHQX1 memory_reg_15__4_ ( .D(n627), .CK(clk), .RN(rstn), .Q(memory[4]) );
  DFFRHQX1 memory_reg_15__3_ ( .D(n628), .CK(clk), .RN(rstn), .Q(memory[3]) );
  DFFRHQX1 memory_reg_15__2_ ( .D(n629), .CK(clk), .RN(rstn), .Q(memory[2]) );
  DFFRHQX1 memory_reg_15__1_ ( .D(n630), .CK(clk), .RN(rstn), .Q(memory[1]) );
  DFFRHQX1 memory_reg_15__0_ ( .D(n631), .CK(clk), .RN(rstn), .Q(memory[0]) );
  DFFRHQX1 memory_reg_0__15_ ( .D(n376), .CK(clk), .RN(rstn), .Q(memory[255])
         );
  DFFRHQX1 memory_reg_0__14_ ( .D(n377), .CK(clk), .RN(rstn), .Q(memory[254])
         );
  DFFRHQX1 memory_reg_0__13_ ( .D(n378), .CK(clk), .RN(rstn), .Q(memory[253])
         );
  DFFRHQX1 memory_reg_0__12_ ( .D(n379), .CK(clk), .RN(rstn), .Q(memory[252])
         );
  DFFRHQX1 memory_reg_0__11_ ( .D(n380), .CK(clk), .RN(rstn), .Q(memory[251])
         );
  DFFRHQX1 memory_reg_0__10_ ( .D(n381), .CK(clk), .RN(rstn), .Q(memory[250])
         );
  DFFRHQX1 memory_reg_0__9_ ( .D(n382), .CK(clk), .RN(rstn), .Q(memory[249])
         );
  DFFRHQX1 memory_reg_0__8_ ( .D(n383), .CK(clk), .RN(rstn), .Q(memory[248])
         );
  DFFRHQX1 memory_reg_0__7_ ( .D(n384), .CK(clk), .RN(rstn), .Q(memory[247])
         );
  DFFRHQX1 memory_reg_0__6_ ( .D(n385), .CK(clk), .RN(rstn), .Q(memory[246])
         );
  DFFRHQX1 memory_reg_0__5_ ( .D(n386), .CK(clk), .RN(rstn), .Q(memory[245])
         );
  DFFRHQX1 memory_reg_0__4_ ( .D(n387), .CK(clk), .RN(rstn), .Q(memory[244])
         );
  DFFRHQX1 memory_reg_0__3_ ( .D(n388), .CK(clk), .RN(rstn), .Q(memory[243])
         );
  DFFRHQX1 memory_reg_0__2_ ( .D(n389), .CK(clk), .RN(rstn), .Q(memory[242])
         );
  DFFRHQX1 memory_reg_0__1_ ( .D(n390), .CK(clk), .RN(rstn), .Q(memory[241])
         );
  DFFRHQX1 memory_reg_0__0_ ( .D(n391), .CK(clk), .RN(rstn), .Q(memory[240])
         );
  DFFRHQX1 memory_reg_4__15_ ( .D(n440), .CK(clk), .RN(rstn), .Q(memory[191])
         );
  DFFRHQX1 memory_reg_4__14_ ( .D(n441), .CK(clk), .RN(rstn), .Q(memory[190])
         );
  DFFRHQX1 memory_reg_4__13_ ( .D(n442), .CK(clk), .RN(rstn), .Q(memory[189])
         );
  DFFRHQX1 memory_reg_4__12_ ( .D(n443), .CK(clk), .RN(rstn), .Q(memory[188])
         );
  DFFRHQX1 memory_reg_4__11_ ( .D(n444), .CK(clk), .RN(rstn), .Q(memory[187])
         );
  DFFRHQX1 memory_reg_4__10_ ( .D(n445), .CK(clk), .RN(rstn), .Q(memory[186])
         );
  DFFRHQX1 memory_reg_4__9_ ( .D(n446), .CK(clk), .RN(rstn), .Q(memory[185])
         );
  DFFRHQX1 memory_reg_4__8_ ( .D(n447), .CK(clk), .RN(rstn), .Q(memory[184])
         );
  DFFRHQX1 memory_reg_4__7_ ( .D(n448), .CK(clk), .RN(rstn), .Q(memory[183])
         );
  DFFRHQX1 memory_reg_4__6_ ( .D(n449), .CK(clk), .RN(rstn), .Q(memory[182])
         );
  DFFRHQX1 memory_reg_4__5_ ( .D(n450), .CK(clk), .RN(rstn), .Q(memory[181])
         );
  DFFRHQX1 memory_reg_4__4_ ( .D(n451), .CK(clk), .RN(rstn), .Q(memory[180])
         );
  DFFRHQX1 memory_reg_4__3_ ( .D(n452), .CK(clk), .RN(rstn), .Q(memory[179])
         );
  DFFRHQX1 memory_reg_4__2_ ( .D(n453), .CK(clk), .RN(rstn), .Q(memory[178])
         );
  DFFRHQX1 memory_reg_4__1_ ( .D(n454), .CK(clk), .RN(rstn), .Q(memory[177])
         );
  DFFRHQX1 memory_reg_4__0_ ( .D(n455), .CK(clk), .RN(rstn), .Q(memory[176])
         );
  DFFRHQX1 memory_reg_8__15_ ( .D(n504), .CK(clk), .RN(rstn), .Q(memory[127])
         );
  DFFRHQX1 memory_reg_8__14_ ( .D(n505), .CK(clk), .RN(rstn), .Q(memory[126])
         );
  DFFRHQX1 memory_reg_8__13_ ( .D(n506), .CK(clk), .RN(rstn), .Q(memory[125])
         );
  DFFRHQX1 memory_reg_8__12_ ( .D(n507), .CK(clk), .RN(rstn), .Q(memory[124])
         );
  DFFRHQX1 memory_reg_8__11_ ( .D(n508), .CK(clk), .RN(rstn), .Q(memory[123])
         );
  DFFRHQX1 memory_reg_8__10_ ( .D(n509), .CK(clk), .RN(rstn), .Q(memory[122])
         );
  DFFRHQX1 memory_reg_8__9_ ( .D(n510), .CK(clk), .RN(rstn), .Q(memory[121])
         );
  DFFRHQX1 memory_reg_8__8_ ( .D(n511), .CK(clk), .RN(rstn), .Q(memory[120])
         );
  DFFRHQX1 memory_reg_8__7_ ( .D(n512), .CK(clk), .RN(rstn), .Q(memory[119])
         );
  DFFRHQX1 memory_reg_8__6_ ( .D(n513), .CK(clk), .RN(rstn), .Q(memory[118])
         );
  DFFRHQX1 memory_reg_8__5_ ( .D(n514), .CK(clk), .RN(rstn), .Q(memory[117])
         );
  DFFRHQX1 memory_reg_8__4_ ( .D(n515), .CK(clk), .RN(rstn), .Q(memory[116])
         );
  DFFRHQX1 memory_reg_8__3_ ( .D(n516), .CK(clk), .RN(rstn), .Q(memory[115])
         );
  DFFRHQX1 memory_reg_8__2_ ( .D(n517), .CK(clk), .RN(rstn), .Q(memory[114])
         );
  DFFRHQX1 memory_reg_8__1_ ( .D(n518), .CK(clk), .RN(rstn), .Q(memory[113])
         );
  DFFRHQX1 memory_reg_8__0_ ( .D(n519), .CK(clk), .RN(rstn), .Q(memory[112])
         );
  DFFRHQX1 memory_reg_12__15_ ( .D(n568), .CK(clk), .RN(rstn), .Q(memory[63])
         );
  DFFRHQX1 memory_reg_12__14_ ( .D(n569), .CK(clk), .RN(rstn), .Q(memory[62])
         );
  DFFRHQX1 memory_reg_12__13_ ( .D(n570), .CK(clk), .RN(rstn), .Q(memory[61])
         );
  DFFRHQX1 memory_reg_12__12_ ( .D(n571), .CK(clk), .RN(rstn), .Q(memory[60])
         );
  DFFRHQX1 memory_reg_12__11_ ( .D(n572), .CK(clk), .RN(rstn), .Q(memory[59])
         );
  DFFRHQX1 memory_reg_12__10_ ( .D(n573), .CK(clk), .RN(rstn), .Q(memory[58])
         );
  DFFRHQX1 memory_reg_12__9_ ( .D(n574), .CK(clk), .RN(rstn), .Q(memory[57])
         );
  DFFRHQX1 memory_reg_12__8_ ( .D(n575), .CK(clk), .RN(rstn), .Q(memory[56])
         );
  DFFRHQX1 memory_reg_12__7_ ( .D(n576), .CK(clk), .RN(rstn), .Q(memory[55])
         );
  DFFRHQX1 memory_reg_12__6_ ( .D(n577), .CK(clk), .RN(rstn), .Q(memory[54])
         );
  DFFRHQX1 memory_reg_12__5_ ( .D(n578), .CK(clk), .RN(rstn), .Q(memory[53])
         );
  DFFRHQX1 memory_reg_12__4_ ( .D(n579), .CK(clk), .RN(rstn), .Q(memory[52])
         );
  DFFRHQX1 memory_reg_12__3_ ( .D(n580), .CK(clk), .RN(rstn), .Q(memory[51])
         );
  DFFRHQX1 memory_reg_12__2_ ( .D(n581), .CK(clk), .RN(rstn), .Q(memory[50])
         );
  DFFRHQX1 memory_reg_12__1_ ( .D(n582), .CK(clk), .RN(rstn), .Q(memory[49])
         );
  DFFRHQX1 memory_reg_12__0_ ( .D(n583), .CK(clk), .RN(rstn), .Q(memory[48])
         );
  DFFRHQX1 memory_reg_2__15_ ( .D(n408), .CK(clk), .RN(rstn), .Q(memory[223])
         );
  DFFRHQX1 memory_reg_2__14_ ( .D(n409), .CK(clk), .RN(rstn), .Q(memory[222])
         );
  DFFRHQX1 memory_reg_2__13_ ( .D(n410), .CK(clk), .RN(rstn), .Q(memory[221])
         );
  DFFRHQX1 memory_reg_2__12_ ( .D(n411), .CK(clk), .RN(rstn), .Q(memory[220])
         );
  DFFRHQX1 memory_reg_2__11_ ( .D(n412), .CK(clk), .RN(rstn), .Q(memory[219])
         );
  DFFRHQX1 memory_reg_2__10_ ( .D(n413), .CK(clk), .RN(rstn), .Q(memory[218])
         );
  DFFRHQX1 memory_reg_2__9_ ( .D(n414), .CK(clk), .RN(rstn), .Q(memory[217])
         );
  DFFRHQX1 memory_reg_2__8_ ( .D(n415), .CK(clk), .RN(rstn), .Q(memory[216])
         );
  DFFRHQX1 memory_reg_2__7_ ( .D(n416), .CK(clk), .RN(rstn), .Q(memory[215])
         );
  DFFRHQX1 memory_reg_2__6_ ( .D(n417), .CK(clk), .RN(rstn), .Q(memory[214])
         );
  DFFRHQX1 memory_reg_2__5_ ( .D(n418), .CK(clk), .RN(rstn), .Q(memory[213])
         );
  DFFRHQX1 memory_reg_2__4_ ( .D(n419), .CK(clk), .RN(rstn), .Q(memory[212])
         );
  DFFRHQX1 memory_reg_2__3_ ( .D(n420), .CK(clk), .RN(rstn), .Q(memory[211])
         );
  DFFRHQX1 memory_reg_2__2_ ( .D(n421), .CK(clk), .RN(rstn), .Q(memory[210])
         );
  DFFRHQX1 memory_reg_2__1_ ( .D(n422), .CK(clk), .RN(rstn), .Q(memory[209])
         );
  DFFRHQX1 memory_reg_2__0_ ( .D(n423), .CK(clk), .RN(rstn), .Q(memory[208])
         );
  DFFRHQX1 memory_reg_6__15_ ( .D(n472), .CK(clk), .RN(rstn), .Q(memory[159])
         );
  DFFRHQX1 memory_reg_6__14_ ( .D(n473), .CK(clk), .RN(rstn), .Q(memory[158])
         );
  DFFRHQX1 memory_reg_6__13_ ( .D(n474), .CK(clk), .RN(rstn), .Q(memory[157])
         );
  DFFRHQX1 memory_reg_6__12_ ( .D(n475), .CK(clk), .RN(rstn), .Q(memory[156])
         );
  DFFRHQX1 memory_reg_6__11_ ( .D(n476), .CK(clk), .RN(rstn), .Q(memory[155])
         );
  DFFRHQX1 memory_reg_6__10_ ( .D(n477), .CK(clk), .RN(rstn), .Q(memory[154])
         );
  DFFRHQX1 memory_reg_6__9_ ( .D(n478), .CK(clk), .RN(rstn), .Q(memory[153])
         );
  DFFRHQX1 memory_reg_6__8_ ( .D(n479), .CK(clk), .RN(rstn), .Q(memory[152])
         );
  DFFRHQX1 memory_reg_6__7_ ( .D(n480), .CK(clk), .RN(rstn), .Q(memory[151])
         );
  DFFRHQX1 memory_reg_6__6_ ( .D(n481), .CK(clk), .RN(rstn), .Q(memory[150])
         );
  DFFRHQX1 memory_reg_6__5_ ( .D(n482), .CK(clk), .RN(rstn), .Q(memory[149])
         );
  DFFRHQX1 memory_reg_6__4_ ( .D(n483), .CK(clk), .RN(rstn), .Q(memory[148])
         );
  DFFRHQX1 memory_reg_6__3_ ( .D(n484), .CK(clk), .RN(rstn), .Q(memory[147])
         );
  DFFRHQX1 memory_reg_6__2_ ( .D(n485), .CK(clk), .RN(rstn), .Q(memory[146])
         );
  DFFRHQX1 memory_reg_6__1_ ( .D(n486), .CK(clk), .RN(rstn), .Q(memory[145])
         );
  DFFRHQX1 memory_reg_6__0_ ( .D(n487), .CK(clk), .RN(rstn), .Q(memory[144])
         );
  DFFRHQX1 memory_reg_10__15_ ( .D(n536), .CK(clk), .RN(rstn), .Q(memory[95])
         );
  DFFRHQX1 memory_reg_10__14_ ( .D(n537), .CK(clk), .RN(rstn), .Q(memory[94])
         );
  DFFRHQX1 memory_reg_10__13_ ( .D(n538), .CK(clk), .RN(rstn), .Q(memory[93])
         );
  DFFRHQX1 memory_reg_10__12_ ( .D(n539), .CK(clk), .RN(rstn), .Q(memory[92])
         );
  DFFRHQX1 memory_reg_10__11_ ( .D(n540), .CK(clk), .RN(rstn), .Q(memory[91])
         );
  DFFRHQX1 memory_reg_10__10_ ( .D(n541), .CK(clk), .RN(rstn), .Q(memory[90])
         );
  DFFRHQX1 memory_reg_10__9_ ( .D(n542), .CK(clk), .RN(rstn), .Q(memory[89])
         );
  DFFRHQX1 memory_reg_10__8_ ( .D(n543), .CK(clk), .RN(rstn), .Q(memory[88])
         );
  DFFRHQX1 memory_reg_10__7_ ( .D(n544), .CK(clk), .RN(rstn), .Q(memory[87])
         );
  DFFRHQX1 memory_reg_10__6_ ( .D(n545), .CK(clk), .RN(rstn), .Q(memory[86])
         );
  DFFRHQX1 memory_reg_10__5_ ( .D(n546), .CK(clk), .RN(rstn), .Q(memory[85])
         );
  DFFRHQX1 memory_reg_10__4_ ( .D(n547), .CK(clk), .RN(rstn), .Q(memory[84])
         );
  DFFRHQX1 memory_reg_10__3_ ( .D(n548), .CK(clk), .RN(rstn), .Q(memory[83])
         );
  DFFRHQX1 memory_reg_10__2_ ( .D(n549), .CK(clk), .RN(rstn), .Q(memory[82])
         );
  DFFRHQX1 memory_reg_10__1_ ( .D(n550), .CK(clk), .RN(rstn), .Q(memory[81])
         );
  DFFRHQX1 memory_reg_10__0_ ( .D(n551), .CK(clk), .RN(rstn), .Q(memory[80])
         );
  DFFRHQX1 memory_reg_14__15_ ( .D(n600), .CK(clk), .RN(rstn), .Q(memory[31])
         );
  DFFRHQX1 memory_reg_14__14_ ( .D(n601), .CK(clk), .RN(rstn), .Q(memory[30])
         );
  DFFRHQX1 memory_reg_14__13_ ( .D(n602), .CK(clk), .RN(rstn), .Q(memory[29])
         );
  DFFRHQX1 memory_reg_14__12_ ( .D(n603), .CK(clk), .RN(rstn), .Q(memory[28])
         );
  DFFRHQX1 memory_reg_14__11_ ( .D(n604), .CK(clk), .RN(rstn), .Q(memory[27])
         );
  DFFRHQX1 memory_reg_14__10_ ( .D(n605), .CK(clk), .RN(rstn), .Q(memory[26])
         );
  DFFRHQX1 memory_reg_14__9_ ( .D(n606), .CK(clk), .RN(rstn), .Q(memory[25])
         );
  DFFRHQX1 memory_reg_14__8_ ( .D(n607), .CK(clk), .RN(rstn), .Q(memory[24])
         );
  DFFRHQX1 memory_reg_14__7_ ( .D(n608), .CK(clk), .RN(rstn), .Q(memory[23])
         );
  DFFRHQX1 memory_reg_14__6_ ( .D(n609), .CK(clk), .RN(rstn), .Q(memory[22])
         );
  DFFRHQX1 memory_reg_14__5_ ( .D(n610), .CK(clk), .RN(rstn), .Q(memory[21])
         );
  DFFRHQX1 memory_reg_14__4_ ( .D(n611), .CK(clk), .RN(rstn), .Q(memory[20])
         );
  DFFRHQX1 memory_reg_14__3_ ( .D(n612), .CK(clk), .RN(rstn), .Q(memory[19])
         );
  DFFRHQX1 memory_reg_14__2_ ( .D(n613), .CK(clk), .RN(rstn), .Q(memory[18])
         );
  DFFRHQX1 memory_reg_14__1_ ( .D(n614), .CK(clk), .RN(rstn), .Q(memory[17])
         );
  DFFRHQX1 memory_reg_14__0_ ( .D(n615), .CK(clk), .RN(rstn), .Q(memory[16])
         );
  NAND2X1 U2 ( .A(n643), .B(n642), .Y(n1) );
  NAND2X1 U3 ( .A(n641), .B(n643), .Y(n2) );
  NAND2X1 U4 ( .A(n640), .B(n642), .Y(n3) );
  NAND2X1 U5 ( .A(n640), .B(n641), .Y(n4) );
  NAND2X1 U6 ( .A(n639), .B(n642), .Y(n5) );
  NAND2X1 U7 ( .A(n639), .B(n641), .Y(n6) );
  NAND2X1 U8 ( .A(n638), .B(n642), .Y(n7) );
  NAND2X1 U9 ( .A(n638), .B(n641), .Y(n8) );
  NAND2X1 U10 ( .A(n635), .B(n643), .Y(n9) );
  NAND2X1 U11 ( .A(n634), .B(n643), .Y(n10) );
  NAND2X1 U12 ( .A(n635), .B(n640), .Y(n11) );
  NAND2X1 U13 ( .A(n634), .B(n640), .Y(n12) );
  NAND2X1 U14 ( .A(n635), .B(n639), .Y(n13) );
  NAND2X1 U15 ( .A(n634), .B(n639), .Y(n14) );
  NAND2X1 U16 ( .A(n635), .B(n638), .Y(n15) );
  NAND2X1 U17 ( .A(n634), .B(n638), .Y(n16) );
  INVX1 U18 ( .A(n357), .Y(n351) );
  INVX1 U19 ( .A(n357), .Y(n352) );
  INVX1 U20 ( .A(n357), .Y(n353) );
  INVX1 U21 ( .A(n358), .Y(n349) );
  INVX1 U22 ( .A(n358), .Y(n350) );
  NOR2X1 U23 ( .A(n359), .B(addr[1]), .Y(n640) );
  NOR2X1 U24 ( .A(n359), .B(n358), .Y(n643) );
  AND2X2 U25 ( .A(n633), .B(addr[0]), .Y(n635) );
  AND2X2 U26 ( .A(n633), .B(n357), .Y(n634) );
  AND2X2 U27 ( .A(n637), .B(n357), .Y(n641) );
  AND2X2 U28 ( .A(n637), .B(addr[0]), .Y(n642) );
  MX4X1 U29 ( .A(memory[176]), .B(memory[160]), .C(memory[144]), .D(
        memory[128]), .S0(n352), .S1(n350), .Y(n19) );
  MX4X1 U30 ( .A(memory[177]), .B(memory[161]), .C(memory[145]), .D(
        memory[129]), .S0(n351), .S1(n349), .Y(n27) );
  MX4X1 U31 ( .A(memory[178]), .B(memory[162]), .C(memory[146]), .D(
        memory[130]), .S0(n351), .S1(n349), .Y(n34) );
  MX4X1 U32 ( .A(memory[179]), .B(memory[163]), .C(memory[147]), .D(
        memory[131]), .S0(n351), .S1(n349), .Y(n41) );
  MX4X1 U33 ( .A(memory[180]), .B(memory[164]), .C(memory[148]), .D(
        memory[132]), .S0(n352), .S1(n350), .Y(n46) );
  MX4X1 U34 ( .A(memory[181]), .B(memory[165]), .C(memory[149]), .D(
        memory[133]), .S0(n352), .S1(n350), .Y(n307) );
  MX4X1 U35 ( .A(memory[182]), .B(memory[166]), .C(memory[150]), .D(
        memory[134]), .S0(n352), .S1(n350), .Y(n311) );
  MX4X1 U36 ( .A(memory[183]), .B(memory[167]), .C(memory[151]), .D(
        memory[135]), .S0(addr[0]), .S1(n350), .Y(n315) );
  MX4X1 U37 ( .A(memory[184]), .B(memory[168]), .C(memory[152]), .D(
        memory[136]), .S0(n353), .S1(n350), .Y(n319) );
  MX4X1 U38 ( .A(memory[185]), .B(memory[169]), .C(memory[153]), .D(
        memory[137]), .S0(n351), .S1(n349), .Y(n323) );
  MX4X1 U39 ( .A(memory[186]), .B(memory[170]), .C(memory[154]), .D(
        memory[138]), .S0(n353), .S1(n350), .Y(n327) );
  MX4X1 U40 ( .A(memory[187]), .B(memory[171]), .C(memory[155]), .D(
        memory[139]), .S0(n353), .S1(addr[1]), .Y(n331) );
  MX4X1 U41 ( .A(memory[188]), .B(memory[172]), .C(memory[156]), .D(
        memory[140]), .S0(n353), .S1(addr[1]), .Y(n335) );
  MX4X1 U42 ( .A(memory[189]), .B(memory[173]), .C(memory[157]), .D(
        memory[141]), .S0(n352), .S1(addr[1]), .Y(n339) );
  MX4X1 U43 ( .A(memory[190]), .B(memory[174]), .C(memory[158]), .D(
        memory[142]), .S0(n353), .S1(addr[1]), .Y(n343) );
  MX4X1 U44 ( .A(memory[191]), .B(memory[175]), .C(memory[159]), .D(
        memory[143]), .S0(addr[0]), .S1(addr[1]), .Y(n347) );
  MX4X1 U45 ( .A(memory[48]), .B(memory[32]), .C(memory[16]), .D(memory[0]), 
        .S0(n351), .S1(n349), .Y(n17) );
  MX4X1 U46 ( .A(memory[49]), .B(memory[33]), .C(memory[17]), .D(memory[1]), 
        .S0(n351), .S1(n349), .Y(n23) );
  MX4X1 U47 ( .A(memory[50]), .B(memory[34]), .C(memory[18]), .D(memory[2]), 
        .S0(n351), .S1(n349), .Y(n30) );
  MX4X1 U48 ( .A(memory[51]), .B(memory[35]), .C(memory[19]), .D(memory[3]), 
        .S0(n351), .S1(n349), .Y(n38) );
  MX4X1 U49 ( .A(memory[52]), .B(memory[36]), .C(memory[20]), .D(memory[4]), 
        .S0(n352), .S1(n350), .Y(n43) );
  MX4X1 U50 ( .A(memory[53]), .B(memory[37]), .C(memory[21]), .D(memory[5]), 
        .S0(n352), .S1(n350), .Y(n305) );
  MX4X1 U51 ( .A(memory[54]), .B(memory[38]), .C(memory[22]), .D(memory[6]), 
        .S0(n352), .S1(n350), .Y(n309) );
  MX4X1 U52 ( .A(memory[55]), .B(memory[39]), .C(memory[23]), .D(memory[7]), 
        .S0(n351), .S1(n349), .Y(n313) );
  MX4X1 U53 ( .A(memory[56]), .B(memory[40]), .C(memory[24]), .D(memory[8]), 
        .S0(n352), .S1(n350), .Y(n317) );
  MX4X1 U54 ( .A(memory[57]), .B(memory[41]), .C(memory[25]), .D(memory[9]), 
        .S0(addr[0]), .S1(n349), .Y(n321) );
  MX4X1 U55 ( .A(memory[58]), .B(memory[42]), .C(memory[26]), .D(memory[10]), 
        .S0(n353), .S1(n349), .Y(n325) );
  MX4X1 U56 ( .A(memory[59]), .B(memory[43]), .C(memory[27]), .D(memory[11]), 
        .S0(n353), .S1(n350), .Y(n329) );
  MX4X1 U57 ( .A(memory[60]), .B(memory[44]), .C(memory[28]), .D(memory[12]), 
        .S0(n353), .S1(n349), .Y(n333) );
  MX4X1 U58 ( .A(memory[61]), .B(memory[45]), .C(memory[29]), .D(memory[13]), 
        .S0(n353), .S1(n349), .Y(n337) );
  MX4X1 U59 ( .A(memory[62]), .B(memory[46]), .C(memory[30]), .D(memory[14]), 
        .S0(n351), .S1(n350), .Y(n341) );
  MX4X1 U60 ( .A(memory[63]), .B(memory[47]), .C(memory[31]), .D(memory[15]), 
        .S0(addr[0]), .S1(addr[1]), .Y(n345) );
  NOR2BX1 U61 ( .AN(N50), .B(n356), .Y(dout[0]) );
  MX4X1 U62 ( .A(n20), .B(n18), .C(n19), .D(n17), .S0(n355), .S1(n354), .Y(N50) );
  MX4X1 U63 ( .A(memory[240]), .B(memory[224]), .C(memory[208]), .D(
        memory[192]), .S0(n353), .S1(addr[1]), .Y(n20) );
  MX4X1 U64 ( .A(memory[112]), .B(memory[96]), .C(memory[80]), .D(memory[64]), 
        .S0(n352), .S1(n349), .Y(n18) );
  NOR2BX1 U65 ( .AN(N49), .B(n356), .Y(dout[1]) );
  MX4X1 U66 ( .A(n28), .B(n25), .C(n27), .D(n23), .S0(n355), .S1(n354), .Y(N49) );
  MX4X1 U67 ( .A(memory[241]), .B(memory[225]), .C(memory[209]), .D(
        memory[193]), .S0(n351), .S1(n349), .Y(n28) );
  MX4X1 U68 ( .A(memory[113]), .B(memory[97]), .C(memory[81]), .D(memory[65]), 
        .S0(n351), .S1(n349), .Y(n25) );
  NOR2BX1 U69 ( .AN(N48), .B(n356), .Y(dout[2]) );
  MX4X1 U70 ( .A(n36), .B(n31), .C(n34), .D(n30), .S0(n355), .S1(n354), .Y(N48) );
  MX4X1 U71 ( .A(memory[242]), .B(memory[226]), .C(memory[210]), .D(
        memory[194]), .S0(n351), .S1(n349), .Y(n36) );
  MX4X1 U72 ( .A(memory[114]), .B(memory[98]), .C(memory[82]), .D(memory[66]), 
        .S0(n351), .S1(n349), .Y(n31) );
  NOR2BX1 U73 ( .AN(N47), .B(n356), .Y(dout[3]) );
  MX4X1 U74 ( .A(n42), .B(n40), .C(n41), .D(n38), .S0(n355), .S1(n354), .Y(N47) );
  MX4X1 U75 ( .A(memory[243]), .B(memory[227]), .C(memory[211]), .D(
        memory[195]), .S0(n351), .S1(n349), .Y(n42) );
  MX4X1 U76 ( .A(memory[115]), .B(memory[99]), .C(memory[83]), .D(memory[67]), 
        .S0(n351), .S1(n349), .Y(n40) );
  NOR2BX1 U77 ( .AN(N46), .B(n356), .Y(dout[4]) );
  MX4X1 U78 ( .A(n304), .B(n44), .C(n46), .D(n43), .S0(n355), .S1(n354), .Y(
        N46) );
  MX4X1 U79 ( .A(memory[244]), .B(memory[228]), .C(memory[212]), .D(
        memory[196]), .S0(n352), .S1(n350), .Y(n304) );
  MX4X1 U80 ( .A(memory[116]), .B(memory[100]), .C(memory[84]), .D(memory[68]), 
        .S0(n352), .S1(n350), .Y(n44) );
  NOR2BX1 U81 ( .AN(N45), .B(n356), .Y(dout[5]) );
  MX4X1 U82 ( .A(n308), .B(n306), .C(n307), .D(n305), .S0(n355), .S1(n354), 
        .Y(N45) );
  MX4X1 U83 ( .A(memory[245]), .B(memory[229]), .C(memory[213]), .D(
        memory[197]), .S0(n352), .S1(n350), .Y(n308) );
  MX4X1 U84 ( .A(memory[117]), .B(memory[101]), .C(memory[85]), .D(memory[69]), 
        .S0(n352), .S1(n350), .Y(n306) );
  NOR2BX1 U85 ( .AN(N44), .B(n356), .Y(dout[6]) );
  MX4X1 U86 ( .A(n312), .B(n310), .C(n311), .D(n309), .S0(n355), .S1(n354), 
        .Y(N44) );
  MX4X1 U87 ( .A(memory[246]), .B(memory[230]), .C(memory[214]), .D(
        memory[198]), .S0(n352), .S1(n350), .Y(n312) );
  MX4X1 U88 ( .A(memory[118]), .B(memory[102]), .C(memory[86]), .D(memory[70]), 
        .S0(n352), .S1(n350), .Y(n310) );
  NOR2BX1 U89 ( .AN(N43), .B(n356), .Y(dout[7]) );
  MX4X1 U90 ( .A(n316), .B(n314), .C(n315), .D(n313), .S0(n355), .S1(n354), 
        .Y(N43) );
  MX4X1 U91 ( .A(memory[247]), .B(memory[231]), .C(memory[215]), .D(
        memory[199]), .S0(n353), .S1(n349), .Y(n316) );
  MX4X1 U92 ( .A(memory[119]), .B(memory[103]), .C(memory[87]), .D(memory[71]), 
        .S0(n353), .S1(n350), .Y(n314) );
  NOR2BX1 U93 ( .AN(N42), .B(n356), .Y(dout[8]) );
  MX4X1 U94 ( .A(n320), .B(n318), .C(n319), .D(n317), .S0(n355), .S1(n354), 
        .Y(N42) );
  MX4X1 U95 ( .A(memory[248]), .B(memory[232]), .C(memory[216]), .D(
        memory[200]), .S0(n351), .S1(n350), .Y(n320) );
  MX4X1 U96 ( .A(memory[120]), .B(memory[104]), .C(memory[88]), .D(memory[72]), 
        .S0(n351), .S1(n349), .Y(n318) );
  NOR2BX1 U97 ( .AN(N41), .B(n356), .Y(dout[9]) );
  MX4X1 U98 ( .A(n324), .B(n322), .C(n323), .D(n321), .S0(n355), .S1(n354), 
        .Y(N41) );
  MX4X1 U99 ( .A(memory[249]), .B(memory[233]), .C(memory[217]), .D(
        memory[201]), .S0(n352), .S1(n349), .Y(n324) );
  MX4X1 U100 ( .A(memory[121]), .B(memory[105]), .C(memory[89]), .D(memory[73]), .S0(n352), .S1(n350), .Y(n322) );
  NOR2BX1 U101 ( .AN(N40), .B(n356), .Y(dout[10]) );
  MX4X1 U102 ( .A(n328), .B(n326), .C(n327), .D(n325), .S0(n355), .S1(n354), 
        .Y(N40) );
  MX4X1 U103 ( .A(memory[250]), .B(memory[234]), .C(memory[218]), .D(
        memory[202]), .S0(n353), .S1(addr[1]), .Y(n328) );
  MX4X1 U104 ( .A(memory[122]), .B(memory[106]), .C(memory[90]), .D(memory[74]), .S0(n353), .S1(addr[1]), .Y(n326) );
  NOR2BX1 U105 ( .AN(N39), .B(n356), .Y(dout[11]) );
  MX4X1 U106 ( .A(n332), .B(n330), .C(n331), .D(n329), .S0(n355), .S1(n354), 
        .Y(N39) );
  MX4X1 U107 ( .A(memory[251]), .B(memory[235]), .C(memory[219]), .D(
        memory[203]), .S0(n353), .S1(addr[1]), .Y(n332) );
  MX4X1 U108 ( .A(memory[123]), .B(memory[107]), .C(memory[91]), .D(memory[75]), .S0(n353), .S1(addr[1]), .Y(n330) );
  NOR2BX1 U109 ( .AN(N38), .B(n356), .Y(dout[12]) );
  MX4X1 U110 ( .A(n336), .B(n334), .C(n335), .D(n333), .S0(n355), .S1(n354), 
        .Y(N38) );
  MX4X1 U111 ( .A(memory[252]), .B(memory[236]), .C(memory[220]), .D(
        memory[204]), .S0(n353), .S1(addr[1]), .Y(n336) );
  MX4X1 U112 ( .A(memory[124]), .B(memory[108]), .C(memory[92]), .D(memory[76]), .S0(n353), .S1(addr[1]), .Y(n334) );
  NOR2BX1 U113 ( .AN(N37), .B(n356), .Y(dout[13]) );
  MX4X1 U114 ( .A(n340), .B(n338), .C(n339), .D(n337), .S0(n355), .S1(n354), 
        .Y(N37) );
  MX4X1 U115 ( .A(memory[253]), .B(memory[237]), .C(memory[221]), .D(
        memory[205]), .S0(addr[0]), .S1(addr[1]), .Y(n340) );
  MX4X1 U116 ( .A(memory[125]), .B(memory[109]), .C(memory[93]), .D(memory[77]), .S0(addr[0]), .S1(addr[1]), .Y(n338) );
  NOR2BX1 U117 ( .AN(N36), .B(n356), .Y(dout[14]) );
  MX4X1 U118 ( .A(n344), .B(n342), .C(n343), .D(n341), .S0(n355), .S1(n354), 
        .Y(N36) );
  MX4X1 U119 ( .A(memory[254]), .B(memory[238]), .C(memory[222]), .D(
        memory[206]), .S0(addr[0]), .S1(addr[1]), .Y(n344) );
  MX4X1 U120 ( .A(memory[126]), .B(memory[110]), .C(memory[94]), .D(memory[78]), .S0(addr[0]), .S1(addr[1]), .Y(n342) );
  NOR2BX1 U121 ( .AN(N35), .B(n356), .Y(dout[15]) );
  MX4X1 U122 ( .A(n348), .B(n346), .C(n347), .D(n345), .S0(n355), .S1(n354), 
        .Y(N35) );
  MX4X1 U123 ( .A(memory[255]), .B(memory[239]), .C(memory[223]), .D(
        memory[207]), .S0(addr[0]), .S1(addr[1]), .Y(n348) );
  MX4X1 U124 ( .A(memory[127]), .B(memory[111]), .C(memory[95]), .D(memory[79]), .S0(addr[0]), .S1(addr[1]), .Y(n346) );
  INVX1 U125 ( .A(addr[1]), .Y(n358) );
  INVX1 U126 ( .A(addr[0]), .Y(n357) );
  NOR2X1 U127 ( .A(n358), .B(addr[2]), .Y(n639) );
  NOR2X1 U128 ( .A(addr[1]), .B(addr[2]), .Y(n638) );
  BUFX3 U129 ( .A(addr[3]), .Y(n355) );
  OAI2BB2X1 U130 ( .B0(n1), .B1(n375), .A0N(memory[0]), .A1N(n1), .Y(n631) );
  OAI2BB2X1 U131 ( .B0(n1), .B1(n374), .A0N(memory[1]), .A1N(n1), .Y(n630) );
  OAI2BB2X1 U132 ( .B0(n1), .B1(n373), .A0N(memory[2]), .A1N(n1), .Y(n629) );
  OAI2BB2X1 U133 ( .B0(n1), .B1(n372), .A0N(memory[3]), .A1N(n1), .Y(n628) );
  OAI2BB2X1 U134 ( .B0(n1), .B1(n371), .A0N(memory[4]), .A1N(n1), .Y(n627) );
  OAI2BB2X1 U135 ( .B0(n1), .B1(n370), .A0N(memory[5]), .A1N(n1), .Y(n626) );
  OAI2BB2X1 U136 ( .B0(n1), .B1(n369), .A0N(memory[6]), .A1N(n1), .Y(n625) );
  OAI2BB2X1 U137 ( .B0(n1), .B1(n368), .A0N(memory[7]), .A1N(n1), .Y(n624) );
  OAI2BB2X1 U138 ( .B0(n1), .B1(n367), .A0N(memory[8]), .A1N(n1), .Y(n623) );
  OAI2BB2X1 U139 ( .B0(n1), .B1(n366), .A0N(memory[9]), .A1N(n1), .Y(n622) );
  OAI2BB2X1 U140 ( .B0(n1), .B1(n365), .A0N(memory[10]), .A1N(n1), .Y(n621) );
  OAI2BB2X1 U141 ( .B0(n1), .B1(n364), .A0N(memory[11]), .A1N(n1), .Y(n620) );
  OAI2BB2X1 U142 ( .B0(n1), .B1(n363), .A0N(memory[12]), .A1N(n1), .Y(n619) );
  OAI2BB2X1 U143 ( .B0(n1), .B1(n362), .A0N(memory[13]), .A1N(n1), .Y(n618) );
  OAI2BB2X1 U144 ( .B0(n1), .B1(n361), .A0N(memory[14]), .A1N(n1), .Y(n617) );
  OAI2BB2X1 U145 ( .B0(n1), .B1(n360), .A0N(memory[15]), .A1N(n1), .Y(n616) );
  OAI2BB2X1 U146 ( .B0(n375), .B1(n2), .A0N(memory[16]), .A1N(n2), .Y(n615) );
  OAI2BB2X1 U147 ( .B0(n374), .B1(n2), .A0N(memory[17]), .A1N(n2), .Y(n614) );
  OAI2BB2X1 U148 ( .B0(n373), .B1(n2), .A0N(memory[18]), .A1N(n2), .Y(n613) );
  OAI2BB2X1 U149 ( .B0(n372), .B1(n2), .A0N(memory[19]), .A1N(n2), .Y(n612) );
  OAI2BB2X1 U150 ( .B0(n371), .B1(n2), .A0N(memory[20]), .A1N(n2), .Y(n611) );
  OAI2BB2X1 U151 ( .B0(n370), .B1(n2), .A0N(memory[21]), .A1N(n2), .Y(n610) );
  OAI2BB2X1 U152 ( .B0(n369), .B1(n2), .A0N(memory[22]), .A1N(n2), .Y(n609) );
  OAI2BB2X1 U153 ( .B0(n368), .B1(n2), .A0N(memory[23]), .A1N(n2), .Y(n608) );
  OAI2BB2X1 U154 ( .B0(n363), .B1(n2), .A0N(memory[28]), .A1N(n2), .Y(n603) );
  OAI2BB2X1 U155 ( .B0(n362), .B1(n2), .A0N(memory[29]), .A1N(n2), .Y(n602) );
  OAI2BB2X1 U156 ( .B0(n361), .B1(n2), .A0N(memory[30]), .A1N(n2), .Y(n601) );
  OAI2BB2X1 U157 ( .B0(n360), .B1(n2), .A0N(memory[31]), .A1N(n2), .Y(n600) );
  OAI2BB2X1 U158 ( .B0(n375), .B1(n3), .A0N(memory[32]), .A1N(n3), .Y(n599) );
  OAI2BB2X1 U159 ( .B0(n374), .B1(n3), .A0N(memory[33]), .A1N(n3), .Y(n598) );
  OAI2BB2X1 U160 ( .B0(n373), .B1(n3), .A0N(memory[34]), .A1N(n3), .Y(n597) );
  OAI2BB2X1 U161 ( .B0(n372), .B1(n3), .A0N(memory[35]), .A1N(n3), .Y(n596) );
  OAI2BB2X1 U162 ( .B0(n371), .B1(n3), .A0N(memory[36]), .A1N(n3), .Y(n595) );
  OAI2BB2X1 U163 ( .B0(n370), .B1(n3), .A0N(memory[37]), .A1N(n3), .Y(n594) );
  OAI2BB2X1 U164 ( .B0(n369), .B1(n3), .A0N(memory[38]), .A1N(n3), .Y(n593) );
  OAI2BB2X1 U165 ( .B0(n368), .B1(n3), .A0N(memory[39]), .A1N(n3), .Y(n592) );
  OAI2BB2X1 U166 ( .B0(n363), .B1(n3), .A0N(memory[44]), .A1N(n3), .Y(n587) );
  OAI2BB2X1 U167 ( .B0(n362), .B1(n3), .A0N(memory[45]), .A1N(n3), .Y(n586) );
  OAI2BB2X1 U168 ( .B0(n361), .B1(n3), .A0N(memory[46]), .A1N(n3), .Y(n585) );
  OAI2BB2X1 U169 ( .B0(n360), .B1(n3), .A0N(memory[47]), .A1N(n3), .Y(n584) );
  OAI2BB2X1 U170 ( .B0(n375), .B1(n4), .A0N(memory[48]), .A1N(n4), .Y(n583) );
  OAI2BB2X1 U171 ( .B0(n374), .B1(n4), .A0N(memory[49]), .A1N(n4), .Y(n582) );
  OAI2BB2X1 U172 ( .B0(n373), .B1(n4), .A0N(memory[50]), .A1N(n4), .Y(n581) );
  OAI2BB2X1 U173 ( .B0(n372), .B1(n4), .A0N(memory[51]), .A1N(n4), .Y(n580) );
  OAI2BB2X1 U174 ( .B0(n371), .B1(n4), .A0N(memory[52]), .A1N(n4), .Y(n579) );
  OAI2BB2X1 U175 ( .B0(n370), .B1(n4), .A0N(memory[53]), .A1N(n4), .Y(n578) );
  OAI2BB2X1 U176 ( .B0(n369), .B1(n4), .A0N(memory[54]), .A1N(n4), .Y(n577) );
  OAI2BB2X1 U177 ( .B0(n368), .B1(n4), .A0N(memory[55]), .A1N(n4), .Y(n576) );
  OAI2BB2X1 U178 ( .B0(n363), .B1(n4), .A0N(memory[60]), .A1N(n4), .Y(n571) );
  OAI2BB2X1 U179 ( .B0(n362), .B1(n4), .A0N(memory[61]), .A1N(n4), .Y(n570) );
  OAI2BB2X1 U180 ( .B0(n361), .B1(n4), .A0N(memory[62]), .A1N(n4), .Y(n569) );
  OAI2BB2X1 U181 ( .B0(n360), .B1(n4), .A0N(memory[63]), .A1N(n4), .Y(n568) );
  OAI2BB2X1 U182 ( .B0(n375), .B1(n5), .A0N(memory[64]), .A1N(n5), .Y(n567) );
  OAI2BB2X1 U183 ( .B0(n374), .B1(n5), .A0N(memory[65]), .A1N(n5), .Y(n566) );
  OAI2BB2X1 U184 ( .B0(n373), .B1(n5), .A0N(memory[66]), .A1N(n5), .Y(n565) );
  OAI2BB2X1 U185 ( .B0(n372), .B1(n5), .A0N(memory[67]), .A1N(n5), .Y(n564) );
  OAI2BB2X1 U186 ( .B0(n371), .B1(n5), .A0N(memory[68]), .A1N(n5), .Y(n563) );
  OAI2BB2X1 U187 ( .B0(n370), .B1(n5), .A0N(memory[69]), .A1N(n5), .Y(n562) );
  OAI2BB2X1 U188 ( .B0(n369), .B1(n5), .A0N(memory[70]), .A1N(n5), .Y(n561) );
  OAI2BB2X1 U189 ( .B0(n368), .B1(n5), .A0N(memory[71]), .A1N(n5), .Y(n560) );
  OAI2BB2X1 U190 ( .B0(n363), .B1(n5), .A0N(memory[76]), .A1N(n5), .Y(n555) );
  OAI2BB2X1 U191 ( .B0(n362), .B1(n5), .A0N(memory[77]), .A1N(n5), .Y(n554) );
  OAI2BB2X1 U192 ( .B0(n361), .B1(n5), .A0N(memory[78]), .A1N(n5), .Y(n553) );
  OAI2BB2X1 U193 ( .B0(n360), .B1(n5), .A0N(memory[79]), .A1N(n5), .Y(n552) );
  OAI2BB2X1 U194 ( .B0(n375), .B1(n6), .A0N(memory[80]), .A1N(n6), .Y(n551) );
  OAI2BB2X1 U195 ( .B0(n374), .B1(n6), .A0N(memory[81]), .A1N(n6), .Y(n550) );
  OAI2BB2X1 U196 ( .B0(n373), .B1(n6), .A0N(memory[82]), .A1N(n6), .Y(n549) );
  OAI2BB2X1 U197 ( .B0(n372), .B1(n6), .A0N(memory[83]), .A1N(n6), .Y(n548) );
  OAI2BB2X1 U198 ( .B0(n371), .B1(n6), .A0N(memory[84]), .A1N(n6), .Y(n547) );
  OAI2BB2X1 U199 ( .B0(n370), .B1(n6), .A0N(memory[85]), .A1N(n6), .Y(n546) );
  OAI2BB2X1 U200 ( .B0(n369), .B1(n6), .A0N(memory[86]), .A1N(n6), .Y(n545) );
  OAI2BB2X1 U201 ( .B0(n368), .B1(n6), .A0N(memory[87]), .A1N(n6), .Y(n544) );
  OAI2BB2X1 U202 ( .B0(n363), .B1(n6), .A0N(memory[92]), .A1N(n6), .Y(n539) );
  OAI2BB2X1 U203 ( .B0(n362), .B1(n6), .A0N(memory[93]), .A1N(n6), .Y(n538) );
  OAI2BB2X1 U204 ( .B0(n361), .B1(n6), .A0N(memory[94]), .A1N(n6), .Y(n537) );
  OAI2BB2X1 U205 ( .B0(n360), .B1(n6), .A0N(memory[95]), .A1N(n6), .Y(n536) );
  OAI2BB2X1 U206 ( .B0(n375), .B1(n7), .A0N(memory[96]), .A1N(n7), .Y(n535) );
  OAI2BB2X1 U207 ( .B0(n374), .B1(n7), .A0N(memory[97]), .A1N(n7), .Y(n534) );
  OAI2BB2X1 U208 ( .B0(n373), .B1(n7), .A0N(memory[98]), .A1N(n7), .Y(n533) );
  OAI2BB2X1 U209 ( .B0(n372), .B1(n7), .A0N(memory[99]), .A1N(n7), .Y(n532) );
  OAI2BB2X1 U210 ( .B0(n371), .B1(n7), .A0N(memory[100]), .A1N(n7), .Y(n531)
         );
  OAI2BB2X1 U211 ( .B0(n370), .B1(n7), .A0N(memory[101]), .A1N(n7), .Y(n530)
         );
  OAI2BB2X1 U212 ( .B0(n369), .B1(n7), .A0N(memory[102]), .A1N(n7), .Y(n529)
         );
  OAI2BB2X1 U213 ( .B0(n368), .B1(n7), .A0N(memory[103]), .A1N(n7), .Y(n528)
         );
  OAI2BB2X1 U214 ( .B0(n363), .B1(n7), .A0N(memory[108]), .A1N(n7), .Y(n523)
         );
  OAI2BB2X1 U215 ( .B0(n362), .B1(n7), .A0N(memory[109]), .A1N(n7), .Y(n522)
         );
  OAI2BB2X1 U216 ( .B0(n361), .B1(n7), .A0N(memory[110]), .A1N(n7), .Y(n521)
         );
  OAI2BB2X1 U217 ( .B0(n360), .B1(n7), .A0N(memory[111]), .A1N(n7), .Y(n520)
         );
  OAI2BB2X1 U218 ( .B0(n375), .B1(n8), .A0N(memory[112]), .A1N(n8), .Y(n519)
         );
  OAI2BB2X1 U219 ( .B0(n374), .B1(n8), .A0N(memory[113]), .A1N(n8), .Y(n518)
         );
  OAI2BB2X1 U220 ( .B0(n373), .B1(n8), .A0N(memory[114]), .A1N(n8), .Y(n517)
         );
  OAI2BB2X1 U221 ( .B0(n372), .B1(n8), .A0N(memory[115]), .A1N(n8), .Y(n516)
         );
  OAI2BB2X1 U222 ( .B0(n371), .B1(n8), .A0N(memory[116]), .A1N(n8), .Y(n515)
         );
  OAI2BB2X1 U223 ( .B0(n370), .B1(n8), .A0N(memory[117]), .A1N(n8), .Y(n514)
         );
  OAI2BB2X1 U224 ( .B0(n369), .B1(n8), .A0N(memory[118]), .A1N(n8), .Y(n513)
         );
  OAI2BB2X1 U225 ( .B0(n368), .B1(n8), .A0N(memory[119]), .A1N(n8), .Y(n512)
         );
  OAI2BB2X1 U226 ( .B0(n363), .B1(n8), .A0N(memory[124]), .A1N(n8), .Y(n507)
         );
  OAI2BB2X1 U227 ( .B0(n362), .B1(n8), .A0N(memory[125]), .A1N(n8), .Y(n506)
         );
  OAI2BB2X1 U228 ( .B0(n361), .B1(n8), .A0N(memory[126]), .A1N(n8), .Y(n505)
         );
  OAI2BB2X1 U229 ( .B0(n360), .B1(n8), .A0N(memory[127]), .A1N(n8), .Y(n504)
         );
  OAI2BB2X1 U230 ( .B0(n375), .B1(n9), .A0N(memory[128]), .A1N(n9), .Y(n503)
         );
  OAI2BB2X1 U231 ( .B0(n374), .B1(n9), .A0N(memory[129]), .A1N(n9), .Y(n502)
         );
  OAI2BB2X1 U232 ( .B0(n373), .B1(n9), .A0N(memory[130]), .A1N(n9), .Y(n501)
         );
  OAI2BB2X1 U233 ( .B0(n372), .B1(n9), .A0N(memory[131]), .A1N(n9), .Y(n500)
         );
  OAI2BB2X1 U234 ( .B0(n371), .B1(n9), .A0N(memory[132]), .A1N(n9), .Y(n499)
         );
  OAI2BB2X1 U235 ( .B0(n370), .B1(n9), .A0N(memory[133]), .A1N(n9), .Y(n498)
         );
  OAI2BB2X1 U236 ( .B0(n369), .B1(n9), .A0N(memory[134]), .A1N(n9), .Y(n497)
         );
  OAI2BB2X1 U237 ( .B0(n368), .B1(n9), .A0N(memory[135]), .A1N(n9), .Y(n496)
         );
  OAI2BB2X1 U238 ( .B0(n363), .B1(n9), .A0N(memory[140]), .A1N(n9), .Y(n491)
         );
  OAI2BB2X1 U239 ( .B0(n362), .B1(n9), .A0N(memory[141]), .A1N(n9), .Y(n490)
         );
  OAI2BB2X1 U240 ( .B0(n361), .B1(n9), .A0N(memory[142]), .A1N(n9), .Y(n489)
         );
  OAI2BB2X1 U241 ( .B0(n360), .B1(n9), .A0N(memory[143]), .A1N(n9), .Y(n488)
         );
  OAI2BB2X1 U242 ( .B0(n375), .B1(n10), .A0N(memory[144]), .A1N(n10), .Y(n487)
         );
  OAI2BB2X1 U243 ( .B0(n374), .B1(n10), .A0N(memory[145]), .A1N(n10), .Y(n486)
         );
  OAI2BB2X1 U244 ( .B0(n373), .B1(n10), .A0N(memory[146]), .A1N(n10), .Y(n485)
         );
  OAI2BB2X1 U245 ( .B0(n372), .B1(n10), .A0N(memory[147]), .A1N(n10), .Y(n484)
         );
  OAI2BB2X1 U246 ( .B0(n371), .B1(n10), .A0N(memory[148]), .A1N(n10), .Y(n483)
         );
  OAI2BB2X1 U247 ( .B0(n370), .B1(n10), .A0N(memory[149]), .A1N(n10), .Y(n482)
         );
  OAI2BB2X1 U248 ( .B0(n369), .B1(n10), .A0N(memory[150]), .A1N(n10), .Y(n481)
         );
  OAI2BB2X1 U249 ( .B0(n368), .B1(n10), .A0N(memory[151]), .A1N(n10), .Y(n480)
         );
  OAI2BB2X1 U250 ( .B0(n363), .B1(n10), .A0N(memory[156]), .A1N(n10), .Y(n475)
         );
  OAI2BB2X1 U251 ( .B0(n362), .B1(n10), .A0N(memory[157]), .A1N(n10), .Y(n474)
         );
  OAI2BB2X1 U252 ( .B0(n361), .B1(n10), .A0N(memory[158]), .A1N(n10), .Y(n473)
         );
  OAI2BB2X1 U253 ( .B0(n360), .B1(n10), .A0N(memory[159]), .A1N(n10), .Y(n472)
         );
  OAI2BB2X1 U254 ( .B0(n375), .B1(n11), .A0N(memory[160]), .A1N(n11), .Y(n471)
         );
  OAI2BB2X1 U255 ( .B0(n374), .B1(n11), .A0N(memory[161]), .A1N(n11), .Y(n470)
         );
  OAI2BB2X1 U256 ( .B0(n373), .B1(n11), .A0N(memory[162]), .A1N(n11), .Y(n469)
         );
  OAI2BB2X1 U257 ( .B0(n372), .B1(n11), .A0N(memory[163]), .A1N(n11), .Y(n468)
         );
  OAI2BB2X1 U258 ( .B0(n371), .B1(n11), .A0N(memory[164]), .A1N(n11), .Y(n467)
         );
  OAI2BB2X1 U259 ( .B0(n370), .B1(n11), .A0N(memory[165]), .A1N(n11), .Y(n466)
         );
  OAI2BB2X1 U260 ( .B0(n369), .B1(n11), .A0N(memory[166]), .A1N(n11), .Y(n465)
         );
  OAI2BB2X1 U261 ( .B0(n368), .B1(n11), .A0N(memory[167]), .A1N(n11), .Y(n464)
         );
  OAI2BB2X1 U262 ( .B0(n363), .B1(n11), .A0N(memory[172]), .A1N(n11), .Y(n459)
         );
  OAI2BB2X1 U263 ( .B0(n362), .B1(n11), .A0N(memory[173]), .A1N(n11), .Y(n458)
         );
  OAI2BB2X1 U264 ( .B0(n361), .B1(n11), .A0N(memory[174]), .A1N(n11), .Y(n457)
         );
  OAI2BB2X1 U265 ( .B0(n360), .B1(n11), .A0N(memory[175]), .A1N(n11), .Y(n456)
         );
  OAI2BB2X1 U266 ( .B0(n375), .B1(n12), .A0N(memory[176]), .A1N(n12), .Y(n455)
         );
  OAI2BB2X1 U267 ( .B0(n374), .B1(n12), .A0N(memory[177]), .A1N(n12), .Y(n454)
         );
  OAI2BB2X1 U268 ( .B0(n373), .B1(n12), .A0N(memory[178]), .A1N(n12), .Y(n453)
         );
  OAI2BB2X1 U269 ( .B0(n372), .B1(n12), .A0N(memory[179]), .A1N(n12), .Y(n452)
         );
  OAI2BB2X1 U270 ( .B0(n371), .B1(n12), .A0N(memory[180]), .A1N(n12), .Y(n451)
         );
  OAI2BB2X1 U271 ( .B0(n370), .B1(n12), .A0N(memory[181]), .A1N(n12), .Y(n450)
         );
  OAI2BB2X1 U272 ( .B0(n369), .B1(n12), .A0N(memory[182]), .A1N(n12), .Y(n449)
         );
  OAI2BB2X1 U273 ( .B0(n368), .B1(n12), .A0N(memory[183]), .A1N(n12), .Y(n448)
         );
  OAI2BB2X1 U274 ( .B0(n363), .B1(n12), .A0N(memory[188]), .A1N(n12), .Y(n443)
         );
  OAI2BB2X1 U275 ( .B0(n362), .B1(n12), .A0N(memory[189]), .A1N(n12), .Y(n442)
         );
  OAI2BB2X1 U276 ( .B0(n361), .B1(n12), .A0N(memory[190]), .A1N(n12), .Y(n441)
         );
  OAI2BB2X1 U277 ( .B0(n360), .B1(n12), .A0N(memory[191]), .A1N(n12), .Y(n440)
         );
  OAI2BB2X1 U278 ( .B0(n375), .B1(n13), .A0N(memory[192]), .A1N(n13), .Y(n439)
         );
  OAI2BB2X1 U279 ( .B0(n374), .B1(n13), .A0N(memory[193]), .A1N(n13), .Y(n438)
         );
  OAI2BB2X1 U280 ( .B0(n373), .B1(n13), .A0N(memory[194]), .A1N(n13), .Y(n437)
         );
  OAI2BB2X1 U281 ( .B0(n372), .B1(n13), .A0N(memory[195]), .A1N(n13), .Y(n436)
         );
  OAI2BB2X1 U282 ( .B0(n371), .B1(n13), .A0N(memory[196]), .A1N(n13), .Y(n435)
         );
  OAI2BB2X1 U283 ( .B0(n370), .B1(n13), .A0N(memory[197]), .A1N(n13), .Y(n434)
         );
  OAI2BB2X1 U284 ( .B0(n369), .B1(n13), .A0N(memory[198]), .A1N(n13), .Y(n433)
         );
  OAI2BB2X1 U285 ( .B0(n368), .B1(n13), .A0N(memory[199]), .A1N(n13), .Y(n432)
         );
  OAI2BB2X1 U286 ( .B0(n363), .B1(n13), .A0N(memory[204]), .A1N(n13), .Y(n427)
         );
  OAI2BB2X1 U287 ( .B0(n362), .B1(n13), .A0N(memory[205]), .A1N(n13), .Y(n426)
         );
  OAI2BB2X1 U288 ( .B0(n361), .B1(n13), .A0N(memory[206]), .A1N(n13), .Y(n425)
         );
  OAI2BB2X1 U289 ( .B0(n360), .B1(n13), .A0N(memory[207]), .A1N(n13), .Y(n424)
         );
  OAI2BB2X1 U290 ( .B0(n375), .B1(n14), .A0N(memory[208]), .A1N(n14), .Y(n423)
         );
  OAI2BB2X1 U291 ( .B0(n374), .B1(n14), .A0N(memory[209]), .A1N(n14), .Y(n422)
         );
  OAI2BB2X1 U292 ( .B0(n373), .B1(n14), .A0N(memory[210]), .A1N(n14), .Y(n421)
         );
  OAI2BB2X1 U293 ( .B0(n372), .B1(n14), .A0N(memory[211]), .A1N(n14), .Y(n420)
         );
  OAI2BB2X1 U294 ( .B0(n371), .B1(n14), .A0N(memory[212]), .A1N(n14), .Y(n419)
         );
  OAI2BB2X1 U295 ( .B0(n370), .B1(n14), .A0N(memory[213]), .A1N(n14), .Y(n418)
         );
  OAI2BB2X1 U296 ( .B0(n369), .B1(n14), .A0N(memory[214]), .A1N(n14), .Y(n417)
         );
  OAI2BB2X1 U297 ( .B0(n368), .B1(n14), .A0N(memory[215]), .A1N(n14), .Y(n416)
         );
  OAI2BB2X1 U298 ( .B0(n363), .B1(n14), .A0N(memory[220]), .A1N(n14), .Y(n411)
         );
  OAI2BB2X1 U299 ( .B0(n362), .B1(n14), .A0N(memory[221]), .A1N(n14), .Y(n410)
         );
  OAI2BB2X1 U300 ( .B0(n361), .B1(n14), .A0N(memory[222]), .A1N(n14), .Y(n409)
         );
  OAI2BB2X1 U301 ( .B0(n360), .B1(n14), .A0N(memory[223]), .A1N(n14), .Y(n408)
         );
  OAI2BB2X1 U302 ( .B0(n375), .B1(n15), .A0N(memory[224]), .A1N(n15), .Y(n407)
         );
  OAI2BB2X1 U303 ( .B0(n374), .B1(n15), .A0N(memory[225]), .A1N(n15), .Y(n406)
         );
  OAI2BB2X1 U304 ( .B0(n373), .B1(n15), .A0N(memory[226]), .A1N(n15), .Y(n405)
         );
  OAI2BB2X1 U305 ( .B0(n372), .B1(n15), .A0N(memory[227]), .A1N(n15), .Y(n404)
         );
  OAI2BB2X1 U306 ( .B0(n371), .B1(n15), .A0N(memory[228]), .A1N(n15), .Y(n403)
         );
  OAI2BB2X1 U307 ( .B0(n370), .B1(n15), .A0N(memory[229]), .A1N(n15), .Y(n402)
         );
  OAI2BB2X1 U308 ( .B0(n369), .B1(n15), .A0N(memory[230]), .A1N(n15), .Y(n401)
         );
  OAI2BB2X1 U309 ( .B0(n368), .B1(n15), .A0N(memory[231]), .A1N(n15), .Y(n400)
         );
  OAI2BB2X1 U310 ( .B0(n363), .B1(n15), .A0N(memory[236]), .A1N(n15), .Y(n395)
         );
  OAI2BB2X1 U311 ( .B0(n362), .B1(n15), .A0N(memory[237]), .A1N(n15), .Y(n394)
         );
  OAI2BB2X1 U312 ( .B0(n361), .B1(n15), .A0N(memory[238]), .A1N(n15), .Y(n393)
         );
  OAI2BB2X1 U313 ( .B0(n360), .B1(n15), .A0N(memory[239]), .A1N(n15), .Y(n392)
         );
  OAI2BB2X1 U314 ( .B0(n375), .B1(n16), .A0N(memory[240]), .A1N(n16), .Y(n391)
         );
  OAI2BB2X1 U315 ( .B0(n374), .B1(n16), .A0N(memory[241]), .A1N(n16), .Y(n390)
         );
  OAI2BB2X1 U316 ( .B0(n373), .B1(n16), .A0N(memory[242]), .A1N(n16), .Y(n389)
         );
  OAI2BB2X1 U317 ( .B0(n372), .B1(n16), .A0N(memory[243]), .A1N(n16), .Y(n388)
         );
  OAI2BB2X1 U318 ( .B0(n371), .B1(n16), .A0N(memory[244]), .A1N(n16), .Y(n387)
         );
  OAI2BB2X1 U319 ( .B0(n370), .B1(n16), .A0N(memory[245]), .A1N(n16), .Y(n386)
         );
  OAI2BB2X1 U320 ( .B0(n369), .B1(n16), .A0N(memory[246]), .A1N(n16), .Y(n385)
         );
  OAI2BB2X1 U321 ( .B0(n368), .B1(n16), .A0N(memory[247]), .A1N(n16), .Y(n384)
         );
  OAI2BB2X1 U322 ( .B0(n363), .B1(n16), .A0N(memory[252]), .A1N(n16), .Y(n379)
         );
  OAI2BB2X1 U323 ( .B0(n362), .B1(n16), .A0N(memory[253]), .A1N(n16), .Y(n378)
         );
  OAI2BB2X1 U324 ( .B0(n361), .B1(n16), .A0N(memory[254]), .A1N(n16), .Y(n377)
         );
  OAI2BB2X1 U325 ( .B0(n360), .B1(n16), .A0N(memory[255]), .A1N(n16), .Y(n376)
         );
  OAI2BB2X1 U326 ( .B0(n367), .B1(n2), .A0N(memory[24]), .A1N(n2), .Y(n607) );
  OAI2BB2X1 U327 ( .B0(n366), .B1(n2), .A0N(memory[25]), .A1N(n2), .Y(n606) );
  OAI2BB2X1 U328 ( .B0(n365), .B1(n2), .A0N(memory[26]), .A1N(n2), .Y(n605) );
  OAI2BB2X1 U329 ( .B0(n364), .B1(n2), .A0N(memory[27]), .A1N(n2), .Y(n604) );
  OAI2BB2X1 U330 ( .B0(n367), .B1(n3), .A0N(memory[40]), .A1N(n3), .Y(n591) );
  OAI2BB2X1 U331 ( .B0(n366), .B1(n3), .A0N(memory[41]), .A1N(n3), .Y(n590) );
  OAI2BB2X1 U332 ( .B0(n365), .B1(n3), .A0N(memory[42]), .A1N(n3), .Y(n589) );
  OAI2BB2X1 U333 ( .B0(n364), .B1(n3), .A0N(memory[43]), .A1N(n3), .Y(n588) );
  OAI2BB2X1 U334 ( .B0(n367), .B1(n4), .A0N(memory[56]), .A1N(n4), .Y(n575) );
  OAI2BB2X1 U335 ( .B0(n366), .B1(n4), .A0N(memory[57]), .A1N(n4), .Y(n574) );
  OAI2BB2X1 U336 ( .B0(n365), .B1(n4), .A0N(memory[58]), .A1N(n4), .Y(n573) );
  OAI2BB2X1 U337 ( .B0(n364), .B1(n4), .A0N(memory[59]), .A1N(n4), .Y(n572) );
  OAI2BB2X1 U338 ( .B0(n367), .B1(n5), .A0N(memory[72]), .A1N(n5), .Y(n559) );
  OAI2BB2X1 U339 ( .B0(n366), .B1(n5), .A0N(memory[73]), .A1N(n5), .Y(n558) );
  OAI2BB2X1 U340 ( .B0(n365), .B1(n5), .A0N(memory[74]), .A1N(n5), .Y(n557) );
  OAI2BB2X1 U341 ( .B0(n364), .B1(n5), .A0N(memory[75]), .A1N(n5), .Y(n556) );
  OAI2BB2X1 U342 ( .B0(n367), .B1(n6), .A0N(memory[88]), .A1N(n6), .Y(n543) );
  OAI2BB2X1 U343 ( .B0(n366), .B1(n6), .A0N(memory[89]), .A1N(n6), .Y(n542) );
  OAI2BB2X1 U344 ( .B0(n365), .B1(n6), .A0N(memory[90]), .A1N(n6), .Y(n541) );
  OAI2BB2X1 U345 ( .B0(n364), .B1(n6), .A0N(memory[91]), .A1N(n6), .Y(n540) );
  OAI2BB2X1 U346 ( .B0(n367), .B1(n7), .A0N(memory[104]), .A1N(n7), .Y(n527)
         );
  OAI2BB2X1 U347 ( .B0(n366), .B1(n7), .A0N(memory[105]), .A1N(n7), .Y(n526)
         );
  OAI2BB2X1 U348 ( .B0(n365), .B1(n7), .A0N(memory[106]), .A1N(n7), .Y(n525)
         );
  OAI2BB2X1 U349 ( .B0(n364), .B1(n7), .A0N(memory[107]), .A1N(n7), .Y(n524)
         );
  OAI2BB2X1 U350 ( .B0(n367), .B1(n8), .A0N(memory[120]), .A1N(n8), .Y(n511)
         );
  OAI2BB2X1 U351 ( .B0(n366), .B1(n8), .A0N(memory[121]), .A1N(n8), .Y(n510)
         );
  OAI2BB2X1 U352 ( .B0(n365), .B1(n8), .A0N(memory[122]), .A1N(n8), .Y(n509)
         );
  OAI2BB2X1 U353 ( .B0(n364), .B1(n8), .A0N(memory[123]), .A1N(n8), .Y(n508)
         );
  OAI2BB2X1 U354 ( .B0(n367), .B1(n9), .A0N(memory[136]), .A1N(n9), .Y(n495)
         );
  OAI2BB2X1 U355 ( .B0(n366), .B1(n9), .A0N(memory[137]), .A1N(n9), .Y(n494)
         );
  OAI2BB2X1 U356 ( .B0(n365), .B1(n9), .A0N(memory[138]), .A1N(n9), .Y(n493)
         );
  OAI2BB2X1 U357 ( .B0(n364), .B1(n9), .A0N(memory[139]), .A1N(n9), .Y(n492)
         );
  OAI2BB2X1 U358 ( .B0(n367), .B1(n10), .A0N(memory[152]), .A1N(n10), .Y(n479)
         );
  OAI2BB2X1 U359 ( .B0(n366), .B1(n10), .A0N(memory[153]), .A1N(n10), .Y(n478)
         );
  OAI2BB2X1 U360 ( .B0(n365), .B1(n10), .A0N(memory[154]), .A1N(n10), .Y(n477)
         );
  OAI2BB2X1 U361 ( .B0(n364), .B1(n10), .A0N(memory[155]), .A1N(n10), .Y(n476)
         );
  OAI2BB2X1 U362 ( .B0(n367), .B1(n11), .A0N(memory[168]), .A1N(n11), .Y(n463)
         );
  OAI2BB2X1 U363 ( .B0(n366), .B1(n11), .A0N(memory[169]), .A1N(n11), .Y(n462)
         );
  OAI2BB2X1 U364 ( .B0(n365), .B1(n11), .A0N(memory[170]), .A1N(n11), .Y(n461)
         );
  OAI2BB2X1 U365 ( .B0(n364), .B1(n11), .A0N(memory[171]), .A1N(n11), .Y(n460)
         );
  OAI2BB2X1 U366 ( .B0(n367), .B1(n12), .A0N(memory[184]), .A1N(n12), .Y(n447)
         );
  OAI2BB2X1 U367 ( .B0(n366), .B1(n12), .A0N(memory[185]), .A1N(n12), .Y(n446)
         );
  OAI2BB2X1 U368 ( .B0(n365), .B1(n12), .A0N(memory[186]), .A1N(n12), .Y(n445)
         );
  OAI2BB2X1 U369 ( .B0(n364), .B1(n12), .A0N(memory[187]), .A1N(n12), .Y(n444)
         );
  OAI2BB2X1 U370 ( .B0(n367), .B1(n13), .A0N(memory[200]), .A1N(n13), .Y(n431)
         );
  OAI2BB2X1 U371 ( .B0(n366), .B1(n13), .A0N(memory[201]), .A1N(n13), .Y(n430)
         );
  OAI2BB2X1 U372 ( .B0(n365), .B1(n13), .A0N(memory[202]), .A1N(n13), .Y(n429)
         );
  OAI2BB2X1 U373 ( .B0(n364), .B1(n13), .A0N(memory[203]), .A1N(n13), .Y(n428)
         );
  OAI2BB2X1 U374 ( .B0(n367), .B1(n14), .A0N(memory[216]), .A1N(n14), .Y(n415)
         );
  OAI2BB2X1 U375 ( .B0(n366), .B1(n14), .A0N(memory[217]), .A1N(n14), .Y(n414)
         );
  OAI2BB2X1 U376 ( .B0(n365), .B1(n14), .A0N(memory[218]), .A1N(n14), .Y(n413)
         );
  OAI2BB2X1 U377 ( .B0(n364), .B1(n14), .A0N(memory[219]), .A1N(n14), .Y(n412)
         );
  OAI2BB2X1 U378 ( .B0(n367), .B1(n15), .A0N(memory[232]), .A1N(n15), .Y(n399)
         );
  OAI2BB2X1 U379 ( .B0(n366), .B1(n15), .A0N(memory[233]), .A1N(n15), .Y(n398)
         );
  OAI2BB2X1 U380 ( .B0(n365), .B1(n15), .A0N(memory[234]), .A1N(n15), .Y(n397)
         );
  OAI2BB2X1 U381 ( .B0(n364), .B1(n15), .A0N(memory[235]), .A1N(n15), .Y(n396)
         );
  OAI2BB2X1 U382 ( .B0(n367), .B1(n16), .A0N(memory[248]), .A1N(n16), .Y(n383)
         );
  OAI2BB2X1 U383 ( .B0(n366), .B1(n16), .A0N(memory[249]), .A1N(n16), .Y(n382)
         );
  OAI2BB2X1 U384 ( .B0(n365), .B1(n16), .A0N(memory[250]), .A1N(n16), .Y(n381)
         );
  OAI2BB2X1 U385 ( .B0(n364), .B1(n16), .A0N(memory[251]), .A1N(n16), .Y(n380)
         );
  BUFX3 U386 ( .A(n632), .Y(n356) );
  NAND2BX1 U387 ( .AN(wr_rd), .B(en), .Y(n632) );
  NOR2BX1 U388 ( .AN(n636), .B(addr[3]), .Y(n633) );
  BUFX3 U389 ( .A(addr[2]), .Y(n354) );
  INVX1 U390 ( .A(addr[2]), .Y(n359) );
  AND2X2 U391 ( .A(wr_rd), .B(en), .Y(n636) );
  AND2X2 U392 ( .A(addr[3]), .B(n636), .Y(n637) );
  INVX1 U393 ( .A(din[0]), .Y(n375) );
  INVX1 U394 ( .A(din[1]), .Y(n374) );
  INVX1 U395 ( .A(din[2]), .Y(n373) );
  INVX1 U396 ( .A(din[3]), .Y(n372) );
  INVX1 U397 ( .A(din[4]), .Y(n371) );
  INVX1 U398 ( .A(din[5]), .Y(n370) );
  INVX1 U399 ( .A(din[6]), .Y(n369) );
  INVX1 U400 ( .A(din[7]), .Y(n368) );
  INVX1 U401 ( .A(din[8]), .Y(n367) );
  INVX1 U402 ( .A(din[9]), .Y(n366) );
  INVX1 U403 ( .A(din[10]), .Y(n365) );
  INVX1 U404 ( .A(din[11]), .Y(n364) );
  INVX1 U405 ( .A(din[12]), .Y(n363) );
  INVX1 U406 ( .A(din[13]), .Y(n362) );
  INVX1 U407 ( .A(din[14]), .Y(n361) );
  INVX1 U408 ( .A(din[15]), .Y(n360) );
endmodule


module s2p_1 ( clk, rstn, start, mode, din, dout, s2p_ready, mode_out );
  input [1:0] mode;
  input [15:0] din;
  output [255:0] dout;
  output [1:0] mode_out;
  input clk, rstn, start;
  output s2p_ready;
  wire   N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43,
         N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57,
         N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71,
         N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85,
         N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99,
         N100, N101, N102, N103, N104, N105, N106, N107, N108, N109, N110,
         N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121,
         N122, N123, N124, N125, N126, N127, N128, N129, N131, N132, N133,
         N134, N135, N136, N137, N138, N139, N140, N141, N142, N143, N144,
         N145, N146, N147, N148, N149, N150, N151, N152, N153, N154, N155,
         N156, N157, N158, N159, N160, N161, N162, N163, N164, N165, N166,
         N167, N168, N169, N170, N171, N172, N173, N174, N175, N176, N177,
         N178, N179, N180, N181, N182, N183, N184, N185, N186, N187, N188,
         N189, N190, N191, N192, N193, N194, N195, N196, N197, N198, N199,
         N200, N201, N202, N203, N204, N205, N206, N207, N208, N209, N210,
         N211, N212, N213, N214, N215, N216, N217, N218, N219, N220, N221,
         N222, N223, N224, N225, N226, N227, N228, N229, N231, N232, N233,
         N234, N235, N236, N237, N238, N239, N240, N241, N242, N243, N244,
         N245, N246, N247, N248, N249, N250, N251, N252, N253, N254, N255,
         N256, N257, N258, N259, N260, N261, N262, N263, N264, N265, N266,
         N267, N268, N269, N270, N271, N272, N273, N274, N275, N276, N277,
         N278, N279, N280, N281, N282, N283, N284, N285, N286, N287, N288,
         N302, N303, N304, N1114, N1115, N1116, N1117, N1118, N1119, n1, n2,
         n3, n4, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n732, n738,
         n739, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
         n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
         n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
         n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
         n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
         n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
         n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
         n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
         n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
         n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
         n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
         n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
         n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
         n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
         n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
         n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427,
         n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437,
         n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
         n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
         n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
         n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
         n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487,
         n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497,
         n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507,
         n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517,
         n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527,
         n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537,
         n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547,
         n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557,
         n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567,
         n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577,
         n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587,
         n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597,
         n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607,
         n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617,
         n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627,
         n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637,
         n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647,
         n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657,
         n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667,
         n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677,
         n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687,
         n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
         n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707,
         n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
         n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727,
         n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735;
  wire   [1:0] mode_reg;
  wire   [63:0] dout4_reg;
  wire   [127:0] dout8_reg;
  wire   [255:0] dout16_reg;
  wire   [4:0] count;
  wire   [4:2] r71_carry;

  OAI2BB2X4 U3 ( .B0(n349), .B1(n351), .A0N(n351), .A1N(mode_out[0]), .Y(
        mode_out[0]) );
  OAI2BB2X4 U4 ( .B0(n351), .B1(n348), .A0N(n351), .A1N(mode_out[1]), .Y(
        mode_out[1]) );
  TLATX1 dout_reg_16_ ( .G(n327), .D(N47), .Q(dout[16]) );
  TLATX1 dout_reg_111_ ( .G(n319), .D(N143), .Q(dout[111]) );
  TLATX1 dout_reg_79_ ( .G(n318), .D(N110), .Q(dout[79]) );
  TLATX1 dout_reg_47_ ( .G(n328), .D(N78), .Q(dout[47]) );
  TLATX1 dout_reg_31_ ( .G(n326), .D(N62), .Q(dout[31]) );
  TLATX1 dout_reg_110_ ( .G(N30), .D(N142), .Q(dout[110]) );
  TLATX1 dout_reg_78_ ( .G(n318), .D(N109), .Q(dout[78]) );
  TLATX1 dout_reg_46_ ( .G(n322), .D(N77), .Q(dout[46]) );
  TLATX1 dout_reg_30_ ( .G(n322), .D(N61), .Q(dout[30]) );
  TLATX1 dout_reg_109_ ( .G(n326), .D(N141), .Q(dout[109]) );
  TLATX1 dout_reg_77_ ( .G(N30), .D(N108), .Q(dout[77]) );
  TLATX1 dout_reg_45_ ( .G(n318), .D(N76), .Q(dout[45]) );
  TLATX1 dout_reg_29_ ( .G(n328), .D(N60), .Q(dout[29]) );
  TLATX1 dout_reg_108_ ( .G(n330), .D(N140), .Q(dout[108]) );
  TLATX1 dout_reg_76_ ( .G(n324), .D(N107), .Q(dout[76]) );
  TLATX1 dout_reg_44_ ( .G(n328), .D(N75), .Q(dout[44]) );
  TLATX1 dout_reg_28_ ( .G(n326), .D(N59), .Q(dout[28]) );
  TLATX1 dout_reg_107_ ( .G(N30), .D(N139), .Q(dout[107]) );
  TLATX1 dout_reg_75_ ( .G(n318), .D(N106), .Q(dout[75]) );
  TLATX1 dout_reg_43_ ( .G(n330), .D(N74), .Q(dout[43]) );
  TLATX1 dout_reg_27_ ( .G(n324), .D(N58), .Q(dout[27]) );
  TLATX1 dout_reg_106_ ( .G(n323), .D(N138), .Q(dout[106]) );
  TLATX1 dout_reg_74_ ( .G(n321), .D(N105), .Q(dout[74]) );
  TLATX1 dout_reg_42_ ( .G(n329), .D(N73), .Q(dout[42]) );
  TLATX1 dout_reg_26_ ( .G(n320), .D(N57), .Q(dout[26]) );
  TLATX1 dout_reg_105_ ( .G(N30), .D(N137), .Q(dout[105]) );
  TLATX1 dout_reg_73_ ( .G(N30), .D(N104), .Q(dout[73]) );
  TLATX1 dout_reg_41_ ( .G(n327), .D(N72), .Q(dout[41]) );
  TLATX1 dout_reg_25_ ( .G(n325), .D(N56), .Q(dout[25]) );
  TLATX1 dout_reg_104_ ( .G(n322), .D(N136), .Q(dout[104]) );
  TLATX1 dout_reg_72_ ( .G(n328), .D(N103), .Q(dout[72]) );
  TLATX1 dout_reg_40_ ( .G(n326), .D(N71), .Q(dout[40]) );
  TLATX1 dout_reg_24_ ( .G(N30), .D(N55), .Q(dout[24]) );
  TLATX1 dout_reg_103_ ( .G(n330), .D(N135), .Q(dout[103]) );
  TLATX1 dout_reg_71_ ( .G(n330), .D(N102), .Q(dout[71]) );
  TLATX1 dout_reg_39_ ( .G(n330), .D(N70), .Q(dout[39]) );
  TLATX1 dout_reg_23_ ( .G(n330), .D(N54), .Q(dout[23]) );
  TLATX1 dout_reg_102_ ( .G(n330), .D(N134), .Q(dout[102]) );
  TLATX1 dout_reg_70_ ( .G(n330), .D(N101), .Q(dout[70]) );
  TLATX1 dout_reg_38_ ( .G(n320), .D(N69), .Q(dout[38]) );
  TLATX1 dout_reg_22_ ( .G(n327), .D(N53), .Q(dout[22]) );
  TLATX1 dout_reg_101_ ( .G(n325), .D(N133), .Q(dout[101]) );
  TLATX1 dout_reg_69_ ( .G(n322), .D(N100), .Q(dout[69]) );
  TLATX1 dout_reg_37_ ( .G(n328), .D(N68), .Q(dout[37]) );
  TLATX1 dout_reg_21_ ( .G(n326), .D(N52), .Q(dout[21]) );
  TLATX1 dout_reg_100_ ( .G(n329), .D(N132), .Q(dout[100]) );
  TLATX1 dout_reg_68_ ( .G(n329), .D(N99), .Q(dout[68]) );
  TLATX1 dout_reg_36_ ( .G(n329), .D(N67), .Q(dout[36]) );
  TLATX1 dout_reg_20_ ( .G(n329), .D(N51), .Q(dout[20]) );
  TLATX1 dout_reg_99_ ( .G(n329), .D(N131), .Q(dout[99]) );
  TLATX1 dout_reg_67_ ( .G(n329), .D(N98), .Q(dout[67]) );
  TLATX1 dout_reg_35_ ( .G(n328), .D(N66), .Q(dout[35]) );
  TLATX1 dout_reg_19_ ( .G(n328), .D(N50), .Q(dout[19]) );
  TLATX1 dout_reg_98_ ( .G(n328), .D(N129), .Q(dout[98]) );
  TLATX1 dout_reg_66_ ( .G(n328), .D(N97), .Q(dout[66]) );
  TLATX1 dout_reg_34_ ( .G(n328), .D(N65), .Q(dout[34]) );
  TLATX1 dout_reg_18_ ( .G(n328), .D(N49), .Q(dout[18]) );
  TLATX1 dout_reg_97_ ( .G(n327), .D(N128), .Q(dout[97]) );
  TLATX1 dout_reg_65_ ( .G(n327), .D(N96), .Q(dout[65]) );
  TLATX1 dout_reg_33_ ( .G(n327), .D(N64), .Q(dout[33]) );
  TLATX1 dout_reg_17_ ( .G(n327), .D(N48), .Q(dout[17]) );
  TLATX1 dout_reg_96_ ( .G(n327), .D(N127), .Q(dout[96]) );
  TLATX1 dout_reg_64_ ( .G(n327), .D(N95), .Q(dout[64]) );
  TLATX1 dout_reg_32_ ( .G(n325), .D(N63), .Q(dout[32]) );
  TLATX1 dout_reg_143_ ( .G(n322), .D(N175), .Q(dout[143]) );
  TLATX1 dout_reg_142_ ( .G(n328), .D(N174), .Q(dout[142]) );
  TLATX1 dout_reg_141_ ( .G(n326), .D(N173), .Q(dout[141]) );
  TLATX1 dout_reg_140_ ( .G(n326), .D(N172), .Q(dout[140]) );
  TLATX1 dout_reg_139_ ( .G(n326), .D(N171), .Q(dout[139]) );
  TLATX1 dout_reg_138_ ( .G(n325), .D(N170), .Q(dout[138]) );
  TLATX1 dout_reg_137_ ( .G(n325), .D(N169), .Q(dout[137]) );
  TLATX1 dout_reg_136_ ( .G(n325), .D(N168), .Q(dout[136]) );
  TLATX1 dout_reg_135_ ( .G(n324), .D(N167), .Q(dout[135]) );
  TLATX1 dout_reg_134_ ( .G(n324), .D(N166), .Q(dout[134]) );
  TLATX1 dout_reg_133_ ( .G(n324), .D(N165), .Q(dout[133]) );
  TLATX1 dout_reg_132_ ( .G(n323), .D(N164), .Q(dout[132]) );
  TLATX1 dout_reg_131_ ( .G(n323), .D(N163), .Q(dout[131]) );
  TLATX1 dout_reg_130_ ( .G(n323), .D(N162), .Q(dout[130]) );
  TLATX1 dout_reg_129_ ( .G(n322), .D(N161), .Q(dout[129]) );
  TLATX1 dout_reg_128_ ( .G(n322), .D(N160), .Q(dout[128]) );
  TLATX1 dout_reg_15_ ( .G(n330), .D(N46), .Q(dout[15]) );
  TLATX1 dout_reg_14_ ( .G(n324), .D(N45), .Q(dout[14]) );
  TLATX1 dout_reg_13_ ( .G(n323), .D(N44), .Q(dout[13]) );
  TLATX1 dout_reg_12_ ( .G(n323), .D(N43), .Q(dout[12]) );
  TLATX1 dout_reg_11_ ( .G(n321), .D(N42), .Q(dout[11]) );
  TLATX1 dout_reg_10_ ( .G(N30), .D(N41), .Q(dout[10]) );
  TLATX1 dout_reg_9_ ( .G(n318), .D(N40), .Q(dout[9]) );
  TLATX1 dout_reg_8_ ( .G(n330), .D(N39), .Q(dout[8]) );
  TLATX1 dout_reg_7_ ( .G(n330), .D(N38), .Q(dout[7]) );
  TLATX1 dout_reg_6_ ( .G(n320), .D(N37), .Q(dout[6]) );
  TLATX1 dout_reg_5_ ( .G(n327), .D(N36), .Q(dout[5]) );
  TLATX1 dout_reg_4_ ( .G(n329), .D(N35), .Q(dout[4]) );
  TLATX1 dout_reg_3_ ( .G(n328), .D(N34), .Q(dout[3]) );
  TLATX1 dout_reg_2_ ( .G(n328), .D(N33), .Q(dout[2]) );
  TLATX1 dout_reg_1_ ( .G(n327), .D(N32), .Q(dout[1]) );
  TLATX1 dout_reg_0_ ( .G(n326), .D(N31), .Q(dout[0]) );
  TLATX1 dout_reg_255_ ( .G(n322), .D(N288), .Q(dout[255]) );
  TLATX1 dout_reg_254_ ( .G(n321), .D(N287), .Q(dout[254]) );
  TLATX1 dout_reg_253_ ( .G(n321), .D(N286), .Q(dout[253]) );
  TLATX1 dout_reg_252_ ( .G(n321), .D(N285), .Q(dout[252]) );
  TLATX1 dout_reg_251_ ( .G(n321), .D(N284), .Q(dout[251]) );
  TLATX1 dout_reg_250_ ( .G(n329), .D(N283), .Q(dout[250]) );
  TLATX1 dout_reg_249_ ( .G(n319), .D(N282), .Q(dout[249]) );
  TLATX1 dout_reg_248_ ( .G(n320), .D(N281), .Q(dout[248]) );
  TLATX1 dout_reg_247_ ( .G(n320), .D(N280), .Q(dout[247]) );
  TLATX1 dout_reg_246_ ( .G(n320), .D(N279), .Q(dout[246]) );
  TLATX1 dout_reg_245_ ( .G(n319), .D(N278), .Q(dout[245]) );
  TLATX1 dout_reg_244_ ( .G(n319), .D(N277), .Q(dout[244]) );
  TLATX1 dout_reg_243_ ( .G(n319), .D(N276), .Q(dout[243]) );
  TLATX1 dout_reg_242_ ( .G(n318), .D(N275), .Q(dout[242]) );
  TLATX1 dout_reg_241_ ( .G(n318), .D(N274), .Q(dout[241]) );
  TLATX1 dout_reg_240_ ( .G(n318), .D(N273), .Q(dout[240]) );
  TLATX1 dout_reg_127_ ( .G(N30), .D(N159), .Q(dout[127]) );
  TLATX1 dout_reg_95_ ( .G(N30), .D(N126), .Q(dout[95]) );
  TLATX1 dout_reg_63_ ( .G(n323), .D(N94), .Q(dout[63]) );
  TLATX1 dout_reg_126_ ( .G(n321), .D(N158), .Q(dout[126]) );
  TLATX1 dout_reg_94_ ( .G(n329), .D(N125), .Q(dout[94]) );
  TLATX1 dout_reg_62_ ( .G(n327), .D(N93), .Q(dout[62]) );
  TLATX1 dout_reg_125_ ( .G(n321), .D(N157), .Q(dout[125]) );
  TLATX1 dout_reg_93_ ( .G(n329), .D(N124), .Q(dout[93]) );
  TLATX1 dout_reg_61_ ( .G(n325), .D(N92), .Q(dout[61]) );
  TLATX1 dout_reg_124_ ( .G(n320), .D(N156), .Q(dout[124]) );
  TLATX1 dout_reg_92_ ( .G(n319), .D(N123), .Q(dout[92]) );
  TLATX1 dout_reg_60_ ( .G(n329), .D(N91), .Q(dout[60]) );
  TLATX1 dout_reg_123_ ( .G(n322), .D(N155), .Q(dout[123]) );
  TLATX1 dout_reg_91_ ( .G(n320), .D(N122), .Q(dout[91]) );
  TLATX1 dout_reg_59_ ( .G(n319), .D(N90), .Q(dout[59]) );
  TLATX1 dout_reg_122_ ( .G(N30), .D(N154), .Q(dout[122]) );
  TLATX1 dout_reg_90_ ( .G(N30), .D(N121), .Q(dout[90]) );
  TLATX1 dout_reg_58_ ( .G(N30), .D(N89), .Q(dout[58]) );
  TLATX1 dout_reg_121_ ( .G(N30), .D(N153), .Q(dout[121]) );
  TLATX1 dout_reg_89_ ( .G(N30), .D(N120), .Q(dout[89]) );
  TLATX1 dout_reg_57_ ( .G(n324), .D(N88), .Q(dout[57]) );
  TLATX1 dout_reg_120_ ( .G(n323), .D(N152), .Q(dout[120]) );
  TLATX1 dout_reg_88_ ( .G(n321), .D(N119), .Q(dout[88]) );
  TLATX1 dout_reg_56_ ( .G(n329), .D(N87), .Q(dout[56]) );
  TLATX1 dout_reg_119_ ( .G(n330), .D(N151), .Q(dout[119]) );
  TLATX1 dout_reg_87_ ( .G(n330), .D(N118), .Q(dout[87]) );
  TLATX1 dout_reg_55_ ( .G(n330), .D(N86), .Q(dout[55]) );
  TLATX1 dout_reg_118_ ( .G(n330), .D(N150), .Q(dout[118]) );
  TLATX1 dout_reg_86_ ( .G(n330), .D(N117), .Q(dout[86]) );
  TLATX1 dout_reg_54_ ( .G(n323), .D(N85), .Q(dout[54]) );
  TLATX1 dout_reg_117_ ( .G(n327), .D(N149), .Q(dout[117]) );
  TLATX1 dout_reg_85_ ( .G(n330), .D(N116), .Q(dout[85]) );
  TLATX1 dout_reg_53_ ( .G(n324), .D(N84), .Q(dout[53]) );
  TLATX1 dout_reg_116_ ( .G(n329), .D(N148), .Q(dout[116]) );
  TLATX1 dout_reg_84_ ( .G(n329), .D(N115), .Q(dout[84]) );
  TLATX1 dout_reg_52_ ( .G(n329), .D(N83), .Q(dout[52]) );
  TLATX1 dout_reg_115_ ( .G(n329), .D(N147), .Q(dout[115]) );
  TLATX1 dout_reg_83_ ( .G(n329), .D(N114), .Q(dout[83]) );
  TLATX1 dout_reg_51_ ( .G(n328), .D(N82), .Q(dout[51]) );
  TLATX1 dout_reg_114_ ( .G(n328), .D(N146), .Q(dout[114]) );
  TLATX1 dout_reg_82_ ( .G(n328), .D(N113), .Q(dout[82]) );
  TLATX1 dout_reg_50_ ( .G(n328), .D(N81), .Q(dout[50]) );
  TLATX1 dout_reg_113_ ( .G(n327), .D(N145), .Q(dout[113]) );
  TLATX1 dout_reg_81_ ( .G(n327), .D(N112), .Q(dout[81]) );
  TLATX1 dout_reg_49_ ( .G(n327), .D(N80), .Q(dout[49]) );
  TLATX1 dout_reg_112_ ( .G(n327), .D(N144), .Q(dout[112]) );
  TLATX1 dout_reg_80_ ( .G(n327), .D(N111), .Q(dout[80]) );
  TLATX1 dout_reg_48_ ( .G(N30), .D(N79), .Q(dout[48]) );
  TLATX1 dout_reg_175_ ( .G(n318), .D(N207), .Q(dout[175]) );
  TLATX1 dout_reg_174_ ( .G(n319), .D(N206), .Q(dout[174]) );
  TLATX1 dout_reg_173_ ( .G(n326), .D(N205), .Q(dout[173]) );
  TLATX1 dout_reg_172_ ( .G(n326), .D(N204), .Q(dout[172]) );
  TLATX1 dout_reg_171_ ( .G(n326), .D(N203), .Q(dout[171]) );
  TLATX1 dout_reg_170_ ( .G(n325), .D(N202), .Q(dout[170]) );
  TLATX1 dout_reg_169_ ( .G(n325), .D(N201), .Q(dout[169]) );
  TLATX1 dout_reg_168_ ( .G(n325), .D(N200), .Q(dout[168]) );
  TLATX1 dout_reg_167_ ( .G(n324), .D(N199), .Q(dout[167]) );
  TLATX1 dout_reg_166_ ( .G(n324), .D(N198), .Q(dout[166]) );
  TLATX1 dout_reg_165_ ( .G(n324), .D(N197), .Q(dout[165]) );
  TLATX1 dout_reg_164_ ( .G(n323), .D(N196), .Q(dout[164]) );
  TLATX1 dout_reg_163_ ( .G(n323), .D(N195), .Q(dout[163]) );
  TLATX1 dout_reg_162_ ( .G(n323), .D(N194), .Q(dout[162]) );
  TLATX1 dout_reg_161_ ( .G(n322), .D(N193), .Q(dout[161]) );
  TLATX1 dout_reg_160_ ( .G(n322), .D(N192), .Q(dout[160]) );
  TLATX1 dout_reg_239_ ( .G(n322), .D(N272), .Q(dout[239]) );
  TLATX1 dout_reg_207_ ( .G(n322), .D(N240), .Q(dout[207]) );
  TLATX1 dout_reg_238_ ( .G(n321), .D(N271), .Q(dout[238]) );
  TLATX1 dout_reg_206_ ( .G(n321), .D(N239), .Q(dout[206]) );
  TLATX1 dout_reg_237_ ( .G(n321), .D(N270), .Q(dout[237]) );
  TLATX1 dout_reg_205_ ( .G(n321), .D(N238), .Q(dout[205]) );
  TLATX1 dout_reg_236_ ( .G(n321), .D(N269), .Q(dout[236]) );
  TLATX1 dout_reg_204_ ( .G(n321), .D(N237), .Q(dout[204]) );
  TLATX1 dout_reg_235_ ( .G(n320), .D(N268), .Q(dout[235]) );
  TLATX1 dout_reg_203_ ( .G(n319), .D(N236), .Q(dout[203]) );
  TLATX1 dout_reg_234_ ( .G(n327), .D(N267), .Q(dout[234]) );
  TLATX1 dout_reg_202_ ( .G(n325), .D(N235), .Q(dout[202]) );
  TLATX1 dout_reg_233_ ( .G(n322), .D(N266), .Q(dout[233]) );
  TLATX1 dout_reg_201_ ( .G(n328), .D(N234), .Q(dout[201]) );
  TLATX1 dout_reg_232_ ( .G(n320), .D(N265), .Q(dout[232]) );
  TLATX1 dout_reg_200_ ( .G(n320), .D(N233), .Q(dout[200]) );
  TLATX1 dout_reg_231_ ( .G(n320), .D(N264), .Q(dout[231]) );
  TLATX1 dout_reg_199_ ( .G(n320), .D(N232), .Q(dout[199]) );
  TLATX1 dout_reg_230_ ( .G(n320), .D(N263), .Q(dout[230]) );
  TLATX1 dout_reg_198_ ( .G(n320), .D(N231), .Q(dout[198]) );
  TLATX1 dout_reg_229_ ( .G(n319), .D(N262), .Q(dout[229]) );
  TLATX1 dout_reg_197_ ( .G(n319), .D(N229), .Q(dout[197]) );
  TLATX1 dout_reg_228_ ( .G(n319), .D(N261), .Q(dout[228]) );
  TLATX1 dout_reg_196_ ( .G(n319), .D(N228), .Q(dout[196]) );
  TLATX1 dout_reg_227_ ( .G(n319), .D(N260), .Q(dout[227]) );
  TLATX1 dout_reg_195_ ( .G(n319), .D(N227), .Q(dout[195]) );
  TLATX1 dout_reg_226_ ( .G(n318), .D(N259), .Q(dout[226]) );
  TLATX1 dout_reg_194_ ( .G(n318), .D(N226), .Q(dout[194]) );
  TLATX1 dout_reg_225_ ( .G(n318), .D(N258), .Q(dout[225]) );
  TLATX1 dout_reg_193_ ( .G(n318), .D(N225), .Q(dout[193]) );
  TLATX1 dout_reg_224_ ( .G(n318), .D(N257), .Q(dout[224]) );
  TLATX1 dout_reg_192_ ( .G(n318), .D(N224), .Q(dout[192]) );
  TLATX1 dout_reg_191_ ( .G(n325), .D(N223), .Q(dout[191]) );
  TLATX1 dout_reg_159_ ( .G(n325), .D(N191), .Q(dout[159]) );
  TLATX1 dout_reg_190_ ( .G(n330), .D(N222), .Q(dout[190]) );
  TLATX1 dout_reg_158_ ( .G(n324), .D(N190), .Q(dout[158]) );
  TLATX1 dout_reg_189_ ( .G(n326), .D(N221), .Q(dout[189]) );
  TLATX1 dout_reg_157_ ( .G(n326), .D(N189), .Q(dout[157]) );
  TLATX1 dout_reg_188_ ( .G(n326), .D(N220), .Q(dout[188]) );
  TLATX1 dout_reg_156_ ( .G(n326), .D(N188), .Q(dout[156]) );
  TLATX1 dout_reg_187_ ( .G(n326), .D(N219), .Q(dout[187]) );
  TLATX1 dout_reg_155_ ( .G(n326), .D(N187), .Q(dout[155]) );
  TLATX1 dout_reg_186_ ( .G(n325), .D(N218), .Q(dout[186]) );
  TLATX1 dout_reg_154_ ( .G(n325), .D(N186), .Q(dout[154]) );
  TLATX1 dout_reg_185_ ( .G(n325), .D(N217), .Q(dout[185]) );
  TLATX1 dout_reg_153_ ( .G(n325), .D(N185), .Q(dout[153]) );
  TLATX1 dout_reg_184_ ( .G(n325), .D(N216), .Q(dout[184]) );
  TLATX1 dout_reg_152_ ( .G(n325), .D(N184), .Q(dout[152]) );
  TLATX1 dout_reg_183_ ( .G(n324), .D(N215), .Q(dout[183]) );
  TLATX1 dout_reg_151_ ( .G(n324), .D(N183), .Q(dout[151]) );
  TLATX1 dout_reg_182_ ( .G(n324), .D(N214), .Q(dout[182]) );
  TLATX1 dout_reg_150_ ( .G(n324), .D(N182), .Q(dout[150]) );
  TLATX1 dout_reg_181_ ( .G(n324), .D(N213), .Q(dout[181]) );
  TLATX1 dout_reg_149_ ( .G(n324), .D(N181), .Q(dout[149]) );
  TLATX1 dout_reg_180_ ( .G(n323), .D(N212), .Q(dout[180]) );
  TLATX1 dout_reg_148_ ( .G(n323), .D(N180), .Q(dout[148]) );
  TLATX1 dout_reg_179_ ( .G(n323), .D(N211), .Q(dout[179]) );
  TLATX1 dout_reg_147_ ( .G(n323), .D(N179), .Q(dout[147]) );
  TLATX1 dout_reg_178_ ( .G(n323), .D(N210), .Q(dout[178]) );
  TLATX1 dout_reg_146_ ( .G(n323), .D(N178), .Q(dout[146]) );
  TLATX1 dout_reg_177_ ( .G(n322), .D(N209), .Q(dout[177]) );
  TLATX1 dout_reg_145_ ( .G(n322), .D(N177), .Q(dout[145]) );
  TLATX1 dout_reg_176_ ( .G(n322), .D(N208), .Q(dout[176]) );
  TLATX1 dout_reg_144_ ( .G(n322), .D(N176), .Q(dout[144]) );
  TLATX1 dout_reg_223_ ( .G(n322), .D(N256), .Q(dout[223]) );
  TLATX1 dout_reg_222_ ( .G(n321), .D(N255), .Q(dout[222]) );
  TLATX1 dout_reg_221_ ( .G(n321), .D(N254), .Q(dout[221]) );
  TLATX1 dout_reg_220_ ( .G(n321), .D(N253), .Q(dout[220]) );
  TLATX1 dout_reg_219_ ( .G(n326), .D(N252), .Q(dout[219]) );
  TLATX1 dout_reg_218_ ( .G(N30), .D(N251), .Q(dout[218]) );
  TLATX1 dout_reg_217_ ( .G(N30), .D(N250), .Q(dout[217]) );
  TLATX1 dout_reg_216_ ( .G(n320), .D(N249), .Q(dout[216]) );
  TLATX1 dout_reg_215_ ( .G(n320), .D(N248), .Q(dout[215]) );
  TLATX1 dout_reg_214_ ( .G(n320), .D(N247), .Q(dout[214]) );
  TLATX1 dout_reg_213_ ( .G(n319), .D(N246), .Q(dout[213]) );
  TLATX1 dout_reg_212_ ( .G(n319), .D(N245), .Q(dout[212]) );
  TLATX1 dout_reg_211_ ( .G(n319), .D(N244), .Q(dout[211]) );
  TLATX1 dout_reg_210_ ( .G(n318), .D(N243), .Q(dout[210]) );
  TLATX1 dout_reg_209_ ( .G(n318), .D(N242), .Q(dout[209]) );
  TLATX1 dout_reg_208_ ( .G(n318), .D(N241), .Q(dout[208]) );
  DFFRHQX1 dout16_reg_reg_207_ ( .D(n1478), .CK(clk), .RN(rstn), .Q(
        dout16_reg[207]) );
  DFFRHQX1 dout16_reg_reg_223_ ( .D(n1494), .CK(clk), .RN(rstn), .Q(
        dout16_reg[223]) );
  DFFRHQX1 dout16_reg_reg_239_ ( .D(n1510), .CK(clk), .RN(rstn), .Q(
        dout16_reg[239]) );
  DFFRHQX1 dout16_reg_reg_255_ ( .D(n1526), .CK(clk), .RN(rstn), .Q(
        dout16_reg[255]) );
  DFFRHQX1 dout16_reg_reg_206_ ( .D(n1477), .CK(clk), .RN(rstn), .Q(
        dout16_reg[206]) );
  DFFRHQX1 dout16_reg_reg_222_ ( .D(n1493), .CK(clk), .RN(rstn), .Q(
        dout16_reg[222]) );
  DFFRHQX1 dout16_reg_reg_238_ ( .D(n1509), .CK(clk), .RN(rstn), .Q(
        dout16_reg[238]) );
  DFFRHQX1 dout16_reg_reg_254_ ( .D(n1525), .CK(clk), .RN(rstn), .Q(
        dout16_reg[254]) );
  DFFRHQX1 dout16_reg_reg_205_ ( .D(n1476), .CK(clk), .RN(rstn), .Q(
        dout16_reg[205]) );
  DFFRHQX1 dout16_reg_reg_221_ ( .D(n1492), .CK(clk), .RN(rstn), .Q(
        dout16_reg[221]) );
  DFFRHQX1 dout16_reg_reg_237_ ( .D(n1508), .CK(clk), .RN(rstn), .Q(
        dout16_reg[237]) );
  DFFRHQX1 dout16_reg_reg_253_ ( .D(n1524), .CK(clk), .RN(rstn), .Q(
        dout16_reg[253]) );
  DFFRHQX1 dout16_reg_reg_204_ ( .D(n1475), .CK(clk), .RN(rstn), .Q(
        dout16_reg[204]) );
  DFFRHQX1 dout16_reg_reg_220_ ( .D(n1491), .CK(clk), .RN(rstn), .Q(
        dout16_reg[220]) );
  DFFRHQX1 dout16_reg_reg_236_ ( .D(n1507), .CK(clk), .RN(rstn), .Q(
        dout16_reg[236]) );
  DFFRHQX1 dout16_reg_reg_252_ ( .D(n1523), .CK(clk), .RN(rstn), .Q(
        dout16_reg[252]) );
  DFFRHQX1 dout16_reg_reg_203_ ( .D(n1474), .CK(clk), .RN(rstn), .Q(
        dout16_reg[203]) );
  DFFRHQX1 dout16_reg_reg_219_ ( .D(n1490), .CK(clk), .RN(rstn), .Q(
        dout16_reg[219]) );
  DFFRHQX1 dout16_reg_reg_235_ ( .D(n1506), .CK(clk), .RN(rstn), .Q(
        dout16_reg[235]) );
  DFFRHQX1 dout16_reg_reg_251_ ( .D(n1522), .CK(clk), .RN(rstn), .Q(
        dout16_reg[251]) );
  DFFRHQX1 dout16_reg_reg_202_ ( .D(n1473), .CK(clk), .RN(rstn), .Q(
        dout16_reg[202]) );
  DFFRHQX1 dout16_reg_reg_218_ ( .D(n1489), .CK(clk), .RN(rstn), .Q(
        dout16_reg[218]) );
  DFFRHQX1 dout16_reg_reg_234_ ( .D(n1505), .CK(clk), .RN(rstn), .Q(
        dout16_reg[234]) );
  DFFRHQX1 dout16_reg_reg_250_ ( .D(n1521), .CK(clk), .RN(rstn), .Q(
        dout16_reg[250]) );
  DFFRHQX1 dout16_reg_reg_201_ ( .D(n1472), .CK(clk), .RN(rstn), .Q(
        dout16_reg[201]) );
  DFFRHQX1 dout16_reg_reg_217_ ( .D(n1488), .CK(clk), .RN(rstn), .Q(
        dout16_reg[217]) );
  DFFRHQX1 dout16_reg_reg_233_ ( .D(n1504), .CK(clk), .RN(rstn), .Q(
        dout16_reg[233]) );
  DFFRHQX1 dout16_reg_reg_249_ ( .D(n1520), .CK(clk), .RN(rstn), .Q(
        dout16_reg[249]) );
  DFFRHQX1 dout16_reg_reg_200_ ( .D(n1471), .CK(clk), .RN(rstn), .Q(
        dout16_reg[200]) );
  DFFRHQX1 dout16_reg_reg_216_ ( .D(n1487), .CK(clk), .RN(rstn), .Q(
        dout16_reg[216]) );
  DFFRHQX1 dout16_reg_reg_232_ ( .D(n1503), .CK(clk), .RN(rstn), .Q(
        dout16_reg[232]) );
  DFFRHQX1 dout16_reg_reg_248_ ( .D(n1519), .CK(clk), .RN(rstn), .Q(
        dout16_reg[248]) );
  DFFRHQX1 dout16_reg_reg_199_ ( .D(n1470), .CK(clk), .RN(rstn), .Q(
        dout16_reg[199]) );
  DFFRHQX1 dout16_reg_reg_215_ ( .D(n1486), .CK(clk), .RN(rstn), .Q(
        dout16_reg[215]) );
  DFFRHQX1 dout16_reg_reg_231_ ( .D(n1502), .CK(clk), .RN(rstn), .Q(
        dout16_reg[231]) );
  DFFRHQX1 dout16_reg_reg_247_ ( .D(n1518), .CK(clk), .RN(rstn), .Q(
        dout16_reg[247]) );
  DFFRHQX1 dout16_reg_reg_198_ ( .D(n1469), .CK(clk), .RN(rstn), .Q(
        dout16_reg[198]) );
  DFFRHQX1 dout16_reg_reg_214_ ( .D(n1485), .CK(clk), .RN(rstn), .Q(
        dout16_reg[214]) );
  DFFRHQX1 dout16_reg_reg_230_ ( .D(n1501), .CK(clk), .RN(rstn), .Q(
        dout16_reg[230]) );
  DFFRHQX1 dout16_reg_reg_246_ ( .D(n1517), .CK(clk), .RN(rstn), .Q(
        dout16_reg[246]) );
  DFFRHQX1 dout16_reg_reg_197_ ( .D(n1468), .CK(clk), .RN(rstn), .Q(
        dout16_reg[197]) );
  DFFRHQX1 dout16_reg_reg_213_ ( .D(n1484), .CK(clk), .RN(rstn), .Q(
        dout16_reg[213]) );
  DFFRHQX1 dout16_reg_reg_229_ ( .D(n1500), .CK(clk), .RN(rstn), .Q(
        dout16_reg[229]) );
  DFFRHQX1 dout16_reg_reg_245_ ( .D(n1516), .CK(clk), .RN(rstn), .Q(
        dout16_reg[245]) );
  DFFRHQX1 dout16_reg_reg_196_ ( .D(n1467), .CK(clk), .RN(rstn), .Q(
        dout16_reg[196]) );
  DFFRHQX1 dout16_reg_reg_212_ ( .D(n1483), .CK(clk), .RN(rstn), .Q(
        dout16_reg[212]) );
  DFFRHQX1 dout16_reg_reg_228_ ( .D(n1499), .CK(clk), .RN(rstn), .Q(
        dout16_reg[228]) );
  DFFRHQX1 dout16_reg_reg_244_ ( .D(n1515), .CK(clk), .RN(rstn), .Q(
        dout16_reg[244]) );
  DFFRHQX1 dout16_reg_reg_195_ ( .D(n1466), .CK(clk), .RN(rstn), .Q(
        dout16_reg[195]) );
  DFFRHQX1 dout16_reg_reg_211_ ( .D(n1482), .CK(clk), .RN(rstn), .Q(
        dout16_reg[211]) );
  DFFRHQX1 dout16_reg_reg_227_ ( .D(n1498), .CK(clk), .RN(rstn), .Q(
        dout16_reg[227]) );
  DFFRHQX1 dout16_reg_reg_243_ ( .D(n1514), .CK(clk), .RN(rstn), .Q(
        dout16_reg[243]) );
  DFFRHQX1 dout16_reg_reg_194_ ( .D(n1465), .CK(clk), .RN(rstn), .Q(
        dout16_reg[194]) );
  DFFRHQX1 dout16_reg_reg_210_ ( .D(n1481), .CK(clk), .RN(rstn), .Q(
        dout16_reg[210]) );
  DFFRHQX1 dout16_reg_reg_226_ ( .D(n1497), .CK(clk), .RN(rstn), .Q(
        dout16_reg[226]) );
  DFFRHQX1 dout16_reg_reg_242_ ( .D(n1513), .CK(clk), .RN(rstn), .Q(
        dout16_reg[242]) );
  DFFRHQX1 dout16_reg_reg_193_ ( .D(n1464), .CK(clk), .RN(rstn), .Q(
        dout16_reg[193]) );
  DFFRHQX1 dout16_reg_reg_209_ ( .D(n1480), .CK(clk), .RN(rstn), .Q(
        dout16_reg[209]) );
  DFFRHQX1 dout16_reg_reg_225_ ( .D(n1496), .CK(clk), .RN(rstn), .Q(
        dout16_reg[225]) );
  DFFRHQX1 dout16_reg_reg_241_ ( .D(n1512), .CK(clk), .RN(rstn), .Q(
        dout16_reg[241]) );
  DFFRHQX1 dout16_reg_reg_192_ ( .D(n1463), .CK(clk), .RN(rstn), .Q(
        dout16_reg[192]) );
  DFFRHQX1 dout16_reg_reg_208_ ( .D(n1479), .CK(clk), .RN(rstn), .Q(
        dout16_reg[208]) );
  DFFRHQX1 dout16_reg_reg_224_ ( .D(n1495), .CK(clk), .RN(rstn), .Q(
        dout16_reg[224]) );
  DFFRHQX1 dout16_reg_reg_240_ ( .D(n1511), .CK(clk), .RN(rstn), .Q(
        dout16_reg[240]) );
  DFFRHQX1 dout8_reg_reg_79_ ( .D(n1606), .CK(clk), .RN(rstn), .Q(
        dout8_reg[79]) );
  DFFRHQX1 dout8_reg_reg_95_ ( .D(n1622), .CK(clk), .RN(rstn), .Q(
        dout8_reg[95]) );
  DFFRHQX1 dout8_reg_reg_111_ ( .D(n1638), .CK(clk), .RN(rstn), .Q(
        dout8_reg[111]) );
  DFFRHQX1 dout8_reg_reg_127_ ( .D(n1654), .CK(clk), .RN(rstn), .Q(
        dout8_reg[127]) );
  DFFRHQX1 dout8_reg_reg_78_ ( .D(n1605), .CK(clk), .RN(rstn), .Q(
        dout8_reg[78]) );
  DFFRHQX1 dout8_reg_reg_94_ ( .D(n1621), .CK(clk), .RN(rstn), .Q(
        dout8_reg[94]) );
  DFFRHQX1 dout8_reg_reg_110_ ( .D(n1637), .CK(clk), .RN(rstn), .Q(
        dout8_reg[110]) );
  DFFRHQX1 dout8_reg_reg_126_ ( .D(n1653), .CK(clk), .RN(rstn), .Q(
        dout8_reg[126]) );
  DFFRHQX1 dout8_reg_reg_77_ ( .D(n1604), .CK(clk), .RN(rstn), .Q(
        dout8_reg[77]) );
  DFFRHQX1 dout8_reg_reg_93_ ( .D(n1620), .CK(clk), .RN(rstn), .Q(
        dout8_reg[93]) );
  DFFRHQX1 dout8_reg_reg_109_ ( .D(n1636), .CK(clk), .RN(rstn), .Q(
        dout8_reg[109]) );
  DFFRHQX1 dout8_reg_reg_125_ ( .D(n1652), .CK(clk), .RN(rstn), .Q(
        dout8_reg[125]) );
  DFFRHQX1 dout8_reg_reg_76_ ( .D(n1603), .CK(clk), .RN(rstn), .Q(
        dout8_reg[76]) );
  DFFRHQX1 dout8_reg_reg_92_ ( .D(n1619), .CK(clk), .RN(rstn), .Q(
        dout8_reg[92]) );
  DFFRHQX1 dout8_reg_reg_108_ ( .D(n1635), .CK(clk), .RN(rstn), .Q(
        dout8_reg[108]) );
  DFFRHQX1 dout8_reg_reg_124_ ( .D(n1651), .CK(clk), .RN(rstn), .Q(
        dout8_reg[124]) );
  DFFRHQX1 dout8_reg_reg_75_ ( .D(n1602), .CK(clk), .RN(rstn), .Q(
        dout8_reg[75]) );
  DFFRHQX1 dout8_reg_reg_91_ ( .D(n1618), .CK(clk), .RN(rstn), .Q(
        dout8_reg[91]) );
  DFFRHQX1 dout8_reg_reg_107_ ( .D(n1634), .CK(clk), .RN(rstn), .Q(
        dout8_reg[107]) );
  DFFRHQX1 dout8_reg_reg_123_ ( .D(n1650), .CK(clk), .RN(rstn), .Q(
        dout8_reg[123]) );
  DFFRHQX1 dout8_reg_reg_74_ ( .D(n1601), .CK(clk), .RN(rstn), .Q(
        dout8_reg[74]) );
  DFFRHQX1 dout8_reg_reg_90_ ( .D(n1617), .CK(clk), .RN(rstn), .Q(
        dout8_reg[90]) );
  DFFRHQX1 dout8_reg_reg_106_ ( .D(n1633), .CK(clk), .RN(rstn), .Q(
        dout8_reg[106]) );
  DFFRHQX1 dout8_reg_reg_122_ ( .D(n1649), .CK(clk), .RN(rstn), .Q(
        dout8_reg[122]) );
  DFFRHQX1 dout8_reg_reg_73_ ( .D(n1600), .CK(clk), .RN(rstn), .Q(
        dout8_reg[73]) );
  DFFRHQX1 dout8_reg_reg_89_ ( .D(n1616), .CK(clk), .RN(rstn), .Q(
        dout8_reg[89]) );
  DFFRHQX1 dout8_reg_reg_105_ ( .D(n1632), .CK(clk), .RN(rstn), .Q(
        dout8_reg[105]) );
  DFFRHQX1 dout8_reg_reg_121_ ( .D(n1648), .CK(clk), .RN(rstn), .Q(
        dout8_reg[121]) );
  DFFRHQX1 dout8_reg_reg_72_ ( .D(n1599), .CK(clk), .RN(rstn), .Q(
        dout8_reg[72]) );
  DFFRHQX1 dout8_reg_reg_88_ ( .D(n1615), .CK(clk), .RN(rstn), .Q(
        dout8_reg[88]) );
  DFFRHQX1 dout8_reg_reg_104_ ( .D(n1631), .CK(clk), .RN(rstn), .Q(
        dout8_reg[104]) );
  DFFRHQX1 dout8_reg_reg_120_ ( .D(n1647), .CK(clk), .RN(rstn), .Q(
        dout8_reg[120]) );
  DFFRHQX1 dout8_reg_reg_71_ ( .D(n1598), .CK(clk), .RN(rstn), .Q(
        dout8_reg[71]) );
  DFFRHQX1 dout8_reg_reg_87_ ( .D(n1614), .CK(clk), .RN(rstn), .Q(
        dout8_reg[87]) );
  DFFRHQX1 dout8_reg_reg_103_ ( .D(n1630), .CK(clk), .RN(rstn), .Q(
        dout8_reg[103]) );
  DFFRHQX1 dout8_reg_reg_119_ ( .D(n1646), .CK(clk), .RN(rstn), .Q(
        dout8_reg[119]) );
  DFFRHQX1 dout8_reg_reg_70_ ( .D(n1597), .CK(clk), .RN(rstn), .Q(
        dout8_reg[70]) );
  DFFRHQX1 dout8_reg_reg_86_ ( .D(n1613), .CK(clk), .RN(rstn), .Q(
        dout8_reg[86]) );
  DFFRHQX1 dout8_reg_reg_102_ ( .D(n1629), .CK(clk), .RN(rstn), .Q(
        dout8_reg[102]) );
  DFFRHQX1 dout8_reg_reg_118_ ( .D(n1645), .CK(clk), .RN(rstn), .Q(
        dout8_reg[118]) );
  DFFRHQX1 dout8_reg_reg_69_ ( .D(n1596), .CK(clk), .RN(rstn), .Q(
        dout8_reg[69]) );
  DFFRHQX1 dout8_reg_reg_85_ ( .D(n1612), .CK(clk), .RN(rstn), .Q(
        dout8_reg[85]) );
  DFFRHQX1 dout8_reg_reg_101_ ( .D(n1628), .CK(clk), .RN(rstn), .Q(
        dout8_reg[101]) );
  DFFRHQX1 dout8_reg_reg_117_ ( .D(n1644), .CK(clk), .RN(rstn), .Q(
        dout8_reg[117]) );
  DFFRHQX1 dout8_reg_reg_68_ ( .D(n1595), .CK(clk), .RN(rstn), .Q(
        dout8_reg[68]) );
  DFFRHQX1 dout8_reg_reg_84_ ( .D(n1611), .CK(clk), .RN(rstn), .Q(
        dout8_reg[84]) );
  DFFRHQX1 dout8_reg_reg_100_ ( .D(n1627), .CK(clk), .RN(rstn), .Q(
        dout8_reg[100]) );
  DFFRHQX1 dout8_reg_reg_116_ ( .D(n1643), .CK(clk), .RN(rstn), .Q(
        dout8_reg[116]) );
  DFFRHQX1 dout8_reg_reg_67_ ( .D(n1594), .CK(clk), .RN(rstn), .Q(
        dout8_reg[67]) );
  DFFRHQX1 dout8_reg_reg_83_ ( .D(n1610), .CK(clk), .RN(rstn), .Q(
        dout8_reg[83]) );
  DFFRHQX1 dout8_reg_reg_99_ ( .D(n1626), .CK(clk), .RN(rstn), .Q(
        dout8_reg[99]) );
  DFFRHQX1 dout8_reg_reg_115_ ( .D(n1642), .CK(clk), .RN(rstn), .Q(
        dout8_reg[115]) );
  DFFRHQX1 dout8_reg_reg_66_ ( .D(n1593), .CK(clk), .RN(rstn), .Q(
        dout8_reg[66]) );
  DFFRHQX1 dout8_reg_reg_82_ ( .D(n1609), .CK(clk), .RN(rstn), .Q(
        dout8_reg[82]) );
  DFFRHQX1 dout8_reg_reg_98_ ( .D(n1625), .CK(clk), .RN(rstn), .Q(
        dout8_reg[98]) );
  DFFRHQX1 dout8_reg_reg_114_ ( .D(n1641), .CK(clk), .RN(rstn), .Q(
        dout8_reg[114]) );
  DFFRHQX1 dout8_reg_reg_65_ ( .D(n1592), .CK(clk), .RN(rstn), .Q(
        dout8_reg[65]) );
  DFFRHQX1 dout8_reg_reg_81_ ( .D(n1608), .CK(clk), .RN(rstn), .Q(
        dout8_reg[81]) );
  DFFRHQX1 dout8_reg_reg_97_ ( .D(n1624), .CK(clk), .RN(rstn), .Q(
        dout8_reg[97]) );
  DFFRHQX1 dout8_reg_reg_113_ ( .D(n1640), .CK(clk), .RN(rstn), .Q(
        dout8_reg[113]) );
  DFFRHQX1 dout8_reg_reg_64_ ( .D(n1591), .CK(clk), .RN(rstn), .Q(
        dout8_reg[64]) );
  DFFRHQX1 dout8_reg_reg_80_ ( .D(n1607), .CK(clk), .RN(rstn), .Q(
        dout8_reg[80]) );
  DFFRHQX1 dout8_reg_reg_96_ ( .D(n1623), .CK(clk), .RN(rstn), .Q(
        dout8_reg[96]) );
  DFFRHQX1 dout8_reg_reg_112_ ( .D(n1639), .CK(clk), .RN(rstn), .Q(
        dout8_reg[112]) );
  DFFRHQX1 dout4_reg_reg_15_ ( .D(n1670), .CK(clk), .RN(rstn), .Q(
        dout4_reg[15]) );
  DFFRHQX1 dout4_reg_reg_31_ ( .D(n1686), .CK(clk), .RN(rstn), .Q(
        dout4_reg[31]) );
  DFFRHQX1 dout4_reg_reg_47_ ( .D(n1702), .CK(clk), .RN(rstn), .Q(
        dout4_reg[47]) );
  DFFRHQX1 dout4_reg_reg_63_ ( .D(n1718), .CK(clk), .RN(rstn), .Q(
        dout4_reg[63]) );
  DFFRHQX1 dout4_reg_reg_14_ ( .D(n1669), .CK(clk), .RN(rstn), .Q(
        dout4_reg[14]) );
  DFFRHQX1 dout4_reg_reg_30_ ( .D(n1685), .CK(clk), .RN(rstn), .Q(
        dout4_reg[30]) );
  DFFRHQX1 dout4_reg_reg_46_ ( .D(n1701), .CK(clk), .RN(rstn), .Q(
        dout4_reg[46]) );
  DFFRHQX1 dout4_reg_reg_62_ ( .D(n1717), .CK(clk), .RN(rstn), .Q(
        dout4_reg[62]) );
  DFFRHQX1 dout4_reg_reg_13_ ( .D(n1668), .CK(clk), .RN(rstn), .Q(
        dout4_reg[13]) );
  DFFRHQX1 dout4_reg_reg_29_ ( .D(n1684), .CK(clk), .RN(rstn), .Q(
        dout4_reg[29]) );
  DFFRHQX1 dout4_reg_reg_45_ ( .D(n1700), .CK(clk), .RN(rstn), .Q(
        dout4_reg[45]) );
  DFFRHQX1 dout4_reg_reg_61_ ( .D(n1716), .CK(clk), .RN(rstn), .Q(
        dout4_reg[61]) );
  DFFRHQX1 dout4_reg_reg_12_ ( .D(n1667), .CK(clk), .RN(rstn), .Q(
        dout4_reg[12]) );
  DFFRHQX1 dout4_reg_reg_28_ ( .D(n1683), .CK(clk), .RN(rstn), .Q(
        dout4_reg[28]) );
  DFFRHQX1 dout4_reg_reg_44_ ( .D(n1699), .CK(clk), .RN(rstn), .Q(
        dout4_reg[44]) );
  DFFRHQX1 dout4_reg_reg_60_ ( .D(n1715), .CK(clk), .RN(rstn), .Q(
        dout4_reg[60]) );
  DFFRHQX1 dout4_reg_reg_11_ ( .D(n1666), .CK(clk), .RN(rstn), .Q(
        dout4_reg[11]) );
  DFFRHQX1 dout4_reg_reg_27_ ( .D(n1682), .CK(clk), .RN(rstn), .Q(
        dout4_reg[27]) );
  DFFRHQX1 dout4_reg_reg_43_ ( .D(n1698), .CK(clk), .RN(rstn), .Q(
        dout4_reg[43]) );
  DFFRHQX1 dout4_reg_reg_59_ ( .D(n1714), .CK(clk), .RN(rstn), .Q(
        dout4_reg[59]) );
  DFFRHQX1 dout4_reg_reg_10_ ( .D(n1665), .CK(clk), .RN(rstn), .Q(
        dout4_reg[10]) );
  DFFRHQX1 dout4_reg_reg_26_ ( .D(n1681), .CK(clk), .RN(rstn), .Q(
        dout4_reg[26]) );
  DFFRHQX1 dout4_reg_reg_42_ ( .D(n1697), .CK(clk), .RN(rstn), .Q(
        dout4_reg[42]) );
  DFFRHQX1 dout4_reg_reg_58_ ( .D(n1713), .CK(clk), .RN(rstn), .Q(
        dout4_reg[58]) );
  DFFRHQX1 dout4_reg_reg_9_ ( .D(n1664), .CK(clk), .RN(rstn), .Q(dout4_reg[9])
         );
  DFFRHQX1 dout4_reg_reg_25_ ( .D(n1680), .CK(clk), .RN(rstn), .Q(
        dout4_reg[25]) );
  DFFRHQX1 dout4_reg_reg_41_ ( .D(n1696), .CK(clk), .RN(rstn), .Q(
        dout4_reg[41]) );
  DFFRHQX1 dout4_reg_reg_57_ ( .D(n1712), .CK(clk), .RN(rstn), .Q(
        dout4_reg[57]) );
  DFFRHQX1 dout4_reg_reg_8_ ( .D(n1663), .CK(clk), .RN(rstn), .Q(dout4_reg[8])
         );
  DFFRHQX1 dout4_reg_reg_24_ ( .D(n1679), .CK(clk), .RN(rstn), .Q(
        dout4_reg[24]) );
  DFFRHQX1 dout4_reg_reg_40_ ( .D(n1695), .CK(clk), .RN(rstn), .Q(
        dout4_reg[40]) );
  DFFRHQX1 dout4_reg_reg_56_ ( .D(n1711), .CK(clk), .RN(rstn), .Q(
        dout4_reg[56]) );
  DFFRHQX1 dout4_reg_reg_7_ ( .D(n1662), .CK(clk), .RN(rstn), .Q(dout4_reg[7])
         );
  DFFRHQX1 dout4_reg_reg_23_ ( .D(n1678), .CK(clk), .RN(rstn), .Q(
        dout4_reg[23]) );
  DFFRHQX1 dout4_reg_reg_39_ ( .D(n1694), .CK(clk), .RN(rstn), .Q(
        dout4_reg[39]) );
  DFFRHQX1 dout4_reg_reg_55_ ( .D(n1710), .CK(clk), .RN(rstn), .Q(
        dout4_reg[55]) );
  DFFRHQX1 dout4_reg_reg_6_ ( .D(n1661), .CK(clk), .RN(rstn), .Q(dout4_reg[6])
         );
  DFFRHQX1 dout4_reg_reg_22_ ( .D(n1677), .CK(clk), .RN(rstn), .Q(
        dout4_reg[22]) );
  DFFRHQX1 dout4_reg_reg_38_ ( .D(n1693), .CK(clk), .RN(rstn), .Q(
        dout4_reg[38]) );
  DFFRHQX1 dout4_reg_reg_54_ ( .D(n1709), .CK(clk), .RN(rstn), .Q(
        dout4_reg[54]) );
  DFFRHQX1 dout4_reg_reg_5_ ( .D(n1660), .CK(clk), .RN(rstn), .Q(dout4_reg[5])
         );
  DFFRHQX1 dout4_reg_reg_21_ ( .D(n1676), .CK(clk), .RN(rstn), .Q(
        dout4_reg[21]) );
  DFFRHQX1 dout4_reg_reg_37_ ( .D(n1692), .CK(clk), .RN(rstn), .Q(
        dout4_reg[37]) );
  DFFRHQX1 dout4_reg_reg_53_ ( .D(n1708), .CK(clk), .RN(rstn), .Q(
        dout4_reg[53]) );
  DFFRHQX1 dout4_reg_reg_4_ ( .D(n1659), .CK(clk), .RN(rstn), .Q(dout4_reg[4])
         );
  DFFRHQX1 dout4_reg_reg_20_ ( .D(n1675), .CK(clk), .RN(rstn), .Q(
        dout4_reg[20]) );
  DFFRHQX1 dout4_reg_reg_36_ ( .D(n1691), .CK(clk), .RN(rstn), .Q(
        dout4_reg[36]) );
  DFFRHQX1 dout4_reg_reg_52_ ( .D(n1707), .CK(clk), .RN(rstn), .Q(
        dout4_reg[52]) );
  DFFRHQX1 dout4_reg_reg_3_ ( .D(n1658), .CK(clk), .RN(rstn), .Q(dout4_reg[3])
         );
  DFFRHQX1 dout4_reg_reg_19_ ( .D(n1674), .CK(clk), .RN(rstn), .Q(
        dout4_reg[19]) );
  DFFRHQX1 dout4_reg_reg_35_ ( .D(n1690), .CK(clk), .RN(rstn), .Q(
        dout4_reg[35]) );
  DFFRHQX1 dout4_reg_reg_51_ ( .D(n1706), .CK(clk), .RN(rstn), .Q(
        dout4_reg[51]) );
  DFFRHQX1 dout4_reg_reg_2_ ( .D(n1657), .CK(clk), .RN(rstn), .Q(dout4_reg[2])
         );
  DFFRHQX1 dout4_reg_reg_18_ ( .D(n1673), .CK(clk), .RN(rstn), .Q(
        dout4_reg[18]) );
  DFFRHQX1 dout4_reg_reg_34_ ( .D(n1689), .CK(clk), .RN(rstn), .Q(
        dout4_reg[34]) );
  DFFRHQX1 dout4_reg_reg_50_ ( .D(n1705), .CK(clk), .RN(rstn), .Q(
        dout4_reg[50]) );
  DFFRHQX1 dout4_reg_reg_1_ ( .D(n1656), .CK(clk), .RN(rstn), .Q(dout4_reg[1])
         );
  DFFRHQX1 dout4_reg_reg_17_ ( .D(n1672), .CK(clk), .RN(rstn), .Q(
        dout4_reg[17]) );
  DFFRHQX1 dout4_reg_reg_33_ ( .D(n1688), .CK(clk), .RN(rstn), .Q(
        dout4_reg[33]) );
  DFFRHQX1 dout4_reg_reg_49_ ( .D(n1704), .CK(clk), .RN(rstn), .Q(
        dout4_reg[49]) );
  DFFRHQX1 dout4_reg_reg_0_ ( .D(n1655), .CK(clk), .RN(rstn), .Q(dout4_reg[0])
         );
  DFFRHQX1 dout4_reg_reg_16_ ( .D(n1671), .CK(clk), .RN(rstn), .Q(
        dout4_reg[16]) );
  DFFRHQX1 dout4_reg_reg_32_ ( .D(n1687), .CK(clk), .RN(rstn), .Q(
        dout4_reg[32]) );
  DFFRHQX1 dout4_reg_reg_48_ ( .D(n1703), .CK(clk), .RN(rstn), .Q(
        dout4_reg[48]) );
  DFFRHQX1 count_reg_4_ ( .D(N1118), .CK(clk), .RN(rstn), .Q(count[4]) );
  DFFRHQX1 dout16_reg_reg_15_ ( .D(n1286), .CK(clk), .RN(rstn), .Q(
        dout16_reg[15]) );
  DFFRHQX1 dout16_reg_reg_31_ ( .D(n1302), .CK(clk), .RN(rstn), .Q(
        dout16_reg[31]) );
  DFFRHQX1 dout16_reg_reg_47_ ( .D(n1318), .CK(clk), .RN(rstn), .Q(
        dout16_reg[47]) );
  DFFRHQX1 dout16_reg_reg_63_ ( .D(n1334), .CK(clk), .RN(rstn), .Q(
        dout16_reg[63]) );
  DFFRHQX1 dout16_reg_reg_79_ ( .D(n1350), .CK(clk), .RN(rstn), .Q(
        dout16_reg[79]) );
  DFFRHQX1 dout16_reg_reg_95_ ( .D(n1366), .CK(clk), .RN(rstn), .Q(
        dout16_reg[95]) );
  DFFRHQX1 dout16_reg_reg_111_ ( .D(n1382), .CK(clk), .RN(rstn), .Q(
        dout16_reg[111]) );
  DFFRHQX1 dout16_reg_reg_127_ ( .D(n1398), .CK(clk), .RN(rstn), .Q(
        dout16_reg[127]) );
  DFFRHQX1 dout16_reg_reg_143_ ( .D(n1414), .CK(clk), .RN(rstn), .Q(
        dout16_reg[143]) );
  DFFRHQX1 dout16_reg_reg_159_ ( .D(n1430), .CK(clk), .RN(rstn), .Q(
        dout16_reg[159]) );
  DFFRHQX1 dout16_reg_reg_175_ ( .D(n1446), .CK(clk), .RN(rstn), .Q(
        dout16_reg[175]) );
  DFFRHQX1 dout16_reg_reg_191_ ( .D(n1462), .CK(clk), .RN(rstn), .Q(
        dout16_reg[191]) );
  DFFRHQX1 dout16_reg_reg_14_ ( .D(n1285), .CK(clk), .RN(rstn), .Q(
        dout16_reg[14]) );
  DFFRHQX1 dout16_reg_reg_30_ ( .D(n1301), .CK(clk), .RN(rstn), .Q(
        dout16_reg[30]) );
  DFFRHQX1 dout16_reg_reg_46_ ( .D(n1317), .CK(clk), .RN(rstn), .Q(
        dout16_reg[46]) );
  DFFRHQX1 dout16_reg_reg_62_ ( .D(n1333), .CK(clk), .RN(rstn), .Q(
        dout16_reg[62]) );
  DFFRHQX1 dout16_reg_reg_78_ ( .D(n1349), .CK(clk), .RN(rstn), .Q(
        dout16_reg[78]) );
  DFFRHQX1 dout16_reg_reg_94_ ( .D(n1365), .CK(clk), .RN(rstn), .Q(
        dout16_reg[94]) );
  DFFRHQX1 dout16_reg_reg_110_ ( .D(n1381), .CK(clk), .RN(rstn), .Q(
        dout16_reg[110]) );
  DFFRHQX1 dout16_reg_reg_126_ ( .D(n1397), .CK(clk), .RN(rstn), .Q(
        dout16_reg[126]) );
  DFFRHQX1 dout16_reg_reg_142_ ( .D(n1413), .CK(clk), .RN(rstn), .Q(
        dout16_reg[142]) );
  DFFRHQX1 dout16_reg_reg_158_ ( .D(n1429), .CK(clk), .RN(rstn), .Q(
        dout16_reg[158]) );
  DFFRHQX1 dout16_reg_reg_174_ ( .D(n1445), .CK(clk), .RN(rstn), .Q(
        dout16_reg[174]) );
  DFFRHQX1 dout16_reg_reg_190_ ( .D(n1461), .CK(clk), .RN(rstn), .Q(
        dout16_reg[190]) );
  DFFRHQX1 dout16_reg_reg_13_ ( .D(n1284), .CK(clk), .RN(rstn), .Q(
        dout16_reg[13]) );
  DFFRHQX1 dout16_reg_reg_29_ ( .D(n1300), .CK(clk), .RN(rstn), .Q(
        dout16_reg[29]) );
  DFFRHQX1 dout16_reg_reg_45_ ( .D(n1316), .CK(clk), .RN(rstn), .Q(
        dout16_reg[45]) );
  DFFRHQX1 dout16_reg_reg_61_ ( .D(n1332), .CK(clk), .RN(rstn), .Q(
        dout16_reg[61]) );
  DFFRHQX1 dout16_reg_reg_77_ ( .D(n1348), .CK(clk), .RN(rstn), .Q(
        dout16_reg[77]) );
  DFFRHQX1 dout16_reg_reg_93_ ( .D(n1364), .CK(clk), .RN(rstn), .Q(
        dout16_reg[93]) );
  DFFRHQX1 dout16_reg_reg_109_ ( .D(n1380), .CK(clk), .RN(rstn), .Q(
        dout16_reg[109]) );
  DFFRHQX1 dout16_reg_reg_125_ ( .D(n1396), .CK(clk), .RN(rstn), .Q(
        dout16_reg[125]) );
  DFFRHQX1 dout16_reg_reg_141_ ( .D(n1412), .CK(clk), .RN(rstn), .Q(
        dout16_reg[141]) );
  DFFRHQX1 dout16_reg_reg_157_ ( .D(n1428), .CK(clk), .RN(rstn), .Q(
        dout16_reg[157]) );
  DFFRHQX1 dout16_reg_reg_173_ ( .D(n1444), .CK(clk), .RN(rstn), .Q(
        dout16_reg[173]) );
  DFFRHQX1 dout16_reg_reg_189_ ( .D(n1460), .CK(clk), .RN(rstn), .Q(
        dout16_reg[189]) );
  DFFRHQX1 dout16_reg_reg_12_ ( .D(n1283), .CK(clk), .RN(rstn), .Q(
        dout16_reg[12]) );
  DFFRHQX1 dout16_reg_reg_28_ ( .D(n1299), .CK(clk), .RN(rstn), .Q(
        dout16_reg[28]) );
  DFFRHQX1 dout16_reg_reg_44_ ( .D(n1315), .CK(clk), .RN(rstn), .Q(
        dout16_reg[44]) );
  DFFRHQX1 dout16_reg_reg_60_ ( .D(n1331), .CK(clk), .RN(rstn), .Q(
        dout16_reg[60]) );
  DFFRHQX1 dout16_reg_reg_76_ ( .D(n1347), .CK(clk), .RN(rstn), .Q(
        dout16_reg[76]) );
  DFFRHQX1 dout16_reg_reg_92_ ( .D(n1363), .CK(clk), .RN(rstn), .Q(
        dout16_reg[92]) );
  DFFRHQX1 dout16_reg_reg_108_ ( .D(n1379), .CK(clk), .RN(rstn), .Q(
        dout16_reg[108]) );
  DFFRHQX1 dout16_reg_reg_124_ ( .D(n1395), .CK(clk), .RN(rstn), .Q(
        dout16_reg[124]) );
  DFFRHQX1 dout16_reg_reg_140_ ( .D(n1411), .CK(clk), .RN(rstn), .Q(
        dout16_reg[140]) );
  DFFRHQX1 dout16_reg_reg_156_ ( .D(n1427), .CK(clk), .RN(rstn), .Q(
        dout16_reg[156]) );
  DFFRHQX1 dout16_reg_reg_172_ ( .D(n1443), .CK(clk), .RN(rstn), .Q(
        dout16_reg[172]) );
  DFFRHQX1 dout16_reg_reg_188_ ( .D(n1459), .CK(clk), .RN(rstn), .Q(
        dout16_reg[188]) );
  DFFRHQX1 dout16_reg_reg_11_ ( .D(n1282), .CK(clk), .RN(rstn), .Q(
        dout16_reg[11]) );
  DFFRHQX1 dout16_reg_reg_27_ ( .D(n1298), .CK(clk), .RN(rstn), .Q(
        dout16_reg[27]) );
  DFFRHQX1 dout16_reg_reg_43_ ( .D(n1314), .CK(clk), .RN(rstn), .Q(
        dout16_reg[43]) );
  DFFRHQX1 dout16_reg_reg_59_ ( .D(n1330), .CK(clk), .RN(rstn), .Q(
        dout16_reg[59]) );
  DFFRHQX1 dout16_reg_reg_75_ ( .D(n1346), .CK(clk), .RN(rstn), .Q(
        dout16_reg[75]) );
  DFFRHQX1 dout16_reg_reg_91_ ( .D(n1362), .CK(clk), .RN(rstn), .Q(
        dout16_reg[91]) );
  DFFRHQX1 dout16_reg_reg_107_ ( .D(n1378), .CK(clk), .RN(rstn), .Q(
        dout16_reg[107]) );
  DFFRHQX1 dout16_reg_reg_123_ ( .D(n1394), .CK(clk), .RN(rstn), .Q(
        dout16_reg[123]) );
  DFFRHQX1 dout16_reg_reg_139_ ( .D(n1410), .CK(clk), .RN(rstn), .Q(
        dout16_reg[139]) );
  DFFRHQX1 dout16_reg_reg_155_ ( .D(n1426), .CK(clk), .RN(rstn), .Q(
        dout16_reg[155]) );
  DFFRHQX1 dout16_reg_reg_171_ ( .D(n1442), .CK(clk), .RN(rstn), .Q(
        dout16_reg[171]) );
  DFFRHQX1 dout16_reg_reg_187_ ( .D(n1458), .CK(clk), .RN(rstn), .Q(
        dout16_reg[187]) );
  DFFRHQX1 dout16_reg_reg_10_ ( .D(n1281), .CK(clk), .RN(rstn), .Q(
        dout16_reg[10]) );
  DFFRHQX1 dout16_reg_reg_26_ ( .D(n1297), .CK(clk), .RN(rstn), .Q(
        dout16_reg[26]) );
  DFFRHQX1 dout16_reg_reg_42_ ( .D(n1313), .CK(clk), .RN(rstn), .Q(
        dout16_reg[42]) );
  DFFRHQX1 dout16_reg_reg_58_ ( .D(n1329), .CK(clk), .RN(rstn), .Q(
        dout16_reg[58]) );
  DFFRHQX1 dout16_reg_reg_74_ ( .D(n1345), .CK(clk), .RN(rstn), .Q(
        dout16_reg[74]) );
  DFFRHQX1 dout16_reg_reg_90_ ( .D(n1361), .CK(clk), .RN(rstn), .Q(
        dout16_reg[90]) );
  DFFRHQX1 dout16_reg_reg_106_ ( .D(n1377), .CK(clk), .RN(rstn), .Q(
        dout16_reg[106]) );
  DFFRHQX1 dout16_reg_reg_122_ ( .D(n1393), .CK(clk), .RN(rstn), .Q(
        dout16_reg[122]) );
  DFFRHQX1 dout16_reg_reg_138_ ( .D(n1409), .CK(clk), .RN(rstn), .Q(
        dout16_reg[138]) );
  DFFRHQX1 dout16_reg_reg_154_ ( .D(n1425), .CK(clk), .RN(rstn), .Q(
        dout16_reg[154]) );
  DFFRHQX1 dout16_reg_reg_170_ ( .D(n1441), .CK(clk), .RN(rstn), .Q(
        dout16_reg[170]) );
  DFFRHQX1 dout16_reg_reg_186_ ( .D(n1457), .CK(clk), .RN(rstn), .Q(
        dout16_reg[186]) );
  DFFRHQX1 dout16_reg_reg_9_ ( .D(n1280), .CK(clk), .RN(rstn), .Q(
        dout16_reg[9]) );
  DFFRHQX1 dout16_reg_reg_25_ ( .D(n1296), .CK(clk), .RN(rstn), .Q(
        dout16_reg[25]) );
  DFFRHQX1 dout16_reg_reg_41_ ( .D(n1312), .CK(clk), .RN(rstn), .Q(
        dout16_reg[41]) );
  DFFRHQX1 dout16_reg_reg_57_ ( .D(n1328), .CK(clk), .RN(rstn), .Q(
        dout16_reg[57]) );
  DFFRHQX1 dout16_reg_reg_73_ ( .D(n1344), .CK(clk), .RN(rstn), .Q(
        dout16_reg[73]) );
  DFFRHQX1 dout16_reg_reg_89_ ( .D(n1360), .CK(clk), .RN(rstn), .Q(
        dout16_reg[89]) );
  DFFRHQX1 dout16_reg_reg_105_ ( .D(n1376), .CK(clk), .RN(rstn), .Q(
        dout16_reg[105]) );
  DFFRHQX1 dout16_reg_reg_121_ ( .D(n1392), .CK(clk), .RN(rstn), .Q(
        dout16_reg[121]) );
  DFFRHQX1 dout16_reg_reg_137_ ( .D(n1408), .CK(clk), .RN(rstn), .Q(
        dout16_reg[137]) );
  DFFRHQX1 dout16_reg_reg_153_ ( .D(n1424), .CK(clk), .RN(rstn), .Q(
        dout16_reg[153]) );
  DFFRHQX1 dout16_reg_reg_169_ ( .D(n1440), .CK(clk), .RN(rstn), .Q(
        dout16_reg[169]) );
  DFFRHQX1 dout16_reg_reg_185_ ( .D(n1456), .CK(clk), .RN(rstn), .Q(
        dout16_reg[185]) );
  DFFRHQX1 dout16_reg_reg_8_ ( .D(n1279), .CK(clk), .RN(rstn), .Q(
        dout16_reg[8]) );
  DFFRHQX1 dout16_reg_reg_24_ ( .D(n1295), .CK(clk), .RN(rstn), .Q(
        dout16_reg[24]) );
  DFFRHQX1 dout16_reg_reg_40_ ( .D(n1311), .CK(clk), .RN(rstn), .Q(
        dout16_reg[40]) );
  DFFRHQX1 dout16_reg_reg_56_ ( .D(n1327), .CK(clk), .RN(rstn), .Q(
        dout16_reg[56]) );
  DFFRHQX1 dout16_reg_reg_72_ ( .D(n1343), .CK(clk), .RN(rstn), .Q(
        dout16_reg[72]) );
  DFFRHQX1 dout16_reg_reg_88_ ( .D(n1359), .CK(clk), .RN(rstn), .Q(
        dout16_reg[88]) );
  DFFRHQX1 dout16_reg_reg_104_ ( .D(n1375), .CK(clk), .RN(rstn), .Q(
        dout16_reg[104]) );
  DFFRHQX1 dout16_reg_reg_120_ ( .D(n1391), .CK(clk), .RN(rstn), .Q(
        dout16_reg[120]) );
  DFFRHQX1 dout16_reg_reg_136_ ( .D(n1407), .CK(clk), .RN(rstn), .Q(
        dout16_reg[136]) );
  DFFRHQX1 dout16_reg_reg_152_ ( .D(n1423), .CK(clk), .RN(rstn), .Q(
        dout16_reg[152]) );
  DFFRHQX1 dout16_reg_reg_168_ ( .D(n1439), .CK(clk), .RN(rstn), .Q(
        dout16_reg[168]) );
  DFFRHQX1 dout16_reg_reg_184_ ( .D(n1455), .CK(clk), .RN(rstn), .Q(
        dout16_reg[184]) );
  DFFRHQX1 dout16_reg_reg_7_ ( .D(n1278), .CK(clk), .RN(rstn), .Q(
        dout16_reg[7]) );
  DFFRHQX1 dout16_reg_reg_23_ ( .D(n1294), .CK(clk), .RN(rstn), .Q(
        dout16_reg[23]) );
  DFFRHQX1 dout16_reg_reg_39_ ( .D(n1310), .CK(clk), .RN(rstn), .Q(
        dout16_reg[39]) );
  DFFRHQX1 dout16_reg_reg_55_ ( .D(n1326), .CK(clk), .RN(rstn), .Q(
        dout16_reg[55]) );
  DFFRHQX1 dout16_reg_reg_71_ ( .D(n1342), .CK(clk), .RN(rstn), .Q(
        dout16_reg[71]) );
  DFFRHQX1 dout16_reg_reg_87_ ( .D(n1358), .CK(clk), .RN(rstn), .Q(
        dout16_reg[87]) );
  DFFRHQX1 dout16_reg_reg_103_ ( .D(n1374), .CK(clk), .RN(rstn), .Q(
        dout16_reg[103]) );
  DFFRHQX1 dout16_reg_reg_119_ ( .D(n1390), .CK(clk), .RN(rstn), .Q(
        dout16_reg[119]) );
  DFFRHQX1 dout16_reg_reg_135_ ( .D(n1406), .CK(clk), .RN(rstn), .Q(
        dout16_reg[135]) );
  DFFRHQX1 dout16_reg_reg_151_ ( .D(n1422), .CK(clk), .RN(rstn), .Q(
        dout16_reg[151]) );
  DFFRHQX1 dout16_reg_reg_167_ ( .D(n1438), .CK(clk), .RN(rstn), .Q(
        dout16_reg[167]) );
  DFFRHQX1 dout16_reg_reg_183_ ( .D(n1454), .CK(clk), .RN(rstn), .Q(
        dout16_reg[183]) );
  DFFRHQX1 dout16_reg_reg_6_ ( .D(n1277), .CK(clk), .RN(rstn), .Q(
        dout16_reg[6]) );
  DFFRHQX1 dout16_reg_reg_22_ ( .D(n1293), .CK(clk), .RN(rstn), .Q(
        dout16_reg[22]) );
  DFFRHQX1 dout16_reg_reg_38_ ( .D(n1309), .CK(clk), .RN(rstn), .Q(
        dout16_reg[38]) );
  DFFRHQX1 dout16_reg_reg_54_ ( .D(n1325), .CK(clk), .RN(rstn), .Q(
        dout16_reg[54]) );
  DFFRHQX1 dout16_reg_reg_70_ ( .D(n1341), .CK(clk), .RN(rstn), .Q(
        dout16_reg[70]) );
  DFFRHQX1 dout16_reg_reg_86_ ( .D(n1357), .CK(clk), .RN(rstn), .Q(
        dout16_reg[86]) );
  DFFRHQX1 dout16_reg_reg_102_ ( .D(n1373), .CK(clk), .RN(rstn), .Q(
        dout16_reg[102]) );
  DFFRHQX1 dout16_reg_reg_118_ ( .D(n1389), .CK(clk), .RN(rstn), .Q(
        dout16_reg[118]) );
  DFFRHQX1 dout16_reg_reg_134_ ( .D(n1405), .CK(clk), .RN(rstn), .Q(
        dout16_reg[134]) );
  DFFRHQX1 dout16_reg_reg_150_ ( .D(n1421), .CK(clk), .RN(rstn), .Q(
        dout16_reg[150]) );
  DFFRHQX1 dout16_reg_reg_166_ ( .D(n1437), .CK(clk), .RN(rstn), .Q(
        dout16_reg[166]) );
  DFFRHQX1 dout16_reg_reg_182_ ( .D(n1453), .CK(clk), .RN(rstn), .Q(
        dout16_reg[182]) );
  DFFRHQX1 dout16_reg_reg_5_ ( .D(n1276), .CK(clk), .RN(rstn), .Q(
        dout16_reg[5]) );
  DFFRHQX1 dout16_reg_reg_21_ ( .D(n1292), .CK(clk), .RN(rstn), .Q(
        dout16_reg[21]) );
  DFFRHQX1 dout16_reg_reg_37_ ( .D(n1308), .CK(clk), .RN(rstn), .Q(
        dout16_reg[37]) );
  DFFRHQX1 dout16_reg_reg_53_ ( .D(n1324), .CK(clk), .RN(rstn), .Q(
        dout16_reg[53]) );
  DFFRHQX1 dout16_reg_reg_69_ ( .D(n1340), .CK(clk), .RN(rstn), .Q(
        dout16_reg[69]) );
  DFFRHQX1 dout16_reg_reg_85_ ( .D(n1356), .CK(clk), .RN(rstn), .Q(
        dout16_reg[85]) );
  DFFRHQX1 dout16_reg_reg_101_ ( .D(n1372), .CK(clk), .RN(rstn), .Q(
        dout16_reg[101]) );
  DFFRHQX1 dout16_reg_reg_117_ ( .D(n1388), .CK(clk), .RN(rstn), .Q(
        dout16_reg[117]) );
  DFFRHQX1 dout16_reg_reg_133_ ( .D(n1404), .CK(clk), .RN(rstn), .Q(
        dout16_reg[133]) );
  DFFRHQX1 dout16_reg_reg_149_ ( .D(n1420), .CK(clk), .RN(rstn), .Q(
        dout16_reg[149]) );
  DFFRHQX1 dout16_reg_reg_165_ ( .D(n1436), .CK(clk), .RN(rstn), .Q(
        dout16_reg[165]) );
  DFFRHQX1 dout16_reg_reg_181_ ( .D(n1452), .CK(clk), .RN(rstn), .Q(
        dout16_reg[181]) );
  DFFRHQX1 dout16_reg_reg_4_ ( .D(n1275), .CK(clk), .RN(rstn), .Q(
        dout16_reg[4]) );
  DFFRHQX1 dout16_reg_reg_20_ ( .D(n1291), .CK(clk), .RN(rstn), .Q(
        dout16_reg[20]) );
  DFFRHQX1 dout16_reg_reg_36_ ( .D(n1307), .CK(clk), .RN(rstn), .Q(
        dout16_reg[36]) );
  DFFRHQX1 dout16_reg_reg_52_ ( .D(n1323), .CK(clk), .RN(rstn), .Q(
        dout16_reg[52]) );
  DFFRHQX1 dout16_reg_reg_68_ ( .D(n1339), .CK(clk), .RN(rstn), .Q(
        dout16_reg[68]) );
  DFFRHQX1 dout16_reg_reg_84_ ( .D(n1355), .CK(clk), .RN(rstn), .Q(
        dout16_reg[84]) );
  DFFRHQX1 dout16_reg_reg_100_ ( .D(n1371), .CK(clk), .RN(rstn), .Q(
        dout16_reg[100]) );
  DFFRHQX1 dout16_reg_reg_116_ ( .D(n1387), .CK(clk), .RN(rstn), .Q(
        dout16_reg[116]) );
  DFFRHQX1 dout16_reg_reg_132_ ( .D(n1403), .CK(clk), .RN(rstn), .Q(
        dout16_reg[132]) );
  DFFRHQX1 dout16_reg_reg_148_ ( .D(n1419), .CK(clk), .RN(rstn), .Q(
        dout16_reg[148]) );
  DFFRHQX1 dout16_reg_reg_164_ ( .D(n1435), .CK(clk), .RN(rstn), .Q(
        dout16_reg[164]) );
  DFFRHQX1 dout16_reg_reg_180_ ( .D(n1451), .CK(clk), .RN(rstn), .Q(
        dout16_reg[180]) );
  DFFRHQX1 dout16_reg_reg_3_ ( .D(n1274), .CK(clk), .RN(rstn), .Q(
        dout16_reg[3]) );
  DFFRHQX1 dout16_reg_reg_19_ ( .D(n1290), .CK(clk), .RN(rstn), .Q(
        dout16_reg[19]) );
  DFFRHQX1 dout16_reg_reg_35_ ( .D(n1306), .CK(clk), .RN(rstn), .Q(
        dout16_reg[35]) );
  DFFRHQX1 dout16_reg_reg_51_ ( .D(n1322), .CK(clk), .RN(rstn), .Q(
        dout16_reg[51]) );
  DFFRHQX1 dout16_reg_reg_67_ ( .D(n1338), .CK(clk), .RN(rstn), .Q(
        dout16_reg[67]) );
  DFFRHQX1 dout16_reg_reg_83_ ( .D(n1354), .CK(clk), .RN(rstn), .Q(
        dout16_reg[83]) );
  DFFRHQX1 dout16_reg_reg_99_ ( .D(n1370), .CK(clk), .RN(rstn), .Q(
        dout16_reg[99]) );
  DFFRHQX1 dout16_reg_reg_115_ ( .D(n1386), .CK(clk), .RN(rstn), .Q(
        dout16_reg[115]) );
  DFFRHQX1 dout16_reg_reg_131_ ( .D(n1402), .CK(clk), .RN(rstn), .Q(
        dout16_reg[131]) );
  DFFRHQX1 dout16_reg_reg_147_ ( .D(n1418), .CK(clk), .RN(rstn), .Q(
        dout16_reg[147]) );
  DFFRHQX1 dout16_reg_reg_163_ ( .D(n1434), .CK(clk), .RN(rstn), .Q(
        dout16_reg[163]) );
  DFFRHQX1 dout16_reg_reg_179_ ( .D(n1450), .CK(clk), .RN(rstn), .Q(
        dout16_reg[179]) );
  DFFRHQX1 dout16_reg_reg_2_ ( .D(n1273), .CK(clk), .RN(rstn), .Q(
        dout16_reg[2]) );
  DFFRHQX1 dout16_reg_reg_18_ ( .D(n1289), .CK(clk), .RN(rstn), .Q(
        dout16_reg[18]) );
  DFFRHQX1 dout16_reg_reg_34_ ( .D(n1305), .CK(clk), .RN(rstn), .Q(
        dout16_reg[34]) );
  DFFRHQX1 dout16_reg_reg_50_ ( .D(n1321), .CK(clk), .RN(rstn), .Q(
        dout16_reg[50]) );
  DFFRHQX1 dout16_reg_reg_66_ ( .D(n1337), .CK(clk), .RN(rstn), .Q(
        dout16_reg[66]) );
  DFFRHQX1 dout16_reg_reg_82_ ( .D(n1353), .CK(clk), .RN(rstn), .Q(
        dout16_reg[82]) );
  DFFRHQX1 dout16_reg_reg_98_ ( .D(n1369), .CK(clk), .RN(rstn), .Q(
        dout16_reg[98]) );
  DFFRHQX1 dout16_reg_reg_114_ ( .D(n1385), .CK(clk), .RN(rstn), .Q(
        dout16_reg[114]) );
  DFFRHQX1 dout16_reg_reg_130_ ( .D(n1401), .CK(clk), .RN(rstn), .Q(
        dout16_reg[130]) );
  DFFRHQX1 dout16_reg_reg_146_ ( .D(n1417), .CK(clk), .RN(rstn), .Q(
        dout16_reg[146]) );
  DFFRHQX1 dout16_reg_reg_162_ ( .D(n1433), .CK(clk), .RN(rstn), .Q(
        dout16_reg[162]) );
  DFFRHQX1 dout16_reg_reg_178_ ( .D(n1449), .CK(clk), .RN(rstn), .Q(
        dout16_reg[178]) );
  DFFRHQX1 dout16_reg_reg_1_ ( .D(n1272), .CK(clk), .RN(rstn), .Q(
        dout16_reg[1]) );
  DFFRHQX1 dout16_reg_reg_17_ ( .D(n1288), .CK(clk), .RN(rstn), .Q(
        dout16_reg[17]) );
  DFFRHQX1 dout16_reg_reg_33_ ( .D(n1304), .CK(clk), .RN(rstn), .Q(
        dout16_reg[33]) );
  DFFRHQX1 dout16_reg_reg_49_ ( .D(n1320), .CK(clk), .RN(rstn), .Q(
        dout16_reg[49]) );
  DFFRHQX1 dout16_reg_reg_65_ ( .D(n1336), .CK(clk), .RN(rstn), .Q(
        dout16_reg[65]) );
  DFFRHQX1 dout16_reg_reg_81_ ( .D(n1352), .CK(clk), .RN(rstn), .Q(
        dout16_reg[81]) );
  DFFRHQX1 dout16_reg_reg_97_ ( .D(n1368), .CK(clk), .RN(rstn), .Q(
        dout16_reg[97]) );
  DFFRHQX1 dout16_reg_reg_113_ ( .D(n1384), .CK(clk), .RN(rstn), .Q(
        dout16_reg[113]) );
  DFFRHQX1 dout16_reg_reg_129_ ( .D(n1400), .CK(clk), .RN(rstn), .Q(
        dout16_reg[129]) );
  DFFRHQX1 dout16_reg_reg_145_ ( .D(n1416), .CK(clk), .RN(rstn), .Q(
        dout16_reg[145]) );
  DFFRHQX1 dout16_reg_reg_161_ ( .D(n1432), .CK(clk), .RN(rstn), .Q(
        dout16_reg[161]) );
  DFFRHQX1 dout16_reg_reg_177_ ( .D(n1448), .CK(clk), .RN(rstn), .Q(
        dout16_reg[177]) );
  DFFRHQX1 dout16_reg_reg_0_ ( .D(n1271), .CK(clk), .RN(rstn), .Q(
        dout16_reg[0]) );
  DFFRHQX1 dout16_reg_reg_16_ ( .D(n1287), .CK(clk), .RN(rstn), .Q(
        dout16_reg[16]) );
  DFFRHQX1 dout16_reg_reg_32_ ( .D(n1303), .CK(clk), .RN(rstn), .Q(
        dout16_reg[32]) );
  DFFRHQX1 dout16_reg_reg_48_ ( .D(n1319), .CK(clk), .RN(rstn), .Q(
        dout16_reg[48]) );
  DFFRHQX1 dout16_reg_reg_64_ ( .D(n1335), .CK(clk), .RN(rstn), .Q(
        dout16_reg[64]) );
  DFFRHQX1 dout16_reg_reg_80_ ( .D(n1351), .CK(clk), .RN(rstn), .Q(
        dout16_reg[80]) );
  DFFRHQX1 dout16_reg_reg_96_ ( .D(n1367), .CK(clk), .RN(rstn), .Q(
        dout16_reg[96]) );
  DFFRHQX1 dout16_reg_reg_112_ ( .D(n1383), .CK(clk), .RN(rstn), .Q(
        dout16_reg[112]) );
  DFFRHQX1 dout16_reg_reg_128_ ( .D(n1399), .CK(clk), .RN(rstn), .Q(
        dout16_reg[128]) );
  DFFRHQX1 dout16_reg_reg_144_ ( .D(n1415), .CK(clk), .RN(rstn), .Q(
        dout16_reg[144]) );
  DFFRHQX1 dout16_reg_reg_160_ ( .D(n1431), .CK(clk), .RN(rstn), .Q(
        dout16_reg[160]) );
  DFFRHQX1 dout16_reg_reg_176_ ( .D(n1447), .CK(clk), .RN(rstn), .Q(
        dout16_reg[176]) );
  DFFRHQX1 dout8_reg_reg_15_ ( .D(n1542), .CK(clk), .RN(rstn), .Q(
        dout8_reg[15]) );
  DFFRHQX1 dout8_reg_reg_31_ ( .D(n1558), .CK(clk), .RN(rstn), .Q(
        dout8_reg[31]) );
  DFFRHQX1 dout8_reg_reg_47_ ( .D(n1574), .CK(clk), .RN(rstn), .Q(
        dout8_reg[47]) );
  DFFRHQX1 dout8_reg_reg_63_ ( .D(n1590), .CK(clk), .RN(rstn), .Q(
        dout8_reg[63]) );
  DFFRHQX1 dout8_reg_reg_14_ ( .D(n1541), .CK(clk), .RN(rstn), .Q(
        dout8_reg[14]) );
  DFFRHQX1 dout8_reg_reg_30_ ( .D(n1557), .CK(clk), .RN(rstn), .Q(
        dout8_reg[30]) );
  DFFRHQX1 dout8_reg_reg_46_ ( .D(n1573), .CK(clk), .RN(rstn), .Q(
        dout8_reg[46]) );
  DFFRHQX1 dout8_reg_reg_62_ ( .D(n1589), .CK(clk), .RN(rstn), .Q(
        dout8_reg[62]) );
  DFFRHQX1 dout8_reg_reg_13_ ( .D(n1540), .CK(clk), .RN(rstn), .Q(
        dout8_reg[13]) );
  DFFRHQX1 dout8_reg_reg_29_ ( .D(n1556), .CK(clk), .RN(rstn), .Q(
        dout8_reg[29]) );
  DFFRHQX1 dout8_reg_reg_45_ ( .D(n1572), .CK(clk), .RN(rstn), .Q(
        dout8_reg[45]) );
  DFFRHQX1 dout8_reg_reg_61_ ( .D(n1588), .CK(clk), .RN(rstn), .Q(
        dout8_reg[61]) );
  DFFRHQX1 dout8_reg_reg_12_ ( .D(n1539), .CK(clk), .RN(rstn), .Q(
        dout8_reg[12]) );
  DFFRHQX1 dout8_reg_reg_28_ ( .D(n1555), .CK(clk), .RN(rstn), .Q(
        dout8_reg[28]) );
  DFFRHQX1 dout8_reg_reg_44_ ( .D(n1571), .CK(clk), .RN(rstn), .Q(
        dout8_reg[44]) );
  DFFRHQX1 dout8_reg_reg_60_ ( .D(n1587), .CK(clk), .RN(rstn), .Q(
        dout8_reg[60]) );
  DFFRHQX1 dout8_reg_reg_11_ ( .D(n1538), .CK(clk), .RN(rstn), .Q(
        dout8_reg[11]) );
  DFFRHQX1 dout8_reg_reg_27_ ( .D(n1554), .CK(clk), .RN(rstn), .Q(
        dout8_reg[27]) );
  DFFRHQX1 dout8_reg_reg_43_ ( .D(n1570), .CK(clk), .RN(rstn), .Q(
        dout8_reg[43]) );
  DFFRHQX1 dout8_reg_reg_59_ ( .D(n1586), .CK(clk), .RN(rstn), .Q(
        dout8_reg[59]) );
  DFFRHQX1 dout8_reg_reg_10_ ( .D(n1537), .CK(clk), .RN(rstn), .Q(
        dout8_reg[10]) );
  DFFRHQX1 dout8_reg_reg_26_ ( .D(n1553), .CK(clk), .RN(rstn), .Q(
        dout8_reg[26]) );
  DFFRHQX1 dout8_reg_reg_42_ ( .D(n1569), .CK(clk), .RN(rstn), .Q(
        dout8_reg[42]) );
  DFFRHQX1 dout8_reg_reg_58_ ( .D(n1585), .CK(clk), .RN(rstn), .Q(
        dout8_reg[58]) );
  DFFRHQX1 dout8_reg_reg_9_ ( .D(n1536), .CK(clk), .RN(rstn), .Q(dout8_reg[9])
         );
  DFFRHQX1 dout8_reg_reg_25_ ( .D(n1552), .CK(clk), .RN(rstn), .Q(
        dout8_reg[25]) );
  DFFRHQX1 dout8_reg_reg_41_ ( .D(n1568), .CK(clk), .RN(rstn), .Q(
        dout8_reg[41]) );
  DFFRHQX1 dout8_reg_reg_57_ ( .D(n1584), .CK(clk), .RN(rstn), .Q(
        dout8_reg[57]) );
  DFFRHQX1 dout8_reg_reg_8_ ( .D(n1535), .CK(clk), .RN(rstn), .Q(dout8_reg[8])
         );
  DFFRHQX1 dout8_reg_reg_24_ ( .D(n1551), .CK(clk), .RN(rstn), .Q(
        dout8_reg[24]) );
  DFFRHQX1 dout8_reg_reg_40_ ( .D(n1567), .CK(clk), .RN(rstn), .Q(
        dout8_reg[40]) );
  DFFRHQX1 dout8_reg_reg_56_ ( .D(n1583), .CK(clk), .RN(rstn), .Q(
        dout8_reg[56]) );
  DFFRHQX1 dout8_reg_reg_7_ ( .D(n1534), .CK(clk), .RN(rstn), .Q(dout8_reg[7])
         );
  DFFRHQX1 dout8_reg_reg_23_ ( .D(n1550), .CK(clk), .RN(rstn), .Q(
        dout8_reg[23]) );
  DFFRHQX1 dout8_reg_reg_39_ ( .D(n1566), .CK(clk), .RN(rstn), .Q(
        dout8_reg[39]) );
  DFFRHQX1 dout8_reg_reg_55_ ( .D(n1582), .CK(clk), .RN(rstn), .Q(
        dout8_reg[55]) );
  DFFRHQX1 dout8_reg_reg_6_ ( .D(n1533), .CK(clk), .RN(rstn), .Q(dout8_reg[6])
         );
  DFFRHQX1 dout8_reg_reg_22_ ( .D(n1549), .CK(clk), .RN(rstn), .Q(
        dout8_reg[22]) );
  DFFRHQX1 dout8_reg_reg_38_ ( .D(n1565), .CK(clk), .RN(rstn), .Q(
        dout8_reg[38]) );
  DFFRHQX1 dout8_reg_reg_54_ ( .D(n1581), .CK(clk), .RN(rstn), .Q(
        dout8_reg[54]) );
  DFFRHQX1 dout8_reg_reg_5_ ( .D(n1532), .CK(clk), .RN(rstn), .Q(dout8_reg[5])
         );
  DFFRHQX1 dout8_reg_reg_21_ ( .D(n1548), .CK(clk), .RN(rstn), .Q(
        dout8_reg[21]) );
  DFFRHQX1 dout8_reg_reg_37_ ( .D(n1564), .CK(clk), .RN(rstn), .Q(
        dout8_reg[37]) );
  DFFRHQX1 dout8_reg_reg_53_ ( .D(n1580), .CK(clk), .RN(rstn), .Q(
        dout8_reg[53]) );
  DFFRHQX1 dout8_reg_reg_4_ ( .D(n1531), .CK(clk), .RN(rstn), .Q(dout8_reg[4])
         );
  DFFRHQX1 dout8_reg_reg_20_ ( .D(n1547), .CK(clk), .RN(rstn), .Q(
        dout8_reg[20]) );
  DFFRHQX1 dout8_reg_reg_36_ ( .D(n1563), .CK(clk), .RN(rstn), .Q(
        dout8_reg[36]) );
  DFFRHQX1 dout8_reg_reg_52_ ( .D(n1579), .CK(clk), .RN(rstn), .Q(
        dout8_reg[52]) );
  DFFRHQX1 dout8_reg_reg_3_ ( .D(n1530), .CK(clk), .RN(rstn), .Q(dout8_reg[3])
         );
  DFFRHQX1 dout8_reg_reg_19_ ( .D(n1546), .CK(clk), .RN(rstn), .Q(
        dout8_reg[19]) );
  DFFRHQX1 dout8_reg_reg_35_ ( .D(n1562), .CK(clk), .RN(rstn), .Q(
        dout8_reg[35]) );
  DFFRHQX1 dout8_reg_reg_51_ ( .D(n1578), .CK(clk), .RN(rstn), .Q(
        dout8_reg[51]) );
  DFFRHQX1 dout8_reg_reg_2_ ( .D(n1529), .CK(clk), .RN(rstn), .Q(dout8_reg[2])
         );
  DFFRHQX1 dout8_reg_reg_18_ ( .D(n1545), .CK(clk), .RN(rstn), .Q(
        dout8_reg[18]) );
  DFFRHQX1 dout8_reg_reg_34_ ( .D(n1561), .CK(clk), .RN(rstn), .Q(
        dout8_reg[34]) );
  DFFRHQX1 dout8_reg_reg_50_ ( .D(n1577), .CK(clk), .RN(rstn), .Q(
        dout8_reg[50]) );
  DFFRHQX1 dout8_reg_reg_1_ ( .D(n1528), .CK(clk), .RN(rstn), .Q(dout8_reg[1])
         );
  DFFRHQX1 dout8_reg_reg_17_ ( .D(n1544), .CK(clk), .RN(rstn), .Q(
        dout8_reg[17]) );
  DFFRHQX1 dout8_reg_reg_33_ ( .D(n1560), .CK(clk), .RN(rstn), .Q(
        dout8_reg[33]) );
  DFFRHQX1 dout8_reg_reg_49_ ( .D(n1576), .CK(clk), .RN(rstn), .Q(
        dout8_reg[49]) );
  DFFRHQX1 dout8_reg_reg_0_ ( .D(n1527), .CK(clk), .RN(rstn), .Q(dout8_reg[0])
         );
  DFFRHQX1 dout8_reg_reg_16_ ( .D(n1543), .CK(clk), .RN(rstn), .Q(
        dout8_reg[16]) );
  DFFRHQX1 dout8_reg_reg_32_ ( .D(n1559), .CK(clk), .RN(rstn), .Q(
        dout8_reg[32]) );
  DFFRHQX1 dout8_reg_reg_48_ ( .D(n1575), .CK(clk), .RN(rstn), .Q(
        dout8_reg[48]) );
  DFFRHQX1 count_reg_0_ ( .D(N1114), .CK(clk), .RN(rstn), .Q(count[0]) );
  DFFRHQX1 count_reg_1_ ( .D(N1115), .CK(clk), .RN(rstn), .Q(count[1]) );
  DFFRHQX1 count_reg_3_ ( .D(N1117), .CK(clk), .RN(rstn), .Q(count[3]) );
  DFFRHQX1 count_reg_2_ ( .D(N1116), .CK(clk), .RN(rstn), .Q(count[2]) );
  DFFRHQX1 mode_reg_reg_0_ ( .D(mode[0]), .CK(clk), .RN(rstn), .Q(mode_reg[0])
         );
  DFFRHQX1 s2p_ready_reg ( .D(N1119), .CK(clk), .RN(rstn), .Q(s2p_ready) );
  DFFRXL mode_reg_reg_1_ ( .D(mode[1]), .CK(clk), .RN(rstn), .Q(mode_reg[1]), 
        .QN(n348) );
  AND2X2 U5 ( .A(n1730), .B(n1268), .Y(n1) );
  AND2X2 U6 ( .A(n1729), .B(start), .Y(n2) );
  AND2X2 U7 ( .A(start), .B(n1734), .Y(n3) );
  INVX1 U8 ( .A(n3), .Y(n313) );
  INVX1 U9 ( .A(n3), .Y(n314) );
  INVX1 U10 ( .A(n307), .Y(n303) );
  INVX1 U11 ( .A(n307), .Y(n304) );
  INVX1 U12 ( .A(n307), .Y(n305) );
  INVX1 U13 ( .A(n307), .Y(n306) );
  INVX1 U14 ( .A(n2), .Y(n284) );
  INVX1 U15 ( .A(n2), .Y(n280) );
  INVX1 U16 ( .A(n2), .Y(n278) );
  INVX1 U17 ( .A(n2), .Y(n279) );
  INVX1 U18 ( .A(n2), .Y(n281) );
  INVX1 U19 ( .A(n2), .Y(n282) );
  INVX1 U20 ( .A(n2), .Y(n283) );
  INVX1 U21 ( .A(n2), .Y(n285) );
  INVX1 U22 ( .A(n2), .Y(n286) );
  INVX1 U23 ( .A(n2), .Y(n287) );
  INVX1 U24 ( .A(n2), .Y(n288) );
  INVX1 U25 ( .A(n317), .Y(n315) );
  INVX1 U26 ( .A(n317), .Y(n316) );
  INVX1 U27 ( .A(n312), .Y(n310) );
  INVX1 U28 ( .A(n312), .Y(n308) );
  INVX1 U29 ( .A(n312), .Y(n309) );
  INVX1 U30 ( .A(n312), .Y(n311) );
  INVX1 U31 ( .A(n1), .Y(n293) );
  INVX1 U32 ( .A(n1), .Y(n302) );
  INVX1 U33 ( .A(n1), .Y(n296) );
  INVX1 U34 ( .A(n1), .Y(n294) );
  INVX1 U35 ( .A(n1), .Y(n292) );
  INVX1 U36 ( .A(n1), .Y(n291) );
  INVX1 U37 ( .A(n1), .Y(n290) );
  INVX1 U38 ( .A(n1), .Y(n301) );
  INVX1 U39 ( .A(n1), .Y(n300) );
  INVX1 U40 ( .A(n1), .Y(n299) );
  INVX1 U41 ( .A(n1), .Y(n298) );
  INVX1 U42 ( .A(n1), .Y(n297) );
  INVX1 U43 ( .A(n1), .Y(n295) );
  INVX1 U44 ( .A(n268), .Y(n266) );
  INVX1 U45 ( .A(n268), .Y(n267) );
  INVX1 U46 ( .A(n331), .Y(n319) );
  INVX1 U47 ( .A(n331), .Y(n320) );
  INVX1 U48 ( .A(n331), .Y(n321) );
  INVX1 U49 ( .A(n331), .Y(n322) );
  INVX1 U50 ( .A(n331), .Y(n323) );
  INVX1 U51 ( .A(n331), .Y(n324) );
  INVX1 U52 ( .A(n331), .Y(n325) );
  INVX1 U53 ( .A(n331), .Y(n326) );
  INVX1 U54 ( .A(n331), .Y(n327) );
  INVX1 U55 ( .A(n331), .Y(n328) );
  INVX1 U56 ( .A(n331), .Y(n329) );
  INVX1 U57 ( .A(n331), .Y(n330) );
  INVX1 U58 ( .A(n1), .Y(n289) );
  INVX1 U59 ( .A(start), .Y(n1265) );
  INVX1 U60 ( .A(n1735), .Y(n317) );
  INVX1 U61 ( .A(n1733), .Y(n312) );
  INVX1 U62 ( .A(n1732), .Y(n307) );
  INVX1 U63 ( .A(n277), .Y(n270) );
  INVX1 U64 ( .A(n277), .Y(n269) );
  INVX1 U65 ( .A(n277), .Y(n271) );
  INVX1 U66 ( .A(n277), .Y(n272) );
  INVX1 U67 ( .A(n277), .Y(n273) );
  INVX1 U68 ( .A(n277), .Y(n276) );
  INVX1 U69 ( .A(n277), .Y(n275) );
  INVX1 U70 ( .A(n265), .Y(n264) );
  INVX1 U71 ( .A(n277), .Y(n274) );
  INVX1 U72 ( .A(n265), .Y(n261) );
  INVX1 U73 ( .A(n265), .Y(n263) );
  INVX1 U74 ( .A(n265), .Y(n262) );
  INVX1 U75 ( .A(n331), .Y(n318) );
  INVX1 U76 ( .A(N30), .Y(n331) );
  INVX1 U77 ( .A(n1727), .Y(n268) );
  OAI22X1 U78 ( .A0(n1733), .A1(n640), .B0(n336), .B1(n1732), .Y(n1538) );
  OAI22X1 U79 ( .A0(n1733), .A1(n632), .B0(n335), .B1(n1732), .Y(n1539) );
  OAI22X1 U80 ( .A0(n1733), .A1(n624), .B0(n334), .B1(n1732), .Y(n1540) );
  OAI22X1 U81 ( .A0(n1733), .A1(n616), .B0(n333), .B1(n1732), .Y(n1541) );
  OAI22X1 U82 ( .A0(n1733), .A1(n608), .B0(n332), .B1(n1732), .Y(n1542) );
  OAI22X1 U83 ( .A0(n295), .A1(n448), .B0(n338), .B1(n286), .Y(n1280) );
  OAI22X1 U84 ( .A0(n295), .A1(n432), .B0(n337), .B1(n282), .Y(n1281) );
  OAI22X1 U85 ( .A0(n295), .A1(n416), .B0(n336), .B1(n286), .Y(n1282) );
  OAI22X1 U86 ( .A0(n295), .A1(n400), .B0(n335), .B1(n282), .Y(n1283) );
  OAI22X1 U87 ( .A0(n295), .A1(n384), .B0(n334), .B1(n288), .Y(n1284) );
  OAI22X1 U88 ( .A0(n295), .A1(n368), .B0(n333), .B1(n285), .Y(n1285) );
  OAI22X1 U89 ( .A0(n295), .A1(n352), .B0(n332), .B1(n286), .Y(n1286) );
  OAI22X1 U90 ( .A0(n315), .A1(n1261), .B0(n313), .B1(n347), .Y(n1655) );
  OAI22X1 U91 ( .A0(n1735), .A1(n1257), .B0(n313), .B1(n346), .Y(n1656) );
  OAI22X1 U92 ( .A0(n316), .A1(n1253), .B0(n313), .B1(n345), .Y(n1657) );
  OAI22X1 U93 ( .A0(n315), .A1(n1249), .B0(n313), .B1(n344), .Y(n1658) );
  OAI22X1 U94 ( .A0(n315), .A1(n1245), .B0(n313), .B1(n343), .Y(n1659) );
  OAI22X1 U95 ( .A0(n315), .A1(n1241), .B0(n313), .B1(n342), .Y(n1660) );
  OAI22X1 U96 ( .A0(n316), .A1(n1237), .B0(n313), .B1(n341), .Y(n1661) );
  OAI22X1 U97 ( .A0(n315), .A1(n1233), .B0(n313), .B1(n340), .Y(n1662) );
  OAI22X1 U98 ( .A0(n316), .A1(n1229), .B0(n313), .B1(n339), .Y(n1663) );
  OAI22X1 U99 ( .A0(n316), .A1(n1225), .B0(n313), .B1(n338), .Y(n1664) );
  OAI22X1 U100 ( .A0(n1735), .A1(n1221), .B0(n313), .B1(n337), .Y(n1665) );
  OAI22X1 U101 ( .A0(n1735), .A1(n1217), .B0(n313), .B1(n336), .Y(n1666) );
  OAI22X1 U102 ( .A0(n1735), .A1(n1213), .B0(n313), .B1(n335), .Y(n1667) );
  OAI22X1 U103 ( .A0(n1735), .A1(n1209), .B0(n314), .B1(n334), .Y(n1668) );
  OAI22X1 U104 ( .A0(n1735), .A1(n1205), .B0(n314), .B1(n333), .Y(n1669) );
  OAI22X1 U105 ( .A0(n316), .A1(n1201), .B0(n314), .B1(n332), .Y(n1670) );
  OAI22X1 U106 ( .A0(n309), .A1(n728), .B0(n347), .B1(n306), .Y(n1527) );
  OAI22X1 U107 ( .A0(n1733), .A1(n720), .B0(n346), .B1(n1732), .Y(n1528) );
  OAI22X1 U108 ( .A0(n1733), .A1(n712), .B0(n345), .B1(n1732), .Y(n1529) );
  OAI22X1 U109 ( .A0(n1733), .A1(n704), .B0(n344), .B1(n1732), .Y(n1530) );
  OAI22X1 U110 ( .A0(n1733), .A1(n696), .B0(n343), .B1(n1732), .Y(n1531) );
  OAI22X1 U111 ( .A0(n1733), .A1(n688), .B0(n342), .B1(n303), .Y(n1532) );
  OAI22X1 U112 ( .A0(n1733), .A1(n680), .B0(n341), .B1(n306), .Y(n1533) );
  OAI22X1 U113 ( .A0(n1733), .A1(n672), .B0(n340), .B1(n304), .Y(n1534) );
  OAI22X1 U114 ( .A0(n1733), .A1(n664), .B0(n339), .B1(n304), .Y(n1535) );
  OAI22X1 U115 ( .A0(n1733), .A1(n656), .B0(n338), .B1(n305), .Y(n1536) );
  OAI22X1 U116 ( .A0(n1733), .A1(n648), .B0(n337), .B1(n303), .Y(n1537) );
  OAI22X1 U117 ( .A0(n289), .A1(n592), .B0(n347), .B1(n286), .Y(n1271) );
  OAI22X1 U118 ( .A0(n289), .A1(n576), .B0(n346), .B1(n282), .Y(n1272) );
  OAI22X1 U119 ( .A0(n289), .A1(n560), .B0(n345), .B1(n285), .Y(n1273) );
  OAI22X1 U120 ( .A0(n295), .A1(n544), .B0(n344), .B1(n285), .Y(n1274) );
  OAI22X1 U121 ( .A0(n302), .A1(n528), .B0(n343), .B1(n282), .Y(n1275) );
  OAI22X1 U122 ( .A0(n293), .A1(n512), .B0(n342), .B1(n285), .Y(n1276) );
  OAI22X1 U123 ( .A0(n295), .A1(n496), .B0(n341), .B1(n282), .Y(n1277) );
  OAI22X1 U124 ( .A0(n295), .A1(n480), .B0(n340), .B1(n278), .Y(n1278) );
  OAI22X1 U125 ( .A0(n295), .A1(n464), .B0(n339), .B1(n285), .Y(n1279) );
  INVX1 U126 ( .A(din[1]), .Y(n346) );
  INVX1 U127 ( .A(din[2]), .Y(n345) );
  INVX1 U128 ( .A(din[3]), .Y(n344) );
  INVX1 U129 ( .A(din[4]), .Y(n343) );
  INVX1 U130 ( .A(din[5]), .Y(n342) );
  INVX1 U131 ( .A(din[6]), .Y(n341) );
  INVX1 U132 ( .A(din[7]), .Y(n340) );
  INVX1 U133 ( .A(din[8]), .Y(n339) );
  INVX1 U134 ( .A(din[9]), .Y(n338) );
  INVX1 U135 ( .A(din[10]), .Y(n337) );
  INVX1 U136 ( .A(din[11]), .Y(n336) );
  INVX1 U137 ( .A(din[12]), .Y(n335) );
  INVX1 U138 ( .A(din[0]), .Y(n347) );
  INVX1 U139 ( .A(din[13]), .Y(n334) );
  INVX1 U140 ( .A(din[14]), .Y(n333) );
  INVX1 U141 ( .A(din[15]), .Y(n332) );
  OAI211X1 U142 ( .A0(n1267), .A1(n1270), .B0(n1269), .C0(start), .Y(n1735) );
  NAND2X1 U143 ( .A(start), .B(n1720), .Y(n1721) );
  OAI222XL U144 ( .A0(n1722), .A1(n1266), .B0(n1723), .B1(n1268), .C0(n1724), 
        .C1(n1269), .Y(n1720) );
  OAI22X1 U145 ( .A0(n308), .A1(n738), .B0(n304), .B1(n732), .Y(n1591) );
  OAI22X1 U146 ( .A0(n309), .A1(n732), .B0(n305), .B1(n730), .Y(n1575) );
  OAI22X1 U147 ( .A0(n310), .A1(n730), .B0(n306), .B1(n729), .Y(n1559) );
  OAI22X1 U148 ( .A0(n1733), .A1(n729), .B0(n1732), .B1(n728), .Y(n1543) );
  OAI22X1 U149 ( .A0(n310), .A1(n724), .B0(n304), .B1(n723), .Y(n1592) );
  OAI22X1 U150 ( .A0(n309), .A1(n723), .B0(n305), .B1(n722), .Y(n1576) );
  OAI22X1 U151 ( .A0(n310), .A1(n722), .B0(n306), .B1(n721), .Y(n1560) );
  OAI22X1 U152 ( .A0(n1733), .A1(n721), .B0(n1732), .B1(n720), .Y(n1544) );
  OAI22X1 U153 ( .A0(n311), .A1(n716), .B0(n304), .B1(n715), .Y(n1593) );
  OAI22X1 U154 ( .A0(n309), .A1(n715), .B0(n303), .B1(n714), .Y(n1577) );
  OAI22X1 U155 ( .A0(n310), .A1(n714), .B0(n306), .B1(n713), .Y(n1561) );
  OAI22X1 U156 ( .A0(n1733), .A1(n713), .B0(n1732), .B1(n712), .Y(n1545) );
  OAI22X1 U157 ( .A0(n308), .A1(n708), .B0(n304), .B1(n707), .Y(n1594) );
  OAI22X1 U158 ( .A0(n309), .A1(n707), .B0(n306), .B1(n706), .Y(n1578) );
  OAI22X1 U159 ( .A0(n310), .A1(n706), .B0(n306), .B1(n705), .Y(n1562) );
  OAI22X1 U160 ( .A0(n1733), .A1(n705), .B0(n1732), .B1(n704), .Y(n1546) );
  OAI22X1 U161 ( .A0(n308), .A1(n700), .B0(n304), .B1(n699), .Y(n1595) );
  OAI22X1 U162 ( .A0(n309), .A1(n699), .B0(n305), .B1(n698), .Y(n1579) );
  OAI22X1 U163 ( .A0(n310), .A1(n698), .B0(n306), .B1(n697), .Y(n1563) );
  OAI22X1 U164 ( .A0(n311), .A1(n697), .B0(n1732), .B1(n696), .Y(n1547) );
  OAI22X1 U165 ( .A0(n308), .A1(n692), .B0(n304), .B1(n691), .Y(n1596) );
  OAI22X1 U166 ( .A0(n309), .A1(n691), .B0(n304), .B1(n690), .Y(n1580) );
  OAI22X1 U167 ( .A0(n310), .A1(n690), .B0(n305), .B1(n689), .Y(n1564) );
  OAI22X1 U168 ( .A0(n311), .A1(n689), .B0(n1732), .B1(n688), .Y(n1548) );
  OAI22X1 U169 ( .A0(n308), .A1(n684), .B0(n304), .B1(n683), .Y(n1597) );
  OAI22X1 U170 ( .A0(n309), .A1(n683), .B0(n303), .B1(n682), .Y(n1581) );
  OAI22X1 U171 ( .A0(n310), .A1(n682), .B0(n305), .B1(n681), .Y(n1565) );
  OAI22X1 U172 ( .A0(n311), .A1(n681), .B0(n1732), .B1(n680), .Y(n1549) );
  OAI22X1 U173 ( .A0(n308), .A1(n676), .B0(n304), .B1(n675), .Y(n1598) );
  OAI22X1 U174 ( .A0(n309), .A1(n675), .B0(n306), .B1(n674), .Y(n1582) );
  OAI22X1 U175 ( .A0(n310), .A1(n674), .B0(n305), .B1(n673), .Y(n1566) );
  OAI22X1 U176 ( .A0(n311), .A1(n673), .B0(n1732), .B1(n672), .Y(n1550) );
  OAI22X1 U177 ( .A0(n308), .A1(n668), .B0(n304), .B1(n667), .Y(n1599) );
  OAI22X1 U178 ( .A0(n310), .A1(n667), .B0(n305), .B1(n666), .Y(n1583) );
  OAI22X1 U179 ( .A0(n310), .A1(n666), .B0(n305), .B1(n665), .Y(n1567) );
  OAI22X1 U180 ( .A0(n311), .A1(n665), .B0(n306), .B1(n664), .Y(n1551) );
  OAI22X1 U181 ( .A0(n308), .A1(n660), .B0(n304), .B1(n659), .Y(n1600) );
  OAI22X1 U182 ( .A0(n309), .A1(n659), .B0(n304), .B1(n658), .Y(n1584) );
  OAI22X1 U183 ( .A0(n310), .A1(n658), .B0(n305), .B1(n657), .Y(n1568) );
  OAI22X1 U184 ( .A0(n311), .A1(n657), .B0(n306), .B1(n656), .Y(n1552) );
  OAI22X1 U185 ( .A0(n308), .A1(n652), .B0(n304), .B1(n651), .Y(n1601) );
  OAI22X1 U186 ( .A0(n1733), .A1(n651), .B0(n305), .B1(n650), .Y(n1585) );
  OAI22X1 U187 ( .A0(n310), .A1(n650), .B0(n305), .B1(n649), .Y(n1569) );
  OAI22X1 U188 ( .A0(n311), .A1(n649), .B0(n306), .B1(n648), .Y(n1553) );
  OAI22X1 U189 ( .A0(n308), .A1(n644), .B0(n304), .B1(n643), .Y(n1602) );
  OAI22X1 U190 ( .A0(n1733), .A1(n643), .B0(n304), .B1(n642), .Y(n1586) );
  OAI22X1 U191 ( .A0(n310), .A1(n642), .B0(n305), .B1(n641), .Y(n1570) );
  OAI22X1 U192 ( .A0(n311), .A1(n641), .B0(n306), .B1(n640), .Y(n1554) );
  OAI22X1 U193 ( .A0(n308), .A1(n636), .B0(n306), .B1(n635), .Y(n1603) );
  OAI22X1 U194 ( .A0(n1733), .A1(n635), .B0(n303), .B1(n634), .Y(n1587) );
  OAI22X1 U195 ( .A0(n309), .A1(n634), .B0(n305), .B1(n633), .Y(n1571) );
  OAI22X1 U196 ( .A0(n311), .A1(n633), .B0(n306), .B1(n632), .Y(n1555) );
  OAI22X1 U197 ( .A0(n308), .A1(n628), .B0(n303), .B1(n627), .Y(n1604) );
  OAI22X1 U198 ( .A0(n1733), .A1(n627), .B0(n306), .B1(n626), .Y(n1588) );
  OAI22X1 U199 ( .A0(n309), .A1(n626), .B0(n305), .B1(n625), .Y(n1572) );
  OAI22X1 U200 ( .A0(n311), .A1(n625), .B0(n306), .B1(n624), .Y(n1556) );
  OAI22X1 U201 ( .A0(n308), .A1(n620), .B0(n306), .B1(n619), .Y(n1605) );
  OAI22X1 U202 ( .A0(n1733), .A1(n619), .B0(n305), .B1(n618), .Y(n1589) );
  OAI22X1 U203 ( .A0(n309), .A1(n618), .B0(n305), .B1(n617), .Y(n1573) );
  OAI22X1 U204 ( .A0(n311), .A1(n617), .B0(n306), .B1(n616), .Y(n1557) );
  OAI22X1 U205 ( .A0(n310), .A1(n612), .B0(n304), .B1(n611), .Y(n1606) );
  OAI22X1 U206 ( .A0(n1733), .A1(n611), .B0(n304), .B1(n610), .Y(n1590) );
  OAI22X1 U207 ( .A0(n309), .A1(n610), .B0(n305), .B1(n609), .Y(n1574) );
  OAI22X1 U208 ( .A0(n311), .A1(n609), .B0(n306), .B1(n608), .Y(n1558) );
  OAI22X1 U209 ( .A0(n294), .A1(n604), .B0(n279), .B1(n603), .Y(n1463) );
  OAI22X1 U210 ( .A0(n293), .A1(n603), .B0(n281), .B1(n602), .Y(n1447) );
  OAI22X1 U211 ( .A0(n291), .A1(n602), .B0(n287), .B1(n601), .Y(n1431) );
  OAI22X1 U212 ( .A0(n290), .A1(n601), .B0(n282), .B1(n600), .Y(n1415) );
  OAI22X1 U213 ( .A0(n294), .A1(n600), .B0(n283), .B1(n599), .Y(n1399) );
  OAI22X1 U214 ( .A0(n302), .A1(n599), .B0(n285), .B1(n598), .Y(n1383) );
  OAI22X1 U215 ( .A0(n300), .A1(n598), .B0(n286), .B1(n597), .Y(n1367) );
  OAI22X1 U216 ( .A0(n299), .A1(n597), .B0(n287), .B1(n596), .Y(n1351) );
  OAI22X1 U217 ( .A0(n290), .A1(n596), .B0(n283), .B1(n595), .Y(n1335) );
  OAI22X1 U218 ( .A0(n298), .A1(n595), .B0(n283), .B1(n594), .Y(n1319) );
  OAI22X1 U219 ( .A0(n297), .A1(n594), .B0(n281), .B1(n593), .Y(n1303) );
  OAI22X1 U220 ( .A0(n295), .A1(n593), .B0(n283), .B1(n592), .Y(n1287) );
  OAI22X1 U221 ( .A0(n294), .A1(n588), .B0(n288), .B1(n587), .Y(n1464) );
  OAI22X1 U222 ( .A0(n293), .A1(n587), .B0(n281), .B1(n586), .Y(n1448) );
  OAI22X1 U223 ( .A0(n291), .A1(n586), .B0(n280), .B1(n585), .Y(n1432) );
  OAI22X1 U224 ( .A0(n290), .A1(n585), .B0(n282), .B1(n584), .Y(n1416) );
  OAI22X1 U225 ( .A0(n289), .A1(n584), .B0(n283), .B1(n583), .Y(n1400) );
  OAI22X1 U226 ( .A0(n301), .A1(n583), .B0(n284), .B1(n582), .Y(n1384) );
  OAI22X1 U227 ( .A0(n300), .A1(n582), .B0(n286), .B1(n581), .Y(n1368) );
  OAI22X1 U228 ( .A0(n299), .A1(n581), .B0(n287), .B1(n580), .Y(n1352) );
  OAI22X1 U229 ( .A0(n300), .A1(n580), .B0(n278), .B1(n579), .Y(n1336) );
  OAI22X1 U230 ( .A0(n298), .A1(n579), .B0(n279), .B1(n578), .Y(n1320) );
  OAI22X1 U231 ( .A0(n297), .A1(n578), .B0(n287), .B1(n577), .Y(n1304) );
  OAI22X1 U232 ( .A0(n295), .A1(n577), .B0(n279), .B1(n576), .Y(n1288) );
  OAI22X1 U233 ( .A0(n294), .A1(n572), .B0(n278), .B1(n571), .Y(n1465) );
  OAI22X1 U234 ( .A0(n293), .A1(n571), .B0(n280), .B1(n570), .Y(n1449) );
  OAI22X1 U235 ( .A0(n291), .A1(n570), .B0(n285), .B1(n569), .Y(n1433) );
  OAI22X1 U236 ( .A0(n290), .A1(n569), .B0(n282), .B1(n568), .Y(n1417) );
  OAI22X1 U237 ( .A0(n289), .A1(n568), .B0(n283), .B1(n567), .Y(n1401) );
  OAI22X1 U238 ( .A0(n302), .A1(n567), .B0(n284), .B1(n566), .Y(n1385) );
  OAI22X1 U239 ( .A0(n300), .A1(n566), .B0(n286), .B1(n565), .Y(n1369) );
  OAI22X1 U240 ( .A0(n299), .A1(n565), .B0(n287), .B1(n564), .Y(n1353) );
  OAI22X1 U241 ( .A0(n301), .A1(n564), .B0(n280), .B1(n563), .Y(n1337) );
  OAI22X1 U242 ( .A0(n298), .A1(n563), .B0(n288), .B1(n562), .Y(n1321) );
  OAI22X1 U243 ( .A0(n297), .A1(n562), .B0(n284), .B1(n561), .Y(n1305) );
  OAI22X1 U244 ( .A0(n296), .A1(n561), .B0(n281), .B1(n560), .Y(n1289) );
  OAI22X1 U245 ( .A0(n294), .A1(n556), .B0(n280), .B1(n555), .Y(n1466) );
  OAI22X1 U246 ( .A0(n293), .A1(n555), .B0(n280), .B1(n554), .Y(n1450) );
  OAI22X1 U247 ( .A0(n291), .A1(n554), .B0(n283), .B1(n553), .Y(n1434) );
  OAI22X1 U248 ( .A0(n290), .A1(n553), .B0(n282), .B1(n552), .Y(n1418) );
  OAI22X1 U249 ( .A0(n289), .A1(n552), .B0(n283), .B1(n551), .Y(n1402) );
  OAI22X1 U250 ( .A0(n302), .A1(n551), .B0(n284), .B1(n550), .Y(n1386) );
  OAI22X1 U251 ( .A0(n300), .A1(n550), .B0(n286), .B1(n549), .Y(n1370) );
  OAI22X1 U252 ( .A0(n299), .A1(n549), .B0(n287), .B1(n548), .Y(n1354) );
  OAI22X1 U253 ( .A0(n292), .A1(n548), .B0(n281), .B1(n547), .Y(n1338) );
  OAI22X1 U254 ( .A0(n298), .A1(n547), .B0(n278), .B1(n546), .Y(n1322) );
  OAI22X1 U255 ( .A0(n297), .A1(n546), .B0(n288), .B1(n545), .Y(n1306) );
  OAI22X1 U256 ( .A0(n296), .A1(n545), .B0(n287), .B1(n544), .Y(n1290) );
  OAI22X1 U257 ( .A0(n294), .A1(n540), .B0(n281), .B1(n539), .Y(n1467) );
  OAI22X1 U258 ( .A0(n293), .A1(n539), .B0(n280), .B1(n538), .Y(n1451) );
  OAI22X1 U259 ( .A0(n292), .A1(n538), .B0(n280), .B1(n537), .Y(n1435) );
  OAI22X1 U260 ( .A0(n290), .A1(n537), .B0(n282), .B1(n536), .Y(n1419) );
  OAI22X1 U261 ( .A0(n289), .A1(n536), .B0(n283), .B1(n535), .Y(n1403) );
  OAI22X1 U262 ( .A0(n302), .A1(n535), .B0(n284), .B1(n534), .Y(n1387) );
  OAI22X1 U263 ( .A0(n300), .A1(n534), .B0(n285), .B1(n533), .Y(n1371) );
  OAI22X1 U264 ( .A0(n299), .A1(n533), .B0(n287), .B1(n532), .Y(n1355) );
  OAI22X1 U265 ( .A0(n290), .A1(n532), .B0(n280), .B1(n531), .Y(n1339) );
  OAI22X1 U266 ( .A0(n298), .A1(n531), .B0(n280), .B1(n530), .Y(n1323) );
  OAI22X1 U267 ( .A0(n297), .A1(n530), .B0(n288), .B1(n529), .Y(n1307) );
  OAI22X1 U268 ( .A0(n296), .A1(n529), .B0(n287), .B1(n528), .Y(n1291) );
  OAI22X1 U269 ( .A0(n294), .A1(n524), .B0(n283), .B1(n523), .Y(n1468) );
  OAI22X1 U270 ( .A0(n293), .A1(n523), .B0(n280), .B1(n522), .Y(n1452) );
  OAI22X1 U271 ( .A0(n292), .A1(n522), .B0(n281), .B1(n521), .Y(n1436) );
  OAI22X1 U272 ( .A0(n290), .A1(n521), .B0(n282), .B1(n520), .Y(n1420) );
  OAI22X1 U273 ( .A0(n289), .A1(n520), .B0(n283), .B1(n519), .Y(n1404) );
  OAI22X1 U274 ( .A0(n302), .A1(n519), .B0(n284), .B1(n518), .Y(n1388) );
  OAI22X1 U275 ( .A0(n301), .A1(n518), .B0(n285), .B1(n517), .Y(n1372) );
  OAI22X1 U276 ( .A0(n299), .A1(n517), .B0(n287), .B1(n516), .Y(n1356) );
  OAI22X1 U277 ( .A0(n294), .A1(n516), .B0(n287), .B1(n515), .Y(n1340) );
  OAI22X1 U278 ( .A0(n298), .A1(n515), .B0(n281), .B1(n514), .Y(n1324) );
  OAI22X1 U279 ( .A0(n297), .A1(n514), .B0(n288), .B1(n513), .Y(n1308) );
  OAI22X1 U280 ( .A0(n296), .A1(n513), .B0(n283), .B1(n512), .Y(n1292) );
  OAI22X1 U281 ( .A0(n294), .A1(n508), .B0(n287), .B1(n507), .Y(n1469) );
  OAI22X1 U282 ( .A0(n293), .A1(n507), .B0(n280), .B1(n506), .Y(n1453) );
  OAI22X1 U283 ( .A0(n292), .A1(n506), .B0(n281), .B1(n505), .Y(n1437) );
  OAI22X1 U284 ( .A0(n290), .A1(n505), .B0(n282), .B1(n504), .Y(n1421) );
  OAI22X1 U285 ( .A0(n289), .A1(n504), .B0(n283), .B1(n503), .Y(n1405) );
  OAI22X1 U286 ( .A0(n302), .A1(n503), .B0(n284), .B1(n502), .Y(n1389) );
  OAI22X1 U287 ( .A0(n301), .A1(n502), .B0(n285), .B1(n501), .Y(n1373) );
  OAI22X1 U288 ( .A0(n299), .A1(n501), .B0(n287), .B1(n500), .Y(n1357) );
  OAI22X1 U289 ( .A0(n295), .A1(n500), .B0(n281), .B1(n499), .Y(n1341) );
  OAI22X1 U290 ( .A0(n301), .A1(n499), .B0(n285), .B1(n498), .Y(n1325) );
  OAI22X1 U291 ( .A0(n297), .A1(n498), .B0(n288), .B1(n497), .Y(n1309) );
  OAI22X1 U292 ( .A0(n296), .A1(n497), .B0(n283), .B1(n496), .Y(n1293) );
  OAI22X1 U293 ( .A0(n297), .A1(n492), .B0(n286), .B1(n491), .Y(n1470) );
  OAI22X1 U294 ( .A0(n293), .A1(n491), .B0(n280), .B1(n490), .Y(n1454) );
  OAI22X1 U295 ( .A0(n292), .A1(n490), .B0(n281), .B1(n489), .Y(n1438) );
  OAI22X1 U296 ( .A0(n290), .A1(n489), .B0(n282), .B1(n488), .Y(n1422) );
  OAI22X1 U297 ( .A0(n289), .A1(n488), .B0(n283), .B1(n487), .Y(n1406) );
  OAI22X1 U298 ( .A0(n302), .A1(n487), .B0(n284), .B1(n486), .Y(n1390) );
  OAI22X1 U299 ( .A0(n301), .A1(n486), .B0(n285), .B1(n485), .Y(n1374) );
  OAI22X1 U300 ( .A0(n299), .A1(n485), .B0(n286), .B1(n484), .Y(n1358) );
  OAI22X1 U301 ( .A0(n302), .A1(n484), .B0(n285), .B1(n483), .Y(n1342) );
  OAI22X1 U302 ( .A0(n292), .A1(n483), .B0(n282), .B1(n482), .Y(n1326) );
  OAI22X1 U303 ( .A0(n297), .A1(n482), .B0(n288), .B1(n481), .Y(n1310) );
  OAI22X1 U304 ( .A0(n296), .A1(n481), .B0(n279), .B1(n480), .Y(n1294) );
  OAI22X1 U305 ( .A0(n289), .A1(n476), .B0(n284), .B1(n475), .Y(n1471) );
  OAI22X1 U306 ( .A0(n293), .A1(n475), .B0(n280), .B1(n474), .Y(n1455) );
  OAI22X1 U307 ( .A0(n292), .A1(n474), .B0(n281), .B1(n473), .Y(n1439) );
  OAI22X1 U308 ( .A0(n291), .A1(n473), .B0(n281), .B1(n472), .Y(n1423) );
  OAI22X1 U309 ( .A0(n289), .A1(n472), .B0(n283), .B1(n471), .Y(n1407) );
  OAI22X1 U310 ( .A0(n302), .A1(n471), .B0(n284), .B1(n470), .Y(n1391) );
  OAI22X1 U311 ( .A0(n301), .A1(n470), .B0(n285), .B1(n469), .Y(n1375) );
  OAI22X1 U312 ( .A0(n299), .A1(n469), .B0(n286), .B1(n468), .Y(n1359) );
  OAI22X1 U313 ( .A0(n289), .A1(n468), .B0(n286), .B1(n467), .Y(n1343) );
  OAI22X1 U314 ( .A0(n294), .A1(n467), .B0(n286), .B1(n466), .Y(n1327) );
  OAI22X1 U315 ( .A0(n297), .A1(n466), .B0(n288), .B1(n465), .Y(n1311) );
  OAI22X1 U316 ( .A0(n296), .A1(n465), .B0(n282), .B1(n464), .Y(n1295) );
  OAI22X1 U317 ( .A0(n295), .A1(n460), .B0(n279), .B1(n459), .Y(n1472) );
  OAI22X1 U318 ( .A0(n293), .A1(n459), .B0(n280), .B1(n458), .Y(n1456) );
  OAI22X1 U319 ( .A0(n292), .A1(n458), .B0(n281), .B1(n457), .Y(n1440) );
  OAI22X1 U320 ( .A0(n291), .A1(n457), .B0(n287), .B1(n456), .Y(n1424) );
  OAI22X1 U321 ( .A0(n289), .A1(n456), .B0(n283), .B1(n455), .Y(n1408) );
  OAI22X1 U322 ( .A0(n302), .A1(n455), .B0(n284), .B1(n454), .Y(n1392) );
  OAI22X1 U323 ( .A0(n301), .A1(n454), .B0(n285), .B1(n453), .Y(n1376) );
  OAI22X1 U324 ( .A0(n300), .A1(n453), .B0(n286), .B1(n452), .Y(n1360) );
  OAI22X1 U325 ( .A0(n296), .A1(n452), .B0(n283), .B1(n451), .Y(n1344) );
  OAI22X1 U326 ( .A0(n296), .A1(n451), .B0(n287), .B1(n450), .Y(n1328) );
  OAI22X1 U327 ( .A0(n297), .A1(n450), .B0(n288), .B1(n449), .Y(n1312) );
  OAI22X1 U328 ( .A0(n296), .A1(n449), .B0(n285), .B1(n448), .Y(n1296) );
  OAI22X1 U329 ( .A0(n293), .A1(n444), .B0(n288), .B1(n443), .Y(n1473) );
  OAI22X1 U330 ( .A0(n293), .A1(n443), .B0(n280), .B1(n442), .Y(n1457) );
  OAI22X1 U331 ( .A0(n292), .A1(n442), .B0(n281), .B1(n441), .Y(n1441) );
  OAI22X1 U332 ( .A0(n291), .A1(n441), .B0(n286), .B1(n440), .Y(n1425) );
  OAI22X1 U333 ( .A0(n289), .A1(n440), .B0(n283), .B1(n439), .Y(n1409) );
  OAI22X1 U334 ( .A0(n302), .A1(n439), .B0(n284), .B1(n438), .Y(n1393) );
  OAI22X1 U335 ( .A0(n301), .A1(n438), .B0(n285), .B1(n437), .Y(n1377) );
  OAI22X1 U336 ( .A0(n300), .A1(n437), .B0(n286), .B1(n436), .Y(n1361) );
  OAI22X1 U337 ( .A0(n298), .A1(n436), .B0(n287), .B1(n435), .Y(n1345) );
  OAI22X1 U338 ( .A0(n295), .A1(n435), .B0(n284), .B1(n434), .Y(n1329) );
  OAI22X1 U339 ( .A0(n298), .A1(n434), .B0(n288), .B1(n433), .Y(n1313) );
  OAI22X1 U340 ( .A0(n296), .A1(n433), .B0(n286), .B1(n432), .Y(n1297) );
  OAI22X1 U341 ( .A0(n291), .A1(n428), .B0(n284), .B1(n427), .Y(n1474) );
  OAI22X1 U342 ( .A0(n293), .A1(n427), .B0(n280), .B1(n426), .Y(n1458) );
  OAI22X1 U343 ( .A0(n292), .A1(n426), .B0(n281), .B1(n425), .Y(n1442) );
  OAI22X1 U344 ( .A0(n291), .A1(n425), .B0(n284), .B1(n424), .Y(n1426) );
  OAI22X1 U345 ( .A0(n289), .A1(n424), .B0(n282), .B1(n423), .Y(n1410) );
  OAI22X1 U346 ( .A0(n302), .A1(n423), .B0(n284), .B1(n422), .Y(n1394) );
  OAI22X1 U347 ( .A0(n301), .A1(n422), .B0(n285), .B1(n421), .Y(n1378) );
  OAI22X1 U348 ( .A0(n300), .A1(n421), .B0(n286), .B1(n420), .Y(n1362) );
  OAI22X1 U349 ( .A0(n297), .A1(n420), .B0(n287), .B1(n419), .Y(n1346) );
  OAI22X1 U350 ( .A0(n289), .A1(n419), .B0(n283), .B1(n418), .Y(n1330) );
  OAI22X1 U351 ( .A0(n298), .A1(n418), .B0(n288), .B1(n417), .Y(n1314) );
  OAI22X1 U352 ( .A0(n296), .A1(n417), .B0(n280), .B1(n416), .Y(n1298) );
  OAI22X1 U353 ( .A0(n291), .A1(n412), .B0(n279), .B1(n411), .Y(n1475) );
  OAI22X1 U354 ( .A0(n294), .A1(n411), .B0(n280), .B1(n410), .Y(n1459) );
  OAI22X1 U355 ( .A0(n292), .A1(n410), .B0(n281), .B1(n409), .Y(n1443) );
  OAI22X1 U356 ( .A0(n291), .A1(n409), .B0(n279), .B1(n408), .Y(n1427) );
  OAI22X1 U357 ( .A0(n290), .A1(n408), .B0(n282), .B1(n407), .Y(n1411) );
  OAI22X1 U358 ( .A0(n300), .A1(n407), .B0(n284), .B1(n406), .Y(n1395) );
  OAI22X1 U359 ( .A0(n301), .A1(n406), .B0(n285), .B1(n405), .Y(n1379) );
  OAI22X1 U360 ( .A0(n300), .A1(n405), .B0(n286), .B1(n404), .Y(n1363) );
  OAI22X1 U361 ( .A0(n293), .A1(n404), .B0(n287), .B1(n403), .Y(n1347) );
  OAI22X1 U362 ( .A0(n301), .A1(n403), .B0(n279), .B1(n402), .Y(n1331) );
  OAI22X1 U363 ( .A0(n298), .A1(n402), .B0(n288), .B1(n401), .Y(n1315) );
  OAI22X1 U364 ( .A0(n296), .A1(n401), .B0(n281), .B1(n400), .Y(n1299) );
  OAI22X1 U365 ( .A0(n299), .A1(n396), .B0(n279), .B1(n395), .Y(n1476) );
  OAI22X1 U366 ( .A0(n294), .A1(n395), .B0(n280), .B1(n394), .Y(n1460) );
  OAI22X1 U367 ( .A0(n292), .A1(n394), .B0(n281), .B1(n393), .Y(n1444) );
  OAI22X1 U368 ( .A0(n291), .A1(n393), .B0(n288), .B1(n392), .Y(n1428) );
  OAI22X1 U369 ( .A0(n290), .A1(n392), .B0(n282), .B1(n391), .Y(n1412) );
  OAI22X1 U370 ( .A0(n302), .A1(n391), .B0(n284), .B1(n390), .Y(n1396) );
  OAI22X1 U371 ( .A0(n301), .A1(n390), .B0(n285), .B1(n389), .Y(n1380) );
  OAI22X1 U372 ( .A0(n300), .A1(n389), .B0(n286), .B1(n388), .Y(n1364) );
  OAI22X1 U373 ( .A0(n299), .A1(n388), .B0(n287), .B1(n387), .Y(n1348) );
  OAI22X1 U374 ( .A0(n292), .A1(n387), .B0(n284), .B1(n386), .Y(n1332) );
  OAI22X1 U375 ( .A0(n298), .A1(n386), .B0(n288), .B1(n385), .Y(n1316) );
  OAI22X1 U376 ( .A0(n296), .A1(n385), .B0(n287), .B1(n384), .Y(n1300) );
  OAI22X1 U377 ( .A0(n302), .A1(n380), .B0(n279), .B1(n379), .Y(n1477) );
  OAI22X1 U378 ( .A0(n294), .A1(n379), .B0(n280), .B1(n378), .Y(n1461) );
  OAI22X1 U379 ( .A0(n292), .A1(n378), .B0(n281), .B1(n377), .Y(n1445) );
  OAI22X1 U380 ( .A0(n291), .A1(n377), .B0(n278), .B1(n376), .Y(n1429) );
  OAI22X1 U381 ( .A0(n290), .A1(n376), .B0(n282), .B1(n375), .Y(n1413) );
  OAI22X1 U382 ( .A0(n301), .A1(n375), .B0(n283), .B1(n374), .Y(n1397) );
  OAI22X1 U383 ( .A0(n301), .A1(n374), .B0(n285), .B1(n373), .Y(n1381) );
  OAI22X1 U384 ( .A0(n300), .A1(n373), .B0(n286), .B1(n372), .Y(n1365) );
  OAI22X1 U385 ( .A0(n299), .A1(n372), .B0(n287), .B1(n371), .Y(n1349) );
  OAI22X1 U386 ( .A0(n294), .A1(n371), .B0(n279), .B1(n370), .Y(n1333) );
  OAI22X1 U387 ( .A0(n298), .A1(n370), .B0(n288), .B1(n369), .Y(n1317) );
  OAI22X1 U388 ( .A0(n297), .A1(n369), .B0(n284), .B1(n368), .Y(n1301) );
  OAI22X1 U389 ( .A0(n301), .A1(n364), .B0(n279), .B1(n363), .Y(n1478) );
  OAI22X1 U390 ( .A0(n294), .A1(n363), .B0(n278), .B1(n362), .Y(n1462) );
  OAI22X1 U391 ( .A0(n292), .A1(n362), .B0(n281), .B1(n361), .Y(n1446) );
  OAI22X1 U392 ( .A0(n291), .A1(n361), .B0(n282), .B1(n360), .Y(n1430) );
  OAI22X1 U393 ( .A0(n290), .A1(n360), .B0(n282), .B1(n359), .Y(n1414) );
  OAI22X1 U394 ( .A0(n292), .A1(n359), .B0(n283), .B1(n358), .Y(n1398) );
  OAI22X1 U395 ( .A0(n301), .A1(n358), .B0(n285), .B1(n357), .Y(n1382) );
  OAI22X1 U396 ( .A0(n300), .A1(n357), .B0(n286), .B1(n356), .Y(n1366) );
  OAI22X1 U397 ( .A0(n299), .A1(n356), .B0(n287), .B1(n355), .Y(n1350) );
  OAI22X1 U398 ( .A0(n296), .A1(n355), .B0(n288), .B1(n354), .Y(n1334) );
  OAI22X1 U399 ( .A0(n298), .A1(n354), .B0(n288), .B1(n353), .Y(n1318) );
  OAI22X1 U400 ( .A0(n297), .A1(n353), .B0(n283), .B1(n352), .Y(n1302) );
  OAI22X1 U401 ( .A0(n1735), .A1(n1264), .B0(n313), .B1(n1263), .Y(n1703) );
  OAI22X1 U402 ( .A0(n1735), .A1(n1263), .B0(n313), .B1(n1262), .Y(n1687) );
  OAI22X1 U403 ( .A0(n1735), .A1(n1262), .B0(n314), .B1(n1261), .Y(n1671) );
  OAI22X1 U404 ( .A0(n1735), .A1(n1260), .B0(n314), .B1(n1259), .Y(n1704) );
  OAI22X1 U405 ( .A0(n1735), .A1(n1259), .B0(n314), .B1(n1258), .Y(n1688) );
  OAI22X1 U406 ( .A0(n316), .A1(n1258), .B0(n314), .B1(n1257), .Y(n1672) );
  OAI22X1 U407 ( .A0(n1735), .A1(n1256), .B0(n313), .B1(n1255), .Y(n1705) );
  OAI22X1 U408 ( .A0(n1735), .A1(n1255), .B0(n314), .B1(n1254), .Y(n1689) );
  OAI22X1 U409 ( .A0(n316), .A1(n1254), .B0(n314), .B1(n1253), .Y(n1673) );
  OAI22X1 U410 ( .A0(n1735), .A1(n1252), .B0(n314), .B1(n1251), .Y(n1706) );
  OAI22X1 U411 ( .A0(n1735), .A1(n1251), .B0(n313), .B1(n1250), .Y(n1690) );
  OAI22X1 U412 ( .A0(n316), .A1(n1250), .B0(n314), .B1(n1249), .Y(n1674) );
  OAI22X1 U413 ( .A0(n315), .A1(n1248), .B0(n313), .B1(n1247), .Y(n1707) );
  OAI22X1 U414 ( .A0(n1735), .A1(n1247), .B0(n314), .B1(n1246), .Y(n1691) );
  OAI22X1 U415 ( .A0(n316), .A1(n1246), .B0(n314), .B1(n1245), .Y(n1675) );
  OAI22X1 U416 ( .A0(n315), .A1(n1244), .B0(n314), .B1(n1243), .Y(n1708) );
  OAI22X1 U417 ( .A0(n1735), .A1(n1243), .B0(n313), .B1(n1242), .Y(n1692) );
  OAI22X1 U418 ( .A0(n316), .A1(n1242), .B0(n314), .B1(n1241), .Y(n1676) );
  OAI22X1 U419 ( .A0(n315), .A1(n1240), .B0(n313), .B1(n1239), .Y(n1709) );
  OAI22X1 U420 ( .A0(n1735), .A1(n1239), .B0(n313), .B1(n1238), .Y(n1693) );
  OAI22X1 U421 ( .A0(n316), .A1(n1238), .B0(n314), .B1(n1237), .Y(n1677) );
  OAI22X1 U422 ( .A0(n1735), .A1(n1236), .B0(n314), .B1(n1235), .Y(n1710) );
  OAI22X1 U423 ( .A0(n1735), .A1(n1235), .B0(n313), .B1(n1234), .Y(n1694) );
  OAI22X1 U424 ( .A0(n316), .A1(n1234), .B0(n314), .B1(n1233), .Y(n1678) );
  OAI22X1 U425 ( .A0(n315), .A1(n1232), .B0(n313), .B1(n1231), .Y(n1711) );
  OAI22X1 U426 ( .A0(n1735), .A1(n1231), .B0(n314), .B1(n1230), .Y(n1695) );
  OAI22X1 U427 ( .A0(n316), .A1(n1230), .B0(n314), .B1(n1229), .Y(n1679) );
  OAI22X1 U428 ( .A0(n315), .A1(n1228), .B0(n314), .B1(n1227), .Y(n1712) );
  OAI22X1 U429 ( .A0(n1735), .A1(n1227), .B0(n313), .B1(n1226), .Y(n1696) );
  OAI22X1 U430 ( .A0(n316), .A1(n1226), .B0(n314), .B1(n1225), .Y(n1680) );
  OAI22X1 U431 ( .A0(n315), .A1(n1224), .B0(n314), .B1(n1223), .Y(n1713) );
  OAI22X1 U432 ( .A0(n1735), .A1(n1223), .B0(n314), .B1(n1222), .Y(n1697) );
  OAI22X1 U433 ( .A0(n316), .A1(n1222), .B0(n314), .B1(n1221), .Y(n1681) );
  OAI22X1 U434 ( .A0(n315), .A1(n1220), .B0(n313), .B1(n1219), .Y(n1714) );
  OAI22X1 U435 ( .A0(n1735), .A1(n1219), .B0(n313), .B1(n1218), .Y(n1698) );
  OAI22X1 U436 ( .A0(n316), .A1(n1218), .B0(n314), .B1(n1217), .Y(n1682) );
  OAI22X1 U437 ( .A0(n315), .A1(n1216), .B0(n313), .B1(n1215), .Y(n1715) );
  OAI22X1 U438 ( .A0(n1735), .A1(n1215), .B0(n314), .B1(n1214), .Y(n1699) );
  OAI22X1 U439 ( .A0(n1735), .A1(n1214), .B0(n313), .B1(n1213), .Y(n1683) );
  OAI22X1 U440 ( .A0(n315), .A1(n1212), .B0(n314), .B1(n1211), .Y(n1716) );
  OAI22X1 U441 ( .A0(n1735), .A1(n1211), .B0(n313), .B1(n1210), .Y(n1700) );
  OAI22X1 U442 ( .A0(n1735), .A1(n1210), .B0(n314), .B1(n1209), .Y(n1684) );
  OAI22X1 U443 ( .A0(n315), .A1(n1208), .B0(n313), .B1(n1207), .Y(n1717) );
  OAI22X1 U444 ( .A0(n1735), .A1(n1207), .B0(n314), .B1(n1206), .Y(n1701) );
  OAI22X1 U445 ( .A0(n1735), .A1(n1206), .B0(n313), .B1(n1205), .Y(n1685) );
  OAI22X1 U446 ( .A0(n315), .A1(n1204), .B0(n314), .B1(n1203), .Y(n1718) );
  OAI22X1 U447 ( .A0(n1203), .A1(n1735), .B0(n314), .B1(n1202), .Y(n1702) );
  OAI22X1 U448 ( .A0(n315), .A1(n1202), .B0(n313), .B1(n1201), .Y(n1686) );
  OAI22X1 U449 ( .A0(n308), .A1(n1200), .B0(n303), .B1(n1199), .Y(n1639) );
  OAI22X1 U450 ( .A0(n309), .A1(n1199), .B0(n305), .B1(n739), .Y(n1623) );
  OAI22X1 U451 ( .A0(n308), .A1(n739), .B0(n305), .B1(n738), .Y(n1607) );
  OAI22X1 U452 ( .A0(n311), .A1(n727), .B0(n303), .B1(n726), .Y(n1640) );
  OAI22X1 U453 ( .A0(n308), .A1(n726), .B0(n303), .B1(n725), .Y(n1624) );
  OAI22X1 U454 ( .A0(n309), .A1(n725), .B0(n303), .B1(n724), .Y(n1608) );
  OAI22X1 U455 ( .A0(n309), .A1(n719), .B0(n303), .B1(n718), .Y(n1641) );
  OAI22X1 U456 ( .A0(n308), .A1(n718), .B0(n304), .B1(n717), .Y(n1625) );
  OAI22X1 U457 ( .A0(n311), .A1(n717), .B0(n306), .B1(n716), .Y(n1609) );
  OAI22X1 U458 ( .A0(n308), .A1(n711), .B0(n305), .B1(n710), .Y(n1642) );
  OAI22X1 U459 ( .A0(n310), .A1(n710), .B0(n1732), .B1(n709), .Y(n1626) );
  OAI22X1 U460 ( .A0(n308), .A1(n709), .B0(n303), .B1(n708), .Y(n1610) );
  OAI22X1 U461 ( .A0(n311), .A1(n703), .B0(n303), .B1(n702), .Y(n1643) );
  OAI22X1 U462 ( .A0(n309), .A1(n702), .B0(n1732), .B1(n701), .Y(n1627) );
  OAI22X1 U463 ( .A0(n310), .A1(n701), .B0(n305), .B1(n700), .Y(n1611) );
  OAI22X1 U464 ( .A0(n310), .A1(n695), .B0(n306), .B1(n694), .Y(n1644) );
  OAI22X1 U465 ( .A0(n311), .A1(n694), .B0(n1732), .B1(n693), .Y(n1628) );
  OAI22X1 U466 ( .A0(n309), .A1(n693), .B0(n304), .B1(n692), .Y(n1612) );
  OAI22X1 U467 ( .A0(n309), .A1(n687), .B0(n303), .B1(n686), .Y(n1645) );
  OAI22X1 U468 ( .A0(n311), .A1(n686), .B0(n303), .B1(n685), .Y(n1629) );
  OAI22X1 U469 ( .A0(n309), .A1(n685), .B0(n305), .B1(n684), .Y(n1613) );
  OAI22X1 U470 ( .A0(n308), .A1(n679), .B0(n304), .B1(n678), .Y(n1646) );
  OAI22X1 U471 ( .A0(n308), .A1(n678), .B0(n303), .B1(n677), .Y(n1630) );
  OAI22X1 U472 ( .A0(n311), .A1(n677), .B0(n304), .B1(n676), .Y(n1614) );
  OAI22X1 U473 ( .A0(n308), .A1(n671), .B0(n306), .B1(n670), .Y(n1647) );
  OAI22X1 U474 ( .A0(n310), .A1(n670), .B0(n303), .B1(n669), .Y(n1631) );
  OAI22X1 U475 ( .A0(n309), .A1(n669), .B0(n1732), .B1(n668), .Y(n1615) );
  OAI22X1 U476 ( .A0(n311), .A1(n663), .B0(n304), .B1(n662), .Y(n1648) );
  OAI22X1 U477 ( .A0(n309), .A1(n662), .B0(n303), .B1(n661), .Y(n1632) );
  OAI22X1 U478 ( .A0(n308), .A1(n661), .B0(n1732), .B1(n660), .Y(n1616) );
  OAI22X1 U479 ( .A0(n309), .A1(n655), .B0(n304), .B1(n654), .Y(n1649) );
  OAI22X1 U480 ( .A0(n1733), .A1(n654), .B0(n303), .B1(n653), .Y(n1633) );
  OAI22X1 U481 ( .A0(n310), .A1(n653), .B0(n1732), .B1(n652), .Y(n1617) );
  OAI22X1 U482 ( .A0(n310), .A1(n647), .B0(n305), .B1(n646), .Y(n1650) );
  OAI22X1 U483 ( .A0(n308), .A1(n646), .B0(n303), .B1(n645), .Y(n1634) );
  OAI22X1 U484 ( .A0(n311), .A1(n645), .B0(n1732), .B1(n644), .Y(n1618) );
  OAI22X1 U485 ( .A0(n311), .A1(n639), .B0(n306), .B1(n638), .Y(n1651) );
  OAI22X1 U486 ( .A0(n311), .A1(n638), .B0(n303), .B1(n637), .Y(n1635) );
  OAI22X1 U487 ( .A0(n1733), .A1(n637), .B0(n1732), .B1(n636), .Y(n1619) );
  OAI22X1 U488 ( .A0(n310), .A1(n631), .B0(n1732), .B1(n630), .Y(n1652) );
  OAI22X1 U489 ( .A0(n308), .A1(n630), .B0(n303), .B1(n629), .Y(n1636) );
  OAI22X1 U490 ( .A0(n1733), .A1(n629), .B0(n1732), .B1(n628), .Y(n1620) );
  OAI22X1 U491 ( .A0(n310), .A1(n623), .B0(n1732), .B1(n622), .Y(n1653) );
  OAI22X1 U492 ( .A0(n310), .A1(n622), .B0(n303), .B1(n621), .Y(n1637) );
  OAI22X1 U493 ( .A0(n1733), .A1(n621), .B0(n1732), .B1(n620), .Y(n1621) );
  OAI22X1 U494 ( .A0(n311), .A1(n615), .B0(n1732), .B1(n614), .Y(n1654) );
  OAI22X1 U495 ( .A0(n614), .A1(n1733), .B0(n303), .B1(n613), .Y(n1638) );
  OAI22X1 U496 ( .A0(n1733), .A1(n613), .B0(n1732), .B1(n612), .Y(n1622) );
  OAI22X1 U497 ( .A0(n292), .A1(n607), .B0(n279), .B1(n606), .Y(n1511) );
  OAI22X1 U498 ( .A0(n299), .A1(n606), .B0(n284), .B1(n605), .Y(n1495) );
  OAI22X1 U499 ( .A0(n300), .A1(n605), .B0(n279), .B1(n604), .Y(n1479) );
  OAI22X1 U500 ( .A0(n298), .A1(n591), .B0(n281), .B1(n590), .Y(n1512) );
  OAI22X1 U501 ( .A0(n294), .A1(n590), .B0(n281), .B1(n589), .Y(n1496) );
  OAI22X1 U502 ( .A0(n290), .A1(n589), .B0(n279), .B1(n588), .Y(n1480) );
  OAI22X1 U503 ( .A0(n290), .A1(n575), .B0(n282), .B1(n574), .Y(n1513) );
  OAI22X1 U504 ( .A0(n290), .A1(n574), .B0(n279), .B1(n573), .Y(n1497) );
  OAI22X1 U505 ( .A0(n298), .A1(n573), .B0(n279), .B1(n572), .Y(n1481) );
  OAI22X1 U506 ( .A0(n297), .A1(n559), .B0(n278), .B1(n558), .Y(n1514) );
  OAI22X1 U507 ( .A0(n296), .A1(n558), .B0(n281), .B1(n557), .Y(n1498) );
  OAI22X1 U508 ( .A0(n299), .A1(n557), .B0(n279), .B1(n556), .Y(n1482) );
  OAI22X1 U509 ( .A0(n293), .A1(n543), .B0(n278), .B1(n542), .Y(n1515) );
  OAI22X1 U510 ( .A0(n291), .A1(n542), .B0(n288), .B1(n541), .Y(n1499) );
  OAI22X1 U511 ( .A0(n302), .A1(n541), .B0(n279), .B1(n540), .Y(n1483) );
  OAI22X1 U512 ( .A0(n289), .A1(n527), .B0(n278), .B1(n526), .Y(n1516) );
  OAI22X1 U513 ( .A0(n298), .A1(n526), .B0(n278), .B1(n525), .Y(n1500) );
  OAI22X1 U514 ( .A0(n300), .A1(n525), .B0(n279), .B1(n524), .Y(n1484) );
  OAI22X1 U515 ( .A0(n295), .A1(n511), .B0(n278), .B1(n510), .Y(n1517) );
  OAI22X1 U516 ( .A0(n293), .A1(n510), .B0(n288), .B1(n509), .Y(n1501) );
  OAI22X1 U517 ( .A0(n300), .A1(n509), .B0(n279), .B1(n508), .Y(n1485) );
  OAI22X1 U518 ( .A0(n299), .A1(n495), .B0(n278), .B1(n494), .Y(n1518) );
  OAI22X1 U519 ( .A0(n302), .A1(n494), .B0(n278), .B1(n493), .Y(n1502) );
  OAI22X1 U520 ( .A0(n301), .A1(n493), .B0(n279), .B1(n492), .Y(n1486) );
  OAI22X1 U521 ( .A0(n290), .A1(n479), .B0(n278), .B1(n478), .Y(n1519) );
  OAI22X1 U522 ( .A0(n296), .A1(n478), .B0(n280), .B1(n477), .Y(n1503) );
  OAI22X1 U523 ( .A0(n292), .A1(n477), .B0(n279), .B1(n476), .Y(n1487) );
  OAI22X1 U524 ( .A0(n302), .A1(n463), .B0(n278), .B1(n462), .Y(n1520) );
  OAI22X1 U525 ( .A0(n294), .A1(n462), .B0(n284), .B1(n461), .Y(n1504) );
  OAI22X1 U526 ( .A0(n296), .A1(n461), .B0(n287), .B1(n460), .Y(n1488) );
  OAI22X1 U527 ( .A0(n294), .A1(n447), .B0(n278), .B1(n446), .Y(n1521) );
  OAI22X1 U528 ( .A0(n299), .A1(n446), .B0(n283), .B1(n445), .Y(n1505) );
  OAI22X1 U529 ( .A0(n295), .A1(n445), .B0(n282), .B1(n444), .Y(n1489) );
  OAI22X1 U530 ( .A0(n300), .A1(n431), .B0(n278), .B1(n430), .Y(n1522) );
  OAI22X1 U531 ( .A0(n300), .A1(n430), .B0(n288), .B1(n429), .Y(n1506) );
  OAI22X1 U532 ( .A0(n299), .A1(n429), .B0(n284), .B1(n428), .Y(n1490) );
  OAI22X1 U533 ( .A0(n298), .A1(n415), .B0(n278), .B1(n414), .Y(n1523) );
  OAI22X1 U534 ( .A0(n301), .A1(n414), .B0(n278), .B1(n413), .Y(n1507) );
  OAI22X1 U535 ( .A0(n297), .A1(n413), .B0(n280), .B1(n412), .Y(n1491) );
  OAI22X1 U536 ( .A0(n297), .A1(n399), .B0(n278), .B1(n398), .Y(n1524) );
  OAI22X1 U537 ( .A0(n292), .A1(n398), .B0(n280), .B1(n397), .Y(n1508) );
  OAI22X1 U538 ( .A0(n293), .A1(n397), .B0(n285), .B1(n396), .Y(n1492) );
  OAI22X1 U539 ( .A0(n291), .A1(n383), .B0(n278), .B1(n382), .Y(n1525) );
  OAI22X1 U540 ( .A0(n290), .A1(n382), .B0(n284), .B1(n381), .Y(n1509) );
  OAI22X1 U541 ( .A0(n298), .A1(n381), .B0(n286), .B1(n380), .Y(n1493) );
  OAI22X1 U542 ( .A0(n299), .A1(n367), .B0(n278), .B1(n366), .Y(n1526) );
  OAI22X1 U543 ( .A0(n366), .A1(n291), .B0(n287), .B1(n365), .Y(n1510) );
  OAI22X1 U544 ( .A0(n297), .A1(n365), .B0(n280), .B1(n364), .Y(n1494) );
  NAND2X1 U545 ( .A(n1731), .B(start), .Y(n1732) );
  NAND2X1 U546 ( .A(n1730), .B(n1266), .Y(n1733) );
  NOR2BX1 U547 ( .AN(N304), .B(n1721), .Y(N1117) );
  NOR2BX1 U548 ( .AN(N303), .B(n1721), .Y(N1116) );
  NOR2BX1 U549 ( .AN(N302), .B(n1721), .Y(N1115) );
  INVX1 U550 ( .A(n1731), .Y(n1266) );
  INVX1 U551 ( .A(n1729), .Y(n1268) );
  NOR2X1 U552 ( .A(n1725), .B(n1265), .Y(N1119) );
  AOI222X1 U553 ( .A0(n1724), .A1(n1734), .B0(n1723), .B1(n1729), .C0(n1722), 
        .C1(n1731), .Y(n1725) );
  INVX1 U554 ( .A(n1734), .Y(n1269) );
  OAI222XL U555 ( .A0(n604), .A1(n274), .B0(n1261), .B1(n266), .C0(n738), .C1(
        n262), .Y(N224) );
  OAI222XL U556 ( .A0(n605), .A1(n276), .B0(n1262), .B1(n1727), .C0(n739), 
        .C1(n264), .Y(N241) );
  OAI222XL U557 ( .A0(n606), .A1(n276), .B0(n1263), .B1(n266), .C0(n1199), 
        .C1(n264), .Y(N257) );
  OAI222XL U558 ( .A0(n607), .A1(n275), .B0(n1264), .B1(n267), .C0(n1200), 
        .C1(n264), .Y(N273) );
  OAI222XL U559 ( .A0(n588), .A1(n274), .B0(n1257), .B1(n266), .C0(n724), .C1(
        n1726), .Y(N225) );
  OAI222XL U560 ( .A0(n589), .A1(n276), .B0(n1258), .B1(n267), .C0(n725), .C1(
        n264), .Y(N242) );
  OAI222XL U561 ( .A0(n590), .A1(n276), .B0(n1259), .B1(n266), .C0(n726), .C1(
        n264), .Y(N258) );
  OAI222XL U562 ( .A0(n591), .A1(n275), .B0(n1260), .B1(n267), .C0(n727), .C1(
        n263), .Y(N274) );
  OAI222XL U563 ( .A0(n572), .A1(n274), .B0(n1253), .B1(n266), .C0(n716), .C1(
        n264), .Y(N226) );
  OAI222XL U564 ( .A0(n573), .A1(n276), .B0(n1254), .B1(n266), .C0(n717), .C1(
        n264), .Y(N243) );
  OAI222XL U565 ( .A0(n574), .A1(n275), .B0(n1255), .B1(n1727), .C0(n718), 
        .C1(n264), .Y(N259) );
  OAI222XL U566 ( .A0(n575), .A1(n275), .B0(n1256), .B1(n267), .C0(n719), .C1(
        n261), .Y(N275) );
  OAI222XL U567 ( .A0(n556), .A1(n274), .B0(n1249), .B1(n266), .C0(n708), .C1(
        n263), .Y(N227) );
  OAI222XL U568 ( .A0(n557), .A1(n276), .B0(n1250), .B1(n1727), .C0(n709), 
        .C1(n264), .Y(N244) );
  OAI222XL U569 ( .A0(n558), .A1(n275), .B0(n1251), .B1(n267), .C0(n710), .C1(
        n262), .Y(N260) );
  OAI222XL U570 ( .A0(n559), .A1(n275), .B0(n1252), .B1(n267), .C0(n711), .C1(
        n264), .Y(N276) );
  OAI222XL U571 ( .A0(n540), .A1(n274), .B0(n1245), .B1(n266), .C0(n700), .C1(
        n261), .Y(N228) );
  OAI222XL U572 ( .A0(n541), .A1(n276), .B0(n1246), .B1(n267), .C0(n701), .C1(
        n264), .Y(N245) );
  OAI222XL U573 ( .A0(n542), .A1(n275), .B0(n1247), .B1(n1727), .C0(n702), 
        .C1(n264), .Y(N261) );
  OAI222XL U574 ( .A0(n543), .A1(n275), .B0(n1248), .B1(n267), .C0(n703), .C1(
        n263), .Y(N277) );
  OAI222XL U575 ( .A0(n524), .A1(n274), .B0(n1241), .B1(n266), .C0(n692), .C1(
        n262), .Y(N229) );
  OAI222XL U576 ( .A0(n525), .A1(n276), .B0(n1242), .B1(n266), .C0(n693), .C1(
        n264), .Y(N246) );
  OAI222XL U577 ( .A0(n526), .A1(n275), .B0(n1243), .B1(n1727), .C0(n694), 
        .C1(n261), .Y(N262) );
  OAI222XL U578 ( .A0(n527), .A1(n275), .B0(n1244), .B1(n267), .C0(n695), .C1(
        n262), .Y(N278) );
  OAI222XL U579 ( .A0(n508), .A1(n274), .B0(n1237), .B1(n266), .C0(n684), .C1(
        n1726), .Y(N231) );
  OAI222XL U580 ( .A0(n509), .A1(n276), .B0(n1238), .B1(n1727), .C0(n685), 
        .C1(n264), .Y(N247) );
  OAI222XL U581 ( .A0(n510), .A1(n275), .B0(n1239), .B1(n1727), .C0(n686), 
        .C1(n1726), .Y(N263) );
  OAI222XL U582 ( .A0(n511), .A1(n275), .B0(n1240), .B1(n267), .C0(n687), .C1(
        n263), .Y(N279) );
  OAI222XL U583 ( .A0(n492), .A1(n274), .B0(n1233), .B1(n266), .C0(n676), .C1(
        n264), .Y(N232) );
  OAI222XL U584 ( .A0(n493), .A1(n276), .B0(n1234), .B1(n267), .C0(n677), .C1(
        n264), .Y(N248) );
  OAI222XL U585 ( .A0(n494), .A1(n275), .B0(n1235), .B1(n1727), .C0(n678), 
        .C1(n264), .Y(N264) );
  OAI222XL U586 ( .A0(n495), .A1(n275), .B0(n1236), .B1(n267), .C0(n679), .C1(
        n263), .Y(N280) );
  OAI222XL U587 ( .A0(n476), .A1(n274), .B0(n1229), .B1(n266), .C0(n668), .C1(
        n263), .Y(N233) );
  OAI222XL U588 ( .A0(n477), .A1(n276), .B0(n1230), .B1(n266), .C0(n669), .C1(
        n264), .Y(N249) );
  OAI222XL U589 ( .A0(n478), .A1(n274), .B0(n1231), .B1(n1727), .C0(n670), 
        .C1(n261), .Y(N265) );
  OAI222XL U590 ( .A0(n479), .A1(n275), .B0(n1232), .B1(n267), .C0(n671), .C1(
        n1726), .Y(N281) );
  OAI222XL U591 ( .A0(n460), .A1(n274), .B0(n1225), .B1(n266), .C0(n660), .C1(
        n261), .Y(N234) );
  OAI222XL U592 ( .A0(n461), .A1(n276), .B0(n1226), .B1(n1727), .C0(n661), 
        .C1(n264), .Y(N250) );
  OAI222XL U593 ( .A0(n462), .A1(n275), .B0(n1227), .B1(n1727), .C0(n662), 
        .C1(n262), .Y(N266) );
  OAI222XL U594 ( .A0(n463), .A1(n274), .B0(n1228), .B1(n267), .C0(n663), .C1(
        n1726), .Y(N282) );
  OAI222XL U595 ( .A0(n444), .A1(n274), .B0(n1221), .B1(n266), .C0(n652), .C1(
        n262), .Y(N235) );
  OAI222XL U596 ( .A0(n445), .A1(n276), .B0(n1222), .B1(n1727), .C0(n653), 
        .C1(n264), .Y(N251) );
  OAI222XL U597 ( .A0(n446), .A1(n275), .B0(n1223), .B1(n1727), .C0(n654), 
        .C1(n1726), .Y(N267) );
  OAI222XL U598 ( .A0(n447), .A1(n274), .B0(n1224), .B1(n267), .C0(n655), .C1(
        n1726), .Y(N283) );
  OAI222XL U599 ( .A0(n428), .A1(n274), .B0(n1217), .B1(n266), .C0(n644), .C1(
        n1726), .Y(N236) );
  OAI222XL U600 ( .A0(n429), .A1(n276), .B0(n1218), .B1(n267), .C0(n645), .C1(
        n264), .Y(N252) );
  OAI222XL U601 ( .A0(n430), .A1(n275), .B0(n1219), .B1(n267), .C0(n646), .C1(
        n261), .Y(N268) );
  OAI222XL U602 ( .A0(n431), .A1(n274), .B0(n1220), .B1(n267), .C0(n647), .C1(
        n1726), .Y(N284) );
  OAI222XL U603 ( .A0(n412), .A1(n276), .B0(n1213), .B1(n266), .C0(n636), .C1(
        n264), .Y(N237) );
  OAI222XL U604 ( .A0(n413), .A1(n276), .B0(n1214), .B1(n266), .C0(n637), .C1(
        n264), .Y(N253) );
  OAI222XL U605 ( .A0(n414), .A1(n275), .B0(n1215), .B1(n266), .C0(n638), .C1(
        n264), .Y(N269) );
  OAI222XL U606 ( .A0(n415), .A1(n274), .B0(n1216), .B1(n1727), .C0(n639), 
        .C1(n1726), .Y(N285) );
  OAI222XL U607 ( .A0(n396), .A1(n276), .B0(n1209), .B1(n1727), .C0(n628), 
        .C1(n263), .Y(N238) );
  OAI222XL U608 ( .A0(n397), .A1(n276), .B0(n1210), .B1(n267), .C0(n629), .C1(
        n264), .Y(N254) );
  OAI222XL U609 ( .A0(n398), .A1(n275), .B0(n1211), .B1(n266), .C0(n630), .C1(
        n263), .Y(N270) );
  OAI222XL U610 ( .A0(n399), .A1(n274), .B0(n1212), .B1(n1727), .C0(n631), 
        .C1(n1726), .Y(N286) );
  OAI222XL U611 ( .A0(n380), .A1(n276), .B0(n1205), .B1(n267), .C0(n620), .C1(
        n264), .Y(N239) );
  OAI222XL U612 ( .A0(n381), .A1(n276), .B0(n1206), .B1(n1727), .C0(n621), 
        .C1(n264), .Y(N255) );
  OAI222XL U613 ( .A0(n382), .A1(n275), .B0(n1207), .B1(n267), .C0(n622), .C1(
        n261), .Y(N271) );
  OAI222XL U614 ( .A0(n383), .A1(n274), .B0(n1208), .B1(n1727), .C0(n623), 
        .C1(n1726), .Y(N287) );
  OAI222XL U615 ( .A0(n364), .A1(n276), .B0(n1201), .B1(n266), .C0(n612), .C1(
        n264), .Y(N240) );
  OAI222XL U616 ( .A0(n365), .A1(n276), .B0(n1202), .B1(n267), .C0(n613), .C1(
        n264), .Y(N256) );
  OAI222XL U617 ( .A0(n366), .A1(n275), .B0(n1203), .B1(n1727), .C0(n614), 
        .C1(n262), .Y(N272) );
  OAI222XL U618 ( .A0(n367), .A1(n274), .B0(n1204), .B1(n1727), .C0(n615), 
        .C1(n1726), .Y(N288) );
  OAI21XL U619 ( .A0(n349), .A1(n348), .B0(n351), .Y(N30) );
  OAI22X1 U620 ( .A0(n728), .A1(n261), .B0(n600), .B1(n270), .Y(N160) );
  OAI22X1 U621 ( .A0(n729), .A1(n262), .B0(n601), .B1(n273), .Y(N176) );
  OAI22X1 U622 ( .A0(n730), .A1(n262), .B0(n602), .B1(n1728), .Y(N192) );
  OAI22X1 U623 ( .A0(n732), .A1(n263), .B0(n603), .B1(n270), .Y(N208) );
  OAI22X1 U624 ( .A0(n720), .A1(n261), .B0(n584), .B1(n276), .Y(N161) );
  OAI22X1 U625 ( .A0(n721), .A1(n262), .B0(n585), .B1(n269), .Y(N177) );
  OAI22X1 U626 ( .A0(n722), .A1(n1726), .B0(n586), .B1(n273), .Y(N193) );
  OAI22X1 U627 ( .A0(n723), .A1(n263), .B0(n587), .B1(n270), .Y(N209) );
  OAI22X1 U628 ( .A0(n712), .A1(n261), .B0(n568), .B1(n274), .Y(N162) );
  OAI22X1 U629 ( .A0(n713), .A1(n262), .B0(n569), .B1(n274), .Y(N178) );
  OAI22X1 U630 ( .A0(n714), .A1(n263), .B0(n570), .B1(n272), .Y(N194) );
  OAI22X1 U631 ( .A0(n715), .A1(n263), .B0(n571), .B1(n270), .Y(N210) );
  OAI22X1 U632 ( .A0(n704), .A1(n261), .B0(n552), .B1(n1728), .Y(N163) );
  OAI22X1 U633 ( .A0(n705), .A1(n262), .B0(n553), .B1(n1728), .Y(N179) );
  OAI22X1 U634 ( .A0(n706), .A1(n261), .B0(n554), .B1(n273), .Y(N195) );
  OAI22X1 U635 ( .A0(n707), .A1(n263), .B0(n555), .B1(n269), .Y(N211) );
  OAI22X1 U636 ( .A0(n696), .A1(n261), .B0(n536), .B1(n275), .Y(N164) );
  OAI22X1 U637 ( .A0(n697), .A1(n262), .B0(n537), .B1(n272), .Y(N180) );
  OAI22X1 U638 ( .A0(n698), .A1(n1726), .B0(n538), .B1(n271), .Y(N196) );
  OAI22X1 U639 ( .A0(n699), .A1(n263), .B0(n539), .B1(n269), .Y(N212) );
  OAI22X1 U640 ( .A0(n688), .A1(n261), .B0(n520), .B1(n271), .Y(N165) );
  OAI22X1 U641 ( .A0(n689), .A1(n262), .B0(n521), .B1(n271), .Y(N181) );
  OAI22X1 U642 ( .A0(n690), .A1(n1726), .B0(n522), .B1(n276), .Y(N197) );
  OAI22X1 U643 ( .A0(n691), .A1(n263), .B0(n523), .B1(n269), .Y(N213) );
  OAI22X1 U644 ( .A0(n680), .A1(n261), .B0(n504), .B1(n271), .Y(N166) );
  OAI22X1 U645 ( .A0(n681), .A1(n262), .B0(n505), .B1(n270), .Y(N182) );
  OAI22X1 U646 ( .A0(n682), .A1(n1726), .B0(n506), .B1(n270), .Y(N198) );
  OAI22X1 U647 ( .A0(n683), .A1(n263), .B0(n507), .B1(n269), .Y(N214) );
  OAI22X1 U648 ( .A0(n672), .A1(n261), .B0(n488), .B1(n276), .Y(N167) );
  OAI22X1 U649 ( .A0(n673), .A1(n262), .B0(n489), .B1(n276), .Y(N183) );
  OAI22X1 U650 ( .A0(n674), .A1(n1726), .B0(n490), .B1(n270), .Y(N199) );
  OAI22X1 U651 ( .A0(n675), .A1(n263), .B0(n491), .B1(n269), .Y(N215) );
  OAI22X1 U652 ( .A0(n664), .A1(n261), .B0(n472), .B1(n275), .Y(N168) );
  OAI22X1 U653 ( .A0(n665), .A1(n262), .B0(n473), .B1(n275), .Y(N184) );
  OAI22X1 U654 ( .A0(n666), .A1(n1726), .B0(n474), .B1(n270), .Y(N200) );
  OAI22X1 U655 ( .A0(n667), .A1(n263), .B0(n475), .B1(n269), .Y(N216) );
  OAI22X1 U656 ( .A0(n656), .A1(n261), .B0(n456), .B1(n273), .Y(N169) );
  OAI22X1 U657 ( .A0(n657), .A1(n1726), .B0(n457), .B1(n269), .Y(N185) );
  OAI22X1 U658 ( .A0(n658), .A1(n1726), .B0(n458), .B1(n270), .Y(N201) );
  OAI22X1 U659 ( .A0(n659), .A1(n263), .B0(n459), .B1(n269), .Y(N217) );
  OAI22X1 U660 ( .A0(n648), .A1(n261), .B0(n440), .B1(n272), .Y(N170) );
  OAI22X1 U661 ( .A0(n649), .A1(n1726), .B0(n441), .B1(n269), .Y(N186) );
  OAI22X1 U662 ( .A0(n650), .A1(n263), .B0(n442), .B1(n270), .Y(N202) );
  OAI22X1 U663 ( .A0(n651), .A1(n263), .B0(n443), .B1(n269), .Y(N218) );
  OAI22X1 U664 ( .A0(n640), .A1(n261), .B0(n424), .B1(n269), .Y(N171) );
  OAI22X1 U665 ( .A0(n641), .A1(n263), .B0(n425), .B1(n270), .Y(N187) );
  OAI22X1 U666 ( .A0(n642), .A1(n261), .B0(n426), .B1(n270), .Y(N203) );
  OAI22X1 U667 ( .A0(n643), .A1(n263), .B0(n427), .B1(n269), .Y(N219) );
  OAI22X1 U668 ( .A0(n632), .A1(n262), .B0(n408), .B1(n273), .Y(N172) );
  OAI22X1 U669 ( .A0(n633), .A1(n261), .B0(n409), .B1(n275), .Y(N188) );
  OAI22X1 U670 ( .A0(n634), .A1(n262), .B0(n410), .B1(n270), .Y(N204) );
  OAI22X1 U671 ( .A0(n635), .A1(n263), .B0(n411), .B1(n269), .Y(N220) );
  OAI22X1 U672 ( .A0(n624), .A1(n262), .B0(n392), .B1(n269), .Y(N173) );
  OAI22X1 U673 ( .A0(n625), .A1(n262), .B0(n393), .B1(n1728), .Y(N189) );
  OAI22X1 U674 ( .A0(n626), .A1(n261), .B0(n394), .B1(n270), .Y(N205) );
  OAI22X1 U675 ( .A0(n627), .A1(n261), .B0(n395), .B1(n269), .Y(N221) );
  OAI22X1 U676 ( .A0(n616), .A1(n262), .B0(n376), .B1(n274), .Y(N174) );
  OAI22X1 U677 ( .A0(n617), .A1(n264), .B0(n377), .B1(n273), .Y(N190) );
  OAI22X1 U678 ( .A0(n618), .A1(n1726), .B0(n378), .B1(n270), .Y(N206) );
  OAI22X1 U679 ( .A0(n619), .A1(n262), .B0(n379), .B1(n269), .Y(N222) );
  OAI22X1 U680 ( .A0(n608), .A1(n262), .B0(n360), .B1(n1728), .Y(N175) );
  OAI22X1 U681 ( .A0(n609), .A1(n1726), .B0(n361), .B1(n272), .Y(N191) );
  OAI22X1 U682 ( .A0(n610), .A1(n263), .B0(n362), .B1(n270), .Y(N207) );
  OAI22X1 U683 ( .A0(n611), .A1(n1726), .B0(n363), .B1(n269), .Y(N223) );
  NOR2X1 U684 ( .A(n592), .B(n271), .Y(N31) );
  NOR2X1 U685 ( .A(n593), .B(n271), .Y(N47) );
  NOR2X1 U686 ( .A(n594), .B(n272), .Y(N63) );
  NOR2X1 U687 ( .A(n595), .B(n269), .Y(N79) );
  NOR2X1 U688 ( .A(n596), .B(n269), .Y(N95) );
  NOR2X1 U689 ( .A(n597), .B(n276), .Y(N111) );
  NOR2X1 U690 ( .A(n598), .B(n273), .Y(N127) );
  NOR2X1 U691 ( .A(n599), .B(n1728), .Y(N144) );
  NOR2X1 U692 ( .A(n576), .B(n1728), .Y(N32) );
  NOR2X1 U693 ( .A(n577), .B(n271), .Y(N48) );
  NOR2X1 U694 ( .A(n578), .B(n272), .Y(N64) );
  NOR2X1 U695 ( .A(n579), .B(n274), .Y(N80) );
  NOR2X1 U696 ( .A(n580), .B(n270), .Y(N96) );
  NOR2X1 U697 ( .A(n581), .B(n271), .Y(N112) );
  NOR2X1 U698 ( .A(n582), .B(n273), .Y(N128) );
  NOR2X1 U699 ( .A(n583), .B(n1728), .Y(N145) );
  NOR2X1 U700 ( .A(n560), .B(n272), .Y(N33) );
  NOR2X1 U701 ( .A(n561), .B(n271), .Y(N49) );
  NOR2X1 U702 ( .A(n562), .B(n272), .Y(N65) );
  NOR2X1 U703 ( .A(n563), .B(n1728), .Y(N81) );
  NOR2X1 U704 ( .A(n564), .B(n271), .Y(N97) );
  NOR2X1 U705 ( .A(n565), .B(n270), .Y(N113) );
  NOR2X1 U706 ( .A(n566), .B(n273), .Y(N129) );
  NOR2X1 U707 ( .A(n567), .B(n1728), .Y(N146) );
  NOR2X1 U708 ( .A(n544), .B(n271), .Y(N34) );
  NOR2X1 U709 ( .A(n545), .B(n271), .Y(N50) );
  NOR2X1 U710 ( .A(n546), .B(n272), .Y(N66) );
  NOR2X1 U711 ( .A(n547), .B(n272), .Y(N82) );
  NOR2X1 U712 ( .A(n548), .B(n276), .Y(N98) );
  NOR2X1 U713 ( .A(n549), .B(n270), .Y(N114) );
  NOR2X1 U714 ( .A(n550), .B(n273), .Y(N131) );
  NOR2X1 U715 ( .A(n551), .B(n1728), .Y(N147) );
  NOR2X1 U716 ( .A(n528), .B(n275), .Y(N35) );
  NOR2X1 U717 ( .A(n529), .B(n271), .Y(N51) );
  NOR2X1 U718 ( .A(n530), .B(n272), .Y(N67) );
  NOR2X1 U719 ( .A(n531), .B(n273), .Y(N83) );
  NOR2X1 U720 ( .A(n532), .B(n273), .Y(N99) );
  NOR2X1 U721 ( .A(n533), .B(n273), .Y(N115) );
  NOR2X1 U722 ( .A(n534), .B(n272), .Y(N132) );
  NOR2X1 U723 ( .A(n535), .B(n1728), .Y(N148) );
  NOR2X1 U724 ( .A(n512), .B(n269), .Y(N36) );
  NOR2X1 U725 ( .A(n513), .B(n271), .Y(N52) );
  NOR2X1 U726 ( .A(n514), .B(n272), .Y(N68) );
  NOR2X1 U727 ( .A(n515), .B(n270), .Y(N84) );
  NOR2X1 U728 ( .A(n516), .B(n274), .Y(N100) );
  NOR2X1 U729 ( .A(n517), .B(n273), .Y(N116) );
  NOR2X1 U730 ( .A(n518), .B(n272), .Y(N133) );
  NOR2X1 U731 ( .A(n519), .B(n274), .Y(N149) );
  NOR2X1 U732 ( .A(n496), .B(n1728), .Y(N37) );
  NOR2X1 U733 ( .A(n497), .B(n271), .Y(N53) );
  NOR2X1 U734 ( .A(n498), .B(n275), .Y(N69) );
  NOR2X1 U735 ( .A(n499), .B(n1728), .Y(N85) );
  NOR2X1 U736 ( .A(n500), .B(n271), .Y(N101) );
  NOR2X1 U737 ( .A(n501), .B(n273), .Y(N117) );
  NOR2X1 U738 ( .A(n502), .B(n270), .Y(N134) );
  NOR2X1 U739 ( .A(n503), .B(n1728), .Y(N150) );
  NOR2X1 U740 ( .A(n480), .B(n272), .Y(N38) );
  NOR2X1 U741 ( .A(n481), .B(n271), .Y(N54) );
  NOR2X1 U742 ( .A(n482), .B(n273), .Y(N70) );
  NOR2X1 U743 ( .A(n483), .B(n273), .Y(N86) );
  NOR2X1 U744 ( .A(n484), .B(n274), .Y(N102) );
  NOR2X1 U745 ( .A(n485), .B(n273), .Y(N118) );
  NOR2X1 U746 ( .A(n486), .B(n270), .Y(N135) );
  NOR2X1 U747 ( .A(n487), .B(n1728), .Y(N151) );
  NOR2X1 U748 ( .A(n464), .B(n271), .Y(N39) );
  NOR2X1 U749 ( .A(n465), .B(n272), .Y(N55) );
  NOR2X1 U750 ( .A(n466), .B(n272), .Y(N71) );
  NOR2X1 U751 ( .A(n467), .B(n272), .Y(N87) );
  NOR2X1 U752 ( .A(n468), .B(n269), .Y(N103) );
  NOR2X1 U753 ( .A(n469), .B(n273), .Y(N119) );
  NOR2X1 U754 ( .A(n470), .B(n1728), .Y(N136) );
  NOR2X1 U755 ( .A(n471), .B(n1728), .Y(N152) );
  NOR2X1 U756 ( .A(n448), .B(n270), .Y(N40) );
  NOR2X1 U757 ( .A(n449), .B(n272), .Y(N56) );
  NOR2X1 U758 ( .A(n450), .B(n271), .Y(N72) );
  NOR2X1 U759 ( .A(n451), .B(n272), .Y(N88) );
  NOR2X1 U760 ( .A(n452), .B(n270), .Y(N104) );
  NOR2X1 U761 ( .A(n453), .B(n273), .Y(N120) );
  NOR2X1 U762 ( .A(n454), .B(n273), .Y(N137) );
  NOR2X1 U763 ( .A(n455), .B(n1728), .Y(N153) );
  NOR2X1 U764 ( .A(n432), .B(n271), .Y(N41) );
  NOR2X1 U765 ( .A(n433), .B(n272), .Y(N57) );
  NOR2X1 U766 ( .A(n434), .B(n270), .Y(N73) );
  NOR2X1 U767 ( .A(n435), .B(n271), .Y(N89) );
  NOR2X1 U768 ( .A(n436), .B(n274), .Y(N105) );
  NOR2X1 U769 ( .A(n437), .B(n273), .Y(N121) );
  NOR2X1 U770 ( .A(n438), .B(n269), .Y(N138) );
  NOR2X1 U771 ( .A(n439), .B(n1728), .Y(N154) );
  NOR2X1 U772 ( .A(n416), .B(n271), .Y(N42) );
  NOR2X1 U773 ( .A(n417), .B(n272), .Y(N58) );
  NOR2X1 U774 ( .A(n418), .B(n276), .Y(N74) );
  NOR2X1 U775 ( .A(n419), .B(n272), .Y(N90) );
  NOR2X1 U776 ( .A(n420), .B(n271), .Y(N106) );
  NOR2X1 U777 ( .A(n421), .B(n273), .Y(N122) );
  NOR2X1 U778 ( .A(n422), .B(n270), .Y(N139) );
  NOR2X1 U779 ( .A(n423), .B(n1728), .Y(N155) );
  NOR2X1 U780 ( .A(n400), .B(n271), .Y(N43) );
  NOR2X1 U781 ( .A(n401), .B(n272), .Y(N59) );
  NOR2X1 U782 ( .A(n402), .B(n276), .Y(N75) );
  NOR2X1 U783 ( .A(n403), .B(n275), .Y(N91) );
  NOR2X1 U784 ( .A(n404), .B(n1728), .Y(N107) );
  NOR2X1 U785 ( .A(n405), .B(n273), .Y(N123) );
  NOR2X1 U786 ( .A(n406), .B(n1728), .Y(N140) );
  NOR2X1 U787 ( .A(n407), .B(n1728), .Y(N156) );
  NOR2X1 U788 ( .A(n384), .B(n271), .Y(N44) );
  NOR2X1 U789 ( .A(n385), .B(n272), .Y(N60) );
  NOR2X1 U790 ( .A(n386), .B(n269), .Y(N76) );
  NOR2X1 U791 ( .A(n387), .B(n269), .Y(N92) );
  NOR2X1 U792 ( .A(n388), .B(n273), .Y(N108) );
  NOR2X1 U793 ( .A(n389), .B(n273), .Y(N124) );
  NOR2X1 U794 ( .A(n390), .B(n275), .Y(N141) );
  NOR2X1 U795 ( .A(n391), .B(n1728), .Y(N157) );
  NOR2X1 U796 ( .A(n368), .B(n271), .Y(N45) );
  NOR2X1 U797 ( .A(n369), .B(n272), .Y(N61) );
  NOR2X1 U798 ( .A(n370), .B(n274), .Y(N77) );
  NOR2X1 U799 ( .A(n371), .B(n270), .Y(N93) );
  NOR2X1 U800 ( .A(n372), .B(n272), .Y(N109) );
  NOR2X1 U801 ( .A(n373), .B(n269), .Y(N125) );
  NOR2X1 U802 ( .A(n374), .B(n1728), .Y(N142) );
  NOR2X1 U803 ( .A(n375), .B(n274), .Y(N158) );
  NOR2X1 U804 ( .A(n352), .B(n271), .Y(N46) );
  NOR2X1 U805 ( .A(n353), .B(n272), .Y(N62) );
  NOR2X1 U806 ( .A(n354), .B(n1728), .Y(N78) );
  NOR2X1 U807 ( .A(n355), .B(n269), .Y(N94) );
  NOR2X1 U808 ( .A(n356), .B(n271), .Y(N110) );
  NOR2X1 U809 ( .A(n357), .B(n273), .Y(N126) );
  NOR2X1 U810 ( .A(n358), .B(n273), .Y(N143) );
  NOR2X1 U811 ( .A(n359), .B(n1728), .Y(N159) );
  NAND2X1 U812 ( .A(n349), .B(n348), .Y(n1727) );
  INVX1 U813 ( .A(n1728), .Y(n277) );
  INVX1 U814 ( .A(n1726), .Y(n265) );
  INVX1 U815 ( .A(s2p_ready), .Y(n351) );
  NOR2X1 U816 ( .A(n1270), .B(mode[0]), .Y(n1729) );
  NOR2X1 U817 ( .A(n1267), .B(mode[1]), .Y(n1731) );
  AOI21X1 U818 ( .A0(mode[0]), .A1(mode[1]), .B0(n1265), .Y(n1730) );
  INVX1 U819 ( .A(mode_reg[0]), .Y(n349) );
  INVX1 U820 ( .A(mode[0]), .Y(n1267) );
  INVX1 U821 ( .A(mode[1]), .Y(n1270) );
  NOR2X1 U822 ( .A(n4), .B(n1721), .Y(N1118) );
  XNOR2X1 U823 ( .A(r71_carry[4]), .B(count[4]), .Y(n4) );
  NOR2X1 U824 ( .A(count[0]), .B(n1721), .Y(N1114) );
  NAND3BX1 U825 ( .AN(count[4]), .B(count[0]), .C(count[1]), .Y(n1719) );
  NOR2X1 U826 ( .A(mode[0]), .B(mode[1]), .Y(n1734) );
  NOR3X1 U827 ( .A(count[2]), .B(count[3]), .C(n1719), .Y(n1724) );
  NOR3X1 U828 ( .A(n1719), .B(count[3]), .C(n350), .Y(n1722) );
  NOR3BX1 U829 ( .AN(count[3]), .B(n350), .C(n1719), .Y(n1723) );
  INVX1 U830 ( .A(dout16_reg[176]), .Y(n603) );
  INVX1 U831 ( .A(dout16_reg[160]), .Y(n602) );
  INVX1 U832 ( .A(dout16_reg[144]), .Y(n601) );
  INVX1 U833 ( .A(dout16_reg[128]), .Y(n600) );
  INVX1 U834 ( .A(dout16_reg[177]), .Y(n587) );
  INVX1 U835 ( .A(dout16_reg[161]), .Y(n586) );
  INVX1 U836 ( .A(dout16_reg[145]), .Y(n585) );
  INVX1 U837 ( .A(dout16_reg[129]), .Y(n584) );
  INVX1 U838 ( .A(dout16_reg[178]), .Y(n571) );
  INVX1 U839 ( .A(dout16_reg[162]), .Y(n570) );
  INVX1 U840 ( .A(dout16_reg[146]), .Y(n569) );
  INVX1 U841 ( .A(dout16_reg[130]), .Y(n568) );
  INVX1 U842 ( .A(dout16_reg[179]), .Y(n555) );
  INVX1 U843 ( .A(dout16_reg[163]), .Y(n554) );
  INVX1 U844 ( .A(dout16_reg[147]), .Y(n553) );
  INVX1 U845 ( .A(dout16_reg[131]), .Y(n552) );
  INVX1 U846 ( .A(dout16_reg[180]), .Y(n539) );
  INVX1 U847 ( .A(dout16_reg[164]), .Y(n538) );
  INVX1 U848 ( .A(dout16_reg[148]), .Y(n537) );
  INVX1 U849 ( .A(dout16_reg[132]), .Y(n536) );
  INVX1 U850 ( .A(dout16_reg[181]), .Y(n523) );
  INVX1 U851 ( .A(dout16_reg[165]), .Y(n522) );
  INVX1 U852 ( .A(dout16_reg[149]), .Y(n521) );
  INVX1 U853 ( .A(dout16_reg[133]), .Y(n520) );
  INVX1 U854 ( .A(dout16_reg[182]), .Y(n507) );
  INVX1 U855 ( .A(dout16_reg[166]), .Y(n506) );
  INVX1 U856 ( .A(dout16_reg[150]), .Y(n505) );
  INVX1 U857 ( .A(dout16_reg[134]), .Y(n504) );
  INVX1 U858 ( .A(dout16_reg[183]), .Y(n491) );
  INVX1 U859 ( .A(dout16_reg[167]), .Y(n490) );
  INVX1 U860 ( .A(dout16_reg[151]), .Y(n489) );
  INVX1 U861 ( .A(dout16_reg[135]), .Y(n488) );
  INVX1 U862 ( .A(dout16_reg[184]), .Y(n475) );
  INVX1 U863 ( .A(dout16_reg[168]), .Y(n474) );
  INVX1 U864 ( .A(dout16_reg[152]), .Y(n473) );
  INVX1 U865 ( .A(dout16_reg[136]), .Y(n472) );
  INVX1 U866 ( .A(dout16_reg[185]), .Y(n459) );
  INVX1 U867 ( .A(dout16_reg[169]), .Y(n458) );
  INVX1 U868 ( .A(dout16_reg[153]), .Y(n457) );
  INVX1 U869 ( .A(dout16_reg[137]), .Y(n456) );
  INVX1 U870 ( .A(dout16_reg[186]), .Y(n443) );
  INVX1 U871 ( .A(dout16_reg[170]), .Y(n442) );
  INVX1 U872 ( .A(dout16_reg[154]), .Y(n441) );
  INVX1 U873 ( .A(dout16_reg[138]), .Y(n440) );
  INVX1 U874 ( .A(dout16_reg[187]), .Y(n427) );
  INVX1 U875 ( .A(dout16_reg[171]), .Y(n426) );
  INVX1 U876 ( .A(dout16_reg[155]), .Y(n425) );
  INVX1 U877 ( .A(dout16_reg[139]), .Y(n424) );
  INVX1 U878 ( .A(dout16_reg[188]), .Y(n411) );
  INVX1 U879 ( .A(dout16_reg[172]), .Y(n410) );
  INVX1 U880 ( .A(dout16_reg[156]), .Y(n409) );
  INVX1 U881 ( .A(dout16_reg[140]), .Y(n408) );
  INVX1 U882 ( .A(dout16_reg[189]), .Y(n395) );
  INVX1 U883 ( .A(dout16_reg[173]), .Y(n394) );
  INVX1 U884 ( .A(dout16_reg[157]), .Y(n393) );
  INVX1 U885 ( .A(dout16_reg[141]), .Y(n392) );
  INVX1 U886 ( .A(dout16_reg[190]), .Y(n379) );
  INVX1 U887 ( .A(dout16_reg[174]), .Y(n378) );
  INVX1 U888 ( .A(dout16_reg[158]), .Y(n377) );
  INVX1 U889 ( .A(dout16_reg[142]), .Y(n376) );
  INVX1 U890 ( .A(dout16_reg[191]), .Y(n363) );
  INVX1 U891 ( .A(dout16_reg[175]), .Y(n362) );
  INVX1 U892 ( .A(dout16_reg[159]), .Y(n361) );
  INVX1 U893 ( .A(dout16_reg[143]), .Y(n360) );
  INVX1 U894 ( .A(dout8_reg[48]), .Y(n732) );
  INVX1 U895 ( .A(dout8_reg[32]), .Y(n730) );
  INVX1 U896 ( .A(dout8_reg[16]), .Y(n729) );
  INVX1 U897 ( .A(dout8_reg[0]), .Y(n728) );
  INVX1 U898 ( .A(dout8_reg[49]), .Y(n723) );
  INVX1 U899 ( .A(dout8_reg[33]), .Y(n722) );
  INVX1 U900 ( .A(dout8_reg[17]), .Y(n721) );
  INVX1 U901 ( .A(dout8_reg[1]), .Y(n720) );
  INVX1 U902 ( .A(dout8_reg[50]), .Y(n715) );
  INVX1 U903 ( .A(dout8_reg[34]), .Y(n714) );
  INVX1 U904 ( .A(dout8_reg[18]), .Y(n713) );
  INVX1 U905 ( .A(dout8_reg[2]), .Y(n712) );
  INVX1 U906 ( .A(dout8_reg[51]), .Y(n707) );
  INVX1 U907 ( .A(dout8_reg[35]), .Y(n706) );
  INVX1 U908 ( .A(dout8_reg[19]), .Y(n705) );
  INVX1 U909 ( .A(dout8_reg[3]), .Y(n704) );
  INVX1 U910 ( .A(dout8_reg[52]), .Y(n699) );
  INVX1 U911 ( .A(dout8_reg[36]), .Y(n698) );
  INVX1 U912 ( .A(dout8_reg[20]), .Y(n697) );
  INVX1 U913 ( .A(dout8_reg[4]), .Y(n696) );
  INVX1 U914 ( .A(dout8_reg[53]), .Y(n691) );
  INVX1 U915 ( .A(dout8_reg[37]), .Y(n690) );
  INVX1 U916 ( .A(dout8_reg[21]), .Y(n689) );
  INVX1 U917 ( .A(dout8_reg[5]), .Y(n688) );
  INVX1 U918 ( .A(dout8_reg[54]), .Y(n683) );
  INVX1 U919 ( .A(dout8_reg[38]), .Y(n682) );
  INVX1 U920 ( .A(dout8_reg[22]), .Y(n681) );
  INVX1 U921 ( .A(dout8_reg[6]), .Y(n680) );
  INVX1 U922 ( .A(dout8_reg[55]), .Y(n675) );
  INVX1 U923 ( .A(dout8_reg[39]), .Y(n674) );
  INVX1 U924 ( .A(dout8_reg[23]), .Y(n673) );
  INVX1 U925 ( .A(dout8_reg[7]), .Y(n672) );
  INVX1 U926 ( .A(dout8_reg[56]), .Y(n667) );
  INVX1 U927 ( .A(dout8_reg[40]), .Y(n666) );
  INVX1 U928 ( .A(dout8_reg[24]), .Y(n665) );
  INVX1 U929 ( .A(dout8_reg[8]), .Y(n664) );
  INVX1 U930 ( .A(dout8_reg[57]), .Y(n659) );
  INVX1 U931 ( .A(dout8_reg[41]), .Y(n658) );
  INVX1 U932 ( .A(dout8_reg[25]), .Y(n657) );
  INVX1 U933 ( .A(dout8_reg[9]), .Y(n656) );
  INVX1 U934 ( .A(dout8_reg[58]), .Y(n651) );
  INVX1 U935 ( .A(dout8_reg[42]), .Y(n650) );
  INVX1 U936 ( .A(dout8_reg[26]), .Y(n649) );
  INVX1 U937 ( .A(dout8_reg[10]), .Y(n648) );
  INVX1 U938 ( .A(dout8_reg[59]), .Y(n643) );
  INVX1 U939 ( .A(dout8_reg[43]), .Y(n642) );
  INVX1 U940 ( .A(dout8_reg[27]), .Y(n641) );
  INVX1 U941 ( .A(dout8_reg[11]), .Y(n640) );
  INVX1 U942 ( .A(dout8_reg[60]), .Y(n635) );
  INVX1 U943 ( .A(dout8_reg[44]), .Y(n634) );
  INVX1 U944 ( .A(dout8_reg[28]), .Y(n633) );
  INVX1 U945 ( .A(dout8_reg[12]), .Y(n632) );
  INVX1 U946 ( .A(dout8_reg[61]), .Y(n627) );
  INVX1 U947 ( .A(dout8_reg[45]), .Y(n626) );
  INVX1 U948 ( .A(dout8_reg[29]), .Y(n625) );
  INVX1 U949 ( .A(dout8_reg[13]), .Y(n624) );
  INVX1 U950 ( .A(dout8_reg[62]), .Y(n619) );
  INVX1 U951 ( .A(dout8_reg[46]), .Y(n618) );
  INVX1 U952 ( .A(dout8_reg[30]), .Y(n617) );
  INVX1 U953 ( .A(dout8_reg[14]), .Y(n616) );
  INVX1 U954 ( .A(dout8_reg[63]), .Y(n611) );
  INVX1 U955 ( .A(dout8_reg[47]), .Y(n610) );
  INVX1 U956 ( .A(dout8_reg[31]), .Y(n609) );
  INVX1 U957 ( .A(dout8_reg[15]), .Y(n608) );
  INVX1 U958 ( .A(dout16_reg[112]), .Y(n599) );
  INVX1 U959 ( .A(dout16_reg[96]), .Y(n598) );
  INVX1 U960 ( .A(dout16_reg[80]), .Y(n597) );
  INVX1 U961 ( .A(dout16_reg[64]), .Y(n596) );
  INVX1 U962 ( .A(dout16_reg[48]), .Y(n595) );
  INVX1 U963 ( .A(dout16_reg[32]), .Y(n594) );
  INVX1 U964 ( .A(dout16_reg[16]), .Y(n593) );
  INVX1 U965 ( .A(dout16_reg[0]), .Y(n592) );
  INVX1 U966 ( .A(dout16_reg[113]), .Y(n583) );
  INVX1 U967 ( .A(dout16_reg[97]), .Y(n582) );
  INVX1 U968 ( .A(dout16_reg[81]), .Y(n581) );
  INVX1 U969 ( .A(dout16_reg[65]), .Y(n580) );
  INVX1 U970 ( .A(dout16_reg[49]), .Y(n579) );
  INVX1 U971 ( .A(dout16_reg[33]), .Y(n578) );
  INVX1 U972 ( .A(dout16_reg[17]), .Y(n577) );
  INVX1 U973 ( .A(dout16_reg[1]), .Y(n576) );
  INVX1 U974 ( .A(dout16_reg[114]), .Y(n567) );
  INVX1 U975 ( .A(dout16_reg[98]), .Y(n566) );
  INVX1 U976 ( .A(dout16_reg[82]), .Y(n565) );
  INVX1 U977 ( .A(dout16_reg[66]), .Y(n564) );
  INVX1 U978 ( .A(dout16_reg[50]), .Y(n563) );
  INVX1 U979 ( .A(dout16_reg[34]), .Y(n562) );
  INVX1 U980 ( .A(dout16_reg[18]), .Y(n561) );
  INVX1 U981 ( .A(dout16_reg[2]), .Y(n560) );
  INVX1 U982 ( .A(dout16_reg[115]), .Y(n551) );
  INVX1 U983 ( .A(dout16_reg[99]), .Y(n550) );
  INVX1 U984 ( .A(dout16_reg[83]), .Y(n549) );
  INVX1 U985 ( .A(dout16_reg[67]), .Y(n548) );
  INVX1 U986 ( .A(dout16_reg[51]), .Y(n547) );
  INVX1 U987 ( .A(dout16_reg[35]), .Y(n546) );
  INVX1 U988 ( .A(dout16_reg[19]), .Y(n545) );
  INVX1 U989 ( .A(dout16_reg[3]), .Y(n544) );
  INVX1 U990 ( .A(dout16_reg[116]), .Y(n535) );
  INVX1 U991 ( .A(dout16_reg[100]), .Y(n534) );
  INVX1 U992 ( .A(dout16_reg[84]), .Y(n533) );
  INVX1 U993 ( .A(dout16_reg[68]), .Y(n532) );
  INVX1 U994 ( .A(dout16_reg[52]), .Y(n531) );
  INVX1 U995 ( .A(dout16_reg[36]), .Y(n530) );
  INVX1 U996 ( .A(dout16_reg[20]), .Y(n529) );
  INVX1 U997 ( .A(dout16_reg[4]), .Y(n528) );
  INVX1 U998 ( .A(dout16_reg[117]), .Y(n519) );
  INVX1 U999 ( .A(dout16_reg[101]), .Y(n518) );
  INVX1 U1000 ( .A(dout16_reg[85]), .Y(n517) );
  INVX1 U1001 ( .A(dout16_reg[69]), .Y(n516) );
  INVX1 U1002 ( .A(dout16_reg[53]), .Y(n515) );
  INVX1 U1003 ( .A(dout16_reg[37]), .Y(n514) );
  INVX1 U1004 ( .A(dout16_reg[21]), .Y(n513) );
  INVX1 U1005 ( .A(dout16_reg[5]), .Y(n512) );
  INVX1 U1006 ( .A(dout16_reg[118]), .Y(n503) );
  INVX1 U1007 ( .A(dout16_reg[102]), .Y(n502) );
  INVX1 U1008 ( .A(dout16_reg[86]), .Y(n501) );
  INVX1 U1009 ( .A(dout16_reg[70]), .Y(n500) );
  INVX1 U1010 ( .A(dout16_reg[54]), .Y(n499) );
  INVX1 U1011 ( .A(dout16_reg[38]), .Y(n498) );
  INVX1 U1012 ( .A(dout16_reg[22]), .Y(n497) );
  INVX1 U1013 ( .A(dout16_reg[6]), .Y(n496) );
  INVX1 U1014 ( .A(dout16_reg[119]), .Y(n487) );
  INVX1 U1015 ( .A(dout16_reg[103]), .Y(n486) );
  INVX1 U1016 ( .A(dout16_reg[87]), .Y(n485) );
  INVX1 U1017 ( .A(dout16_reg[71]), .Y(n484) );
  INVX1 U1018 ( .A(dout16_reg[55]), .Y(n483) );
  INVX1 U1019 ( .A(dout16_reg[39]), .Y(n482) );
  INVX1 U1020 ( .A(dout16_reg[23]), .Y(n481) );
  INVX1 U1021 ( .A(dout16_reg[7]), .Y(n480) );
  INVX1 U1022 ( .A(dout16_reg[120]), .Y(n471) );
  INVX1 U1023 ( .A(dout16_reg[104]), .Y(n470) );
  INVX1 U1024 ( .A(dout16_reg[88]), .Y(n469) );
  INVX1 U1025 ( .A(dout16_reg[72]), .Y(n468) );
  INVX1 U1026 ( .A(dout16_reg[56]), .Y(n467) );
  INVX1 U1027 ( .A(dout16_reg[40]), .Y(n466) );
  INVX1 U1028 ( .A(dout16_reg[24]), .Y(n465) );
  INVX1 U1029 ( .A(dout16_reg[8]), .Y(n464) );
  INVX1 U1030 ( .A(dout16_reg[121]), .Y(n455) );
  INVX1 U1031 ( .A(dout16_reg[105]), .Y(n454) );
  INVX1 U1032 ( .A(dout16_reg[89]), .Y(n453) );
  INVX1 U1033 ( .A(dout16_reg[73]), .Y(n452) );
  INVX1 U1034 ( .A(dout16_reg[57]), .Y(n451) );
  INVX1 U1035 ( .A(dout16_reg[41]), .Y(n450) );
  INVX1 U1036 ( .A(dout16_reg[25]), .Y(n449) );
  INVX1 U1037 ( .A(dout16_reg[9]), .Y(n448) );
  INVX1 U1038 ( .A(dout16_reg[122]), .Y(n439) );
  INVX1 U1039 ( .A(dout16_reg[106]), .Y(n438) );
  INVX1 U1040 ( .A(dout16_reg[90]), .Y(n437) );
  INVX1 U1041 ( .A(dout16_reg[74]), .Y(n436) );
  INVX1 U1042 ( .A(dout16_reg[58]), .Y(n435) );
  INVX1 U1043 ( .A(dout16_reg[42]), .Y(n434) );
  INVX1 U1044 ( .A(dout16_reg[26]), .Y(n433) );
  INVX1 U1045 ( .A(dout16_reg[10]), .Y(n432) );
  INVX1 U1046 ( .A(dout16_reg[123]), .Y(n423) );
  INVX1 U1047 ( .A(dout16_reg[107]), .Y(n422) );
  INVX1 U1048 ( .A(dout16_reg[91]), .Y(n421) );
  INVX1 U1049 ( .A(dout16_reg[75]), .Y(n420) );
  INVX1 U1050 ( .A(dout16_reg[59]), .Y(n419) );
  INVX1 U1051 ( .A(dout16_reg[43]), .Y(n418) );
  INVX1 U1052 ( .A(dout16_reg[27]), .Y(n417) );
  INVX1 U1053 ( .A(dout16_reg[11]), .Y(n416) );
  INVX1 U1054 ( .A(dout16_reg[124]), .Y(n407) );
  INVX1 U1055 ( .A(dout16_reg[108]), .Y(n406) );
  INVX1 U1056 ( .A(dout16_reg[92]), .Y(n405) );
  INVX1 U1057 ( .A(dout16_reg[76]), .Y(n404) );
  INVX1 U1058 ( .A(dout16_reg[60]), .Y(n403) );
  INVX1 U1059 ( .A(dout16_reg[44]), .Y(n402) );
  INVX1 U1060 ( .A(dout16_reg[28]), .Y(n401) );
  INVX1 U1061 ( .A(dout16_reg[12]), .Y(n400) );
  INVX1 U1062 ( .A(dout16_reg[125]), .Y(n391) );
  INVX1 U1063 ( .A(dout16_reg[109]), .Y(n390) );
  INVX1 U1064 ( .A(dout16_reg[93]), .Y(n389) );
  INVX1 U1065 ( .A(dout16_reg[77]), .Y(n388) );
  INVX1 U1066 ( .A(dout16_reg[61]), .Y(n387) );
  INVX1 U1067 ( .A(dout16_reg[45]), .Y(n386) );
  INVX1 U1068 ( .A(dout16_reg[29]), .Y(n385) );
  INVX1 U1069 ( .A(dout16_reg[13]), .Y(n384) );
  INVX1 U1070 ( .A(dout16_reg[126]), .Y(n375) );
  INVX1 U1071 ( .A(dout16_reg[110]), .Y(n374) );
  INVX1 U1072 ( .A(dout16_reg[94]), .Y(n373) );
  INVX1 U1073 ( .A(dout16_reg[78]), .Y(n372) );
  INVX1 U1074 ( .A(dout16_reg[62]), .Y(n371) );
  INVX1 U1075 ( .A(dout16_reg[46]), .Y(n370) );
  INVX1 U1076 ( .A(dout16_reg[30]), .Y(n369) );
  INVX1 U1077 ( .A(dout16_reg[14]), .Y(n368) );
  INVX1 U1078 ( .A(dout16_reg[127]), .Y(n359) );
  INVX1 U1079 ( .A(dout16_reg[111]), .Y(n358) );
  INVX1 U1080 ( .A(dout16_reg[95]), .Y(n357) );
  INVX1 U1081 ( .A(dout16_reg[79]), .Y(n356) );
  INVX1 U1082 ( .A(dout16_reg[63]), .Y(n355) );
  INVX1 U1083 ( .A(dout16_reg[47]), .Y(n354) );
  INVX1 U1084 ( .A(dout16_reg[31]), .Y(n353) );
  INVX1 U1085 ( .A(dout16_reg[15]), .Y(n352) );
  INVX1 U1086 ( .A(count[2]), .Y(n350) );
  ADDHXL U1087 ( .A(count[2]), .B(r71_carry[2]), .CO(r71_carry[3]), .S(N303)
         );
  ADDHXL U1088 ( .A(count[1]), .B(count[0]), .CO(r71_carry[2]), .S(N302) );
  ADDHXL U1089 ( .A(count[3]), .B(r71_carry[3]), .CO(r71_carry[4]), .S(N304)
         );
  INVX1 U1090 ( .A(dout16_reg[239]), .Y(n366) );
  INVX1 U1091 ( .A(dout8_reg[111]), .Y(n614) );
  INVX1 U1092 ( .A(dout4_reg[47]), .Y(n1203) );
  INVX1 U1093 ( .A(dout16_reg[224]), .Y(n606) );
  INVX1 U1094 ( .A(dout16_reg[208]), .Y(n605) );
  INVX1 U1095 ( .A(dout16_reg[192]), .Y(n604) );
  INVX1 U1096 ( .A(dout16_reg[225]), .Y(n590) );
  INVX1 U1097 ( .A(dout16_reg[209]), .Y(n589) );
  INVX1 U1098 ( .A(dout16_reg[193]), .Y(n588) );
  INVX1 U1099 ( .A(dout16_reg[226]), .Y(n574) );
  INVX1 U1100 ( .A(dout16_reg[210]), .Y(n573) );
  INVX1 U1101 ( .A(dout16_reg[194]), .Y(n572) );
  INVX1 U1102 ( .A(dout16_reg[227]), .Y(n558) );
  INVX1 U1103 ( .A(dout16_reg[211]), .Y(n557) );
  INVX1 U1104 ( .A(dout16_reg[195]), .Y(n556) );
  INVX1 U1105 ( .A(dout16_reg[228]), .Y(n542) );
  INVX1 U1106 ( .A(dout16_reg[212]), .Y(n541) );
  INVX1 U1107 ( .A(dout16_reg[196]), .Y(n540) );
  INVX1 U1108 ( .A(dout16_reg[229]), .Y(n526) );
  INVX1 U1109 ( .A(dout16_reg[213]), .Y(n525) );
  INVX1 U1110 ( .A(dout16_reg[197]), .Y(n524) );
  INVX1 U1111 ( .A(dout16_reg[230]), .Y(n510) );
  INVX1 U1112 ( .A(dout16_reg[214]), .Y(n509) );
  INVX1 U1113 ( .A(dout16_reg[198]), .Y(n508) );
  INVX1 U1114 ( .A(dout16_reg[231]), .Y(n494) );
  INVX1 U1115 ( .A(dout16_reg[215]), .Y(n493) );
  INVX1 U1116 ( .A(dout16_reg[199]), .Y(n492) );
  INVX1 U1117 ( .A(dout16_reg[232]), .Y(n478) );
  INVX1 U1118 ( .A(dout16_reg[216]), .Y(n477) );
  INVX1 U1119 ( .A(dout16_reg[200]), .Y(n476) );
  INVX1 U1120 ( .A(dout16_reg[233]), .Y(n462) );
  INVX1 U1121 ( .A(dout16_reg[217]), .Y(n461) );
  INVX1 U1122 ( .A(dout16_reg[201]), .Y(n460) );
  INVX1 U1123 ( .A(dout16_reg[234]), .Y(n446) );
  INVX1 U1124 ( .A(dout16_reg[218]), .Y(n445) );
  INVX1 U1125 ( .A(dout16_reg[202]), .Y(n444) );
  INVX1 U1126 ( .A(dout16_reg[235]), .Y(n430) );
  INVX1 U1127 ( .A(dout16_reg[219]), .Y(n429) );
  INVX1 U1128 ( .A(dout16_reg[203]), .Y(n428) );
  INVX1 U1129 ( .A(dout16_reg[236]), .Y(n414) );
  INVX1 U1130 ( .A(dout16_reg[220]), .Y(n413) );
  INVX1 U1131 ( .A(dout16_reg[204]), .Y(n412) );
  INVX1 U1132 ( .A(dout16_reg[237]), .Y(n398) );
  INVX1 U1133 ( .A(dout16_reg[221]), .Y(n397) );
  INVX1 U1134 ( .A(dout16_reg[205]), .Y(n396) );
  INVX1 U1135 ( .A(dout16_reg[238]), .Y(n382) );
  INVX1 U1136 ( .A(dout16_reg[222]), .Y(n381) );
  INVX1 U1137 ( .A(dout16_reg[206]), .Y(n380) );
  INVX1 U1138 ( .A(dout16_reg[223]), .Y(n365) );
  INVX1 U1139 ( .A(dout16_reg[207]), .Y(n364) );
  INVX1 U1140 ( .A(dout8_reg[96]), .Y(n1199) );
  INVX1 U1141 ( .A(dout8_reg[80]), .Y(n739) );
  INVX1 U1142 ( .A(dout8_reg[64]), .Y(n738) );
  INVX1 U1143 ( .A(dout8_reg[97]), .Y(n726) );
  INVX1 U1144 ( .A(dout8_reg[81]), .Y(n725) );
  INVX1 U1145 ( .A(dout8_reg[65]), .Y(n724) );
  INVX1 U1146 ( .A(dout8_reg[98]), .Y(n718) );
  INVX1 U1147 ( .A(dout8_reg[82]), .Y(n717) );
  INVX1 U1148 ( .A(dout8_reg[66]), .Y(n716) );
  INVX1 U1149 ( .A(dout8_reg[99]), .Y(n710) );
  INVX1 U1150 ( .A(dout8_reg[83]), .Y(n709) );
  INVX1 U1151 ( .A(dout8_reg[67]), .Y(n708) );
  INVX1 U1152 ( .A(dout8_reg[100]), .Y(n702) );
  INVX1 U1153 ( .A(dout8_reg[84]), .Y(n701) );
  INVX1 U1154 ( .A(dout8_reg[68]), .Y(n700) );
  INVX1 U1155 ( .A(dout8_reg[101]), .Y(n694) );
  INVX1 U1156 ( .A(dout8_reg[85]), .Y(n693) );
  INVX1 U1157 ( .A(dout8_reg[69]), .Y(n692) );
  INVX1 U1158 ( .A(dout8_reg[102]), .Y(n686) );
  INVX1 U1159 ( .A(dout8_reg[86]), .Y(n685) );
  INVX1 U1160 ( .A(dout8_reg[70]), .Y(n684) );
  INVX1 U1161 ( .A(dout8_reg[103]), .Y(n678) );
  INVX1 U1162 ( .A(dout8_reg[87]), .Y(n677) );
  INVX1 U1163 ( .A(dout8_reg[71]), .Y(n676) );
  INVX1 U1164 ( .A(dout8_reg[104]), .Y(n670) );
  INVX1 U1165 ( .A(dout8_reg[88]), .Y(n669) );
  INVX1 U1166 ( .A(dout8_reg[72]), .Y(n668) );
  INVX1 U1167 ( .A(dout8_reg[105]), .Y(n662) );
  INVX1 U1168 ( .A(dout8_reg[89]), .Y(n661) );
  INVX1 U1169 ( .A(dout8_reg[73]), .Y(n660) );
  INVX1 U1170 ( .A(dout8_reg[106]), .Y(n654) );
  INVX1 U1171 ( .A(dout8_reg[90]), .Y(n653) );
  INVX1 U1172 ( .A(dout8_reg[74]), .Y(n652) );
  INVX1 U1173 ( .A(dout8_reg[107]), .Y(n646) );
  INVX1 U1174 ( .A(dout8_reg[91]), .Y(n645) );
  INVX1 U1175 ( .A(dout8_reg[75]), .Y(n644) );
  INVX1 U1176 ( .A(dout8_reg[108]), .Y(n638) );
  INVX1 U1177 ( .A(dout8_reg[92]), .Y(n637) );
  INVX1 U1178 ( .A(dout8_reg[76]), .Y(n636) );
  INVX1 U1179 ( .A(dout8_reg[109]), .Y(n630) );
  INVX1 U1180 ( .A(dout8_reg[93]), .Y(n629) );
  INVX1 U1181 ( .A(dout8_reg[77]), .Y(n628) );
  INVX1 U1182 ( .A(dout8_reg[110]), .Y(n622) );
  INVX1 U1183 ( .A(dout8_reg[94]), .Y(n621) );
  INVX1 U1184 ( .A(dout8_reg[78]), .Y(n620) );
  INVX1 U1185 ( .A(dout8_reg[95]), .Y(n613) );
  INVX1 U1186 ( .A(dout8_reg[79]), .Y(n612) );
  INVX1 U1187 ( .A(dout4_reg[32]), .Y(n1263) );
  INVX1 U1188 ( .A(dout4_reg[16]), .Y(n1262) );
  INVX1 U1189 ( .A(dout4_reg[0]), .Y(n1261) );
  INVX1 U1190 ( .A(dout4_reg[33]), .Y(n1259) );
  INVX1 U1191 ( .A(dout4_reg[17]), .Y(n1258) );
  INVX1 U1192 ( .A(dout4_reg[1]), .Y(n1257) );
  INVX1 U1193 ( .A(dout4_reg[34]), .Y(n1255) );
  INVX1 U1194 ( .A(dout4_reg[18]), .Y(n1254) );
  INVX1 U1195 ( .A(dout4_reg[2]), .Y(n1253) );
  INVX1 U1196 ( .A(dout4_reg[35]), .Y(n1251) );
  INVX1 U1197 ( .A(dout4_reg[19]), .Y(n1250) );
  INVX1 U1198 ( .A(dout4_reg[3]), .Y(n1249) );
  INVX1 U1199 ( .A(dout4_reg[36]), .Y(n1247) );
  INVX1 U1200 ( .A(dout4_reg[20]), .Y(n1246) );
  INVX1 U1201 ( .A(dout4_reg[4]), .Y(n1245) );
  INVX1 U1202 ( .A(dout4_reg[37]), .Y(n1243) );
  INVX1 U1203 ( .A(dout4_reg[21]), .Y(n1242) );
  INVX1 U1204 ( .A(dout4_reg[5]), .Y(n1241) );
  INVX1 U1205 ( .A(dout4_reg[38]), .Y(n1239) );
  INVX1 U1206 ( .A(dout4_reg[22]), .Y(n1238) );
  INVX1 U1207 ( .A(dout4_reg[6]), .Y(n1237) );
  INVX1 U1208 ( .A(dout4_reg[39]), .Y(n1235) );
  INVX1 U1209 ( .A(dout4_reg[23]), .Y(n1234) );
  INVX1 U1210 ( .A(dout4_reg[7]), .Y(n1233) );
  INVX1 U1211 ( .A(dout4_reg[40]), .Y(n1231) );
  INVX1 U1212 ( .A(dout4_reg[24]), .Y(n1230) );
  INVX1 U1213 ( .A(dout4_reg[8]), .Y(n1229) );
  INVX1 U1214 ( .A(dout4_reg[41]), .Y(n1227) );
  INVX1 U1215 ( .A(dout4_reg[25]), .Y(n1226) );
  INVX1 U1216 ( .A(dout4_reg[9]), .Y(n1225) );
  INVX1 U1217 ( .A(dout4_reg[42]), .Y(n1223) );
  INVX1 U1218 ( .A(dout4_reg[26]), .Y(n1222) );
  INVX1 U1219 ( .A(dout4_reg[10]), .Y(n1221) );
  INVX1 U1220 ( .A(dout4_reg[43]), .Y(n1219) );
  INVX1 U1221 ( .A(dout4_reg[27]), .Y(n1218) );
  INVX1 U1222 ( .A(dout4_reg[11]), .Y(n1217) );
  INVX1 U1223 ( .A(dout4_reg[44]), .Y(n1215) );
  INVX1 U1224 ( .A(dout4_reg[28]), .Y(n1214) );
  INVX1 U1225 ( .A(dout4_reg[12]), .Y(n1213) );
  INVX1 U1226 ( .A(dout4_reg[45]), .Y(n1211) );
  INVX1 U1227 ( .A(dout4_reg[29]), .Y(n1210) );
  INVX1 U1228 ( .A(dout4_reg[13]), .Y(n1209) );
  INVX1 U1229 ( .A(dout4_reg[46]), .Y(n1207) );
  INVX1 U1230 ( .A(dout4_reg[30]), .Y(n1206) );
  INVX1 U1231 ( .A(dout4_reg[14]), .Y(n1205) );
  INVX1 U1232 ( .A(dout4_reg[31]), .Y(n1202) );
  INVX1 U1233 ( .A(dout4_reg[15]), .Y(n1201) );
  INVX1 U1234 ( .A(dout16_reg[240]), .Y(n607) );
  INVX1 U1235 ( .A(dout16_reg[241]), .Y(n591) );
  INVX1 U1236 ( .A(dout16_reg[242]), .Y(n575) );
  INVX1 U1237 ( .A(dout16_reg[243]), .Y(n559) );
  INVX1 U1238 ( .A(dout16_reg[244]), .Y(n543) );
  INVX1 U1239 ( .A(dout16_reg[245]), .Y(n527) );
  INVX1 U1240 ( .A(dout16_reg[246]), .Y(n511) );
  INVX1 U1241 ( .A(dout16_reg[247]), .Y(n495) );
  INVX1 U1242 ( .A(dout16_reg[248]), .Y(n479) );
  INVX1 U1243 ( .A(dout16_reg[249]), .Y(n463) );
  INVX1 U1244 ( .A(dout16_reg[250]), .Y(n447) );
  INVX1 U1245 ( .A(dout16_reg[251]), .Y(n431) );
  INVX1 U1246 ( .A(dout16_reg[252]), .Y(n415) );
  INVX1 U1247 ( .A(dout16_reg[253]), .Y(n399) );
  INVX1 U1248 ( .A(dout16_reg[254]), .Y(n383) );
  INVX1 U1249 ( .A(dout16_reg[255]), .Y(n367) );
  INVX1 U1250 ( .A(dout8_reg[112]), .Y(n1200) );
  INVX1 U1251 ( .A(dout8_reg[113]), .Y(n727) );
  INVX1 U1252 ( .A(dout8_reg[114]), .Y(n719) );
  INVX1 U1253 ( .A(dout8_reg[115]), .Y(n711) );
  INVX1 U1254 ( .A(dout8_reg[116]), .Y(n703) );
  INVX1 U1255 ( .A(dout8_reg[117]), .Y(n695) );
  INVX1 U1256 ( .A(dout8_reg[118]), .Y(n687) );
  INVX1 U1257 ( .A(dout8_reg[119]), .Y(n679) );
  INVX1 U1258 ( .A(dout8_reg[120]), .Y(n671) );
  INVX1 U1259 ( .A(dout8_reg[121]), .Y(n663) );
  INVX1 U1260 ( .A(dout8_reg[122]), .Y(n655) );
  INVX1 U1261 ( .A(dout8_reg[123]), .Y(n647) );
  INVX1 U1262 ( .A(dout8_reg[124]), .Y(n639) );
  INVX1 U1263 ( .A(dout8_reg[125]), .Y(n631) );
  INVX1 U1264 ( .A(dout8_reg[126]), .Y(n623) );
  INVX1 U1265 ( .A(dout8_reg[127]), .Y(n615) );
  INVX1 U1266 ( .A(dout4_reg[48]), .Y(n1264) );
  INVX1 U1267 ( .A(dout4_reg[49]), .Y(n1260) );
  INVX1 U1268 ( .A(dout4_reg[50]), .Y(n1256) );
  INVX1 U1269 ( .A(dout4_reg[51]), .Y(n1252) );
  INVX1 U1270 ( .A(dout4_reg[52]), .Y(n1248) );
  INVX1 U1271 ( .A(dout4_reg[53]), .Y(n1244) );
  INVX1 U1272 ( .A(dout4_reg[54]), .Y(n1240) );
  INVX1 U1273 ( .A(dout4_reg[55]), .Y(n1236) );
  INVX1 U1274 ( .A(dout4_reg[56]), .Y(n1232) );
  INVX1 U1275 ( .A(dout4_reg[57]), .Y(n1228) );
  INVX1 U1276 ( .A(dout4_reg[58]), .Y(n1224) );
  INVX1 U1277 ( .A(dout4_reg[59]), .Y(n1220) );
  INVX1 U1278 ( .A(dout4_reg[60]), .Y(n1216) );
  INVX1 U1279 ( .A(dout4_reg[61]), .Y(n1212) );
  INVX1 U1280 ( .A(dout4_reg[62]), .Y(n1208) );
  INVX1 U1281 ( .A(dout4_reg[63]), .Y(n1204) );
  NAND2X1 U1282 ( .A(mode_reg[1]), .B(n349), .Y(n1728) );
  NAND2X1 U1283 ( .A(mode_reg[0]), .B(n348), .Y(n1726) );
endmodule


module even_odd_1 ( clk, rstn, mode, start, din, dout, even_odd_ready, 
        mode_out );
  input [1:0] mode;
  input [255:0] din;
  output [255:0] dout;
  output [1:0] mode_out;
  input clk, rstn, start;
  output even_odd_ready;
  wire   N275, n2, n19, n20, n149, n150, n151, n152, n154, n155, n157, n158,
         n160, n161, n163, n164, n166, n167, n169, n170, n172, n173, n175,
         n176, n178, n179, n181, n182, n184, n185, n187, n188, n190, n191,
         n193, n194, n196, n197, n199, n201, n203, n205, n207, n209, n211,
         n213, n215, n217, n219, n221, n223, n225, n227, n229, n231, n232,
         n234, n235, n237, n238, n240, n241, n243, n244, n246, n247, n249,
         n250, n252, n253, n255, n256, n258, n259, n261, n262, n264, n265,
         n267, n268, n270, n271, n273, n274, n276, n277, n295, n297, n299,
         n301, n303, n305, n307, n309, n311, n313, n315, n317, n319, n321,
         n323, n325, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170;

  DFFRHQX1 dout_reg_15_ ( .D(n892), .CK(clk), .RN(rstn), .Q(dout[15]) );
  DFFRHQX1 dout_reg_14_ ( .D(n893), .CK(clk), .RN(rstn), .Q(dout[14]) );
  DFFRHQX1 dout_reg_13_ ( .D(n894), .CK(clk), .RN(rstn), .Q(dout[13]) );
  DFFRHQX1 dout_reg_12_ ( .D(n895), .CK(clk), .RN(rstn), .Q(dout[12]) );
  DFFRHQX1 dout_reg_11_ ( .D(n896), .CK(clk), .RN(rstn), .Q(dout[11]) );
  DFFRHQX1 dout_reg_10_ ( .D(n897), .CK(clk), .RN(rstn), .Q(dout[10]) );
  DFFRHQX1 dout_reg_9_ ( .D(n898), .CK(clk), .RN(rstn), .Q(dout[9]) );
  DFFRHQX1 dout_reg_8_ ( .D(n899), .CK(clk), .RN(rstn), .Q(dout[8]) );
  DFFRHQX1 dout_reg_7_ ( .D(n900), .CK(clk), .RN(rstn), .Q(dout[7]) );
  DFFRHQX1 dout_reg_6_ ( .D(n901), .CK(clk), .RN(rstn), .Q(dout[6]) );
  DFFRHQX1 dout_reg_5_ ( .D(n902), .CK(clk), .RN(rstn), .Q(dout[5]) );
  DFFRHQX1 dout_reg_4_ ( .D(n903), .CK(clk), .RN(rstn), .Q(dout[4]) );
  DFFRHQX1 dout_reg_3_ ( .D(n904), .CK(clk), .RN(rstn), .Q(dout[3]) );
  DFFRHQX1 dout_reg_2_ ( .D(n905), .CK(clk), .RN(rstn), .Q(dout[2]) );
  DFFRHQX1 dout_reg_1_ ( .D(n906), .CK(clk), .RN(rstn), .Q(dout[1]) );
  DFFRHQX1 dout_reg_0_ ( .D(n907), .CK(clk), .RN(rstn), .Q(dout[0]) );
  DFFRHQX1 mode_out_reg_1_ ( .D(n650), .CK(clk), .RN(rstn), .Q(mode_out[1]) );
  DFFRHQX1 mode_out_reg_0_ ( .D(n651), .CK(clk), .RN(rstn), .Q(mode_out[0]) );
  DFFRHQX1 dout_reg_255_ ( .D(n652), .CK(clk), .RN(rstn), .Q(dout[255]) );
  DFFRHQX1 dout_reg_254_ ( .D(n653), .CK(clk), .RN(rstn), .Q(dout[254]) );
  DFFRHQX1 dout_reg_253_ ( .D(n654), .CK(clk), .RN(rstn), .Q(dout[253]) );
  DFFRHQX1 dout_reg_252_ ( .D(n655), .CK(clk), .RN(rstn), .Q(dout[252]) );
  DFFRHQX1 dout_reg_251_ ( .D(n656), .CK(clk), .RN(rstn), .Q(dout[251]) );
  DFFRHQX1 dout_reg_250_ ( .D(n657), .CK(clk), .RN(rstn), .Q(dout[250]) );
  DFFRHQX1 dout_reg_249_ ( .D(n658), .CK(clk), .RN(rstn), .Q(dout[249]) );
  DFFRHQX1 dout_reg_248_ ( .D(n659), .CK(clk), .RN(rstn), .Q(dout[248]) );
  DFFRHQX1 dout_reg_247_ ( .D(n660), .CK(clk), .RN(rstn), .Q(dout[247]) );
  DFFRHQX1 dout_reg_246_ ( .D(n661), .CK(clk), .RN(rstn), .Q(dout[246]) );
  DFFRHQX1 dout_reg_245_ ( .D(n662), .CK(clk), .RN(rstn), .Q(dout[245]) );
  DFFRHQX1 dout_reg_244_ ( .D(n663), .CK(clk), .RN(rstn), .Q(dout[244]) );
  DFFRHQX1 dout_reg_243_ ( .D(n664), .CK(clk), .RN(rstn), .Q(dout[243]) );
  DFFRHQX1 dout_reg_242_ ( .D(n665), .CK(clk), .RN(rstn), .Q(dout[242]) );
  DFFRHQX1 dout_reg_241_ ( .D(n666), .CK(clk), .RN(rstn), .Q(dout[241]) );
  DFFRHQX1 dout_reg_240_ ( .D(n667), .CK(clk), .RN(rstn), .Q(dout[240]) );
  DFFRHQX1 dout_reg_127_ ( .D(n780), .CK(clk), .RN(rstn), .Q(dout[127]) );
  DFFRHQX1 dout_reg_126_ ( .D(n781), .CK(clk), .RN(rstn), .Q(dout[126]) );
  DFFRHQX1 dout_reg_125_ ( .D(n782), .CK(clk), .RN(rstn), .Q(dout[125]) );
  DFFRHQX1 dout_reg_124_ ( .D(n783), .CK(clk), .RN(rstn), .Q(dout[124]) );
  DFFRHQX1 dout_reg_123_ ( .D(n784), .CK(clk), .RN(rstn), .Q(dout[123]) );
  DFFRHQX1 dout_reg_122_ ( .D(n785), .CK(clk), .RN(rstn), .Q(dout[122]) );
  DFFRHQX1 dout_reg_121_ ( .D(n786), .CK(clk), .RN(rstn), .Q(dout[121]) );
  DFFRHQX1 dout_reg_120_ ( .D(n787), .CK(clk), .RN(rstn), .Q(dout[120]) );
  DFFRHQX1 dout_reg_119_ ( .D(n788), .CK(clk), .RN(rstn), .Q(dout[119]) );
  DFFRHQX1 dout_reg_118_ ( .D(n789), .CK(clk), .RN(rstn), .Q(dout[118]) );
  DFFRHQX1 dout_reg_117_ ( .D(n790), .CK(clk), .RN(rstn), .Q(dout[117]) );
  DFFRHQX1 dout_reg_116_ ( .D(n791), .CK(clk), .RN(rstn), .Q(dout[116]) );
  DFFRHQX1 dout_reg_115_ ( .D(n792), .CK(clk), .RN(rstn), .Q(dout[115]) );
  DFFRHQX1 dout_reg_114_ ( .D(n793), .CK(clk), .RN(rstn), .Q(dout[114]) );
  DFFRHQX1 dout_reg_113_ ( .D(n794), .CK(clk), .RN(rstn), .Q(dout[113]) );
  DFFRHQX1 dout_reg_112_ ( .D(n795), .CK(clk), .RN(rstn), .Q(dout[112]) );
  DFFRHQX1 dout_reg_111_ ( .D(n796), .CK(clk), .RN(rstn), .Q(dout[111]) );
  DFFRHQX1 dout_reg_110_ ( .D(n797), .CK(clk), .RN(rstn), .Q(dout[110]) );
  DFFRHQX1 dout_reg_109_ ( .D(n798), .CK(clk), .RN(rstn), .Q(dout[109]) );
  DFFRHQX1 dout_reg_108_ ( .D(n799), .CK(clk), .RN(rstn), .Q(dout[108]) );
  DFFRHQX1 dout_reg_107_ ( .D(n800), .CK(clk), .RN(rstn), .Q(dout[107]) );
  DFFRHQX1 dout_reg_106_ ( .D(n801), .CK(clk), .RN(rstn), .Q(dout[106]) );
  DFFRHQX1 dout_reg_105_ ( .D(n802), .CK(clk), .RN(rstn), .Q(dout[105]) );
  DFFRHQX1 dout_reg_104_ ( .D(n803), .CK(clk), .RN(rstn), .Q(dout[104]) );
  DFFRHQX1 dout_reg_103_ ( .D(n804), .CK(clk), .RN(rstn), .Q(dout[103]) );
  DFFRHQX1 dout_reg_102_ ( .D(n805), .CK(clk), .RN(rstn), .Q(dout[102]) );
  DFFRHQX1 dout_reg_101_ ( .D(n806), .CK(clk), .RN(rstn), .Q(dout[101]) );
  DFFRHQX1 dout_reg_100_ ( .D(n807), .CK(clk), .RN(rstn), .Q(dout[100]) );
  DFFRHQX1 dout_reg_99_ ( .D(n808), .CK(clk), .RN(rstn), .Q(dout[99]) );
  DFFRHQX1 dout_reg_98_ ( .D(n809), .CK(clk), .RN(rstn), .Q(dout[98]) );
  DFFRHQX1 dout_reg_97_ ( .D(n810), .CK(clk), .RN(rstn), .Q(dout[97]) );
  DFFRHQX1 dout_reg_96_ ( .D(n811), .CK(clk), .RN(rstn), .Q(dout[96]) );
  DFFRHQX1 dout_reg_95_ ( .D(n812), .CK(clk), .RN(rstn), .Q(dout[95]) );
  DFFRHQX1 dout_reg_94_ ( .D(n813), .CK(clk), .RN(rstn), .Q(dout[94]) );
  DFFRHQX1 dout_reg_93_ ( .D(n814), .CK(clk), .RN(rstn), .Q(dout[93]) );
  DFFRHQX1 dout_reg_92_ ( .D(n815), .CK(clk), .RN(rstn), .Q(dout[92]) );
  DFFRHQX1 dout_reg_91_ ( .D(n816), .CK(clk), .RN(rstn), .Q(dout[91]) );
  DFFRHQX1 dout_reg_90_ ( .D(n817), .CK(clk), .RN(rstn), .Q(dout[90]) );
  DFFRHQX1 dout_reg_89_ ( .D(n818), .CK(clk), .RN(rstn), .Q(dout[89]) );
  DFFRHQX1 dout_reg_88_ ( .D(n819), .CK(clk), .RN(rstn), .Q(dout[88]) );
  DFFRHQX1 dout_reg_87_ ( .D(n820), .CK(clk), .RN(rstn), .Q(dout[87]) );
  DFFRHQX1 dout_reg_86_ ( .D(n821), .CK(clk), .RN(rstn), .Q(dout[86]) );
  DFFRHQX1 dout_reg_85_ ( .D(n822), .CK(clk), .RN(rstn), .Q(dout[85]) );
  DFFRHQX1 dout_reg_84_ ( .D(n823), .CK(clk), .RN(rstn), .Q(dout[84]) );
  DFFRHQX1 dout_reg_83_ ( .D(n824), .CK(clk), .RN(rstn), .Q(dout[83]) );
  DFFRHQX1 dout_reg_82_ ( .D(n825), .CK(clk), .RN(rstn), .Q(dout[82]) );
  DFFRHQX1 dout_reg_81_ ( .D(n826), .CK(clk), .RN(rstn), .Q(dout[81]) );
  DFFRHQX1 dout_reg_80_ ( .D(n827), .CK(clk), .RN(rstn), .Q(dout[80]) );
  DFFRHQX1 dout_reg_79_ ( .D(n828), .CK(clk), .RN(rstn), .Q(dout[79]) );
  DFFRHQX1 dout_reg_78_ ( .D(n829), .CK(clk), .RN(rstn), .Q(dout[78]) );
  DFFRHQX1 dout_reg_77_ ( .D(n830), .CK(clk), .RN(rstn), .Q(dout[77]) );
  DFFRHQX1 dout_reg_76_ ( .D(n831), .CK(clk), .RN(rstn), .Q(dout[76]) );
  DFFRHQX1 dout_reg_75_ ( .D(n832), .CK(clk), .RN(rstn), .Q(dout[75]) );
  DFFRHQX1 dout_reg_74_ ( .D(n833), .CK(clk), .RN(rstn), .Q(dout[74]) );
  DFFRHQX1 dout_reg_73_ ( .D(n834), .CK(clk), .RN(rstn), .Q(dout[73]) );
  DFFRHQX1 dout_reg_72_ ( .D(n835), .CK(clk), .RN(rstn), .Q(dout[72]) );
  DFFRHQX1 dout_reg_71_ ( .D(n836), .CK(clk), .RN(rstn), .Q(dout[71]) );
  DFFRHQX1 dout_reg_70_ ( .D(n837), .CK(clk), .RN(rstn), .Q(dout[70]) );
  DFFRHQX1 dout_reg_69_ ( .D(n838), .CK(clk), .RN(rstn), .Q(dout[69]) );
  DFFRHQX1 dout_reg_68_ ( .D(n839), .CK(clk), .RN(rstn), .Q(dout[68]) );
  DFFRHQX1 dout_reg_67_ ( .D(n840), .CK(clk), .RN(rstn), .Q(dout[67]) );
  DFFRHQX1 dout_reg_66_ ( .D(n841), .CK(clk), .RN(rstn), .Q(dout[66]) );
  DFFRHQX1 dout_reg_65_ ( .D(n842), .CK(clk), .RN(rstn), .Q(dout[65]) );
  DFFRHQX1 dout_reg_64_ ( .D(n843), .CK(clk), .RN(rstn), .Q(dout[64]) );
  DFFRHQX1 dout_reg_63_ ( .D(n844), .CK(clk), .RN(rstn), .Q(dout[63]) );
  DFFRHQX1 dout_reg_62_ ( .D(n845), .CK(clk), .RN(rstn), .Q(dout[62]) );
  DFFRHQX1 dout_reg_61_ ( .D(n846), .CK(clk), .RN(rstn), .Q(dout[61]) );
  DFFRHQX1 dout_reg_60_ ( .D(n847), .CK(clk), .RN(rstn), .Q(dout[60]) );
  DFFRHQX1 dout_reg_59_ ( .D(n848), .CK(clk), .RN(rstn), .Q(dout[59]) );
  DFFRHQX1 dout_reg_58_ ( .D(n849), .CK(clk), .RN(rstn), .Q(dout[58]) );
  DFFRHQX1 dout_reg_57_ ( .D(n850), .CK(clk), .RN(rstn), .Q(dout[57]) );
  DFFRHQX1 dout_reg_56_ ( .D(n851), .CK(clk), .RN(rstn), .Q(dout[56]) );
  DFFRHQX1 dout_reg_55_ ( .D(n852), .CK(clk), .RN(rstn), .Q(dout[55]) );
  DFFRHQX1 dout_reg_54_ ( .D(n853), .CK(clk), .RN(rstn), .Q(dout[54]) );
  DFFRHQX1 dout_reg_53_ ( .D(n854), .CK(clk), .RN(rstn), .Q(dout[53]) );
  DFFRHQX1 dout_reg_52_ ( .D(n855), .CK(clk), .RN(rstn), .Q(dout[52]) );
  DFFRHQX1 dout_reg_51_ ( .D(n856), .CK(clk), .RN(rstn), .Q(dout[51]) );
  DFFRHQX1 dout_reg_50_ ( .D(n857), .CK(clk), .RN(rstn), .Q(dout[50]) );
  DFFRHQX1 dout_reg_49_ ( .D(n858), .CK(clk), .RN(rstn), .Q(dout[49]) );
  DFFRHQX1 dout_reg_48_ ( .D(n859), .CK(clk), .RN(rstn), .Q(dout[48]) );
  DFFRHQX1 dout_reg_47_ ( .D(n860), .CK(clk), .RN(rstn), .Q(dout[47]) );
  DFFRHQX1 dout_reg_46_ ( .D(n861), .CK(clk), .RN(rstn), .Q(dout[46]) );
  DFFRHQX1 dout_reg_45_ ( .D(n862), .CK(clk), .RN(rstn), .Q(dout[45]) );
  DFFRHQX1 dout_reg_44_ ( .D(n863), .CK(clk), .RN(rstn), .Q(dout[44]) );
  DFFRHQX1 dout_reg_43_ ( .D(n864), .CK(clk), .RN(rstn), .Q(dout[43]) );
  DFFRHQX1 dout_reg_42_ ( .D(n865), .CK(clk), .RN(rstn), .Q(dout[42]) );
  DFFRHQX1 dout_reg_41_ ( .D(n866), .CK(clk), .RN(rstn), .Q(dout[41]) );
  DFFRHQX1 dout_reg_40_ ( .D(n867), .CK(clk), .RN(rstn), .Q(dout[40]) );
  DFFRHQX1 dout_reg_39_ ( .D(n868), .CK(clk), .RN(rstn), .Q(dout[39]) );
  DFFRHQX1 dout_reg_38_ ( .D(n869), .CK(clk), .RN(rstn), .Q(dout[38]) );
  DFFRHQX1 dout_reg_37_ ( .D(n870), .CK(clk), .RN(rstn), .Q(dout[37]) );
  DFFRHQX1 dout_reg_36_ ( .D(n871), .CK(clk), .RN(rstn), .Q(dout[36]) );
  DFFRHQX1 dout_reg_35_ ( .D(n872), .CK(clk), .RN(rstn), .Q(dout[35]) );
  DFFRHQX1 dout_reg_34_ ( .D(n873), .CK(clk), .RN(rstn), .Q(dout[34]) );
  DFFRHQX1 dout_reg_33_ ( .D(n874), .CK(clk), .RN(rstn), .Q(dout[33]) );
  DFFRHQX1 dout_reg_32_ ( .D(n875), .CK(clk), .RN(rstn), .Q(dout[32]) );
  DFFRHQX1 dout_reg_31_ ( .D(n876), .CK(clk), .RN(rstn), .Q(dout[31]) );
  DFFRHQX1 dout_reg_30_ ( .D(n877), .CK(clk), .RN(rstn), .Q(dout[30]) );
  DFFRHQX1 dout_reg_29_ ( .D(n878), .CK(clk), .RN(rstn), .Q(dout[29]) );
  DFFRHQX1 dout_reg_28_ ( .D(n879), .CK(clk), .RN(rstn), .Q(dout[28]) );
  DFFRHQX1 dout_reg_27_ ( .D(n880), .CK(clk), .RN(rstn), .Q(dout[27]) );
  DFFRHQX1 dout_reg_26_ ( .D(n881), .CK(clk), .RN(rstn), .Q(dout[26]) );
  DFFRHQX1 dout_reg_25_ ( .D(n882), .CK(clk), .RN(rstn), .Q(dout[25]) );
  DFFRHQX1 dout_reg_24_ ( .D(n883), .CK(clk), .RN(rstn), .Q(dout[24]) );
  DFFRHQX1 dout_reg_23_ ( .D(n884), .CK(clk), .RN(rstn), .Q(dout[23]) );
  DFFRHQX1 dout_reg_22_ ( .D(n885), .CK(clk), .RN(rstn), .Q(dout[22]) );
  DFFRHQX1 dout_reg_21_ ( .D(n886), .CK(clk), .RN(rstn), .Q(dout[21]) );
  DFFRHQX1 dout_reg_20_ ( .D(n887), .CK(clk), .RN(rstn), .Q(dout[20]) );
  DFFRHQX1 dout_reg_19_ ( .D(n888), .CK(clk), .RN(rstn), .Q(dout[19]) );
  DFFRHQX1 dout_reg_18_ ( .D(n889), .CK(clk), .RN(rstn), .Q(dout[18]) );
  DFFRHQX1 dout_reg_17_ ( .D(n890), .CK(clk), .RN(rstn), .Q(dout[17]) );
  DFFRHQX1 dout_reg_16_ ( .D(n891), .CK(clk), .RN(rstn), .Q(dout[16]) );
  DFFRHQX1 dout_reg_223_ ( .D(n684), .CK(clk), .RN(rstn), .Q(dout[223]) );
  DFFRHQX1 dout_reg_222_ ( .D(n685), .CK(clk), .RN(rstn), .Q(dout[222]) );
  DFFRHQX1 dout_reg_221_ ( .D(n686), .CK(clk), .RN(rstn), .Q(dout[221]) );
  DFFRHQX1 dout_reg_220_ ( .D(n687), .CK(clk), .RN(rstn), .Q(dout[220]) );
  DFFRHQX1 dout_reg_219_ ( .D(n688), .CK(clk), .RN(rstn), .Q(dout[219]) );
  DFFRHQX1 dout_reg_218_ ( .D(n689), .CK(clk), .RN(rstn), .Q(dout[218]) );
  DFFRHQX1 dout_reg_217_ ( .D(n690), .CK(clk), .RN(rstn), .Q(dout[217]) );
  DFFRHQX1 dout_reg_216_ ( .D(n691), .CK(clk), .RN(rstn), .Q(dout[216]) );
  DFFRHQX1 dout_reg_215_ ( .D(n692), .CK(clk), .RN(rstn), .Q(dout[215]) );
  DFFRHQX1 dout_reg_214_ ( .D(n693), .CK(clk), .RN(rstn), .Q(dout[214]) );
  DFFRHQX1 dout_reg_213_ ( .D(n694), .CK(clk), .RN(rstn), .Q(dout[213]) );
  DFFRHQX1 dout_reg_212_ ( .D(n695), .CK(clk), .RN(rstn), .Q(dout[212]) );
  DFFRHQX1 dout_reg_211_ ( .D(n696), .CK(clk), .RN(rstn), .Q(dout[211]) );
  DFFRHQX1 dout_reg_210_ ( .D(n697), .CK(clk), .RN(rstn), .Q(dout[210]) );
  DFFRHQX1 dout_reg_209_ ( .D(n698), .CK(clk), .RN(rstn), .Q(dout[209]) );
  DFFRHQX1 dout_reg_208_ ( .D(n699), .CK(clk), .RN(rstn), .Q(dout[208]) );
  DFFRHQX1 dout_reg_143_ ( .D(n764), .CK(clk), .RN(rstn), .Q(dout[143]) );
  DFFRHQX1 dout_reg_191_ ( .D(n716), .CK(clk), .RN(rstn), .Q(dout[191]) );
  DFFRHQX1 dout_reg_175_ ( .D(n732), .CK(clk), .RN(rstn), .Q(dout[175]) );
  DFFRHQX1 dout_reg_159_ ( .D(n748), .CK(clk), .RN(rstn), .Q(dout[159]) );
  DFFRHQX1 dout_reg_142_ ( .D(n765), .CK(clk), .RN(rstn), .Q(dout[142]) );
  DFFRHQX1 dout_reg_141_ ( .D(n766), .CK(clk), .RN(rstn), .Q(dout[141]) );
  DFFRHQX1 dout_reg_239_ ( .D(n668), .CK(clk), .RN(rstn), .Q(dout[239]) );
  DFFRHQX1 dout_reg_207_ ( .D(n700), .CK(clk), .RN(rstn), .Q(dout[207]) );
  DFFRHQX1 dout_reg_190_ ( .D(n717), .CK(clk), .RN(rstn), .Q(dout[190]) );
  DFFRHQX1 dout_reg_189_ ( .D(n718), .CK(clk), .RN(rstn), .Q(dout[189]) );
  DFFRHQX1 dout_reg_174_ ( .D(n733), .CK(clk), .RN(rstn), .Q(dout[174]) );
  DFFRHQX1 dout_reg_173_ ( .D(n734), .CK(clk), .RN(rstn), .Q(dout[173]) );
  DFFRHQX1 dout_reg_158_ ( .D(n749), .CK(clk), .RN(rstn), .Q(dout[158]) );
  DFFRHQX1 dout_reg_157_ ( .D(n750), .CK(clk), .RN(rstn), .Q(dout[157]) );
  DFFRHQX1 dout_reg_238_ ( .D(n669), .CK(clk), .RN(rstn), .Q(dout[238]) );
  DFFRHQX1 dout_reg_237_ ( .D(n670), .CK(clk), .RN(rstn), .Q(dout[237]) );
  DFFRHQX1 dout_reg_206_ ( .D(n701), .CK(clk), .RN(rstn), .Q(dout[206]) );
  DFFRHQX1 dout_reg_205_ ( .D(n702), .CK(clk), .RN(rstn), .Q(dout[205]) );
  DFFRHQX1 dout_reg_140_ ( .D(n767), .CK(clk), .RN(rstn), .Q(dout[140]) );
  DFFRHQX1 dout_reg_139_ ( .D(n768), .CK(clk), .RN(rstn), .Q(dout[139]) );
  DFFRHQX1 dout_reg_138_ ( .D(n769), .CK(clk), .RN(rstn), .Q(dout[138]) );
  DFFRHQX1 dout_reg_137_ ( .D(n770), .CK(clk), .RN(rstn), .Q(dout[137]) );
  DFFRHQX1 dout_reg_188_ ( .D(n719), .CK(clk), .RN(rstn), .Q(dout[188]) );
  DFFRHQX1 dout_reg_187_ ( .D(n720), .CK(clk), .RN(rstn), .Q(dout[187]) );
  DFFRHQX1 dout_reg_186_ ( .D(n721), .CK(clk), .RN(rstn), .Q(dout[186]) );
  DFFRHQX1 dout_reg_185_ ( .D(n722), .CK(clk), .RN(rstn), .Q(dout[185]) );
  DFFRHQX1 dout_reg_172_ ( .D(n735), .CK(clk), .RN(rstn), .Q(dout[172]) );
  DFFRHQX1 dout_reg_171_ ( .D(n736), .CK(clk), .RN(rstn), .Q(dout[171]) );
  DFFRHQX1 dout_reg_170_ ( .D(n737), .CK(clk), .RN(rstn), .Q(dout[170]) );
  DFFRHQX1 dout_reg_169_ ( .D(n738), .CK(clk), .RN(rstn), .Q(dout[169]) );
  DFFRHQX1 dout_reg_156_ ( .D(n751), .CK(clk), .RN(rstn), .Q(dout[156]) );
  DFFRHQX1 dout_reg_155_ ( .D(n752), .CK(clk), .RN(rstn), .Q(dout[155]) );
  DFFRHQX1 dout_reg_154_ ( .D(n753), .CK(clk), .RN(rstn), .Q(dout[154]) );
  DFFRHQX1 dout_reg_153_ ( .D(n754), .CK(clk), .RN(rstn), .Q(dout[153]) );
  DFFRHQX1 dout_reg_236_ ( .D(n671), .CK(clk), .RN(rstn), .Q(dout[236]) );
  DFFRHQX1 dout_reg_235_ ( .D(n672), .CK(clk), .RN(rstn), .Q(dout[235]) );
  DFFRHQX1 dout_reg_234_ ( .D(n673), .CK(clk), .RN(rstn), .Q(dout[234]) );
  DFFRHQX1 dout_reg_233_ ( .D(n674), .CK(clk), .RN(rstn), .Q(dout[233]) );
  DFFRHQX1 dout_reg_204_ ( .D(n703), .CK(clk), .RN(rstn), .Q(dout[204]) );
  DFFRHQX1 dout_reg_203_ ( .D(n704), .CK(clk), .RN(rstn), .Q(dout[203]) );
  DFFRHQX1 dout_reg_202_ ( .D(n705), .CK(clk), .RN(rstn), .Q(dout[202]) );
  DFFRHQX1 dout_reg_201_ ( .D(n706), .CK(clk), .RN(rstn), .Q(dout[201]) );
  DFFRHQX1 dout_reg_136_ ( .D(n771), .CK(clk), .RN(rstn), .Q(dout[136]) );
  DFFRHQX1 dout_reg_135_ ( .D(n772), .CK(clk), .RN(rstn), .Q(dout[135]) );
  DFFRHQX1 dout_reg_134_ ( .D(n773), .CK(clk), .RN(rstn), .Q(dout[134]) );
  DFFRHQX1 dout_reg_133_ ( .D(n774), .CK(clk), .RN(rstn), .Q(dout[133]) );
  DFFRHQX1 dout_reg_132_ ( .D(n775), .CK(clk), .RN(rstn), .Q(dout[132]) );
  DFFRHQX1 dout_reg_131_ ( .D(n776), .CK(clk), .RN(rstn), .Q(dout[131]) );
  DFFRHQX1 dout_reg_130_ ( .D(n777), .CK(clk), .RN(rstn), .Q(dout[130]) );
  DFFRHQX1 dout_reg_184_ ( .D(n723), .CK(clk), .RN(rstn), .Q(dout[184]) );
  DFFRHQX1 dout_reg_183_ ( .D(n724), .CK(clk), .RN(rstn), .Q(dout[183]) );
  DFFRHQX1 dout_reg_182_ ( .D(n725), .CK(clk), .RN(rstn), .Q(dout[182]) );
  DFFRHQX1 dout_reg_181_ ( .D(n726), .CK(clk), .RN(rstn), .Q(dout[181]) );
  DFFRHQX1 dout_reg_180_ ( .D(n727), .CK(clk), .RN(rstn), .Q(dout[180]) );
  DFFRHQX1 dout_reg_179_ ( .D(n728), .CK(clk), .RN(rstn), .Q(dout[179]) );
  DFFRHQX1 dout_reg_178_ ( .D(n729), .CK(clk), .RN(rstn), .Q(dout[178]) );
  DFFRHQX1 dout_reg_168_ ( .D(n739), .CK(clk), .RN(rstn), .Q(dout[168]) );
  DFFRHQX1 dout_reg_167_ ( .D(n740), .CK(clk), .RN(rstn), .Q(dout[167]) );
  DFFRHQX1 dout_reg_166_ ( .D(n741), .CK(clk), .RN(rstn), .Q(dout[166]) );
  DFFRHQX1 dout_reg_165_ ( .D(n742), .CK(clk), .RN(rstn), .Q(dout[165]) );
  DFFRHQX1 dout_reg_164_ ( .D(n743), .CK(clk), .RN(rstn), .Q(dout[164]) );
  DFFRHQX1 dout_reg_163_ ( .D(n744), .CK(clk), .RN(rstn), .Q(dout[163]) );
  DFFRHQX1 dout_reg_162_ ( .D(n745), .CK(clk), .RN(rstn), .Q(dout[162]) );
  DFFRHQX1 dout_reg_152_ ( .D(n755), .CK(clk), .RN(rstn), .Q(dout[152]) );
  DFFRHQX1 dout_reg_151_ ( .D(n756), .CK(clk), .RN(rstn), .Q(dout[151]) );
  DFFRHQX1 dout_reg_150_ ( .D(n757), .CK(clk), .RN(rstn), .Q(dout[150]) );
  DFFRHQX1 dout_reg_149_ ( .D(n758), .CK(clk), .RN(rstn), .Q(dout[149]) );
  DFFRHQX1 dout_reg_148_ ( .D(n759), .CK(clk), .RN(rstn), .Q(dout[148]) );
  DFFRHQX1 dout_reg_147_ ( .D(n760), .CK(clk), .RN(rstn), .Q(dout[147]) );
  DFFRHQX1 dout_reg_146_ ( .D(n761), .CK(clk), .RN(rstn), .Q(dout[146]) );
  DFFRHQX1 dout_reg_224_ ( .D(n683), .CK(clk), .RN(rstn), .Q(dout[224]) );
  DFFRHQX1 dout_reg_192_ ( .D(n715), .CK(clk), .RN(rstn), .Q(dout[192]) );
  DFFRHQX1 dout_reg_226_ ( .D(n681), .CK(clk), .RN(rstn), .Q(dout[226]) );
  DFFRHQX1 dout_reg_225_ ( .D(n682), .CK(clk), .RN(rstn), .Q(dout[225]) );
  DFFRHQX1 dout_reg_194_ ( .D(n713), .CK(clk), .RN(rstn), .Q(dout[194]) );
  DFFRHQX1 dout_reg_193_ ( .D(n714), .CK(clk), .RN(rstn), .Q(dout[193]) );
  DFFRHQX1 dout_reg_227_ ( .D(n680), .CK(clk), .RN(rstn), .Q(dout[227]) );
  DFFRHQX1 dout_reg_195_ ( .D(n712), .CK(clk), .RN(rstn), .Q(dout[195]) );
  DFFRHQX1 dout_reg_128_ ( .D(n779), .CK(clk), .RN(rstn), .Q(dout[128]) );
  DFFRHQX1 dout_reg_176_ ( .D(n731), .CK(clk), .RN(rstn), .Q(dout[176]) );
  DFFRHQX1 dout_reg_160_ ( .D(n747), .CK(clk), .RN(rstn), .Q(dout[160]) );
  DFFRHQX1 dout_reg_144_ ( .D(n763), .CK(clk), .RN(rstn), .Q(dout[144]) );
  DFFRHQX1 dout_reg_129_ ( .D(n778), .CK(clk), .RN(rstn), .Q(dout[129]) );
  DFFRHQX1 dout_reg_177_ ( .D(n730), .CK(clk), .RN(rstn), .Q(dout[177]) );
  DFFRHQX1 dout_reg_161_ ( .D(n746), .CK(clk), .RN(rstn), .Q(dout[161]) );
  DFFRHQX1 dout_reg_145_ ( .D(n762), .CK(clk), .RN(rstn), .Q(dout[145]) );
  DFFRHQX1 dout_reg_229_ ( .D(n678), .CK(clk), .RN(rstn), .Q(dout[229]) );
  DFFRHQX1 dout_reg_228_ ( .D(n679), .CK(clk), .RN(rstn), .Q(dout[228]) );
  DFFRHQX1 dout_reg_197_ ( .D(n710), .CK(clk), .RN(rstn), .Q(dout[197]) );
  DFFRHQX1 dout_reg_196_ ( .D(n711), .CK(clk), .RN(rstn), .Q(dout[196]) );
  DFFRHQX1 dout_reg_230_ ( .D(n677), .CK(clk), .RN(rstn), .Q(dout[230]) );
  DFFRHQX1 dout_reg_198_ ( .D(n709), .CK(clk), .RN(rstn), .Q(dout[198]) );
  DFFRHQX1 dout_reg_232_ ( .D(n675), .CK(clk), .RN(rstn), .Q(dout[232]) );
  DFFRHQX1 dout_reg_231_ ( .D(n676), .CK(clk), .RN(rstn), .Q(dout[231]) );
  DFFRHQX1 dout_reg_200_ ( .D(n707), .CK(clk), .RN(rstn), .Q(dout[200]) );
  DFFRHQX1 dout_reg_199_ ( .D(n708), .CK(clk), .RN(rstn), .Q(dout[199]) );
  DFFRHQX1 even_odd_ready_reg ( .D(N275), .CK(clk), .RN(rstn), .Q(
        even_odd_ready) );
  NAND2X1 U3 ( .A(n929), .B(start), .Y(n2) );
  NAND2X1 U4 ( .A(n1026), .B(start), .Y(n19) );
  AND2X2 U5 ( .A(n927), .B(start), .Y(n20) );
  AND2X2 U6 ( .A(n928), .B(start), .Y(n149) );
  INVX1 U7 ( .A(n19), .Y(n170) );
  INVX1 U8 ( .A(n19), .Y(n172) );
  INVX1 U9 ( .A(n19), .Y(n173) );
  INVX1 U10 ( .A(n19), .Y(n175) );
  INVX1 U11 ( .A(n188), .Y(n187) );
  INVX1 U12 ( .A(n2), .Y(n176) );
  INVX1 U13 ( .A(n2), .Y(n178) );
  INVX1 U14 ( .A(n2), .Y(n179) );
  INVX1 U15 ( .A(n2), .Y(n181) );
  INVX1 U16 ( .A(start), .Y(n154) );
  INVX1 U17 ( .A(start), .Y(n150) );
  INVX1 U18 ( .A(start), .Y(n151) );
  INVX1 U19 ( .A(start), .Y(n152) );
  INVX1 U20 ( .A(n20), .Y(n166) );
  INVX1 U21 ( .A(n20), .Y(n167) );
  INVX1 U22 ( .A(n20), .Y(n169) );
  INVX1 U23 ( .A(n149), .Y(n164) );
  INVX1 U24 ( .A(n149), .Y(n163) );
  INVX1 U25 ( .A(n149), .Y(n161) );
  INVX1 U26 ( .A(n2), .Y(n182) );
  INVX1 U27 ( .A(n2), .Y(n184) );
  INVX1 U28 ( .A(n2), .Y(n185) );
  INVX1 U29 ( .A(start), .Y(n155) );
  INVX1 U30 ( .A(start), .Y(n157) );
  INVX1 U31 ( .A(start), .Y(n158) );
  INVX1 U32 ( .A(start), .Y(n160) );
  OR2X2 U33 ( .A(n927), .B(n928), .Y(n1026) );
  INVX1 U34 ( .A(N275), .Y(n188) );
  AOI2BB1X1 U35 ( .A0N(n929), .A1N(n1026), .B0(n154), .Y(N275) );
  NOR2X1 U36 ( .A(mode[0]), .B(mode[1]), .Y(n927) );
  NOR2X1 U37 ( .A(n910), .B(mode[1]), .Y(n928) );
  INVX1 U38 ( .A(mode[0]), .Y(n910) );
  INVX1 U39 ( .A(n1154), .Y(n891) );
  AOI222X1 U40 ( .A0(n178), .A1(din[32]), .B0(n170), .B1(din[16]), .C0(n154), 
        .C1(dout[16]), .Y(n1154) );
  INVX1 U41 ( .A(n1153), .Y(n890) );
  AOI222X1 U42 ( .A0(n181), .A1(din[33]), .B0(n170), .B1(din[17]), .C0(n157), 
        .C1(dout[17]), .Y(n1153) );
  INVX1 U43 ( .A(n1152), .Y(n889) );
  AOI222X1 U44 ( .A0(n184), .A1(din[34]), .B0(n170), .B1(din[18]), .C0(n154), 
        .C1(dout[18]), .Y(n1152) );
  INVX1 U45 ( .A(n1151), .Y(n888) );
  AOI222X1 U46 ( .A0(n179), .A1(din[35]), .B0(n170), .B1(din[19]), .C0(n154), 
        .C1(dout[19]), .Y(n1151) );
  INVX1 U47 ( .A(n1150), .Y(n887) );
  AOI222X1 U48 ( .A0(n176), .A1(din[36]), .B0(n170), .B1(din[20]), .C0(n154), 
        .C1(dout[20]), .Y(n1150) );
  INVX1 U49 ( .A(n1149), .Y(n886) );
  AOI222X1 U50 ( .A0(n178), .A1(din[37]), .B0(n170), .B1(din[21]), .C0(n154), 
        .C1(dout[21]), .Y(n1149) );
  INVX1 U51 ( .A(n1148), .Y(n885) );
  AOI222X1 U52 ( .A0(n181), .A1(din[38]), .B0(n170), .B1(din[22]), .C0(n154), 
        .C1(dout[22]), .Y(n1148) );
  INVX1 U53 ( .A(n1147), .Y(n884) );
  AOI222X1 U54 ( .A0(n179), .A1(din[39]), .B0(n170), .B1(din[23]), .C0(n154), 
        .C1(dout[23]), .Y(n1147) );
  INVX1 U55 ( .A(n1146), .Y(n883) );
  AOI222X1 U56 ( .A0(n176), .A1(din[40]), .B0(n170), .B1(din[24]), .C0(n154), 
        .C1(dout[24]), .Y(n1146) );
  INVX1 U57 ( .A(n1145), .Y(n882) );
  AOI222X1 U58 ( .A0(n178), .A1(din[41]), .B0(n170), .B1(din[25]), .C0(n154), 
        .C1(dout[25]), .Y(n1145) );
  INVX1 U59 ( .A(n1144), .Y(n881) );
  AOI222X1 U60 ( .A0(n181), .A1(din[42]), .B0(n170), .B1(din[26]), .C0(n155), 
        .C1(dout[26]), .Y(n1144) );
  INVX1 U61 ( .A(n1143), .Y(n880) );
  AOI222X1 U62 ( .A0(n179), .A1(din[43]), .B0(n170), .B1(din[27]), .C0(n155), 
        .C1(dout[27]), .Y(n1143) );
  INVX1 U63 ( .A(n1142), .Y(n879) );
  AOI222X1 U64 ( .A0(n182), .A1(din[44]), .B0(n172), .B1(din[28]), .C0(n155), 
        .C1(dout[28]), .Y(n1142) );
  INVX1 U65 ( .A(n1141), .Y(n878) );
  AOI222X1 U66 ( .A0(n182), .A1(din[45]), .B0(n172), .B1(din[29]), .C0(n155), 
        .C1(dout[29]), .Y(n1141) );
  INVX1 U67 ( .A(n1140), .Y(n877) );
  AOI222X1 U68 ( .A0(n182), .A1(din[46]), .B0(n172), .B1(din[30]), .C0(n155), 
        .C1(dout[30]), .Y(n1140) );
  INVX1 U69 ( .A(n1139), .Y(n876) );
  AOI222X1 U70 ( .A0(n182), .A1(din[47]), .B0(n172), .B1(din[31]), .C0(n155), 
        .C1(dout[31]), .Y(n1139) );
  INVX1 U71 ( .A(n1138), .Y(n875) );
  AOI222X1 U72 ( .A0(n182), .A1(din[64]), .B0(n172), .B1(din[32]), .C0(n155), 
        .C1(dout[32]), .Y(n1138) );
  INVX1 U73 ( .A(n1137), .Y(n874) );
  AOI222X1 U74 ( .A0(n182), .A1(din[65]), .B0(n172), .B1(din[33]), .C0(n155), 
        .C1(dout[33]), .Y(n1137) );
  INVX1 U75 ( .A(n1136), .Y(n873) );
  AOI222X1 U76 ( .A0(n182), .A1(din[66]), .B0(n172), .B1(din[34]), .C0(n155), 
        .C1(dout[34]), .Y(n1136) );
  INVX1 U77 ( .A(n1135), .Y(n872) );
  AOI222X1 U78 ( .A0(n182), .A1(din[67]), .B0(n172), .B1(din[35]), .C0(n155), 
        .C1(dout[35]), .Y(n1135) );
  INVX1 U79 ( .A(n1134), .Y(n871) );
  AOI222X1 U80 ( .A0(n182), .A1(din[68]), .B0(n172), .B1(din[36]), .C0(n155), 
        .C1(dout[36]), .Y(n1134) );
  INVX1 U81 ( .A(n1133), .Y(n870) );
  AOI222X1 U82 ( .A0(n182), .A1(din[69]), .B0(n172), .B1(din[37]), .C0(n155), 
        .C1(dout[37]), .Y(n1133) );
  INVX1 U83 ( .A(n1132), .Y(n869) );
  AOI222X1 U84 ( .A0(n182), .A1(din[70]), .B0(n172), .B1(din[38]), .C0(n155), 
        .C1(dout[38]), .Y(n1132) );
  INVX1 U85 ( .A(n1131), .Y(n868) );
  AOI222X1 U86 ( .A0(n182), .A1(din[71]), .B0(n172), .B1(din[39]), .C0(n155), 
        .C1(dout[39]), .Y(n1131) );
  INVX1 U87 ( .A(n1034), .Y(n771) );
  AOI222X1 U88 ( .A0(n176), .A1(din[24]), .B0(n172), .B1(din[136]), .C0(n160), 
        .C1(dout[136]), .Y(n1034) );
  INVX1 U89 ( .A(n1033), .Y(n770) );
  AOI222X1 U90 ( .A0(n178), .A1(din[25]), .B0(n172), .B1(din[137]), .C0(n154), 
        .C1(dout[137]), .Y(n1033) );
  INVX1 U91 ( .A(n1032), .Y(n769) );
  AOI222X1 U92 ( .A0(n181), .A1(din[26]), .B0(n172), .B1(din[138]), .C0(n154), 
        .C1(dout[138]), .Y(n1032) );
  INVX1 U93 ( .A(n1031), .Y(n768) );
  AOI222X1 U94 ( .A0(n179), .A1(din[27]), .B0(n170), .B1(din[139]), .C0(n154), 
        .C1(dout[139]), .Y(n1031) );
  INVX1 U95 ( .A(n1030), .Y(n767) );
  AOI222X1 U96 ( .A0(n176), .A1(din[28]), .B0(n170), .B1(din[140]), .C0(n154), 
        .C1(dout[140]), .Y(n1030) );
  INVX1 U97 ( .A(n1029), .Y(n766) );
  AOI222X1 U98 ( .A0(n178), .A1(din[29]), .B0(n173), .B1(din[141]), .C0(n154), 
        .C1(dout[141]), .Y(n1029) );
  INVX1 U99 ( .A(n1028), .Y(n765) );
  AOI222X1 U100 ( .A0(n181), .A1(din[30]), .B0(n175), .B1(din[142]), .C0(n154), 
        .C1(dout[142]), .Y(n1028) );
  INVX1 U101 ( .A(n1027), .Y(n764) );
  AOI222X1 U102 ( .A0(n179), .A1(din[31]), .B0(n170), .B1(din[143]), .C0(n154), 
        .C1(dout[143]), .Y(n1027) );
  INVX1 U103 ( .A(n1130), .Y(n867) );
  AOI222X1 U104 ( .A0(n182), .A1(din[72]), .B0(n173), .B1(din[40]), .C0(n155), 
        .C1(dout[40]), .Y(n1130) );
  INVX1 U105 ( .A(n1129), .Y(n866) );
  AOI222X1 U106 ( .A0(n182), .A1(din[73]), .B0(n173), .B1(din[41]), .C0(n155), 
        .C1(dout[41]), .Y(n1129) );
  INVX1 U107 ( .A(n1128), .Y(n865) );
  AOI222X1 U108 ( .A0(n182), .A1(din[74]), .B0(n173), .B1(din[42]), .C0(n155), 
        .C1(dout[42]), .Y(n1128) );
  INVX1 U109 ( .A(n1127), .Y(n864) );
  AOI222X1 U110 ( .A0(n182), .A1(din[75]), .B0(n173), .B1(din[43]), .C0(n155), 
        .C1(dout[43]), .Y(n1127) );
  INVX1 U111 ( .A(n1126), .Y(n863) );
  AOI222X1 U112 ( .A0(n182), .A1(din[76]), .B0(n173), .B1(din[44]), .C0(n155), 
        .C1(dout[44]), .Y(n1126) );
  INVX1 U113 ( .A(n1125), .Y(n862) );
  AOI222X1 U114 ( .A0(n182), .A1(din[77]), .B0(n173), .B1(din[45]), .C0(n155), 
        .C1(dout[45]), .Y(n1125) );
  INVX1 U115 ( .A(n1124), .Y(n861) );
  AOI222X1 U116 ( .A0(n182), .A1(din[78]), .B0(n173), .B1(din[46]), .C0(n155), 
        .C1(dout[46]), .Y(n1124) );
  INVX1 U117 ( .A(n1123), .Y(n860) );
  AOI222X1 U118 ( .A0(n182), .A1(din[79]), .B0(n173), .B1(din[47]), .C0(n155), 
        .C1(dout[47]), .Y(n1123) );
  INVX1 U119 ( .A(n1106), .Y(n843) );
  AOI222X1 U120 ( .A0(n184), .A1(din[128]), .B0(n175), .B1(din[64]), .C0(n154), 
        .C1(dout[64]), .Y(n1106) );
  INVX1 U121 ( .A(n1105), .Y(n842) );
  AOI222X1 U122 ( .A0(n184), .A1(din[129]), .B0(n175), .B1(din[65]), .C0(n157), 
        .C1(dout[65]), .Y(n1105) );
  INVX1 U123 ( .A(n1104), .Y(n841) );
  AOI222X1 U124 ( .A0(n184), .A1(din[130]), .B0(n175), .B1(din[66]), .C0(n157), 
        .C1(dout[66]), .Y(n1104) );
  INVX1 U125 ( .A(n1103), .Y(n840) );
  AOI222X1 U126 ( .A0(n184), .A1(din[131]), .B0(n175), .B1(din[67]), .C0(n157), 
        .C1(dout[67]), .Y(n1103) );
  INVX1 U127 ( .A(n1102), .Y(n839) );
  AOI222X1 U128 ( .A0(n184), .A1(din[132]), .B0(n175), .B1(din[68]), .C0(n157), 
        .C1(dout[68]), .Y(n1102) );
  INVX1 U129 ( .A(n1101), .Y(n838) );
  AOI222X1 U130 ( .A0(n184), .A1(din[133]), .B0(n175), .B1(din[69]), .C0(n157), 
        .C1(dout[69]), .Y(n1101) );
  INVX1 U131 ( .A(n1100), .Y(n837) );
  AOI222X1 U132 ( .A0(n184), .A1(din[134]), .B0(n175), .B1(din[70]), .C0(n157), 
        .C1(dout[70]), .Y(n1100) );
  INVX1 U133 ( .A(n1099), .Y(n836) );
  AOI222X1 U134 ( .A0(n184), .A1(din[135]), .B0(n175), .B1(din[71]), .C0(n157), 
        .C1(dout[71]), .Y(n1099) );
  INVX1 U135 ( .A(n1098), .Y(n835) );
  AOI222X1 U136 ( .A0(n184), .A1(din[136]), .B0(n175), .B1(din[72]), .C0(n157), 
        .C1(dout[72]), .Y(n1098) );
  INVX1 U137 ( .A(n1097), .Y(n834) );
  AOI222X1 U138 ( .A0(n184), .A1(din[137]), .B0(n175), .B1(din[73]), .C0(n157), 
        .C1(dout[73]), .Y(n1097) );
  INVX1 U139 ( .A(n1096), .Y(n833) );
  AOI222X1 U140 ( .A0(n184), .A1(din[138]), .B0(n175), .B1(din[74]), .C0(n157), 
        .C1(dout[74]), .Y(n1096) );
  INVX1 U141 ( .A(n1095), .Y(n832) );
  AOI222X1 U142 ( .A0(n184), .A1(din[139]), .B0(n175), .B1(din[75]), .C0(n157), 
        .C1(dout[75]), .Y(n1095) );
  INVX1 U143 ( .A(n1094), .Y(n831) );
  AOI222X1 U144 ( .A0(n184), .A1(din[140]), .B0(n173), .B1(din[76]), .C0(n157), 
        .C1(dout[76]), .Y(n1094) );
  INVX1 U145 ( .A(n1093), .Y(n830) );
  AOI222X1 U146 ( .A0(n184), .A1(din[141]), .B0(n170), .B1(din[77]), .C0(n157), 
        .C1(dout[77]), .Y(n1093) );
  INVX1 U147 ( .A(n1092), .Y(n829) );
  AOI222X1 U148 ( .A0(n184), .A1(din[142]), .B0(n170), .B1(din[78]), .C0(n157), 
        .C1(dout[78]), .Y(n1092) );
  INVX1 U149 ( .A(n1091), .Y(n828) );
  AOI222X1 U150 ( .A0(n184), .A1(din[143]), .B0(n175), .B1(din[79]), .C0(n157), 
        .C1(dout[79]), .Y(n1091) );
  INVX1 U151 ( .A(n1074), .Y(n811) );
  AOI222X1 U152 ( .A0(n185), .A1(din[192]), .B0(n170), .B1(din[96]), .C0(n158), 
        .C1(dout[96]), .Y(n1074) );
  INVX1 U153 ( .A(n1073), .Y(n810) );
  AOI222X1 U154 ( .A0(n185), .A1(din[193]), .B0(n173), .B1(din[97]), .C0(n158), 
        .C1(dout[97]), .Y(n1073) );
  INVX1 U155 ( .A(n1072), .Y(n809) );
  AOI222X1 U156 ( .A0(n185), .A1(din[194]), .B0(n172), .B1(din[98]), .C0(n158), 
        .C1(dout[98]), .Y(n1072) );
  INVX1 U157 ( .A(n1071), .Y(n808) );
  AOI222X1 U158 ( .A0(n185), .A1(din[195]), .B0(n173), .B1(din[99]), .C0(n158), 
        .C1(dout[99]), .Y(n1071) );
  INVX1 U159 ( .A(n1070), .Y(n807) );
  AOI222X1 U160 ( .A0(n185), .A1(din[196]), .B0(n173), .B1(din[100]), .C0(n158), .C1(dout[100]), .Y(n1070) );
  INVX1 U161 ( .A(n1069), .Y(n806) );
  AOI222X1 U162 ( .A0(n185), .A1(din[197]), .B0(n173), .B1(din[101]), .C0(n158), .C1(dout[101]), .Y(n1069) );
  INVX1 U163 ( .A(n1068), .Y(n805) );
  AOI222X1 U164 ( .A0(n185), .A1(din[198]), .B0(n172), .B1(din[102]), .C0(n158), .C1(dout[102]), .Y(n1068) );
  INVX1 U165 ( .A(n1067), .Y(n804) );
  AOI222X1 U166 ( .A0(n185), .A1(din[199]), .B0(n170), .B1(din[103]), .C0(n158), .C1(dout[103]), .Y(n1067) );
  INVX1 U167 ( .A(n1066), .Y(n803) );
  AOI222X1 U168 ( .A0(n185), .A1(din[200]), .B0(n175), .B1(din[104]), .C0(n158), .C1(dout[104]), .Y(n1066) );
  INVX1 U169 ( .A(n1065), .Y(n802) );
  AOI222X1 U170 ( .A0(n185), .A1(din[201]), .B0(n173), .B1(din[105]), .C0(n158), .C1(dout[105]), .Y(n1065) );
  INVX1 U171 ( .A(n1064), .Y(n801) );
  AOI222X1 U172 ( .A0(n185), .A1(din[202]), .B0(n173), .B1(din[106]), .C0(n158), .C1(dout[106]), .Y(n1064) );
  INVX1 U173 ( .A(n1063), .Y(n800) );
  AOI222X1 U174 ( .A0(n185), .A1(din[203]), .B0(n172), .B1(din[107]), .C0(n158), .C1(dout[107]), .Y(n1063) );
  INVX1 U175 ( .A(n1062), .Y(n799) );
  AOI222X1 U176 ( .A0(n185), .A1(din[204]), .B0(n170), .B1(din[108]), .C0(n158), .C1(dout[108]), .Y(n1062) );
  INVX1 U177 ( .A(n1061), .Y(n798) );
  AOI222X1 U178 ( .A0(n185), .A1(din[205]), .B0(n175), .B1(din[109]), .C0(n158), .C1(dout[109]), .Y(n1061) );
  INVX1 U179 ( .A(n1060), .Y(n797) );
  AOI222X1 U180 ( .A0(n185), .A1(din[206]), .B0(n173), .B1(din[110]), .C0(n158), .C1(dout[110]), .Y(n1060) );
  INVX1 U181 ( .A(n1059), .Y(n796) );
  AOI222X1 U182 ( .A0(n185), .A1(din[207]), .B0(n172), .B1(din[111]), .C0(n158), .C1(dout[111]), .Y(n1059) );
  INVX1 U183 ( .A(n1042), .Y(n779) );
  AOI222X1 U184 ( .A0(din[16]), .A1(n176), .B0(n175), .B1(din[128]), .C0(n160), 
        .C1(dout[128]), .Y(n1042) );
  INVX1 U185 ( .A(n1041), .Y(n778) );
  AOI222X1 U186 ( .A0(n179), .A1(din[17]), .B0(n175), .B1(din[129]), .C0(n160), 
        .C1(dout[129]), .Y(n1041) );
  INVX1 U187 ( .A(n1040), .Y(n777) );
  AOI222X1 U188 ( .A0(n176), .A1(din[18]), .B0(n172), .B1(din[130]), .C0(n160), 
        .C1(dout[130]), .Y(n1040) );
  INVX1 U189 ( .A(n1039), .Y(n776) );
  AOI222X1 U190 ( .A0(n178), .A1(din[19]), .B0(n173), .B1(din[131]), .C0(n160), 
        .C1(dout[131]), .Y(n1039) );
  INVX1 U191 ( .A(n1038), .Y(n775) );
  AOI222X1 U192 ( .A0(n181), .A1(din[20]), .B0(n172), .B1(din[132]), .C0(n160), 
        .C1(dout[132]), .Y(n1038) );
  INVX1 U193 ( .A(n1037), .Y(n774) );
  AOI222X1 U194 ( .A0(n179), .A1(din[21]), .B0(n175), .B1(din[133]), .C0(n160), 
        .C1(dout[133]), .Y(n1037) );
  INVX1 U195 ( .A(n1036), .Y(n773) );
  AOI222X1 U196 ( .A0(n176), .A1(din[22]), .B0(n170), .B1(din[134]), .C0(n160), 
        .C1(dout[134]), .Y(n1036) );
  INVX1 U197 ( .A(n1035), .Y(n772) );
  AOI222X1 U198 ( .A0(n178), .A1(din[23]), .B0(n173), .B1(din[135]), .C0(n160), 
        .C1(dout[135]), .Y(n1035) );
  INVX1 U199 ( .A(n1122), .Y(n859) );
  AOI222X1 U200 ( .A0(n182), .A1(din[96]), .B0(n173), .B1(din[48]), .C0(n155), 
        .C1(dout[48]), .Y(n1122) );
  INVX1 U201 ( .A(n1121), .Y(n858) );
  AOI222X1 U202 ( .A0(n182), .A1(din[97]), .B0(n173), .B1(din[49]), .C0(n155), 
        .C1(dout[49]), .Y(n1121) );
  INVX1 U203 ( .A(n1120), .Y(n857) );
  AOI222X1 U204 ( .A0(n182), .A1(din[98]), .B0(n173), .B1(din[50]), .C0(n155), 
        .C1(dout[50]), .Y(n1120) );
  INVX1 U205 ( .A(n1119), .Y(n856) );
  AOI222X1 U206 ( .A0(n182), .A1(din[99]), .B0(n173), .B1(din[51]), .C0(n155), 
        .C1(dout[51]), .Y(n1119) );
  INVX1 U207 ( .A(n1118), .Y(n855) );
  AOI222X1 U208 ( .A0(n182), .A1(din[100]), .B0(n172), .B1(din[52]), .C0(n155), 
        .C1(dout[52]), .Y(n1118) );
  INVX1 U209 ( .A(n1117), .Y(n854) );
  AOI222X1 U210 ( .A0(n182), .A1(din[101]), .B0(n175), .B1(din[53]), .C0(n155), 
        .C1(dout[53]), .Y(n1117) );
  INVX1 U211 ( .A(n1116), .Y(n853) );
  AOI222X1 U212 ( .A0(n182), .A1(din[102]), .B0(n170), .B1(din[54]), .C0(n155), 
        .C1(dout[54]), .Y(n1116) );
  INVX1 U213 ( .A(n1115), .Y(n852) );
  AOI222X1 U214 ( .A0(n182), .A1(din[103]), .B0(n173), .B1(din[55]), .C0(n155), 
        .C1(dout[55]), .Y(n1115) );
  INVX1 U215 ( .A(n1114), .Y(n851) );
  AOI222X1 U216 ( .A0(n182), .A1(din[104]), .B0(n172), .B1(din[56]), .C0(n155), 
        .C1(dout[56]), .Y(n1114) );
  INVX1 U217 ( .A(n1113), .Y(n850) );
  AOI222X1 U218 ( .A0(n182), .A1(din[105]), .B0(n175), .B1(din[57]), .C0(n155), 
        .C1(dout[57]), .Y(n1113) );
  INVX1 U219 ( .A(n1112), .Y(n849) );
  AOI222X1 U220 ( .A0(n182), .A1(din[106]), .B0(n170), .B1(din[58]), .C0(n157), 
        .C1(dout[58]), .Y(n1112) );
  INVX1 U221 ( .A(n1111), .Y(n848) );
  AOI222X1 U222 ( .A0(n182), .A1(din[107]), .B0(n173), .B1(din[59]), .C0(n157), 
        .C1(dout[59]), .Y(n1111) );
  INVX1 U223 ( .A(n1110), .Y(n847) );
  AOI222X1 U224 ( .A0(n184), .A1(din[108]), .B0(n172), .B1(din[60]), .C0(n157), 
        .C1(dout[60]), .Y(n1110) );
  INVX1 U225 ( .A(n1109), .Y(n846) );
  AOI222X1 U226 ( .A0(n184), .A1(din[109]), .B0(n175), .B1(din[61]), .C0(n157), 
        .C1(dout[61]), .Y(n1109) );
  INVX1 U227 ( .A(n1108), .Y(n845) );
  AOI222X1 U228 ( .A0(n184), .A1(din[110]), .B0(n170), .B1(din[62]), .C0(n157), 
        .C1(dout[62]), .Y(n1108) );
  INVX1 U229 ( .A(n1107), .Y(n844) );
  AOI222X1 U230 ( .A0(n184), .A1(din[111]), .B0(n173), .B1(din[63]), .C0(n157), 
        .C1(dout[63]), .Y(n1107) );
  INVX1 U231 ( .A(n1090), .Y(n827) );
  AOI222X1 U232 ( .A0(n184), .A1(din[160]), .B0(n172), .B1(din[80]), .C0(n157), 
        .C1(dout[80]), .Y(n1090) );
  INVX1 U233 ( .A(n1089), .Y(n826) );
  AOI222X1 U234 ( .A0(n184), .A1(din[161]), .B0(n172), .B1(din[81]), .C0(n157), 
        .C1(dout[81]), .Y(n1089) );
  INVX1 U235 ( .A(n1088), .Y(n825) );
  AOI222X1 U236 ( .A0(n184), .A1(din[162]), .B0(n173), .B1(din[82]), .C0(n157), 
        .C1(dout[82]), .Y(n1088) );
  INVX1 U237 ( .A(n1087), .Y(n824) );
  AOI222X1 U238 ( .A0(n184), .A1(din[163]), .B0(n173), .B1(din[83]), .C0(n157), 
        .C1(dout[83]), .Y(n1087) );
  INVX1 U239 ( .A(n1086), .Y(n823) );
  AOI222X1 U240 ( .A0(n184), .A1(din[164]), .B0(n170), .B1(din[84]), .C0(n157), 
        .C1(dout[84]), .Y(n1086) );
  INVX1 U241 ( .A(n1085), .Y(n822) );
  AOI222X1 U242 ( .A0(n184), .A1(din[165]), .B0(n175), .B1(din[85]), .C0(n157), 
        .C1(dout[85]), .Y(n1085) );
  INVX1 U243 ( .A(n1084), .Y(n821) );
  AOI222X1 U244 ( .A0(n184), .A1(din[166]), .B0(n172), .B1(din[86]), .C0(n157), 
        .C1(dout[86]), .Y(n1084) );
  INVX1 U245 ( .A(n1083), .Y(n820) );
  AOI222X1 U246 ( .A0(n184), .A1(din[167]), .B0(n170), .B1(din[87]), .C0(n157), 
        .C1(dout[87]), .Y(n1083) );
  INVX1 U247 ( .A(n1082), .Y(n819) );
  AOI222X1 U248 ( .A0(n184), .A1(din[168]), .B0(n175), .B1(din[88]), .C0(n157), 
        .C1(dout[88]), .Y(n1082) );
  INVX1 U249 ( .A(n1081), .Y(n818) );
  AOI222X1 U250 ( .A0(n184), .A1(din[169]), .B0(n172), .B1(din[89]), .C0(n157), 
        .C1(dout[89]), .Y(n1081) );
  INVX1 U251 ( .A(n1080), .Y(n817) );
  AOI222X1 U252 ( .A0(n184), .A1(din[170]), .B0(n172), .B1(din[90]), .C0(n158), 
        .C1(dout[90]), .Y(n1080) );
  INVX1 U253 ( .A(n1079), .Y(n816) );
  AOI222X1 U254 ( .A0(n185), .A1(din[171]), .B0(n170), .B1(din[91]), .C0(n158), 
        .C1(dout[91]), .Y(n1079) );
  INVX1 U255 ( .A(n1078), .Y(n815) );
  AOI222X1 U256 ( .A0(n185), .A1(din[172]), .B0(n173), .B1(din[92]), .C0(n158), 
        .C1(dout[92]), .Y(n1078) );
  INVX1 U257 ( .A(n1077), .Y(n814) );
  AOI222X1 U258 ( .A0(n185), .A1(din[173]), .B0(n175), .B1(din[93]), .C0(n158), 
        .C1(dout[93]), .Y(n1077) );
  INVX1 U259 ( .A(n1076), .Y(n813) );
  AOI222X1 U260 ( .A0(n185), .A1(din[174]), .B0(n175), .B1(din[94]), .C0(n158), 
        .C1(dout[94]), .Y(n1076) );
  INVX1 U261 ( .A(n1075), .Y(n812) );
  AOI222X1 U262 ( .A0(n185), .A1(din[175]), .B0(n175), .B1(din[95]), .C0(n158), 
        .C1(dout[95]), .Y(n1075) );
  INVX1 U263 ( .A(n1058), .Y(n795) );
  AOI222X1 U264 ( .A0(n185), .A1(din[224]), .B0(n172), .B1(din[112]), .C0(n158), .C1(dout[112]), .Y(n1058) );
  INVX1 U265 ( .A(n1057), .Y(n794) );
  AOI222X1 U266 ( .A0(n185), .A1(din[225]), .B0(n170), .B1(din[113]), .C0(n158), .C1(dout[113]), .Y(n1057) );
  INVX1 U267 ( .A(n1056), .Y(n793) );
  AOI222X1 U268 ( .A0(n185), .A1(din[226]), .B0(n170), .B1(din[114]), .C0(n158), .C1(dout[114]), .Y(n1056) );
  INVX1 U269 ( .A(n1055), .Y(n792) );
  AOI222X1 U270 ( .A0(n185), .A1(din[227]), .B0(n173), .B1(din[115]), .C0(n158), .C1(dout[115]), .Y(n1055) );
  INVX1 U271 ( .A(n1054), .Y(n791) );
  AOI222X1 U272 ( .A0(n185), .A1(din[228]), .B0(n170), .B1(din[116]), .C0(n158), .C1(dout[116]), .Y(n1054) );
  INVX1 U273 ( .A(n1053), .Y(n790) );
  AOI222X1 U274 ( .A0(n185), .A1(din[229]), .B0(n175), .B1(din[117]), .C0(n158), .C1(dout[117]), .Y(n1053) );
  INVX1 U275 ( .A(n1052), .Y(n789) );
  AOI222X1 U276 ( .A0(n185), .A1(din[230]), .B0(n175), .B1(din[118]), .C0(n158), .C1(dout[118]), .Y(n1052) );
  INVX1 U277 ( .A(n1051), .Y(n788) );
  AOI222X1 U278 ( .A0(n185), .A1(din[231]), .B0(n170), .B1(din[119]), .C0(n158), .C1(dout[119]), .Y(n1051) );
  INVX1 U279 ( .A(n1050), .Y(n787) );
  AOI222X1 U280 ( .A0(n185), .A1(din[232]), .B0(n173), .B1(din[120]), .C0(n158), .C1(dout[120]), .Y(n1050) );
  INVX1 U281 ( .A(n1049), .Y(n786) );
  AOI222X1 U282 ( .A0(n185), .A1(din[233]), .B0(n173), .B1(din[121]), .C0(n158), .C1(dout[121]), .Y(n1049) );
  INVX1 U283 ( .A(n1048), .Y(n785) );
  AOI222X1 U284 ( .A0(n185), .A1(din[234]), .B0(n175), .B1(din[122]), .C0(n160), .C1(dout[122]), .Y(n1048) );
  INVX1 U285 ( .A(n1047), .Y(n784) );
  AOI222X1 U286 ( .A0(n176), .A1(din[235]), .B0(n175), .B1(din[123]), .C0(n160), .C1(dout[123]), .Y(n1047) );
  INVX1 U287 ( .A(n1046), .Y(n783) );
  AOI222X1 U288 ( .A0(n179), .A1(din[236]), .B0(n170), .B1(din[124]), .C0(n160), .C1(dout[124]), .Y(n1046) );
  INVX1 U289 ( .A(n1045), .Y(n782) );
  AOI222X1 U290 ( .A0(n181), .A1(din[237]), .B0(n172), .B1(din[125]), .C0(n160), .C1(dout[125]), .Y(n1045) );
  INVX1 U291 ( .A(n1044), .Y(n781) );
  AOI222X1 U292 ( .A0(n178), .A1(din[238]), .B0(n175), .B1(din[126]), .C0(n160), .C1(dout[126]), .Y(n1044) );
  INVX1 U293 ( .A(n1043), .Y(n780) );
  AOI222X1 U294 ( .A0(n178), .A1(din[239]), .B0(n172), .B1(din[127]), .C0(n160), .C1(dout[127]), .Y(n1043) );
  OAI221XL U295 ( .A0(n646), .A1(n167), .B0(n161), .B1(n265), .C0(n976), .Y(
        n714) );
  AOI22X1 U296 ( .A0(din[49]), .A1(n179), .B0(dout[193]), .B1(n151), .Y(n976)
         );
  OAI221XL U297 ( .A0(n643), .A1(n169), .B0(n161), .B1(n261), .C0(n975), .Y(
        n713) );
  AOI22X1 U298 ( .A0(din[50]), .A1(n181), .B0(dout[194]), .B1(n150), .Y(n975)
         );
  OAI221XL U299 ( .A0(n640), .A1(n169), .B0(n164), .B1(n256), .C0(n974), .Y(
        n712) );
  AOI22X1 U300 ( .A0(din[51]), .A1(n178), .B0(dout[195]), .B1(n160), .Y(n974)
         );
  OAI221XL U301 ( .A0(n637), .A1(n166), .B0(n163), .B1(n252), .C0(n973), .Y(
        n711) );
  AOI22X1 U302 ( .A0(din[52]), .A1(n178), .B0(dout[196]), .B1(n151), .Y(n973)
         );
  OAI221XL U303 ( .A0(n634), .A1(n169), .B0(n164), .B1(n247), .C0(n972), .Y(
        n710) );
  AOI22X1 U304 ( .A0(din[53]), .A1(n178), .B0(dout[197]), .B1(n152), .Y(n972)
         );
  OAI221XL U305 ( .A0(n631), .A1(n169), .B0(n161), .B1(n243), .C0(n971), .Y(
        n709) );
  AOI22X1 U306 ( .A0(din[54]), .A1(n178), .B0(dout[198]), .B1(n151), .Y(n971)
         );
  OAI221XL U307 ( .A0(n628), .A1(n169), .B0(n164), .B1(n238), .C0(n970), .Y(
        n708) );
  AOI22X1 U308 ( .A0(din[55]), .A1(n178), .B0(dout[199]), .B1(n150), .Y(n970)
         );
  OAI221XL U309 ( .A0(n625), .A1(n167), .B0(n163), .B1(n234), .C0(n969), .Y(
        n707) );
  AOI22X1 U310 ( .A0(din[56]), .A1(n178), .B0(dout[200]), .B1(n160), .Y(n969)
         );
  OAI221XL U311 ( .A0(n325), .A1(n169), .B0(n164), .B1(n229), .C0(n968), .Y(
        n706) );
  AOI22X1 U312 ( .A0(din[57]), .A1(n178), .B0(dout[201]), .B1(n160), .Y(n968)
         );
  OAI221XL U313 ( .A0(n319), .A1(n166), .B0(n164), .B1(n223), .C0(n967), .Y(
        n705) );
  AOI22X1 U314 ( .A0(din[58]), .A1(n178), .B0(dout[202]), .B1(n160), .Y(n967)
         );
  OAI221XL U315 ( .A0(n313), .A1(n167), .B0(n164), .B1(n217), .C0(n966), .Y(
        n704) );
  AOI22X1 U316 ( .A0(din[59]), .A1(n178), .B0(dout[203]), .B1(n152), .Y(n966)
         );
  OAI221XL U317 ( .A0(n307), .A1(n169), .B0(n164), .B1(n211), .C0(n965), .Y(
        n703) );
  AOI22X1 U318 ( .A0(din[60]), .A1(n178), .B0(dout[204]), .B1(n151), .Y(n965)
         );
  OAI221XL U319 ( .A0(n301), .A1(n169), .B0(n164), .B1(n205), .C0(n964), .Y(
        n702) );
  AOI22X1 U320 ( .A0(din[61]), .A1(n178), .B0(dout[205]), .B1(n151), .Y(n964)
         );
  OAI221XL U321 ( .A0(n295), .A1(n169), .B0(n164), .B1(n199), .C0(n963), .Y(
        n701) );
  AOI22X1 U322 ( .A0(din[62]), .A1(n178), .B0(dout[206]), .B1(n151), .Y(n963)
         );
  OAI221XL U323 ( .A0(n274), .A1(n169), .B0(n164), .B1(n194), .C0(n962), .Y(
        n700) );
  AOI22X1 U324 ( .A0(din[63]), .A1(n178), .B0(dout[207]), .B1(n151), .Y(n962)
         );
  OAI221XL U325 ( .A0(n167), .A1(n648), .B0(n164), .B1(n267), .C0(n961), .Y(
        n699) );
  AOI22X1 U326 ( .A0(din[112]), .A1(n179), .B0(dout[208]), .B1(n151), .Y(n961)
         );
  OAI221XL U327 ( .A0(n169), .A1(n645), .B0(n164), .B1(n262), .C0(n960), .Y(
        n698) );
  AOI22X1 U328 ( .A0(din[113]), .A1(n179), .B0(dout[209]), .B1(n151), .Y(n960)
         );
  OAI221XL U329 ( .A0(n166), .A1(n642), .B0(n164), .B1(n258), .C0(n959), .Y(
        n697) );
  AOI22X1 U330 ( .A0(din[114]), .A1(n179), .B0(dout[210]), .B1(n151), .Y(n959)
         );
  OAI221XL U331 ( .A0(n167), .A1(n639), .B0(n164), .B1(n253), .C0(n958), .Y(
        n696) );
  AOI22X1 U332 ( .A0(din[115]), .A1(n179), .B0(dout[211]), .B1(n151), .Y(n958)
         );
  OAI221XL U333 ( .A0(n166), .A1(n636), .B0(n164), .B1(n249), .C0(n957), .Y(
        n695) );
  AOI22X1 U334 ( .A0(din[116]), .A1(n179), .B0(dout[212]), .B1(n151), .Y(n957)
         );
  OAI221XL U335 ( .A0(n167), .A1(n633), .B0(n164), .B1(n244), .C0(n956), .Y(
        n694) );
  AOI22X1 U336 ( .A0(din[117]), .A1(n179), .B0(dout[213]), .B1(n151), .Y(n956)
         );
  OAI221XL U337 ( .A0(n169), .A1(n630), .B0(n163), .B1(n240), .C0(n955), .Y(
        n693) );
  AOI22X1 U338 ( .A0(din[118]), .A1(n179), .B0(dout[214]), .B1(n152), .Y(n955)
         );
  OAI221XL U339 ( .A0(n169), .A1(n627), .B0(n163), .B1(n235), .C0(n954), .Y(
        n692) );
  AOI22X1 U340 ( .A0(din[119]), .A1(n179), .B0(dout[215]), .B1(n152), .Y(n954)
         );
  OAI221XL U341 ( .A0(n167), .A1(n624), .B0(n163), .B1(n231), .C0(n953), .Y(
        n691) );
  AOI22X1 U342 ( .A0(din[120]), .A1(n179), .B0(dout[216]), .B1(n152), .Y(n953)
         );
  OAI221XL U343 ( .A0(n166), .A1(n323), .B0(n163), .B1(n225), .C0(n952), .Y(
        n690) );
  AOI22X1 U344 ( .A0(din[121]), .A1(n179), .B0(dout[217]), .B1(n152), .Y(n952)
         );
  OAI221XL U345 ( .A0(n167), .A1(n317), .B0(n163), .B1(n219), .C0(n951), .Y(
        n689) );
  AOI22X1 U346 ( .A0(din[122]), .A1(n179), .B0(dout[218]), .B1(n152), .Y(n951)
         );
  OAI221XL U347 ( .A0(n169), .A1(n311), .B0(n163), .B1(n213), .C0(n950), .Y(
        n688) );
  AOI22X1 U348 ( .A0(din[123]), .A1(n179), .B0(dout[219]), .B1(n152), .Y(n950)
         );
  OAI221XL U349 ( .A0(n169), .A1(n305), .B0(n163), .B1(n207), .C0(n949), .Y(
        n687) );
  AOI22X1 U350 ( .A0(din[124]), .A1(n179), .B0(dout[220]), .B1(n152), .Y(n949)
         );
  OAI221XL U351 ( .A0(n166), .A1(n299), .B0(n163), .B1(n201), .C0(n948), .Y(
        n686) );
  AOI22X1 U352 ( .A0(din[125]), .A1(n181), .B0(dout[221]), .B1(n152), .Y(n948)
         );
  OAI221XL U353 ( .A0(n166), .A1(n277), .B0(n163), .B1(n196), .C0(n947), .Y(
        n685) );
  AOI22X1 U354 ( .A0(din[126]), .A1(n181), .B0(dout[222]), .B1(n151), .Y(n947)
         );
  OAI221XL U355 ( .A0(n167), .A1(n273), .B0(n163), .B1(n191), .C0(n946), .Y(
        n684) );
  AOI22X1 U356 ( .A0(din[127]), .A1(n181), .B0(dout[223]), .B1(n152), .Y(n946)
         );
  OAI221XL U357 ( .A0(n647), .A1(n169), .B0(n163), .B1(n648), .C0(n945), .Y(
        n683) );
  AOI22X1 U358 ( .A0(din[176]), .A1(n181), .B0(dout[224]), .B1(n152), .Y(n945)
         );
  OAI221XL U359 ( .A0(n644), .A1(n167), .B0(n163), .B1(n645), .C0(n944), .Y(
        n682) );
  AOI22X1 U360 ( .A0(din[177]), .A1(n181), .B0(dout[225]), .B1(n152), .Y(n944)
         );
  OAI221XL U361 ( .A0(n641), .A1(n167), .B0(n163), .B1(n642), .C0(n943), .Y(
        n681) );
  AOI22X1 U362 ( .A0(din[178]), .A1(n181), .B0(dout[226]), .B1(n151), .Y(n943)
         );
  OAI221XL U363 ( .A0(n638), .A1(n166), .B0(n161), .B1(n639), .C0(n942), .Y(
        n680) );
  AOI22X1 U364 ( .A0(din[179]), .A1(n181), .B0(dout[227]), .B1(n151), .Y(n942)
         );
  OAI221XL U365 ( .A0(n635), .A1(n169), .B0(n161), .B1(n636), .C0(n941), .Y(
        n679) );
  AOI22X1 U366 ( .A0(din[180]), .A1(n181), .B0(dout[228]), .B1(n151), .Y(n941)
         );
  OAI221XL U367 ( .A0(n632), .A1(n166), .B0(n161), .B1(n633), .C0(n940), .Y(
        n678) );
  AOI22X1 U368 ( .A0(din[181]), .A1(n181), .B0(dout[229]), .B1(n152), .Y(n940)
         );
  OAI221XL U369 ( .A0(n629), .A1(n167), .B0(n161), .B1(n630), .C0(n939), .Y(
        n677) );
  AOI22X1 U370 ( .A0(din[182]), .A1(n181), .B0(dout[230]), .B1(n150), .Y(n939)
         );
  OAI221XL U371 ( .A0(n626), .A1(n166), .B0(n161), .B1(n627), .C0(n938), .Y(
        n676) );
  AOI22X1 U372 ( .A0(din[183]), .A1(n181), .B0(dout[231]), .B1(n150), .Y(n938)
         );
  OAI221XL U373 ( .A0(n623), .A1(n169), .B0(n161), .B1(n624), .C0(n937), .Y(
        n675) );
  AOI22X1 U374 ( .A0(din[184]), .A1(n181), .B0(dout[232]), .B1(n151), .Y(n937)
         );
  OAI221XL U375 ( .A0(n321), .A1(n169), .B0(n161), .B1(n323), .C0(n936), .Y(
        n674) );
  AOI22X1 U376 ( .A0(din[185]), .A1(n181), .B0(dout[233]), .B1(n151), .Y(n936)
         );
  OAI221XL U377 ( .A0(n315), .A1(n167), .B0(n161), .B1(n317), .C0(n935), .Y(
        n673) );
  AOI22X1 U378 ( .A0(din[186]), .A1(n176), .B0(dout[234]), .B1(n150), .Y(n935)
         );
  OAI221XL U379 ( .A0(n309), .A1(n169), .B0(n161), .B1(n311), .C0(n934), .Y(
        n672) );
  AOI22X1 U380 ( .A0(din[187]), .A1(n181), .B0(dout[235]), .B1(n152), .Y(n934)
         );
  OAI221XL U381 ( .A0(n303), .A1(n169), .B0(n161), .B1(n305), .C0(n933), .Y(
        n671) );
  AOI22X1 U382 ( .A0(din[188]), .A1(n178), .B0(dout[236]), .B1(n152), .Y(n933)
         );
  OAI221XL U383 ( .A0(n297), .A1(n167), .B0(n161), .B1(n299), .C0(n932), .Y(
        n670) );
  AOI22X1 U384 ( .A0(din[189]), .A1(n179), .B0(dout[237]), .B1(n150), .Y(n932)
         );
  OAI221XL U385 ( .A0(n276), .A1(n169), .B0(n161), .B1(n277), .C0(n931), .Y(
        n669) );
  AOI22X1 U386 ( .A0(din[190]), .A1(n181), .B0(dout[238]), .B1(n152), .Y(n931)
         );
  OAI221XL U387 ( .A0(n271), .A1(n169), .B0(n161), .B1(n273), .C0(n930), .Y(
        n668) );
  AOI22X1 U388 ( .A0(din[191]), .A1(n179), .B0(dout[239]), .B1(n152), .Y(n930)
         );
  OAI221XL U389 ( .A0(n169), .A1(n270), .B0(n268), .B1(n164), .C0(n1025), .Y(
        n763) );
  AOI22X1 U390 ( .A0(din[80]), .A1(n176), .B0(dout[144]), .B1(n150), .Y(n1025)
         );
  OAI221XL U391 ( .A0(n166), .A1(n265), .B0(n264), .B1(n161), .C0(n1024), .Y(
        n762) );
  AOI22X1 U392 ( .A0(din[81]), .A1(n176), .B0(dout[145]), .B1(n150), .Y(n1024)
         );
  OAI221XL U393 ( .A0(n167), .A1(n261), .B0(n259), .B1(n163), .C0(n1023), .Y(
        n761) );
  AOI22X1 U394 ( .A0(din[82]), .A1(n176), .B0(dout[146]), .B1(n150), .Y(n1023)
         );
  OAI221XL U395 ( .A0(n167), .A1(n256), .B0(n255), .B1(n164), .C0(n1022), .Y(
        n760) );
  AOI22X1 U396 ( .A0(din[83]), .A1(n176), .B0(dout[147]), .B1(n160), .Y(n1022)
         );
  OAI221XL U397 ( .A0(n167), .A1(n252), .B0(n250), .B1(n161), .C0(n1021), .Y(
        n759) );
  AOI22X1 U398 ( .A0(din[84]), .A1(n176), .B0(dout[148]), .B1(n151), .Y(n1021)
         );
  OAI221XL U399 ( .A0(n167), .A1(n247), .B0(n246), .B1(n163), .C0(n1020), .Y(
        n758) );
  AOI22X1 U400 ( .A0(din[85]), .A1(n176), .B0(dout[149]), .B1(n154), .Y(n1020)
         );
  OAI221XL U401 ( .A0(n166), .A1(n243), .B0(n241), .B1(n163), .C0(n1019), .Y(
        n757) );
  AOI22X1 U402 ( .A0(din[86]), .A1(n176), .B0(dout[150]), .B1(n152), .Y(n1019)
         );
  OAI221XL U403 ( .A0(n167), .A1(n238), .B0(n237), .B1(n161), .C0(n1018), .Y(
        n756) );
  AOI22X1 U404 ( .A0(din[87]), .A1(n176), .B0(dout[151]), .B1(n151), .Y(n1018)
         );
  OAI221XL U405 ( .A0(n167), .A1(n234), .B0(n232), .B1(n164), .C0(n1017), .Y(
        n755) );
  AOI22X1 U406 ( .A0(din[88]), .A1(n176), .B0(dout[152]), .B1(n152), .Y(n1017)
         );
  OAI221XL U407 ( .A0(n167), .A1(n229), .B0(n227), .B1(n163), .C0(n1016), .Y(
        n754) );
  AOI22X1 U408 ( .A0(din[89]), .A1(n176), .B0(dout[153]), .B1(n150), .Y(n1016)
         );
  OAI221XL U409 ( .A0(n166), .A1(n223), .B0(n221), .B1(n161), .C0(n1015), .Y(
        n753) );
  AOI22X1 U410 ( .A0(din[90]), .A1(n176), .B0(dout[154]), .B1(n151), .Y(n1015)
         );
  OAI221XL U411 ( .A0(n166), .A1(n217), .B0(n215), .B1(n164), .C0(n1014), .Y(
        n752) );
  AOI22X1 U412 ( .A0(din[91]), .A1(n176), .B0(dout[155]), .B1(n150), .Y(n1014)
         );
  OAI221XL U413 ( .A0(n166), .A1(n211), .B0(n209), .B1(n163), .C0(n1013), .Y(
        n751) );
  AOI22X1 U414 ( .A0(din[92]), .A1(n176), .B0(dout[156]), .B1(n150), .Y(n1013)
         );
  OAI221XL U415 ( .A0(n167), .A1(n205), .B0(n203), .B1(n161), .C0(n1012), .Y(
        n750) );
  AOI22X1 U416 ( .A0(din[93]), .A1(n178), .B0(dout[157]), .B1(n150), .Y(n1012)
         );
  OAI221XL U417 ( .A0(n166), .A1(n199), .B0(n197), .B1(n161), .C0(n1011), .Y(
        n749) );
  AOI22X1 U418 ( .A0(din[94]), .A1(n181), .B0(dout[158]), .B1(n150), .Y(n1011)
         );
  OAI221XL U419 ( .A0(n167), .A1(n194), .B0(n193), .B1(n164), .C0(n1010), .Y(
        n748) );
  AOI22X1 U420 ( .A0(din[95]), .A1(n176), .B0(dout[159]), .B1(n150), .Y(n1010)
         );
  OAI221XL U421 ( .A0(n268), .A1(n166), .B0(n649), .B1(n163), .C0(n1009), .Y(
        n747) );
  AOI22X1 U422 ( .A0(din[144]), .A1(n181), .B0(dout[160]), .B1(n150), .Y(n1009) );
  OAI221XL U423 ( .A0(n264), .A1(n169), .B0(n646), .B1(n164), .C0(n1008), .Y(
        n746) );
  AOI22X1 U424 ( .A0(din[145]), .A1(n181), .B0(dout[161]), .B1(n150), .Y(n1008) );
  OAI221XL U425 ( .A0(n259), .A1(n169), .B0(n643), .B1(n163), .C0(n1007), .Y(
        n745) );
  AOI22X1 U426 ( .A0(din[146]), .A1(n178), .B0(dout[162]), .B1(n150), .Y(n1007) );
  OAI221XL U427 ( .A0(n255), .A1(n167), .B0(n640), .B1(n161), .C0(n1006), .Y(
        n744) );
  AOI22X1 U428 ( .A0(din[147]), .A1(n179), .B0(dout[163]), .B1(n150), .Y(n1006) );
  OAI221XL U429 ( .A0(n250), .A1(n169), .B0(n637), .B1(n164), .C0(n1005), .Y(
        n743) );
  AOI22X1 U430 ( .A0(din[148]), .A1(n181), .B0(dout[164]), .B1(n150), .Y(n1005) );
  OAI221XL U431 ( .A0(n246), .A1(n169), .B0(n634), .B1(n163), .C0(n1004), .Y(
        n742) );
  AOI22X1 U432 ( .A0(din[149]), .A1(n176), .B0(dout[165]), .B1(n150), .Y(n1004) );
  OAI221XL U433 ( .A0(n241), .A1(n166), .B0(n631), .B1(n161), .C0(n1003), .Y(
        n741) );
  AOI22X1 U434 ( .A0(din[150]), .A1(n181), .B0(dout[166]), .B1(n150), .Y(n1003) );
  OAI221XL U435 ( .A0(n237), .A1(n167), .B0(n628), .B1(n164), .C0(n1002), .Y(
        n740) );
  AOI22X1 U436 ( .A0(din[151]), .A1(n179), .B0(dout[167]), .B1(n152), .Y(n1002) );
  OAI221XL U437 ( .A0(n232), .A1(n169), .B0(n625), .B1(n161), .C0(n1001), .Y(
        n739) );
  AOI22X1 U438 ( .A0(din[152]), .A1(n178), .B0(dout[168]), .B1(n152), .Y(n1001) );
  OAI221XL U439 ( .A0(n227), .A1(n167), .B0(n325), .B1(n163), .C0(n1000), .Y(
        n738) );
  AOI22X1 U440 ( .A0(din[153]), .A1(n179), .B0(dout[169]), .B1(n150), .Y(n1000) );
  OAI221XL U441 ( .A0(n221), .A1(n169), .B0(n319), .B1(n161), .C0(n999), .Y(
        n737) );
  AOI22X1 U442 ( .A0(din[154]), .A1(n179), .B0(dout[170]), .B1(n150), .Y(n999)
         );
  OAI221XL U443 ( .A0(n215), .A1(n167), .B0(n313), .B1(n164), .C0(n998), .Y(
        n736) );
  AOI22X1 U444 ( .A0(din[155]), .A1(n181), .B0(dout[171]), .B1(n151), .Y(n998)
         );
  OAI221XL U445 ( .A0(n209), .A1(n167), .B0(n307), .B1(n164), .C0(n997), .Y(
        n735) );
  AOI22X1 U446 ( .A0(din[156]), .A1(n176), .B0(dout[172]), .B1(n160), .Y(n997)
         );
  OAI221XL U447 ( .A0(n203), .A1(n167), .B0(n301), .B1(n161), .C0(n996), .Y(
        n734) );
  AOI22X1 U448 ( .A0(din[157]), .A1(n178), .B0(dout[173]), .B1(n160), .Y(n996)
         );
  OAI221XL U449 ( .A0(n197), .A1(n166), .B0(n295), .B1(n163), .C0(n995), .Y(
        n733) );
  AOI22X1 U450 ( .A0(din[158]), .A1(n178), .B0(dout[174]), .B1(n152), .Y(n995)
         );
  OAI221XL U451 ( .A0(n193), .A1(n167), .B0(n274), .B1(n161), .C0(n994), .Y(
        n732) );
  AOI22X1 U452 ( .A0(din[159]), .A1(n176), .B0(dout[175]), .B1(n160), .Y(n994)
         );
  OAI221XL U453 ( .A0(n166), .A1(n267), .B0(n647), .B1(n164), .C0(n993), .Y(
        n731) );
  AOI22X1 U454 ( .A0(din[208]), .A1(n179), .B0(dout[176]), .B1(n154), .Y(n993)
         );
  OAI221XL U455 ( .A0(n166), .A1(n262), .B0(n644), .B1(n163), .C0(n992), .Y(
        n730) );
  AOI22X1 U456 ( .A0(din[209]), .A1(n176), .B0(dout[177]), .B1(n160), .Y(n992)
         );
  OAI221XL U457 ( .A0(n166), .A1(n258), .B0(n641), .B1(n161), .C0(n991), .Y(
        n729) );
  AOI22X1 U458 ( .A0(din[210]), .A1(n179), .B0(dout[178]), .B1(n151), .Y(n991)
         );
  OAI221XL U459 ( .A0(n166), .A1(n253), .B0(n638), .B1(n164), .C0(n990), .Y(
        n728) );
  AOI22X1 U460 ( .A0(din[211]), .A1(n176), .B0(dout[179]), .B1(n152), .Y(n990)
         );
  OAI221XL U461 ( .A0(n166), .A1(n249), .B0(n635), .B1(n161), .C0(n989), .Y(
        n727) );
  AOI22X1 U462 ( .A0(din[212]), .A1(n178), .B0(dout[180]), .B1(n151), .Y(n989)
         );
  OAI221XL U463 ( .A0(n166), .A1(n244), .B0(n632), .B1(n164), .C0(n988), .Y(
        n726) );
  AOI22X1 U464 ( .A0(din[213]), .A1(n181), .B0(dout[181]), .B1(n160), .Y(n988)
         );
  OAI221XL U465 ( .A0(n166), .A1(n240), .B0(n629), .B1(n163), .C0(n987), .Y(
        n725) );
  AOI22X1 U466 ( .A0(din[214]), .A1(n176), .B0(dout[182]), .B1(n152), .Y(n987)
         );
  OAI221XL U467 ( .A0(n166), .A1(n235), .B0(n626), .B1(n164), .C0(n986), .Y(
        n724) );
  AOI22X1 U468 ( .A0(din[215]), .A1(n178), .B0(dout[183]), .B1(n160), .Y(n986)
         );
  OAI221XL U469 ( .A0(n166), .A1(n231), .B0(n623), .B1(n163), .C0(n985), .Y(
        n723) );
  AOI22X1 U470 ( .A0(din[216]), .A1(n181), .B0(dout[184]), .B1(n150), .Y(n985)
         );
  OAI221XL U471 ( .A0(n167), .A1(n225), .B0(n321), .B1(n164), .C0(n984), .Y(
        n722) );
  AOI22X1 U472 ( .A0(din[217]), .A1(n181), .B0(dout[185]), .B1(n190), .Y(n984)
         );
  OAI221XL U473 ( .A0(n166), .A1(n219), .B0(n315), .B1(n163), .C0(n983), .Y(
        n721) );
  AOI22X1 U474 ( .A0(din[218]), .A1(n179), .B0(dout[186]), .B1(n160), .Y(n983)
         );
  OAI221XL U475 ( .A0(n169), .A1(n213), .B0(n309), .B1(n163), .C0(n982), .Y(
        n720) );
  AOI22X1 U476 ( .A0(din[219]), .A1(n179), .B0(dout[187]), .B1(n150), .Y(n982)
         );
  OAI221XL U477 ( .A0(n166), .A1(n207), .B0(n303), .B1(n163), .C0(n981), .Y(
        n719) );
  AOI22X1 U478 ( .A0(din[220]), .A1(n176), .B0(dout[188]), .B1(n151), .Y(n981)
         );
  OAI221XL U479 ( .A0(n167), .A1(n201), .B0(n297), .B1(n161), .C0(n980), .Y(
        n718) );
  AOI22X1 U480 ( .A0(din[221]), .A1(n178), .B0(dout[189]), .B1(n152), .Y(n980)
         );
  OAI221XL U481 ( .A0(n169), .A1(n196), .B0(n276), .B1(n164), .C0(n979), .Y(
        n717) );
  AOI22X1 U482 ( .A0(din[222]), .A1(n176), .B0(dout[190]), .B1(n160), .Y(n979)
         );
  OAI221XL U483 ( .A0(n166), .A1(n191), .B0(n271), .B1(n163), .C0(n978), .Y(
        n716) );
  AOI22X1 U484 ( .A0(din[223]), .A1(n178), .B0(dout[191]), .B1(n160), .Y(n978)
         );
  OAI221XL U485 ( .A0(n649), .A1(n166), .B0(n270), .B1(n161), .C0(n977), .Y(
        n715) );
  AOI22X1 U486 ( .A0(din[48]), .A1(n176), .B0(dout[192]), .B1(n152), .Y(n977)
         );
  INVX1 U487 ( .A(start), .Y(n190) );
  INVX1 U488 ( .A(mode[1]), .Y(n908) );
  NOR2X1 U489 ( .A(n908), .B(mode[0]), .Y(n929) );
  INVX1 U490 ( .A(n1170), .Y(n907) );
  AOI22X1 U491 ( .A0(din[0]), .A1(n187), .B0(dout[0]), .B1(n150), .Y(n1170) );
  INVX1 U492 ( .A(n1169), .Y(n906) );
  AOI22X1 U493 ( .A0(din[1]), .A1(n187), .B0(dout[1]), .B1(n150), .Y(n1169) );
  INVX1 U494 ( .A(n1168), .Y(n905) );
  AOI22X1 U495 ( .A0(din[2]), .A1(n187), .B0(dout[2]), .B1(n154), .Y(n1168) );
  INVX1 U496 ( .A(n1167), .Y(n904) );
  AOI22X1 U497 ( .A0(din[3]), .A1(n187), .B0(dout[3]), .B1(n154), .Y(n1167) );
  INVX1 U498 ( .A(n1166), .Y(n903) );
  AOI22X1 U499 ( .A0(din[4]), .A1(n187), .B0(dout[4]), .B1(n154), .Y(n1166) );
  INVX1 U500 ( .A(n1165), .Y(n902) );
  AOI22X1 U501 ( .A0(din[5]), .A1(n187), .B0(dout[5]), .B1(n154), .Y(n1165) );
  INVX1 U502 ( .A(n1164), .Y(n901) );
  AOI22X1 U503 ( .A0(din[6]), .A1(n187), .B0(dout[6]), .B1(n154), .Y(n1164) );
  INVX1 U504 ( .A(n1163), .Y(n900) );
  AOI22X1 U505 ( .A0(din[7]), .A1(n187), .B0(dout[7]), .B1(n154), .Y(n1163) );
  INVX1 U506 ( .A(n1162), .Y(n899) );
  AOI22X1 U507 ( .A0(din[8]), .A1(n187), .B0(dout[8]), .B1(n154), .Y(n1162) );
  INVX1 U508 ( .A(n1161), .Y(n898) );
  AOI22X1 U509 ( .A0(din[9]), .A1(n187), .B0(dout[9]), .B1(n150), .Y(n1161) );
  INVX1 U510 ( .A(n1160), .Y(n897) );
  AOI22X1 U511 ( .A0(din[10]), .A1(n187), .B0(dout[10]), .B1(n154), .Y(n1160)
         );
  INVX1 U512 ( .A(n1159), .Y(n896) );
  AOI22X1 U513 ( .A0(din[11]), .A1(n187), .B0(dout[11]), .B1(n160), .Y(n1159)
         );
  INVX1 U514 ( .A(n1158), .Y(n895) );
  AOI22X1 U515 ( .A0(din[12]), .A1(n187), .B0(dout[12]), .B1(n151), .Y(n1158)
         );
  INVX1 U516 ( .A(n1157), .Y(n894) );
  AOI22X1 U517 ( .A0(din[13]), .A1(N275), .B0(dout[13]), .B1(n150), .Y(n1157)
         );
  INVX1 U518 ( .A(n1156), .Y(n893) );
  AOI22X1 U519 ( .A0(din[14]), .A1(N275), .B0(dout[14]), .B1(n152), .Y(n1156)
         );
  INVX1 U520 ( .A(n1155), .Y(n892) );
  AOI22X1 U521 ( .A0(din[15]), .A1(N275), .B0(dout[15]), .B1(n152), .Y(n1155)
         );
  INVX1 U522 ( .A(n926), .Y(n667) );
  AOI22X1 U523 ( .A0(din[240]), .A1(N275), .B0(dout[240]), .B1(n151), .Y(n926)
         );
  INVX1 U524 ( .A(n925), .Y(n666) );
  AOI22X1 U525 ( .A0(din[241]), .A1(N275), .B0(dout[241]), .B1(n151), .Y(n925)
         );
  INVX1 U526 ( .A(n924), .Y(n665) );
  AOI22X1 U527 ( .A0(din[242]), .A1(N275), .B0(dout[242]), .B1(n152), .Y(n924)
         );
  INVX1 U528 ( .A(n923), .Y(n664) );
  AOI22X1 U529 ( .A0(din[243]), .A1(N275), .B0(dout[243]), .B1(n190), .Y(n923)
         );
  INVX1 U530 ( .A(n922), .Y(n663) );
  AOI22X1 U531 ( .A0(din[244]), .A1(N275), .B0(dout[244]), .B1(n151), .Y(n922)
         );
  INVX1 U532 ( .A(n921), .Y(n662) );
  AOI22X1 U533 ( .A0(din[245]), .A1(N275), .B0(dout[245]), .B1(n190), .Y(n921)
         );
  INVX1 U534 ( .A(n920), .Y(n661) );
  AOI22X1 U535 ( .A0(din[246]), .A1(N275), .B0(dout[246]), .B1(n150), .Y(n920)
         );
  INVX1 U536 ( .A(n919), .Y(n660) );
  AOI22X1 U537 ( .A0(din[247]), .A1(N275), .B0(dout[247]), .B1(n152), .Y(n919)
         );
  INVX1 U538 ( .A(n918), .Y(n659) );
  AOI22X1 U539 ( .A0(din[248]), .A1(N275), .B0(dout[248]), .B1(n151), .Y(n918)
         );
  INVX1 U540 ( .A(n917), .Y(n658) );
  AOI22X1 U541 ( .A0(din[249]), .A1(N275), .B0(dout[249]), .B1(n152), .Y(n917)
         );
  INVX1 U542 ( .A(n916), .Y(n657) );
  AOI22X1 U543 ( .A0(din[250]), .A1(n187), .B0(dout[250]), .B1(n190), .Y(n916)
         );
  INVX1 U544 ( .A(n915), .Y(n656) );
  AOI22X1 U545 ( .A0(din[251]), .A1(n187), .B0(dout[251]), .B1(n150), .Y(n915)
         );
  INVX1 U546 ( .A(n914), .Y(n655) );
  AOI22X1 U547 ( .A0(din[252]), .A1(N275), .B0(dout[252]), .B1(n160), .Y(n914)
         );
  INVX1 U548 ( .A(n913), .Y(n654) );
  AOI22X1 U549 ( .A0(din[253]), .A1(N275), .B0(dout[253]), .B1(n160), .Y(n913)
         );
  INVX1 U550 ( .A(n912), .Y(n653) );
  AOI22X1 U551 ( .A0(din[254]), .A1(N275), .B0(dout[254]), .B1(n190), .Y(n912)
         );
  INVX1 U552 ( .A(n911), .Y(n652) );
  AOI22X1 U553 ( .A0(din[255]), .A1(N275), .B0(dout[255]), .B1(n151), .Y(n911)
         );
  OAI21XL U554 ( .A0(n910), .A1(n908), .B0(start), .Y(n909) );
  OAI2BB2X1 U555 ( .B0(n910), .B1(n909), .A0N(mode_out[0]), .A1N(n909), .Y(
        n651) );
  OAI2BB2X1 U556 ( .B0(n908), .B1(n909), .A0N(mode_out[1]), .A1N(n909), .Y(
        n650) );
  INVX1 U557 ( .A(din[144]), .Y(n270) );
  INVX1 U558 ( .A(din[145]), .Y(n265) );
  INVX1 U559 ( .A(din[146]), .Y(n261) );
  INVX1 U560 ( .A(din[147]), .Y(n256) );
  INVX1 U561 ( .A(din[148]), .Y(n252) );
  INVX1 U562 ( .A(din[149]), .Y(n247) );
  INVX1 U563 ( .A(din[150]), .Y(n243) );
  INVX1 U564 ( .A(din[151]), .Y(n238) );
  INVX1 U565 ( .A(din[152]), .Y(n234) );
  INVX1 U566 ( .A(din[153]), .Y(n229) );
  INVX1 U567 ( .A(din[154]), .Y(n223) );
  INVX1 U568 ( .A(din[155]), .Y(n217) );
  INVX1 U569 ( .A(din[156]), .Y(n211) );
  INVX1 U570 ( .A(din[157]), .Y(n205) );
  INVX1 U571 ( .A(din[158]), .Y(n199) );
  INVX1 U572 ( .A(din[159]), .Y(n194) );
  INVX1 U573 ( .A(din[176]), .Y(n267) );
  INVX1 U574 ( .A(din[177]), .Y(n262) );
  INVX1 U575 ( .A(din[178]), .Y(n258) );
  INVX1 U576 ( .A(din[179]), .Y(n253) );
  INVX1 U577 ( .A(din[180]), .Y(n249) );
  INVX1 U578 ( .A(din[181]), .Y(n244) );
  INVX1 U579 ( .A(din[182]), .Y(n240) );
  INVX1 U580 ( .A(din[183]), .Y(n235) );
  INVX1 U581 ( .A(din[184]), .Y(n231) );
  INVX1 U582 ( .A(din[185]), .Y(n225) );
  INVX1 U583 ( .A(din[186]), .Y(n219) );
  INVX1 U584 ( .A(din[187]), .Y(n213) );
  INVX1 U585 ( .A(din[188]), .Y(n207) );
  INVX1 U586 ( .A(din[189]), .Y(n201) );
  INVX1 U587 ( .A(din[190]), .Y(n196) );
  INVX1 U588 ( .A(din[191]), .Y(n191) );
  INVX1 U589 ( .A(din[208]), .Y(n648) );
  INVX1 U590 ( .A(din[209]), .Y(n645) );
  INVX1 U591 ( .A(din[210]), .Y(n642) );
  INVX1 U592 ( .A(din[211]), .Y(n639) );
  INVX1 U593 ( .A(din[212]), .Y(n636) );
  INVX1 U594 ( .A(din[213]), .Y(n633) );
  INVX1 U595 ( .A(din[214]), .Y(n630) );
  INVX1 U596 ( .A(din[215]), .Y(n627) );
  INVX1 U597 ( .A(din[216]), .Y(n624) );
  INVX1 U598 ( .A(din[217]), .Y(n323) );
  INVX1 U599 ( .A(din[218]), .Y(n317) );
  INVX1 U600 ( .A(din[219]), .Y(n311) );
  INVX1 U601 ( .A(din[220]), .Y(n305) );
  INVX1 U602 ( .A(din[221]), .Y(n299) );
  INVX1 U603 ( .A(din[222]), .Y(n277) );
  INVX1 U604 ( .A(din[223]), .Y(n273) );
  INVX1 U605 ( .A(din[160]), .Y(n268) );
  INVX1 U606 ( .A(din[161]), .Y(n264) );
  INVX1 U607 ( .A(din[162]), .Y(n259) );
  INVX1 U608 ( .A(din[163]), .Y(n255) );
  INVX1 U609 ( .A(din[164]), .Y(n250) );
  INVX1 U610 ( .A(din[165]), .Y(n246) );
  INVX1 U611 ( .A(din[166]), .Y(n241) );
  INVX1 U612 ( .A(din[167]), .Y(n237) );
  INVX1 U613 ( .A(din[168]), .Y(n232) );
  INVX1 U614 ( .A(din[169]), .Y(n227) );
  INVX1 U615 ( .A(din[170]), .Y(n221) );
  INVX1 U616 ( .A(din[171]), .Y(n215) );
  INVX1 U617 ( .A(din[172]), .Y(n209) );
  INVX1 U618 ( .A(din[173]), .Y(n203) );
  INVX1 U619 ( .A(din[174]), .Y(n197) );
  INVX1 U620 ( .A(din[175]), .Y(n193) );
  INVX1 U621 ( .A(din[192]), .Y(n649) );
  INVX1 U622 ( .A(din[193]), .Y(n646) );
  INVX1 U623 ( .A(din[194]), .Y(n643) );
  INVX1 U624 ( .A(din[195]), .Y(n640) );
  INVX1 U625 ( .A(din[196]), .Y(n637) );
  INVX1 U626 ( .A(din[197]), .Y(n634) );
  INVX1 U627 ( .A(din[198]), .Y(n631) );
  INVX1 U628 ( .A(din[199]), .Y(n628) );
  INVX1 U629 ( .A(din[200]), .Y(n625) );
  INVX1 U630 ( .A(din[201]), .Y(n325) );
  INVX1 U631 ( .A(din[202]), .Y(n319) );
  INVX1 U632 ( .A(din[203]), .Y(n313) );
  INVX1 U633 ( .A(din[204]), .Y(n307) );
  INVX1 U634 ( .A(din[205]), .Y(n301) );
  INVX1 U635 ( .A(din[206]), .Y(n295) );
  INVX1 U636 ( .A(din[207]), .Y(n274) );
  INVX1 U637 ( .A(din[224]), .Y(n647) );
  INVX1 U638 ( .A(din[225]), .Y(n644) );
  INVX1 U639 ( .A(din[226]), .Y(n641) );
  INVX1 U640 ( .A(din[227]), .Y(n638) );
  INVX1 U641 ( .A(din[228]), .Y(n635) );
  INVX1 U642 ( .A(din[229]), .Y(n632) );
  INVX1 U643 ( .A(din[230]), .Y(n629) );
  INVX1 U644 ( .A(din[231]), .Y(n626) );
  INVX1 U645 ( .A(din[232]), .Y(n623) );
  INVX1 U646 ( .A(din[233]), .Y(n321) );
  INVX1 U647 ( .A(din[234]), .Y(n315) );
  INVX1 U648 ( .A(din[235]), .Y(n309) );
  INVX1 U649 ( .A(din[236]), .Y(n303) );
  INVX1 U650 ( .A(din[237]), .Y(n297) );
  INVX1 U651 ( .A(din[238]), .Y(n276) );
  INVX1 U652 ( .A(din[239]), .Y(n271) );
endmodule


module idct4_shift12_add2048_DW01_add_4 ( A, B, SUM );
  input [24:0] A;
  input [24:0] B;
  output [24:0] SUM;
  wire   n2;
  wire   [24:1] carry;

  XOR3X2 U1_24 ( .A(A[24]), .B(B[24]), .C(carry[24]), .Y(SUM[24]) );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_5 ( .A(1'b0), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(1'b0), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(1'b0), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(1'b0), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_1 ( .A(1'b0), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  CLKINVX8 U1 ( .A(n2), .Y(carry[1]) );
  CLKINVX8 U2 ( .A(B[0]), .Y(SUM[0]) );
  INVX1 U4 ( .A(B[0]), .Y(n2) );
endmodule


module idct4_shift12_add2048_DW01_add_5 ( A, B, SUM );
  input [24:0] A;
  input [24:0] B;
  output [24:0] SUM;
  wire   n2;
  wire   [24:1] carry;

  XOR3X2 U1_24 ( .A(A[24]), .B(B[24]), .C(carry[24]), .Y(SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(1'b0), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(1'b0), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(1'b0), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(1'b0), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_1 ( .A(1'b0), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  CLKINVX8 U1 ( .A(n2), .Y(carry[1]) );
  CLKINVX8 U2 ( .A(B[0]), .Y(SUM[0]) );
  INVX1 U4 ( .A(B[0]), .Y(n2) );
endmodule


module idct4_shift12_add2048_DW01_add_6 ( A, B, SUM );
  input [24:0] A;
  input [24:0] B;
  output [24:0] SUM;

  wire   [24:1] carry;

  XOR3X2 U1_24 ( .A(A[24]), .B(B[24]), .C(carry[24]), .Y(SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_1 ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(SUM[1]) );
  ADDFX2 U1_5 ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(SUM[5]) );
  ADDFX2 U1_4 ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(SUM[4]) );
  ADDFX2 U1_3 ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(SUM[3]) );
  ADDFX2 U1_2 ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(SUM[2]) );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(1'b0), .CO(carry[7]), .S(SUM[6]) );
  XOR2X1 U1 ( .A(B[0]), .B(1'b0), .Y(SUM[0]) );
endmodule


module idct4_shift12_add2048_DW01_add_7 ( A, B, SUM );
  input [24:0] A;
  input [24:0] B;
  output [24:0] SUM;

  wire   [24:1] carry;

  XOR3X2 U1_24 ( .A(A[24]), .B(B[24]), .C(carry[24]), .Y(SUM[24]) );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_1 ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(SUM[1]) );
  ADDFX2 U1_5 ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(SUM[5]) );
  ADDFX2 U1_4 ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(SUM[4]) );
  ADDFX2 U1_3 ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(SUM[3]) );
  ADDFX2 U1_2 ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(SUM[2]) );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(1'b0), .CO(carry[7]), .S(SUM[6]) );
  XOR2X1 U1 ( .A(B[0]), .B(1'b0), .Y(SUM[0]) );
endmodule


module idct4_shift12_add2048_DW01_add_8 ( A, B, SUM );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;

  wire   [23:1] carry;

  XOR3X2 U1_23 ( .A(A[23]), .B(B[23]), .C(carry[23]), .Y(SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_1 ( .A(A[1]), .B(1'b0), .CI(1'b0), .S(SUM[1]) );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(1'b0), .CO(carry[3]), .S(SUM[2]) );
  XOR2X1 U1 ( .A(1'b0), .B(A[0]), .Y(SUM[0]) );
endmodule


module idct4_shift12_add2048_DW01_add_9 ( A, B, SUM );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  wire   n2;
  wire   [23:1] carry;

  XOR3X2 U1_23 ( .A(A[23]), .B(B[23]), .C(carry[23]), .Y(SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_1 ( .A(1'b0), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  CLKINVX8 U1 ( .A(n2), .Y(carry[1]) );
  CLKINVX8 U2 ( .A(B[0]), .Y(SUM[0]) );
  INVX1 U4 ( .A(B[0]), .Y(n2) );
endmodule


module idct4_shift12_add2048_DW01_add_12 ( A, B, SUM );
  input [22:0] A;
  input [22:0] B;
  output [22:0] SUM;

  wire   [22:1] carry;

  XOR3X2 U1_22 ( .A(A[22]), .B(B[22]), .C(carry[22]), .Y(SUM[22]) );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(1'b0), .CO(carry[2]), .S(SUM[1]) );
  XOR2X1 U1 ( .A(1'b0), .B(A[0]), .Y(SUM[0]) );
endmodule


module idct4_shift12_add2048_DW01_add_13 ( A, B, SUM );
  input [22:0] A;
  input [22:0] B;
  output [22:0] SUM;

  wire   [22:1] carry;

  XOR3X2 U1_22 ( .A(A[22]), .B(B[22]), .C(carry[22]), .Y(SUM[22]) );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(1'b0), .CO(carry[2]), .S(SUM[1]) );
  XOR2X1 U1 ( .A(1'b0), .B(A[0]), .Y(SUM[0]) );
endmodule


module idct4_shift12_add2048 ( clk, rstn, mode, start, x0, x1, x2, x3, y0, y1, 
        y2, y3, idct4_ready );
  input [1:0] mode;
  input [15:0] x0;
  input [15:0] x1;
  input [15:0] x2;
  input [15:0] x3;
  output [24:0] y0;
  output [24:0] y1;
  output [24:0] y2;
  output [24:0] y3;
  input clk, rstn, start;
  output idct4_ready;
  wire   idct4_ready_delay1, idct4_ready_delay2, idct4_ready_delay3, N14, N15,
         N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29,
         N30, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48,
         N49, N50, N51, N52, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68,
         N69, N70, N71, N72, N73, N74, N80, N81, N82, N83, N84, N85, N86, N87,
         N88, N89, N90, N91, N92, N93, N94, N95, N103, N104, N105, N106, N107,
         N108, N109, N110, N111, N112, N113, N114, N115, N116, N117, N118,
         N124, N125, N126, N127, N128, N129, N130, N131, N132, N133, N134,
         N135, N136, N137, N138, N139, N141, N142, N143, N144, N145, N146,
         N147, N148, N149, N150, N151, N152, N153, N154, N155, N156, N157,
         N158, N159, N160, N161, N162, N163, N164, N165, N166, N167, N168,
         N169, N170, N171, N172, N173, N174, N175, N176, N177, N178, N179,
         N180, N181, N182, N183, N184, N185, N186, N193, N194, N195, N196,
         N197, N198, N199, N200, N201, N202, N203, N204, N205, N206, N207,
         N208, N209, N261, N262, N263, N264, N265, N266, N267, N268, N269,
         N270, N271, N272, N273, N274, N275, N276, N277, N325, N326, N327,
         N328, N329, N330, N331, N332, N333, N334, N335, N336, N337, N338,
         N339, N340, N341, N342, N343, N344, N345, N346, N347, N348, N349,
         N350, N351, N352, N353, N354, N355, N356, N357, N358, N359, N360,
         N361, N362, N363, N364, N365, N366, N367, N368, N369, N370, N371,
         N372, N373, N374, N375, N376, N377, N378, N379, N380, N381, N382,
         N383, N384, N385, N386, N387, N388, N389, N390, N391, N392, N393,
         N394, N395, N396, N397, N398, N399, N400, N401, N402, N403, N404,
         N405, N406, N407, N408, N409, N410, N411, N412, N413, N414, N415,
         N416, N417, N418, N419, N420, N421, N422, N472, N473, N474, N475,
         N476, N477, N478, N479, N480, N481, N482, N483, N484, N485, N486,
         N487, N488, N489, N490, N491, N492, N493, N494, N495, N496, N546,
         N547, N548, N549, N550, N551, N552, N553, N554, N555, N556, N557,
         N558, N559, N560, N561, N562, N563, N564, N565, N566, N567, N568,
         N569, N570, N571, N572, N573, N574, N575, N576, N577, N578, N579,
         N580, N581, N582, N583, N584, N585, N586, N587, N588, N589, N590,
         N591, N592, N593, N594, N595, N596, N597, N598, N599, N600, N601,
         N602, N603, N604, N605, N606, N607, N608, N609, N610, N611, N612,
         N613, N614, N615, N616, N617, N618, N619, N620, N621, N622, N623,
         N624, N625, N626, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, add_125_carry_13_, add_125_carry_14_,
         add_125_carry_15_, add_125_carry_16_, add_125_carry_17_,
         add_125_carry_18_, add_125_carry_19_, add_125_carry_20_,
         add_125_carry_21_, add_125_carry_22_, add_125_carry_23_,
         add_125_carry_24_, add_125_carry_25_, add_124_carry_13_,
         add_124_carry_14_, add_124_carry_15_, add_124_carry_16_,
         add_124_carry_17_, add_124_carry_18_, add_124_carry_19_,
         add_124_carry_20_, add_124_carry_21_, add_124_carry_22_,
         add_124_carry_23_, add_124_carry_24_, add_124_carry_25_,
         add_123_carry_13_, add_123_carry_14_, add_123_carry_15_,
         add_123_carry_16_, add_123_carry_17_, add_123_carry_18_,
         add_123_carry_19_, add_123_carry_20_, add_123_carry_21_,
         add_123_carry_22_, add_123_carry_23_, add_123_carry_24_,
         add_123_carry_25_, add_122_carry_13_, add_122_carry_14_,
         add_122_carry_15_, add_122_carry_16_, add_122_carry_17_,
         add_122_carry_18_, add_122_carry_19_, add_122_carry_20_,
         add_122_carry_21_, add_122_carry_22_, add_122_carry_23_,
         add_122_carry_24_, add_122_carry_25_, add_1_root_add_112_2_B_6_,
         add_1_root_add_112_2_B_7_, add_1_root_add_112_2_B_8_,
         add_1_root_add_112_2_B_9_, add_1_root_add_112_2_B_10_,
         add_1_root_add_112_2_B_11_, add_1_root_add_112_2_B_12_,
         add_1_root_add_112_2_B_13_, add_1_root_add_112_2_B_14_,
         add_1_root_add_112_2_B_15_, add_1_root_add_112_2_B_16_,
         add_1_root_add_112_2_B_17_, add_1_root_add_112_2_B_18_,
         add_1_root_add_112_2_B_19_, add_1_root_add_112_2_B_20_,
         add_1_root_add_112_2_B_21_, add_88_carry_10_, add_88_carry_11_,
         add_88_carry_12_, add_88_carry_13_, add_88_carry_14_,
         add_88_carry_15_, add_88_carry_16_, add_88_carry_17_,
         add_88_carry_18_, add_88_carry_5_, add_88_carry_6_, add_88_carry_7_,
         add_88_carry_8_, add_88_carry_9_, add_87_carry_10_, add_87_carry_11_,
         add_87_carry_12_, add_87_carry_13_, add_87_carry_14_,
         add_87_carry_15_, add_87_carry_16_, add_87_carry_17_,
         add_87_carry_18_, add_87_carry_19_, add_87_carry_20_, add_87_carry_7_,
         add_87_carry_8_, add_87_carry_9_, add_86_carry_10_, add_86_carry_11_,
         add_86_carry_12_, add_86_carry_13_, add_86_carry_14_,
         add_86_carry_15_, add_86_carry_16_, add_86_carry_17_,
         add_86_carry_18_, add_86_carry_5_, add_86_carry_6_, add_86_carry_7_,
         add_86_carry_8_, add_86_carry_9_, add_85_carry_10_, add_85_carry_11_,
         add_85_carry_12_, add_85_carry_13_, add_85_carry_14_,
         add_85_carry_15_, add_85_carry_16_, add_85_carry_17_,
         add_85_carry_18_, add_85_carry_19_, add_85_carry_20_, add_85_carry_7_,
         add_85_carry_8_, add_85_carry_9_, add_81_carry_10_, add_81_carry_11_,
         add_81_carry_12_, add_81_carry_13_, add_81_carry_14_,
         add_81_carry_15_, add_81_carry_16_, add_81_carry_17_,
         add_81_carry_18_, add_81_carry_19_, add_81_carry_6_, add_81_carry_7_,
         add_81_carry_8_, add_81_carry_9_, add_80_carry_10_, add_80_carry_11_,
         add_80_carry_12_, add_80_carry_13_, add_80_carry_14_,
         add_80_carry_15_, add_80_carry_16_, add_80_carry_17_,
         add_80_carry_18_, add_80_carry_19_, add_80_carry_6_, add_80_carry_7_,
         add_80_carry_8_, add_80_carry_9_, n1, n2, n3, n4, n8, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108;
  wire   [1:0] mode_delay2;
  wire   [1:0] mode_delay1;
  wire   [20:0] x1_o0_tmp2;
  wire   [20:0] x3_o1_tmp2;
  wire   [21:6] x0_e;
  wire   [21:6] x2_e;
  wire   [21:0] x1_o1;
  wire   [21:0] x3_o0;
  wire   [22:0] x1_o0;
  wire   [22:0] x3_o1;
  wire   [21:2] x3_o0_tmp;
  wire   [21:2] x1_o1_tmp;
  wire   [21:6] x2_e_tmp;
  wire   [21:6] x0_e_tmp;
  wire   [22:0] x3_o1_tmp1;
  wire   [22:0] x1_o0_tmp1;
  wire   [22:0] e0;
  wire   [23:0] o0;
  wire   [22:0] e1;
  wire   [23:0] o1;
  wire   [24:0] y0_tmp;
  wire   [24:0] y1_tmp;
  wire   [24:0] y2_tmp;
  wire   [24:0] y3_tmp;
  wire   [22:7] add_1_root_add_112_2_carry;
  wire   [22:7] add_111_carry;

  idct4_shift12_add2048_DW01_add_4 add_1_root_add_119_2 ( .A({e0[22], e0[22], 
        e0[22:6], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({n85, n85, n86, n87, 
        n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, 
        n102, n103, n104, n105, n106, n107, n108}), .SUM({N570, N569, N568, 
        N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, 
        N555, N554, N553, N552, N551, N550, N549, N548, N547, N546}) );
  idct4_shift12_add2048_DW01_add_5 add_1_root_add_118_2 ( .A({e1[22], e1[22], 
        e1[22:6], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({n61, n61, n62, n63, 
        n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
        n78, n79, n80, n81, n82, n83, n84}), .SUM({N496, N495, N494, N493, 
        N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, 
        N480, N479, N478, N477, N476, N475, N474, N473, N472}) );
  idct4_shift12_add2048_DW01_add_6 add_117 ( .A({e1[22], e1[22], e1[22:6], 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({o1[23], o1}), .SUM({N422, 
        N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, 
        N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398}) );
  idct4_shift12_add2048_DW01_add_7 add_116 ( .A({e0[22], e0[22], e0[22:6], 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({o0[23], o0}), .SUM({N397, 
        N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, 
        N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373}) );
  idct4_shift12_add2048_DW01_add_8 add_114 ( .A({x1_o0[22], x1_o0}), .B({
        x3_o0[21], x3_o0[21], x3_o0[21:2], 1'b0, 1'b0}), .SUM({N372, N371, 
        N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, 
        N358, N357, N356, N355, N354, N353, N352, N351, N350, N349}) );
  idct4_shift12_add2048_DW01_add_9 add_1_root_add_113_2 ( .A({x1_o1[21], 
        x1_o1[21], x1_o1[21:2], 1'b0, 1'b0}), .B({n38, n38, n39, n40, n41, n42, 
        n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, 
        n57, n58, n59, n60}), .SUM({N348, N347, N346, N345, N344, N343, N342, 
        N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, 
        N329, N328, N327, N326, N325}) );
  idct4_shift12_add2048_DW01_add_12 add_90 ( .A(x3_o1_tmp1), .B({
        x3_o1_tmp2[20], x3_o1_tmp2[20], x3_o1_tmp2[20:1], 1'b0}), .SUM({N186, 
        N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, 
        N173, N172, N171, N170, N169, N168, N167, N166, N165, N164}) );
  idct4_shift12_add2048_DW01_add_13 add_89 ( .A(x1_o0_tmp1), .B({
        x1_o0_tmp2[20], x1_o0_tmp2[20], x1_o0_tmp2[20:1], 1'b0}), .SUM({N163, 
        N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, 
        N150, N149, N148, N147, N146, N145, N144, N143, N142, N141}) );
  DFFRHQX1 x3_o1_tmp1_reg_22_ ( .D(N52), .CK(clk), .RN(rstn), .Q(
        x3_o1_tmp1[22]) );
  DFFRHQX1 x3_o1_tmp1_reg_21_ ( .D(N118), .CK(clk), .RN(rstn), .Q(
        x3_o1_tmp1[21]) );
  DFFRHQX1 x3_o1_tmp1_reg_20_ ( .D(N117), .CK(clk), .RN(rstn), .Q(
        x3_o1_tmp1[20]) );
  DFFRHQX1 x3_o1_tmp1_reg_19_ ( .D(N116), .CK(clk), .RN(rstn), .Q(
        x3_o1_tmp1[19]) );
  DFFRHQX1 x1_o0_tmp1_reg_22_ ( .D(N30), .CK(clk), .RN(rstn), .Q(
        x1_o0_tmp1[22]) );
  DFFRHQX1 x1_o0_tmp1_reg_21_ ( .D(N74), .CK(clk), .RN(rstn), .Q(
        x1_o0_tmp1[21]) );
  DFFRHQX1 x1_o0_tmp1_reg_20_ ( .D(N73), .CK(clk), .RN(rstn), .Q(
        x1_o0_tmp1[20]) );
  DFFRHQX1 x1_o0_tmp1_reg_19_ ( .D(N72), .CK(clk), .RN(rstn), .Q(
        x1_o0_tmp1[19]) );
  DFFRHQX1 x1_o0_reg_20_ ( .D(N161), .CK(clk), .RN(rstn), .Q(x1_o0[20]) );
  DFFRHQX1 x1_o0_reg_21_ ( .D(N162), .CK(clk), .RN(rstn), .Q(x1_o0[21]) );
  DFFRHQX1 x1_o1_reg_20_ ( .D(x1_o1_tmp[20]), .CK(clk), .RN(rstn), .Q(
        x1_o1[20]) );
  DFFRHQX1 x3_o1_reg_22_ ( .D(N186), .CK(clk), .RN(rstn), .Q(x3_o1[22]) );
  DFFRHQX1 x3_o1_reg_21_ ( .D(N185), .CK(clk), .RN(rstn), .Q(x3_o1[21]) );
  DFFRHQX1 x3_o1_reg_20_ ( .D(N184), .CK(clk), .RN(rstn), .Q(x3_o1[20]) );
  DFFRHQX1 x1_o0_reg_22_ ( .D(N163), .CK(clk), .RN(rstn), .Q(x1_o0[22]) );
  DFFRHQX1 x0_e_reg_20_ ( .D(x0_e_tmp[20]), .CK(clk), .RN(rstn), .Q(x0_e[20])
         );
  DFFRHQX1 x0_e_reg_19_ ( .D(x0_e_tmp[19]), .CK(clk), .RN(rstn), .Q(x0_e[19])
         );
  DFFRHQX1 e1_reg_21_ ( .D(N276), .CK(clk), .RN(rstn), .Q(e1[21]) );
  DFFRHQX1 e0_reg_21_ ( .D(N208), .CK(clk), .RN(rstn), .Q(e0[21]) );
  DFFRHQX1 x3_o1_tmp2_reg_19_ ( .D(N139), .CK(clk), .RN(rstn), .Q(
        x3_o1_tmp2[19]) );
  DFFRHQX1 x1_o0_tmp2_reg_19_ ( .D(N95), .CK(clk), .RN(rstn), .Q(
        x1_o0_tmp2[19]) );
  DFFRHQX1 x3_o0_reg_20_ ( .D(x3_o0_tmp[20]), .CK(clk), .RN(rstn), .Q(
        x3_o0[20]) );
  DFFRHQX1 x3_o1_tmp1_reg_0_ ( .D(x3[0]), .CK(clk), .RN(rstn), .Q(
        x3_o1_tmp1[0]) );
  DFFRHQX1 x1_o0_tmp1_reg_0_ ( .D(x1[0]), .CK(clk), .RN(rstn), .Q(
        x1_o0_tmp1[0]) );
  DFFRHQX1 x1_o0_reg_0_ ( .D(N141), .CK(clk), .RN(rstn), .Q(x1_o0[0]) );
  DFFRHQX1 x1_o1_reg_21_ ( .D(x1_o1_tmp[21]), .CK(clk), .RN(rstn), .Q(
        x1_o1[21]) );
  DFFRHQX1 x0_e_reg_21_ ( .D(x0_e_tmp[21]), .CK(clk), .RN(rstn), .Q(x0_e[21])
         );
  DFFRHQX1 x2_e_reg_20_ ( .D(x2_e_tmp[20]), .CK(clk), .RN(rstn), .Q(x2_e[20])
         );
  DFFRHQX1 o1_reg_22_ ( .D(N347), .CK(clk), .RN(rstn), .Q(o1[22]) );
  DFFRHQX1 o0_reg_22_ ( .D(N371), .CK(clk), .RN(rstn), .Q(o0[22]) );
  DFFRHQX1 e1_reg_22_ ( .D(N277), .CK(clk), .RN(rstn), .Q(e1[22]) );
  DFFRHQX1 e0_reg_22_ ( .D(N209), .CK(clk), .RN(rstn), .Q(e0[22]) );
  DFFRHQX1 x2_e_reg_21_ ( .D(x2_e_tmp[21]), .CK(clk), .RN(rstn), .Q(x2_e[21])
         );
  DFFRHQX1 o1_reg_23_ ( .D(N348), .CK(clk), .RN(rstn), .Q(o1[23]) );
  DFFRHQX1 o0_reg_23_ ( .D(N372), .CK(clk), .RN(rstn), .Q(o0[23]) );
  DFFRHQX1 x3_o1_tmp2_reg_20_ ( .D(N52), .CK(clk), .RN(rstn), .Q(
        x3_o1_tmp2[20]) );
  DFFRHQX1 x1_o0_tmp2_reg_20_ ( .D(N30), .CK(clk), .RN(rstn), .Q(
        x1_o0_tmp2[20]) );
  DFFRHQX1 x3_o0_reg_21_ ( .D(x3_o0_tmp[21]), .CK(clk), .RN(rstn), .Q(
        x3_o0[21]) );
  DFFRHQX1 x3_o1_tmp1_reg_18_ ( .D(N115), .CK(clk), .RN(rstn), .Q(
        x3_o1_tmp1[18]) );
  DFFRHQX1 x3_o1_tmp1_reg_17_ ( .D(N114), .CK(clk), .RN(rstn), .Q(
        x3_o1_tmp1[17]) );
  DFFRHQX1 x3_o1_tmp1_reg_16_ ( .D(N113), .CK(clk), .RN(rstn), .Q(
        x3_o1_tmp1[16]) );
  DFFRHQX1 x3_o1_tmp1_reg_15_ ( .D(N112), .CK(clk), .RN(rstn), .Q(
        x3_o1_tmp1[15]) );
  DFFRHQX1 x1_o0_tmp1_reg_18_ ( .D(N71), .CK(clk), .RN(rstn), .Q(
        x1_o0_tmp1[18]) );
  DFFRHQX1 x1_o0_tmp1_reg_17_ ( .D(N70), .CK(clk), .RN(rstn), .Q(
        x1_o0_tmp1[17]) );
  DFFRHQX1 x1_o0_tmp1_reg_16_ ( .D(N69), .CK(clk), .RN(rstn), .Q(
        x1_o0_tmp1[16]) );
  DFFRHQX1 x1_o0_tmp1_reg_15_ ( .D(N68), .CK(clk), .RN(rstn), .Q(
        x1_o0_tmp1[15]) );
  DFFRHQX1 x1_o0_reg_16_ ( .D(N157), .CK(clk), .RN(rstn), .Q(x1_o0[16]) );
  DFFRHQX1 x1_o0_reg_17_ ( .D(N158), .CK(clk), .RN(rstn), .Q(x1_o0[17]) );
  DFFRHQX1 x1_o0_reg_18_ ( .D(N159), .CK(clk), .RN(rstn), .Q(x1_o0[18]) );
  DFFRHQX1 x1_o0_reg_19_ ( .D(N160), .CK(clk), .RN(rstn), .Q(x1_o0[19]) );
  DFFRHQX1 x1_o1_reg_19_ ( .D(x1_o1_tmp[19]), .CK(clk), .RN(rstn), .Q(
        x1_o1[19]) );
  DFFRHQX1 x1_o1_reg_18_ ( .D(x1_o1_tmp[18]), .CK(clk), .RN(rstn), .Q(
        x1_o1[18]) );
  DFFRHQX1 x1_o1_reg_17_ ( .D(x1_o1_tmp[17]), .CK(clk), .RN(rstn), .Q(
        x1_o1[17]) );
  DFFRHQX1 x1_o1_reg_16_ ( .D(x1_o1_tmp[16]), .CK(clk), .RN(rstn), .Q(
        x1_o1[16]) );
  DFFRHQX1 x3_o1_reg_19_ ( .D(N183), .CK(clk), .RN(rstn), .Q(x3_o1[19]) );
  DFFRHQX1 x3_o1_reg_18_ ( .D(N182), .CK(clk), .RN(rstn), .Q(x3_o1[18]) );
  DFFRHQX1 x3_o1_reg_17_ ( .D(N181), .CK(clk), .RN(rstn), .Q(x3_o1[17]) );
  DFFRHQX1 x3_o1_reg_16_ ( .D(N180), .CK(clk), .RN(rstn), .Q(x3_o1[16]) );
  DFFRHQX1 x0_e_reg_18_ ( .D(x0_e_tmp[18]), .CK(clk), .RN(rstn), .Q(x0_e[18])
         );
  DFFRHQX1 x0_e_reg_17_ ( .D(x0_e_tmp[17]), .CK(clk), .RN(rstn), .Q(x0_e[17])
         );
  DFFRHQX1 x0_e_reg_16_ ( .D(x0_e_tmp[16]), .CK(clk), .RN(rstn), .Q(x0_e[16])
         );
  DFFRHQX1 x0_e_reg_15_ ( .D(x0_e_tmp[15]), .CK(clk), .RN(rstn), .Q(x0_e[15])
         );
  DFFRHQX1 e1_reg_20_ ( .D(N275), .CK(clk), .RN(rstn), .Q(e1[20]) );
  DFFRHQX1 e1_reg_19_ ( .D(N274), .CK(clk), .RN(rstn), .Q(e1[19]) );
  DFFRHQX1 e1_reg_18_ ( .D(N273), .CK(clk), .RN(rstn), .Q(e1[18]) );
  DFFRHQX1 e1_reg_17_ ( .D(N272), .CK(clk), .RN(rstn), .Q(e1[17]) );
  DFFRHQX1 e0_reg_20_ ( .D(N207), .CK(clk), .RN(rstn), .Q(e0[20]) );
  DFFRHQX1 e0_reg_19_ ( .D(N206), .CK(clk), .RN(rstn), .Q(e0[19]) );
  DFFRHQX1 e0_reg_18_ ( .D(N205), .CK(clk), .RN(rstn), .Q(e0[18]) );
  DFFRHQX1 e0_reg_17_ ( .D(N204), .CK(clk), .RN(rstn), .Q(e0[17]) );
  DFFRHQX1 x3_o1_tmp2_reg_18_ ( .D(N138), .CK(clk), .RN(rstn), .Q(
        x3_o1_tmp2[18]) );
  DFFRHQX1 x3_o1_tmp2_reg_17_ ( .D(N137), .CK(clk), .RN(rstn), .Q(
        x3_o1_tmp2[17]) );
  DFFRHQX1 x3_o1_tmp2_reg_16_ ( .D(N136), .CK(clk), .RN(rstn), .Q(
        x3_o1_tmp2[16]) );
  DFFRHQX1 x3_o1_tmp2_reg_15_ ( .D(N135), .CK(clk), .RN(rstn), .Q(
        x3_o1_tmp2[15]) );
  DFFRHQX1 x3_o1_tmp2_reg_14_ ( .D(N134), .CK(clk), .RN(rstn), .Q(
        x3_o1_tmp2[14]) );
  DFFRHQX1 x1_o0_tmp2_reg_18_ ( .D(N94), .CK(clk), .RN(rstn), .Q(
        x1_o0_tmp2[18]) );
  DFFRHQX1 x1_o0_tmp2_reg_17_ ( .D(N93), .CK(clk), .RN(rstn), .Q(
        x1_o0_tmp2[17]) );
  DFFRHQX1 x1_o0_tmp2_reg_16_ ( .D(N92), .CK(clk), .RN(rstn), .Q(
        x1_o0_tmp2[16]) );
  DFFRHQX1 x1_o0_tmp2_reg_15_ ( .D(N91), .CK(clk), .RN(rstn), .Q(
        x1_o0_tmp2[15]) );
  DFFRHQX1 x1_o0_tmp2_reg_14_ ( .D(N90), .CK(clk), .RN(rstn), .Q(
        x1_o0_tmp2[14]) );
  DFFRHQX1 x3_o0_reg_19_ ( .D(x3_o0_tmp[19]), .CK(clk), .RN(rstn), .Q(
        x3_o0[19]) );
  DFFRHQX1 x3_o0_reg_18_ ( .D(x3_o0_tmp[18]), .CK(clk), .RN(rstn), .Q(
        x3_o0[18]) );
  DFFRHQX1 x3_o0_reg_17_ ( .D(x3_o0_tmp[17]), .CK(clk), .RN(rstn), .Q(
        x3_o0[17]) );
  DFFRHQX1 x3_o0_reg_16_ ( .D(x3_o0_tmp[16]), .CK(clk), .RN(rstn), .Q(
        x3_o0[16]) );
  DFFRHQX1 x3_o0_reg_15_ ( .D(x3_o0_tmp[15]), .CK(clk), .RN(rstn), .Q(
        x3_o0[15]) );
  DFFRHQX1 x2_e_reg_19_ ( .D(x2_e_tmp[19]), .CK(clk), .RN(rstn), .Q(x2_e[19])
         );
  DFFRHQX1 x2_e_reg_18_ ( .D(x2_e_tmp[18]), .CK(clk), .RN(rstn), .Q(x2_e[18])
         );
  DFFRHQX1 x2_e_reg_17_ ( .D(x2_e_tmp[17]), .CK(clk), .RN(rstn), .Q(x2_e[17])
         );
  DFFRHQX1 x2_e_reg_16_ ( .D(x2_e_tmp[16]), .CK(clk), .RN(rstn), .Q(x2_e[16])
         );
  DFFRHQX1 x2_e_reg_15_ ( .D(x2_e_tmp[15]), .CK(clk), .RN(rstn), .Q(x2_e[15])
         );
  DFFRHQX1 o1_reg_21_ ( .D(N346), .CK(clk), .RN(rstn), .Q(o1[21]) );
  DFFRHQX1 o1_reg_20_ ( .D(N345), .CK(clk), .RN(rstn), .Q(o1[20]) );
  DFFRHQX1 o1_reg_19_ ( .D(N344), .CK(clk), .RN(rstn), .Q(o1[19]) );
  DFFRHQX1 o1_reg_18_ ( .D(N343), .CK(clk), .RN(rstn), .Q(o1[18]) );
  DFFRHQX1 o1_reg_17_ ( .D(N342), .CK(clk), .RN(rstn), .Q(o1[17]) );
  DFFRHQX1 o0_reg_21_ ( .D(N370), .CK(clk), .RN(rstn), .Q(o0[21]) );
  DFFRHQX1 o0_reg_20_ ( .D(N369), .CK(clk), .RN(rstn), .Q(o0[20]) );
  DFFRHQX1 o0_reg_19_ ( .D(N368), .CK(clk), .RN(rstn), .Q(o0[19]) );
  DFFRHQX1 o0_reg_18_ ( .D(N367), .CK(clk), .RN(rstn), .Q(o0[18]) );
  DFFRHQX1 o0_reg_17_ ( .D(N366), .CK(clk), .RN(rstn), .Q(o0[17]) );
  DFFRHQX1 x3_o1_tmp1_reg_14_ ( .D(N111), .CK(clk), .RN(rstn), .Q(
        x3_o1_tmp1[14]) );
  DFFRHQX1 x3_o1_tmp1_reg_13_ ( .D(N110), .CK(clk), .RN(rstn), .Q(
        x3_o1_tmp1[13]) );
  DFFRHQX1 x3_o1_tmp1_reg_12_ ( .D(N109), .CK(clk), .RN(rstn), .Q(
        x3_o1_tmp1[12]) );
  DFFRHQX1 x3_o1_tmp1_reg_11_ ( .D(N108), .CK(clk), .RN(rstn), .Q(
        x3_o1_tmp1[11]) );
  DFFRHQX1 x3_o1_tmp1_reg_10_ ( .D(N107), .CK(clk), .RN(rstn), .Q(
        x3_o1_tmp1[10]) );
  DFFRHQX1 x1_o0_tmp1_reg_14_ ( .D(N67), .CK(clk), .RN(rstn), .Q(
        x1_o0_tmp1[14]) );
  DFFRHQX1 x1_o0_tmp1_reg_13_ ( .D(N66), .CK(clk), .RN(rstn), .Q(
        x1_o0_tmp1[13]) );
  DFFRHQX1 x1_o0_tmp1_reg_12_ ( .D(N65), .CK(clk), .RN(rstn), .Q(
        x1_o0_tmp1[12]) );
  DFFRHQX1 x1_o0_tmp1_reg_11_ ( .D(N64), .CK(clk), .RN(rstn), .Q(
        x1_o0_tmp1[11]) );
  DFFRHQX1 x1_o0_tmp1_reg_10_ ( .D(N63), .CK(clk), .RN(rstn), .Q(
        x1_o0_tmp1[10]) );
  DFFRHQX1 x1_o0_reg_11_ ( .D(N152), .CK(clk), .RN(rstn), .Q(x1_o0[11]) );
  DFFRHQX1 x1_o0_reg_12_ ( .D(N153), .CK(clk), .RN(rstn), .Q(x1_o0[12]) );
  DFFRHQX1 x1_o0_reg_13_ ( .D(N154), .CK(clk), .RN(rstn), .Q(x1_o0[13]) );
  DFFRHQX1 x1_o0_reg_14_ ( .D(N155), .CK(clk), .RN(rstn), .Q(x1_o0[14]) );
  DFFRHQX1 x1_o0_reg_15_ ( .D(N156), .CK(clk), .RN(rstn), .Q(x1_o0[15]) );
  DFFRHQX1 x1_o1_reg_15_ ( .D(x1_o1_tmp[15]), .CK(clk), .RN(rstn), .Q(
        x1_o1[15]) );
  DFFRHQX1 x1_o1_reg_14_ ( .D(x1_o1_tmp[14]), .CK(clk), .RN(rstn), .Q(
        x1_o1[14]) );
  DFFRHQX1 x1_o1_reg_13_ ( .D(x1_o1_tmp[13]), .CK(clk), .RN(rstn), .Q(
        x1_o1[13]) );
  DFFRHQX1 x1_o1_reg_12_ ( .D(x1_o1_tmp[12]), .CK(clk), .RN(rstn), .Q(
        x1_o1[12]) );
  DFFRHQX1 x1_o1_reg_11_ ( .D(x1_o1_tmp[11]), .CK(clk), .RN(rstn), .Q(
        x1_o1[11]) );
  DFFRHQX1 x3_o1_reg_15_ ( .D(N179), .CK(clk), .RN(rstn), .Q(x3_o1[15]) );
  DFFRHQX1 x3_o1_reg_14_ ( .D(N178), .CK(clk), .RN(rstn), .Q(x3_o1[14]) );
  DFFRHQX1 x3_o1_reg_13_ ( .D(N177), .CK(clk), .RN(rstn), .Q(x3_o1[13]) );
  DFFRHQX1 x3_o1_reg_12_ ( .D(N176), .CK(clk), .RN(rstn), .Q(x3_o1[12]) );
  DFFRHQX1 x0_e_reg_14_ ( .D(x0_e_tmp[14]), .CK(clk), .RN(rstn), .Q(x0_e[14])
         );
  DFFRHQX1 x0_e_reg_13_ ( .D(x0_e_tmp[13]), .CK(clk), .RN(rstn), .Q(x0_e[13])
         );
  DFFRHQX1 x0_e_reg_12_ ( .D(x0_e_tmp[12]), .CK(clk), .RN(rstn), .Q(x0_e[12])
         );
  DFFRHQX1 x0_e_reg_11_ ( .D(x0_e_tmp[11]), .CK(clk), .RN(rstn), .Q(x0_e[11])
         );
  DFFRHQX1 e1_reg_16_ ( .D(N271), .CK(clk), .RN(rstn), .Q(e1[16]) );
  DFFRHQX1 e1_reg_15_ ( .D(N270), .CK(clk), .RN(rstn), .Q(e1[15]) );
  DFFRHQX1 e1_reg_14_ ( .D(N269), .CK(clk), .RN(rstn), .Q(e1[14]) );
  DFFRHQX1 e1_reg_13_ ( .D(N268), .CK(clk), .RN(rstn), .Q(e1[13]) );
  DFFRHQX1 e0_reg_16_ ( .D(N203), .CK(clk), .RN(rstn), .Q(e0[16]) );
  DFFRHQX1 e0_reg_15_ ( .D(N202), .CK(clk), .RN(rstn), .Q(e0[15]) );
  DFFRHQX1 e0_reg_14_ ( .D(N201), .CK(clk), .RN(rstn), .Q(e0[14]) );
  DFFRHQX1 e0_reg_13_ ( .D(N200), .CK(clk), .RN(rstn), .Q(e0[13]) );
  DFFRHQX1 x3_o1_tmp2_reg_13_ ( .D(N133), .CK(clk), .RN(rstn), .Q(
        x3_o1_tmp2[13]) );
  DFFRHQX1 x3_o1_tmp2_reg_12_ ( .D(N132), .CK(clk), .RN(rstn), .Q(
        x3_o1_tmp2[12]) );
  DFFRHQX1 x3_o1_tmp2_reg_11_ ( .D(N131), .CK(clk), .RN(rstn), .Q(
        x3_o1_tmp2[11]) );
  DFFRHQX1 x3_o1_tmp2_reg_10_ ( .D(N130), .CK(clk), .RN(rstn), .Q(
        x3_o1_tmp2[10]) );
  DFFRHQX1 x1_o0_tmp2_reg_13_ ( .D(N89), .CK(clk), .RN(rstn), .Q(
        x1_o0_tmp2[13]) );
  DFFRHQX1 x1_o0_tmp2_reg_12_ ( .D(N88), .CK(clk), .RN(rstn), .Q(
        x1_o0_tmp2[12]) );
  DFFRHQX1 x1_o0_tmp2_reg_11_ ( .D(N87), .CK(clk), .RN(rstn), .Q(
        x1_o0_tmp2[11]) );
  DFFRHQX1 x1_o0_tmp2_reg_10_ ( .D(N86), .CK(clk), .RN(rstn), .Q(
        x1_o0_tmp2[10]) );
  DFFRHQX1 x3_o0_reg_14_ ( .D(x3_o0_tmp[14]), .CK(clk), .RN(rstn), .Q(
        x3_o0[14]) );
  DFFRHQX1 x3_o0_reg_13_ ( .D(x3_o0_tmp[13]), .CK(clk), .RN(rstn), .Q(
        x3_o0[13]) );
  DFFRHQX1 x3_o0_reg_12_ ( .D(x3_o0_tmp[12]), .CK(clk), .RN(rstn), .Q(
        x3_o0[12]) );
  DFFRHQX1 x3_o0_reg_11_ ( .D(x3_o0_tmp[11]), .CK(clk), .RN(rstn), .Q(
        x3_o0[11]) );
  DFFRHQX1 x2_e_reg_14_ ( .D(x2_e_tmp[14]), .CK(clk), .RN(rstn), .Q(x2_e[14])
         );
  DFFRHQX1 x2_e_reg_13_ ( .D(x2_e_tmp[13]), .CK(clk), .RN(rstn), .Q(x2_e[13])
         );
  DFFRHQX1 x2_e_reg_12_ ( .D(x2_e_tmp[12]), .CK(clk), .RN(rstn), .Q(x2_e[12])
         );
  DFFRHQX1 x2_e_reg_11_ ( .D(x2_e_tmp[11]), .CK(clk), .RN(rstn), .Q(x2_e[11])
         );
  DFFRHQX1 o1_reg_16_ ( .D(N341), .CK(clk), .RN(rstn), .Q(o1[16]) );
  DFFRHQX1 o1_reg_15_ ( .D(N340), .CK(clk), .RN(rstn), .Q(o1[15]) );
  DFFRHQX1 o1_reg_14_ ( .D(N339), .CK(clk), .RN(rstn), .Q(o1[14]) );
  DFFRHQX1 o1_reg_13_ ( .D(N338), .CK(clk), .RN(rstn), .Q(o1[13]) );
  DFFRHQX1 o0_reg_16_ ( .D(N365), .CK(clk), .RN(rstn), .Q(o0[16]) );
  DFFRHQX1 o0_reg_15_ ( .D(N364), .CK(clk), .RN(rstn), .Q(o0[15]) );
  DFFRHQX1 o0_reg_14_ ( .D(N363), .CK(clk), .RN(rstn), .Q(o0[14]) );
  DFFRHQX1 o0_reg_13_ ( .D(N362), .CK(clk), .RN(rstn), .Q(o0[13]) );
  DFFRHQX1 x3_o1_tmp1_reg_9_ ( .D(N106), .CK(clk), .RN(rstn), .Q(x3_o1_tmp1[9]) );
  DFFRHQX1 x3_o1_tmp1_reg_8_ ( .D(N105), .CK(clk), .RN(rstn), .Q(x3_o1_tmp1[8]) );
  DFFRHQX1 x3_o1_tmp1_reg_7_ ( .D(N104), .CK(clk), .RN(rstn), .Q(x3_o1_tmp1[7]) );
  DFFRHQX1 x3_o1_tmp1_reg_6_ ( .D(N103), .CK(clk), .RN(rstn), .Q(x3_o1_tmp1[6]) );
  DFFRHQX1 x1_o0_tmp1_reg_9_ ( .D(N62), .CK(clk), .RN(rstn), .Q(x1_o0_tmp1[9])
         );
  DFFRHQX1 x1_o0_tmp1_reg_8_ ( .D(N61), .CK(clk), .RN(rstn), .Q(x1_o0_tmp1[8])
         );
  DFFRHQX1 x1_o0_tmp1_reg_7_ ( .D(N60), .CK(clk), .RN(rstn), .Q(x1_o0_tmp1[7])
         );
  DFFRHQX1 x1_o0_tmp1_reg_6_ ( .D(N59), .CK(clk), .RN(rstn), .Q(x1_o0_tmp1[6])
         );
  DFFRHQX1 x1_o0_reg_7_ ( .D(N148), .CK(clk), .RN(rstn), .Q(x1_o0[7]) );
  DFFRHQX1 x1_o0_reg_8_ ( .D(N149), .CK(clk), .RN(rstn), .Q(x1_o0[8]) );
  DFFRHQX1 x1_o0_reg_9_ ( .D(N150), .CK(clk), .RN(rstn), .Q(x1_o0[9]) );
  DFFRHQX1 x1_o0_reg_10_ ( .D(N151), .CK(clk), .RN(rstn), .Q(x1_o0[10]) );
  DFFRHQX1 x1_o1_reg_10_ ( .D(x1_o1_tmp[10]), .CK(clk), .RN(rstn), .Q(
        x1_o1[10]) );
  DFFRHQX1 x1_o1_reg_9_ ( .D(x1_o1_tmp[9]), .CK(clk), .RN(rstn), .Q(x1_o1[9])
         );
  DFFRHQX1 x1_o1_reg_8_ ( .D(x1_o1_tmp[8]), .CK(clk), .RN(rstn), .Q(x1_o1[8])
         );
  DFFRHQX1 x1_o1_reg_7_ ( .D(x1_o1_tmp[7]), .CK(clk), .RN(rstn), .Q(x1_o1[7])
         );
  DFFRHQX1 x0_e_reg_6_ ( .D(x0_e_tmp[6]), .CK(clk), .RN(rstn), .Q(x0_e[6]) );
  DFFRHQX1 y1_tmp_reg_10_ ( .D(N408), .CK(clk), .RN(rstn), .Q(y1_tmp[10]) );
  DFFRHQX1 y2_tmp_reg_10_ ( .D(N482), .CK(clk), .RN(rstn), .Q(y2_tmp[10]) );
  DFFRHQX1 y0_tmp_reg_10_ ( .D(N383), .CK(clk), .RN(rstn), .Q(y0_tmp[10]) );
  DFFRHQX1 y3_tmp_reg_10_ ( .D(N556), .CK(clk), .RN(rstn), .Q(y3_tmp[10]) );
  DFFRHQX1 y1_tmp_reg_24_ ( .D(N422), .CK(clk), .RN(rstn), .Q(y1_tmp[24]) );
  DFFRHQX1 y2_tmp_reg_24_ ( .D(N496), .CK(clk), .RN(rstn), .Q(y2_tmp[24]) );
  DFFRHQX1 y0_tmp_reg_24_ ( .D(N397), .CK(clk), .RN(rstn), .Q(y0_tmp[24]) );
  DFFRHQX1 y3_tmp_reg_24_ ( .D(N570), .CK(clk), .RN(rstn), .Q(y3_tmp[24]) );
  DFFRHQX1 idct4_ready_reg ( .D(idct4_ready_delay3), .CK(clk), .RN(rstn), .Q(
        idct4_ready) );
  DFFRHQX1 x3_o1_reg_11_ ( .D(N175), .CK(clk), .RN(rstn), .Q(x3_o1[11]) );
  DFFRHQX1 x3_o1_reg_10_ ( .D(N174), .CK(clk), .RN(rstn), .Q(x3_o1[10]) );
  DFFRHQX1 x3_o1_reg_9_ ( .D(N173), .CK(clk), .RN(rstn), .Q(x3_o1[9]) );
  DFFRHQX1 x3_o1_reg_8_ ( .D(N172), .CK(clk), .RN(rstn), .Q(x3_o1[8]) );
  DFFRHQX1 x3_o1_reg_7_ ( .D(N171), .CK(clk), .RN(rstn), .Q(x3_o1[7]) );
  DFFRHQX1 x0_e_reg_10_ ( .D(x0_e_tmp[10]), .CK(clk), .RN(rstn), .Q(x0_e[10])
         );
  DFFRHQX1 x0_e_reg_9_ ( .D(x0_e_tmp[9]), .CK(clk), .RN(rstn), .Q(x0_e[9]) );
  DFFRHQX1 x0_e_reg_8_ ( .D(x0_e_tmp[8]), .CK(clk), .RN(rstn), .Q(x0_e[8]) );
  DFFRHQX1 x0_e_reg_7_ ( .D(x0_e_tmp[7]), .CK(clk), .RN(rstn), .Q(x0_e[7]) );
  DFFRHQX1 e1_reg_12_ ( .D(N267), .CK(clk), .RN(rstn), .Q(e1[12]) );
  DFFRHQX1 e1_reg_11_ ( .D(N266), .CK(clk), .RN(rstn), .Q(e1[11]) );
  DFFRHQX1 e1_reg_10_ ( .D(N265), .CK(clk), .RN(rstn), .Q(e1[10]) );
  DFFRHQX1 e1_reg_9_ ( .D(N264), .CK(clk), .RN(rstn), .Q(e1[9]) );
  DFFRHQX1 e1_reg_8_ ( .D(N263), .CK(clk), .RN(rstn), .Q(e1[8]) );
  DFFRHQX1 e0_reg_12_ ( .D(N199), .CK(clk), .RN(rstn), .Q(e0[12]) );
  DFFRHQX1 e0_reg_11_ ( .D(N198), .CK(clk), .RN(rstn), .Q(e0[11]) );
  DFFRHQX1 e0_reg_10_ ( .D(N197), .CK(clk), .RN(rstn), .Q(e0[10]) );
  DFFRHQX1 e0_reg_9_ ( .D(N196), .CK(clk), .RN(rstn), .Q(e0[9]) );
  DFFRHQX1 e0_reg_8_ ( .D(N195), .CK(clk), .RN(rstn), .Q(e0[8]) );
  DFFRHQX1 x3_o1_tmp2_reg_9_ ( .D(N129), .CK(clk), .RN(rstn), .Q(x3_o1_tmp2[9]) );
  DFFRHQX1 x3_o1_tmp2_reg_8_ ( .D(N128), .CK(clk), .RN(rstn), .Q(x3_o1_tmp2[8]) );
  DFFRHQX1 x3_o1_tmp2_reg_7_ ( .D(N127), .CK(clk), .RN(rstn), .Q(x3_o1_tmp2[7]) );
  DFFRHQX1 x3_o1_tmp2_reg_6_ ( .D(N126), .CK(clk), .RN(rstn), .Q(x3_o1_tmp2[6]) );
  DFFRHQX1 x1_o0_tmp2_reg_9_ ( .D(N85), .CK(clk), .RN(rstn), .Q(x1_o0_tmp2[9])
         );
  DFFRHQX1 x1_o0_tmp2_reg_8_ ( .D(N84), .CK(clk), .RN(rstn), .Q(x1_o0_tmp2[8])
         );
  DFFRHQX1 x1_o0_tmp2_reg_7_ ( .D(N83), .CK(clk), .RN(rstn), .Q(x1_o0_tmp2[7])
         );
  DFFRHQX1 x1_o0_tmp2_reg_6_ ( .D(N82), .CK(clk), .RN(rstn), .Q(x1_o0_tmp2[6])
         );
  DFFRHQX1 x3_o0_reg_10_ ( .D(x3_o0_tmp[10]), .CK(clk), .RN(rstn), .Q(
        x3_o0[10]) );
  DFFRHQX1 x3_o0_reg_9_ ( .D(x3_o0_tmp[9]), .CK(clk), .RN(rstn), .Q(x3_o0[9])
         );
  DFFRHQX1 x3_o0_reg_8_ ( .D(x3_o0_tmp[8]), .CK(clk), .RN(rstn), .Q(x3_o0[8])
         );
  DFFRHQX1 x3_o0_reg_7_ ( .D(x3_o0_tmp[7]), .CK(clk), .RN(rstn), .Q(x3_o0[7])
         );
  DFFRHQX1 x2_e_reg_6_ ( .D(x2_e_tmp[6]), .CK(clk), .RN(rstn), .Q(x2_e[6]) );
  DFFRHQX1 x2_e_reg_10_ ( .D(x2_e_tmp[10]), .CK(clk), .RN(rstn), .Q(x2_e[10])
         );
  DFFRHQX1 x2_e_reg_9_ ( .D(x2_e_tmp[9]), .CK(clk), .RN(rstn), .Q(x2_e[9]) );
  DFFRHQX1 x2_e_reg_8_ ( .D(x2_e_tmp[8]), .CK(clk), .RN(rstn), .Q(x2_e[8]) );
  DFFRHQX1 x2_e_reg_7_ ( .D(x2_e_tmp[7]), .CK(clk), .RN(rstn), .Q(x2_e[7]) );
  DFFRHQX1 o1_reg_12_ ( .D(N337), .CK(clk), .RN(rstn), .Q(o1[12]) );
  DFFRHQX1 o1_reg_11_ ( .D(N336), .CK(clk), .RN(rstn), .Q(o1[11]) );
  DFFRHQX1 o1_reg_10_ ( .D(N335), .CK(clk), .RN(rstn), .Q(o1[10]) );
  DFFRHQX1 o1_reg_9_ ( .D(N334), .CK(clk), .RN(rstn), .Q(o1[9]) );
  DFFRHQX1 o0_reg_12_ ( .D(N361), .CK(clk), .RN(rstn), .Q(o0[12]) );
  DFFRHQX1 o0_reg_11_ ( .D(N360), .CK(clk), .RN(rstn), .Q(o0[11]) );
  DFFRHQX1 o0_reg_10_ ( .D(N359), .CK(clk), .RN(rstn), .Q(o0[10]) );
  DFFRHQX1 o0_reg_9_ ( .D(N358), .CK(clk), .RN(rstn), .Q(o0[9]) );
  DFFRHQX1 x3_o1_tmp1_reg_5_ ( .D(x3[5]), .CK(clk), .RN(rstn), .Q(
        x3_o1_tmp1[5]) );
  DFFRHQX1 x3_o1_tmp1_reg_4_ ( .D(x3[4]), .CK(clk), .RN(rstn), .Q(
        x3_o1_tmp1[4]) );
  DFFRHQX1 x3_o1_tmp1_reg_3_ ( .D(x3[3]), .CK(clk), .RN(rstn), .Q(
        x3_o1_tmp1[3]) );
  DFFRHQX1 x3_o1_tmp1_reg_2_ ( .D(x3[2]), .CK(clk), .RN(rstn), .Q(
        x3_o1_tmp1[2]) );
  DFFRHQX1 x1_o0_tmp1_reg_5_ ( .D(x1[5]), .CK(clk), .RN(rstn), .Q(
        x1_o0_tmp1[5]) );
  DFFRHQX1 x1_o0_tmp1_reg_4_ ( .D(x1[4]), .CK(clk), .RN(rstn), .Q(
        x1_o0_tmp1[4]) );
  DFFRHQX1 x1_o0_tmp1_reg_3_ ( .D(x1[3]), .CK(clk), .RN(rstn), .Q(
        x1_o0_tmp1[3]) );
  DFFRHQX1 x1_o0_tmp1_reg_2_ ( .D(x1[2]), .CK(clk), .RN(rstn), .Q(
        x1_o0_tmp1[2]) );
  DFFRHQX1 x1_o0_reg_3_ ( .D(N144), .CK(clk), .RN(rstn), .Q(x1_o0[3]) );
  DFFRHQX1 x1_o0_reg_4_ ( .D(N145), .CK(clk), .RN(rstn), .Q(x1_o0[4]) );
  DFFRHQX1 x1_o0_reg_5_ ( .D(N146), .CK(clk), .RN(rstn), .Q(x1_o0[5]) );
  DFFRHQX1 x1_o0_reg_6_ ( .D(N147), .CK(clk), .RN(rstn), .Q(x1_o0[6]) );
  DFFRHQX1 x1_o1_reg_6_ ( .D(x1_o1_tmp[6]), .CK(clk), .RN(rstn), .Q(x1_o1[6])
         );
  DFFRHQX1 x1_o1_reg_5_ ( .D(x1_o1_tmp[5]), .CK(clk), .RN(rstn), .Q(x1_o1[5])
         );
  DFFRHQX1 x1_o1_reg_4_ ( .D(x1_o1_tmp[4]), .CK(clk), .RN(rstn), .Q(x1_o1[4])
         );
  DFFRHQX1 x1_o1_reg_3_ ( .D(x1_o1_tmp[3]), .CK(clk), .RN(rstn), .Q(x1_o1[3])
         );
  DFFRHQX1 y1_tmp_reg_23_ ( .D(N421), .CK(clk), .RN(rstn), .Q(y1_tmp[23]) );
  DFFRHQX1 y1_tmp_reg_22_ ( .D(N420), .CK(clk), .RN(rstn), .Q(y1_tmp[22]) );
  DFFRHQX1 y1_tmp_reg_21_ ( .D(N419), .CK(clk), .RN(rstn), .Q(y1_tmp[21]) );
  DFFRHQX1 y1_tmp_reg_20_ ( .D(N418), .CK(clk), .RN(rstn), .Q(y1_tmp[20]) );
  DFFRHQX1 y2_tmp_reg_23_ ( .D(N495), .CK(clk), .RN(rstn), .Q(y2_tmp[23]) );
  DFFRHQX1 y2_tmp_reg_22_ ( .D(N494), .CK(clk), .RN(rstn), .Q(y2_tmp[22]) );
  DFFRHQX1 y2_tmp_reg_21_ ( .D(N493), .CK(clk), .RN(rstn), .Q(y2_tmp[21]) );
  DFFRHQX1 y2_tmp_reg_20_ ( .D(N492), .CK(clk), .RN(rstn), .Q(y2_tmp[20]) );
  DFFRHQX1 y0_tmp_reg_20_ ( .D(N393), .CK(clk), .RN(rstn), .Q(y0_tmp[20]) );
  DFFRHQX1 y0_tmp_reg_21_ ( .D(N394), .CK(clk), .RN(rstn), .Q(y0_tmp[21]) );
  DFFRHQX1 y0_tmp_reg_22_ ( .D(N395), .CK(clk), .RN(rstn), .Q(y0_tmp[22]) );
  DFFRHQX1 y0_tmp_reg_23_ ( .D(N396), .CK(clk), .RN(rstn), .Q(y0_tmp[23]) );
  DFFRHQX1 y3_tmp_reg_20_ ( .D(N566), .CK(clk), .RN(rstn), .Q(y3_tmp[20]) );
  DFFRHQX1 y3_tmp_reg_21_ ( .D(N567), .CK(clk), .RN(rstn), .Q(y3_tmp[21]) );
  DFFRHQX1 y3_tmp_reg_22_ ( .D(N568), .CK(clk), .RN(rstn), .Q(y3_tmp[22]) );
  DFFRHQX1 y3_tmp_reg_23_ ( .D(N569), .CK(clk), .RN(rstn), .Q(y3_tmp[23]) );
  DFFRHQX1 y1_tmp_reg_9_ ( .D(N407), .CK(clk), .RN(rstn), .Q(y1_tmp[9]) );
  DFFRHQX1 y1_tmp_reg_8_ ( .D(N406), .CK(clk), .RN(rstn), .Q(y1_tmp[8]) );
  DFFRHQX1 y1_tmp_reg_7_ ( .D(N405), .CK(clk), .RN(rstn), .Q(y1_tmp[7]) );
  DFFRHQX1 y1_tmp_reg_6_ ( .D(N404), .CK(clk), .RN(rstn), .Q(y1_tmp[6]) );
  DFFRHQX1 y2_tmp_reg_9_ ( .D(N481), .CK(clk), .RN(rstn), .Q(y2_tmp[9]) );
  DFFRHQX1 y2_tmp_reg_8_ ( .D(N480), .CK(clk), .RN(rstn), .Q(y2_tmp[8]) );
  DFFRHQX1 y2_tmp_reg_7_ ( .D(N479), .CK(clk), .RN(rstn), .Q(y2_tmp[7]) );
  DFFRHQX1 y2_tmp_reg_6_ ( .D(N478), .CK(clk), .RN(rstn), .Q(y2_tmp[6]) );
  DFFRHQX1 y0_tmp_reg_6_ ( .D(N379), .CK(clk), .RN(rstn), .Q(y0_tmp[6]) );
  DFFRHQX1 y0_tmp_reg_7_ ( .D(N380), .CK(clk), .RN(rstn), .Q(y0_tmp[7]) );
  DFFRHQX1 y0_tmp_reg_8_ ( .D(N381), .CK(clk), .RN(rstn), .Q(y0_tmp[8]) );
  DFFRHQX1 y0_tmp_reg_9_ ( .D(N382), .CK(clk), .RN(rstn), .Q(y0_tmp[9]) );
  DFFRHQX1 y3_tmp_reg_6_ ( .D(N552), .CK(clk), .RN(rstn), .Q(y3_tmp[6]) );
  DFFRHQX1 y3_tmp_reg_7_ ( .D(N553), .CK(clk), .RN(rstn), .Q(y3_tmp[7]) );
  DFFRHQX1 y3_tmp_reg_8_ ( .D(N554), .CK(clk), .RN(rstn), .Q(y3_tmp[8]) );
  DFFRHQX1 y3_tmp_reg_9_ ( .D(N555), .CK(clk), .RN(rstn), .Q(y3_tmp[9]) );
  DFFRHQX1 x3_o1_reg_6_ ( .D(N170), .CK(clk), .RN(rstn), .Q(x3_o1[6]) );
  DFFRHQX1 x3_o1_reg_5_ ( .D(N169), .CK(clk), .RN(rstn), .Q(x3_o1[5]) );
  DFFRHQX1 x3_o1_reg_4_ ( .D(N168), .CK(clk), .RN(rstn), .Q(x3_o1[4]) );
  DFFRHQX1 x3_o1_reg_3_ ( .D(N167), .CK(clk), .RN(rstn), .Q(x3_o1[3]) );
  DFFRHQX1 e1_reg_7_ ( .D(N262), .CK(clk), .RN(rstn), .Q(e1[7]) );
  DFFRHQX1 e1_reg_6_ ( .D(N261), .CK(clk), .RN(rstn), .Q(e1[6]) );
  DFFRHQX1 e0_reg_7_ ( .D(N194), .CK(clk), .RN(rstn), .Q(e0[7]) );
  DFFRHQX1 e0_reg_6_ ( .D(N193), .CK(clk), .RN(rstn), .Q(e0[6]) );
  DFFRHQX1 x3_o1_tmp2_reg_5_ ( .D(N125), .CK(clk), .RN(rstn), .Q(x3_o1_tmp2[5]) );
  DFFRHQX1 x3_o1_tmp2_reg_4_ ( .D(N124), .CK(clk), .RN(rstn), .Q(x3_o1_tmp2[4]) );
  DFFRHQX1 x3_o1_tmp2_reg_3_ ( .D(x3[2]), .CK(clk), .RN(rstn), .Q(
        x3_o1_tmp2[3]) );
  DFFRHQX1 x3_o1_tmp2_reg_2_ ( .D(x3[1]), .CK(clk), .RN(rstn), .Q(
        x3_o1_tmp2[2]) );
  DFFRHQX1 x3_o1_tmp2_reg_1_ ( .D(x3[0]), .CK(clk), .RN(rstn), .Q(
        x3_o1_tmp2[1]) );
  DFFRHQX1 x1_o0_tmp2_reg_5_ ( .D(N81), .CK(clk), .RN(rstn), .Q(x1_o0_tmp2[5])
         );
  DFFRHQX1 x1_o0_tmp2_reg_4_ ( .D(N80), .CK(clk), .RN(rstn), .Q(x1_o0_tmp2[4])
         );
  DFFRHQX1 x1_o0_tmp2_reg_3_ ( .D(x1[2]), .CK(clk), .RN(rstn), .Q(
        x1_o0_tmp2[3]) );
  DFFRHQX1 x1_o0_tmp2_reg_2_ ( .D(x1[1]), .CK(clk), .RN(rstn), .Q(
        x1_o0_tmp2[2]) );
  DFFRHQX1 x1_o0_tmp2_reg_1_ ( .D(x1[0]), .CK(clk), .RN(rstn), .Q(
        x1_o0_tmp2[1]) );
  DFFRHQX1 x3_o0_reg_6_ ( .D(x3_o0_tmp[6]), .CK(clk), .RN(rstn), .Q(x3_o0[6])
         );
  DFFRHQX1 x3_o0_reg_5_ ( .D(x3_o0_tmp[5]), .CK(clk), .RN(rstn), .Q(x3_o0[5])
         );
  DFFRHQX1 x3_o0_reg_4_ ( .D(x3_o0_tmp[4]), .CK(clk), .RN(rstn), .Q(x3_o0[4])
         );
  DFFRHQX1 x3_o0_reg_3_ ( .D(x3_o0_tmp[3]), .CK(clk), .RN(rstn), .Q(x3_o0[3])
         );
  DFFRHQX1 x3_o0_reg_2_ ( .D(x3_o0_tmp[2]), .CK(clk), .RN(rstn), .Q(x3_o0[2])
         );
  DFFRHQX1 o1_reg_8_ ( .D(N333), .CK(clk), .RN(rstn), .Q(o1[8]) );
  DFFRHQX1 o1_reg_7_ ( .D(N332), .CK(clk), .RN(rstn), .Q(o1[7]) );
  DFFRHQX1 o1_reg_6_ ( .D(N331), .CK(clk), .RN(rstn), .Q(o1[6]) );
  DFFRHQX1 o1_reg_5_ ( .D(N330), .CK(clk), .RN(rstn), .Q(o1[5]) );
  DFFRHQX1 o1_reg_4_ ( .D(N329), .CK(clk), .RN(rstn), .Q(o1[4]) );
  DFFRHQX1 o0_reg_8_ ( .D(N357), .CK(clk), .RN(rstn), .Q(o0[8]) );
  DFFRHQX1 o0_reg_7_ ( .D(N356), .CK(clk), .RN(rstn), .Q(o0[7]) );
  DFFRHQX1 o0_reg_6_ ( .D(N355), .CK(clk), .RN(rstn), .Q(o0[6]) );
  DFFRHQX1 o0_reg_5_ ( .D(N354), .CK(clk), .RN(rstn), .Q(o0[5]) );
  DFFRHQX1 o0_reg_4_ ( .D(N353), .CK(clk), .RN(rstn), .Q(o0[4]) );
  DFFRHQX1 x3_o1_tmp1_reg_1_ ( .D(x3[1]), .CK(clk), .RN(rstn), .Q(
        x3_o1_tmp1[1]) );
  DFFRHQX1 x1_o0_tmp1_reg_1_ ( .D(x1[1]), .CK(clk), .RN(rstn), .Q(
        x1_o0_tmp1[1]) );
  DFFRHQX1 x1_o0_reg_1_ ( .D(N142), .CK(clk), .RN(rstn), .Q(x1_o0[1]) );
  DFFRHQX1 x1_o0_reg_2_ ( .D(N143), .CK(clk), .RN(rstn), .Q(x1_o0[2]) );
  DFFRHQX1 x1_o1_reg_2_ ( .D(x1_o1_tmp[2]), .CK(clk), .RN(rstn), .Q(x1_o1[2])
         );
  DFFRHQX1 y1_tmp_reg_19_ ( .D(N417), .CK(clk), .RN(rstn), .Q(y1_tmp[19]) );
  DFFRHQX1 y1_tmp_reg_18_ ( .D(N416), .CK(clk), .RN(rstn), .Q(y1_tmp[18]) );
  DFFRHQX1 y1_tmp_reg_17_ ( .D(N415), .CK(clk), .RN(rstn), .Q(y1_tmp[17]) );
  DFFRHQX1 y1_tmp_reg_16_ ( .D(N414), .CK(clk), .RN(rstn), .Q(y1_tmp[16]) );
  DFFRHQX1 y1_tmp_reg_15_ ( .D(N413), .CK(clk), .RN(rstn), .Q(y1_tmp[15]) );
  DFFRHQX1 y2_tmp_reg_19_ ( .D(N491), .CK(clk), .RN(rstn), .Q(y2_tmp[19]) );
  DFFRHQX1 y2_tmp_reg_18_ ( .D(N490), .CK(clk), .RN(rstn), .Q(y2_tmp[18]) );
  DFFRHQX1 y2_tmp_reg_17_ ( .D(N489), .CK(clk), .RN(rstn), .Q(y2_tmp[17]) );
  DFFRHQX1 y2_tmp_reg_16_ ( .D(N488), .CK(clk), .RN(rstn), .Q(y2_tmp[16]) );
  DFFRHQX1 y2_tmp_reg_15_ ( .D(N487), .CK(clk), .RN(rstn), .Q(y2_tmp[15]) );
  DFFRHQX1 y0_tmp_reg_15_ ( .D(N388), .CK(clk), .RN(rstn), .Q(y0_tmp[15]) );
  DFFRHQX1 y0_tmp_reg_16_ ( .D(N389), .CK(clk), .RN(rstn), .Q(y0_tmp[16]) );
  DFFRHQX1 y0_tmp_reg_17_ ( .D(N390), .CK(clk), .RN(rstn), .Q(y0_tmp[17]) );
  DFFRHQX1 y0_tmp_reg_18_ ( .D(N391), .CK(clk), .RN(rstn), .Q(y0_tmp[18]) );
  DFFRHQX1 y0_tmp_reg_19_ ( .D(N392), .CK(clk), .RN(rstn), .Q(y0_tmp[19]) );
  DFFRHQX1 y3_tmp_reg_15_ ( .D(N561), .CK(clk), .RN(rstn), .Q(y3_tmp[15]) );
  DFFRHQX1 y3_tmp_reg_16_ ( .D(N562), .CK(clk), .RN(rstn), .Q(y3_tmp[16]) );
  DFFRHQX1 y3_tmp_reg_17_ ( .D(N563), .CK(clk), .RN(rstn), .Q(y3_tmp[17]) );
  DFFRHQX1 y3_tmp_reg_18_ ( .D(N564), .CK(clk), .RN(rstn), .Q(y3_tmp[18]) );
  DFFRHQX1 y3_tmp_reg_19_ ( .D(N565), .CK(clk), .RN(rstn), .Q(y3_tmp[19]) );
  DFFRHQX1 y1_tmp_reg_5_ ( .D(N403), .CK(clk), .RN(rstn), .Q(y1_tmp[5]) );
  DFFRHQX1 y1_tmp_reg_4_ ( .D(N402), .CK(clk), .RN(rstn), .Q(y1_tmp[4]) );
  DFFRHQX1 y1_tmp_reg_3_ ( .D(N401), .CK(clk), .RN(rstn), .Q(y1_tmp[3]) );
  DFFRHQX1 y1_tmp_reg_2_ ( .D(N400), .CK(clk), .RN(rstn), .Q(y1_tmp[2]) );
  DFFRHQX1 y2_tmp_reg_5_ ( .D(N477), .CK(clk), .RN(rstn), .Q(y2_tmp[5]) );
  DFFRHQX1 y2_tmp_reg_4_ ( .D(N476), .CK(clk), .RN(rstn), .Q(y2_tmp[4]) );
  DFFRHQX1 y2_tmp_reg_3_ ( .D(N475), .CK(clk), .RN(rstn), .Q(y2_tmp[3]) );
  DFFRHQX1 y2_tmp_reg_2_ ( .D(N474), .CK(clk), .RN(rstn), .Q(y2_tmp[2]) );
  DFFRHQX1 y0_tmp_reg_2_ ( .D(N375), .CK(clk), .RN(rstn), .Q(y0_tmp[2]) );
  DFFRHQX1 y0_tmp_reg_3_ ( .D(N376), .CK(clk), .RN(rstn), .Q(y0_tmp[3]) );
  DFFRHQX1 y0_tmp_reg_4_ ( .D(N377), .CK(clk), .RN(rstn), .Q(y0_tmp[4]) );
  DFFRHQX1 y0_tmp_reg_5_ ( .D(N378), .CK(clk), .RN(rstn), .Q(y0_tmp[5]) );
  DFFRHQX1 y3_tmp_reg_2_ ( .D(N548), .CK(clk), .RN(rstn), .Q(y3_tmp[2]) );
  DFFRHQX1 y3_tmp_reg_3_ ( .D(N549), .CK(clk), .RN(rstn), .Q(y3_tmp[3]) );
  DFFRHQX1 y3_tmp_reg_4_ ( .D(N550), .CK(clk), .RN(rstn), .Q(y3_tmp[4]) );
  DFFRHQX1 y3_tmp_reg_5_ ( .D(N551), .CK(clk), .RN(rstn), .Q(y3_tmp[5]) );
  DFFRHQX1 x3_o1_reg_2_ ( .D(N166), .CK(clk), .RN(rstn), .Q(x3_o1[2]) );
  DFFRHQX1 x3_o1_reg_1_ ( .D(N165), .CK(clk), .RN(rstn), .Q(x3_o1[1]) );
  DFFRHQX1 x3_o1_reg_0_ ( .D(N164), .CK(clk), .RN(rstn), .Q(x3_o1[0]) );
  DFFRHQX1 o1_reg_0_ ( .D(N325), .CK(clk), .RN(rstn), .Q(o1[0]) );
  DFFRHQX1 o0_reg_0_ ( .D(N349), .CK(clk), .RN(rstn), .Q(o0[0]) );
  DFFRHQX1 o1_reg_3_ ( .D(N328), .CK(clk), .RN(rstn), .Q(o1[3]) );
  DFFRHQX1 o1_reg_2_ ( .D(N327), .CK(clk), .RN(rstn), .Q(o1[2]) );
  DFFRHQX1 o1_reg_1_ ( .D(N326), .CK(clk), .RN(rstn), .Q(o1[1]) );
  DFFRHQX1 o0_reg_3_ ( .D(N352), .CK(clk), .RN(rstn), .Q(o0[3]) );
  DFFRHQX1 o0_reg_2_ ( .D(N351), .CK(clk), .RN(rstn), .Q(o0[2]) );
  DFFRHQX1 o0_reg_1_ ( .D(N350), .CK(clk), .RN(rstn), .Q(o0[1]) );
  DFFRHQX1 y1_tmp_reg_14_ ( .D(N412), .CK(clk), .RN(rstn), .Q(y1_tmp[14]) );
  DFFRHQX1 y1_tmp_reg_13_ ( .D(N411), .CK(clk), .RN(rstn), .Q(y1_tmp[13]) );
  DFFRHQX1 y2_tmp_reg_14_ ( .D(N486), .CK(clk), .RN(rstn), .Q(y2_tmp[14]) );
  DFFRHQX1 y2_tmp_reg_13_ ( .D(N485), .CK(clk), .RN(rstn), .Q(y2_tmp[13]) );
  DFFRHQX1 y0_tmp_reg_13_ ( .D(N386), .CK(clk), .RN(rstn), .Q(y0_tmp[13]) );
  DFFRHQX1 y0_tmp_reg_14_ ( .D(N387), .CK(clk), .RN(rstn), .Q(y0_tmp[14]) );
  DFFRHQX1 y3_tmp_reg_13_ ( .D(N559), .CK(clk), .RN(rstn), .Q(y3_tmp[13]) );
  DFFRHQX1 y3_tmp_reg_14_ ( .D(N560), .CK(clk), .RN(rstn), .Q(y3_tmp[14]) );
  DFFRHQX1 y1_tmp_reg_1_ ( .D(N399), .CK(clk), .RN(rstn), .Q(y1_tmp[1]) );
  DFFRHQX1 y1_tmp_reg_0_ ( .D(N398), .CK(clk), .RN(rstn), .Q(y1_tmp[0]) );
  DFFRHQX1 y2_tmp_reg_1_ ( .D(N473), .CK(clk), .RN(rstn), .Q(y2_tmp[1]) );
  DFFRHQX1 y2_tmp_reg_0_ ( .D(N472), .CK(clk), .RN(rstn), .Q(y2_tmp[0]) );
  DFFRHQX1 y0_tmp_reg_0_ ( .D(N373), .CK(clk), .RN(rstn), .Q(y0_tmp[0]) );
  DFFRHQX1 y0_tmp_reg_1_ ( .D(N374), .CK(clk), .RN(rstn), .Q(y0_tmp[1]) );
  DFFRHQX1 y3_tmp_reg_0_ ( .D(N546), .CK(clk), .RN(rstn), .Q(y3_tmp[0]) );
  DFFRHQX1 y3_tmp_reg_1_ ( .D(N547), .CK(clk), .RN(rstn), .Q(y3_tmp[1]) );
  DFFRHQX1 y1_tmp_reg_12_ ( .D(N410), .CK(clk), .RN(rstn), .Q(y1_tmp[12]) );
  DFFRHQX1 y2_tmp_reg_12_ ( .D(N484), .CK(clk), .RN(rstn), .Q(y2_tmp[12]) );
  DFFRHQX1 y0_tmp_reg_12_ ( .D(N385), .CK(clk), .RN(rstn), .Q(y0_tmp[12]) );
  DFFRHQX1 y3_tmp_reg_12_ ( .D(N558), .CK(clk), .RN(rstn), .Q(y3_tmp[12]) );
  DFFRHQX1 y1_tmp_reg_11_ ( .D(N409), .CK(clk), .RN(rstn), .Q(y1_tmp[11]) );
  DFFRHQX1 y2_tmp_reg_11_ ( .D(N483), .CK(clk), .RN(rstn), .Q(y2_tmp[11]) );
  DFFRHQX1 y0_tmp_reg_11_ ( .D(N384), .CK(clk), .RN(rstn), .Q(y0_tmp[11]) );
  DFFRHQX1 y3_tmp_reg_11_ ( .D(N557), .CK(clk), .RN(rstn), .Q(y3_tmp[11]) );
  DFFRHQX1 mode_delay2_reg_1_ ( .D(mode_delay1[1]), .CK(clk), .RN(rstn), .Q(
        mode_delay2[1]) );
  DFFRHQX1 mode_delay2_reg_0_ ( .D(mode_delay1[0]), .CK(clk), .RN(rstn), .Q(
        mode_delay2[0]) );
  DFFRHQX1 x1_o1_tmp_reg_21_ ( .D(N30), .CK(clk), .RN(rstn), .Q(x1_o1_tmp[21])
         );
  DFFRHQX1 x1_o1_tmp_reg_20_ ( .D(N29), .CK(clk), .RN(rstn), .Q(x1_o1_tmp[20])
         );
  DFFRHQX1 x1_o1_tmp_reg_19_ ( .D(N28), .CK(clk), .RN(rstn), .Q(x1_o1_tmp[19])
         );
  DFFRHQX1 x1_o1_tmp_reg_18_ ( .D(N27), .CK(clk), .RN(rstn), .Q(x1_o1_tmp[18])
         );
  DFFRHQX1 x1_o1_tmp_reg_17_ ( .D(N26), .CK(clk), .RN(rstn), .Q(x1_o1_tmp[17])
         );
  DFFRHQX1 x1_o1_tmp_reg_16_ ( .D(N25), .CK(clk), .RN(rstn), .Q(x1_o1_tmp[16])
         );
  DFFRHQX1 x1_o1_tmp_reg_15_ ( .D(N24), .CK(clk), .RN(rstn), .Q(x1_o1_tmp[15])
         );
  DFFRHQX1 x1_o1_tmp_reg_14_ ( .D(N23), .CK(clk), .RN(rstn), .Q(x1_o1_tmp[14])
         );
  DFFRHQX1 x1_o1_tmp_reg_13_ ( .D(N22), .CK(clk), .RN(rstn), .Q(x1_o1_tmp[13])
         );
  DFFRHQX1 x1_o1_tmp_reg_12_ ( .D(N21), .CK(clk), .RN(rstn), .Q(x1_o1_tmp[12])
         );
  DFFRHQX1 x1_o1_tmp_reg_11_ ( .D(N20), .CK(clk), .RN(rstn), .Q(x1_o1_tmp[11])
         );
  DFFRHQX1 x1_o1_tmp_reg_10_ ( .D(N19), .CK(clk), .RN(rstn), .Q(x1_o1_tmp[10])
         );
  DFFRHQX1 x1_o1_tmp_reg_9_ ( .D(N18), .CK(clk), .RN(rstn), .Q(x1_o1_tmp[9])
         );
  DFFRHQX1 x1_o1_tmp_reg_8_ ( .D(N17), .CK(clk), .RN(rstn), .Q(x1_o1_tmp[8])
         );
  DFFRHQX1 x1_o1_tmp_reg_7_ ( .D(N16), .CK(clk), .RN(rstn), .Q(x1_o1_tmp[7])
         );
  DFFRHQX1 x1_o1_tmp_reg_6_ ( .D(N15), .CK(clk), .RN(rstn), .Q(x1_o1_tmp[6])
         );
  DFFRHQX1 x1_o1_tmp_reg_5_ ( .D(N14), .CK(clk), .RN(rstn), .Q(x1_o1_tmp[5])
         );
  DFFRHQX1 x3_o0_tmp_reg_21_ ( .D(N52), .CK(clk), .RN(rstn), .Q(x3_o0_tmp[21])
         );
  DFFRHQX1 x3_o0_tmp_reg_20_ ( .D(N51), .CK(clk), .RN(rstn), .Q(x3_o0_tmp[20])
         );
  DFFRHQX1 x3_o0_tmp_reg_19_ ( .D(N50), .CK(clk), .RN(rstn), .Q(x3_o0_tmp[19])
         );
  DFFRHQX1 x3_o0_tmp_reg_18_ ( .D(N49), .CK(clk), .RN(rstn), .Q(x3_o0_tmp[18])
         );
  DFFRHQX1 x3_o0_tmp_reg_17_ ( .D(N48), .CK(clk), .RN(rstn), .Q(x3_o0_tmp[17])
         );
  DFFRHQX1 x3_o0_tmp_reg_16_ ( .D(N47), .CK(clk), .RN(rstn), .Q(x3_o0_tmp[16])
         );
  DFFRHQX1 x3_o0_tmp_reg_15_ ( .D(N46), .CK(clk), .RN(rstn), .Q(x3_o0_tmp[15])
         );
  DFFRHQX1 x3_o0_tmp_reg_14_ ( .D(N45), .CK(clk), .RN(rstn), .Q(x3_o0_tmp[14])
         );
  DFFRHQX1 x3_o0_tmp_reg_13_ ( .D(N44), .CK(clk), .RN(rstn), .Q(x3_o0_tmp[13])
         );
  DFFRHQX1 x3_o0_tmp_reg_12_ ( .D(N43), .CK(clk), .RN(rstn), .Q(x3_o0_tmp[12])
         );
  DFFRHQX1 x3_o0_tmp_reg_11_ ( .D(N42), .CK(clk), .RN(rstn), .Q(x3_o0_tmp[11])
         );
  DFFRHQX1 x3_o0_tmp_reg_10_ ( .D(N41), .CK(clk), .RN(rstn), .Q(x3_o0_tmp[10])
         );
  DFFRHQX1 x3_o0_tmp_reg_9_ ( .D(N40), .CK(clk), .RN(rstn), .Q(x3_o0_tmp[9])
         );
  DFFRHQX1 x3_o0_tmp_reg_8_ ( .D(N39), .CK(clk), .RN(rstn), .Q(x3_o0_tmp[8])
         );
  DFFRHQX1 x3_o0_tmp_reg_7_ ( .D(N38), .CK(clk), .RN(rstn), .Q(x3_o0_tmp[7])
         );
  DFFRHQX1 x3_o0_tmp_reg_6_ ( .D(N37), .CK(clk), .RN(rstn), .Q(x3_o0_tmp[6])
         );
  DFFRHQX1 x3_o0_tmp_reg_5_ ( .D(N36), .CK(clk), .RN(rstn), .Q(x3_o0_tmp[5])
         );
  DFFRHQX1 mode_delay1_reg_1_ ( .D(mode[1]), .CK(clk), .RN(rstn), .Q(
        mode_delay1[1]) );
  DFFRHQX1 mode_delay1_reg_0_ ( .D(mode[0]), .CK(clk), .RN(rstn), .Q(
        mode_delay1[0]) );
  DFFRHQX1 idct4_ready_delay3_reg ( .D(idct4_ready_delay2), .CK(clk), .RN(rstn), .Q(idct4_ready_delay3) );
  DFFRHQX1 x1_o1_tmp_reg_4_ ( .D(x1[2]), .CK(clk), .RN(rstn), .Q(x1_o1_tmp[4])
         );
  DFFRHQX1 x1_o1_tmp_reg_3_ ( .D(x1[1]), .CK(clk), .RN(rstn), .Q(x1_o1_tmp[3])
         );
  DFFRHQX1 x1_o1_tmp_reg_2_ ( .D(x1[0]), .CK(clk), .RN(rstn), .Q(x1_o1_tmp[2])
         );
  DFFRHQX1 x2_e_tmp_reg_21_ ( .D(x2[15]), .CK(clk), .RN(rstn), .Q(x2_e_tmp[21]) );
  DFFRHQX1 x2_e_tmp_reg_20_ ( .D(x2[14]), .CK(clk), .RN(rstn), .Q(x2_e_tmp[20]) );
  DFFRHQX1 x2_e_tmp_reg_19_ ( .D(x2[13]), .CK(clk), .RN(rstn), .Q(x2_e_tmp[19]) );
  DFFRHQX1 x2_e_tmp_reg_18_ ( .D(x2[12]), .CK(clk), .RN(rstn), .Q(x2_e_tmp[18]) );
  DFFRHQX1 x2_e_tmp_reg_17_ ( .D(x2[11]), .CK(clk), .RN(rstn), .Q(x2_e_tmp[17]) );
  DFFRHQX1 x2_e_tmp_reg_16_ ( .D(x2[10]), .CK(clk), .RN(rstn), .Q(x2_e_tmp[16]) );
  DFFRHQX1 x2_e_tmp_reg_15_ ( .D(x2[9]), .CK(clk), .RN(rstn), .Q(x2_e_tmp[15])
         );
  DFFRHQX1 x2_e_tmp_reg_14_ ( .D(x2[8]), .CK(clk), .RN(rstn), .Q(x2_e_tmp[14])
         );
  DFFRHQX1 x2_e_tmp_reg_13_ ( .D(x2[7]), .CK(clk), .RN(rstn), .Q(x2_e_tmp[13])
         );
  DFFRHQX1 x2_e_tmp_reg_12_ ( .D(x2[6]), .CK(clk), .RN(rstn), .Q(x2_e_tmp[12])
         );
  DFFRHQX1 x2_e_tmp_reg_11_ ( .D(x2[5]), .CK(clk), .RN(rstn), .Q(x2_e_tmp[11])
         );
  DFFRHQX1 x2_e_tmp_reg_10_ ( .D(x2[4]), .CK(clk), .RN(rstn), .Q(x2_e_tmp[10])
         );
  DFFRHQX1 x2_e_tmp_reg_9_ ( .D(x2[3]), .CK(clk), .RN(rstn), .Q(x2_e_tmp[9])
         );
  DFFRHQX1 x2_e_tmp_reg_8_ ( .D(x2[2]), .CK(clk), .RN(rstn), .Q(x2_e_tmp[8])
         );
  DFFRHQX1 x2_e_tmp_reg_7_ ( .D(x2[1]), .CK(clk), .RN(rstn), .Q(x2_e_tmp[7])
         );
  DFFRHQX1 x2_e_tmp_reg_6_ ( .D(x2[0]), .CK(clk), .RN(rstn), .Q(x2_e_tmp[6])
         );
  DFFRHQX1 x0_e_tmp_reg_21_ ( .D(x0[15]), .CK(clk), .RN(rstn), .Q(x0_e_tmp[21]) );
  DFFRHQX1 x0_e_tmp_reg_20_ ( .D(x0[14]), .CK(clk), .RN(rstn), .Q(x0_e_tmp[20]) );
  DFFRHQX1 x0_e_tmp_reg_19_ ( .D(x0[13]), .CK(clk), .RN(rstn), .Q(x0_e_tmp[19]) );
  DFFRHQX1 x0_e_tmp_reg_18_ ( .D(x0[12]), .CK(clk), .RN(rstn), .Q(x0_e_tmp[18]) );
  DFFRHQX1 x0_e_tmp_reg_17_ ( .D(x0[11]), .CK(clk), .RN(rstn), .Q(x0_e_tmp[17]) );
  DFFRHQX1 x0_e_tmp_reg_16_ ( .D(x0[10]), .CK(clk), .RN(rstn), .Q(x0_e_tmp[16]) );
  DFFRHQX1 x0_e_tmp_reg_15_ ( .D(x0[9]), .CK(clk), .RN(rstn), .Q(x0_e_tmp[15])
         );
  DFFRHQX1 x0_e_tmp_reg_14_ ( .D(x0[8]), .CK(clk), .RN(rstn), .Q(x0_e_tmp[14])
         );
  DFFRHQX1 x0_e_tmp_reg_13_ ( .D(x0[7]), .CK(clk), .RN(rstn), .Q(x0_e_tmp[13])
         );
  DFFRHQX1 x0_e_tmp_reg_12_ ( .D(x0[6]), .CK(clk), .RN(rstn), .Q(x0_e_tmp[12])
         );
  DFFRHQX1 x0_e_tmp_reg_11_ ( .D(x0[5]), .CK(clk), .RN(rstn), .Q(x0_e_tmp[11])
         );
  DFFRHQX1 x0_e_tmp_reg_10_ ( .D(x0[4]), .CK(clk), .RN(rstn), .Q(x0_e_tmp[10])
         );
  DFFRHQX1 x0_e_tmp_reg_9_ ( .D(x0[3]), .CK(clk), .RN(rstn), .Q(x0_e_tmp[9])
         );
  DFFRHQX1 x0_e_tmp_reg_8_ ( .D(x0[2]), .CK(clk), .RN(rstn), .Q(x0_e_tmp[8])
         );
  DFFRHQX1 x0_e_tmp_reg_7_ ( .D(x0[1]), .CK(clk), .RN(rstn), .Q(x0_e_tmp[7])
         );
  DFFRHQX1 x0_e_tmp_reg_6_ ( .D(x0[0]), .CK(clk), .RN(rstn), .Q(x0_e_tmp[6])
         );
  DFFRHQX1 x3_o0_tmp_reg_4_ ( .D(x3[2]), .CK(clk), .RN(rstn), .Q(x3_o0_tmp[4])
         );
  DFFRHQX1 x3_o0_tmp_reg_3_ ( .D(x3[1]), .CK(clk), .RN(rstn), .Q(x3_o0_tmp[3])
         );
  DFFRHQX1 x3_o0_tmp_reg_2_ ( .D(x3[0]), .CK(clk), .RN(rstn), .Q(x3_o0_tmp[2])
         );
  DFFRHQX1 idct4_ready_delay1_reg ( .D(start), .CK(clk), .RN(rstn), .Q(
        idct4_ready_delay1) );
  DFFRHQX1 idct4_ready_delay2_reg ( .D(idct4_ready_delay1), .CK(clk), .RN(rstn), .Q(idct4_ready_delay2) );
  INVX1 U3 ( .A(n36), .Y(n20) );
  INVX1 U4 ( .A(n36), .Y(n22) );
  INVX1 U5 ( .A(n37), .Y(n19) );
  INVX1 U6 ( .A(n13), .Y(n36) );
  INVX1 U7 ( .A(n12), .Y(n33) );
  INVX1 U8 ( .A(n4), .Y(n29) );
  INVX1 U9 ( .A(n4), .Y(n27) );
  INVX1 U10 ( .A(n37), .Y(n21) );
  INVX1 U11 ( .A(n3), .Y(n24) );
  INVX1 U15 ( .A(n2), .Y(n25) );
  INVX1 U18 ( .A(n13), .Y(n35) );
  INVX1 U19 ( .A(n13), .Y(n34) );
  INVX1 U20 ( .A(n2), .Y(n26) );
  INVX1 U21 ( .A(n11), .Y(n31) );
  INVX1 U22 ( .A(n8), .Y(n30) );
  INVX1 U23 ( .A(n12), .Y(n32) );
  INVX1 U24 ( .A(n4), .Y(n28) );
  INVX1 U25 ( .A(n1), .Y(n23) );
  INVX1 U26 ( .A(n15), .Y(n13) );
  INVX1 U27 ( .A(n15), .Y(n12) );
  INVX1 U28 ( .A(n16), .Y(n4) );
  INVX1 U29 ( .A(n14), .Y(n37) );
  INVX1 U30 ( .A(n15), .Y(n14) );
  INVX1 U31 ( .A(n16), .Y(n8) );
  INVX1 U32 ( .A(n17), .Y(n2) );
  INVX1 U33 ( .A(n16), .Y(n11) );
  INVX1 U34 ( .A(n17), .Y(n3) );
  INVX1 U35 ( .A(n196), .Y(n15) );
  INVX1 U36 ( .A(n196), .Y(n16) );
  INVX1 U37 ( .A(n18), .Y(n1) );
  INVX1 U38 ( .A(n196), .Y(n18) );
  INVX1 U39 ( .A(n196), .Y(n17) );
  NOR2X1 U40 ( .A(mode_delay2[0]), .B(mode_delay2[1]), .Y(n196) );
  INVX1 U41 ( .A(n204), .Y(y3[1]) );
  AOI22X1 U42 ( .A0(N614), .A1(n19), .B0(y3_tmp[1]), .B1(n25), .Y(n204) );
  INVX1 U43 ( .A(n223), .Y(y2[0]) );
  AOI22X1 U44 ( .A0(N599), .A1(n20), .B0(y2_tmp[0]), .B1(n33), .Y(n223) );
  INVX1 U45 ( .A(n209), .Y(y3[0]) );
  AOI22X1 U46 ( .A0(N613), .A1(n19), .B0(y3_tmp[0]), .B1(n29), .Y(n209) );
  INVX1 U47 ( .A(n251), .Y(y0[0]) );
  AOI22X1 U48 ( .A0(N571), .A1(n19), .B0(y0_tmp[0]), .B1(n23), .Y(n251) );
  INVX1 U49 ( .A(n237), .Y(y1[0]) );
  AOI22X1 U50 ( .A0(N585), .A1(n22), .B0(y1_tmp[0]), .B1(n27), .Y(n237) );
  INVX1 U51 ( .A(n218), .Y(y2[1]) );
  AOI22X1 U52 ( .A0(N600), .A1(n20), .B0(y2_tmp[1]), .B1(n35), .Y(n218) );
  INVX1 U53 ( .A(n217), .Y(y2[2]) );
  AOI22X1 U54 ( .A0(N601), .A1(n20), .B0(y2_tmp[2]), .B1(n35), .Y(n217) );
  INVX1 U55 ( .A(n232), .Y(y1[1]) );
  AOI22X1 U56 ( .A0(N586), .A1(n22), .B0(y1_tmp[1]), .B1(n31), .Y(n232) );
  INVX1 U57 ( .A(n246), .Y(y0[1]) );
  AOI22X1 U58 ( .A0(N572), .A1(n22), .B0(y0_tmp[1]), .B1(n26), .Y(n246) );
  NAND2X1 U59 ( .A(N626), .B(n8), .Y(n205) );
  NAND2X1 U60 ( .A(N612), .B(n8), .Y(n219) );
  NAND2X1 U61 ( .A(N584), .B(n8), .Y(n247) );
  NAND2X1 U62 ( .A(N598), .B(n8), .Y(n233) );
  INVX1 U63 ( .A(n199), .Y(y3[6]) );
  AOI22X1 U64 ( .A0(N619), .A1(n19), .B0(y3_tmp[6]), .B1(n32), .Y(n199) );
  INVX1 U65 ( .A(n198), .Y(y3[7]) );
  AOI22X1 U66 ( .A0(N620), .A1(n19), .B0(y3_tmp[7]), .B1(n28), .Y(n198) );
  INVX1 U67 ( .A(n213), .Y(y2[6]) );
  AOI22X1 U68 ( .A0(N605), .A1(n20), .B0(y2_tmp[6]), .B1(n30), .Y(n213) );
  INVX1 U69 ( .A(n212), .Y(y2[7]) );
  AOI22X1 U70 ( .A0(N606), .A1(n20), .B0(y2_tmp[7]), .B1(n30), .Y(n212) );
  INVX1 U71 ( .A(n227), .Y(y1[6]) );
  AOI22X1 U72 ( .A0(N591), .A1(n21), .B0(y1_tmp[6]), .B1(n28), .Y(n227) );
  INVX1 U73 ( .A(n226), .Y(y1[7]) );
  AOI22X1 U74 ( .A0(N592), .A1(n21), .B0(y1_tmp[7]), .B1(n32), .Y(n226) );
  INVX1 U75 ( .A(n241), .Y(y0[6]) );
  AOI22X1 U76 ( .A0(N577), .A1(n22), .B0(y0_tmp[6]), .B1(n30), .Y(n241) );
  INVX1 U77 ( .A(n240), .Y(y0[7]) );
  AOI22X1 U78 ( .A0(N578), .A1(n21), .B0(y0_tmp[7]), .B1(n28), .Y(n240) );
  INVX1 U79 ( .A(n202), .Y(y3[3]) );
  AOI22X1 U80 ( .A0(N616), .A1(n19), .B0(y3_tmp[3]), .B1(n24), .Y(n202) );
  INVX1 U81 ( .A(n208), .Y(y3[10]) );
  AOI22X1 U82 ( .A0(N623), .A1(n19), .B0(y3_tmp[10]), .B1(n28), .Y(n208) );
  INVX1 U83 ( .A(n222), .Y(y2[10]) );
  AOI22X1 U84 ( .A0(N609), .A1(n20), .B0(y2_tmp[10]), .B1(n28), .Y(n222) );
  INVX1 U85 ( .A(n230), .Y(y1[3]) );
  AOI22X1 U86 ( .A0(N588), .A1(n21), .B0(y1_tmp[3]), .B1(n34), .Y(n230) );
  INVX1 U87 ( .A(n236), .Y(y1[10]) );
  AOI22X1 U88 ( .A0(N595), .A1(n22), .B0(y1_tmp[10]), .B1(n28), .Y(n236) );
  INVX1 U89 ( .A(n250), .Y(y0[10]) );
  AOI22X1 U90 ( .A0(N581), .A1(n22), .B0(y0_tmp[10]), .B1(n28), .Y(n250) );
  OAI2BB1X1 U91 ( .A0N(y3_tmp[13]), .A1N(n29), .B0(n205), .Y(y3[13]) );
  OAI2BB1X1 U92 ( .A0N(y3_tmp[14]), .A1N(n37), .B0(n205), .Y(y3[14]) );
  OAI2BB1X1 U93 ( .A0N(y3_tmp[15]), .A1N(n30), .B0(n205), .Y(y3[15]) );
  OAI2BB1X1 U94 ( .A0N(y2_tmp[13]), .A1N(n30), .B0(n219), .Y(y2[13]) );
  OAI2BB1X1 U95 ( .A0N(y2_tmp[14]), .A1N(n24), .B0(n219), .Y(y2[14]) );
  OAI2BB1X1 U96 ( .A0N(y2_tmp[15]), .A1N(n23), .B0(n219), .Y(y2[15]) );
  OAI2BB1X1 U97 ( .A0N(y1_tmp[13]), .A1N(n28), .B0(n233), .Y(y1[13]) );
  OAI2BB1X1 U98 ( .A0N(y1_tmp[14]), .A1N(n30), .B0(n233), .Y(y1[14]) );
  OAI2BB1X1 U99 ( .A0N(y1_tmp[15]), .A1N(n28), .B0(n233), .Y(y1[15]) );
  OAI2BB1X1 U100 ( .A0N(y0_tmp[13]), .A1N(n37), .B0(n247), .Y(y0[13]) );
  OAI2BB1X1 U101 ( .A0N(y0_tmp[14]), .A1N(n34), .B0(n247), .Y(y0[14]) );
  OAI2BB1X1 U102 ( .A0N(y0_tmp[15]), .A1N(n35), .B0(n247), .Y(y0[15]) );
  INVX1 U103 ( .A(n203), .Y(y3[2]) );
  AOI22X1 U104 ( .A0(N615), .A1(n19), .B0(y3_tmp[2]), .B1(n24), .Y(n203) );
  INVX1 U105 ( .A(n201), .Y(y3[4]) );
  AOI22X1 U106 ( .A0(N617), .A1(n19), .B0(y3_tmp[4]), .B1(n32), .Y(n201) );
  INVX1 U107 ( .A(n200), .Y(y3[5]) );
  AOI22X1 U108 ( .A0(N618), .A1(n19), .B0(y3_tmp[5]), .B1(n23), .Y(n200) );
  INVX1 U109 ( .A(n197), .Y(y3[8]) );
  AOI22X1 U110 ( .A0(N621), .A1(n19), .B0(y3_tmp[8]), .B1(n28), .Y(n197) );
  INVX1 U111 ( .A(n195), .Y(y3[9]) );
  AOI22X1 U112 ( .A0(N622), .A1(n21), .B0(y3_tmp[9]), .B1(n28), .Y(n195) );
  INVX1 U113 ( .A(n207), .Y(y3[11]) );
  AOI22X1 U114 ( .A0(N624), .A1(n19), .B0(y3_tmp[11]), .B1(n28), .Y(n207) );
  INVX1 U115 ( .A(n206), .Y(y3[12]) );
  AOI22X1 U116 ( .A0(N625), .A1(n19), .B0(y3_tmp[12]), .B1(n25), .Y(n206) );
  INVX1 U117 ( .A(n216), .Y(y2[3]) );
  AOI22X1 U118 ( .A0(N602), .A1(n20), .B0(y2_tmp[3]), .B1(n34), .Y(n216) );
  INVX1 U119 ( .A(n215), .Y(y2[4]) );
  AOI22X1 U120 ( .A0(N603), .A1(n20), .B0(y2_tmp[4]), .B1(n32), .Y(n215) );
  INVX1 U121 ( .A(n214), .Y(y2[5]) );
  AOI22X1 U122 ( .A0(N604), .A1(n20), .B0(y2_tmp[5]), .B1(n28), .Y(n214) );
  INVX1 U123 ( .A(n211), .Y(y2[8]) );
  AOI22X1 U124 ( .A0(N607), .A1(n20), .B0(y2_tmp[8]), .B1(n28), .Y(n211) );
  INVX1 U125 ( .A(n210), .Y(y2[9]) );
  AOI22X1 U126 ( .A0(N608), .A1(n20), .B0(y2_tmp[9]), .B1(n28), .Y(n210) );
  INVX1 U127 ( .A(n221), .Y(y2[11]) );
  AOI22X1 U128 ( .A0(N610), .A1(n20), .B0(y2_tmp[11]), .B1(n28), .Y(n221) );
  INVX1 U129 ( .A(n220), .Y(y2[12]) );
  AOI22X1 U130 ( .A0(N611), .A1(n20), .B0(y2_tmp[12]), .B1(n34), .Y(n220) );
  INVX1 U131 ( .A(n231), .Y(y1[2]) );
  AOI22X1 U132 ( .A0(N587), .A1(n21), .B0(y1_tmp[2]), .B1(n31), .Y(n231) );
  INVX1 U133 ( .A(n229), .Y(y1[4]) );
  AOI22X1 U134 ( .A0(N589), .A1(n21), .B0(y1_tmp[4]), .B1(n32), .Y(n229) );
  INVX1 U135 ( .A(n228), .Y(y1[5]) );
  AOI22X1 U136 ( .A0(N590), .A1(n21), .B0(y1_tmp[5]), .B1(n32), .Y(n228) );
  INVX1 U137 ( .A(n225), .Y(y1[8]) );
  AOI22X1 U138 ( .A0(N593), .A1(n21), .B0(y1_tmp[8]), .B1(n32), .Y(n225) );
  INVX1 U139 ( .A(n224), .Y(y1[9]) );
  AOI22X1 U140 ( .A0(N594), .A1(n21), .B0(y1_tmp[9]), .B1(n33), .Y(n224) );
  INVX1 U141 ( .A(n235), .Y(y1[11]) );
  AOI22X1 U142 ( .A0(N596), .A1(n22), .B0(y1_tmp[11]), .B1(n28), .Y(n235) );
  INVX1 U143 ( .A(n234), .Y(y1[12]) );
  AOI22X1 U144 ( .A0(N597), .A1(n21), .B0(y1_tmp[12]), .B1(n29), .Y(n234) );
  INVX1 U145 ( .A(n245), .Y(y0[2]) );
  AOI22X1 U146 ( .A0(N573), .A1(n21), .B0(y0_tmp[2]), .B1(n26), .Y(n245) );
  INVX1 U147 ( .A(n244), .Y(y0[3]) );
  AOI22X1 U148 ( .A0(N574), .A1(n22), .B0(y0_tmp[3]), .B1(n34), .Y(n244) );
  INVX1 U149 ( .A(n243), .Y(y0[4]) );
  AOI22X1 U150 ( .A0(N575), .A1(n22), .B0(y0_tmp[4]), .B1(n32), .Y(n243) );
  INVX1 U151 ( .A(n242), .Y(y0[5]) );
  AOI22X1 U152 ( .A0(N576), .A1(n21), .B0(y0_tmp[5]), .B1(n28), .Y(n242) );
  INVX1 U153 ( .A(n239), .Y(y0[8]) );
  AOI22X1 U154 ( .A0(N579), .A1(n22), .B0(y0_tmp[8]), .B1(n28), .Y(n239) );
  INVX1 U155 ( .A(n238), .Y(y0[9]) );
  AOI22X1 U156 ( .A0(N580), .A1(n22), .B0(y0_tmp[9]), .B1(n27), .Y(n238) );
  INVX1 U157 ( .A(n249), .Y(y0[11]) );
  AOI22X1 U158 ( .A0(N582), .A1(n22), .B0(y0_tmp[11]), .B1(n28), .Y(n249) );
  INVX1 U159 ( .A(n248), .Y(y0[12]) );
  AOI22X1 U160 ( .A0(N583), .A1(n22), .B0(y0_tmp[12]), .B1(n30), .Y(n248) );
  OAI2BB1X1 U161 ( .A0N(y3_tmp[16]), .A1N(n28), .B0(n205), .Y(y3[16]) );
  OAI2BB1X1 U162 ( .A0N(y3_tmp[17]), .A1N(n31), .B0(n205), .Y(y3[17]) );
  OAI2BB1X1 U163 ( .A0N(y3_tmp[18]), .A1N(n32), .B0(n205), .Y(y3[18]) );
  OAI2BB1X1 U164 ( .A0N(y3_tmp[19]), .A1N(n28), .B0(n205), .Y(y3[19]) );
  OAI2BB1X1 U165 ( .A0N(y2_tmp[16]), .A1N(n30), .B0(n219), .Y(y2[16]) );
  OAI2BB1X1 U166 ( .A0N(y2_tmp[17]), .A1N(n28), .B0(n219), .Y(y2[17]) );
  OAI2BB1X1 U167 ( .A0N(y2_tmp[18]), .A1N(n28), .B0(n219), .Y(y2[18]) );
  OAI2BB1X1 U168 ( .A0N(y2_tmp[19]), .A1N(n28), .B0(n219), .Y(y2[19]) );
  OAI2BB1X1 U169 ( .A0N(y0_tmp[16]), .A1N(n33), .B0(n247), .Y(y0[16]) );
  OAI2BB1X1 U170 ( .A0N(y0_tmp[17]), .A1N(n28), .B0(n247), .Y(y0[17]) );
  OAI2BB1X1 U171 ( .A0N(y0_tmp[18]), .A1N(n28), .B0(n247), .Y(y0[18]) );
  OAI2BB1X1 U172 ( .A0N(y0_tmp[19]), .A1N(n27), .B0(n247), .Y(y0[19]) );
  OAI2BB1X1 U173 ( .A0N(y1_tmp[16]), .A1N(n26), .B0(n233), .Y(y1[16]) );
  OAI2BB1X1 U174 ( .A0N(y1_tmp[17]), .A1N(n28), .B0(n233), .Y(y1[17]) );
  OAI2BB1X1 U175 ( .A0N(y1_tmp[18]), .A1N(n25), .B0(n233), .Y(y1[18]) );
  OAI2BB1X1 U176 ( .A0N(y1_tmp[19]), .A1N(n28), .B0(n233), .Y(y1[19]) );
  INVX1 U177 ( .A(o0[0]), .Y(n108) );
  INVX1 U178 ( .A(o1[0]), .Y(n84) );
  INVX1 U179 ( .A(x3_o1[0]), .Y(n60) );
  INVX1 U180 ( .A(o0[1]), .Y(n107) );
  INVX1 U181 ( .A(o1[1]), .Y(n83) );
  INVX1 U182 ( .A(o0[22]), .Y(n86) );
  INVX1 U183 ( .A(o0[21]), .Y(n87) );
  INVX1 U184 ( .A(o0[20]), .Y(n88) );
  INVX1 U185 ( .A(o0[19]), .Y(n89) );
  INVX1 U186 ( .A(o0[18]), .Y(n90) );
  INVX1 U187 ( .A(o0[17]), .Y(n91) );
  INVX1 U188 ( .A(o0[16]), .Y(n92) );
  INVX1 U189 ( .A(o0[15]), .Y(n93) );
  INVX1 U190 ( .A(o0[14]), .Y(n94) );
  INVX1 U191 ( .A(o0[13]), .Y(n95) );
  INVX1 U192 ( .A(o0[12]), .Y(n96) );
  INVX1 U193 ( .A(o0[11]), .Y(n97) );
  INVX1 U194 ( .A(o0[10]), .Y(n98) );
  INVX1 U195 ( .A(o0[9]), .Y(n99) );
  INVX1 U196 ( .A(o0[8]), .Y(n100) );
  INVX1 U197 ( .A(o0[7]), .Y(n101) );
  INVX1 U198 ( .A(o0[6]), .Y(n102) );
  INVX1 U199 ( .A(o0[5]), .Y(n103) );
  INVX1 U200 ( .A(o0[4]), .Y(n104) );
  INVX1 U201 ( .A(o0[3]), .Y(n105) );
  INVX1 U202 ( .A(o0[2]), .Y(n106) );
  INVX1 U203 ( .A(o1[2]), .Y(n82) );
  INVX1 U204 ( .A(o1[3]), .Y(n81) );
  INVX1 U205 ( .A(o1[4]), .Y(n80) );
  INVX1 U206 ( .A(o1[5]), .Y(n79) );
  INVX1 U207 ( .A(o1[6]), .Y(n78) );
  INVX1 U208 ( .A(o1[7]), .Y(n77) );
  INVX1 U209 ( .A(o1[8]), .Y(n76) );
  INVX1 U210 ( .A(o1[9]), .Y(n75) );
  INVX1 U211 ( .A(o1[10]), .Y(n74) );
  INVX1 U212 ( .A(o1[11]), .Y(n73) );
  INVX1 U213 ( .A(o1[12]), .Y(n72) );
  INVX1 U214 ( .A(o1[13]), .Y(n71) );
  INVX1 U215 ( .A(o1[14]), .Y(n70) );
  INVX1 U216 ( .A(o1[15]), .Y(n69) );
  INVX1 U217 ( .A(o1[16]), .Y(n68) );
  INVX1 U218 ( .A(o1[17]), .Y(n67) );
  INVX1 U219 ( .A(o1[18]), .Y(n66) );
  INVX1 U220 ( .A(o1[19]), .Y(n65) );
  INVX1 U221 ( .A(o1[20]), .Y(n64) );
  INVX1 U222 ( .A(o1[21]), .Y(n63) );
  INVX1 U223 ( .A(o1[22]), .Y(n62) );
  INVX1 U224 ( .A(x3_o1[2]), .Y(n58) );
  INVX1 U225 ( .A(x3_o1[3]), .Y(n57) );
  INVX1 U226 ( .A(x3_o1[4]), .Y(n56) );
  INVX1 U227 ( .A(x3_o1[5]), .Y(n55) );
  INVX1 U228 ( .A(x3_o1[6]), .Y(n54) );
  INVX1 U229 ( .A(x3_o1[7]), .Y(n53) );
  INVX1 U230 ( .A(x3_o1[8]), .Y(n52) );
  INVX1 U231 ( .A(x3_o1[9]), .Y(n51) );
  INVX1 U232 ( .A(x3_o1[10]), .Y(n50) );
  INVX1 U233 ( .A(x3_o1[11]), .Y(n49) );
  INVX1 U234 ( .A(x3_o1[12]), .Y(n48) );
  INVX1 U235 ( .A(x3_o1[13]), .Y(n47) );
  INVX1 U236 ( .A(x3_o1[14]), .Y(n46) );
  INVX1 U237 ( .A(x3_o1[15]), .Y(n45) );
  INVX1 U238 ( .A(x3_o1[16]), .Y(n44) );
  INVX1 U239 ( .A(x3_o1[17]), .Y(n43) );
  INVX1 U240 ( .A(x3_o1[18]), .Y(n42) );
  INVX1 U241 ( .A(x3_o1[19]), .Y(n41) );
  INVX1 U242 ( .A(x3_o1[20]), .Y(n40) );
  INVX1 U243 ( .A(x3_o1[21]), .Y(n39) );
  INVX1 U244 ( .A(x3_o1[1]), .Y(n59) );
  ADDFX2 U245 ( .A(x1[1]), .B(x1[7]), .CI(add_85_carry_7_), .CO(
        add_85_carry_8_), .S(N60) );
  ADDFX2 U246 ( .A(x3[1]), .B(x3[7]), .CI(add_87_carry_7_), .CO(
        add_87_carry_8_), .S(N104) );
  ADDFX2 U247 ( .A(x3[1]), .B(x3[4]), .CI(add_81_carry_6_), .CO(
        add_81_carry_7_), .S(N37) );
  ADDFX2 U248 ( .A(x1[1]), .B(x1[4]), .CI(add_80_carry_6_), .CO(
        add_80_carry_7_), .S(N15) );
  ADDFX2 U249 ( .A(x1[1]), .B(x1[4]), .CI(add_86_carry_5_), .CO(
        add_86_carry_6_), .S(N81) );
  ADDFX2 U250 ( .A(x3[1]), .B(x3[4]), .CI(add_88_carry_5_), .CO(
        add_88_carry_6_), .S(N125) );
  ADDFX2 U251 ( .A(x0_e[7]), .B(add_1_root_add_112_2_B_7_), .CI(
        add_1_root_add_112_2_carry[7]), .CO(add_1_root_add_112_2_carry[8]), 
        .S(N262) );
  INVX1 U252 ( .A(x2_e[7]), .Y(add_1_root_add_112_2_B_7_) );
  ADDFX2 U253 ( .A(x0_e[7]), .B(x2_e[7]), .CI(add_111_carry[7]), .CO(
        add_111_carry[8]), .S(N194) );
  ADDFX2 U254 ( .A(x0_e[8]), .B(x2_e[8]), .CI(add_111_carry[8]), .CO(
        add_111_carry[9]), .S(N195) );
  ADDFX2 U255 ( .A(x0_e[9]), .B(x2_e[9]), .CI(add_111_carry[9]), .CO(
        add_111_carry[10]), .S(N196) );
  ADDFX2 U256 ( .A(x0_e[10]), .B(x2_e[10]), .CI(add_111_carry[10]), .CO(
        add_111_carry[11]), .S(N197) );
  ADDFX2 U257 ( .A(x0_e[11]), .B(x2_e[11]), .CI(add_111_carry[11]), .CO(
        add_111_carry[12]), .S(N198) );
  ADDFX2 U258 ( .A(x0_e[12]), .B(x2_e[12]), .CI(add_111_carry[12]), .CO(
        add_111_carry[13]), .S(N199) );
  ADDFX2 U259 ( .A(x0_e[13]), .B(x2_e[13]), .CI(add_111_carry[13]), .CO(
        add_111_carry[14]), .S(N200) );
  ADDFX2 U260 ( .A(x0_e[14]), .B(x2_e[14]), .CI(add_111_carry[14]), .CO(
        add_111_carry[15]), .S(N201) );
  ADDFX2 U261 ( .A(x0_e[15]), .B(x2_e[15]), .CI(add_111_carry[15]), .CO(
        add_111_carry[16]), .S(N202) );
  ADDFX2 U262 ( .A(x0_e[16]), .B(x2_e[16]), .CI(add_111_carry[16]), .CO(
        add_111_carry[17]), .S(N203) );
  ADDFX2 U263 ( .A(x0_e[17]), .B(x2_e[17]), .CI(add_111_carry[17]), .CO(
        add_111_carry[18]), .S(N204) );
  ADDFX2 U264 ( .A(x0_e[18]), .B(x2_e[18]), .CI(add_111_carry[18]), .CO(
        add_111_carry[19]), .S(N205) );
  ADDFX2 U265 ( .A(x0_e[19]), .B(x2_e[19]), .CI(add_111_carry[19]), .CO(
        add_111_carry[20]), .S(N206) );
  ADDFX2 U266 ( .A(x0_e[20]), .B(x2_e[20]), .CI(add_111_carry[20]), .CO(
        add_111_carry[21]), .S(N207) );
  ADDFX2 U267 ( .A(x0_e[21]), .B(x2_e[21]), .CI(add_111_carry[21]), .CO(
        add_111_carry[22]), .S(N208) );
  ADDFX2 U268 ( .A(x0_e[8]), .B(add_1_root_add_112_2_B_8_), .CI(
        add_1_root_add_112_2_carry[8]), .CO(add_1_root_add_112_2_carry[9]), 
        .S(N263) );
  INVX1 U269 ( .A(x2_e[8]), .Y(add_1_root_add_112_2_B_8_) );
  ADDFX2 U270 ( .A(x0_e[9]), .B(add_1_root_add_112_2_B_9_), .CI(
        add_1_root_add_112_2_carry[9]), .CO(add_1_root_add_112_2_carry[10]), 
        .S(N264) );
  INVX1 U271 ( .A(x2_e[9]), .Y(add_1_root_add_112_2_B_9_) );
  ADDFX2 U272 ( .A(x0_e[10]), .B(add_1_root_add_112_2_B_10_), .CI(
        add_1_root_add_112_2_carry[10]), .CO(add_1_root_add_112_2_carry[11]), 
        .S(N265) );
  INVX1 U273 ( .A(x2_e[10]), .Y(add_1_root_add_112_2_B_10_) );
  ADDFX2 U274 ( .A(x0_e[11]), .B(add_1_root_add_112_2_B_11_), .CI(
        add_1_root_add_112_2_carry[11]), .CO(add_1_root_add_112_2_carry[12]), 
        .S(N266) );
  INVX1 U275 ( .A(x2_e[11]), .Y(add_1_root_add_112_2_B_11_) );
  ADDFX2 U276 ( .A(x0_e[12]), .B(add_1_root_add_112_2_B_12_), .CI(
        add_1_root_add_112_2_carry[12]), .CO(add_1_root_add_112_2_carry[13]), 
        .S(N267) );
  INVX1 U277 ( .A(x2_e[12]), .Y(add_1_root_add_112_2_B_12_) );
  ADDFX2 U278 ( .A(x0_e[13]), .B(add_1_root_add_112_2_B_13_), .CI(
        add_1_root_add_112_2_carry[13]), .CO(add_1_root_add_112_2_carry[14]), 
        .S(N268) );
  INVX1 U279 ( .A(x2_e[13]), .Y(add_1_root_add_112_2_B_13_) );
  ADDFX2 U280 ( .A(x0_e[14]), .B(add_1_root_add_112_2_B_14_), .CI(
        add_1_root_add_112_2_carry[14]), .CO(add_1_root_add_112_2_carry[15]), 
        .S(N269) );
  INVX1 U281 ( .A(x2_e[14]), .Y(add_1_root_add_112_2_B_14_) );
  ADDFX2 U282 ( .A(x0_e[15]), .B(add_1_root_add_112_2_B_15_), .CI(
        add_1_root_add_112_2_carry[15]), .CO(add_1_root_add_112_2_carry[16]), 
        .S(N270) );
  INVX1 U283 ( .A(x2_e[15]), .Y(add_1_root_add_112_2_B_15_) );
  ADDFX2 U284 ( .A(x0_e[16]), .B(add_1_root_add_112_2_B_16_), .CI(
        add_1_root_add_112_2_carry[16]), .CO(add_1_root_add_112_2_carry[17]), 
        .S(N271) );
  INVX1 U285 ( .A(x2_e[16]), .Y(add_1_root_add_112_2_B_16_) );
  ADDFX2 U286 ( .A(x0_e[17]), .B(add_1_root_add_112_2_B_17_), .CI(
        add_1_root_add_112_2_carry[17]), .CO(add_1_root_add_112_2_carry[18]), 
        .S(N272) );
  INVX1 U287 ( .A(x2_e[17]), .Y(add_1_root_add_112_2_B_17_) );
  ADDFX2 U288 ( .A(x0_e[18]), .B(add_1_root_add_112_2_B_18_), .CI(
        add_1_root_add_112_2_carry[18]), .CO(add_1_root_add_112_2_carry[19]), 
        .S(N273) );
  INVX1 U289 ( .A(x2_e[18]), .Y(add_1_root_add_112_2_B_18_) );
  ADDFX2 U290 ( .A(x0_e[19]), .B(add_1_root_add_112_2_B_19_), .CI(
        add_1_root_add_112_2_carry[19]), .CO(add_1_root_add_112_2_carry[20]), 
        .S(N274) );
  INVX1 U291 ( .A(x2_e[19]), .Y(add_1_root_add_112_2_B_19_) );
  ADDFX2 U292 ( .A(x0_e[20]), .B(add_1_root_add_112_2_B_20_), .CI(
        add_1_root_add_112_2_carry[20]), .CO(add_1_root_add_112_2_carry[21]), 
        .S(N275) );
  INVX1 U293 ( .A(x2_e[20]), .Y(add_1_root_add_112_2_B_20_) );
  ADDFX2 U294 ( .A(x0_e[21]), .B(add_1_root_add_112_2_B_21_), .CI(
        add_1_root_add_112_2_carry[21]), .CO(add_1_root_add_112_2_carry[22]), 
        .S(N276) );
  ADDFX2 U295 ( .A(x1[2]), .B(x1[8]), .CI(add_85_carry_8_), .CO(
        add_85_carry_9_), .S(N61) );
  ADDFX2 U296 ( .A(x1[3]), .B(x1[9]), .CI(add_85_carry_9_), .CO(
        add_85_carry_10_), .S(N62) );
  ADDFX2 U297 ( .A(x1[4]), .B(x1[10]), .CI(add_85_carry_10_), .CO(
        add_85_carry_11_), .S(N63) );
  ADDFX2 U298 ( .A(x1[5]), .B(x1[11]), .CI(add_85_carry_11_), .CO(
        add_85_carry_12_), .S(N64) );
  ADDFX2 U299 ( .A(x1[6]), .B(x1[12]), .CI(add_85_carry_12_), .CO(
        add_85_carry_13_), .S(N65) );
  ADDFX2 U300 ( .A(x1[7]), .B(x1[13]), .CI(add_85_carry_13_), .CO(
        add_85_carry_14_), .S(N66) );
  ADDFX2 U301 ( .A(x1[8]), .B(x1[14]), .CI(add_85_carry_14_), .CO(
        add_85_carry_15_), .S(N67) );
  ADDFX2 U302 ( .A(x1[9]), .B(N30), .CI(add_85_carry_15_), .CO(
        add_85_carry_16_), .S(N68) );
  ADDFX2 U303 ( .A(x1[10]), .B(N30), .CI(add_85_carry_16_), .CO(
        add_85_carry_17_), .S(N69) );
  ADDFX2 U304 ( .A(x1[11]), .B(N30), .CI(add_85_carry_17_), .CO(
        add_85_carry_18_), .S(N70) );
  ADDFX2 U305 ( .A(x1[12]), .B(N30), .CI(add_85_carry_18_), .CO(
        add_85_carry_19_), .S(N71) );
  ADDFX2 U306 ( .A(x1[13]), .B(N30), .CI(add_85_carry_19_), .CO(
        add_85_carry_20_), .S(N72) );
  ADDFX2 U307 ( .A(x3[2]), .B(x3[5]), .CI(add_81_carry_7_), .CO(
        add_81_carry_8_), .S(N38) );
  ADDFX2 U308 ( .A(x3[3]), .B(x3[6]), .CI(add_81_carry_8_), .CO(
        add_81_carry_9_), .S(N39) );
  ADDFX2 U309 ( .A(x3[4]), .B(x3[7]), .CI(add_81_carry_9_), .CO(
        add_81_carry_10_), .S(N40) );
  ADDFX2 U310 ( .A(x3[5]), .B(x3[8]), .CI(add_81_carry_10_), .CO(
        add_81_carry_11_), .S(N41) );
  ADDFX2 U311 ( .A(x3[6]), .B(x3[9]), .CI(add_81_carry_11_), .CO(
        add_81_carry_12_), .S(N42) );
  ADDFX2 U312 ( .A(x3[7]), .B(x3[10]), .CI(add_81_carry_12_), .CO(
        add_81_carry_13_), .S(N43) );
  ADDFX2 U313 ( .A(x3[8]), .B(x3[11]), .CI(add_81_carry_13_), .CO(
        add_81_carry_14_), .S(N44) );
  ADDFX2 U314 ( .A(x3[9]), .B(x3[12]), .CI(add_81_carry_14_), .CO(
        add_81_carry_15_), .S(N45) );
  ADDFX2 U315 ( .A(x3[10]), .B(x3[13]), .CI(add_81_carry_15_), .CO(
        add_81_carry_16_), .S(N46) );
  ADDFX2 U316 ( .A(x3[11]), .B(x3[14]), .CI(add_81_carry_16_), .CO(
        add_81_carry_17_), .S(N47) );
  ADDFX2 U317 ( .A(x3[12]), .B(N52), .CI(add_81_carry_17_), .CO(
        add_81_carry_18_), .S(N48) );
  ADDFX2 U318 ( .A(x3[13]), .B(N52), .CI(add_81_carry_18_), .CO(
        add_81_carry_19_), .S(N49) );
  ADDFX2 U319 ( .A(x1[2]), .B(x1[5]), .CI(add_80_carry_7_), .CO(
        add_80_carry_8_), .S(N16) );
  ADDFX2 U320 ( .A(x1[3]), .B(x1[6]), .CI(add_80_carry_8_), .CO(
        add_80_carry_9_), .S(N17) );
  ADDFX2 U321 ( .A(x1[4]), .B(x1[7]), .CI(add_80_carry_9_), .CO(
        add_80_carry_10_), .S(N18) );
  ADDFX2 U322 ( .A(x1[5]), .B(x1[8]), .CI(add_80_carry_10_), .CO(
        add_80_carry_11_), .S(N19) );
  ADDFX2 U323 ( .A(x1[6]), .B(x1[9]), .CI(add_80_carry_11_), .CO(
        add_80_carry_12_), .S(N20) );
  ADDFX2 U324 ( .A(x1[7]), .B(x1[10]), .CI(add_80_carry_12_), .CO(
        add_80_carry_13_), .S(N21) );
  ADDFX2 U325 ( .A(x1[8]), .B(x1[11]), .CI(add_80_carry_13_), .CO(
        add_80_carry_14_), .S(N22) );
  ADDFX2 U326 ( .A(x1[9]), .B(x1[12]), .CI(add_80_carry_14_), .CO(
        add_80_carry_15_), .S(N23) );
  ADDFX2 U327 ( .A(x1[10]), .B(x1[13]), .CI(add_80_carry_15_), .CO(
        add_80_carry_16_), .S(N24) );
  ADDFX2 U328 ( .A(x1[11]), .B(x1[14]), .CI(add_80_carry_16_), .CO(
        add_80_carry_17_), .S(N25) );
  ADDFX2 U329 ( .A(x1[12]), .B(N30), .CI(add_80_carry_17_), .CO(
        add_80_carry_18_), .S(N26) );
  ADDFX2 U330 ( .A(x1[13]), .B(N30), .CI(add_80_carry_18_), .CO(
        add_80_carry_19_), .S(N27) );
  ADDFX2 U331 ( .A(x1[2]), .B(x1[5]), .CI(add_86_carry_6_), .CO(
        add_86_carry_7_), .S(N82) );
  ADDFX2 U332 ( .A(x1[3]), .B(x1[6]), .CI(add_86_carry_7_), .CO(
        add_86_carry_8_), .S(N83) );
  ADDFX2 U333 ( .A(x1[4]), .B(x1[7]), .CI(add_86_carry_8_), .CO(
        add_86_carry_9_), .S(N84) );
  ADDFX2 U334 ( .A(x1[5]), .B(x1[8]), .CI(add_86_carry_9_), .CO(
        add_86_carry_10_), .S(N85) );
  ADDFX2 U335 ( .A(x1[6]), .B(x1[9]), .CI(add_86_carry_10_), .CO(
        add_86_carry_11_), .S(N86) );
  ADDFX2 U336 ( .A(x1[7]), .B(x1[10]), .CI(add_86_carry_11_), .CO(
        add_86_carry_12_), .S(N87) );
  ADDFX2 U337 ( .A(x1[8]), .B(x1[11]), .CI(add_86_carry_12_), .CO(
        add_86_carry_13_), .S(N88) );
  ADDFX2 U338 ( .A(x1[9]), .B(x1[12]), .CI(add_86_carry_13_), .CO(
        add_86_carry_14_), .S(N89) );
  ADDFX2 U339 ( .A(x1[10]), .B(x1[13]), .CI(add_86_carry_14_), .CO(
        add_86_carry_15_), .S(N90) );
  ADDFX2 U340 ( .A(x1[11]), .B(x1[14]), .CI(add_86_carry_15_), .CO(
        add_86_carry_16_), .S(N91) );
  ADDFX2 U341 ( .A(x1[12]), .B(N30), .CI(add_86_carry_16_), .CO(
        add_86_carry_17_), .S(N92) );
  ADDFX2 U342 ( .A(x1[13]), .B(N30), .CI(add_86_carry_17_), .CO(
        add_86_carry_18_), .S(N93) );
  ADDFX2 U343 ( .A(x3[2]), .B(x3[8]), .CI(add_87_carry_8_), .CO(
        add_87_carry_9_), .S(N105) );
  ADDFX2 U344 ( .A(x3[3]), .B(x3[9]), .CI(add_87_carry_9_), .CO(
        add_87_carry_10_), .S(N106) );
  ADDFX2 U345 ( .A(x3[4]), .B(x3[10]), .CI(add_87_carry_10_), .CO(
        add_87_carry_11_), .S(N107) );
  ADDFX2 U346 ( .A(x3[5]), .B(x3[11]), .CI(add_87_carry_11_), .CO(
        add_87_carry_12_), .S(N108) );
  ADDFX2 U347 ( .A(x3[6]), .B(x3[12]), .CI(add_87_carry_12_), .CO(
        add_87_carry_13_), .S(N109) );
  ADDFX2 U348 ( .A(x3[7]), .B(x3[13]), .CI(add_87_carry_13_), .CO(
        add_87_carry_14_), .S(N110) );
  ADDFX2 U349 ( .A(x3[8]), .B(x3[14]), .CI(add_87_carry_14_), .CO(
        add_87_carry_15_), .S(N111) );
  ADDFX2 U350 ( .A(x3[9]), .B(N52), .CI(add_87_carry_15_), .CO(
        add_87_carry_16_), .S(N112) );
  ADDFX2 U351 ( .A(x3[10]), .B(N52), .CI(add_87_carry_16_), .CO(
        add_87_carry_17_), .S(N113) );
  ADDFX2 U352 ( .A(x3[11]), .B(N52), .CI(add_87_carry_17_), .CO(
        add_87_carry_18_), .S(N114) );
  ADDFX2 U353 ( .A(x3[12]), .B(N52), .CI(add_87_carry_18_), .CO(
        add_87_carry_19_), .S(N115) );
  ADDFX2 U354 ( .A(x3[13]), .B(N52), .CI(add_87_carry_19_), .CO(
        add_87_carry_20_), .S(N116) );
  ADDFX2 U355 ( .A(x3[2]), .B(x3[5]), .CI(add_88_carry_6_), .CO(
        add_88_carry_7_), .S(N126) );
  ADDFX2 U356 ( .A(x3[3]), .B(x3[6]), .CI(add_88_carry_7_), .CO(
        add_88_carry_8_), .S(N127) );
  ADDFX2 U357 ( .A(x3[4]), .B(x3[7]), .CI(add_88_carry_8_), .CO(
        add_88_carry_9_), .S(N128) );
  ADDFX2 U358 ( .A(x3[5]), .B(x3[8]), .CI(add_88_carry_9_), .CO(
        add_88_carry_10_), .S(N129) );
  ADDFX2 U359 ( .A(x3[6]), .B(x3[9]), .CI(add_88_carry_10_), .CO(
        add_88_carry_11_), .S(N130) );
  ADDFX2 U360 ( .A(x3[7]), .B(x3[10]), .CI(add_88_carry_11_), .CO(
        add_88_carry_12_), .S(N131) );
  ADDFX2 U361 ( .A(x3[8]), .B(x3[11]), .CI(add_88_carry_12_), .CO(
        add_88_carry_13_), .S(N132) );
  ADDFX2 U362 ( .A(x3[9]), .B(x3[12]), .CI(add_88_carry_13_), .CO(
        add_88_carry_14_), .S(N133) );
  ADDFX2 U363 ( .A(x3[10]), .B(x3[13]), .CI(add_88_carry_14_), .CO(
        add_88_carry_15_), .S(N134) );
  ADDFX2 U364 ( .A(x3[11]), .B(x3[14]), .CI(add_88_carry_15_), .CO(
        add_88_carry_16_), .S(N135) );
  ADDFX2 U365 ( .A(x3[12]), .B(N52), .CI(add_88_carry_16_), .CO(
        add_88_carry_17_), .S(N136) );
  ADDFX2 U366 ( .A(x3[13]), .B(N52), .CI(add_88_carry_17_), .CO(
        add_88_carry_18_), .S(N137) );
  XOR3X2 U367 ( .A(x0_e[21]), .B(x2_e[21]), .C(add_111_carry[22]), .Y(N209) );
  XOR3X2 U368 ( .A(x0_e[21]), .B(add_1_root_add_112_2_B_21_), .C(
        add_1_root_add_112_2_carry[22]), .Y(N277) );
  ADDFX2 U369 ( .A(x1[14]), .B(N30), .CI(add_85_carry_20_), .CO(N74), .S(N73)
         );
  ADDFX2 U370 ( .A(x3[14]), .B(N52), .CI(add_81_carry_19_), .CO(N51), .S(N50)
         );
  ADDFX2 U371 ( .A(x1[14]), .B(N30), .CI(add_80_carry_19_), .CO(N29), .S(N28)
         );
  ADDFX2 U372 ( .A(x1[14]), .B(N30), .CI(add_86_carry_18_), .CO(N95), .S(N94)
         );
  ADDFX2 U373 ( .A(x3[14]), .B(N52), .CI(add_87_carry_20_), .CO(N118), .S(N117) );
  ADDFX2 U374 ( .A(x3[14]), .B(N52), .CI(add_88_carry_18_), .CO(N139), .S(N138) );
  INVX1 U375 ( .A(x2_e[6]), .Y(add_1_root_add_112_2_B_6_) );
  NOR2BX1 U376 ( .AN(y3_tmp[20]), .B(n8), .Y(y3[20]) );
  NOR2BX1 U377 ( .AN(y3_tmp[21]), .B(n8), .Y(y3[21]) );
  NOR2BX1 U378 ( .AN(y2_tmp[20]), .B(n8), .Y(y2[20]) );
  NOR2BX1 U379 ( .AN(y2_tmp[21]), .B(n8), .Y(y2[21]) );
  NOR2BX1 U380 ( .AN(y2_tmp[22]), .B(n8), .Y(y2[22]) );
  NOR2BX1 U381 ( .AN(y1_tmp[20]), .B(n8), .Y(y1[20]) );
  NOR2BX1 U382 ( .AN(y1_tmp[21]), .B(n8), .Y(y1[21]) );
  NOR2BX1 U383 ( .AN(y3_tmp[22]), .B(n8), .Y(y3[22]) );
  NOR2BX1 U384 ( .AN(y0_tmp[20]), .B(n8), .Y(y0[20]) );
  NOR2BX1 U385 ( .AN(y0_tmp[21]), .B(n8), .Y(y0[21]) );
  NOR2BX1 U386 ( .AN(y0_tmp[22]), .B(n3), .Y(y0[22]) );
  NOR2BX1 U387 ( .AN(y1_tmp[22]), .B(n8), .Y(y1[22]) );
  NOR2BX1 U388 ( .AN(y2_tmp[24]), .B(n3), .Y(y2[24]) );
  NOR2BX1 U389 ( .AN(y0_tmp[24]), .B(n8), .Y(y0[24]) );
  NOR2BX1 U390 ( .AN(y1_tmp[24]), .B(n3), .Y(y1[24]) );
  NOR2BX1 U391 ( .AN(y3_tmp[24]), .B(n8), .Y(y3[24]) );
  NOR2BX1 U392 ( .AN(y3_tmp[23]), .B(n8), .Y(y3[23]) );
  NOR2BX1 U393 ( .AN(y2_tmp[23]), .B(n3), .Y(y2[23]) );
  NOR2BX1 U394 ( .AN(y0_tmp[23]), .B(n8), .Y(y0[23]) );
  NOR2BX1 U395 ( .AN(y1_tmp[23]), .B(n3), .Y(y1[23]) );
  BUFX3 U396 ( .A(x1[15]), .Y(N30) );
  BUFX3 U397 ( .A(x3[15]), .Y(N52) );
  INVX1 U398 ( .A(o0[23]), .Y(n85) );
  INVX1 U399 ( .A(o1[23]), .Y(n61) );
  INVX1 U400 ( .A(x2_e[21]), .Y(add_1_root_add_112_2_B_21_) );
  INVX1 U401 ( .A(x3_o1[22]), .Y(n38) );
  XOR2X1 U420 ( .A(y3_tmp[24]), .B(add_125_carry_25_), .Y(N626) );
  AND2X1 U421 ( .A(add_125_carry_24_), .B(y3_tmp[24]), .Y(add_125_carry_25_)
         );
  XOR2X1 U422 ( .A(y3_tmp[24]), .B(add_125_carry_24_), .Y(N625) );
  AND2X1 U423 ( .A(add_125_carry_23_), .B(y3_tmp[23]), .Y(add_125_carry_24_)
         );
  XOR2X1 U424 ( .A(y3_tmp[23]), .B(add_125_carry_23_), .Y(N624) );
  AND2X1 U425 ( .A(add_125_carry_22_), .B(y3_tmp[22]), .Y(add_125_carry_23_)
         );
  XOR2X1 U426 ( .A(y3_tmp[22]), .B(add_125_carry_22_), .Y(N623) );
  AND2X1 U427 ( .A(add_125_carry_21_), .B(y3_tmp[21]), .Y(add_125_carry_22_)
         );
  XOR2X1 U428 ( .A(y3_tmp[21]), .B(add_125_carry_21_), .Y(N622) );
  AND2X1 U429 ( .A(add_125_carry_20_), .B(y3_tmp[20]), .Y(add_125_carry_21_)
         );
  XOR2X1 U430 ( .A(y3_tmp[20]), .B(add_125_carry_20_), .Y(N621) );
  AND2X1 U431 ( .A(add_125_carry_19_), .B(y3_tmp[19]), .Y(add_125_carry_20_)
         );
  XOR2X1 U432 ( .A(y3_tmp[19]), .B(add_125_carry_19_), .Y(N620) );
  AND2X1 U433 ( .A(add_125_carry_18_), .B(y3_tmp[18]), .Y(add_125_carry_19_)
         );
  XOR2X1 U434 ( .A(y3_tmp[18]), .B(add_125_carry_18_), .Y(N619) );
  AND2X1 U435 ( .A(add_125_carry_17_), .B(y3_tmp[17]), .Y(add_125_carry_18_)
         );
  XOR2X1 U436 ( .A(y3_tmp[17]), .B(add_125_carry_17_), .Y(N618) );
  AND2X1 U437 ( .A(add_125_carry_16_), .B(y3_tmp[16]), .Y(add_125_carry_17_)
         );
  XOR2X1 U438 ( .A(y3_tmp[16]), .B(add_125_carry_16_), .Y(N617) );
  AND2X1 U439 ( .A(add_125_carry_15_), .B(y3_tmp[15]), .Y(add_125_carry_16_)
         );
  XOR2X1 U440 ( .A(y3_tmp[15]), .B(add_125_carry_15_), .Y(N616) );
  AND2X1 U441 ( .A(add_125_carry_14_), .B(y3_tmp[14]), .Y(add_125_carry_15_)
         );
  XOR2X1 U442 ( .A(y3_tmp[14]), .B(add_125_carry_14_), .Y(N615) );
  AND2X1 U443 ( .A(add_125_carry_13_), .B(y3_tmp[13]), .Y(add_125_carry_14_)
         );
  XOR2X1 U444 ( .A(y3_tmp[13]), .B(add_125_carry_13_), .Y(N614) );
  AND2X1 U445 ( .A(y3_tmp[11]), .B(y3_tmp[12]), .Y(add_125_carry_13_) );
  XOR2X1 U446 ( .A(y3_tmp[12]), .B(y3_tmp[11]), .Y(N613) );
  XOR2X1 U447 ( .A(y2_tmp[24]), .B(add_124_carry_25_), .Y(N612) );
  AND2X1 U448 ( .A(add_124_carry_24_), .B(y2_tmp[24]), .Y(add_124_carry_25_)
         );
  XOR2X1 U449 ( .A(y2_tmp[24]), .B(add_124_carry_24_), .Y(N611) );
  AND2X1 U450 ( .A(add_124_carry_23_), .B(y2_tmp[23]), .Y(add_124_carry_24_)
         );
  XOR2X1 U451 ( .A(y2_tmp[23]), .B(add_124_carry_23_), .Y(N610) );
  AND2X1 U452 ( .A(add_124_carry_22_), .B(y2_tmp[22]), .Y(add_124_carry_23_)
         );
  XOR2X1 U453 ( .A(y2_tmp[22]), .B(add_124_carry_22_), .Y(N609) );
  AND2X1 U454 ( .A(add_124_carry_21_), .B(y2_tmp[21]), .Y(add_124_carry_22_)
         );
  XOR2X1 U455 ( .A(y2_tmp[21]), .B(add_124_carry_21_), .Y(N608) );
  AND2X1 U456 ( .A(add_124_carry_20_), .B(y2_tmp[20]), .Y(add_124_carry_21_)
         );
  XOR2X1 U457 ( .A(y2_tmp[20]), .B(add_124_carry_20_), .Y(N607) );
  AND2X1 U458 ( .A(add_124_carry_19_), .B(y2_tmp[19]), .Y(add_124_carry_20_)
         );
  XOR2X1 U459 ( .A(y2_tmp[19]), .B(add_124_carry_19_), .Y(N606) );
  AND2X1 U460 ( .A(add_124_carry_18_), .B(y2_tmp[18]), .Y(add_124_carry_19_)
         );
  XOR2X1 U461 ( .A(y2_tmp[18]), .B(add_124_carry_18_), .Y(N605) );
  AND2X1 U462 ( .A(add_124_carry_17_), .B(y2_tmp[17]), .Y(add_124_carry_18_)
         );
  XOR2X1 U463 ( .A(y2_tmp[17]), .B(add_124_carry_17_), .Y(N604) );
  AND2X1 U464 ( .A(add_124_carry_16_), .B(y2_tmp[16]), .Y(add_124_carry_17_)
         );
  XOR2X1 U465 ( .A(y2_tmp[16]), .B(add_124_carry_16_), .Y(N603) );
  AND2X1 U466 ( .A(add_124_carry_15_), .B(y2_tmp[15]), .Y(add_124_carry_16_)
         );
  XOR2X1 U467 ( .A(y2_tmp[15]), .B(add_124_carry_15_), .Y(N602) );
  AND2X1 U468 ( .A(add_124_carry_14_), .B(y2_tmp[14]), .Y(add_124_carry_15_)
         );
  XOR2X1 U469 ( .A(y2_tmp[14]), .B(add_124_carry_14_), .Y(N601) );
  AND2X1 U470 ( .A(add_124_carry_13_), .B(y2_tmp[13]), .Y(add_124_carry_14_)
         );
  XOR2X1 U471 ( .A(y2_tmp[13]), .B(add_124_carry_13_), .Y(N600) );
  AND2X1 U472 ( .A(y2_tmp[11]), .B(y2_tmp[12]), .Y(add_124_carry_13_) );
  XOR2X1 U473 ( .A(y2_tmp[12]), .B(y2_tmp[11]), .Y(N599) );
  XOR2X1 U474 ( .A(y0_tmp[24]), .B(add_122_carry_25_), .Y(N584) );
  AND2X1 U475 ( .A(add_122_carry_24_), .B(y0_tmp[24]), .Y(add_122_carry_25_)
         );
  XOR2X1 U476 ( .A(y0_tmp[24]), .B(add_122_carry_24_), .Y(N583) );
  AND2X1 U477 ( .A(add_122_carry_23_), .B(y0_tmp[23]), .Y(add_122_carry_24_)
         );
  XOR2X1 U478 ( .A(y0_tmp[23]), .B(add_122_carry_23_), .Y(N582) );
  AND2X1 U479 ( .A(add_122_carry_22_), .B(y0_tmp[22]), .Y(add_122_carry_23_)
         );
  XOR2X1 U480 ( .A(y0_tmp[22]), .B(add_122_carry_22_), .Y(N581) );
  AND2X1 U481 ( .A(add_122_carry_21_), .B(y0_tmp[21]), .Y(add_122_carry_22_)
         );
  XOR2X1 U482 ( .A(y0_tmp[21]), .B(add_122_carry_21_), .Y(N580) );
  AND2X1 U483 ( .A(add_122_carry_20_), .B(y0_tmp[20]), .Y(add_122_carry_21_)
         );
  XOR2X1 U484 ( .A(y0_tmp[20]), .B(add_122_carry_20_), .Y(N579) );
  AND2X1 U485 ( .A(add_122_carry_19_), .B(y0_tmp[19]), .Y(add_122_carry_20_)
         );
  XOR2X1 U486 ( .A(y0_tmp[19]), .B(add_122_carry_19_), .Y(N578) );
  AND2X1 U487 ( .A(add_122_carry_18_), .B(y0_tmp[18]), .Y(add_122_carry_19_)
         );
  XOR2X1 U488 ( .A(y0_tmp[18]), .B(add_122_carry_18_), .Y(N577) );
  AND2X1 U489 ( .A(add_122_carry_17_), .B(y0_tmp[17]), .Y(add_122_carry_18_)
         );
  XOR2X1 U490 ( .A(y0_tmp[17]), .B(add_122_carry_17_), .Y(N576) );
  AND2X1 U491 ( .A(add_122_carry_16_), .B(y0_tmp[16]), .Y(add_122_carry_17_)
         );
  XOR2X1 U492 ( .A(y0_tmp[16]), .B(add_122_carry_16_), .Y(N575) );
  AND2X1 U493 ( .A(add_122_carry_15_), .B(y0_tmp[15]), .Y(add_122_carry_16_)
         );
  XOR2X1 U494 ( .A(y0_tmp[15]), .B(add_122_carry_15_), .Y(N574) );
  AND2X1 U495 ( .A(add_122_carry_14_), .B(y0_tmp[14]), .Y(add_122_carry_15_)
         );
  XOR2X1 U496 ( .A(y0_tmp[14]), .B(add_122_carry_14_), .Y(N573) );
  AND2X1 U497 ( .A(add_122_carry_13_), .B(y0_tmp[13]), .Y(add_122_carry_14_)
         );
  XOR2X1 U498 ( .A(y0_tmp[13]), .B(add_122_carry_13_), .Y(N572) );
  AND2X1 U499 ( .A(y0_tmp[11]), .B(y0_tmp[12]), .Y(add_122_carry_13_) );
  XOR2X1 U500 ( .A(y0_tmp[12]), .B(y0_tmp[11]), .Y(N571) );
  XOR2X1 U501 ( .A(y1_tmp[24]), .B(add_123_carry_25_), .Y(N598) );
  AND2X1 U502 ( .A(add_123_carry_24_), .B(y1_tmp[24]), .Y(add_123_carry_25_)
         );
  XOR2X1 U503 ( .A(y1_tmp[24]), .B(add_123_carry_24_), .Y(N597) );
  AND2X1 U504 ( .A(add_123_carry_23_), .B(y1_tmp[23]), .Y(add_123_carry_24_)
         );
  XOR2X1 U505 ( .A(y1_tmp[23]), .B(add_123_carry_23_), .Y(N596) );
  AND2X1 U506 ( .A(add_123_carry_22_), .B(y1_tmp[22]), .Y(add_123_carry_23_)
         );
  XOR2X1 U507 ( .A(y1_tmp[22]), .B(add_123_carry_22_), .Y(N595) );
  AND2X1 U508 ( .A(add_123_carry_21_), .B(y1_tmp[21]), .Y(add_123_carry_22_)
         );
  XOR2X1 U509 ( .A(y1_tmp[21]), .B(add_123_carry_21_), .Y(N594) );
  AND2X1 U510 ( .A(add_123_carry_20_), .B(y1_tmp[20]), .Y(add_123_carry_21_)
         );
  XOR2X1 U511 ( .A(y1_tmp[20]), .B(add_123_carry_20_), .Y(N593) );
  AND2X1 U512 ( .A(add_123_carry_19_), .B(y1_tmp[19]), .Y(add_123_carry_20_)
         );
  XOR2X1 U513 ( .A(y1_tmp[19]), .B(add_123_carry_19_), .Y(N592) );
  AND2X1 U514 ( .A(add_123_carry_18_), .B(y1_tmp[18]), .Y(add_123_carry_19_)
         );
  XOR2X1 U515 ( .A(y1_tmp[18]), .B(add_123_carry_18_), .Y(N591) );
  AND2X1 U516 ( .A(add_123_carry_17_), .B(y1_tmp[17]), .Y(add_123_carry_18_)
         );
  XOR2X1 U517 ( .A(y1_tmp[17]), .B(add_123_carry_17_), .Y(N590) );
  AND2X1 U518 ( .A(add_123_carry_16_), .B(y1_tmp[16]), .Y(add_123_carry_17_)
         );
  XOR2X1 U519 ( .A(y1_tmp[16]), .B(add_123_carry_16_), .Y(N589) );
  AND2X1 U520 ( .A(add_123_carry_15_), .B(y1_tmp[15]), .Y(add_123_carry_16_)
         );
  XOR2X1 U521 ( .A(y1_tmp[15]), .B(add_123_carry_15_), .Y(N588) );
  AND2X1 U522 ( .A(add_123_carry_14_), .B(y1_tmp[14]), .Y(add_123_carry_15_)
         );
  XOR2X1 U523 ( .A(y1_tmp[14]), .B(add_123_carry_14_), .Y(N587) );
  AND2X1 U524 ( .A(add_123_carry_13_), .B(y1_tmp[13]), .Y(add_123_carry_14_)
         );
  XOR2X1 U525 ( .A(y1_tmp[13]), .B(add_123_carry_13_), .Y(N586) );
  AND2X1 U526 ( .A(y1_tmp[11]), .B(y1_tmp[12]), .Y(add_123_carry_13_) );
  XOR2X1 U527 ( .A(y1_tmp[12]), .B(y1_tmp[11]), .Y(N585) );
  AND2X1 U528 ( .A(x0_e[6]), .B(x2_e[6]), .Y(add_111_carry[7]) );
  XOR2X1 U529 ( .A(x2_e[6]), .B(x0_e[6]), .Y(N193) );
  OR2X1 U530 ( .A(add_1_root_add_112_2_B_6_), .B(x0_e[6]), .Y(
        add_1_root_add_112_2_carry[7]) );
  XNOR2X1 U531 ( .A(x0_e[6]), .B(add_1_root_add_112_2_B_6_), .Y(N261) );
  AND2X1 U532 ( .A(x1[0]), .B(x1[6]), .Y(add_85_carry_7_) );
  XOR2X1 U533 ( .A(x1[6]), .B(x1[0]), .Y(N59) );
  AND2X1 U534 ( .A(x3[0]), .B(x3[3]), .Y(add_81_carry_6_) );
  XOR2X1 U535 ( .A(x3[3]), .B(x3[0]), .Y(N36) );
  AND2X1 U536 ( .A(x1[0]), .B(x1[3]), .Y(add_80_carry_6_) );
  XOR2X1 U537 ( .A(x1[3]), .B(x1[0]), .Y(N14) );
  AND2X1 U538 ( .A(x1[0]), .B(x1[3]), .Y(add_86_carry_5_) );
  XOR2X1 U539 ( .A(x1[3]), .B(x1[0]), .Y(N80) );
  AND2X1 U540 ( .A(x3[0]), .B(x3[6]), .Y(add_87_carry_7_) );
  XOR2X1 U541 ( .A(x3[6]), .B(x3[0]), .Y(N103) );
  AND2X1 U542 ( .A(x3[0]), .B(x3[3]), .Y(add_88_carry_5_) );
  XOR2X1 U543 ( .A(x3[3]), .B(x3[0]), .Y(N124) );
endmodule


module idct8_shift12_add2048_DW01_add_8 ( A, B, SUM );
  input [25:0] A;
  input [25:0] B;
  output [25:0] SUM;
  wire   n1, n2;
  wire   [25:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  XOR3X2 U1_25 ( .A(A[25]), .B(B[25]), .C(carry[25]), .Y(SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  INVX1 U1 ( .A(A[0]), .Y(n2) );
  XNOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  NAND2X1 U3 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U4 ( .A(B[0]), .Y(n1) );
endmodule


module idct8_shift12_add2048_DW01_add_9 ( A, B, SUM );
  input [25:0] A;
  input [25:0] B;
  output [25:0] SUM;
  wire   n1, n2;
  wire   [25:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  XOR3X2 U1_25 ( .A(A[25]), .B(B[25]), .C(carry[25]), .Y(SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  INVX1 U1 ( .A(A[0]), .Y(n2) );
  XNOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  NAND2X1 U3 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U4 ( .A(B[0]), .Y(n1) );
endmodule


module idct8_shift12_add2048_DW01_add_10 ( A, B, SUM );
  input [25:0] A;
  input [25:0] B;
  output [25:0] SUM;
  wire   n1, n2;
  wire   [25:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  XOR3X2 U1_25 ( .A(A[25]), .B(B[25]), .C(carry[25]), .Y(SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  INVX1 U1 ( .A(A[0]), .Y(n2) );
  XNOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  NAND2X1 U3 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U4 ( .A(B[0]), .Y(n1) );
endmodule


module idct8_shift12_add2048_DW01_add_11 ( A, B, SUM );
  input [25:0] A;
  input [25:0] B;
  output [25:0] SUM;
  wire   n1, n2;
  wire   [25:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  XOR3X2 U1_25 ( .A(A[25]), .B(B[25]), .C(carry[25]), .Y(SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  INVX1 U1 ( .A(A[0]), .Y(n2) );
  XNOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  NAND2X1 U3 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U4 ( .A(B[0]), .Y(n1) );
endmodule


module idct8_shift12_add2048_DW01_add_12 ( A, B, SUM );
  input [25:0] A;
  input [25:0] B;
  output [25:0] SUM;
  wire   n1;
  wire   [25:2] carry;

  XOR3X2 U1_25 ( .A(A[25]), .B(B[25]), .C(carry[25]), .Y(SUM[25]) );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module idct8_shift12_add2048_DW01_add_13 ( A, B, SUM );
  input [25:0] A;
  input [25:0] B;
  output [25:0] SUM;
  wire   n1;
  wire   [25:2] carry;

  XOR3X2 U1_25 ( .A(A[25]), .B(B[25]), .C(carry[25]), .Y(SUM[25]) );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module idct8_shift12_add2048_DW01_add_14 ( A, B, SUM );
  input [25:0] A;
  input [25:0] B;
  output [25:0] SUM;
  wire   n1;
  wire   [25:2] carry;

  XOR3X2 U1_25 ( .A(A[25]), .B(B[25]), .C(carry[25]), .Y(SUM[25]) );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module idct8_shift12_add2048_DW01_add_15 ( A, B, SUM );
  input [25:0] A;
  input [25:0] B;
  output [25:0] SUM;
  wire   n1;
  wire   [25:2] carry;

  XOR3X2 U1_25 ( .A(A[25]), .B(B[25]), .C(carry[25]), .Y(SUM[25]) );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module idct8_shift12_add2048_DW01_add_16 ( A, B, SUM );
  input [24:0] A;
  input [24:0] B;
  output [24:0] SUM;
  wire   n1;
  wire   [24:2] carry;

  XOR3X2 U1_24 ( .A(A[24]), .B(B[24]), .C(carry[24]), .Y(SUM[24]) );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module idct8_shift12_add2048_DW01_add_17 ( A, B, SUM );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  wire   n1;
  wire   [23:2] carry;

  XOR3X2 U1_23 ( .A(A[23]), .B(B[23]), .C(carry[23]), .Y(SUM[23]) );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module idct8_shift12_add2048_DW01_add_18 ( A, B, SUM );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;

  wire   [23:1] carry;

  XOR3X2 U1_23 ( .A(A[23]), .B(B[23]), .C(carry[23]), .Y(SUM[23]) );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(1'b0), .CO(carry[2]), .S(SUM[1]) );
  XOR2X1 U1 ( .A(1'b0), .B(A[0]), .Y(SUM[0]) );
endmodule


module idct8_shift12_add2048_DW01_add_19 ( A, B, SUM );
  input [24:0] A;
  input [24:0] B;
  output [24:0] SUM;
  wire   n1;
  wire   [24:2] carry;

  XOR3X2 U1_24 ( .A(A[24]), .B(B[24]), .C(carry[24]), .Y(SUM[24]) );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module idct8_shift12_add2048_DW01_add_20 ( A, B, SUM );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  wire   n1, n2;
  wire   [23:1] carry;

  XOR3X2 U1_23 ( .A(A[23]), .B(B[23]), .C(carry[23]), .Y(SUM[23]) );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  INVX1 U1 ( .A(B[0]), .Y(n1) );
  NAND2X1 U2 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U3 ( .A(A[0]), .Y(n2) );
  XNOR2X1 U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module idct8_shift12_add2048_DW01_add_21 ( A, B, SUM );
  input [24:0] A;
  input [24:0] B;
  output [24:0] SUM;
  wire   n1;
  wire   [24:2] carry;

  XOR3X2 U1_24 ( .A(A[24]), .B(B[24]), .C(carry[24]), .Y(SUM[24]) );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module idct8_shift12_add2048_DW01_add_22 ( A, B, SUM );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  wire   n1;
  wire   [23:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  XOR3X2 U1_23 ( .A(A[23]), .B(B[23]), .C(carry[23]), .Y(SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  CLKINVX8 U1 ( .A(n1), .Y(carry[1]) );
  CLKINVX8 U2 ( .A(B[0]), .Y(SUM[0]) );
  INVX1 U3 ( .A(B[0]), .Y(n1) );
endmodule


module idct8_shift12_add2048_DW01_add_23 ( A, B, SUM );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  wire   n1;
  wire   [23:2] carry;

  XOR3X2 U1_23 ( .A(A[23]), .B(B[23]), .C(carry[23]), .Y(SUM[23]) );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module idct8_shift12_add2048_DW01_add_24 ( A, B, SUM );
  input [24:0] A;
  input [24:0] B;
  output [24:0] SUM;
  wire   n1;
  wire   [24:2] carry;

  XOR3X2 U1_24 ( .A(A[24]), .B(B[24]), .C(carry[24]), .Y(SUM[24]) );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module idct8_shift12_add2048_DW01_add_25 ( A, B, SUM );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  wire   n1, n2;
  wire   [23:1] carry;

  XOR3X2 U1_23 ( .A(A[23]), .B(B[23]), .C(carry[23]), .Y(SUM[23]) );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  INVX1 U1 ( .A(B[0]), .Y(n1) );
  NAND2X1 U2 ( .A(n1), .B(n2), .Y(carry[1]) );
  INVX1 U3 ( .A(A[0]), .Y(n2) );
  XNOR2X1 U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module idct8_shift12_add2048_DW01_add_26 ( A, B, SUM );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  wire   n1;
  wire   [23:1] carry;

  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  XOR3X2 U1_23 ( .A(A[23]), .B(B[23]), .C(carry[23]), .Y(SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  CLKINVX8 U1 ( .A(n1), .Y(carry[1]) );
  CLKINVX8 U2 ( .A(B[0]), .Y(SUM[0]) );
  INVX1 U3 ( .A(B[0]), .Y(n1) );
endmodule


module idct8_shift12_add2048_DW01_add_27 ( A, B, SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n1;
  wire   [20:6] carry;

  XOR3X2 U1_20 ( .A(A[20]), .B(B[20]), .C(carry[20]), .Y(SUM[20]) );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(n1), .CO(carry[6]), .S(SUM[5]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  AND2X2 U1 ( .A(B[4]), .B(A[4]), .Y(n1) );
  XOR2X1 U2 ( .A(B[4]), .B(A[4]), .Y(SUM[4]) );
  BUFX3 U3 ( .A(B[3]), .Y(SUM[3]) );
  BUFX3 U4 ( .A(B[2]), .Y(SUM[2]) );
  BUFX3 U5 ( .A(B[1]), .Y(SUM[1]) );
endmodule


module idct8_shift12_add2048_DW01_add_28 ( A, B, SUM );
  input [21:0] A;
  input [21:0] B;
  output [21:0] SUM;
  wire   n1;
  wire   [21:7] carry;

  XOR3X2 U1_21 ( .A(A[21]), .B(B[21]), .C(carry[21]), .Y(SUM[21]) );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(n1), .CO(carry[7]), .S(SUM[6]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  AND2X2 U1 ( .A(B[5]), .B(A[5]), .Y(n1) );
  XOR2X1 U2 ( .A(B[5]), .B(A[5]), .Y(SUM[5]) );
  BUFX3 U3 ( .A(B[4]), .Y(SUM[4]) );
  BUFX3 U4 ( .A(B[3]), .Y(SUM[3]) );
  BUFX3 U5 ( .A(B[2]), .Y(SUM[2]) );
  BUFX3 U6 ( .A(B[1]), .Y(SUM[1]) );
endmodule


module idct8_shift12_add2048_DW01_add_29 ( A, B, SUM );
  input [22:0] A;
  input [22:0] B;
  output [22:0] SUM;

  wire   [22:1] carry;

  XOR3X2 U1_22 ( .A(A[22]), .B(B[22]), .C(carry[22]), .Y(SUM[22]) );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(1'b0), .CO(carry[2]), .S(SUM[1]) );
  XOR2X1 U1 ( .A(1'b0), .B(A[0]), .Y(SUM[0]) );
endmodule


module idct8_shift12_add2048_DW01_add_30 ( A, B, SUM );
  input [22:0] A;
  input [22:0] B;
  output [22:0] SUM;

  wire   [22:1] carry;

  XOR3X2 U1_22 ( .A(A[22]), .B(B[22]), .C(carry[22]), .Y(SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_1 ( .A(A[1]), .B(1'b0), .CI(1'b0), .S(SUM[1]) );
  ADDFX2 U1_2 ( .A(A[2]), .B(1'b0), .CI(1'b0), .S(SUM[2]) );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(1'b0), .CO(carry[4]), .S(SUM[3]) );
  XOR2X1 U1 ( .A(1'b0), .B(A[0]), .Y(SUM[0]) );
endmodule


module idct8_shift12_add2048_DW01_add_31 ( A, B, SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n1;
  wire   [20:6] carry;

  XOR3X2 U1_20 ( .A(A[20]), .B(B[20]), .C(carry[20]), .Y(SUM[20]) );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(n1), .CO(carry[6]), .S(SUM[5]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  AND2X2 U1 ( .A(B[4]), .B(A[4]), .Y(n1) );
  XOR2X1 U2 ( .A(B[4]), .B(A[4]), .Y(SUM[4]) );
  BUFX3 U3 ( .A(B[3]), .Y(SUM[3]) );
  BUFX3 U4 ( .A(B[2]), .Y(SUM[2]) );
  BUFX3 U5 ( .A(B[1]), .Y(SUM[1]) );
endmodule


module idct8_shift12_add2048_DW01_add_32 ( A, B, SUM );
  input [21:0] A;
  input [21:0] B;
  output [21:0] SUM;
  wire   n1;
  wire   [21:7] carry;

  XOR3X2 U1_21 ( .A(A[21]), .B(B[21]), .C(carry[21]), .Y(SUM[21]) );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(n1), .CO(carry[7]), .S(SUM[6]) );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  AND2X2 U1 ( .A(B[5]), .B(A[5]), .Y(n1) );
  XOR2X1 U2 ( .A(B[5]), .B(A[5]), .Y(SUM[5]) );
  BUFX3 U3 ( .A(B[4]), .Y(SUM[4]) );
  BUFX3 U4 ( .A(B[3]), .Y(SUM[3]) );
  BUFX3 U5 ( .A(B[2]), .Y(SUM[2]) );
  BUFX3 U6 ( .A(B[1]), .Y(SUM[1]) );
endmodule


module idct8_shift12_add2048_DW01_add_33 ( A, B, SUM );
  input [22:0] A;
  input [22:0] B;
  output [22:0] SUM;

  wire   [22:1] carry;

  XOR3X2 U1_22 ( .A(A[22]), .B(B[22]), .C(carry[22]), .Y(SUM[22]) );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(1'b0), .CO(carry[2]), .S(SUM[1]) );
  XOR2X1 U1 ( .A(1'b0), .B(A[0]), .Y(SUM[0]) );
endmodule


module idct8_shift12_add2048_DW01_add_34 ( A, B, SUM );
  input [22:0] A;
  input [22:0] B;
  output [22:0] SUM;

  wire   [22:1] carry;

  XOR3X2 U1_22 ( .A(A[22]), .B(B[22]), .C(carry[22]), .Y(SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_1 ( .A(A[1]), .B(1'b0), .CI(1'b0), .S(SUM[1]) );
  ADDFX2 U1_2 ( .A(A[2]), .B(1'b0), .CI(1'b0), .S(SUM[2]) );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(1'b0), .CO(carry[4]), .S(SUM[3]) );
  XOR2X1 U1 ( .A(1'b0), .B(A[0]), .Y(SUM[0]) );
endmodule


module idct8_shift12_add2048_DW01_add_35 ( A, B, SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n1;
  wire   [20:6] carry;

  XOR3X2 U1_20 ( .A(A[20]), .B(B[20]), .C(carry[20]), .Y(SUM[20]) );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(n1), .CO(carry[6]), .S(SUM[5]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  AND2X2 U1 ( .A(B[4]), .B(A[4]), .Y(n1) );
  XOR2X1 U2 ( .A(B[4]), .B(A[4]), .Y(SUM[4]) );
  BUFX3 U3 ( .A(B[3]), .Y(SUM[3]) );
  BUFX3 U4 ( .A(B[2]), .Y(SUM[2]) );
  BUFX3 U5 ( .A(B[1]), .Y(SUM[1]) );
endmodule


module idct8_shift12_add2048_DW01_add_36 ( A, B, SUM );
  input [21:0] A;
  input [21:0] B;
  output [21:0] SUM;
  wire   n1;
  wire   [21:7] carry;

  XOR3X2 U1_21 ( .A(A[21]), .B(B[21]), .C(carry[21]), .Y(SUM[21]) );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(n1), .CO(carry[7]), .S(SUM[6]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  AND2X2 U1 ( .A(B[5]), .B(A[5]), .Y(n1) );
  XOR2X1 U2 ( .A(B[5]), .B(A[5]), .Y(SUM[5]) );
  BUFX3 U3 ( .A(B[4]), .Y(SUM[4]) );
  BUFX3 U4 ( .A(B[3]), .Y(SUM[3]) );
  BUFX3 U5 ( .A(B[2]), .Y(SUM[2]) );
  BUFX3 U6 ( .A(B[1]), .Y(SUM[1]) );
endmodule


module idct8_shift12_add2048_DW01_add_37 ( A, B, SUM );
  input [22:0] A;
  input [22:0] B;
  output [22:0] SUM;

  wire   [22:1] carry;

  XOR3X2 U1_22 ( .A(A[22]), .B(B[22]), .C(carry[22]), .Y(SUM[22]) );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(1'b0), .CO(carry[2]), .S(SUM[1]) );
  XOR2X1 U1 ( .A(1'b0), .B(A[0]), .Y(SUM[0]) );
endmodule


module idct8_shift12_add2048_DW01_add_38 ( A, B, SUM );
  input [22:0] A;
  input [22:0] B;
  output [22:0] SUM;

  wire   [22:1] carry;

  XOR3X2 U1_22 ( .A(A[22]), .B(B[22]), .C(carry[22]), .Y(SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_1 ( .A(A[1]), .B(1'b0), .CI(1'b0), .S(SUM[1]) );
  ADDFX2 U1_2 ( .A(A[2]), .B(1'b0), .CI(1'b0), .S(SUM[2]) );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(1'b0), .CO(carry[4]), .S(SUM[3]) );
  XOR2X1 U1 ( .A(1'b0), .B(A[0]), .Y(SUM[0]) );
endmodule


module idct8_shift12_add2048_DW01_add_39 ( A, B, SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n1;
  wire   [20:6] carry;

  XOR3X2 U1_20 ( .A(A[20]), .B(B[20]), .C(carry[20]), .Y(SUM[20]) );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(n1), .CO(carry[6]), .S(SUM[5]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  AND2X2 U1 ( .A(B[4]), .B(A[4]), .Y(n1) );
  XOR2X1 U2 ( .A(B[4]), .B(A[4]), .Y(SUM[4]) );
  BUFX3 U3 ( .A(B[1]), .Y(SUM[1]) );
  BUFX3 U4 ( .A(B[2]), .Y(SUM[2]) );
  BUFX3 U5 ( .A(B[3]), .Y(SUM[3]) );
endmodule


module idct8_shift12_add2048_DW01_add_40 ( A, B, SUM );
  input [21:0] A;
  input [21:0] B;
  output [21:0] SUM;
  wire   n1;
  wire   [21:7] carry;

  XOR3X2 U1_21 ( .A(A[21]), .B(B[21]), .C(carry[21]), .Y(SUM[21]) );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(n1), .CO(carry[7]), .S(SUM[6]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  AND2X2 U1 ( .A(B[5]), .B(A[5]), .Y(n1) );
  XOR2X1 U2 ( .A(B[5]), .B(A[5]), .Y(SUM[5]) );
  BUFX3 U3 ( .A(B[1]), .Y(SUM[1]) );
  BUFX3 U4 ( .A(B[2]), .Y(SUM[2]) );
  BUFX3 U5 ( .A(B[3]), .Y(SUM[3]) );
  BUFX3 U6 ( .A(B[4]), .Y(SUM[4]) );
endmodule


module idct8_shift12_add2048_DW01_add_41 ( A, B, SUM );
  input [22:0] A;
  input [22:0] B;
  output [22:0] SUM;

  wire   [22:1] carry;

  XOR3X2 U1_22 ( .A(A[22]), .B(B[22]), .C(carry[22]), .Y(SUM[22]) );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(1'b0), .CO(carry[2]), .S(SUM[1]) );
  XOR2X1 U1 ( .A(1'b0), .B(A[0]), .Y(SUM[0]) );
endmodule


module idct8_shift12_add2048_DW01_add_42 ( A, B, SUM );
  input [22:0] A;
  input [22:0] B;
  output [22:0] SUM;

  wire   [22:1] carry;

  XOR3X2 U1_22 ( .A(A[22]), .B(B[22]), .C(carry[22]), .Y(SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_1 ( .A(A[1]), .B(1'b0), .CI(1'b0), .S(SUM[1]) );
  ADDFX2 U1_2 ( .A(A[2]), .B(1'b0), .CI(1'b0), .S(SUM[2]) );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(1'b0), .CO(carry[4]), .S(SUM[3]) );
  XOR2X1 U1 ( .A(1'b0), .B(A[0]), .Y(SUM[0]) );
endmodule


module idct8_shift12_add2048_DW01_add_59 ( A, B, SUM );
  input [24:0] A;
  input [24:0] B;
  output [24:0] SUM;

  wire   [23:1] carry;

  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  XOR3X2 U1_23 ( .A(A[23]), .B(B[23]), .C(carry[23]), .Y(SUM[23]) );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(1'b0), .CO(carry[2]), .S(SUM[1]) );
  XOR2X1 U1 ( .A(B[0]), .B(1'b0), .Y(SUM[0]) );
endmodule


module idct8_shift12_add2048_DW01_sub_0 ( B, DIFF );
  input [23:0] B;
  output [23:0] DIFF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46;

  AND2X2 U1 ( .A(n35), .B(n21), .Y(n1) );
  AND2X2 U2 ( .A(n34), .B(n1), .Y(n2) );
  AND2X2 U3 ( .A(n33), .B(n2), .Y(n3) );
  AND2X2 U4 ( .A(n32), .B(n3), .Y(n4) );
  AND2X2 U5 ( .A(n31), .B(n4), .Y(n5) );
  AND2X2 U6 ( .A(n30), .B(n5), .Y(n6) );
  AND2X2 U7 ( .A(n29), .B(n6), .Y(n7) );
  AND2X2 U8 ( .A(n28), .B(n7), .Y(n8) );
  AND2X2 U9 ( .A(n27), .B(n8), .Y(n9) );
  AND2X2 U10 ( .A(n26), .B(n9), .Y(n10) );
  AND2X2 U11 ( .A(n25), .B(n10), .Y(n11) );
  XOR2X1 U12 ( .A(n25), .B(n10), .Y(DIFF[21]) );
  XOR2X1 U13 ( .A(n24), .B(n11), .Y(DIFF[22]) );
  AND2X2 U14 ( .A(n45), .B(n46), .Y(n12) );
  AND2X2 U15 ( .A(n44), .B(n12), .Y(n13) );
  AND2X2 U16 ( .A(n43), .B(n13), .Y(n14) );
  AND2X2 U17 ( .A(n42), .B(n14), .Y(n15) );
  AND2X2 U18 ( .A(n41), .B(n15), .Y(n16) );
  AND2X2 U19 ( .A(n40), .B(n16), .Y(n17) );
  AND2X2 U20 ( .A(n39), .B(n17), .Y(n18) );
  AND2X2 U21 ( .A(n38), .B(n18), .Y(n19) );
  AND2X2 U22 ( .A(n37), .B(n19), .Y(n20) );
  AND2X2 U23 ( .A(n36), .B(n20), .Y(n21) );
  XOR2X1 U24 ( .A(n29), .B(n6), .Y(DIFF[17]) );
  XOR2X1 U25 ( .A(n28), .B(n7), .Y(DIFF[18]) );
  XOR2X1 U26 ( .A(n27), .B(n8), .Y(DIFF[19]) );
  XOR2X1 U27 ( .A(n26), .B(n9), .Y(DIFF[20]) );
  XOR2X1 U28 ( .A(n34), .B(n1), .Y(DIFF[12]) );
  XOR2X1 U29 ( .A(n33), .B(n2), .Y(DIFF[13]) );
  XOR2X1 U30 ( .A(n32), .B(n3), .Y(DIFF[14]) );
  XOR2X1 U31 ( .A(n31), .B(n4), .Y(DIFF[15]) );
  XOR2X1 U32 ( .A(n30), .B(n5), .Y(DIFF[16]) );
  XOR2X1 U33 ( .A(n38), .B(n18), .Y(DIFF[8]) );
  XOR2X1 U34 ( .A(n37), .B(n19), .Y(DIFF[9]) );
  XOR2X1 U35 ( .A(n36), .B(n20), .Y(DIFF[10]) );
  XOR2X1 U36 ( .A(n35), .B(n21), .Y(DIFF[11]) );
  XOR2X1 U37 ( .A(n43), .B(n13), .Y(DIFF[3]) );
  XOR2X1 U38 ( .A(n42), .B(n14), .Y(DIFF[4]) );
  XOR2X1 U39 ( .A(n41), .B(n15), .Y(DIFF[5]) );
  XOR2X1 U40 ( .A(n40), .B(n16), .Y(DIFF[6]) );
  XOR2X1 U41 ( .A(n39), .B(n17), .Y(DIFF[7]) );
  XOR2X1 U42 ( .A(n44), .B(n12), .Y(DIFF[2]) );
  XOR2X1 U43 ( .A(n45), .B(n46), .Y(DIFF[1]) );
  INVX1 U44 ( .A(B[11]), .Y(n35) );
  INVX1 U45 ( .A(B[12]), .Y(n34) );
  INVX1 U46 ( .A(B[13]), .Y(n33) );
  INVX1 U47 ( .A(B[14]), .Y(n32) );
  INVX1 U48 ( .A(B[15]), .Y(n31) );
  INVX1 U49 ( .A(B[16]), .Y(n30) );
  INVX1 U50 ( .A(B[17]), .Y(n29) );
  INVX1 U51 ( .A(B[18]), .Y(n28) );
  INVX1 U52 ( .A(B[19]), .Y(n27) );
  INVX1 U53 ( .A(B[20]), .Y(n26) );
  INVX1 U54 ( .A(B[21]), .Y(n25) );
  INVX1 U55 ( .A(B[22]), .Y(n24) );
  XOR2X1 U56 ( .A(B[23]), .B(n23), .Y(DIFF[23]) );
  NAND2X1 U57 ( .A(n24), .B(n11), .Y(n23) );
  INVX1 U58 ( .A(B[0]), .Y(n46) );
  INVX1 U59 ( .A(B[1]), .Y(n45) );
  INVX1 U60 ( .A(B[2]), .Y(n44) );
  INVX1 U61 ( .A(B[3]), .Y(n43) );
  INVX1 U62 ( .A(B[4]), .Y(n42) );
  INVX1 U63 ( .A(B[5]), .Y(n41) );
  INVX1 U64 ( .A(B[6]), .Y(n40) );
  INVX1 U65 ( .A(B[7]), .Y(n39) );
  INVX1 U66 ( .A(B[8]), .Y(n38) );
  INVX1 U67 ( .A(B[9]), .Y(n37) );
  INVX1 U68 ( .A(B[10]), .Y(n36) );
  BUFX3 U69 ( .A(B[0]), .Y(DIFF[0]) );
endmodule


module idct8_shift12_add2048 ( clk, rstn, mode, start, x0, x1, x2, x3, x4, x5, 
        x6, x7, y0, y1, y2, y3, y4, y5, y6, y7, idct8_ready );
  input [1:0] mode;
  input [24:0] x0;
  input [24:0] x1;
  input [24:0] x2;
  input [24:0] x3;
  input [15:0] x4;
  input [15:0] x5;
  input [15:0] x6;
  input [15:0] x7;
  output [25:0] y0;
  output [25:0] y1;
  output [25:0] y2;
  output [25:0] y3;
  output [25:0] y4;
  output [25:0] y5;
  output [25:0] y6;
  output [25:0] y7;
  input clk, rstn, start;
  output idct8_ready;
  wire   N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36,
         N37, N38, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55,
         N56, N57, N58, N59, N60, N64, N65, N66, N67, N68, N69, N70, N71, N72,
         N73, N74, N75, N76, N77, N78, N79, N80, N85, N86, N87, N88, N89, N90,
         N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N108, N109,
         N110, N111, N112, N113, N114, N115, N116, N117, N118, N119, N120,
         N121, N122, N123, N129, N130, N131, N132, N133, N134, N135, N136,
         N137, N138, N139, N140, N141, N142, N143, N144, N145, N149, N150,
         N151, N152, N153, N154, N155, N156, N157, N158, N159, N160, N161,
         N162, N163, N164, N165, N170, N171, N172, N173, N174, N175, N176,
         N177, N178, N179, N180, N181, N182, N183, N184, N185, N186, N193,
         N194, N195, N196, N197, N198, N199, N200, N201, N202, N203, N204,
         N205, N206, N207, N208, N214, N215, N216, N217, N218, N219, N220,
         N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N234,
         N235, N236, N237, N238, N239, N240, N241, N242, N243, N244, N245,
         N246, N247, N248, N249, N250, N255, N256, N257, N258, N259, N260,
         N261, N262, N263, N264, N265, N266, N267, N268, N269, N270, N271,
         N278, N279, N280, N281, N282, N283, N284, N285, N286, N287, N288,
         N289, N290, N291, N292, N293, N299, N300, N301, N302, N303, N304,
         N305, N306, N307, N308, N309, N310, N311, N312, N313, N314, N315,
         N319, N320, N321, N322, N323, N324, N325, N326, N327, N328, N329,
         N330, N331, N332, N333, N334, N335, N340, N341, N342, N343, N344,
         N345, N346, N347, N348, N349, N350, N351, N352, N353, N354, N355,
         N356, N357, N358, N359, N360, N361, N362, N363, N364, N365, N366,
         N367, N368, N369, N370, N371, N372, N373, N374, N375, N376, N377,
         N378, N379, N380, N381, N382, N383, N384, N385, N386, N387, N388,
         N389, N390, N391, N392, N393, N394, N395, N396, N397, N398, N399,
         N400, N401, N402, N404, N405, N406, N407, N408, N409, N410, N411,
         N412, N413, N414, N415, N416, N417, N418, N419, N420, N421, N422,
         N423, N424, N426, N427, N428, N429, N430, N431, N432, N433, N434,
         N435, N436, N437, N438, N439, N440, N441, N442, N443, N444, N445,
         N446, N447, N448, N449, N450, N451, N452, N453, N454, N455, N456,
         N457, N458, N459, N460, N461, N462, N463, N464, N465, N466, N467,
         N468, N469, N470, N471, N472, N473, N474, N475, N476, N477, N478,
         N479, N480, N481, N482, N483, N484, N485, N486, N487, N488, N489,
         N490, N491, N493, N494, N495, N496, N497, N498, N499, N500, N501,
         N502, N503, N504, N505, N506, N507, N508, N509, N510, N511, N512,
         N513, N515, N516, N517, N518, N519, N520, N521, N522, N523, N524,
         N525, N526, N527, N528, N529, N530, N531, N532, N533, N534, N535,
         N536, N537, N538, N539, N540, N541, N542, N543, N544, N545, N546,
         N547, N548, N549, N550, N551, N552, N553, N554, N555, N556, N557,
         N558, N559, N560, N561, N562, N563, N564, N565, N566, N567, N568,
         N569, N570, N571, N572, N573, N574, N575, N576, N577, N578, N579,
         N580, N582, N583, N584, N585, N586, N587, N588, N589, N590, N591,
         N592, N593, N594, N595, N596, N597, N598, N599, N600, N601, N602,
         N604, N605, N606, N607, N608, N609, N610, N611, N612, N613, N614,
         N615, N616, N617, N618, N619, N620, N621, N622, N623, N624, N625,
         N626, N627, N628, N629, N630, N631, N632, N633, N634, N635, N636,
         N637, N638, N639, N640, N641, N642, N643, N644, N645, N646, N647,
         N648, N649, N650, N651, N652, N653, N654, N655, N656, N657, N658,
         N659, N660, N661, N662, N663, N664, N665, N666, N667, N668, N669,
         N671, N672, N673, N674, N675, N676, N677, N678, N679, N680, N681,
         N682, N683, N684, N685, N686, N687, N688, N689, N690, N691, N693,
         N694, N695, N696, N697, N698, N699, N700, N701, N702, N703, N704,
         N705, N706, N707, N708, N709, N710, N711, N712, N760, N761, N762,
         N763, N764, N765, N766, N767, N768, N769, N770, N771, N772, N773,
         N774, N775, N776, N777, N778, N779, N780, N781, N782, N783, N830,
         N831, N832, N833, N834, N835, N836, N837, N838, N839, N840, N841,
         N842, N843, N844, N845, N846, N847, N848, N849, N850, N851, N852,
         N853, N854, N855, N856, N857, N858, N859, N860, N861, N862, N863,
         N864, N865, N866, N867, N868, N869, N870, N871, N872, N873, N874,
         N875, N876, N877, N878, N879, N880, N881, N882, N883, N884, N885,
         N886, N887, N888, N889, N890, N891, N892, N893, N894, N895, N896,
         N897, N898, N899, N900, N901, N902, N950, N951, N952, N953, N954,
         N955, N956, N957, N958, N959, N960, N961, N962, N963, N964, N965,
         N966, N967, N968, N969, N970, N971, N972, N973, N974, N975, N976,
         N977, N978, N979, N980, N981, N982, N983, N984, N985, N986, N987,
         N988, N989, N990, N991, N992, N993, N994, N995, N996, N997, N998,
         N1045, N1046, N1047, N1048, N1049, N1050, N1051, N1052, N1053, N1054,
         N1055, N1056, N1057, N1058, N1059, N1060, N1061, N1062, N1063, N1064,
         N1065, N1066, N1067, N1068, N1093, N1094, N1095, N1096, N1097, N1098,
         N1099, N1100, N1101, N1102, N1103, N1104, N1105, N1106, N1107, N1108,
         N1109, N1110, N1111, N1112, N1113, N1114, N1115, N1116, N1117, N1118,
         N1119, N1120, N1121, N1122, N1123, N1124, N1125, N1126, N1127, N1128,
         N1129, N1130, N1131, N1132, N1133, N1134, N1135, N1136, N1137, N1138,
         N1139, N1140, N1141, N1142, N1143, N1144, N1145, N1146, N1147, N1148,
         N1149, N1150, N1151, N1152, N1153, N1154, N1155, N1156, N1157, N1158,
         N1159, N1160, N1161, N1162, N1163, N1164, N1165, N1166, N1167, N1168,
         N1169, N1170, N1171, N1172, N1173, N1174, N1175, N1176, N1177, N1178,
         N1179, N1180, N1181, N1182, N1183, N1184, N1185, N1186, N1187, N1188,
         N1189, N1190, N1191, N1192, N1193, N1194, N1195, N1196, N1197, N1198,
         N1199, N1200, N1201, N1202, N1203, N1204, N1205, N1206, N1207, N1208,
         N1209, N1210, N1211, N1212, N1213, N1214, N1215, N1216, N1217, N1218,
         N1219, N1220, N1221, N1222, N1223, N1224, N1225, N1226, N1227, N1228,
         N1229, N1230, N1231, N1232, N1233, N1234, N1235, N1236, N1237, N1238,
         N1239, N1240, N1241, N1242, N1243, N1244, N1245, N1246, N1247, N1248,
         N1249, N1250, N1251, N1252, N1253, N1254, N1255, N1256, N1257, N1258,
         N1259, N1260, N1261, N1262, N1263, N1264, N1265, N1266, N1267, N1268,
         N1269, N1270, N1271, N1272, N1273, N1274, N1275, N1276, N1277, N1278,
         N1279, N1280, N1281, N1282, N1283, N1284, N1285, N1286, N1287, N1288,
         N1289, N1290, N1291, N1292, N1293, N1294, N1295, N1296, N1297, N1298,
         N1299, N1300, N1301, N1302, N1303, N1304, N1305, N1306, N1307, N1308,
         N1309, N1310, N1311, N1312, N1313, N1314, N1315, N1316, N1317, N1318,
         N1370, N1371, N1372, N1373, N1374, N1375, N1376, N1377, N1378, N1379,
         N1380, N1381, N1382, N1383, N1384, N1385, N1386, N1387, N1388, N1389,
         N1390, N1391, N1392, N1393, N1394, N1395, N1447, N1448, N1449, N1450,
         N1451, N1452, N1453, N1454, N1455, N1456, N1457, N1458, N1459, N1460,
         N1461, N1462, N1463, N1464, N1465, N1466, N1467, N1468, N1469, N1470,
         N1471, N1472, N1524, N1525, N1526, N1527, N1528, N1529, N1530, N1531,
         N1532, N1533, N1534, N1535, N1536, N1537, N1538, N1539, N1540, N1541,
         N1542, N1543, N1544, N1545, N1546, N1547, N1548, N1549, N1601, N1602,
         N1603, N1604, N1605, N1606, N1607, N1608, N1609, N1610, N1611, N1612,
         N1613, N1614, N1615, N1616, N1617, N1618, N1619, N1620, N1621, N1622,
         N1623, N1624, N1625, N1626, N1627, N1628, N1629, N1630, N1631, N1632,
         N1633, N1634, N1635, N1636, N1637, N1638, N1639, N1640, N1641, N1642,
         N1643, N1644, N1645, N1646, N1647, N1648, N1649, N1650, N1651, N1652,
         N1653, N1654, N1655, N1656, N1657, N1658, N1659, N1660, N1661, N1662,
         N1663, N1664, N1665, N1666, N1667, N1668, N1669, N1670, N1671, N1672,
         N1673, N1674, N1675, N1676, N1677, N1678, N1679, N1680, N1681, N1682,
         N1683, N1684, N1685, N1686, N1687, N1688, N1689, N1690, N1691, N1692,
         N1693, N1694, N1695, N1696, N1697, N1698, N1699, N1700, N1701, N1702,
         N1703, N1704, N1705, N1706, N1707, N1708, N1709, N1710, N1711, N1712,
         N1713, N1714, N1715, N1716, N1717, N1718, N1719, N1720, N1721, N1722,
         N1723, N1724, N1725, N1726, N1727, N1728, N1729, N1730, N1731, N1732,
         N1733, N1734, N1735, N1736, N1737, N1738, N1739, N1740, N1741, N1742,
         N1743, N1744, N1745, N1746, N1747, N1748, N1749, N1750, N1751, N1752,
         N1753, N1754, N1755, N1756, N1757, N1758, N1759, N1760, N1761, N1762,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, N1092, N1091, N1090, N1089, N1088,
         N1087, N1086, N1085, N1084, N1083, N1082, N1081, N1080, N1079, N1078,
         N1077, N1076, N1075, N1074, N1073, N1072, N1071, N1070, N1069,
         add_187_carry_13_, add_187_carry_14_, add_187_carry_15_,
         add_187_carry_16_, add_187_carry_17_, add_187_carry_18_,
         add_187_carry_19_, add_187_carry_20_, add_187_carry_21_,
         add_187_carry_22_, add_187_carry_23_, add_187_carry_24_,
         add_187_carry_25_, add_187_carry_26_, add_187_carry_27_,
         add_186_carry_13_, add_186_carry_14_, add_186_carry_15_,
         add_186_carry_16_, add_186_carry_17_, add_186_carry_18_,
         add_186_carry_19_, add_186_carry_20_, add_186_carry_21_,
         add_186_carry_22_, add_186_carry_23_, add_186_carry_24_,
         add_186_carry_25_, add_186_carry_26_, add_186_carry_27_,
         add_185_carry_13_, add_185_carry_14_, add_185_carry_15_,
         add_185_carry_16_, add_185_carry_17_, add_185_carry_18_,
         add_185_carry_19_, add_185_carry_20_, add_185_carry_21_,
         add_185_carry_22_, add_185_carry_23_, add_185_carry_24_,
         add_185_carry_25_, add_185_carry_26_, add_185_carry_27_,
         add_184_carry_13_, add_184_carry_14_, add_184_carry_15_,
         add_184_carry_16_, add_184_carry_17_, add_184_carry_18_,
         add_184_carry_19_, add_184_carry_20_, add_184_carry_21_,
         add_184_carry_22_, add_184_carry_23_, add_184_carry_24_,
         add_184_carry_25_, add_184_carry_26_, add_184_carry_27_,
         add_183_carry_13_, add_183_carry_14_, add_183_carry_15_,
         add_183_carry_16_, add_183_carry_17_, add_183_carry_18_,
         add_183_carry_19_, add_183_carry_20_, add_183_carry_21_,
         add_183_carry_22_, add_183_carry_23_, add_183_carry_24_,
         add_183_carry_25_, add_183_carry_26_, add_183_carry_27_,
         add_182_carry_13_, add_182_carry_14_, add_182_carry_15_,
         add_182_carry_16_, add_182_carry_17_, add_182_carry_18_,
         add_182_carry_19_, add_182_carry_20_, add_182_carry_21_,
         add_182_carry_22_, add_182_carry_23_, add_182_carry_24_,
         add_182_carry_25_, add_182_carry_26_, add_182_carry_27_,
         add_181_carry_13_, add_181_carry_14_, add_181_carry_15_,
         add_181_carry_16_, add_181_carry_17_, add_181_carry_18_,
         add_181_carry_19_, add_181_carry_20_, add_181_carry_21_,
         add_181_carry_22_, add_181_carry_23_, add_181_carry_24_,
         add_181_carry_25_, add_181_carry_26_, add_181_carry_27_,
         add_180_carry_13_, add_180_carry_14_, add_180_carry_15_,
         add_180_carry_16_, add_180_carry_17_, add_180_carry_18_,
         add_180_carry_19_, add_180_carry_20_, add_180_carry_21_,
         add_180_carry_22_, add_180_carry_23_, add_180_carry_24_,
         add_180_carry_25_, add_180_carry_26_, add_180_carry_27_,
         add_104_carry_10_, add_104_carry_11_, add_104_carry_12_,
         add_104_carry_13_, add_104_carry_14_, add_104_carry_15_,
         add_104_carry_16_, add_104_carry_17_, add_104_carry_18_,
         add_104_carry_5_, add_104_carry_6_, add_104_carry_7_,
         add_104_carry_8_, add_104_carry_9_, add_102_carry_10_,
         add_102_carry_11_, add_102_carry_12_, add_102_carry_13_,
         add_102_carry_14_, add_102_carry_15_, add_102_carry_16_,
         add_102_carry_17_, add_102_carry_4_, add_102_carry_5_,
         add_102_carry_6_, add_102_carry_7_, add_102_carry_8_,
         add_102_carry_9_, add_100_carry_10_, add_100_carry_11_,
         add_100_carry_12_, add_100_carry_13_, add_100_carry_14_,
         add_100_carry_15_, add_100_carry_16_, add_100_carry_17_,
         add_100_carry_18_, add_100_carry_5_, add_100_carry_6_,
         add_100_carry_7_, add_100_carry_8_, add_100_carry_9_,
         add_99_carry_10_, add_99_carry_11_, add_99_carry_12_,
         add_99_carry_13_, add_99_carry_14_, add_99_carry_15_,
         add_99_carry_16_, add_99_carry_17_, add_99_carry_18_,
         add_99_carry_19_, add_99_carry_20_, add_99_carry_7_, add_99_carry_8_,
         add_99_carry_9_, add_95_carry_10_, add_95_carry_11_, add_95_carry_12_,
         add_95_carry_13_, add_95_carry_14_, add_95_carry_15_,
         add_95_carry_16_, add_95_carry_17_, add_95_carry_18_, add_95_carry_5_,
         add_95_carry_6_, add_95_carry_7_, add_95_carry_8_, add_95_carry_9_,
         add_93_carry_10_, add_93_carry_11_, add_93_carry_12_,
         add_93_carry_13_, add_93_carry_14_, add_93_carry_15_,
         add_93_carry_16_, add_93_carry_17_, add_93_carry_4_, add_93_carry_5_,
         add_93_carry_6_, add_93_carry_7_, add_93_carry_8_, add_93_carry_9_,
         add_91_carry_10_, add_91_carry_11_, add_91_carry_12_,
         add_91_carry_13_, add_91_carry_14_, add_91_carry_15_,
         add_91_carry_16_, add_91_carry_17_, add_91_carry_18_, add_91_carry_5_,
         add_91_carry_6_, add_91_carry_7_, add_91_carry_8_, add_91_carry_9_,
         add_90_carry_10_, add_90_carry_11_, add_90_carry_12_,
         add_90_carry_13_, add_90_carry_14_, add_90_carry_15_,
         add_90_carry_16_, add_90_carry_17_, add_90_carry_18_,
         add_90_carry_19_, add_90_carry_20_, add_90_carry_7_, add_90_carry_8_,
         add_90_carry_9_, add_86_carry_10_, add_86_carry_11_, add_86_carry_12_,
         add_86_carry_13_, add_86_carry_14_, add_86_carry_15_,
         add_86_carry_16_, add_86_carry_17_, add_86_carry_18_, add_86_carry_5_,
         add_86_carry_6_, add_86_carry_7_, add_86_carry_8_, add_86_carry_9_,
         add_84_carry_10_, add_84_carry_11_, add_84_carry_12_,
         add_84_carry_13_, add_84_carry_14_, add_84_carry_15_,
         add_84_carry_16_, add_84_carry_17_, add_84_carry_4_, add_84_carry_5_,
         add_84_carry_6_, add_84_carry_7_, add_84_carry_8_, add_84_carry_9_,
         add_82_carry_10_, add_82_carry_11_, add_82_carry_12_,
         add_82_carry_13_, add_82_carry_14_, add_82_carry_15_,
         add_82_carry_16_, add_82_carry_17_, add_82_carry_18_, add_82_carry_5_,
         add_82_carry_6_, add_82_carry_7_, add_82_carry_8_, add_82_carry_9_,
         add_81_carry_10_, add_81_carry_11_, add_81_carry_12_,
         add_81_carry_13_, add_81_carry_14_, add_81_carry_15_,
         add_81_carry_16_, add_81_carry_17_, add_81_carry_18_,
         add_81_carry_19_, add_81_carry_20_, add_81_carry_7_, add_81_carry_8_,
         add_81_carry_9_, add_77_carry_10_, add_77_carry_11_, add_77_carry_12_,
         add_77_carry_13_, add_77_carry_14_, add_77_carry_15_,
         add_77_carry_16_, add_77_carry_17_, add_77_carry_18_, add_77_carry_5_,
         add_77_carry_6_, add_77_carry_7_, add_77_carry_8_, add_77_carry_9_,
         add_75_carry_10_, add_75_carry_11_, add_75_carry_12_,
         add_75_carry_13_, add_75_carry_14_, add_75_carry_15_,
         add_75_carry_16_, add_75_carry_17_, add_75_carry_4_, add_75_carry_5_,
         add_75_carry_6_, add_75_carry_7_, add_75_carry_8_, add_75_carry_9_,
         add_73_carry_10_, add_73_carry_11_, add_73_carry_12_,
         add_73_carry_13_, add_73_carry_14_, add_73_carry_15_,
         add_73_carry_16_, add_73_carry_17_, add_73_carry_18_, add_73_carry_5_,
         add_73_carry_6_, add_73_carry_7_, add_73_carry_8_, add_73_carry_9_,
         add_72_carry_10_, add_72_carry_11_, add_72_carry_12_,
         add_72_carry_13_, add_72_carry_14_, add_72_carry_15_,
         add_72_carry_16_, add_72_carry_17_, add_72_carry_18_,
         add_72_carry_19_, add_72_carry_20_, add_72_carry_7_, add_72_carry_8_,
         add_72_carry_9_, n2, n3, n4, n5, n6, n7, n8, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375;
  wire   [1:0] mode_delay2;
  wire   [1:0] mode_delay1;
  wire   [20:0] x4_89_tmp2;
  wire   [19:0] x4_75_tmp2;
  wire   [20:0] x4_50_tmp1;
  wire   [20:0] x4_50_tmp2;
  wire   [19:0] x4_18_tmp1;
  wire   [16:0] x4_18_tmp2;
  wire   [20:0] x5_89_tmp2;
  wire   [19:0] x5_75_tmp2;
  wire   [20:0] x5_50_tmp1;
  wire   [20:0] x5_50_tmp2;
  wire   [19:0] x5_18_tmp1;
  wire   [16:0] x5_18_tmp2;
  wire   [20:0] x6_89_tmp2;
  wire   [19:0] x6_75_tmp2;
  wire   [20:0] x6_50_tmp1;
  wire   [20:0] x6_50_tmp2;
  wire   [19:0] x6_18_tmp1;
  wire   [16:0] x6_18_tmp2;
  wire   [20:0] x7_89_tmp2;
  wire   [19:0] x7_75_tmp2;
  wire   [20:0] x7_50_tmp1;
  wire   [20:0] x7_50_tmp2;
  wire   [19:0] x7_18_tmp1;
  wire   [16:0] x7_18_tmp2;
  wire   [22:0] x4_89;
  wire   [22:0] x5_89;
  wire   [22:0] x6_89;
  wire   [22:0] x7_89;
  wire   [22:0] x4_75;
  wire   [22:0] x5_75;
  wire   [22:0] x6_75;
  wire   [22:0] x7_75;
  wire   [21:0] x4_50;
  wire   [21:0] x5_50;
  wire   [21:0] x6_50;
  wire   [21:0] x7_50;
  wire   [20:0] x4_18;
  wire   [20:0] x5_18;
  wire   [20:0] x6_18;
  wire   [20:0] x7_18;
  wire   [22:0] x7_75_tmp1;
  wire   [22:0] x6_75_tmp1;
  wire   [22:0] x5_75_tmp1;
  wire   [22:0] x4_75_tmp1;
  wire   [22:0] x7_89_tmp1;
  wire   [22:0] x6_89_tmp1;
  wire   [22:0] x5_89_tmp1;
  wire   [22:0] x4_89_tmp1;
  wire   [23:0] x4_tmp1;
  wire   [23:0] x4_tmp2;
  wire   [23:0] x5_tmp1;
  wire   [23:0] x5_tmp2;
  wire   [23:0] x6_tmp1;
  wire   [23:0] x6_tmp2;
  wire   [23:0] x7_tmp1;
  wire   [23:0] x7_tmp2;
  wire   [24:0] x4_tmp;
  wire   [24:0] x5_tmp;
  wire   [24:0] x6_tmp;
  wire   [24:0] x7_tmp;
  wire   [25:0] y0_tmp;
  wire   [25:0] y1_tmp;
  wire   [25:0] y2_tmp;
  wire   [25:0] y3_tmp;
  wire   [25:0] y4_tmp;
  wire   [25:0] y5_tmp;
  wire   [25:0] y6_tmp;
  wire   [25:0] y7_tmp;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8;

  idct8_shift12_add2048_DW01_add_8 add_1_root_add_177_2 ( .A({x0[24], x0}), 
        .B({n300, n300, n299, n298, n297, n296, n295, n294, n293, n292, n291, 
        n290, n289, n288, n287, n286, n285, n284, n283, n282, n281, n280, n279, 
        n278, n277, n276}), .SUM({N1626, N1625, N1624, N1623, N1622, N1621, 
        N1620, N1619, N1618, N1617, N1616, N1615, N1614, N1613, N1612, N1611, 
        N1610, N1609, N1608, N1607, N1606, N1605, N1604, N1603, N1602, N1601})
         );
  idct8_shift12_add2048_DW01_add_9 add_1_root_add_176_2 ( .A({x1[24], x1}), 
        .B({n326, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, 
        n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, 
        n348, n349, n350}), .SUM({N1549, N1548, N1547, N1546, N1545, N1544, 
        N1543, N1542, N1541, N1540, N1539, N1538, N1537, N1536, N1535, N1534, 
        N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524})
         );
  idct8_shift12_add2048_DW01_add_10 add_1_root_add_175_2 ( .A({x2[24], x2}), 
        .B({n301, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, 
        n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, 
        n323, n324, n325}), .SUM({N1472, N1471, N1470, N1469, N1468, N1467, 
        N1466, N1465, N1464, N1463, N1462, N1461, N1460, N1459, N1458, N1457, 
        N1456, N1455, N1454, N1453, N1452, N1451, N1450, N1449, N1448, N1447})
         );
  idct8_shift12_add2048_DW01_add_11 add_1_root_add_174_2 ( .A({x3[24], x3}), 
        .B({n375, n375, n374, n373, n372, n371, n370, n369, n368, n367, n366, 
        n365, n364, n363, n362, n361, n360, n359, n358, n357, n356, n355, n354, 
        n353, n352, n351}), .SUM({N1395, N1394, N1393, N1392, N1391, N1390, 
        N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, 
        N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370})
         );
  idct8_shift12_add2048_DW01_add_12 add_173 ( .A({x3[24], x3}), .B({x4_tmp[24], 
        x4_tmp}), .SUM({N1318, N1317, N1316, N1315, N1314, N1313, N1312, N1311, 
        N1310, N1309, N1308, N1307, N1306, N1305, N1304, N1303, N1302, N1301, 
        N1300, N1299, N1298, N1297, N1296, N1295, N1294, N1293}) );
  idct8_shift12_add2048_DW01_add_13 add_172 ( .A({x2[24], x2}), .B({x5_tmp[24], 
        x5_tmp}), .SUM({N1292, N1291, N1290, N1289, N1288, N1287, N1286, N1285, 
        N1284, N1283, N1282, N1281, N1280, N1279, N1278, N1277, N1276, N1275, 
        N1274, N1273, N1272, N1271, N1270, N1269, N1268, N1267}) );
  idct8_shift12_add2048_DW01_add_14 add_171 ( .A({x1[24], x1}), .B({x6_tmp[24], 
        x6_tmp}), .SUM({N1266, N1265, N1264, N1263, N1262, N1261, N1260, N1259, 
        N1258, N1257, N1256, N1255, N1254, N1253, N1252, N1251, N1250, N1249, 
        N1248, N1247, N1246, N1245, N1244, N1243, N1242, N1241}) );
  idct8_shift12_add2048_DW01_add_15 add_170 ( .A({x0[24], x0}), .B({x7_tmp[24], 
        x7_tmp}), .SUM({N1240, N1239, N1238, N1237, N1236, N1235, N1234, N1233, 
        N1232, N1231, N1230, N1229, N1228, N1227, N1226, N1225, N1224, N1223, 
        N1222, N1221, N1220, N1219, N1218, N1217, N1216, N1215}) );
  idct8_shift12_add2048_DW01_add_16 add_157 ( .A({x7_tmp1[23], x7_tmp1}), .B({
        x7_tmp2[23], x7_tmp2}), .SUM({N1214, N1213, N1212, N1211, N1210, N1209, 
        N1208, N1207, N1206, N1205, N1204, N1203, N1202, N1201, N1200, N1199, 
        N1198, N1197, N1196, N1195, N1194, N1193, N1192, N1191, N1190}) );
  idct8_shift12_add2048_DW01_add_17 add_156 ( .A({x5_75[22], x5_75}), .B({
        x6_50[21], x6_50[21], x6_50}), .SUM({N1189, N1188, N1187, N1186, N1185, 
        N1184, N1183, N1182, N1181, N1180, N1179, N1178, N1177, N1176, N1175, 
        N1174, N1173, N1172, N1171, N1170, N1169, N1168, N1167, N1166}) );
  idct8_shift12_add2048_DW01_add_18 add_155 ( .A({x4_89[22], x4_89}), .B({
        x7_18[20], x7_18[20], x7_18[20], x7_18[20:1], 1'b0}), .SUM({N1165, 
        N1164, N1163, N1162, N1161, N1160, N1159, N1158, N1157, N1156, N1155, 
        N1154, N1153, N1152, N1151, N1150, N1149, N1148, N1147, N1146, N1145, 
        N1144, N1143, N1142}) );
  idct8_shift12_add2048_DW01_add_19 add_153 ( .A({x6_tmp1[23], x6_tmp1}), .B({
        x6_tmp2[23], x6_tmp2}), .SUM({N1141, N1140, N1139, N1138, N1137, N1136, 
        N1135, N1134, N1133, N1132, N1131, N1130, N1129, N1128, N1127, N1126, 
        N1125, N1124, N1123, N1122, N1121, N1120, N1119, N1118, N1117}) );
  idct8_shift12_add2048_DW01_add_20 add_1_root_add_151_2 ( .A({x4_75[22], 
        x4_75}), .B({n186, n186, n186, n187, n188, n189, n190, n191, n192, 
        n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, 
        n205, n206, n207}), .SUM({N1068, N1067, N1066, N1065, N1064, N1063, 
        N1062, N1061, N1060, N1059, N1058, N1057, N1056, N1055, N1054, N1053, 
        N1052, N1051, N1050, N1049, N1048, N1047, N1046, N1045}) );
  idct8_shift12_add2048_DW01_add_21 add_149 ( .A({x5_tmp1[23], x5_tmp1}), .B({
        x5_tmp2[23], x5_tmp2}), .SUM({N998, N997, N996, N995, N994, N993, N992, 
        N991, N990, N989, N988, N987, N986, N985, N984, N983, N982, N981, N980, 
        N979, N978, N977, N976, N975, N974}) );
  idct8_shift12_add2048_DW01_add_22 add_1_root_add_148_2 ( .A({x6_18[20], 
        x6_18[20], x6_18[20], x6_18[20:1], 1'b0}), .B({n208, n208, n209, n210, 
        n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, 
        n223, n224, n225, n226, n227, n228, n229, n230}), .SUM({N973, N972, 
        N971, N970, N969, N968, N967, N966, N965, N964, N963, N962, N961, N960, 
        N959, N958, N957, N956, N955, N954, N953, N952, N951, N950}) );
  idct8_shift12_add2048_DW01_add_23 add_147 ( .A({x4_50[21], x4_50[21], x4_50}), .B({x7_75[22], x7_75}), .SUM({N902, N901, N900, N899, N898, N897, N896, N895, 
        N894, N893, N892, N891, N890, N889, N888, N887, N886, N885, N884, N883, 
        N882, N881, N880, N879}) );
  idct8_shift12_add2048_DW01_add_24 add_145 ( .A({x4_tmp1[23], x4_tmp1}), .B({
        x4_tmp2[23], x4_tmp2}), .SUM({N878, N877, N876, N875, N874, N873, N872, 
        N871, N870, N869, N868, N867, N866, N865, N864, N863, N862, N861, N860, 
        N859, N858, N857, N856, N855, N854}) );
  idct8_shift12_add2048_DW01_add_25 add_1_root_add_144_2 ( .A({x6_75[22], 
        x6_75}), .B({n254, n254, n254, n255, n256, n257, n258, n259, n260, 
        n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, 
        n273, n274, n275}), .SUM({N853, N852, N851, N850, N849, N848, N847, 
        N846, N845, N844, N843, N842, N841, N840, N839, N838, N837, N836, N835, 
        N834, N833, N832, N831, N830}) );
  idct8_shift12_add2048_DW01_add_26 add_1_root_add_143_2 ( .A({x4_18[20], 
        x4_18[20], x4_18[20], x4_18[20:1], 1'b0}), .B({n231, n231, n232, n233, 
        n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, 
        n246, n247, n248, n249, n250, n251, n252, n253}), .SUM({N783, N782, 
        N781, N780, N779, N778, N777, N776, N775, N774, N773, N772, N771, N770, 
        N769, N768, N767, N766, N765, N764, N763, N762, N761, N760}) );
  idct8_shift12_add2048_DW01_add_27 add_127 ( .A({x7_18_tmp1[19], 
        x7_18_tmp1[19:4], 1'b0, 1'b0, 1'b0, 1'b0}), .B({x7_18_tmp2[16], 
        x7_18_tmp2[16], x7_18_tmp2[16], x7_18_tmp2[16], x7_18_tmp2[16:1], 1'b0}), .SUM({N712, N711, N710, N709, N708, N707, N706, N705, N704, N703, N702, 
        N701, N700, N699, N698, N697, N696, N695, N694, N693, 
        SYNOPSYS_UNCONNECTED__0}) );
  idct8_shift12_add2048_DW01_add_28 add_126 ( .A({x7_50_tmp1[20], 
        x7_50_tmp1[20:5], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({x7_50_tmp2[20], 
        x7_50_tmp2[20:1], 1'b0}), .SUM({N691, N690, N689, N688, N687, N686, 
        N685, N684, N683, N682, N681, N680, N679, N678, N677, N676, N675, N674, 
        N673, N672, N671, SYNOPSYS_UNCONNECTED__1}) );
  idct8_shift12_add2048_DW01_add_29 add_125 ( .A(x7_75_tmp1), .B({
        x7_75_tmp2[19], x7_75_tmp2[19], x7_75_tmp2[19], x7_75_tmp2[19:1], 1'b0}), .SUM({N669, N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, 
        N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647}) );
  idct8_shift12_add2048_DW01_add_30 add_124 ( .A(x7_89_tmp1), .B({
        x7_89_tmp2[20], x7_89_tmp2[20], x7_89_tmp2[20:3], 1'b0, 1'b0, 1'b0}), 
        .SUM({N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, 
        N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624}) );
  idct8_shift12_add2048_DW01_add_31 add_122 ( .A({x6_18_tmp1[19], 
        x6_18_tmp1[19:4], 1'b0, 1'b0, 1'b0, 1'b0}), .B({x6_18_tmp2[16], 
        x6_18_tmp2[16], x6_18_tmp2[16], x6_18_tmp2[16], x6_18_tmp2[16:1], 1'b0}), .SUM({N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, 
        N612, N611, N610, N609, N608, N607, N606, N605, N604, 
        SYNOPSYS_UNCONNECTED__2}) );
  idct8_shift12_add2048_DW01_add_32 add_121 ( .A({x6_50_tmp1[20], 
        x6_50_tmp1[20:5], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({x6_50_tmp2[20], 
        x6_50_tmp2[20:1], 1'b0}), .SUM({N602, N601, N600, N599, N598, N597, 
        N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, 
        N584, N583, N582, SYNOPSYS_UNCONNECTED__3}) );
  idct8_shift12_add2048_DW01_add_33 add_120 ( .A(x6_75_tmp1), .B({
        x6_75_tmp2[19], x6_75_tmp2[19], x6_75_tmp2[19], x6_75_tmp2[19:1], 1'b0}), .SUM({N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, 
        N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558}) );
  idct8_shift12_add2048_DW01_add_34 add_119 ( .A(x6_89_tmp1), .B({
        x6_89_tmp2[20], x6_89_tmp2[20], x6_89_tmp2[20:3], 1'b0, 1'b0, 1'b0}), 
        .SUM({N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, 
        N546, N545, N544, N543, N542, N541, N540, N539, N538, N537, N536, N535}) );
  idct8_shift12_add2048_DW01_add_35 add_117 ( .A({x5_18_tmp1[19], 
        x5_18_tmp1[19:4], 1'b0, 1'b0, 1'b0, 1'b0}), .B({x5_18_tmp2[16], 
        x5_18_tmp2[16], x5_18_tmp2[16], x5_18_tmp2[16], x5_18_tmp2[16:1], 1'b0}), .SUM({N534, N533, N532, N531, N530, N529, N528, N527, N526, N525, N524, 
        N523, N522, N521, N520, N519, N518, N517, N516, N515, 
        SYNOPSYS_UNCONNECTED__4}) );
  idct8_shift12_add2048_DW01_add_36 add_116 ( .A({x5_50_tmp1[20], 
        x5_50_tmp1[20:5], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({x5_50_tmp2[20], 
        x5_50_tmp2[20:1], 1'b0}), .SUM({N513, N512, N511, N510, N509, N508, 
        N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, 
        N495, N494, N493, SYNOPSYS_UNCONNECTED__5}) );
  idct8_shift12_add2048_DW01_add_37 add_115 ( .A(x5_75_tmp1), .B({
        x5_75_tmp2[19], x5_75_tmp2[19], x5_75_tmp2[19], x5_75_tmp2[19:1], 1'b0}), .SUM({N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, 
        N480, N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469}) );
  idct8_shift12_add2048_DW01_add_38 add_114 ( .A(x5_89_tmp1), .B({
        x5_89_tmp2[20], x5_89_tmp2[20], x5_89_tmp2[20:3], 1'b0, 1'b0, 1'b0}), 
        .SUM({N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, 
        N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446}) );
  idct8_shift12_add2048_DW01_add_39 add_112 ( .A({x4_18_tmp1[19], 
        x4_18_tmp1[19:4], 1'b0, 1'b0, 1'b0, 1'b0}), .B({x4_18_tmp2[16], 
        x4_18_tmp2[16], x4_18_tmp2[16], x4_18_tmp2[16], x4_18_tmp2[16:1], 1'b0}), .SUM({N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, 
        N434, N433, N432, N431, N430, N429, N428, N427, N426, 
        SYNOPSYS_UNCONNECTED__6}) );
  idct8_shift12_add2048_DW01_add_40 add_111 ( .A({x4_50_tmp1[20], 
        x4_50_tmp1[20:5], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({x4_50_tmp2[20], 
        x4_50_tmp2[20:1], 1'b0}), .SUM({N424, N423, N422, N421, N420, N419, 
        N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, 
        N406, N405, N404, SYNOPSYS_UNCONNECTED__7}) );
  idct8_shift12_add2048_DW01_add_41 add_110 ( .A(x4_75_tmp1), .B({
        x4_75_tmp2[19], x4_75_tmp2[19], x4_75_tmp2[19], x4_75_tmp2[19:1], 1'b0}), .SUM({N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, 
        N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380}) );
  idct8_shift12_add2048_DW01_add_42 add_109 ( .A(x4_89_tmp1), .B({
        x4_89_tmp2[20], x4_89_tmp2[20], x4_89_tmp2[20:3], 1'b0, 1'b0, 1'b0}), 
        .SUM({N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, 
        N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357}) );
  idct8_shift12_add2048_DW01_add_59 add_152 ( .A({1'b0, x5_18[20], x5_18[20], 
        x5_18[20], x5_18[20:1], 1'b0}), .B({1'b0, x6_89[22], x6_89}), .SUM({
        SYNOPSYS_UNCONNECTED__8, N1092, N1091, N1090, N1089, N1088, N1087, 
        N1086, N1085, N1084, N1083, N1082, N1081, N1080, N1079, N1078, N1077, 
        N1076, N1075, N1074, N1073, N1072, N1071, N1070, N1069}) );
  idct8_shift12_add2048_DW01_sub_0 sub_add_152_2_b0 ( .B({N1092, N1091, N1090, 
        N1089, N1088, N1087, N1086, N1085, N1084, N1083, N1082, N1081, N1080, 
        N1079, N1078, N1077, N1076, N1075, N1074, N1073, N1072, N1071, N1070, 
        N1069}), .DIFF({N1116, N1115, N1114, N1113, N1112, N1111, N1110, N1109, 
        N1108, N1107, N1106, N1105, N1104, N1103, N1102, N1101, N1100, N1099, 
        N1098, N1097, N1096, N1095, N1094, N1093}) );
  DFFRHQX1 x6_50_tmp2_reg_4_ ( .D(N255), .CK(clk), .RN(rstn), .Q(x6_50_tmp2[4]) );
  DFFRHQX1 x6_50_tmp2_reg_3_ ( .D(n42), .CK(clk), .RN(rstn), .Q(x6_50_tmp2[3])
         );
  DFFRHQX1 x6_50_tmp2_reg_2_ ( .D(x6[1]), .CK(clk), .RN(rstn), .Q(
        x6_50_tmp2[2]) );
  DFFRHQX1 x6_50_tmp2_reg_1_ ( .D(x6[0]), .CK(clk), .RN(rstn), .Q(
        x6_50_tmp2[1]) );
  DFFRHQX1 x5_50_tmp2_reg_4_ ( .D(N170), .CK(clk), .RN(rstn), .Q(x5_50_tmp2[4]) );
  DFFRHQX1 x5_50_tmp2_reg_3_ ( .D(n55), .CK(clk), .RN(rstn), .Q(x5_50_tmp2[3])
         );
  DFFRHQX1 x5_50_tmp2_reg_2_ ( .D(x5[1]), .CK(clk), .RN(rstn), .Q(
        x5_50_tmp2[2]) );
  DFFRHQX1 x5_50_tmp2_reg_1_ ( .D(x5[0]), .CK(clk), .RN(rstn), .Q(
        x5_50_tmp2[1]) );
  DFFRHQX1 x7_50_tmp2_reg_4_ ( .D(N340), .CK(clk), .RN(rstn), .Q(x7_50_tmp2[4]) );
  DFFRHQX1 x7_50_tmp2_reg_3_ ( .D(n2), .CK(clk), .RN(rstn), .Q(x7_50_tmp2[3])
         );
  DFFRHQX1 x7_50_tmp2_reg_2_ ( .D(x7[1]), .CK(clk), .RN(rstn), .Q(
        x7_50_tmp2[2]) );
  DFFRHQX1 x7_50_tmp2_reg_1_ ( .D(x7[0]), .CK(clk), .RN(rstn), .Q(
        x7_50_tmp2[1]) );
  DFFRHQX1 x6_18_tmp2_reg_3_ ( .D(n42), .CK(clk), .RN(rstn), .Q(x6_18_tmp2[3])
         );
  DFFRHQX1 x6_18_tmp2_reg_2_ ( .D(x6[1]), .CK(clk), .RN(rstn), .Q(
        x6_18_tmp2[2]) );
  DFFRHQX1 x6_18_tmp2_reg_1_ ( .D(x6[0]), .CK(clk), .RN(rstn), .Q(
        x6_18_tmp2[1]) );
  DFFRHQX1 x5_18_tmp2_reg_3_ ( .D(n55), .CK(clk), .RN(rstn), .Q(x5_18_tmp2[3])
         );
  DFFRHQX1 x5_18_tmp2_reg_2_ ( .D(x5[1]), .CK(clk), .RN(rstn), .Q(
        x5_18_tmp2[2]) );
  DFFRHQX1 x5_18_tmp2_reg_1_ ( .D(x5[0]), .CK(clk), .RN(rstn), .Q(
        x5_18_tmp2[1]) );
  DFFRHQX1 x7_18_tmp2_reg_3_ ( .D(n2), .CK(clk), .RN(rstn), .Q(x7_18_tmp2[3])
         );
  DFFRHQX1 x7_18_tmp2_reg_2_ ( .D(x7[1]), .CK(clk), .RN(rstn), .Q(
        x7_18_tmp2[2]) );
  DFFRHQX1 x7_18_tmp2_reg_1_ ( .D(x7[0]), .CK(clk), .RN(rstn), .Q(
        x7_18_tmp2[1]) );
  DFFRHQX1 x4_50_tmp2_reg_4_ ( .D(N85), .CK(clk), .RN(rstn), .Q(x4_50_tmp2[4])
         );
  DFFRHQX1 x4_50_tmp2_reg_3_ ( .D(n68), .CK(clk), .RN(rstn), .Q(x4_50_tmp2[3])
         );
  DFFRHQX1 x4_50_tmp2_reg_2_ ( .D(x4[1]), .CK(clk), .RN(rstn), .Q(
        x4_50_tmp2[2]) );
  DFFRHQX1 x4_50_tmp2_reg_1_ ( .D(x4[0]), .CK(clk), .RN(rstn), .Q(
        x4_50_tmp2[1]) );
  DFFRHQX1 x4_18_tmp2_reg_3_ ( .D(n68), .CK(clk), .RN(rstn), .Q(x4_18_tmp2[3])
         );
  DFFRHQX1 x4_18_tmp2_reg_2_ ( .D(x4[1]), .CK(clk), .RN(rstn), .Q(
        x4_18_tmp2[2]) );
  DFFRHQX1 x4_18_tmp2_reg_1_ ( .D(x4[0]), .CK(clk), .RN(rstn), .Q(
        x4_18_tmp2[1]) );
  DFFRHQX1 x7_89_tmp1_reg_22_ ( .D(x7[15]), .CK(clk), .RN(rstn), .Q(
        x7_89_tmp1[22]) );
  DFFRHQX1 x7_89_tmp1_reg_21_ ( .D(N293), .CK(clk), .RN(rstn), .Q(
        x7_89_tmp1[21]) );
  DFFRHQX1 x7_89_tmp1_reg_20_ ( .D(N292), .CK(clk), .RN(rstn), .Q(
        x7_89_tmp1[20]) );
  DFFRHQX1 x7_89_tmp1_reg_19_ ( .D(N291), .CK(clk), .RN(rstn), .Q(
        x7_89_tmp1[19]) );
  DFFRHQX1 x6_89_tmp1_reg_22_ ( .D(x6[15]), .CK(clk), .RN(rstn), .Q(
        x6_89_tmp1[22]) );
  DFFRHQX1 x6_89_tmp1_reg_21_ ( .D(N208), .CK(clk), .RN(rstn), .Q(
        x6_89_tmp1[21]) );
  DFFRHQX1 x6_89_tmp1_reg_20_ ( .D(N207), .CK(clk), .RN(rstn), .Q(
        x6_89_tmp1[20]) );
  DFFRHQX1 x6_89_tmp1_reg_19_ ( .D(N206), .CK(clk), .RN(rstn), .Q(
        x6_89_tmp1[19]) );
  DFFRHQX1 x5_89_tmp1_reg_22_ ( .D(x5[15]), .CK(clk), .RN(rstn), .Q(
        x5_89_tmp1[22]) );
  DFFRHQX1 x5_89_tmp1_reg_21_ ( .D(N123), .CK(clk), .RN(rstn), .Q(
        x5_89_tmp1[21]) );
  DFFRHQX1 x5_89_tmp1_reg_20_ ( .D(N122), .CK(clk), .RN(rstn), .Q(
        x5_89_tmp1[20]) );
  DFFRHQX1 x5_89_tmp1_reg_19_ ( .D(N121), .CK(clk), .RN(rstn), .Q(
        x5_89_tmp1[19]) );
  DFFRHQX1 x5_75_tmp1_reg_22_ ( .D(x5[15]), .CK(clk), .RN(rstn), .Q(
        x5_75_tmp1[22]) );
  DFFRHQX1 x5_75_tmp1_reg_21_ ( .D(N123), .CK(clk), .RN(rstn), .Q(
        x5_75_tmp1[21]) );
  DFFRHQX1 x5_75_tmp1_reg_20_ ( .D(N122), .CK(clk), .RN(rstn), .Q(
        x5_75_tmp1[20]) );
  DFFRHQX1 x5_75_tmp1_reg_19_ ( .D(N121), .CK(clk), .RN(rstn), .Q(
        x5_75_tmp1[19]) );
  DFFRHQX1 x4_75_tmp1_reg_22_ ( .D(x4[15]), .CK(clk), .RN(rstn), .Q(
        x4_75_tmp1[22]) );
  DFFRHQX1 x4_75_tmp1_reg_21_ ( .D(N38), .CK(clk), .RN(rstn), .Q(
        x4_75_tmp1[21]) );
  DFFRHQX1 x4_75_tmp1_reg_20_ ( .D(N37), .CK(clk), .RN(rstn), .Q(
        x4_75_tmp1[20]) );
  DFFRHQX1 x4_75_tmp1_reg_19_ ( .D(N36), .CK(clk), .RN(rstn), .Q(
        x4_75_tmp1[19]) );
  DFFRHQX1 x7_75_tmp1_reg_22_ ( .D(x7[15]), .CK(clk), .RN(rstn), .Q(
        x7_75_tmp1[22]) );
  DFFRHQX1 x7_75_tmp1_reg_21_ ( .D(N293), .CK(clk), .RN(rstn), .Q(
        x7_75_tmp1[21]) );
  DFFRHQX1 x7_75_tmp1_reg_20_ ( .D(N292), .CK(clk), .RN(rstn), .Q(
        x7_75_tmp1[20]) );
  DFFRHQX1 x7_75_tmp1_reg_19_ ( .D(N291), .CK(clk), .RN(rstn), .Q(
        x7_75_tmp1[19]) );
  DFFRHQX1 x6_75_tmp1_reg_22_ ( .D(x6[15]), .CK(clk), .RN(rstn), .Q(
        x6_75_tmp1[22]) );
  DFFRHQX1 x6_75_tmp1_reg_21_ ( .D(N208), .CK(clk), .RN(rstn), .Q(
        x6_75_tmp1[21]) );
  DFFRHQX1 x6_75_tmp1_reg_20_ ( .D(N207), .CK(clk), .RN(rstn), .Q(
        x6_75_tmp1[20]) );
  DFFRHQX1 x6_75_tmp1_reg_19_ ( .D(N206), .CK(clk), .RN(rstn), .Q(
        x6_75_tmp1[19]) );
  DFFRHQX1 x4_50_tmp1_reg_19_ ( .D(n80), .CK(clk), .RN(rstn), .Q(
        x4_50_tmp1[19]) );
  DFFRHQX1 x4_50_tmp1_reg_18_ ( .D(n79), .CK(clk), .RN(rstn), .Q(
        x4_50_tmp1[18]) );
  DFFRHQX1 x6_50_tmp1_reg_19_ ( .D(n54), .CK(clk), .RN(rstn), .Q(
        x6_50_tmp1[19]) );
  DFFRHQX1 x6_50_tmp1_reg_18_ ( .D(n53), .CK(clk), .RN(rstn), .Q(
        x6_50_tmp1[18]) );
  DFFRHQX1 x5_50_tmp1_reg_19_ ( .D(n67), .CK(clk), .RN(rstn), .Q(
        x5_50_tmp1[19]) );
  DFFRHQX1 x5_50_tmp1_reg_18_ ( .D(n66), .CK(clk), .RN(rstn), .Q(
        x5_50_tmp1[18]) );
  DFFRHQX1 x7_50_tmp1_reg_19_ ( .D(n41), .CK(clk), .RN(rstn), .Q(
        x7_50_tmp1[19]) );
  DFFRHQX1 x7_50_tmp1_reg_18_ ( .D(n40), .CK(clk), .RN(rstn), .Q(
        x7_50_tmp1[18]) );
  DFFRHQX1 x4_18_tmp1_reg_18_ ( .D(n80), .CK(clk), .RN(rstn), .Q(
        x4_18_tmp1[18]) );
  DFFRHQX1 x4_18_tmp1_reg_17_ ( .D(n79), .CK(clk), .RN(rstn), .Q(
        x4_18_tmp1[17]) );
  DFFRHQX1 x5_18_tmp1_reg_18_ ( .D(n67), .CK(clk), .RN(rstn), .Q(
        x5_18_tmp1[18]) );
  DFFRHQX1 x5_18_tmp1_reg_17_ ( .D(n66), .CK(clk), .RN(rstn), .Q(
        x5_18_tmp1[17]) );
  DFFRHQX1 x6_18_tmp1_reg_18_ ( .D(n54), .CK(clk), .RN(rstn), .Q(
        x6_18_tmp1[18]) );
  DFFRHQX1 x6_18_tmp1_reg_17_ ( .D(n53), .CK(clk), .RN(rstn), .Q(
        x6_18_tmp1[17]) );
  DFFRHQX1 x7_18_tmp1_reg_18_ ( .D(n41), .CK(clk), .RN(rstn), .Q(
        x7_18_tmp1[18]) );
  DFFRHQX1 x7_18_tmp1_reg_17_ ( .D(n40), .CK(clk), .RN(rstn), .Q(
        x7_18_tmp1[17]) );
  DFFRHQX1 x4_89_tmp1_reg_22_ ( .D(x4[15]), .CK(clk), .RN(rstn), .Q(
        x4_89_tmp1[22]) );
  DFFRHQX1 x4_89_tmp1_reg_21_ ( .D(N38), .CK(clk), .RN(rstn), .Q(
        x4_89_tmp1[21]) );
  DFFRHQX1 x4_89_tmp1_reg_20_ ( .D(N37), .CK(clk), .RN(rstn), .Q(
        x4_89_tmp1[20]) );
  DFFRHQX1 x4_89_tmp1_reg_19_ ( .D(N36), .CK(clk), .RN(rstn), .Q(
        x4_89_tmp1[19]) );
  DFFRHQX1 x4_89_reg_21_ ( .D(N378), .CK(clk), .RN(rstn), .Q(x4_89[21]) );
  DFFRHQX1 x4_89_reg_20_ ( .D(N377), .CK(clk), .RN(rstn), .Q(x4_89[20]) );
  DFFRHQX1 x4_75_reg_21_ ( .D(N401), .CK(clk), .RN(rstn), .Q(x4_75[21]) );
  DFFRHQX1 x4_75_reg_20_ ( .D(N400), .CK(clk), .RN(rstn), .Q(x4_75[20]) );
  DFFRHQX1 x5_75_reg_21_ ( .D(N490), .CK(clk), .RN(rstn), .Q(x5_75[21]) );
  DFFRHQX1 x5_75_reg_20_ ( .D(N489), .CK(clk), .RN(rstn), .Q(x5_75[20]) );
  DFFRHQX1 x6_75_reg_21_ ( .D(N579), .CK(clk), .RN(rstn), .Q(x6_75[21]) );
  DFFRHQX1 x6_75_reg_20_ ( .D(N578), .CK(clk), .RN(rstn), .Q(x6_75[20]) );
  DFFRHQX1 x4_50_reg_20_ ( .D(N423), .CK(clk), .RN(rstn), .Q(x4_50[20]) );
  DFFRHQX1 x5_tmp1_reg_22_ ( .D(N901), .CK(clk), .RN(rstn), .Q(x5_tmp1[22]) );
  DFFRHQX1 x5_tmp1_reg_21_ ( .D(N900), .CK(clk), .RN(rstn), .Q(x5_tmp1[21]) );
  DFFRHQX1 x6_tmp1_reg_22_ ( .D(N1067), .CK(clk), .RN(rstn), .Q(x6_tmp1[22])
         );
  DFFRHQX1 x6_tmp1_reg_21_ ( .D(N1066), .CK(clk), .RN(rstn), .Q(x6_tmp1[21])
         );
  DFFRHQX1 x7_tmp1_reg_22_ ( .D(N1164), .CK(clk), .RN(rstn), .Q(x7_tmp1[22])
         );
  DFFRHQX1 x7_tmp1_reg_21_ ( .D(N1163), .CK(clk), .RN(rstn), .Q(x7_tmp1[21])
         );
  DFFRHQX1 x4_tmp1_reg_22_ ( .D(N782), .CK(clk), .RN(rstn), .Q(x4_tmp1[22]) );
  DFFRHQX1 x4_tmp1_reg_21_ ( .D(N781), .CK(clk), .RN(rstn), .Q(x4_tmp1[21]) );
  DFFRHQX1 y6_tmp_reg_10_ ( .D(N1534), .CK(clk), .RN(rstn), .Q(y6_tmp[10]) );
  DFFRHQX1 y6_tmp_reg_9_ ( .D(N1533), .CK(clk), .RN(rstn), .Q(y6_tmp[9]) );
  DFFRHQX1 y6_tmp_reg_8_ ( .D(N1532), .CK(clk), .RN(rstn), .Q(y6_tmp[8]) );
  DFFRHQX1 y6_tmp_reg_7_ ( .D(N1531), .CK(clk), .RN(rstn), .Q(y6_tmp[7]) );
  DFFRHQX1 y6_tmp_reg_6_ ( .D(N1530), .CK(clk), .RN(rstn), .Q(y6_tmp[6]) );
  DFFRHQX1 y6_tmp_reg_5_ ( .D(N1529), .CK(clk), .RN(rstn), .Q(y6_tmp[5]) );
  DFFRHQX1 y6_tmp_reg_4_ ( .D(N1528), .CK(clk), .RN(rstn), .Q(y6_tmp[4]) );
  DFFRHQX1 y6_tmp_reg_3_ ( .D(N1527), .CK(clk), .RN(rstn), .Q(y6_tmp[3]) );
  DFFRHQX1 y6_tmp_reg_2_ ( .D(N1526), .CK(clk), .RN(rstn), .Q(y6_tmp[2]) );
  DFFRHQX1 y6_tmp_reg_1_ ( .D(N1525), .CK(clk), .RN(rstn), .Q(y6_tmp[1]) );
  DFFRHQX1 y6_tmp_reg_0_ ( .D(N1524), .CK(clk), .RN(rstn), .Q(y6_tmp[0]) );
  DFFRHQX1 y7_tmp_reg_10_ ( .D(N1611), .CK(clk), .RN(rstn), .Q(y7_tmp[10]) );
  DFFRHQX1 y7_tmp_reg_9_ ( .D(N1610), .CK(clk), .RN(rstn), .Q(y7_tmp[9]) );
  DFFRHQX1 y7_tmp_reg_8_ ( .D(N1609), .CK(clk), .RN(rstn), .Q(y7_tmp[8]) );
  DFFRHQX1 y7_tmp_reg_7_ ( .D(N1608), .CK(clk), .RN(rstn), .Q(y7_tmp[7]) );
  DFFRHQX1 y7_tmp_reg_6_ ( .D(N1607), .CK(clk), .RN(rstn), .Q(y7_tmp[6]) );
  DFFRHQX1 y7_tmp_reg_5_ ( .D(N1606), .CK(clk), .RN(rstn), .Q(y7_tmp[5]) );
  DFFRHQX1 y7_tmp_reg_4_ ( .D(N1605), .CK(clk), .RN(rstn), .Q(y7_tmp[4]) );
  DFFRHQX1 y7_tmp_reg_3_ ( .D(N1604), .CK(clk), .RN(rstn), .Q(y7_tmp[3]) );
  DFFRHQX1 y7_tmp_reg_2_ ( .D(N1603), .CK(clk), .RN(rstn), .Q(y7_tmp[2]) );
  DFFRHQX1 y7_tmp_reg_1_ ( .D(N1602), .CK(clk), .RN(rstn), .Q(y7_tmp[1]) );
  DFFRHQX1 y7_tmp_reg_0_ ( .D(N1601), .CK(clk), .RN(rstn), .Q(y7_tmp[0]) );
  DFFRHQX1 y0_tmp_reg_10_ ( .D(N1225), .CK(clk), .RN(rstn), .Q(y0_tmp[10]) );
  DFFRHQX1 y0_tmp_reg_9_ ( .D(N1224), .CK(clk), .RN(rstn), .Q(y0_tmp[9]) );
  DFFRHQX1 y0_tmp_reg_8_ ( .D(N1223), .CK(clk), .RN(rstn), .Q(y0_tmp[8]) );
  DFFRHQX1 y0_tmp_reg_7_ ( .D(N1222), .CK(clk), .RN(rstn), .Q(y0_tmp[7]) );
  DFFRHQX1 y0_tmp_reg_6_ ( .D(N1221), .CK(clk), .RN(rstn), .Q(y0_tmp[6]) );
  DFFRHQX1 y0_tmp_reg_5_ ( .D(N1220), .CK(clk), .RN(rstn), .Q(y0_tmp[5]) );
  DFFRHQX1 y0_tmp_reg_4_ ( .D(N1219), .CK(clk), .RN(rstn), .Q(y0_tmp[4]) );
  DFFRHQX1 y0_tmp_reg_3_ ( .D(N1218), .CK(clk), .RN(rstn), .Q(y0_tmp[3]) );
  DFFRHQX1 y0_tmp_reg_2_ ( .D(N1217), .CK(clk), .RN(rstn), .Q(y0_tmp[2]) );
  DFFRHQX1 y0_tmp_reg_1_ ( .D(N1216), .CK(clk), .RN(rstn), .Q(y0_tmp[1]) );
  DFFRHQX1 y0_tmp_reg_0_ ( .D(N1215), .CK(clk), .RN(rstn), .Q(y0_tmp[0]) );
  DFFRHQX1 y1_tmp_reg_10_ ( .D(N1251), .CK(clk), .RN(rstn), .Q(y1_tmp[10]) );
  DFFRHQX1 y1_tmp_reg_9_ ( .D(N1250), .CK(clk), .RN(rstn), .Q(y1_tmp[9]) );
  DFFRHQX1 y1_tmp_reg_8_ ( .D(N1249), .CK(clk), .RN(rstn), .Q(y1_tmp[8]) );
  DFFRHQX1 y1_tmp_reg_7_ ( .D(N1248), .CK(clk), .RN(rstn), .Q(y1_tmp[7]) );
  DFFRHQX1 y1_tmp_reg_6_ ( .D(N1247), .CK(clk), .RN(rstn), .Q(y1_tmp[6]) );
  DFFRHQX1 y1_tmp_reg_5_ ( .D(N1246), .CK(clk), .RN(rstn), .Q(y1_tmp[5]) );
  DFFRHQX1 y1_tmp_reg_4_ ( .D(N1245), .CK(clk), .RN(rstn), .Q(y1_tmp[4]) );
  DFFRHQX1 y1_tmp_reg_3_ ( .D(N1244), .CK(clk), .RN(rstn), .Q(y1_tmp[3]) );
  DFFRHQX1 y1_tmp_reg_2_ ( .D(N1243), .CK(clk), .RN(rstn), .Q(y1_tmp[2]) );
  DFFRHQX1 y1_tmp_reg_1_ ( .D(N1242), .CK(clk), .RN(rstn), .Q(y1_tmp[1]) );
  DFFRHQX1 y1_tmp_reg_0_ ( .D(N1241), .CK(clk), .RN(rstn), .Q(y1_tmp[0]) );
  DFFRHQX1 y2_tmp_reg_10_ ( .D(N1277), .CK(clk), .RN(rstn), .Q(y2_tmp[10]) );
  DFFRHQX1 y2_tmp_reg_9_ ( .D(N1276), .CK(clk), .RN(rstn), .Q(y2_tmp[9]) );
  DFFRHQX1 y2_tmp_reg_8_ ( .D(N1275), .CK(clk), .RN(rstn), .Q(y2_tmp[8]) );
  DFFRHQX1 y2_tmp_reg_7_ ( .D(N1274), .CK(clk), .RN(rstn), .Q(y2_tmp[7]) );
  DFFRHQX1 y2_tmp_reg_6_ ( .D(N1273), .CK(clk), .RN(rstn), .Q(y2_tmp[6]) );
  DFFRHQX1 y2_tmp_reg_5_ ( .D(N1272), .CK(clk), .RN(rstn), .Q(y2_tmp[5]) );
  DFFRHQX1 y2_tmp_reg_4_ ( .D(N1271), .CK(clk), .RN(rstn), .Q(y2_tmp[4]) );
  DFFRHQX1 y2_tmp_reg_3_ ( .D(N1270), .CK(clk), .RN(rstn), .Q(y2_tmp[3]) );
  DFFRHQX1 y2_tmp_reg_2_ ( .D(N1269), .CK(clk), .RN(rstn), .Q(y2_tmp[2]) );
  DFFRHQX1 y2_tmp_reg_1_ ( .D(N1268), .CK(clk), .RN(rstn), .Q(y2_tmp[1]) );
  DFFRHQX1 y2_tmp_reg_0_ ( .D(N1267), .CK(clk), .RN(rstn), .Q(y2_tmp[0]) );
  DFFRHQX1 y3_tmp_reg_10_ ( .D(N1303), .CK(clk), .RN(rstn), .Q(y3_tmp[10]) );
  DFFRHQX1 y3_tmp_reg_9_ ( .D(N1302), .CK(clk), .RN(rstn), .Q(y3_tmp[9]) );
  DFFRHQX1 y3_tmp_reg_8_ ( .D(N1301), .CK(clk), .RN(rstn), .Q(y3_tmp[8]) );
  DFFRHQX1 y3_tmp_reg_7_ ( .D(N1300), .CK(clk), .RN(rstn), .Q(y3_tmp[7]) );
  DFFRHQX1 y3_tmp_reg_6_ ( .D(N1299), .CK(clk), .RN(rstn), .Q(y3_tmp[6]) );
  DFFRHQX1 y3_tmp_reg_5_ ( .D(N1298), .CK(clk), .RN(rstn), .Q(y3_tmp[5]) );
  DFFRHQX1 y3_tmp_reg_4_ ( .D(N1297), .CK(clk), .RN(rstn), .Q(y3_tmp[4]) );
  DFFRHQX1 y3_tmp_reg_3_ ( .D(N1296), .CK(clk), .RN(rstn), .Q(y3_tmp[3]) );
  DFFRHQX1 y3_tmp_reg_2_ ( .D(N1295), .CK(clk), .RN(rstn), .Q(y3_tmp[2]) );
  DFFRHQX1 y3_tmp_reg_1_ ( .D(N1294), .CK(clk), .RN(rstn), .Q(y3_tmp[1]) );
  DFFRHQX1 y3_tmp_reg_0_ ( .D(N1293), .CK(clk), .RN(rstn), .Q(y3_tmp[0]) );
  DFFRHQX1 y4_tmp_reg_10_ ( .D(N1380), .CK(clk), .RN(rstn), .Q(y4_tmp[10]) );
  DFFRHQX1 y4_tmp_reg_9_ ( .D(N1379), .CK(clk), .RN(rstn), .Q(y4_tmp[9]) );
  DFFRHQX1 y4_tmp_reg_8_ ( .D(N1378), .CK(clk), .RN(rstn), .Q(y4_tmp[8]) );
  DFFRHQX1 y4_tmp_reg_7_ ( .D(N1377), .CK(clk), .RN(rstn), .Q(y4_tmp[7]) );
  DFFRHQX1 y4_tmp_reg_6_ ( .D(N1376), .CK(clk), .RN(rstn), .Q(y4_tmp[6]) );
  DFFRHQX1 y4_tmp_reg_5_ ( .D(N1375), .CK(clk), .RN(rstn), .Q(y4_tmp[5]) );
  DFFRHQX1 y4_tmp_reg_4_ ( .D(N1374), .CK(clk), .RN(rstn), .Q(y4_tmp[4]) );
  DFFRHQX1 y4_tmp_reg_3_ ( .D(N1373), .CK(clk), .RN(rstn), .Q(y4_tmp[3]) );
  DFFRHQX1 y4_tmp_reg_2_ ( .D(N1372), .CK(clk), .RN(rstn), .Q(y4_tmp[2]) );
  DFFRHQX1 y4_tmp_reg_1_ ( .D(N1371), .CK(clk), .RN(rstn), .Q(y4_tmp[1]) );
  DFFRHQX1 y4_tmp_reg_0_ ( .D(N1370), .CK(clk), .RN(rstn), .Q(y4_tmp[0]) );
  DFFRHQX1 y5_tmp_reg_10_ ( .D(N1457), .CK(clk), .RN(rstn), .Q(y5_tmp[10]) );
  DFFRHQX1 y5_tmp_reg_9_ ( .D(N1456), .CK(clk), .RN(rstn), .Q(y5_tmp[9]) );
  DFFRHQX1 y5_tmp_reg_8_ ( .D(N1455), .CK(clk), .RN(rstn), .Q(y5_tmp[8]) );
  DFFRHQX1 y5_tmp_reg_7_ ( .D(N1454), .CK(clk), .RN(rstn), .Q(y5_tmp[7]) );
  DFFRHQX1 y5_tmp_reg_6_ ( .D(N1453), .CK(clk), .RN(rstn), .Q(y5_tmp[6]) );
  DFFRHQX1 y5_tmp_reg_5_ ( .D(N1452), .CK(clk), .RN(rstn), .Q(y5_tmp[5]) );
  DFFRHQX1 y5_tmp_reg_4_ ( .D(N1451), .CK(clk), .RN(rstn), .Q(y5_tmp[4]) );
  DFFRHQX1 y5_tmp_reg_3_ ( .D(N1450), .CK(clk), .RN(rstn), .Q(y5_tmp[3]) );
  DFFRHQX1 y5_tmp_reg_2_ ( .D(N1449), .CK(clk), .RN(rstn), .Q(y5_tmp[2]) );
  DFFRHQX1 y5_tmp_reg_1_ ( .D(N1448), .CK(clk), .RN(rstn), .Q(y5_tmp[1]) );
  DFFRHQX1 y5_tmp_reg_0_ ( .D(N1447), .CK(clk), .RN(rstn), .Q(y5_tmp[0]) );
  DFFRHQX1 x7_50_reg_21_ ( .D(N691), .CK(clk), .RN(rstn), .Q(x7_50[21]) );
  DFFRHQX1 x7_50_reg_20_ ( .D(N690), .CK(clk), .RN(rstn), .Q(x7_50[20]) );
  DFFRHQX1 x5_89_reg_22_ ( .D(N468), .CK(clk), .RN(rstn), .Q(x5_89[22]) );
  DFFRHQX1 x5_89_reg_21_ ( .D(N467), .CK(clk), .RN(rstn), .Q(x5_89[21]) );
  DFFRHQX1 x5_89_reg_20_ ( .D(N466), .CK(clk), .RN(rstn), .Q(x5_89[20]) );
  DFFRHQX1 x7_89_reg_22_ ( .D(N646), .CK(clk), .RN(rstn), .Q(x7_89[22]) );
  DFFRHQX1 x7_89_reg_21_ ( .D(N645), .CK(clk), .RN(rstn), .Q(x7_89[21]) );
  DFFRHQX1 x7_89_reg_20_ ( .D(N644), .CK(clk), .RN(rstn), .Q(x7_89[20]) );
  DFFRHQX1 x5_50_reg_21_ ( .D(N513), .CK(clk), .RN(rstn), .Q(x5_50[21]) );
  DFFRHQX1 x5_50_reg_20_ ( .D(N512), .CK(clk), .RN(rstn), .Q(x5_50[20]) );
  DFFRHQX1 x4_50_tmp1_reg_20_ ( .D(x4[15]), .CK(clk), .RN(rstn), .Q(
        x4_50_tmp1[20]) );
  DFFRHQX1 x6_50_tmp1_reg_20_ ( .D(x6[15]), .CK(clk), .RN(rstn), .Q(
        x6_50_tmp1[20]) );
  DFFRHQX1 x5_50_tmp1_reg_20_ ( .D(x5[15]), .CK(clk), .RN(rstn), .Q(
        x5_50_tmp1[20]) );
  DFFRHQX1 x7_50_tmp1_reg_20_ ( .D(x7[15]), .CK(clk), .RN(rstn), .Q(
        x7_50_tmp1[20]) );
  DFFRHQX1 x4_18_tmp1_reg_19_ ( .D(x4[15]), .CK(clk), .RN(rstn), .Q(
        x4_18_tmp1[19]) );
  DFFRHQX1 x5_18_tmp1_reg_19_ ( .D(x5[15]), .CK(clk), .RN(rstn), .Q(
        x5_18_tmp1[19]) );
  DFFRHQX1 x6_18_tmp1_reg_19_ ( .D(x6[15]), .CK(clk), .RN(rstn), .Q(
        x6_18_tmp1[19]) );
  DFFRHQX1 x7_18_tmp1_reg_19_ ( .D(x7[15]), .CK(clk), .RN(rstn), .Q(
        x7_18_tmp1[19]) );
  DFFRHQX1 x4_89_reg_22_ ( .D(N379), .CK(clk), .RN(rstn), .Q(x4_89[22]) );
  DFFRHQX1 x4_75_reg_22_ ( .D(N402), .CK(clk), .RN(rstn), .Q(x4_75[22]) );
  DFFRHQX1 x5_75_reg_22_ ( .D(N491), .CK(clk), .RN(rstn), .Q(x5_75[22]) );
  DFFRHQX1 x6_75_reg_22_ ( .D(N580), .CK(clk), .RN(rstn), .Q(x6_75[22]) );
  DFFRHQX1 x5_tmp1_reg_23_ ( .D(N902), .CK(clk), .RN(rstn), .Q(x5_tmp1[23]) );
  DFFRHQX1 x6_tmp1_reg_23_ ( .D(N1068), .CK(clk), .RN(rstn), .Q(x6_tmp1[23])
         );
  DFFRHQX1 x7_tmp1_reg_23_ ( .D(N1165), .CK(clk), .RN(rstn), .Q(x7_tmp1[23])
         );
  DFFRHQX1 x4_tmp1_reg_23_ ( .D(N783), .CK(clk), .RN(rstn), .Q(x4_tmp1[23]) );
  DFFRHQX1 x6_89_tmp2_reg_19_ ( .D(N229), .CK(clk), .RN(rstn), .Q(
        x6_89_tmp2[19]) );
  DFFRHQX1 x5_89_tmp2_reg_19_ ( .D(N144), .CK(clk), .RN(rstn), .Q(
        x5_89_tmp2[19]) );
  DFFRHQX1 x4_89_tmp2_reg_19_ ( .D(N59), .CK(clk), .RN(rstn), .Q(
        x4_89_tmp2[19]) );
  DFFRHQX1 x7_89_tmp2_reg_19_ ( .D(N314), .CK(clk), .RN(rstn), .Q(
        x7_89_tmp2[19]) );
  DFFRHQX1 x4_50_tmp2_reg_19_ ( .D(N100), .CK(clk), .RN(rstn), .Q(
        x4_50_tmp2[19]) );
  DFFRHQX1 x4_50_tmp2_reg_18_ ( .D(N99), .CK(clk), .RN(rstn), .Q(
        x4_50_tmp2[18]) );
  DFFRHQX1 x6_50_tmp2_reg_19_ ( .D(N270), .CK(clk), .RN(rstn), .Q(
        x6_50_tmp2[19]) );
  DFFRHQX1 x6_50_tmp2_reg_18_ ( .D(N269), .CK(clk), .RN(rstn), .Q(
        x6_50_tmp2[18]) );
  DFFRHQX1 x6_50_reg_20_ ( .D(N601), .CK(clk), .RN(rstn), .Q(x6_50[20]) );
  DFFRHQX1 x5_50_tmp2_reg_19_ ( .D(N185), .CK(clk), .RN(rstn), .Q(
        x5_50_tmp2[19]) );
  DFFRHQX1 x5_50_tmp2_reg_18_ ( .D(N184), .CK(clk), .RN(rstn), .Q(
        x5_50_tmp2[18]) );
  DFFRHQX1 x7_50_tmp2_reg_19_ ( .D(N355), .CK(clk), .RN(rstn), .Q(
        x7_50_tmp2[19]) );
  DFFRHQX1 x7_50_tmp2_reg_18_ ( .D(N354), .CK(clk), .RN(rstn), .Q(
        x7_50_tmp2[18]) );
  DFFRHQX1 x6_89_reg_21_ ( .D(N556), .CK(clk), .RN(rstn), .Q(x6_89[21]) );
  DFFRHQX1 x7_75_reg_21_ ( .D(N668), .CK(clk), .RN(rstn), .Q(x7_75[21]) );
  DFFRHQX1 x7_75_reg_20_ ( .D(N667), .CK(clk), .RN(rstn), .Q(x7_75[20]) );
  DFFRHQX1 x4_tmp2_reg_22_ ( .D(N852), .CK(clk), .RN(rstn), .Q(x4_tmp2[22]) );
  DFFRHQX1 x4_tmp2_reg_21_ ( .D(N851), .CK(clk), .RN(rstn), .Q(x4_tmp2[21]) );
  DFFRHQX1 x5_tmp2_reg_22_ ( .D(N972), .CK(clk), .RN(rstn), .Q(x5_tmp2[22]) );
  DFFRHQX1 x5_tmp2_reg_21_ ( .D(N971), .CK(clk), .RN(rstn), .Q(x5_tmp2[21]) );
  DFFRHQX1 x6_tmp2_reg_22_ ( .D(N1115), .CK(clk), .RN(rstn), .Q(x6_tmp2[22])
         );
  DFFRHQX1 x6_tmp2_reg_21_ ( .D(N1114), .CK(clk), .RN(rstn), .Q(x6_tmp2[21])
         );
  DFFRHQX1 x7_tmp2_reg_22_ ( .D(N1188), .CK(clk), .RN(rstn), .Q(x7_tmp2[22])
         );
  DFFRHQX1 x7_tmp2_reg_21_ ( .D(N1187), .CK(clk), .RN(rstn), .Q(x7_tmp2[21])
         );
  DFFRHQX1 x7_89_tmp1_reg_0_ ( .D(x7[0]), .CK(clk), .RN(rstn), .Q(
        x7_89_tmp1[0]) );
  DFFRHQX1 x6_89_tmp1_reg_0_ ( .D(x6[0]), .CK(clk), .RN(rstn), .Q(
        x6_89_tmp1[0]) );
  DFFRHQX1 x5_89_tmp1_reg_0_ ( .D(x5[0]), .CK(clk), .RN(rstn), .Q(
        x5_89_tmp1[0]) );
  DFFRHQX1 x5_75_tmp1_reg_0_ ( .D(x5[0]), .CK(clk), .RN(rstn), .Q(
        x5_75_tmp1[0]) );
  DFFRHQX1 x4_75_tmp1_reg_0_ ( .D(x4[0]), .CK(clk), .RN(rstn), .Q(
        x4_75_tmp1[0]) );
  DFFRHQX1 x7_75_tmp1_reg_0_ ( .D(x7[0]), .CK(clk), .RN(rstn), .Q(
        x7_75_tmp1[0]) );
  DFFRHQX1 x6_75_tmp1_reg_0_ ( .D(x6[0]), .CK(clk), .RN(rstn), .Q(
        x6_75_tmp1[0]) );
  DFFRHQX1 x4_89_tmp1_reg_0_ ( .D(x4[0]), .CK(clk), .RN(rstn), .Q(
        x4_89_tmp1[0]) );
  DFFRHQX1 x4_89_reg_0_ ( .D(N357), .CK(clk), .RN(rstn), .Q(x4_89[0]) );
  DFFRHQX1 x4_50_reg_21_ ( .D(N424), .CK(clk), .RN(rstn), .Q(x4_50[21]) );
  DFFRHQX1 x7_tmp_reg_23_ ( .D(N1213), .CK(clk), .RN(rstn), .Q(x7_tmp[23]) );
  DFFRHQX1 x5_tmp_reg_23_ ( .D(N997), .CK(clk), .RN(rstn), .Q(x5_tmp[23]) );
  DFFRHQX1 x6_tmp_reg_23_ ( .D(N1140), .CK(clk), .RN(rstn), .Q(x6_tmp[23]) );
  DFFRHQX1 x4_tmp_reg_23_ ( .D(N877), .CK(clk), .RN(rstn), .Q(x4_tmp[23]) );
  DFFRHQX1 x4_50_tmp2_reg_20_ ( .D(N101), .CK(clk), .RN(rstn), .Q(
        x4_50_tmp2[20]) );
  DFFRHQX1 x6_50_tmp2_reg_20_ ( .D(N271), .CK(clk), .RN(rstn), .Q(
        x6_50_tmp2[20]) );
  DFFRHQX1 x5_50_tmp2_reg_20_ ( .D(N186), .CK(clk), .RN(rstn), .Q(
        x5_50_tmp2[20]) );
  DFFRHQX1 x7_50_tmp2_reg_20_ ( .D(N356), .CK(clk), .RN(rstn), .Q(
        x7_50_tmp2[20]) );
  DFFRHQX1 x6_89_reg_22_ ( .D(N557), .CK(clk), .RN(rstn), .Q(x6_89[22]) );
  DFFRHQX1 x7_75_reg_22_ ( .D(N669), .CK(clk), .RN(rstn), .Q(x7_75[22]) );
  DFFRHQX1 x4_tmp2_reg_23_ ( .D(N853), .CK(clk), .RN(rstn), .Q(x4_tmp2[23]) );
  DFFRHQX1 x5_tmp2_reg_23_ ( .D(N973), .CK(clk), .RN(rstn), .Q(x5_tmp2[23]) );
  DFFRHQX1 x6_tmp2_reg_23_ ( .D(N1116), .CK(clk), .RN(rstn), .Q(x6_tmp2[23])
         );
  DFFRHQX1 x7_tmp2_reg_23_ ( .D(N1189), .CK(clk), .RN(rstn), .Q(x7_tmp2[23])
         );
  DFFRHQX1 x7_tmp_reg_24_ ( .D(N1214), .CK(clk), .RN(rstn), .Q(x7_tmp[24]) );
  DFFRHQX1 x5_tmp_reg_24_ ( .D(N998), .CK(clk), .RN(rstn), .Q(x5_tmp[24]) );
  DFFRHQX1 x6_tmp_reg_24_ ( .D(N1141), .CK(clk), .RN(rstn), .Q(x6_tmp[24]) );
  DFFRHQX1 x4_tmp_reg_24_ ( .D(N878), .CK(clk), .RN(rstn), .Q(x4_tmp[24]) );
  DFFRHQX1 x6_89_tmp2_reg_20_ ( .D(N230), .CK(clk), .RN(rstn), .Q(
        x6_89_tmp2[20]) );
  DFFRHQX1 x5_89_tmp2_reg_20_ ( .D(N145), .CK(clk), .RN(rstn), .Q(
        x5_89_tmp2[20]) );
  DFFRHQX1 x4_89_tmp2_reg_20_ ( .D(N60), .CK(clk), .RN(rstn), .Q(
        x4_89_tmp2[20]) );
  DFFRHQX1 x7_89_tmp2_reg_20_ ( .D(N315), .CK(clk), .RN(rstn), .Q(
        x7_89_tmp2[20]) );
  DFFRHQX1 x6_50_reg_21_ ( .D(N602), .CK(clk), .RN(rstn), .Q(x6_50[21]) );
  DFFRHQX1 x7_89_tmp1_reg_18_ ( .D(N290), .CK(clk), .RN(rstn), .Q(
        x7_89_tmp1[18]) );
  DFFRHQX1 x7_89_tmp1_reg_17_ ( .D(N289), .CK(clk), .RN(rstn), .Q(
        x7_89_tmp1[17]) );
  DFFRHQX1 x7_89_tmp1_reg_16_ ( .D(N288), .CK(clk), .RN(rstn), .Q(
        x7_89_tmp1[16]) );
  DFFRHQX1 x7_89_tmp1_reg_15_ ( .D(N287), .CK(clk), .RN(rstn), .Q(
        x7_89_tmp1[15]) );
  DFFRHQX1 x6_89_tmp1_reg_18_ ( .D(N205), .CK(clk), .RN(rstn), .Q(
        x6_89_tmp1[18]) );
  DFFRHQX1 x6_89_tmp1_reg_17_ ( .D(N204), .CK(clk), .RN(rstn), .Q(
        x6_89_tmp1[17]) );
  DFFRHQX1 x6_89_tmp1_reg_16_ ( .D(N203), .CK(clk), .RN(rstn), .Q(
        x6_89_tmp1[16]) );
  DFFRHQX1 x6_89_tmp1_reg_15_ ( .D(N202), .CK(clk), .RN(rstn), .Q(
        x6_89_tmp1[15]) );
  DFFRHQX1 x5_89_tmp1_reg_18_ ( .D(N120), .CK(clk), .RN(rstn), .Q(
        x5_89_tmp1[18]) );
  DFFRHQX1 x5_89_tmp1_reg_17_ ( .D(N119), .CK(clk), .RN(rstn), .Q(
        x5_89_tmp1[17]) );
  DFFRHQX1 x5_89_tmp1_reg_16_ ( .D(N118), .CK(clk), .RN(rstn), .Q(
        x5_89_tmp1[16]) );
  DFFRHQX1 x5_89_tmp1_reg_15_ ( .D(N117), .CK(clk), .RN(rstn), .Q(
        x5_89_tmp1[15]) );
  DFFRHQX1 x5_75_tmp1_reg_18_ ( .D(N120), .CK(clk), .RN(rstn), .Q(
        x5_75_tmp1[18]) );
  DFFRHQX1 x5_75_tmp1_reg_17_ ( .D(N119), .CK(clk), .RN(rstn), .Q(
        x5_75_tmp1[17]) );
  DFFRHQX1 x5_75_tmp1_reg_16_ ( .D(N118), .CK(clk), .RN(rstn), .Q(
        x5_75_tmp1[16]) );
  DFFRHQX1 x5_75_tmp1_reg_15_ ( .D(N117), .CK(clk), .RN(rstn), .Q(
        x5_75_tmp1[15]) );
  DFFRHQX1 x4_75_tmp1_reg_18_ ( .D(N35), .CK(clk), .RN(rstn), .Q(
        x4_75_tmp1[18]) );
  DFFRHQX1 x4_75_tmp1_reg_17_ ( .D(N34), .CK(clk), .RN(rstn), .Q(
        x4_75_tmp1[17]) );
  DFFRHQX1 x4_75_tmp1_reg_16_ ( .D(N33), .CK(clk), .RN(rstn), .Q(
        x4_75_tmp1[16]) );
  DFFRHQX1 x4_75_tmp1_reg_15_ ( .D(N32), .CK(clk), .RN(rstn), .Q(
        x4_75_tmp1[15]) );
  DFFRHQX1 x7_75_tmp1_reg_18_ ( .D(N290), .CK(clk), .RN(rstn), .Q(
        x7_75_tmp1[18]) );
  DFFRHQX1 x7_75_tmp1_reg_17_ ( .D(N289), .CK(clk), .RN(rstn), .Q(
        x7_75_tmp1[17]) );
  DFFRHQX1 x7_75_tmp1_reg_16_ ( .D(N288), .CK(clk), .RN(rstn), .Q(
        x7_75_tmp1[16]) );
  DFFRHQX1 x7_75_tmp1_reg_15_ ( .D(N287), .CK(clk), .RN(rstn), .Q(
        x7_75_tmp1[15]) );
  DFFRHQX1 x6_75_tmp1_reg_18_ ( .D(N205), .CK(clk), .RN(rstn), .Q(
        x6_75_tmp1[18]) );
  DFFRHQX1 x6_75_tmp1_reg_17_ ( .D(N204), .CK(clk), .RN(rstn), .Q(
        x6_75_tmp1[17]) );
  DFFRHQX1 x6_75_tmp1_reg_16_ ( .D(N203), .CK(clk), .RN(rstn), .Q(
        x6_75_tmp1[16]) );
  DFFRHQX1 x6_75_tmp1_reg_15_ ( .D(N202), .CK(clk), .RN(rstn), .Q(
        x6_75_tmp1[15]) );
  DFFRHQX1 x4_50_tmp1_reg_17_ ( .D(n78), .CK(clk), .RN(rstn), .Q(
        x4_50_tmp1[17]) );
  DFFRHQX1 x4_50_tmp1_reg_16_ ( .D(n77), .CK(clk), .RN(rstn), .Q(
        x4_50_tmp1[16]) );
  DFFRHQX1 x4_50_tmp1_reg_15_ ( .D(n76), .CK(clk), .RN(rstn), .Q(
        x4_50_tmp1[15]) );
  DFFRHQX1 x4_50_tmp1_reg_14_ ( .D(n75), .CK(clk), .RN(rstn), .Q(
        x4_50_tmp1[14]) );
  DFFRHQX1 x6_50_tmp1_reg_17_ ( .D(n52), .CK(clk), .RN(rstn), .Q(
        x6_50_tmp1[17]) );
  DFFRHQX1 x6_50_tmp1_reg_16_ ( .D(n51), .CK(clk), .RN(rstn), .Q(
        x6_50_tmp1[16]) );
  DFFRHQX1 x6_50_tmp1_reg_15_ ( .D(n50), .CK(clk), .RN(rstn), .Q(
        x6_50_tmp1[15]) );
  DFFRHQX1 x6_50_tmp1_reg_14_ ( .D(n49), .CK(clk), .RN(rstn), .Q(
        x6_50_tmp1[14]) );
  DFFRHQX1 x5_50_tmp1_reg_17_ ( .D(n65), .CK(clk), .RN(rstn), .Q(
        x5_50_tmp1[17]) );
  DFFRHQX1 x5_50_tmp1_reg_16_ ( .D(n64), .CK(clk), .RN(rstn), .Q(
        x5_50_tmp1[16]) );
  DFFRHQX1 x5_50_tmp1_reg_15_ ( .D(n63), .CK(clk), .RN(rstn), .Q(
        x5_50_tmp1[15]) );
  DFFRHQX1 x5_50_tmp1_reg_14_ ( .D(n62), .CK(clk), .RN(rstn), .Q(
        x5_50_tmp1[14]) );
  DFFRHQX1 x7_50_tmp1_reg_17_ ( .D(n39), .CK(clk), .RN(rstn), .Q(
        x7_50_tmp1[17]) );
  DFFRHQX1 x7_50_tmp1_reg_16_ ( .D(n38), .CK(clk), .RN(rstn), .Q(
        x7_50_tmp1[16]) );
  DFFRHQX1 x7_50_tmp1_reg_15_ ( .D(n37), .CK(clk), .RN(rstn), .Q(
        x7_50_tmp1[15]) );
  DFFRHQX1 x7_50_tmp1_reg_14_ ( .D(n36), .CK(clk), .RN(rstn), .Q(
        x7_50_tmp1[14]) );
  DFFRHQX1 x4_18_tmp1_reg_16_ ( .D(n78), .CK(clk), .RN(rstn), .Q(
        x4_18_tmp1[16]) );
  DFFRHQX1 x4_18_tmp1_reg_15_ ( .D(n77), .CK(clk), .RN(rstn), .Q(
        x4_18_tmp1[15]) );
  DFFRHQX1 x4_18_tmp1_reg_14_ ( .D(n76), .CK(clk), .RN(rstn), .Q(
        x4_18_tmp1[14]) );
  DFFRHQX1 x4_18_tmp1_reg_13_ ( .D(n75), .CK(clk), .RN(rstn), .Q(
        x4_18_tmp1[13]) );
  DFFRHQX1 x5_18_tmp1_reg_16_ ( .D(n65), .CK(clk), .RN(rstn), .Q(
        x5_18_tmp1[16]) );
  DFFRHQX1 x5_18_tmp1_reg_15_ ( .D(n64), .CK(clk), .RN(rstn), .Q(
        x5_18_tmp1[15]) );
  DFFRHQX1 x5_18_tmp1_reg_14_ ( .D(n63), .CK(clk), .RN(rstn), .Q(
        x5_18_tmp1[14]) );
  DFFRHQX1 x5_18_tmp1_reg_13_ ( .D(n62), .CK(clk), .RN(rstn), .Q(
        x5_18_tmp1[13]) );
  DFFRHQX1 x6_18_tmp1_reg_16_ ( .D(n52), .CK(clk), .RN(rstn), .Q(
        x6_18_tmp1[16]) );
  DFFRHQX1 x6_18_tmp1_reg_15_ ( .D(n51), .CK(clk), .RN(rstn), .Q(
        x6_18_tmp1[15]) );
  DFFRHQX1 x6_18_tmp1_reg_14_ ( .D(n50), .CK(clk), .RN(rstn), .Q(
        x6_18_tmp1[14]) );
  DFFRHQX1 x6_18_tmp1_reg_13_ ( .D(n49), .CK(clk), .RN(rstn), .Q(
        x6_18_tmp1[13]) );
  DFFRHQX1 x7_18_tmp1_reg_16_ ( .D(n39), .CK(clk), .RN(rstn), .Q(
        x7_18_tmp1[16]) );
  DFFRHQX1 x7_18_tmp1_reg_15_ ( .D(n38), .CK(clk), .RN(rstn), .Q(
        x7_18_tmp1[15]) );
  DFFRHQX1 x7_18_tmp1_reg_14_ ( .D(n37), .CK(clk), .RN(rstn), .Q(
        x7_18_tmp1[14]) );
  DFFRHQX1 x7_18_tmp1_reg_13_ ( .D(n36), .CK(clk), .RN(rstn), .Q(
        x7_18_tmp1[13]) );
  DFFRHQX1 x5_18_reg_19_ ( .D(N533), .CK(clk), .RN(rstn), .Q(x5_18[19]) );
  DFFRHQX1 x5_18_reg_18_ ( .D(N532), .CK(clk), .RN(rstn), .Q(x5_18[18]) );
  DFFRHQX1 x5_18_reg_17_ ( .D(N531), .CK(clk), .RN(rstn), .Q(x5_18[17]) );
  DFFRHQX1 x6_18_reg_19_ ( .D(N622), .CK(clk), .RN(rstn), .Q(x6_18[19]) );
  DFFRHQX1 x6_18_reg_18_ ( .D(N621), .CK(clk), .RN(rstn), .Q(x6_18[18]) );
  DFFRHQX1 x6_18_reg_17_ ( .D(N620), .CK(clk), .RN(rstn), .Q(x6_18[17]) );
  DFFRHQX1 x6_18_reg_16_ ( .D(N619), .CK(clk), .RN(rstn), .Q(x6_18[16]) );
  DFFRHQX1 x4_18_reg_19_ ( .D(N444), .CK(clk), .RN(rstn), .Q(x4_18[19]) );
  DFFRHQX1 x4_18_reg_18_ ( .D(N443), .CK(clk), .RN(rstn), .Q(x4_18[18]) );
  DFFRHQX1 x4_18_reg_17_ ( .D(N442), .CK(clk), .RN(rstn), .Q(x4_18[17]) );
  DFFRHQX1 x4_18_reg_16_ ( .D(N441), .CK(clk), .RN(rstn), .Q(x4_18[16]) );
  DFFRHQX1 x4_89_tmp1_reg_18_ ( .D(N35), .CK(clk), .RN(rstn), .Q(
        x4_89_tmp1[18]) );
  DFFRHQX1 x4_89_tmp1_reg_17_ ( .D(N34), .CK(clk), .RN(rstn), .Q(
        x4_89_tmp1[17]) );
  DFFRHQX1 x4_89_tmp1_reg_16_ ( .D(N33), .CK(clk), .RN(rstn), .Q(
        x4_89_tmp1[16]) );
  DFFRHQX1 x4_89_tmp1_reg_15_ ( .D(N32), .CK(clk), .RN(rstn), .Q(
        x4_89_tmp1[15]) );
  DFFRHQX1 x4_89_reg_19_ ( .D(N376), .CK(clk), .RN(rstn), .Q(x4_89[19]) );
  DFFRHQX1 x4_89_reg_18_ ( .D(N375), .CK(clk), .RN(rstn), .Q(x4_89[18]) );
  DFFRHQX1 x4_89_reg_17_ ( .D(N374), .CK(clk), .RN(rstn), .Q(x4_89[17]) );
  DFFRHQX1 x4_89_reg_16_ ( .D(N373), .CK(clk), .RN(rstn), .Q(x4_89[16]) );
  DFFRHQX1 x4_75_reg_19_ ( .D(N399), .CK(clk), .RN(rstn), .Q(x4_75[19]) );
  DFFRHQX1 x4_75_reg_18_ ( .D(N398), .CK(clk), .RN(rstn), .Q(x4_75[18]) );
  DFFRHQX1 x4_75_reg_17_ ( .D(N397), .CK(clk), .RN(rstn), .Q(x4_75[17]) );
  DFFRHQX1 x4_75_reg_16_ ( .D(N396), .CK(clk), .RN(rstn), .Q(x4_75[16]) );
  DFFRHQX1 x5_75_reg_19_ ( .D(N488), .CK(clk), .RN(rstn), .Q(x5_75[19]) );
  DFFRHQX1 x5_75_reg_18_ ( .D(N487), .CK(clk), .RN(rstn), .Q(x5_75[18]) );
  DFFRHQX1 x5_75_reg_17_ ( .D(N486), .CK(clk), .RN(rstn), .Q(x5_75[17]) );
  DFFRHQX1 x5_75_reg_16_ ( .D(N485), .CK(clk), .RN(rstn), .Q(x5_75[16]) );
  DFFRHQX1 x6_75_reg_19_ ( .D(N577), .CK(clk), .RN(rstn), .Q(x6_75[19]) );
  DFFRHQX1 x6_75_reg_18_ ( .D(N576), .CK(clk), .RN(rstn), .Q(x6_75[18]) );
  DFFRHQX1 x6_75_reg_17_ ( .D(N575), .CK(clk), .RN(rstn), .Q(x6_75[17]) );
  DFFRHQX1 x6_75_reg_16_ ( .D(N574), .CK(clk), .RN(rstn), .Q(x6_75[16]) );
  DFFRHQX1 x4_50_reg_19_ ( .D(N422), .CK(clk), .RN(rstn), .Q(x4_50[19]) );
  DFFRHQX1 x4_50_reg_18_ ( .D(N421), .CK(clk), .RN(rstn), .Q(x4_50[18]) );
  DFFRHQX1 x4_50_reg_17_ ( .D(N420), .CK(clk), .RN(rstn), .Q(x4_50[17]) );
  DFFRHQX1 x4_50_reg_16_ ( .D(N419), .CK(clk), .RN(rstn), .Q(x4_50[16]) );
  DFFRHQX1 x5_tmp1_reg_20_ ( .D(N899), .CK(clk), .RN(rstn), .Q(x5_tmp1[20]) );
  DFFRHQX1 x5_tmp1_reg_19_ ( .D(N898), .CK(clk), .RN(rstn), .Q(x5_tmp1[19]) );
  DFFRHQX1 x5_tmp1_reg_18_ ( .D(N897), .CK(clk), .RN(rstn), .Q(x5_tmp1[18]) );
  DFFRHQX1 x5_tmp1_reg_17_ ( .D(N896), .CK(clk), .RN(rstn), .Q(x5_tmp1[17]) );
  DFFRHQX1 x6_tmp1_reg_20_ ( .D(N1065), .CK(clk), .RN(rstn), .Q(x6_tmp1[20])
         );
  DFFRHQX1 x6_tmp1_reg_19_ ( .D(N1064), .CK(clk), .RN(rstn), .Q(x6_tmp1[19])
         );
  DFFRHQX1 x6_tmp1_reg_18_ ( .D(N1063), .CK(clk), .RN(rstn), .Q(x6_tmp1[18])
         );
  DFFRHQX1 x6_tmp1_reg_17_ ( .D(N1062), .CK(clk), .RN(rstn), .Q(x6_tmp1[17])
         );
  DFFRHQX1 x7_tmp1_reg_20_ ( .D(N1162), .CK(clk), .RN(rstn), .Q(x7_tmp1[20])
         );
  DFFRHQX1 x7_tmp1_reg_19_ ( .D(N1161), .CK(clk), .RN(rstn), .Q(x7_tmp1[19])
         );
  DFFRHQX1 x7_tmp1_reg_18_ ( .D(N1160), .CK(clk), .RN(rstn), .Q(x7_tmp1[18])
         );
  DFFRHQX1 x7_tmp1_reg_17_ ( .D(N1159), .CK(clk), .RN(rstn), .Q(x7_tmp1[17])
         );
  DFFRHQX1 x4_tmp1_reg_20_ ( .D(N780), .CK(clk), .RN(rstn), .Q(x4_tmp1[20]) );
  DFFRHQX1 x4_tmp1_reg_19_ ( .D(N779), .CK(clk), .RN(rstn), .Q(x4_tmp1[19]) );
  DFFRHQX1 x4_tmp1_reg_18_ ( .D(N778), .CK(clk), .RN(rstn), .Q(x4_tmp1[18]) );
  DFFRHQX1 x4_tmp1_reg_17_ ( .D(N777), .CK(clk), .RN(rstn), .Q(x4_tmp1[17]) );
  DFFRHQX1 y6_tmp_reg_24_ ( .D(N1548), .CK(clk), .RN(rstn), .Q(y6_tmp[24]) );
  DFFRHQX1 y6_tmp_reg_23_ ( .D(N1547), .CK(clk), .RN(rstn), .Q(y6_tmp[23]) );
  DFFRHQX1 y6_tmp_reg_22_ ( .D(N1546), .CK(clk), .RN(rstn), .Q(y6_tmp[22]) );
  DFFRHQX1 y7_tmp_reg_24_ ( .D(N1625), .CK(clk), .RN(rstn), .Q(y7_tmp[24]) );
  DFFRHQX1 y7_tmp_reg_23_ ( .D(N1624), .CK(clk), .RN(rstn), .Q(y7_tmp[23]) );
  DFFRHQX1 y7_tmp_reg_22_ ( .D(N1623), .CK(clk), .RN(rstn), .Q(y7_tmp[22]) );
  DFFRHQX1 y0_tmp_reg_24_ ( .D(N1239), .CK(clk), .RN(rstn), .Q(y0_tmp[24]) );
  DFFRHQX1 y1_tmp_reg_24_ ( .D(N1265), .CK(clk), .RN(rstn), .Q(y1_tmp[24]) );
  DFFRHQX1 y2_tmp_reg_24_ ( .D(N1291), .CK(clk), .RN(rstn), .Q(y2_tmp[24]) );
  DFFRHQX1 y3_tmp_reg_24_ ( .D(N1317), .CK(clk), .RN(rstn), .Q(y3_tmp[24]) );
  DFFRHQX1 y4_tmp_reg_24_ ( .D(N1394), .CK(clk), .RN(rstn), .Q(y4_tmp[24]) );
  DFFRHQX1 y4_tmp_reg_23_ ( .D(N1393), .CK(clk), .RN(rstn), .Q(y4_tmp[23]) );
  DFFRHQX1 y4_tmp_reg_22_ ( .D(N1392), .CK(clk), .RN(rstn), .Q(y4_tmp[22]) );
  DFFRHQX1 y5_tmp_reg_24_ ( .D(N1471), .CK(clk), .RN(rstn), .Q(y5_tmp[24]) );
  DFFRHQX1 y5_tmp_reg_23_ ( .D(N1470), .CK(clk), .RN(rstn), .Q(y5_tmp[23]) );
  DFFRHQX1 y5_tmp_reg_22_ ( .D(N1469), .CK(clk), .RN(rstn), .Q(y5_tmp[22]) );
  DFFRHQX1 x7_50_reg_19_ ( .D(N689), .CK(clk), .RN(rstn), .Q(x7_50[19]) );
  DFFRHQX1 x7_50_reg_18_ ( .D(N688), .CK(clk), .RN(rstn), .Q(x7_50[18]) );
  DFFRHQX1 x7_50_reg_17_ ( .D(N687), .CK(clk), .RN(rstn), .Q(x7_50[17]) );
  DFFRHQX1 x7_50_reg_16_ ( .D(N686), .CK(clk), .RN(rstn), .Q(x7_50[16]) );
  DFFRHQX1 x5_89_reg_19_ ( .D(N465), .CK(clk), .RN(rstn), .Q(x5_89[19]) );
  DFFRHQX1 x5_89_reg_18_ ( .D(N464), .CK(clk), .RN(rstn), .Q(x5_89[18]) );
  DFFRHQX1 x5_89_reg_17_ ( .D(N463), .CK(clk), .RN(rstn), .Q(x5_89[17]) );
  DFFRHQX1 x5_89_reg_16_ ( .D(N462), .CK(clk), .RN(rstn), .Q(x5_89[16]) );
  DFFRHQX1 x7_89_reg_19_ ( .D(N643), .CK(clk), .RN(rstn), .Q(x7_89[19]) );
  DFFRHQX1 x7_89_reg_18_ ( .D(N642), .CK(clk), .RN(rstn), .Q(x7_89[18]) );
  DFFRHQX1 x7_89_reg_17_ ( .D(N641), .CK(clk), .RN(rstn), .Q(x7_89[17]) );
  DFFRHQX1 x7_89_reg_16_ ( .D(N640), .CK(clk), .RN(rstn), .Q(x7_89[16]) );
  DFFRHQX1 x5_50_reg_19_ ( .D(N511), .CK(clk), .RN(rstn), .Q(x5_50[19]) );
  DFFRHQX1 x5_50_reg_18_ ( .D(N510), .CK(clk), .RN(rstn), .Q(x5_50[18]) );
  DFFRHQX1 x5_50_reg_17_ ( .D(N509), .CK(clk), .RN(rstn), .Q(x5_50[17]) );
  DFFRHQX1 x5_50_reg_16_ ( .D(N508), .CK(clk), .RN(rstn), .Q(x5_50[16]) );
  DFFRHQX1 x6_89_tmp2_reg_18_ ( .D(N228), .CK(clk), .RN(rstn), .Q(
        x6_89_tmp2[18]) );
  DFFRHQX1 x6_89_tmp2_reg_17_ ( .D(N227), .CK(clk), .RN(rstn), .Q(
        x6_89_tmp2[17]) );
  DFFRHQX1 x6_89_tmp2_reg_16_ ( .D(N226), .CK(clk), .RN(rstn), .Q(
        x6_89_tmp2[16]) );
  DFFRHQX1 x6_89_tmp2_reg_15_ ( .D(N225), .CK(clk), .RN(rstn), .Q(
        x6_89_tmp2[15]) );
  DFFRHQX1 x6_89_tmp2_reg_14_ ( .D(N224), .CK(clk), .RN(rstn), .Q(
        x6_89_tmp2[14]) );
  DFFRHQX1 x5_89_tmp2_reg_18_ ( .D(N143), .CK(clk), .RN(rstn), .Q(
        x5_89_tmp2[18]) );
  DFFRHQX1 x5_89_tmp2_reg_17_ ( .D(N142), .CK(clk), .RN(rstn), .Q(
        x5_89_tmp2[17]) );
  DFFRHQX1 x5_89_tmp2_reg_16_ ( .D(N141), .CK(clk), .RN(rstn), .Q(
        x5_89_tmp2[16]) );
  DFFRHQX1 x5_89_tmp2_reg_15_ ( .D(N140), .CK(clk), .RN(rstn), .Q(
        x5_89_tmp2[15]) );
  DFFRHQX1 x5_89_tmp2_reg_14_ ( .D(N139), .CK(clk), .RN(rstn), .Q(
        x5_89_tmp2[14]) );
  DFFRHQX1 x4_89_tmp2_reg_18_ ( .D(N58), .CK(clk), .RN(rstn), .Q(
        x4_89_tmp2[18]) );
  DFFRHQX1 x4_89_tmp2_reg_17_ ( .D(N57), .CK(clk), .RN(rstn), .Q(
        x4_89_tmp2[17]) );
  DFFRHQX1 x4_89_tmp2_reg_16_ ( .D(N56), .CK(clk), .RN(rstn), .Q(
        x4_89_tmp2[16]) );
  DFFRHQX1 x4_89_tmp2_reg_15_ ( .D(N55), .CK(clk), .RN(rstn), .Q(
        x4_89_tmp2[15]) );
  DFFRHQX1 x4_89_tmp2_reg_14_ ( .D(N54), .CK(clk), .RN(rstn), .Q(
        x4_89_tmp2[14]) );
  DFFRHQX1 x7_89_tmp2_reg_18_ ( .D(N313), .CK(clk), .RN(rstn), .Q(
        x7_89_tmp2[18]) );
  DFFRHQX1 x7_89_tmp2_reg_17_ ( .D(N312), .CK(clk), .RN(rstn), .Q(
        x7_89_tmp2[17]) );
  DFFRHQX1 x7_89_tmp2_reg_16_ ( .D(N311), .CK(clk), .RN(rstn), .Q(
        x7_89_tmp2[16]) );
  DFFRHQX1 x7_89_tmp2_reg_15_ ( .D(N310), .CK(clk), .RN(rstn), .Q(
        x7_89_tmp2[15]) );
  DFFRHQX1 x7_89_tmp2_reg_14_ ( .D(N309), .CK(clk), .RN(rstn), .Q(
        x7_89_tmp2[14]) );
  DFFRHQX1 x4_75_tmp2_reg_18_ ( .D(N79), .CK(clk), .RN(rstn), .Q(
        x4_75_tmp2[18]) );
  DFFRHQX1 x4_75_tmp2_reg_17_ ( .D(N78), .CK(clk), .RN(rstn), .Q(
        x4_75_tmp2[17]) );
  DFFRHQX1 x4_75_tmp2_reg_16_ ( .D(N77), .CK(clk), .RN(rstn), .Q(
        x4_75_tmp2[16]) );
  DFFRHQX1 x4_75_tmp2_reg_15_ ( .D(N76), .CK(clk), .RN(rstn), .Q(
        x4_75_tmp2[15]) );
  DFFRHQX1 x4_75_tmp2_reg_14_ ( .D(N75), .CK(clk), .RN(rstn), .Q(
        x4_75_tmp2[14]) );
  DFFRHQX1 x5_75_tmp2_reg_18_ ( .D(N164), .CK(clk), .RN(rstn), .Q(
        x5_75_tmp2[18]) );
  DFFRHQX1 x5_75_tmp2_reg_17_ ( .D(N163), .CK(clk), .RN(rstn), .Q(
        x5_75_tmp2[17]) );
  DFFRHQX1 x5_75_tmp2_reg_16_ ( .D(N162), .CK(clk), .RN(rstn), .Q(
        x5_75_tmp2[16]) );
  DFFRHQX1 x5_75_tmp2_reg_15_ ( .D(N161), .CK(clk), .RN(rstn), .Q(
        x5_75_tmp2[15]) );
  DFFRHQX1 x5_75_tmp2_reg_14_ ( .D(N160), .CK(clk), .RN(rstn), .Q(
        x5_75_tmp2[14]) );
  DFFRHQX1 x6_75_tmp2_reg_18_ ( .D(N249), .CK(clk), .RN(rstn), .Q(
        x6_75_tmp2[18]) );
  DFFRHQX1 x6_75_tmp2_reg_17_ ( .D(N248), .CK(clk), .RN(rstn), .Q(
        x6_75_tmp2[17]) );
  DFFRHQX1 x6_75_tmp2_reg_16_ ( .D(N247), .CK(clk), .RN(rstn), .Q(
        x6_75_tmp2[16]) );
  DFFRHQX1 x6_75_tmp2_reg_15_ ( .D(N246), .CK(clk), .RN(rstn), .Q(
        x6_75_tmp2[15]) );
  DFFRHQX1 x6_75_tmp2_reg_14_ ( .D(N245), .CK(clk), .RN(rstn), .Q(
        x6_75_tmp2[14]) );
  DFFRHQX1 x7_75_tmp2_reg_18_ ( .D(N334), .CK(clk), .RN(rstn), .Q(
        x7_75_tmp2[18]) );
  DFFRHQX1 x7_75_tmp2_reg_17_ ( .D(N333), .CK(clk), .RN(rstn), .Q(
        x7_75_tmp2[17]) );
  DFFRHQX1 x7_75_tmp2_reg_16_ ( .D(N332), .CK(clk), .RN(rstn), .Q(
        x7_75_tmp2[16]) );
  DFFRHQX1 x7_75_tmp2_reg_15_ ( .D(N331), .CK(clk), .RN(rstn), .Q(
        x7_75_tmp2[15]) );
  DFFRHQX1 x7_75_tmp2_reg_14_ ( .D(N330), .CK(clk), .RN(rstn), .Q(
        x7_75_tmp2[14]) );
  DFFRHQX1 x4_50_tmp2_reg_17_ ( .D(N98), .CK(clk), .RN(rstn), .Q(
        x4_50_tmp2[17]) );
  DFFRHQX1 x4_50_tmp2_reg_16_ ( .D(N97), .CK(clk), .RN(rstn), .Q(
        x4_50_tmp2[16]) );
  DFFRHQX1 x4_50_tmp2_reg_15_ ( .D(N96), .CK(clk), .RN(rstn), .Q(
        x4_50_tmp2[15]) );
  DFFRHQX1 x4_50_tmp2_reg_14_ ( .D(N95), .CK(clk), .RN(rstn), .Q(
        x4_50_tmp2[14]) );
  DFFRHQX1 x4_50_tmp2_reg_13_ ( .D(N94), .CK(clk), .RN(rstn), .Q(
        x4_50_tmp2[13]) );
  DFFRHQX1 x6_50_tmp2_reg_17_ ( .D(N268), .CK(clk), .RN(rstn), .Q(
        x6_50_tmp2[17]) );
  DFFRHQX1 x6_50_tmp2_reg_16_ ( .D(N267), .CK(clk), .RN(rstn), .Q(
        x6_50_tmp2[16]) );
  DFFRHQX1 x6_50_tmp2_reg_15_ ( .D(N266), .CK(clk), .RN(rstn), .Q(
        x6_50_tmp2[15]) );
  DFFRHQX1 x6_50_tmp2_reg_14_ ( .D(N265), .CK(clk), .RN(rstn), .Q(
        x6_50_tmp2[14]) );
  DFFRHQX1 x6_50_tmp2_reg_13_ ( .D(N264), .CK(clk), .RN(rstn), .Q(
        x6_50_tmp2[13]) );
  DFFRHQX1 x6_50_reg_15_ ( .D(N596), .CK(clk), .RN(rstn), .Q(x6_50[15]) );
  DFFRHQX1 x6_50_reg_16_ ( .D(N597), .CK(clk), .RN(rstn), .Q(x6_50[16]) );
  DFFRHQX1 x6_50_reg_17_ ( .D(N598), .CK(clk), .RN(rstn), .Q(x6_50[17]) );
  DFFRHQX1 x6_50_reg_18_ ( .D(N599), .CK(clk), .RN(rstn), .Q(x6_50[18]) );
  DFFRHQX1 x6_50_reg_19_ ( .D(N600), .CK(clk), .RN(rstn), .Q(x6_50[19]) );
  DFFRHQX1 x5_50_tmp2_reg_17_ ( .D(N183), .CK(clk), .RN(rstn), .Q(
        x5_50_tmp2[17]) );
  DFFRHQX1 x5_50_tmp2_reg_16_ ( .D(N182), .CK(clk), .RN(rstn), .Q(
        x5_50_tmp2[16]) );
  DFFRHQX1 x5_50_tmp2_reg_15_ ( .D(N181), .CK(clk), .RN(rstn), .Q(
        x5_50_tmp2[15]) );
  DFFRHQX1 x5_50_tmp2_reg_14_ ( .D(N180), .CK(clk), .RN(rstn), .Q(
        x5_50_tmp2[14]) );
  DFFRHQX1 x5_50_tmp2_reg_13_ ( .D(N179), .CK(clk), .RN(rstn), .Q(
        x5_50_tmp2[13]) );
  DFFRHQX1 x7_50_tmp2_reg_17_ ( .D(N353), .CK(clk), .RN(rstn), .Q(
        x7_50_tmp2[17]) );
  DFFRHQX1 x7_50_tmp2_reg_16_ ( .D(N352), .CK(clk), .RN(rstn), .Q(
        x7_50_tmp2[16]) );
  DFFRHQX1 x7_50_tmp2_reg_15_ ( .D(N351), .CK(clk), .RN(rstn), .Q(
        x7_50_tmp2[15]) );
  DFFRHQX1 x7_50_tmp2_reg_14_ ( .D(N350), .CK(clk), .RN(rstn), .Q(
        x7_50_tmp2[14]) );
  DFFRHQX1 x7_50_tmp2_reg_13_ ( .D(N349), .CK(clk), .RN(rstn), .Q(
        x7_50_tmp2[13]) );
  DFFRHQX1 x4_18_tmp2_reg_15_ ( .D(n80), .CK(clk), .RN(rstn), .Q(
        x4_18_tmp2[15]) );
  DFFRHQX1 x4_18_tmp2_reg_14_ ( .D(n79), .CK(clk), .RN(rstn), .Q(
        x4_18_tmp2[14]) );
  DFFRHQX1 x4_18_tmp2_reg_13_ ( .D(n78), .CK(clk), .RN(rstn), .Q(
        x4_18_tmp2[13]) );
  DFFRHQX1 x4_18_tmp2_reg_12_ ( .D(n77), .CK(clk), .RN(rstn), .Q(
        x4_18_tmp2[12]) );
  DFFRHQX1 x6_18_tmp2_reg_15_ ( .D(n54), .CK(clk), .RN(rstn), .Q(
        x6_18_tmp2[15]) );
  DFFRHQX1 x6_18_tmp2_reg_14_ ( .D(n53), .CK(clk), .RN(rstn), .Q(
        x6_18_tmp2[14]) );
  DFFRHQX1 x6_18_tmp2_reg_13_ ( .D(n52), .CK(clk), .RN(rstn), .Q(
        x6_18_tmp2[13]) );
  DFFRHQX1 x6_18_tmp2_reg_12_ ( .D(n51), .CK(clk), .RN(rstn), .Q(
        x6_18_tmp2[12]) );
  DFFRHQX1 x5_18_tmp2_reg_15_ ( .D(n67), .CK(clk), .RN(rstn), .Q(
        x5_18_tmp2[15]) );
  DFFRHQX1 x5_18_tmp2_reg_14_ ( .D(n66), .CK(clk), .RN(rstn), .Q(
        x5_18_tmp2[14]) );
  DFFRHQX1 x5_18_tmp2_reg_13_ ( .D(n65), .CK(clk), .RN(rstn), .Q(
        x5_18_tmp2[13]) );
  DFFRHQX1 x5_18_tmp2_reg_12_ ( .D(n64), .CK(clk), .RN(rstn), .Q(
        x5_18_tmp2[12]) );
  DFFRHQX1 x7_18_tmp2_reg_15_ ( .D(n41), .CK(clk), .RN(rstn), .Q(
        x7_18_tmp2[15]) );
  DFFRHQX1 x7_18_tmp2_reg_14_ ( .D(n40), .CK(clk), .RN(rstn), .Q(
        x7_18_tmp2[14]) );
  DFFRHQX1 x7_18_tmp2_reg_13_ ( .D(n39), .CK(clk), .RN(rstn), .Q(
        x7_18_tmp2[13]) );
  DFFRHQX1 x7_18_tmp2_reg_12_ ( .D(n38), .CK(clk), .RN(rstn), .Q(
        x7_18_tmp2[12]) );
  DFFRHQX1 x7_18_reg_19_ ( .D(N711), .CK(clk), .RN(rstn), .Q(x7_18[19]) );
  DFFRHQX1 x7_18_reg_18_ ( .D(N710), .CK(clk), .RN(rstn), .Q(x7_18[18]) );
  DFFRHQX1 x7_18_reg_17_ ( .D(N709), .CK(clk), .RN(rstn), .Q(x7_18[17]) );
  DFFRHQX1 x7_18_reg_16_ ( .D(N708), .CK(clk), .RN(rstn), .Q(x7_18[16]) );
  DFFRHQX1 x7_18_reg_15_ ( .D(N707), .CK(clk), .RN(rstn), .Q(x7_18[15]) );
  DFFRHQX1 x6_89_reg_20_ ( .D(N555), .CK(clk), .RN(rstn), .Q(x6_89[20]) );
  DFFRHQX1 x6_89_reg_19_ ( .D(N554), .CK(clk), .RN(rstn), .Q(x6_89[19]) );
  DFFRHQX1 x6_89_reg_18_ ( .D(N553), .CK(clk), .RN(rstn), .Q(x6_89[18]) );
  DFFRHQX1 x6_89_reg_17_ ( .D(N552), .CK(clk), .RN(rstn), .Q(x6_89[17]) );
  DFFRHQX1 x7_75_reg_19_ ( .D(N666), .CK(clk), .RN(rstn), .Q(x7_75[19]) );
  DFFRHQX1 x7_75_reg_18_ ( .D(N665), .CK(clk), .RN(rstn), .Q(x7_75[18]) );
  DFFRHQX1 x7_75_reg_17_ ( .D(N664), .CK(clk), .RN(rstn), .Q(x7_75[17]) );
  DFFRHQX1 x7_75_reg_16_ ( .D(N663), .CK(clk), .RN(rstn), .Q(x7_75[16]) );
  DFFRHQX1 x7_75_reg_15_ ( .D(N662), .CK(clk), .RN(rstn), .Q(x7_75[15]) );
  DFFRHQX1 x4_tmp2_reg_20_ ( .D(N850), .CK(clk), .RN(rstn), .Q(x4_tmp2[20]) );
  DFFRHQX1 x4_tmp2_reg_19_ ( .D(N849), .CK(clk), .RN(rstn), .Q(x4_tmp2[19]) );
  DFFRHQX1 x4_tmp2_reg_18_ ( .D(N848), .CK(clk), .RN(rstn), .Q(x4_tmp2[18]) );
  DFFRHQX1 x4_tmp2_reg_17_ ( .D(N847), .CK(clk), .RN(rstn), .Q(x4_tmp2[17]) );
  DFFRHQX1 x4_tmp2_reg_16_ ( .D(N846), .CK(clk), .RN(rstn), .Q(x4_tmp2[16]) );
  DFFRHQX1 x5_tmp2_reg_20_ ( .D(N970), .CK(clk), .RN(rstn), .Q(x5_tmp2[20]) );
  DFFRHQX1 x5_tmp2_reg_19_ ( .D(N969), .CK(clk), .RN(rstn), .Q(x5_tmp2[19]) );
  DFFRHQX1 x5_tmp2_reg_18_ ( .D(N968), .CK(clk), .RN(rstn), .Q(x5_tmp2[18]) );
  DFFRHQX1 x5_tmp2_reg_17_ ( .D(N967), .CK(clk), .RN(rstn), .Q(x5_tmp2[17]) );
  DFFRHQX1 x5_tmp2_reg_16_ ( .D(N966), .CK(clk), .RN(rstn), .Q(x5_tmp2[16]) );
  DFFRHQX1 x6_tmp2_reg_20_ ( .D(N1113), .CK(clk), .RN(rstn), .Q(x6_tmp2[20])
         );
  DFFRHQX1 x6_tmp2_reg_19_ ( .D(N1112), .CK(clk), .RN(rstn), .Q(x6_tmp2[19])
         );
  DFFRHQX1 x6_tmp2_reg_18_ ( .D(N1111), .CK(clk), .RN(rstn), .Q(x6_tmp2[18])
         );
  DFFRHQX1 x6_tmp2_reg_17_ ( .D(N1110), .CK(clk), .RN(rstn), .Q(x6_tmp2[17])
         );
  DFFRHQX1 x6_tmp2_reg_16_ ( .D(N1109), .CK(clk), .RN(rstn), .Q(x6_tmp2[16])
         );
  DFFRHQX1 x7_tmp2_reg_20_ ( .D(N1186), .CK(clk), .RN(rstn), .Q(x7_tmp2[20])
         );
  DFFRHQX1 x7_tmp2_reg_19_ ( .D(N1185), .CK(clk), .RN(rstn), .Q(x7_tmp2[19])
         );
  DFFRHQX1 x7_tmp2_reg_18_ ( .D(N1184), .CK(clk), .RN(rstn), .Q(x7_tmp2[18])
         );
  DFFRHQX1 x7_tmp2_reg_17_ ( .D(N1183), .CK(clk), .RN(rstn), .Q(x7_tmp2[17])
         );
  DFFRHQX1 x7_tmp2_reg_16_ ( .D(N1182), .CK(clk), .RN(rstn), .Q(x7_tmp2[16])
         );
  DFFRHQX1 y6_tmp_reg_25_ ( .D(N1549), .CK(clk), .RN(rstn), .Q(y6_tmp[25]) );
  DFFRHQX1 y7_tmp_reg_25_ ( .D(N1626), .CK(clk), .RN(rstn), .Q(y7_tmp[25]) );
  DFFRHQX1 y0_tmp_reg_25_ ( .D(N1240), .CK(clk), .RN(rstn), .Q(y0_tmp[25]) );
  DFFRHQX1 y1_tmp_reg_25_ ( .D(N1266), .CK(clk), .RN(rstn), .Q(y1_tmp[25]) );
  DFFRHQX1 y2_tmp_reg_25_ ( .D(N1292), .CK(clk), .RN(rstn), .Q(y2_tmp[25]) );
  DFFRHQX1 y3_tmp_reg_25_ ( .D(N1318), .CK(clk), .RN(rstn), .Q(y3_tmp[25]) );
  DFFRHQX1 y4_tmp_reg_25_ ( .D(N1395), .CK(clk), .RN(rstn), .Q(y4_tmp[25]) );
  DFFRHQX1 y5_tmp_reg_25_ ( .D(N1472), .CK(clk), .RN(rstn), .Q(y5_tmp[25]) );
  DFFRHQX1 x5_18_reg_20_ ( .D(N534), .CK(clk), .RN(rstn), .Q(x5_18[20]) );
  DFFRHQX1 x6_18_reg_20_ ( .D(N623), .CK(clk), .RN(rstn), .Q(x6_18[20]) );
  DFFRHQX1 x4_18_reg_20_ ( .D(N445), .CK(clk), .RN(rstn), .Q(x4_18[20]) );
  DFFRHQX1 x7_tmp_reg_18_ ( .D(N1208), .CK(clk), .RN(rstn), .Q(x7_tmp[18]) );
  DFFRHQX1 x7_tmp_reg_19_ ( .D(N1209), .CK(clk), .RN(rstn), .Q(x7_tmp[19]) );
  DFFRHQX1 x7_tmp_reg_20_ ( .D(N1210), .CK(clk), .RN(rstn), .Q(x7_tmp[20]) );
  DFFRHQX1 x7_tmp_reg_21_ ( .D(N1211), .CK(clk), .RN(rstn), .Q(x7_tmp[21]) );
  DFFRHQX1 x7_tmp_reg_22_ ( .D(N1212), .CK(clk), .RN(rstn), .Q(x7_tmp[22]) );
  DFFRHQX1 x5_tmp_reg_22_ ( .D(N996), .CK(clk), .RN(rstn), .Q(x5_tmp[22]) );
  DFFRHQX1 x5_tmp_reg_21_ ( .D(N995), .CK(clk), .RN(rstn), .Q(x5_tmp[21]) );
  DFFRHQX1 x5_tmp_reg_20_ ( .D(N994), .CK(clk), .RN(rstn), .Q(x5_tmp[20]) );
  DFFRHQX1 x5_tmp_reg_19_ ( .D(N993), .CK(clk), .RN(rstn), .Q(x5_tmp[19]) );
  DFFRHQX1 x5_tmp_reg_18_ ( .D(N992), .CK(clk), .RN(rstn), .Q(x5_tmp[18]) );
  DFFRHQX1 x6_tmp_reg_22_ ( .D(N1139), .CK(clk), .RN(rstn), .Q(x6_tmp[22]) );
  DFFRHQX1 x6_tmp_reg_21_ ( .D(N1138), .CK(clk), .RN(rstn), .Q(x6_tmp[21]) );
  DFFRHQX1 x6_tmp_reg_20_ ( .D(N1137), .CK(clk), .RN(rstn), .Q(x6_tmp[20]) );
  DFFRHQX1 x6_tmp_reg_19_ ( .D(N1136), .CK(clk), .RN(rstn), .Q(x6_tmp[19]) );
  DFFRHQX1 x6_tmp_reg_18_ ( .D(N1135), .CK(clk), .RN(rstn), .Q(x6_tmp[18]) );
  DFFRHQX1 x4_tmp_reg_18_ ( .D(N872), .CK(clk), .RN(rstn), .Q(x4_tmp[18]) );
  DFFRHQX1 x4_tmp_reg_19_ ( .D(N873), .CK(clk), .RN(rstn), .Q(x4_tmp[19]) );
  DFFRHQX1 x4_tmp_reg_20_ ( .D(N874), .CK(clk), .RN(rstn), .Q(x4_tmp[20]) );
  DFFRHQX1 x4_tmp_reg_21_ ( .D(N875), .CK(clk), .RN(rstn), .Q(x4_tmp[21]) );
  DFFRHQX1 x4_tmp_reg_22_ ( .D(N876), .CK(clk), .RN(rstn), .Q(x4_tmp[22]) );
  DFFRHQX1 x4_75_tmp2_reg_19_ ( .D(N80), .CK(clk), .RN(rstn), .Q(
        x4_75_tmp2[19]) );
  DFFRHQX1 x5_75_tmp2_reg_19_ ( .D(N165), .CK(clk), .RN(rstn), .Q(
        x5_75_tmp2[19]) );
  DFFRHQX1 x6_75_tmp2_reg_19_ ( .D(N250), .CK(clk), .RN(rstn), .Q(
        x6_75_tmp2[19]) );
  DFFRHQX1 x7_75_tmp2_reg_19_ ( .D(N335), .CK(clk), .RN(rstn), .Q(
        x7_75_tmp2[19]) );
  DFFRHQX1 x7_18_reg_20_ ( .D(N712), .CK(clk), .RN(rstn), .Q(x7_18[20]) );
  DFFRHQX1 x4_18_tmp2_reg_16_ ( .D(x4[15]), .CK(clk), .RN(rstn), .Q(
        x4_18_tmp2[16]) );
  DFFRHQX1 x6_18_tmp2_reg_16_ ( .D(x6[15]), .CK(clk), .RN(rstn), .Q(
        x6_18_tmp2[16]) );
  DFFRHQX1 x5_18_tmp2_reg_16_ ( .D(x5[15]), .CK(clk), .RN(rstn), .Q(
        x5_18_tmp2[16]) );
  DFFRHQX1 x7_18_tmp2_reg_16_ ( .D(x7[15]), .CK(clk), .RN(rstn), .Q(
        x7_18_tmp2[16]) );
  DFFRHQX1 mode_delay2_reg_1_ ( .D(mode_delay1[1]), .CK(clk), .RN(rstn), .Q(
        mode_delay2[1]) );
  DFFRHQX1 x7_89_tmp1_reg_14_ ( .D(N286), .CK(clk), .RN(rstn), .Q(
        x7_89_tmp1[14]) );
  DFFRHQX1 x7_89_tmp1_reg_13_ ( .D(N285), .CK(clk), .RN(rstn), .Q(
        x7_89_tmp1[13]) );
  DFFRHQX1 x7_89_tmp1_reg_12_ ( .D(N284), .CK(clk), .RN(rstn), .Q(
        x7_89_tmp1[12]) );
  DFFRHQX1 x7_89_tmp1_reg_11_ ( .D(N283), .CK(clk), .RN(rstn), .Q(
        x7_89_tmp1[11]) );
  DFFRHQX1 x7_89_tmp1_reg_10_ ( .D(N282), .CK(clk), .RN(rstn), .Q(
        x7_89_tmp1[10]) );
  DFFRHQX1 x6_89_tmp1_reg_14_ ( .D(N201), .CK(clk), .RN(rstn), .Q(
        x6_89_tmp1[14]) );
  DFFRHQX1 x6_89_tmp1_reg_13_ ( .D(N200), .CK(clk), .RN(rstn), .Q(
        x6_89_tmp1[13]) );
  DFFRHQX1 x6_89_tmp1_reg_12_ ( .D(N199), .CK(clk), .RN(rstn), .Q(
        x6_89_tmp1[12]) );
  DFFRHQX1 x6_89_tmp1_reg_11_ ( .D(N198), .CK(clk), .RN(rstn), .Q(
        x6_89_tmp1[11]) );
  DFFRHQX1 x6_89_tmp1_reg_10_ ( .D(N197), .CK(clk), .RN(rstn), .Q(
        x6_89_tmp1[10]) );
  DFFRHQX1 x5_89_tmp1_reg_14_ ( .D(N116), .CK(clk), .RN(rstn), .Q(
        x5_89_tmp1[14]) );
  DFFRHQX1 x5_89_tmp1_reg_13_ ( .D(N115), .CK(clk), .RN(rstn), .Q(
        x5_89_tmp1[13]) );
  DFFRHQX1 x5_89_tmp1_reg_12_ ( .D(N114), .CK(clk), .RN(rstn), .Q(
        x5_89_tmp1[12]) );
  DFFRHQX1 x5_89_tmp1_reg_11_ ( .D(N113), .CK(clk), .RN(rstn), .Q(
        x5_89_tmp1[11]) );
  DFFRHQX1 x5_89_tmp1_reg_10_ ( .D(N112), .CK(clk), .RN(rstn), .Q(
        x5_89_tmp1[10]) );
  DFFRHQX1 x5_75_tmp1_reg_14_ ( .D(N116), .CK(clk), .RN(rstn), .Q(
        x5_75_tmp1[14]) );
  DFFRHQX1 x5_75_tmp1_reg_13_ ( .D(N115), .CK(clk), .RN(rstn), .Q(
        x5_75_tmp1[13]) );
  DFFRHQX1 x5_75_tmp1_reg_12_ ( .D(N114), .CK(clk), .RN(rstn), .Q(
        x5_75_tmp1[12]) );
  DFFRHQX1 x5_75_tmp1_reg_11_ ( .D(N113), .CK(clk), .RN(rstn), .Q(
        x5_75_tmp1[11]) );
  DFFRHQX1 x5_75_tmp1_reg_10_ ( .D(N112), .CK(clk), .RN(rstn), .Q(
        x5_75_tmp1[10]) );
  DFFRHQX1 x4_75_tmp1_reg_14_ ( .D(N31), .CK(clk), .RN(rstn), .Q(
        x4_75_tmp1[14]) );
  DFFRHQX1 x4_75_tmp1_reg_13_ ( .D(N30), .CK(clk), .RN(rstn), .Q(
        x4_75_tmp1[13]) );
  DFFRHQX1 x4_75_tmp1_reg_12_ ( .D(N29), .CK(clk), .RN(rstn), .Q(
        x4_75_tmp1[12]) );
  DFFRHQX1 x4_75_tmp1_reg_11_ ( .D(N28), .CK(clk), .RN(rstn), .Q(
        x4_75_tmp1[11]) );
  DFFRHQX1 x4_75_tmp1_reg_10_ ( .D(N27), .CK(clk), .RN(rstn), .Q(
        x4_75_tmp1[10]) );
  DFFRHQX1 x7_75_tmp1_reg_14_ ( .D(N286), .CK(clk), .RN(rstn), .Q(
        x7_75_tmp1[14]) );
  DFFRHQX1 x7_75_tmp1_reg_13_ ( .D(N285), .CK(clk), .RN(rstn), .Q(
        x7_75_tmp1[13]) );
  DFFRHQX1 x7_75_tmp1_reg_12_ ( .D(N284), .CK(clk), .RN(rstn), .Q(
        x7_75_tmp1[12]) );
  DFFRHQX1 x7_75_tmp1_reg_11_ ( .D(N283), .CK(clk), .RN(rstn), .Q(
        x7_75_tmp1[11]) );
  DFFRHQX1 x7_75_tmp1_reg_10_ ( .D(N282), .CK(clk), .RN(rstn), .Q(
        x7_75_tmp1[10]) );
  DFFRHQX1 x6_75_tmp1_reg_14_ ( .D(N201), .CK(clk), .RN(rstn), .Q(
        x6_75_tmp1[14]) );
  DFFRHQX1 x6_75_tmp1_reg_13_ ( .D(N200), .CK(clk), .RN(rstn), .Q(
        x6_75_tmp1[13]) );
  DFFRHQX1 x6_75_tmp1_reg_12_ ( .D(N199), .CK(clk), .RN(rstn), .Q(
        x6_75_tmp1[12]) );
  DFFRHQX1 x6_75_tmp1_reg_11_ ( .D(N198), .CK(clk), .RN(rstn), .Q(
        x6_75_tmp1[11]) );
  DFFRHQX1 x6_75_tmp1_reg_10_ ( .D(N197), .CK(clk), .RN(rstn), .Q(
        x6_75_tmp1[10]) );
  DFFRHQX1 x4_50_tmp1_reg_13_ ( .D(n74), .CK(clk), .RN(rstn), .Q(
        x4_50_tmp1[13]) );
  DFFRHQX1 x4_50_tmp1_reg_12_ ( .D(n73), .CK(clk), .RN(rstn), .Q(
        x4_50_tmp1[12]) );
  DFFRHQX1 x4_50_tmp1_reg_11_ ( .D(n72), .CK(clk), .RN(rstn), .Q(
        x4_50_tmp1[11]) );
  DFFRHQX1 x4_50_tmp1_reg_10_ ( .D(n71), .CK(clk), .RN(rstn), .Q(
        x4_50_tmp1[10]) );
  DFFRHQX1 x4_50_tmp1_reg_9_ ( .D(n70), .CK(clk), .RN(rstn), .Q(x4_50_tmp1[9])
         );
  DFFRHQX1 x6_50_tmp1_reg_13_ ( .D(n48), .CK(clk), .RN(rstn), .Q(
        x6_50_tmp1[13]) );
  DFFRHQX1 x6_50_tmp1_reg_12_ ( .D(n47), .CK(clk), .RN(rstn), .Q(
        x6_50_tmp1[12]) );
  DFFRHQX1 x6_50_tmp1_reg_11_ ( .D(n46), .CK(clk), .RN(rstn), .Q(
        x6_50_tmp1[11]) );
  DFFRHQX1 x6_50_tmp1_reg_10_ ( .D(n45), .CK(clk), .RN(rstn), .Q(
        x6_50_tmp1[10]) );
  DFFRHQX1 x6_50_tmp1_reg_9_ ( .D(n44), .CK(clk), .RN(rstn), .Q(x6_50_tmp1[9])
         );
  DFFRHQX1 x5_50_tmp1_reg_13_ ( .D(n61), .CK(clk), .RN(rstn), .Q(
        x5_50_tmp1[13]) );
  DFFRHQX1 x5_50_tmp1_reg_12_ ( .D(n60), .CK(clk), .RN(rstn), .Q(
        x5_50_tmp1[12]) );
  DFFRHQX1 x5_50_tmp1_reg_11_ ( .D(n59), .CK(clk), .RN(rstn), .Q(
        x5_50_tmp1[11]) );
  DFFRHQX1 x5_50_tmp1_reg_10_ ( .D(n58), .CK(clk), .RN(rstn), .Q(
        x5_50_tmp1[10]) );
  DFFRHQX1 x5_50_tmp1_reg_9_ ( .D(n57), .CK(clk), .RN(rstn), .Q(x5_50_tmp1[9])
         );
  DFFRHQX1 x7_50_tmp1_reg_13_ ( .D(n8), .CK(clk), .RN(rstn), .Q(x7_50_tmp1[13]) );
  DFFRHQX1 x7_50_tmp1_reg_12_ ( .D(n7), .CK(clk), .RN(rstn), .Q(x7_50_tmp1[12]) );
  DFFRHQX1 x7_50_tmp1_reg_11_ ( .D(n6), .CK(clk), .RN(rstn), .Q(x7_50_tmp1[11]) );
  DFFRHQX1 x7_50_tmp1_reg_10_ ( .D(n5), .CK(clk), .RN(rstn), .Q(x7_50_tmp1[10]) );
  DFFRHQX1 x7_50_tmp1_reg_9_ ( .D(n4), .CK(clk), .RN(rstn), .Q(x7_50_tmp1[9])
         );
  DFFRHQX1 x4_18_tmp1_reg_12_ ( .D(n74), .CK(clk), .RN(rstn), .Q(
        x4_18_tmp1[12]) );
  DFFRHQX1 x4_18_tmp1_reg_11_ ( .D(n73), .CK(clk), .RN(rstn), .Q(
        x4_18_tmp1[11]) );
  DFFRHQX1 x4_18_tmp1_reg_10_ ( .D(n72), .CK(clk), .RN(rstn), .Q(
        x4_18_tmp1[10]) );
  DFFRHQX1 x4_18_tmp1_reg_9_ ( .D(n71), .CK(clk), .RN(rstn), .Q(x4_18_tmp1[9])
         );
  DFFRHQX1 x4_18_tmp1_reg_8_ ( .D(n70), .CK(clk), .RN(rstn), .Q(x4_18_tmp1[8])
         );
  DFFRHQX1 x5_18_tmp1_reg_12_ ( .D(n61), .CK(clk), .RN(rstn), .Q(
        x5_18_tmp1[12]) );
  DFFRHQX1 x5_18_tmp1_reg_11_ ( .D(n60), .CK(clk), .RN(rstn), .Q(
        x5_18_tmp1[11]) );
  DFFRHQX1 x5_18_tmp1_reg_10_ ( .D(n59), .CK(clk), .RN(rstn), .Q(
        x5_18_tmp1[10]) );
  DFFRHQX1 x5_18_tmp1_reg_9_ ( .D(n58), .CK(clk), .RN(rstn), .Q(x5_18_tmp1[9])
         );
  DFFRHQX1 x5_18_tmp1_reg_8_ ( .D(n57), .CK(clk), .RN(rstn), .Q(x5_18_tmp1[8])
         );
  DFFRHQX1 x6_18_tmp1_reg_12_ ( .D(n48), .CK(clk), .RN(rstn), .Q(
        x6_18_tmp1[12]) );
  DFFRHQX1 x6_18_tmp1_reg_11_ ( .D(n47), .CK(clk), .RN(rstn), .Q(
        x6_18_tmp1[11]) );
  DFFRHQX1 x6_18_tmp1_reg_10_ ( .D(n46), .CK(clk), .RN(rstn), .Q(
        x6_18_tmp1[10]) );
  DFFRHQX1 x6_18_tmp1_reg_9_ ( .D(n45), .CK(clk), .RN(rstn), .Q(x6_18_tmp1[9])
         );
  DFFRHQX1 x6_18_tmp1_reg_8_ ( .D(n44), .CK(clk), .RN(rstn), .Q(x6_18_tmp1[8])
         );
  DFFRHQX1 x7_18_tmp1_reg_12_ ( .D(n8), .CK(clk), .RN(rstn), .Q(x7_18_tmp1[12]) );
  DFFRHQX1 x7_18_tmp1_reg_11_ ( .D(n7), .CK(clk), .RN(rstn), .Q(x7_18_tmp1[11]) );
  DFFRHQX1 x7_18_tmp1_reg_10_ ( .D(n6), .CK(clk), .RN(rstn), .Q(x7_18_tmp1[10]) );
  DFFRHQX1 x7_18_tmp1_reg_9_ ( .D(n5), .CK(clk), .RN(rstn), .Q(x7_18_tmp1[9])
         );
  DFFRHQX1 x7_18_tmp1_reg_8_ ( .D(n4), .CK(clk), .RN(rstn), .Q(x7_18_tmp1[8])
         );
  DFFRHQX1 x5_18_reg_16_ ( .D(N530), .CK(clk), .RN(rstn), .Q(x5_18[16]) );
  DFFRHQX1 x5_18_reg_15_ ( .D(N529), .CK(clk), .RN(rstn), .Q(x5_18[15]) );
  DFFRHQX1 x5_18_reg_14_ ( .D(N528), .CK(clk), .RN(rstn), .Q(x5_18[14]) );
  DFFRHQX1 x5_18_reg_13_ ( .D(N527), .CK(clk), .RN(rstn), .Q(x5_18[13]) );
  DFFRHQX1 x6_18_reg_15_ ( .D(N618), .CK(clk), .RN(rstn), .Q(x6_18[15]) );
  DFFRHQX1 x6_18_reg_14_ ( .D(N617), .CK(clk), .RN(rstn), .Q(x6_18[14]) );
  DFFRHQX1 x6_18_reg_13_ ( .D(N616), .CK(clk), .RN(rstn), .Q(x6_18[13]) );
  DFFRHQX1 x6_18_reg_12_ ( .D(N615), .CK(clk), .RN(rstn), .Q(x6_18[12]) );
  DFFRHQX1 x6_18_reg_11_ ( .D(N614), .CK(clk), .RN(rstn), .Q(x6_18[11]) );
  DFFRHQX1 x4_18_reg_15_ ( .D(N440), .CK(clk), .RN(rstn), .Q(x4_18[15]) );
  DFFRHQX1 x4_18_reg_14_ ( .D(N439), .CK(clk), .RN(rstn), .Q(x4_18[14]) );
  DFFRHQX1 x4_18_reg_13_ ( .D(N438), .CK(clk), .RN(rstn), .Q(x4_18[13]) );
  DFFRHQX1 x4_18_reg_12_ ( .D(N437), .CK(clk), .RN(rstn), .Q(x4_18[12]) );
  DFFRHQX1 x4_18_reg_11_ ( .D(N436), .CK(clk), .RN(rstn), .Q(x4_18[11]) );
  DFFRHQX1 x4_89_tmp1_reg_14_ ( .D(N31), .CK(clk), .RN(rstn), .Q(
        x4_89_tmp1[14]) );
  DFFRHQX1 x4_89_tmp1_reg_13_ ( .D(N30), .CK(clk), .RN(rstn), .Q(
        x4_89_tmp1[13]) );
  DFFRHQX1 x4_89_tmp1_reg_12_ ( .D(N29), .CK(clk), .RN(rstn), .Q(
        x4_89_tmp1[12]) );
  DFFRHQX1 x4_89_tmp1_reg_11_ ( .D(N28), .CK(clk), .RN(rstn), .Q(
        x4_89_tmp1[11]) );
  DFFRHQX1 x4_89_tmp1_reg_10_ ( .D(N27), .CK(clk), .RN(rstn), .Q(
        x4_89_tmp1[10]) );
  DFFRHQX1 x4_89_reg_15_ ( .D(N372), .CK(clk), .RN(rstn), .Q(x4_89[15]) );
  DFFRHQX1 x4_89_reg_14_ ( .D(N371), .CK(clk), .RN(rstn), .Q(x4_89[14]) );
  DFFRHQX1 x4_89_reg_13_ ( .D(N370), .CK(clk), .RN(rstn), .Q(x4_89[13]) );
  DFFRHQX1 x4_89_reg_12_ ( .D(N369), .CK(clk), .RN(rstn), .Q(x4_89[12]) );
  DFFRHQX1 x4_89_reg_11_ ( .D(N368), .CK(clk), .RN(rstn), .Q(x4_89[11]) );
  DFFRHQX1 x4_75_reg_15_ ( .D(N395), .CK(clk), .RN(rstn), .Q(x4_75[15]) );
  DFFRHQX1 x4_75_reg_14_ ( .D(N394), .CK(clk), .RN(rstn), .Q(x4_75[14]) );
  DFFRHQX1 x4_75_reg_13_ ( .D(N393), .CK(clk), .RN(rstn), .Q(x4_75[13]) );
  DFFRHQX1 x4_75_reg_12_ ( .D(N392), .CK(clk), .RN(rstn), .Q(x4_75[12]) );
  DFFRHQX1 x4_75_reg_11_ ( .D(N391), .CK(clk), .RN(rstn), .Q(x4_75[11]) );
  DFFRHQX1 x5_75_reg_15_ ( .D(N484), .CK(clk), .RN(rstn), .Q(x5_75[15]) );
  DFFRHQX1 x5_75_reg_14_ ( .D(N483), .CK(clk), .RN(rstn), .Q(x5_75[14]) );
  DFFRHQX1 x5_75_reg_13_ ( .D(N482), .CK(clk), .RN(rstn), .Q(x5_75[13]) );
  DFFRHQX1 x5_75_reg_12_ ( .D(N481), .CK(clk), .RN(rstn), .Q(x5_75[12]) );
  DFFRHQX1 x5_75_reg_11_ ( .D(N480), .CK(clk), .RN(rstn), .Q(x5_75[11]) );
  DFFRHQX1 x6_75_reg_15_ ( .D(N573), .CK(clk), .RN(rstn), .Q(x6_75[15]) );
  DFFRHQX1 x6_75_reg_14_ ( .D(N572), .CK(clk), .RN(rstn), .Q(x6_75[14]) );
  DFFRHQX1 x6_75_reg_13_ ( .D(N571), .CK(clk), .RN(rstn), .Q(x6_75[13]) );
  DFFRHQX1 x6_75_reg_12_ ( .D(N570), .CK(clk), .RN(rstn), .Q(x6_75[12]) );
  DFFRHQX1 x6_75_reg_11_ ( .D(N569), .CK(clk), .RN(rstn), .Q(x6_75[11]) );
  DFFRHQX1 x4_50_reg_15_ ( .D(N418), .CK(clk), .RN(rstn), .Q(x4_50[15]) );
  DFFRHQX1 x4_50_reg_14_ ( .D(N417), .CK(clk), .RN(rstn), .Q(x4_50[14]) );
  DFFRHQX1 x4_50_reg_13_ ( .D(N416), .CK(clk), .RN(rstn), .Q(x4_50[13]) );
  DFFRHQX1 x4_50_reg_12_ ( .D(N415), .CK(clk), .RN(rstn), .Q(x4_50[12]) );
  DFFRHQX1 x4_50_reg_11_ ( .D(N414), .CK(clk), .RN(rstn), .Q(x4_50[11]) );
  DFFRHQX1 x5_tmp1_reg_16_ ( .D(N895), .CK(clk), .RN(rstn), .Q(x5_tmp1[16]) );
  DFFRHQX1 x5_tmp1_reg_15_ ( .D(N894), .CK(clk), .RN(rstn), .Q(x5_tmp1[15]) );
  DFFRHQX1 x5_tmp1_reg_14_ ( .D(N893), .CK(clk), .RN(rstn), .Q(x5_tmp1[14]) );
  DFFRHQX1 x5_tmp1_reg_13_ ( .D(N892), .CK(clk), .RN(rstn), .Q(x5_tmp1[13]) );
  DFFRHQX1 x5_tmp1_reg_12_ ( .D(N891), .CK(clk), .RN(rstn), .Q(x5_tmp1[12]) );
  DFFRHQX1 x6_tmp1_reg_16_ ( .D(N1061), .CK(clk), .RN(rstn), .Q(x6_tmp1[16])
         );
  DFFRHQX1 x6_tmp1_reg_15_ ( .D(N1060), .CK(clk), .RN(rstn), .Q(x6_tmp1[15])
         );
  DFFRHQX1 x6_tmp1_reg_14_ ( .D(N1059), .CK(clk), .RN(rstn), .Q(x6_tmp1[14])
         );
  DFFRHQX1 x6_tmp1_reg_13_ ( .D(N1058), .CK(clk), .RN(rstn), .Q(x6_tmp1[13])
         );
  DFFRHQX1 x6_tmp1_reg_12_ ( .D(N1057), .CK(clk), .RN(rstn), .Q(x6_tmp1[12])
         );
  DFFRHQX1 x7_tmp1_reg_16_ ( .D(N1158), .CK(clk), .RN(rstn), .Q(x7_tmp1[16])
         );
  DFFRHQX1 x7_tmp1_reg_15_ ( .D(N1157), .CK(clk), .RN(rstn), .Q(x7_tmp1[15])
         );
  DFFRHQX1 x7_tmp1_reg_14_ ( .D(N1156), .CK(clk), .RN(rstn), .Q(x7_tmp1[14])
         );
  DFFRHQX1 x7_tmp1_reg_13_ ( .D(N1155), .CK(clk), .RN(rstn), .Q(x7_tmp1[13])
         );
  DFFRHQX1 x7_tmp1_reg_12_ ( .D(N1154), .CK(clk), .RN(rstn), .Q(x7_tmp1[12])
         );
  DFFRHQX1 x4_tmp1_reg_16_ ( .D(N776), .CK(clk), .RN(rstn), .Q(x4_tmp1[16]) );
  DFFRHQX1 x4_tmp1_reg_15_ ( .D(N775), .CK(clk), .RN(rstn), .Q(x4_tmp1[15]) );
  DFFRHQX1 x4_tmp1_reg_14_ ( .D(N774), .CK(clk), .RN(rstn), .Q(x4_tmp1[14]) );
  DFFRHQX1 x4_tmp1_reg_13_ ( .D(N773), .CK(clk), .RN(rstn), .Q(x4_tmp1[13]) );
  DFFRHQX1 x4_tmp1_reg_12_ ( .D(N772), .CK(clk), .RN(rstn), .Q(x4_tmp1[12]) );
  DFFRHQX1 y6_tmp_reg_21_ ( .D(N1545), .CK(clk), .RN(rstn), .Q(y6_tmp[21]) );
  DFFRHQX1 y6_tmp_reg_20_ ( .D(N1544), .CK(clk), .RN(rstn), .Q(y6_tmp[20]) );
  DFFRHQX1 y6_tmp_reg_19_ ( .D(N1543), .CK(clk), .RN(rstn), .Q(y6_tmp[19]) );
  DFFRHQX1 y6_tmp_reg_18_ ( .D(N1542), .CK(clk), .RN(rstn), .Q(y6_tmp[18]) );
  DFFRHQX1 y6_tmp_reg_17_ ( .D(N1541), .CK(clk), .RN(rstn), .Q(y6_tmp[17]) );
  DFFRHQX1 y7_tmp_reg_21_ ( .D(N1622), .CK(clk), .RN(rstn), .Q(y7_tmp[21]) );
  DFFRHQX1 y7_tmp_reg_20_ ( .D(N1621), .CK(clk), .RN(rstn), .Q(y7_tmp[20]) );
  DFFRHQX1 y7_tmp_reg_19_ ( .D(N1620), .CK(clk), .RN(rstn), .Q(y7_tmp[19]) );
  DFFRHQX1 y7_tmp_reg_18_ ( .D(N1619), .CK(clk), .RN(rstn), .Q(y7_tmp[18]) );
  DFFRHQX1 y0_tmp_reg_23_ ( .D(N1238), .CK(clk), .RN(rstn), .Q(y0_tmp[23]) );
  DFFRHQX1 y0_tmp_reg_22_ ( .D(N1237), .CK(clk), .RN(rstn), .Q(y0_tmp[22]) );
  DFFRHQX1 y0_tmp_reg_21_ ( .D(N1236), .CK(clk), .RN(rstn), .Q(y0_tmp[21]) );
  DFFRHQX1 y0_tmp_reg_20_ ( .D(N1235), .CK(clk), .RN(rstn), .Q(y0_tmp[20]) );
  DFFRHQX1 y0_tmp_reg_19_ ( .D(N1234), .CK(clk), .RN(rstn), .Q(y0_tmp[19]) );
  DFFRHQX1 y1_tmp_reg_23_ ( .D(N1264), .CK(clk), .RN(rstn), .Q(y1_tmp[23]) );
  DFFRHQX1 y1_tmp_reg_22_ ( .D(N1263), .CK(clk), .RN(rstn), .Q(y1_tmp[22]) );
  DFFRHQX1 y1_tmp_reg_21_ ( .D(N1262), .CK(clk), .RN(rstn), .Q(y1_tmp[21]) );
  DFFRHQX1 y1_tmp_reg_20_ ( .D(N1261), .CK(clk), .RN(rstn), .Q(y1_tmp[20]) );
  DFFRHQX1 y1_tmp_reg_19_ ( .D(N1260), .CK(clk), .RN(rstn), .Q(y1_tmp[19]) );
  DFFRHQX1 y2_tmp_reg_23_ ( .D(N1290), .CK(clk), .RN(rstn), .Q(y2_tmp[23]) );
  DFFRHQX1 y2_tmp_reg_22_ ( .D(N1289), .CK(clk), .RN(rstn), .Q(y2_tmp[22]) );
  DFFRHQX1 y2_tmp_reg_21_ ( .D(N1288), .CK(clk), .RN(rstn), .Q(y2_tmp[21]) );
  DFFRHQX1 y2_tmp_reg_20_ ( .D(N1287), .CK(clk), .RN(rstn), .Q(y2_tmp[20]) );
  DFFRHQX1 y2_tmp_reg_19_ ( .D(N1286), .CK(clk), .RN(rstn), .Q(y2_tmp[19]) );
  DFFRHQX1 y3_tmp_reg_23_ ( .D(N1316), .CK(clk), .RN(rstn), .Q(y3_tmp[23]) );
  DFFRHQX1 y3_tmp_reg_22_ ( .D(N1315), .CK(clk), .RN(rstn), .Q(y3_tmp[22]) );
  DFFRHQX1 y3_tmp_reg_21_ ( .D(N1314), .CK(clk), .RN(rstn), .Q(y3_tmp[21]) );
  DFFRHQX1 y3_tmp_reg_20_ ( .D(N1313), .CK(clk), .RN(rstn), .Q(y3_tmp[20]) );
  DFFRHQX1 y3_tmp_reg_19_ ( .D(N1312), .CK(clk), .RN(rstn), .Q(y3_tmp[19]) );
  DFFRHQX1 y4_tmp_reg_21_ ( .D(N1391), .CK(clk), .RN(rstn), .Q(y4_tmp[21]) );
  DFFRHQX1 y4_tmp_reg_20_ ( .D(N1390), .CK(clk), .RN(rstn), .Q(y4_tmp[20]) );
  DFFRHQX1 y4_tmp_reg_19_ ( .D(N1389), .CK(clk), .RN(rstn), .Q(y4_tmp[19]) );
  DFFRHQX1 y4_tmp_reg_18_ ( .D(N1388), .CK(clk), .RN(rstn), .Q(y4_tmp[18]) );
  DFFRHQX1 y4_tmp_reg_17_ ( .D(N1387), .CK(clk), .RN(rstn), .Q(y4_tmp[17]) );
  DFFRHQX1 y5_tmp_reg_21_ ( .D(N1468), .CK(clk), .RN(rstn), .Q(y5_tmp[21]) );
  DFFRHQX1 y5_tmp_reg_20_ ( .D(N1467), .CK(clk), .RN(rstn), .Q(y5_tmp[20]) );
  DFFRHQX1 y5_tmp_reg_19_ ( .D(N1466), .CK(clk), .RN(rstn), .Q(y5_tmp[19]) );
  DFFRHQX1 y5_tmp_reg_18_ ( .D(N1465), .CK(clk), .RN(rstn), .Q(y5_tmp[18]) );
  DFFRHQX1 y5_tmp_reg_17_ ( .D(N1464), .CK(clk), .RN(rstn), .Q(y5_tmp[17]) );
  DFFRHQX1 mode_delay2_reg_0_ ( .D(mode_delay1[0]), .CK(clk), .RN(rstn), .Q(
        mode_delay2[0]) );
  DFFRHQX1 x7_50_reg_15_ ( .D(N685), .CK(clk), .RN(rstn), .Q(x7_50[15]) );
  DFFRHQX1 x7_50_reg_14_ ( .D(N684), .CK(clk), .RN(rstn), .Q(x7_50[14]) );
  DFFRHQX1 x7_50_reg_13_ ( .D(N683), .CK(clk), .RN(rstn), .Q(x7_50[13]) );
  DFFRHQX1 x7_50_reg_12_ ( .D(N682), .CK(clk), .RN(rstn), .Q(x7_50[12]) );
  DFFRHQX1 x5_89_reg_15_ ( .D(N461), .CK(clk), .RN(rstn), .Q(x5_89[15]) );
  DFFRHQX1 x5_89_reg_14_ ( .D(N460), .CK(clk), .RN(rstn), .Q(x5_89[14]) );
  DFFRHQX1 x5_89_reg_13_ ( .D(N459), .CK(clk), .RN(rstn), .Q(x5_89[13]) );
  DFFRHQX1 x5_89_reg_12_ ( .D(N458), .CK(clk), .RN(rstn), .Q(x5_89[12]) );
  DFFRHQX1 x7_89_reg_15_ ( .D(N639), .CK(clk), .RN(rstn), .Q(x7_89[15]) );
  DFFRHQX1 x7_89_reg_14_ ( .D(N638), .CK(clk), .RN(rstn), .Q(x7_89[14]) );
  DFFRHQX1 x7_89_reg_13_ ( .D(N637), .CK(clk), .RN(rstn), .Q(x7_89[13]) );
  DFFRHQX1 x7_89_reg_12_ ( .D(N636), .CK(clk), .RN(rstn), .Q(x7_89[12]) );
  DFFRHQX1 x5_50_reg_15_ ( .D(N507), .CK(clk), .RN(rstn), .Q(x5_50[15]) );
  DFFRHQX1 x5_50_reg_14_ ( .D(N506), .CK(clk), .RN(rstn), .Q(x5_50[14]) );
  DFFRHQX1 x5_50_reg_13_ ( .D(N505), .CK(clk), .RN(rstn), .Q(x5_50[13]) );
  DFFRHQX1 x5_50_reg_12_ ( .D(N504), .CK(clk), .RN(rstn), .Q(x5_50[12]) );
  DFFRHQX1 x6_89_tmp2_reg_13_ ( .D(N223), .CK(clk), .RN(rstn), .Q(
        x6_89_tmp2[13]) );
  DFFRHQX1 x6_89_tmp2_reg_12_ ( .D(N222), .CK(clk), .RN(rstn), .Q(
        x6_89_tmp2[12]) );
  DFFRHQX1 x6_89_tmp2_reg_11_ ( .D(N221), .CK(clk), .RN(rstn), .Q(
        x6_89_tmp2[11]) );
  DFFRHQX1 x6_89_tmp2_reg_10_ ( .D(N220), .CK(clk), .RN(rstn), .Q(
        x6_89_tmp2[10]) );
  DFFRHQX1 x5_89_tmp2_reg_13_ ( .D(N138), .CK(clk), .RN(rstn), .Q(
        x5_89_tmp2[13]) );
  DFFRHQX1 x5_89_tmp2_reg_12_ ( .D(N137), .CK(clk), .RN(rstn), .Q(
        x5_89_tmp2[12]) );
  DFFRHQX1 x5_89_tmp2_reg_11_ ( .D(N136), .CK(clk), .RN(rstn), .Q(
        x5_89_tmp2[11]) );
  DFFRHQX1 x5_89_tmp2_reg_10_ ( .D(N135), .CK(clk), .RN(rstn), .Q(
        x5_89_tmp2[10]) );
  DFFRHQX1 x4_89_tmp2_reg_13_ ( .D(N53), .CK(clk), .RN(rstn), .Q(
        x4_89_tmp2[13]) );
  DFFRHQX1 x4_89_tmp2_reg_12_ ( .D(N52), .CK(clk), .RN(rstn), .Q(
        x4_89_tmp2[12]) );
  DFFRHQX1 x4_89_tmp2_reg_11_ ( .D(N51), .CK(clk), .RN(rstn), .Q(
        x4_89_tmp2[11]) );
  DFFRHQX1 x4_89_tmp2_reg_10_ ( .D(N50), .CK(clk), .RN(rstn), .Q(
        x4_89_tmp2[10]) );
  DFFRHQX1 x7_89_tmp2_reg_13_ ( .D(N308), .CK(clk), .RN(rstn), .Q(
        x7_89_tmp2[13]) );
  DFFRHQX1 x7_89_tmp2_reg_12_ ( .D(N307), .CK(clk), .RN(rstn), .Q(
        x7_89_tmp2[12]) );
  DFFRHQX1 x7_89_tmp2_reg_11_ ( .D(N306), .CK(clk), .RN(rstn), .Q(
        x7_89_tmp2[11]) );
  DFFRHQX1 x7_89_tmp2_reg_10_ ( .D(N305), .CK(clk), .RN(rstn), .Q(
        x7_89_tmp2[10]) );
  DFFRHQX1 x4_75_tmp2_reg_13_ ( .D(N74), .CK(clk), .RN(rstn), .Q(
        x4_75_tmp2[13]) );
  DFFRHQX1 x4_75_tmp2_reg_12_ ( .D(N73), .CK(clk), .RN(rstn), .Q(
        x4_75_tmp2[12]) );
  DFFRHQX1 x4_75_tmp2_reg_11_ ( .D(N72), .CK(clk), .RN(rstn), .Q(
        x4_75_tmp2[11]) );
  DFFRHQX1 x4_75_tmp2_reg_10_ ( .D(N71), .CK(clk), .RN(rstn), .Q(
        x4_75_tmp2[10]) );
  DFFRHQX1 x5_75_tmp2_reg_13_ ( .D(N159), .CK(clk), .RN(rstn), .Q(
        x5_75_tmp2[13]) );
  DFFRHQX1 x5_75_tmp2_reg_12_ ( .D(N158), .CK(clk), .RN(rstn), .Q(
        x5_75_tmp2[12]) );
  DFFRHQX1 x5_75_tmp2_reg_11_ ( .D(N157), .CK(clk), .RN(rstn), .Q(
        x5_75_tmp2[11]) );
  DFFRHQX1 x5_75_tmp2_reg_10_ ( .D(N156), .CK(clk), .RN(rstn), .Q(
        x5_75_tmp2[10]) );
  DFFRHQX1 x6_75_tmp2_reg_13_ ( .D(N244), .CK(clk), .RN(rstn), .Q(
        x6_75_tmp2[13]) );
  DFFRHQX1 x6_75_tmp2_reg_12_ ( .D(N243), .CK(clk), .RN(rstn), .Q(
        x6_75_tmp2[12]) );
  DFFRHQX1 x6_75_tmp2_reg_11_ ( .D(N242), .CK(clk), .RN(rstn), .Q(
        x6_75_tmp2[11]) );
  DFFRHQX1 x6_75_tmp2_reg_10_ ( .D(N241), .CK(clk), .RN(rstn), .Q(
        x6_75_tmp2[10]) );
  DFFRHQX1 x7_75_tmp2_reg_13_ ( .D(N329), .CK(clk), .RN(rstn), .Q(
        x7_75_tmp2[13]) );
  DFFRHQX1 x7_75_tmp2_reg_12_ ( .D(N328), .CK(clk), .RN(rstn), .Q(
        x7_75_tmp2[12]) );
  DFFRHQX1 x7_75_tmp2_reg_11_ ( .D(N327), .CK(clk), .RN(rstn), .Q(
        x7_75_tmp2[11]) );
  DFFRHQX1 x7_75_tmp2_reg_10_ ( .D(N326), .CK(clk), .RN(rstn), .Q(
        x7_75_tmp2[10]) );
  DFFRHQX1 x4_50_tmp2_reg_12_ ( .D(N93), .CK(clk), .RN(rstn), .Q(
        x4_50_tmp2[12]) );
  DFFRHQX1 x4_50_tmp2_reg_11_ ( .D(N92), .CK(clk), .RN(rstn), .Q(
        x4_50_tmp2[11]) );
  DFFRHQX1 x4_50_tmp2_reg_10_ ( .D(N91), .CK(clk), .RN(rstn), .Q(
        x4_50_tmp2[10]) );
  DFFRHQX1 x4_50_tmp2_reg_9_ ( .D(N90), .CK(clk), .RN(rstn), .Q(x4_50_tmp2[9])
         );
  DFFRHQX1 x6_50_tmp2_reg_12_ ( .D(N263), .CK(clk), .RN(rstn), .Q(
        x6_50_tmp2[12]) );
  DFFRHQX1 x6_50_tmp2_reg_11_ ( .D(N262), .CK(clk), .RN(rstn), .Q(
        x6_50_tmp2[11]) );
  DFFRHQX1 x6_50_tmp2_reg_10_ ( .D(N261), .CK(clk), .RN(rstn), .Q(
        x6_50_tmp2[10]) );
  DFFRHQX1 x6_50_tmp2_reg_9_ ( .D(N260), .CK(clk), .RN(rstn), .Q(x6_50_tmp2[9]) );
  DFFRHQX1 x6_50_reg_11_ ( .D(N592), .CK(clk), .RN(rstn), .Q(x6_50[11]) );
  DFFRHQX1 x6_50_reg_12_ ( .D(N593), .CK(clk), .RN(rstn), .Q(x6_50[12]) );
  DFFRHQX1 x6_50_reg_13_ ( .D(N594), .CK(clk), .RN(rstn), .Q(x6_50[13]) );
  DFFRHQX1 x6_50_reg_14_ ( .D(N595), .CK(clk), .RN(rstn), .Q(x6_50[14]) );
  DFFRHQX1 x5_50_tmp2_reg_12_ ( .D(N178), .CK(clk), .RN(rstn), .Q(
        x5_50_tmp2[12]) );
  DFFRHQX1 x5_50_tmp2_reg_11_ ( .D(N177), .CK(clk), .RN(rstn), .Q(
        x5_50_tmp2[11]) );
  DFFRHQX1 x5_50_tmp2_reg_10_ ( .D(N176), .CK(clk), .RN(rstn), .Q(
        x5_50_tmp2[10]) );
  DFFRHQX1 x5_50_tmp2_reg_9_ ( .D(N175), .CK(clk), .RN(rstn), .Q(x5_50_tmp2[9]) );
  DFFRHQX1 x7_50_tmp2_reg_12_ ( .D(N348), .CK(clk), .RN(rstn), .Q(
        x7_50_tmp2[12]) );
  DFFRHQX1 x7_50_tmp2_reg_11_ ( .D(N347), .CK(clk), .RN(rstn), .Q(
        x7_50_tmp2[11]) );
  DFFRHQX1 x7_50_tmp2_reg_10_ ( .D(N346), .CK(clk), .RN(rstn), .Q(
        x7_50_tmp2[10]) );
  DFFRHQX1 x7_50_tmp2_reg_9_ ( .D(N345), .CK(clk), .RN(rstn), .Q(x7_50_tmp2[9]) );
  DFFRHQX1 x4_18_tmp2_reg_11_ ( .D(n76), .CK(clk), .RN(rstn), .Q(
        x4_18_tmp2[11]) );
  DFFRHQX1 x4_18_tmp2_reg_10_ ( .D(n75), .CK(clk), .RN(rstn), .Q(
        x4_18_tmp2[10]) );
  DFFRHQX1 x4_18_tmp2_reg_9_ ( .D(n74), .CK(clk), .RN(rstn), .Q(x4_18_tmp2[9])
         );
  DFFRHQX1 x4_18_tmp2_reg_8_ ( .D(n73), .CK(clk), .RN(rstn), .Q(x4_18_tmp2[8])
         );
  DFFRHQX1 x6_18_tmp2_reg_11_ ( .D(n50), .CK(clk), .RN(rstn), .Q(
        x6_18_tmp2[11]) );
  DFFRHQX1 x6_18_tmp2_reg_10_ ( .D(n49), .CK(clk), .RN(rstn), .Q(
        x6_18_tmp2[10]) );
  DFFRHQX1 x6_18_tmp2_reg_9_ ( .D(n48), .CK(clk), .RN(rstn), .Q(x6_18_tmp2[9])
         );
  DFFRHQX1 x6_18_tmp2_reg_8_ ( .D(n47), .CK(clk), .RN(rstn), .Q(x6_18_tmp2[8])
         );
  DFFRHQX1 x5_18_tmp2_reg_11_ ( .D(n63), .CK(clk), .RN(rstn), .Q(
        x5_18_tmp2[11]) );
  DFFRHQX1 x5_18_tmp2_reg_10_ ( .D(n62), .CK(clk), .RN(rstn), .Q(
        x5_18_tmp2[10]) );
  DFFRHQX1 x5_18_tmp2_reg_9_ ( .D(n61), .CK(clk), .RN(rstn), .Q(x5_18_tmp2[9])
         );
  DFFRHQX1 x5_18_tmp2_reg_8_ ( .D(n60), .CK(clk), .RN(rstn), .Q(x5_18_tmp2[8])
         );
  DFFRHQX1 x7_18_tmp2_reg_11_ ( .D(n37), .CK(clk), .RN(rstn), .Q(
        x7_18_tmp2[11]) );
  DFFRHQX1 x7_18_tmp2_reg_10_ ( .D(n36), .CK(clk), .RN(rstn), .Q(
        x7_18_tmp2[10]) );
  DFFRHQX1 x7_18_tmp2_reg_9_ ( .D(n8), .CK(clk), .RN(rstn), .Q(x7_18_tmp2[9])
         );
  DFFRHQX1 x7_18_tmp2_reg_8_ ( .D(n7), .CK(clk), .RN(rstn), .Q(x7_18_tmp2[8])
         );
  DFFRHQX1 x7_18_reg_14_ ( .D(N706), .CK(clk), .RN(rstn), .Q(x7_18[14]) );
  DFFRHQX1 x7_18_reg_13_ ( .D(N705), .CK(clk), .RN(rstn), .Q(x7_18[13]) );
  DFFRHQX1 x7_18_reg_12_ ( .D(N704), .CK(clk), .RN(rstn), .Q(x7_18[12]) );
  DFFRHQX1 x7_18_reg_11_ ( .D(N703), .CK(clk), .RN(rstn), .Q(x7_18[11]) );
  DFFRHQX1 x6_89_reg_16_ ( .D(N551), .CK(clk), .RN(rstn), .Q(x6_89[16]) );
  DFFRHQX1 x6_89_reg_15_ ( .D(N550), .CK(clk), .RN(rstn), .Q(x6_89[15]) );
  DFFRHQX1 x6_89_reg_14_ ( .D(N549), .CK(clk), .RN(rstn), .Q(x6_89[14]) );
  DFFRHQX1 x6_89_reg_13_ ( .D(N548), .CK(clk), .RN(rstn), .Q(x6_89[13]) );
  DFFRHQX1 x6_89_reg_12_ ( .D(N547), .CK(clk), .RN(rstn), .Q(x6_89[12]) );
  DFFRHQX1 x7_75_reg_14_ ( .D(N661), .CK(clk), .RN(rstn), .Q(x7_75[14]) );
  DFFRHQX1 x7_75_reg_13_ ( .D(N660), .CK(clk), .RN(rstn), .Q(x7_75[13]) );
  DFFRHQX1 x7_75_reg_12_ ( .D(N659), .CK(clk), .RN(rstn), .Q(x7_75[12]) );
  DFFRHQX1 x7_75_reg_11_ ( .D(N658), .CK(clk), .RN(rstn), .Q(x7_75[11]) );
  DFFRHQX1 x4_tmp2_reg_15_ ( .D(N845), .CK(clk), .RN(rstn), .Q(x4_tmp2[15]) );
  DFFRHQX1 x4_tmp2_reg_14_ ( .D(N844), .CK(clk), .RN(rstn), .Q(x4_tmp2[14]) );
  DFFRHQX1 x4_tmp2_reg_13_ ( .D(N843), .CK(clk), .RN(rstn), .Q(x4_tmp2[13]) );
  DFFRHQX1 x4_tmp2_reg_12_ ( .D(N842), .CK(clk), .RN(rstn), .Q(x4_tmp2[12]) );
  DFFRHQX1 x5_tmp2_reg_15_ ( .D(N965), .CK(clk), .RN(rstn), .Q(x5_tmp2[15]) );
  DFFRHQX1 x5_tmp2_reg_14_ ( .D(N964), .CK(clk), .RN(rstn), .Q(x5_tmp2[14]) );
  DFFRHQX1 x5_tmp2_reg_13_ ( .D(N963), .CK(clk), .RN(rstn), .Q(x5_tmp2[13]) );
  DFFRHQX1 x5_tmp2_reg_12_ ( .D(N962), .CK(clk), .RN(rstn), .Q(x5_tmp2[12]) );
  DFFRHQX1 x6_tmp2_reg_15_ ( .D(N1108), .CK(clk), .RN(rstn), .Q(x6_tmp2[15])
         );
  DFFRHQX1 x6_tmp2_reg_14_ ( .D(N1107), .CK(clk), .RN(rstn), .Q(x6_tmp2[14])
         );
  DFFRHQX1 x6_tmp2_reg_13_ ( .D(N1106), .CK(clk), .RN(rstn), .Q(x6_tmp2[13])
         );
  DFFRHQX1 x6_tmp2_reg_12_ ( .D(N1105), .CK(clk), .RN(rstn), .Q(x6_tmp2[12])
         );
  DFFRHQX1 x7_tmp2_reg_15_ ( .D(N1181), .CK(clk), .RN(rstn), .Q(x7_tmp2[15])
         );
  DFFRHQX1 x7_tmp2_reg_14_ ( .D(N1180), .CK(clk), .RN(rstn), .Q(x7_tmp2[14])
         );
  DFFRHQX1 x7_tmp2_reg_13_ ( .D(N1179), .CK(clk), .RN(rstn), .Q(x7_tmp2[13])
         );
  DFFRHQX1 x7_tmp2_reg_12_ ( .D(N1178), .CK(clk), .RN(rstn), .Q(x7_tmp2[12])
         );
  DFFRHQX1 x7_tmp_reg_14_ ( .D(N1204), .CK(clk), .RN(rstn), .Q(x7_tmp[14]) );
  DFFRHQX1 x7_tmp_reg_15_ ( .D(N1205), .CK(clk), .RN(rstn), .Q(x7_tmp[15]) );
  DFFRHQX1 x7_tmp_reg_16_ ( .D(N1206), .CK(clk), .RN(rstn), .Q(x7_tmp[16]) );
  DFFRHQX1 x7_tmp_reg_17_ ( .D(N1207), .CK(clk), .RN(rstn), .Q(x7_tmp[17]) );
  DFFRHQX1 x5_tmp_reg_17_ ( .D(N991), .CK(clk), .RN(rstn), .Q(x5_tmp[17]) );
  DFFRHQX1 x5_tmp_reg_16_ ( .D(N990), .CK(clk), .RN(rstn), .Q(x5_tmp[16]) );
  DFFRHQX1 x5_tmp_reg_15_ ( .D(N989), .CK(clk), .RN(rstn), .Q(x5_tmp[15]) );
  DFFRHQX1 x5_tmp_reg_14_ ( .D(N988), .CK(clk), .RN(rstn), .Q(x5_tmp[14]) );
  DFFRHQX1 x6_tmp_reg_17_ ( .D(N1134), .CK(clk), .RN(rstn), .Q(x6_tmp[17]) );
  DFFRHQX1 x6_tmp_reg_16_ ( .D(N1133), .CK(clk), .RN(rstn), .Q(x6_tmp[16]) );
  DFFRHQX1 x6_tmp_reg_15_ ( .D(N1132), .CK(clk), .RN(rstn), .Q(x6_tmp[15]) );
  DFFRHQX1 x6_tmp_reg_14_ ( .D(N1131), .CK(clk), .RN(rstn), .Q(x6_tmp[14]) );
  DFFRHQX1 x4_tmp_reg_14_ ( .D(N868), .CK(clk), .RN(rstn), .Q(x4_tmp[14]) );
  DFFRHQX1 x4_tmp_reg_15_ ( .D(N869), .CK(clk), .RN(rstn), .Q(x4_tmp[15]) );
  DFFRHQX1 x4_tmp_reg_16_ ( .D(N870), .CK(clk), .RN(rstn), .Q(x4_tmp[16]) );
  DFFRHQX1 x4_tmp_reg_17_ ( .D(N871), .CK(clk), .RN(rstn), .Q(x4_tmp[17]) );
  DFFRHQX1 x7_89_tmp1_reg_9_ ( .D(N281), .CK(clk), .RN(rstn), .Q(x7_89_tmp1[9]) );
  DFFRHQX1 x7_89_tmp1_reg_8_ ( .D(N280), .CK(clk), .RN(rstn), .Q(x7_89_tmp1[8]) );
  DFFRHQX1 x7_89_tmp1_reg_7_ ( .D(N279), .CK(clk), .RN(rstn), .Q(x7_89_tmp1[7]) );
  DFFRHQX1 x7_89_tmp1_reg_6_ ( .D(N278), .CK(clk), .RN(rstn), .Q(x7_89_tmp1[6]) );
  DFFRHQX1 x6_89_tmp1_reg_9_ ( .D(N196), .CK(clk), .RN(rstn), .Q(x6_89_tmp1[9]) );
  DFFRHQX1 x6_89_tmp1_reg_8_ ( .D(N195), .CK(clk), .RN(rstn), .Q(x6_89_tmp1[8]) );
  DFFRHQX1 x6_89_tmp1_reg_7_ ( .D(N194), .CK(clk), .RN(rstn), .Q(x6_89_tmp1[7]) );
  DFFRHQX1 x6_89_tmp1_reg_6_ ( .D(N193), .CK(clk), .RN(rstn), .Q(x6_89_tmp1[6]) );
  DFFRHQX1 x5_89_tmp1_reg_9_ ( .D(N111), .CK(clk), .RN(rstn), .Q(x5_89_tmp1[9]) );
  DFFRHQX1 x5_89_tmp1_reg_8_ ( .D(N110), .CK(clk), .RN(rstn), .Q(x5_89_tmp1[8]) );
  DFFRHQX1 x5_89_tmp1_reg_7_ ( .D(N109), .CK(clk), .RN(rstn), .Q(x5_89_tmp1[7]) );
  DFFRHQX1 x5_89_tmp1_reg_6_ ( .D(N108), .CK(clk), .RN(rstn), .Q(x5_89_tmp1[6]) );
  DFFRHQX1 x5_75_tmp1_reg_9_ ( .D(N111), .CK(clk), .RN(rstn), .Q(x5_75_tmp1[9]) );
  DFFRHQX1 x5_75_tmp1_reg_8_ ( .D(N110), .CK(clk), .RN(rstn), .Q(x5_75_tmp1[8]) );
  DFFRHQX1 x5_75_tmp1_reg_7_ ( .D(N109), .CK(clk), .RN(rstn), .Q(x5_75_tmp1[7]) );
  DFFRHQX1 x5_75_tmp1_reg_6_ ( .D(N108), .CK(clk), .RN(rstn), .Q(x5_75_tmp1[6]) );
  DFFRHQX1 x4_75_tmp1_reg_9_ ( .D(N26), .CK(clk), .RN(rstn), .Q(x4_75_tmp1[9])
         );
  DFFRHQX1 x4_75_tmp1_reg_8_ ( .D(N25), .CK(clk), .RN(rstn), .Q(x4_75_tmp1[8])
         );
  DFFRHQX1 x4_75_tmp1_reg_7_ ( .D(N24), .CK(clk), .RN(rstn), .Q(x4_75_tmp1[7])
         );
  DFFRHQX1 x4_75_tmp1_reg_6_ ( .D(N23), .CK(clk), .RN(rstn), .Q(x4_75_tmp1[6])
         );
  DFFRHQX1 x7_75_tmp1_reg_9_ ( .D(N281), .CK(clk), .RN(rstn), .Q(x7_75_tmp1[9]) );
  DFFRHQX1 x7_75_tmp1_reg_8_ ( .D(N280), .CK(clk), .RN(rstn), .Q(x7_75_tmp1[8]) );
  DFFRHQX1 x7_75_tmp1_reg_7_ ( .D(N279), .CK(clk), .RN(rstn), .Q(x7_75_tmp1[7]) );
  DFFRHQX1 x7_75_tmp1_reg_6_ ( .D(N278), .CK(clk), .RN(rstn), .Q(x7_75_tmp1[6]) );
  DFFRHQX1 x6_75_tmp1_reg_9_ ( .D(N196), .CK(clk), .RN(rstn), .Q(x6_75_tmp1[9]) );
  DFFRHQX1 x6_75_tmp1_reg_8_ ( .D(N195), .CK(clk), .RN(rstn), .Q(x6_75_tmp1[8]) );
  DFFRHQX1 x6_75_tmp1_reg_7_ ( .D(N194), .CK(clk), .RN(rstn), .Q(x6_75_tmp1[7]) );
  DFFRHQX1 x6_75_tmp1_reg_6_ ( .D(N193), .CK(clk), .RN(rstn), .Q(x6_75_tmp1[6]) );
  DFFRHQX1 x4_50_tmp1_reg_8_ ( .D(n69), .CK(clk), .RN(rstn), .Q(x4_50_tmp1[8])
         );
  DFFRHQX1 x4_50_tmp1_reg_7_ ( .D(n68), .CK(clk), .RN(rstn), .Q(x4_50_tmp1[7])
         );
  DFFRHQX1 x4_50_tmp1_reg_6_ ( .D(x4[1]), .CK(clk), .RN(rstn), .Q(
        x4_50_tmp1[6]) );
  DFFRHQX1 x6_50_tmp1_reg_8_ ( .D(n43), .CK(clk), .RN(rstn), .Q(x6_50_tmp1[8])
         );
  DFFRHQX1 x6_50_tmp1_reg_7_ ( .D(n42), .CK(clk), .RN(rstn), .Q(x6_50_tmp1[7])
         );
  DFFRHQX1 x6_50_tmp1_reg_6_ ( .D(x6[1]), .CK(clk), .RN(rstn), .Q(
        x6_50_tmp1[6]) );
  DFFRHQX1 x5_50_tmp1_reg_8_ ( .D(n56), .CK(clk), .RN(rstn), .Q(x5_50_tmp1[8])
         );
  DFFRHQX1 x5_50_tmp1_reg_7_ ( .D(n55), .CK(clk), .RN(rstn), .Q(x5_50_tmp1[7])
         );
  DFFRHQX1 x5_50_tmp1_reg_6_ ( .D(x5[1]), .CK(clk), .RN(rstn), .Q(
        x5_50_tmp1[6]) );
  DFFRHQX1 x7_50_tmp1_reg_8_ ( .D(n3), .CK(clk), .RN(rstn), .Q(x7_50_tmp1[8])
         );
  DFFRHQX1 x7_50_tmp1_reg_7_ ( .D(n2), .CK(clk), .RN(rstn), .Q(x7_50_tmp1[7])
         );
  DFFRHQX1 x7_50_tmp1_reg_6_ ( .D(x7[1]), .CK(clk), .RN(rstn), .Q(
        x7_50_tmp1[6]) );
  DFFRHQX1 x4_18_tmp1_reg_7_ ( .D(n69), .CK(clk), .RN(rstn), .Q(x4_18_tmp1[7])
         );
  DFFRHQX1 x4_18_tmp1_reg_6_ ( .D(n68), .CK(clk), .RN(rstn), .Q(x4_18_tmp1[6])
         );
  DFFRHQX1 x4_18_tmp1_reg_5_ ( .D(x4[1]), .CK(clk), .RN(rstn), .Q(
        x4_18_tmp1[5]) );
  DFFRHQX1 x5_18_tmp1_reg_7_ ( .D(n56), .CK(clk), .RN(rstn), .Q(x5_18_tmp1[7])
         );
  DFFRHQX1 x5_18_tmp1_reg_6_ ( .D(n55), .CK(clk), .RN(rstn), .Q(x5_18_tmp1[6])
         );
  DFFRHQX1 x5_18_tmp1_reg_5_ ( .D(x5[1]), .CK(clk), .RN(rstn), .Q(
        x5_18_tmp1[5]) );
  DFFRHQX1 x6_18_tmp1_reg_7_ ( .D(n43), .CK(clk), .RN(rstn), .Q(x6_18_tmp1[7])
         );
  DFFRHQX1 x6_18_tmp1_reg_6_ ( .D(n42), .CK(clk), .RN(rstn), .Q(x6_18_tmp1[6])
         );
  DFFRHQX1 x6_18_tmp1_reg_5_ ( .D(x6[1]), .CK(clk), .RN(rstn), .Q(
        x6_18_tmp1[5]) );
  DFFRHQX1 x7_18_tmp1_reg_7_ ( .D(n3), .CK(clk), .RN(rstn), .Q(x7_18_tmp1[7])
         );
  DFFRHQX1 x7_18_tmp1_reg_6_ ( .D(n2), .CK(clk), .RN(rstn), .Q(x7_18_tmp1[6])
         );
  DFFRHQX1 x7_18_tmp1_reg_5_ ( .D(x7[1]), .CK(clk), .RN(rstn), .Q(
        x7_18_tmp1[5]) );
  DFFRHQX1 x5_18_reg_12_ ( .D(N526), .CK(clk), .RN(rstn), .Q(x5_18[12]) );
  DFFRHQX1 x5_18_reg_11_ ( .D(N525), .CK(clk), .RN(rstn), .Q(x5_18[11]) );
  DFFRHQX1 x5_18_reg_10_ ( .D(N524), .CK(clk), .RN(rstn), .Q(x5_18[10]) );
  DFFRHQX1 x5_18_reg_9_ ( .D(N523), .CK(clk), .RN(rstn), .Q(x5_18[9]) );
  DFFRHQX1 x5_18_reg_8_ ( .D(N522), .CK(clk), .RN(rstn), .Q(x5_18[8]) );
  DFFRHQX1 x6_18_reg_10_ ( .D(N613), .CK(clk), .RN(rstn), .Q(x6_18[10]) );
  DFFRHQX1 x6_18_reg_9_ ( .D(N612), .CK(clk), .RN(rstn), .Q(x6_18[9]) );
  DFFRHQX1 x6_18_reg_8_ ( .D(N611), .CK(clk), .RN(rstn), .Q(x6_18[8]) );
  DFFRHQX1 x6_18_reg_7_ ( .D(N610), .CK(clk), .RN(rstn), .Q(x6_18[7]) );
  DFFRHQX1 x4_18_reg_10_ ( .D(N435), .CK(clk), .RN(rstn), .Q(x4_18[10]) );
  DFFRHQX1 x4_18_reg_9_ ( .D(N434), .CK(clk), .RN(rstn), .Q(x4_18[9]) );
  DFFRHQX1 x4_18_reg_8_ ( .D(N433), .CK(clk), .RN(rstn), .Q(x4_18[8]) );
  DFFRHQX1 x4_18_reg_7_ ( .D(N432), .CK(clk), .RN(rstn), .Q(x4_18[7]) );
  DFFRHQX1 x4_89_tmp1_reg_9_ ( .D(N26), .CK(clk), .RN(rstn), .Q(x4_89_tmp1[9])
         );
  DFFRHQX1 x4_89_tmp1_reg_8_ ( .D(N25), .CK(clk), .RN(rstn), .Q(x4_89_tmp1[8])
         );
  DFFRHQX1 x4_89_tmp1_reg_7_ ( .D(N24), .CK(clk), .RN(rstn), .Q(x4_89_tmp1[7])
         );
  DFFRHQX1 x4_89_tmp1_reg_6_ ( .D(N23), .CK(clk), .RN(rstn), .Q(x4_89_tmp1[6])
         );
  DFFRHQX1 x4_89_reg_10_ ( .D(N367), .CK(clk), .RN(rstn), .Q(x4_89[10]) );
  DFFRHQX1 x4_89_reg_9_ ( .D(N366), .CK(clk), .RN(rstn), .Q(x4_89[9]) );
  DFFRHQX1 x4_89_reg_8_ ( .D(N365), .CK(clk), .RN(rstn), .Q(x4_89[8]) );
  DFFRHQX1 x4_89_reg_7_ ( .D(N364), .CK(clk), .RN(rstn), .Q(x4_89[7]) );
  DFFRHQX1 x4_75_reg_10_ ( .D(N390), .CK(clk), .RN(rstn), .Q(x4_75[10]) );
  DFFRHQX1 x4_75_reg_9_ ( .D(N389), .CK(clk), .RN(rstn), .Q(x4_75[9]) );
  DFFRHQX1 x4_75_reg_8_ ( .D(N388), .CK(clk), .RN(rstn), .Q(x4_75[8]) );
  DFFRHQX1 x4_75_reg_7_ ( .D(N387), .CK(clk), .RN(rstn), .Q(x4_75[7]) );
  DFFRHQX1 x5_75_reg_10_ ( .D(N479), .CK(clk), .RN(rstn), .Q(x5_75[10]) );
  DFFRHQX1 x5_75_reg_9_ ( .D(N478), .CK(clk), .RN(rstn), .Q(x5_75[9]) );
  DFFRHQX1 x5_75_reg_8_ ( .D(N477), .CK(clk), .RN(rstn), .Q(x5_75[8]) );
  DFFRHQX1 x5_75_reg_7_ ( .D(N476), .CK(clk), .RN(rstn), .Q(x5_75[7]) );
  DFFRHQX1 x6_75_reg_10_ ( .D(N568), .CK(clk), .RN(rstn), .Q(x6_75[10]) );
  DFFRHQX1 x6_75_reg_9_ ( .D(N567), .CK(clk), .RN(rstn), .Q(x6_75[9]) );
  DFFRHQX1 x6_75_reg_8_ ( .D(N566), .CK(clk), .RN(rstn), .Q(x6_75[8]) );
  DFFRHQX1 x6_75_reg_7_ ( .D(N565), .CK(clk), .RN(rstn), .Q(x6_75[7]) );
  DFFRHQX1 x4_50_reg_10_ ( .D(N413), .CK(clk), .RN(rstn), .Q(x4_50[10]) );
  DFFRHQX1 x4_50_reg_9_ ( .D(N412), .CK(clk), .RN(rstn), .Q(x4_50[9]) );
  DFFRHQX1 x4_50_reg_8_ ( .D(N411), .CK(clk), .RN(rstn), .Q(x4_50[8]) );
  DFFRHQX1 x4_50_reg_7_ ( .D(N410), .CK(clk), .RN(rstn), .Q(x4_50[7]) );
  DFFRHQX1 x5_tmp1_reg_11_ ( .D(N890), .CK(clk), .RN(rstn), .Q(x5_tmp1[11]) );
  DFFRHQX1 x5_tmp1_reg_10_ ( .D(N889), .CK(clk), .RN(rstn), .Q(x5_tmp1[10]) );
  DFFRHQX1 x5_tmp1_reg_9_ ( .D(N888), .CK(clk), .RN(rstn), .Q(x5_tmp1[9]) );
  DFFRHQX1 x5_tmp1_reg_8_ ( .D(N887), .CK(clk), .RN(rstn), .Q(x5_tmp1[8]) );
  DFFRHQX1 x6_tmp1_reg_11_ ( .D(N1056), .CK(clk), .RN(rstn), .Q(x6_tmp1[11])
         );
  DFFRHQX1 x6_tmp1_reg_10_ ( .D(N1055), .CK(clk), .RN(rstn), .Q(x6_tmp1[10])
         );
  DFFRHQX1 x6_tmp1_reg_9_ ( .D(N1054), .CK(clk), .RN(rstn), .Q(x6_tmp1[9]) );
  DFFRHQX1 x6_tmp1_reg_8_ ( .D(N1053), .CK(clk), .RN(rstn), .Q(x6_tmp1[8]) );
  DFFRHQX1 x7_tmp1_reg_11_ ( .D(N1153), .CK(clk), .RN(rstn), .Q(x7_tmp1[11])
         );
  DFFRHQX1 x7_tmp1_reg_10_ ( .D(N1152), .CK(clk), .RN(rstn), .Q(x7_tmp1[10])
         );
  DFFRHQX1 x7_tmp1_reg_9_ ( .D(N1151), .CK(clk), .RN(rstn), .Q(x7_tmp1[9]) );
  DFFRHQX1 x7_tmp1_reg_8_ ( .D(N1150), .CK(clk), .RN(rstn), .Q(x7_tmp1[8]) );
  DFFRHQX1 x4_tmp1_reg_11_ ( .D(N771), .CK(clk), .RN(rstn), .Q(x4_tmp1[11]) );
  DFFRHQX1 x4_tmp1_reg_10_ ( .D(N770), .CK(clk), .RN(rstn), .Q(x4_tmp1[10]) );
  DFFRHQX1 x4_tmp1_reg_9_ ( .D(N769), .CK(clk), .RN(rstn), .Q(x4_tmp1[9]) );
  DFFRHQX1 x4_tmp1_reg_8_ ( .D(N768), .CK(clk), .RN(rstn), .Q(x4_tmp1[8]) );
  DFFRHQX1 y7_tmp_reg_17_ ( .D(N1618), .CK(clk), .RN(rstn), .Q(y7_tmp[17]) );
  DFFRHQX1 y0_tmp_reg_18_ ( .D(N1233), .CK(clk), .RN(rstn), .Q(y0_tmp[18]) );
  DFFRHQX1 y0_tmp_reg_17_ ( .D(N1232), .CK(clk), .RN(rstn), .Q(y0_tmp[17]) );
  DFFRHQX1 y1_tmp_reg_18_ ( .D(N1259), .CK(clk), .RN(rstn), .Q(y1_tmp[18]) );
  DFFRHQX1 y1_tmp_reg_17_ ( .D(N1258), .CK(clk), .RN(rstn), .Q(y1_tmp[17]) );
  DFFRHQX1 y2_tmp_reg_18_ ( .D(N1285), .CK(clk), .RN(rstn), .Q(y2_tmp[18]) );
  DFFRHQX1 y2_tmp_reg_17_ ( .D(N1284), .CK(clk), .RN(rstn), .Q(y2_tmp[17]) );
  DFFRHQX1 y3_tmp_reg_18_ ( .D(N1311), .CK(clk), .RN(rstn), .Q(y3_tmp[18]) );
  DFFRHQX1 y3_tmp_reg_17_ ( .D(N1310), .CK(clk), .RN(rstn), .Q(y3_tmp[17]) );
  DFFRHQX1 idct8_ready_reg ( .D(start), .CK(clk), .RN(rstn), .Q(idct8_ready)
         );
  DFFRHQX1 x7_50_reg_11_ ( .D(N681), .CK(clk), .RN(rstn), .Q(x7_50[11]) );
  DFFRHQX1 x7_50_reg_10_ ( .D(N680), .CK(clk), .RN(rstn), .Q(x7_50[10]) );
  DFFRHQX1 x7_50_reg_9_ ( .D(N679), .CK(clk), .RN(rstn), .Q(x7_50[9]) );
  DFFRHQX1 x7_50_reg_8_ ( .D(N678), .CK(clk), .RN(rstn), .Q(x7_50[8]) );
  DFFRHQX1 x7_50_reg_7_ ( .D(N677), .CK(clk), .RN(rstn), .Q(x7_50[7]) );
  DFFRHQX1 x5_89_reg_11_ ( .D(N457), .CK(clk), .RN(rstn), .Q(x5_89[11]) );
  DFFRHQX1 x5_89_reg_10_ ( .D(N456), .CK(clk), .RN(rstn), .Q(x5_89[10]) );
  DFFRHQX1 x5_89_reg_9_ ( .D(N455), .CK(clk), .RN(rstn), .Q(x5_89[9]) );
  DFFRHQX1 x5_89_reg_8_ ( .D(N454), .CK(clk), .RN(rstn), .Q(x5_89[8]) );
  DFFRHQX1 x5_89_reg_7_ ( .D(N453), .CK(clk), .RN(rstn), .Q(x5_89[7]) );
  DFFRHQX1 x7_89_reg_11_ ( .D(N635), .CK(clk), .RN(rstn), .Q(x7_89[11]) );
  DFFRHQX1 x7_89_reg_10_ ( .D(N634), .CK(clk), .RN(rstn), .Q(x7_89[10]) );
  DFFRHQX1 x7_89_reg_9_ ( .D(N633), .CK(clk), .RN(rstn), .Q(x7_89[9]) );
  DFFRHQX1 x7_89_reg_8_ ( .D(N632), .CK(clk), .RN(rstn), .Q(x7_89[8]) );
  DFFRHQX1 x7_89_reg_7_ ( .D(N631), .CK(clk), .RN(rstn), .Q(x7_89[7]) );
  DFFRHQX1 x5_50_reg_11_ ( .D(N503), .CK(clk), .RN(rstn), .Q(x5_50[11]) );
  DFFRHQX1 x5_50_reg_10_ ( .D(N502), .CK(clk), .RN(rstn), .Q(x5_50[10]) );
  DFFRHQX1 x5_50_reg_9_ ( .D(N501), .CK(clk), .RN(rstn), .Q(x5_50[9]) );
  DFFRHQX1 x5_50_reg_8_ ( .D(N500), .CK(clk), .RN(rstn), .Q(x5_50[8]) );
  DFFRHQX1 x5_50_reg_7_ ( .D(N499), .CK(clk), .RN(rstn), .Q(x5_50[7]) );
  DFFRHQX1 y6_tmp_reg_16_ ( .D(N1540), .CK(clk), .RN(rstn), .Q(y6_tmp[16]) );
  DFFRHQX1 y6_tmp_reg_15_ ( .D(N1539), .CK(clk), .RN(rstn), .Q(y6_tmp[15]) );
  DFFRHQX1 y6_tmp_reg_14_ ( .D(N1538), .CK(clk), .RN(rstn), .Q(y6_tmp[14]) );
  DFFRHQX1 y6_tmp_reg_13_ ( .D(N1537), .CK(clk), .RN(rstn), .Q(y6_tmp[13]) );
  DFFRHQX1 y7_tmp_reg_16_ ( .D(N1617), .CK(clk), .RN(rstn), .Q(y7_tmp[16]) );
  DFFRHQX1 y7_tmp_reg_15_ ( .D(N1616), .CK(clk), .RN(rstn), .Q(y7_tmp[15]) );
  DFFRHQX1 y7_tmp_reg_14_ ( .D(N1615), .CK(clk), .RN(rstn), .Q(y7_tmp[14]) );
  DFFRHQX1 y7_tmp_reg_13_ ( .D(N1614), .CK(clk), .RN(rstn), .Q(y7_tmp[13]) );
  DFFRHQX1 y0_tmp_reg_16_ ( .D(N1231), .CK(clk), .RN(rstn), .Q(y0_tmp[16]) );
  DFFRHQX1 y0_tmp_reg_15_ ( .D(N1230), .CK(clk), .RN(rstn), .Q(y0_tmp[15]) );
  DFFRHQX1 y1_tmp_reg_16_ ( .D(N1257), .CK(clk), .RN(rstn), .Q(y1_tmp[16]) );
  DFFRHQX1 y1_tmp_reg_15_ ( .D(N1256), .CK(clk), .RN(rstn), .Q(y1_tmp[15]) );
  DFFRHQX1 y2_tmp_reg_16_ ( .D(N1283), .CK(clk), .RN(rstn), .Q(y2_tmp[16]) );
  DFFRHQX1 y2_tmp_reg_15_ ( .D(N1282), .CK(clk), .RN(rstn), .Q(y2_tmp[15]) );
  DFFRHQX1 y3_tmp_reg_16_ ( .D(N1309), .CK(clk), .RN(rstn), .Q(y3_tmp[16]) );
  DFFRHQX1 y3_tmp_reg_15_ ( .D(N1308), .CK(clk), .RN(rstn), .Q(y3_tmp[15]) );
  DFFRHQX1 y4_tmp_reg_16_ ( .D(N1386), .CK(clk), .RN(rstn), .Q(y4_tmp[16]) );
  DFFRHQX1 y4_tmp_reg_15_ ( .D(N1385), .CK(clk), .RN(rstn), .Q(y4_tmp[15]) );
  DFFRHQX1 y4_tmp_reg_14_ ( .D(N1384), .CK(clk), .RN(rstn), .Q(y4_tmp[14]) );
  DFFRHQX1 y4_tmp_reg_13_ ( .D(N1383), .CK(clk), .RN(rstn), .Q(y4_tmp[13]) );
  DFFRHQX1 y5_tmp_reg_16_ ( .D(N1463), .CK(clk), .RN(rstn), .Q(y5_tmp[16]) );
  DFFRHQX1 y5_tmp_reg_15_ ( .D(N1462), .CK(clk), .RN(rstn), .Q(y5_tmp[15]) );
  DFFRHQX1 y5_tmp_reg_14_ ( .D(N1461), .CK(clk), .RN(rstn), .Q(y5_tmp[14]) );
  DFFRHQX1 y5_tmp_reg_13_ ( .D(N1460), .CK(clk), .RN(rstn), .Q(y5_tmp[13]) );
  DFFRHQX1 x6_89_tmp2_reg_9_ ( .D(N219), .CK(clk), .RN(rstn), .Q(x6_89_tmp2[9]) );
  DFFRHQX1 x6_89_tmp2_reg_8_ ( .D(N218), .CK(clk), .RN(rstn), .Q(x6_89_tmp2[8]) );
  DFFRHQX1 x6_89_tmp2_reg_7_ ( .D(N217), .CK(clk), .RN(rstn), .Q(x6_89_tmp2[7]) );
  DFFRHQX1 x6_89_tmp2_reg_6_ ( .D(N216), .CK(clk), .RN(rstn), .Q(x6_89_tmp2[6]) );
  DFFRHQX1 x5_89_tmp2_reg_9_ ( .D(N134), .CK(clk), .RN(rstn), .Q(x5_89_tmp2[9]) );
  DFFRHQX1 x5_89_tmp2_reg_8_ ( .D(N133), .CK(clk), .RN(rstn), .Q(x5_89_tmp2[8]) );
  DFFRHQX1 x5_89_tmp2_reg_7_ ( .D(N132), .CK(clk), .RN(rstn), .Q(x5_89_tmp2[7]) );
  DFFRHQX1 x5_89_tmp2_reg_6_ ( .D(N131), .CK(clk), .RN(rstn), .Q(x5_89_tmp2[6]) );
  DFFRHQX1 x4_89_tmp2_reg_9_ ( .D(N49), .CK(clk), .RN(rstn), .Q(x4_89_tmp2[9])
         );
  DFFRHQX1 x4_89_tmp2_reg_8_ ( .D(N48), .CK(clk), .RN(rstn), .Q(x4_89_tmp2[8])
         );
  DFFRHQX1 x4_89_tmp2_reg_7_ ( .D(N47), .CK(clk), .RN(rstn), .Q(x4_89_tmp2[7])
         );
  DFFRHQX1 x4_89_tmp2_reg_6_ ( .D(N46), .CK(clk), .RN(rstn), .Q(x4_89_tmp2[6])
         );
  DFFRHQX1 x7_89_tmp2_reg_9_ ( .D(N304), .CK(clk), .RN(rstn), .Q(x7_89_tmp2[9]) );
  DFFRHQX1 x7_89_tmp2_reg_8_ ( .D(N303), .CK(clk), .RN(rstn), .Q(x7_89_tmp2[8]) );
  DFFRHQX1 x7_89_tmp2_reg_7_ ( .D(N302), .CK(clk), .RN(rstn), .Q(x7_89_tmp2[7]) );
  DFFRHQX1 x7_89_tmp2_reg_6_ ( .D(N301), .CK(clk), .RN(rstn), .Q(x7_89_tmp2[6]) );
  DFFRHQX1 x4_75_tmp2_reg_9_ ( .D(N70), .CK(clk), .RN(rstn), .Q(x4_75_tmp2[9])
         );
  DFFRHQX1 x4_75_tmp2_reg_8_ ( .D(N69), .CK(clk), .RN(rstn), .Q(x4_75_tmp2[8])
         );
  DFFRHQX1 x4_75_tmp2_reg_7_ ( .D(N68), .CK(clk), .RN(rstn), .Q(x4_75_tmp2[7])
         );
  DFFRHQX1 x4_75_tmp2_reg_6_ ( .D(N67), .CK(clk), .RN(rstn), .Q(x4_75_tmp2[6])
         );
  DFFRHQX1 x5_75_tmp2_reg_9_ ( .D(N155), .CK(clk), .RN(rstn), .Q(x5_75_tmp2[9]) );
  DFFRHQX1 x5_75_tmp2_reg_8_ ( .D(N154), .CK(clk), .RN(rstn), .Q(x5_75_tmp2[8]) );
  DFFRHQX1 x5_75_tmp2_reg_7_ ( .D(N153), .CK(clk), .RN(rstn), .Q(x5_75_tmp2[7]) );
  DFFRHQX1 x5_75_tmp2_reg_6_ ( .D(N152), .CK(clk), .RN(rstn), .Q(x5_75_tmp2[6]) );
  DFFRHQX1 x6_75_tmp2_reg_9_ ( .D(N240), .CK(clk), .RN(rstn), .Q(x6_75_tmp2[9]) );
  DFFRHQX1 x6_75_tmp2_reg_8_ ( .D(N239), .CK(clk), .RN(rstn), .Q(x6_75_tmp2[8]) );
  DFFRHQX1 x6_75_tmp2_reg_7_ ( .D(N238), .CK(clk), .RN(rstn), .Q(x6_75_tmp2[7]) );
  DFFRHQX1 x6_75_tmp2_reg_6_ ( .D(N237), .CK(clk), .RN(rstn), .Q(x6_75_tmp2[6]) );
  DFFRHQX1 x7_75_tmp2_reg_9_ ( .D(N325), .CK(clk), .RN(rstn), .Q(x7_75_tmp2[9]) );
  DFFRHQX1 x7_75_tmp2_reg_8_ ( .D(N324), .CK(clk), .RN(rstn), .Q(x7_75_tmp2[8]) );
  DFFRHQX1 x7_75_tmp2_reg_7_ ( .D(N323), .CK(clk), .RN(rstn), .Q(x7_75_tmp2[7]) );
  DFFRHQX1 x7_75_tmp2_reg_6_ ( .D(N322), .CK(clk), .RN(rstn), .Q(x7_75_tmp2[6]) );
  DFFRHQX1 x4_50_tmp2_reg_8_ ( .D(N89), .CK(clk), .RN(rstn), .Q(x4_50_tmp2[8])
         );
  DFFRHQX1 x4_50_tmp2_reg_7_ ( .D(N88), .CK(clk), .RN(rstn), .Q(x4_50_tmp2[7])
         );
  DFFRHQX1 x4_50_tmp2_reg_6_ ( .D(N87), .CK(clk), .RN(rstn), .Q(x4_50_tmp2[6])
         );
  DFFRHQX1 x6_50_tmp2_reg_8_ ( .D(N259), .CK(clk), .RN(rstn), .Q(x6_50_tmp2[8]) );
  DFFRHQX1 x6_50_tmp2_reg_7_ ( .D(N258), .CK(clk), .RN(rstn), .Q(x6_50_tmp2[7]) );
  DFFRHQX1 x6_50_tmp2_reg_6_ ( .D(N257), .CK(clk), .RN(rstn), .Q(x6_50_tmp2[6]) );
  DFFRHQX1 x6_50_reg_7_ ( .D(N588), .CK(clk), .RN(rstn), .Q(x6_50[7]) );
  DFFRHQX1 x6_50_reg_8_ ( .D(N589), .CK(clk), .RN(rstn), .Q(x6_50[8]) );
  DFFRHQX1 x6_50_reg_9_ ( .D(N590), .CK(clk), .RN(rstn), .Q(x6_50[9]) );
  DFFRHQX1 x6_50_reg_10_ ( .D(N591), .CK(clk), .RN(rstn), .Q(x6_50[10]) );
  DFFRHQX1 x5_50_tmp2_reg_8_ ( .D(N174), .CK(clk), .RN(rstn), .Q(x5_50_tmp2[8]) );
  DFFRHQX1 x5_50_tmp2_reg_7_ ( .D(N173), .CK(clk), .RN(rstn), .Q(x5_50_tmp2[7]) );
  DFFRHQX1 x5_50_tmp2_reg_6_ ( .D(N172), .CK(clk), .RN(rstn), .Q(x5_50_tmp2[6]) );
  DFFRHQX1 x7_50_tmp2_reg_8_ ( .D(N344), .CK(clk), .RN(rstn), .Q(x7_50_tmp2[8]) );
  DFFRHQX1 x7_50_tmp2_reg_7_ ( .D(N343), .CK(clk), .RN(rstn), .Q(x7_50_tmp2[7]) );
  DFFRHQX1 x7_50_tmp2_reg_6_ ( .D(N342), .CK(clk), .RN(rstn), .Q(x7_50_tmp2[6]) );
  DFFRHQX1 x4_18_tmp2_reg_7_ ( .D(n72), .CK(clk), .RN(rstn), .Q(x4_18_tmp2[7])
         );
  DFFRHQX1 x4_18_tmp2_reg_6_ ( .D(n71), .CK(clk), .RN(rstn), .Q(x4_18_tmp2[6])
         );
  DFFRHQX1 x4_18_tmp2_reg_5_ ( .D(n70), .CK(clk), .RN(rstn), .Q(x4_18_tmp2[5])
         );
  DFFRHQX1 x6_18_tmp2_reg_7_ ( .D(n46), .CK(clk), .RN(rstn), .Q(x6_18_tmp2[7])
         );
  DFFRHQX1 x6_18_tmp2_reg_6_ ( .D(n45), .CK(clk), .RN(rstn), .Q(x6_18_tmp2[6])
         );
  DFFRHQX1 x6_18_tmp2_reg_5_ ( .D(n44), .CK(clk), .RN(rstn), .Q(x6_18_tmp2[5])
         );
  DFFRHQX1 x5_18_tmp2_reg_7_ ( .D(n59), .CK(clk), .RN(rstn), .Q(x5_18_tmp2[7])
         );
  DFFRHQX1 x5_18_tmp2_reg_6_ ( .D(n58), .CK(clk), .RN(rstn), .Q(x5_18_tmp2[6])
         );
  DFFRHQX1 x5_18_tmp2_reg_5_ ( .D(n57), .CK(clk), .RN(rstn), .Q(x5_18_tmp2[5])
         );
  DFFRHQX1 x7_18_tmp2_reg_7_ ( .D(n6), .CK(clk), .RN(rstn), .Q(x7_18_tmp2[7])
         );
  DFFRHQX1 x7_18_tmp2_reg_6_ ( .D(n5), .CK(clk), .RN(rstn), .Q(x7_18_tmp2[6])
         );
  DFFRHQX1 x7_18_tmp2_reg_5_ ( .D(n4), .CK(clk), .RN(rstn), .Q(x7_18_tmp2[5])
         );
  DFFRHQX1 x7_18_reg_10_ ( .D(N702), .CK(clk), .RN(rstn), .Q(x7_18[10]) );
  DFFRHQX1 x7_18_reg_9_ ( .D(N701), .CK(clk), .RN(rstn), .Q(x7_18[9]) );
  DFFRHQX1 x7_18_reg_8_ ( .D(N700), .CK(clk), .RN(rstn), .Q(x7_18[8]) );
  DFFRHQX1 x7_18_reg_7_ ( .D(N699), .CK(clk), .RN(rstn), .Q(x7_18[7]) );
  DFFRHQX1 x6_89_reg_11_ ( .D(N546), .CK(clk), .RN(rstn), .Q(x6_89[11]) );
  DFFRHQX1 x6_89_reg_10_ ( .D(N545), .CK(clk), .RN(rstn), .Q(x6_89[10]) );
  DFFRHQX1 x6_89_reg_9_ ( .D(N544), .CK(clk), .RN(rstn), .Q(x6_89[9]) );
  DFFRHQX1 x6_89_reg_8_ ( .D(N543), .CK(clk), .RN(rstn), .Q(x6_89[8]) );
  DFFRHQX1 x7_75_reg_10_ ( .D(N657), .CK(clk), .RN(rstn), .Q(x7_75[10]) );
  DFFRHQX1 x7_75_reg_9_ ( .D(N656), .CK(clk), .RN(rstn), .Q(x7_75[9]) );
  DFFRHQX1 x7_75_reg_8_ ( .D(N655), .CK(clk), .RN(rstn), .Q(x7_75[8]) );
  DFFRHQX1 x7_75_reg_7_ ( .D(N654), .CK(clk), .RN(rstn), .Q(x7_75[7]) );
  DFFRHQX1 x4_tmp2_reg_11_ ( .D(N841), .CK(clk), .RN(rstn), .Q(x4_tmp2[11]) );
  DFFRHQX1 x4_tmp2_reg_10_ ( .D(N840), .CK(clk), .RN(rstn), .Q(x4_tmp2[10]) );
  DFFRHQX1 x4_tmp2_reg_9_ ( .D(N839), .CK(clk), .RN(rstn), .Q(x4_tmp2[9]) );
  DFFRHQX1 x4_tmp2_reg_8_ ( .D(N838), .CK(clk), .RN(rstn), .Q(x4_tmp2[8]) );
  DFFRHQX1 x5_tmp2_reg_11_ ( .D(N961), .CK(clk), .RN(rstn), .Q(x5_tmp2[11]) );
  DFFRHQX1 x5_tmp2_reg_10_ ( .D(N960), .CK(clk), .RN(rstn), .Q(x5_tmp2[10]) );
  DFFRHQX1 x5_tmp2_reg_9_ ( .D(N959), .CK(clk), .RN(rstn), .Q(x5_tmp2[9]) );
  DFFRHQX1 x5_tmp2_reg_8_ ( .D(N958), .CK(clk), .RN(rstn), .Q(x5_tmp2[8]) );
  DFFRHQX1 x6_tmp2_reg_11_ ( .D(N1104), .CK(clk), .RN(rstn), .Q(x6_tmp2[11])
         );
  DFFRHQX1 x6_tmp2_reg_10_ ( .D(N1103), .CK(clk), .RN(rstn), .Q(x6_tmp2[10])
         );
  DFFRHQX1 x6_tmp2_reg_9_ ( .D(N1102), .CK(clk), .RN(rstn), .Q(x6_tmp2[9]) );
  DFFRHQX1 x6_tmp2_reg_8_ ( .D(N1101), .CK(clk), .RN(rstn), .Q(x6_tmp2[8]) );
  DFFRHQX1 x7_tmp2_reg_11_ ( .D(N1177), .CK(clk), .RN(rstn), .Q(x7_tmp2[11])
         );
  DFFRHQX1 x7_tmp2_reg_10_ ( .D(N1176), .CK(clk), .RN(rstn), .Q(x7_tmp2[10])
         );
  DFFRHQX1 x7_tmp2_reg_9_ ( .D(N1175), .CK(clk), .RN(rstn), .Q(x7_tmp2[9]) );
  DFFRHQX1 x7_tmp2_reg_8_ ( .D(N1174), .CK(clk), .RN(rstn), .Q(x7_tmp2[8]) );
  DFFRHQX1 x4_50_tmp2_reg_5_ ( .D(N86), .CK(clk), .RN(rstn), .Q(x4_50_tmp2[5])
         );
  DFFRHQX1 x6_50_tmp2_reg_5_ ( .D(N256), .CK(clk), .RN(rstn), .Q(x6_50_tmp2[5]) );
  DFFRHQX1 x5_50_tmp2_reg_5_ ( .D(N171), .CK(clk), .RN(rstn), .Q(x5_50_tmp2[5]) );
  DFFRHQX1 x7_50_tmp2_reg_5_ ( .D(N341), .CK(clk), .RN(rstn), .Q(x7_50_tmp2[5]) );
  DFFRHQX1 x4_18_tmp2_reg_4_ ( .D(n69), .CK(clk), .RN(rstn), .Q(x4_18_tmp2[4])
         );
  DFFRHQX1 x6_18_tmp2_reg_4_ ( .D(n43), .CK(clk), .RN(rstn), .Q(x6_18_tmp2[4])
         );
  DFFRHQX1 x5_18_tmp2_reg_4_ ( .D(n56), .CK(clk), .RN(rstn), .Q(x5_18_tmp2[4])
         );
  DFFRHQX1 x7_18_tmp2_reg_4_ ( .D(n3), .CK(clk), .RN(rstn), .Q(x7_18_tmp2[4])
         );
  DFFRHQX1 x4_50_tmp1_reg_5_ ( .D(x4[0]), .CK(clk), .RN(rstn), .Q(
        x4_50_tmp1[5]) );
  DFFRHQX1 x6_50_tmp1_reg_5_ ( .D(x6[0]), .CK(clk), .RN(rstn), .Q(
        x6_50_tmp1[5]) );
  DFFRHQX1 x5_50_tmp1_reg_5_ ( .D(x5[0]), .CK(clk), .RN(rstn), .Q(
        x5_50_tmp1[5]) );
  DFFRHQX1 x7_50_tmp1_reg_5_ ( .D(x7[0]), .CK(clk), .RN(rstn), .Q(
        x7_50_tmp1[5]) );
  DFFRHQX1 x4_18_tmp1_reg_4_ ( .D(x4[0]), .CK(clk), .RN(rstn), .Q(
        x4_18_tmp1[4]) );
  DFFRHQX1 x5_18_tmp1_reg_4_ ( .D(x5[0]), .CK(clk), .RN(rstn), .Q(
        x5_18_tmp1[4]) );
  DFFRHQX1 x6_18_tmp1_reg_4_ ( .D(x6[0]), .CK(clk), .RN(rstn), .Q(
        x6_18_tmp1[4]) );
  DFFRHQX1 x7_18_tmp1_reg_4_ ( .D(x7[0]), .CK(clk), .RN(rstn), .Q(
        x7_18_tmp1[4]) );
  DFFRHQX1 x7_tmp_reg_10_ ( .D(N1200), .CK(clk), .RN(rstn), .Q(x7_tmp[10]) );
  DFFRHQX1 x7_tmp_reg_11_ ( .D(N1201), .CK(clk), .RN(rstn), .Q(x7_tmp[11]) );
  DFFRHQX1 x7_tmp_reg_12_ ( .D(N1202), .CK(clk), .RN(rstn), .Q(x7_tmp[12]) );
  DFFRHQX1 x7_tmp_reg_13_ ( .D(N1203), .CK(clk), .RN(rstn), .Q(x7_tmp[13]) );
  DFFRHQX1 x5_tmp_reg_13_ ( .D(N987), .CK(clk), .RN(rstn), .Q(x5_tmp[13]) );
  DFFRHQX1 x5_tmp_reg_12_ ( .D(N986), .CK(clk), .RN(rstn), .Q(x5_tmp[12]) );
  DFFRHQX1 x5_tmp_reg_11_ ( .D(N985), .CK(clk), .RN(rstn), .Q(x5_tmp[11]) );
  DFFRHQX1 x5_tmp_reg_10_ ( .D(N984), .CK(clk), .RN(rstn), .Q(x5_tmp[10]) );
  DFFRHQX1 x6_tmp_reg_13_ ( .D(N1130), .CK(clk), .RN(rstn), .Q(x6_tmp[13]) );
  DFFRHQX1 x6_tmp_reg_12_ ( .D(N1129), .CK(clk), .RN(rstn), .Q(x6_tmp[12]) );
  DFFRHQX1 x6_tmp_reg_11_ ( .D(N1128), .CK(clk), .RN(rstn), .Q(x6_tmp[11]) );
  DFFRHQX1 x6_tmp_reg_10_ ( .D(N1127), .CK(clk), .RN(rstn), .Q(x6_tmp[10]) );
  DFFRHQX1 x4_tmp_reg_10_ ( .D(N864), .CK(clk), .RN(rstn), .Q(x4_tmp[10]) );
  DFFRHQX1 x4_tmp_reg_11_ ( .D(N865), .CK(clk), .RN(rstn), .Q(x4_tmp[11]) );
  DFFRHQX1 x4_tmp_reg_12_ ( .D(N866), .CK(clk), .RN(rstn), .Q(x4_tmp[12]) );
  DFFRHQX1 x4_tmp_reg_13_ ( .D(N867), .CK(clk), .RN(rstn), .Q(x4_tmp[13]) );
  DFFRHQX1 x7_89_tmp1_reg_5_ ( .D(n5), .CK(clk), .RN(rstn), .Q(x7_89_tmp1[5])
         );
  DFFRHQX1 x7_89_tmp1_reg_4_ ( .D(n4), .CK(clk), .RN(rstn), .Q(x7_89_tmp1[4])
         );
  DFFRHQX1 x7_89_tmp1_reg_3_ ( .D(n3), .CK(clk), .RN(rstn), .Q(x7_89_tmp1[3])
         );
  DFFRHQX1 x7_89_tmp1_reg_2_ ( .D(n2), .CK(clk), .RN(rstn), .Q(x7_89_tmp1[2])
         );
  DFFRHQX1 x6_89_tmp1_reg_5_ ( .D(n45), .CK(clk), .RN(rstn), .Q(x6_89_tmp1[5])
         );
  DFFRHQX1 x6_89_tmp1_reg_4_ ( .D(n44), .CK(clk), .RN(rstn), .Q(x6_89_tmp1[4])
         );
  DFFRHQX1 x6_89_tmp1_reg_3_ ( .D(n43), .CK(clk), .RN(rstn), .Q(x6_89_tmp1[3])
         );
  DFFRHQX1 x6_89_tmp1_reg_2_ ( .D(n42), .CK(clk), .RN(rstn), .Q(x6_89_tmp1[2])
         );
  DFFRHQX1 x5_89_tmp1_reg_5_ ( .D(n58), .CK(clk), .RN(rstn), .Q(x5_89_tmp1[5])
         );
  DFFRHQX1 x5_89_tmp1_reg_4_ ( .D(n57), .CK(clk), .RN(rstn), .Q(x5_89_tmp1[4])
         );
  DFFRHQX1 x5_89_tmp1_reg_3_ ( .D(n56), .CK(clk), .RN(rstn), .Q(x5_89_tmp1[3])
         );
  DFFRHQX1 x5_89_tmp1_reg_2_ ( .D(n55), .CK(clk), .RN(rstn), .Q(x5_89_tmp1[2])
         );
  DFFRHQX1 x5_75_tmp1_reg_5_ ( .D(n58), .CK(clk), .RN(rstn), .Q(x5_75_tmp1[5])
         );
  DFFRHQX1 x5_75_tmp1_reg_4_ ( .D(n57), .CK(clk), .RN(rstn), .Q(x5_75_tmp1[4])
         );
  DFFRHQX1 x5_75_tmp1_reg_3_ ( .D(n56), .CK(clk), .RN(rstn), .Q(x5_75_tmp1[3])
         );
  DFFRHQX1 x5_75_tmp1_reg_2_ ( .D(n55), .CK(clk), .RN(rstn), .Q(x5_75_tmp1[2])
         );
  DFFRHQX1 x4_75_tmp1_reg_5_ ( .D(n71), .CK(clk), .RN(rstn), .Q(x4_75_tmp1[5])
         );
  DFFRHQX1 x4_75_tmp1_reg_4_ ( .D(n70), .CK(clk), .RN(rstn), .Q(x4_75_tmp1[4])
         );
  DFFRHQX1 x4_75_tmp1_reg_3_ ( .D(n69), .CK(clk), .RN(rstn), .Q(x4_75_tmp1[3])
         );
  DFFRHQX1 x4_75_tmp1_reg_2_ ( .D(n68), .CK(clk), .RN(rstn), .Q(x4_75_tmp1[2])
         );
  DFFRHQX1 x7_75_tmp1_reg_5_ ( .D(n5), .CK(clk), .RN(rstn), .Q(x7_75_tmp1[5])
         );
  DFFRHQX1 x7_75_tmp1_reg_4_ ( .D(n4), .CK(clk), .RN(rstn), .Q(x7_75_tmp1[4])
         );
  DFFRHQX1 x7_75_tmp1_reg_3_ ( .D(n3), .CK(clk), .RN(rstn), .Q(x7_75_tmp1[3])
         );
  DFFRHQX1 x7_75_tmp1_reg_2_ ( .D(n2), .CK(clk), .RN(rstn), .Q(x7_75_tmp1[2])
         );
  DFFRHQX1 x6_75_tmp1_reg_5_ ( .D(n45), .CK(clk), .RN(rstn), .Q(x6_75_tmp1[5])
         );
  DFFRHQX1 x6_75_tmp1_reg_4_ ( .D(n44), .CK(clk), .RN(rstn), .Q(x6_75_tmp1[4])
         );
  DFFRHQX1 x6_75_tmp1_reg_3_ ( .D(n43), .CK(clk), .RN(rstn), .Q(x6_75_tmp1[3])
         );
  DFFRHQX1 x6_75_tmp1_reg_2_ ( .D(n42), .CK(clk), .RN(rstn), .Q(x6_75_tmp1[2])
         );
  DFFRHQX1 x5_18_reg_7_ ( .D(N521), .CK(clk), .RN(rstn), .Q(x5_18[7]) );
  DFFRHQX1 x5_18_reg_6_ ( .D(N520), .CK(clk), .RN(rstn), .Q(x5_18[6]) );
  DFFRHQX1 x5_18_reg_5_ ( .D(N519), .CK(clk), .RN(rstn), .Q(x5_18[5]) );
  DFFRHQX1 x5_18_reg_4_ ( .D(N518), .CK(clk), .RN(rstn), .Q(x5_18[4]) );
  DFFRHQX1 x6_18_reg_6_ ( .D(N609), .CK(clk), .RN(rstn), .Q(x6_18[6]) );
  DFFRHQX1 x6_18_reg_5_ ( .D(N608), .CK(clk), .RN(rstn), .Q(x6_18[5]) );
  DFFRHQX1 x6_18_reg_4_ ( .D(N607), .CK(clk), .RN(rstn), .Q(x6_18[4]) );
  DFFRHQX1 x6_18_reg_3_ ( .D(N606), .CK(clk), .RN(rstn), .Q(x6_18[3]) );
  DFFRHQX1 x4_18_reg_6_ ( .D(N431), .CK(clk), .RN(rstn), .Q(x4_18[6]) );
  DFFRHQX1 x4_18_reg_5_ ( .D(N430), .CK(clk), .RN(rstn), .Q(x4_18[5]) );
  DFFRHQX1 x4_18_reg_4_ ( .D(N429), .CK(clk), .RN(rstn), .Q(x4_18[4]) );
  DFFRHQX1 x4_18_reg_3_ ( .D(N428), .CK(clk), .RN(rstn), .Q(x4_18[3]) );
  DFFRHQX1 x4_89_tmp1_reg_5_ ( .D(n71), .CK(clk), .RN(rstn), .Q(x4_89_tmp1[5])
         );
  DFFRHQX1 x4_89_tmp1_reg_4_ ( .D(n70), .CK(clk), .RN(rstn), .Q(x4_89_tmp1[4])
         );
  DFFRHQX1 x4_89_tmp1_reg_3_ ( .D(n69), .CK(clk), .RN(rstn), .Q(x4_89_tmp1[3])
         );
  DFFRHQX1 x4_89_tmp1_reg_2_ ( .D(n68), .CK(clk), .RN(rstn), .Q(x4_89_tmp1[2])
         );
  DFFRHQX1 x4_89_reg_6_ ( .D(N363), .CK(clk), .RN(rstn), .Q(x4_89[6]) );
  DFFRHQX1 x4_89_reg_5_ ( .D(N362), .CK(clk), .RN(rstn), .Q(x4_89[5]) );
  DFFRHQX1 x4_89_reg_4_ ( .D(N361), .CK(clk), .RN(rstn), .Q(x4_89[4]) );
  DFFRHQX1 x4_89_reg_3_ ( .D(N360), .CK(clk), .RN(rstn), .Q(x4_89[3]) );
  DFFRHQX1 x4_75_reg_6_ ( .D(N386), .CK(clk), .RN(rstn), .Q(x4_75[6]) );
  DFFRHQX1 x4_75_reg_5_ ( .D(N385), .CK(clk), .RN(rstn), .Q(x4_75[5]) );
  DFFRHQX1 x4_75_reg_4_ ( .D(N384), .CK(clk), .RN(rstn), .Q(x4_75[4]) );
  DFFRHQX1 x4_75_reg_3_ ( .D(N383), .CK(clk), .RN(rstn), .Q(x4_75[3]) );
  DFFRHQX1 x5_75_reg_6_ ( .D(N475), .CK(clk), .RN(rstn), .Q(x5_75[6]) );
  DFFRHQX1 x5_75_reg_5_ ( .D(N474), .CK(clk), .RN(rstn), .Q(x5_75[5]) );
  DFFRHQX1 x5_75_reg_4_ ( .D(N473), .CK(clk), .RN(rstn), .Q(x5_75[4]) );
  DFFRHQX1 x5_75_reg_3_ ( .D(N472), .CK(clk), .RN(rstn), .Q(x5_75[3]) );
  DFFRHQX1 x6_75_reg_6_ ( .D(N564), .CK(clk), .RN(rstn), .Q(x6_75[6]) );
  DFFRHQX1 x6_75_reg_5_ ( .D(N563), .CK(clk), .RN(rstn), .Q(x6_75[5]) );
  DFFRHQX1 x6_75_reg_4_ ( .D(N562), .CK(clk), .RN(rstn), .Q(x6_75[4]) );
  DFFRHQX1 x6_75_reg_3_ ( .D(N561), .CK(clk), .RN(rstn), .Q(x6_75[3]) );
  DFFRHQX1 x4_50_reg_6_ ( .D(N409), .CK(clk), .RN(rstn), .Q(x4_50[6]) );
  DFFRHQX1 x4_50_reg_5_ ( .D(N408), .CK(clk), .RN(rstn), .Q(x4_50[5]) );
  DFFRHQX1 x4_50_reg_4_ ( .D(N407), .CK(clk), .RN(rstn), .Q(x4_50[4]) );
  DFFRHQX1 x4_50_reg_3_ ( .D(N406), .CK(clk), .RN(rstn), .Q(x4_50[3]) );
  DFFRHQX1 x5_tmp1_reg_7_ ( .D(N886), .CK(clk), .RN(rstn), .Q(x5_tmp1[7]) );
  DFFRHQX1 x5_tmp1_reg_6_ ( .D(N885), .CK(clk), .RN(rstn), .Q(x5_tmp1[6]) );
  DFFRHQX1 x5_tmp1_reg_5_ ( .D(N884), .CK(clk), .RN(rstn), .Q(x5_tmp1[5]) );
  DFFRHQX1 x5_tmp1_reg_4_ ( .D(N883), .CK(clk), .RN(rstn), .Q(x5_tmp1[4]) );
  DFFRHQX1 x6_tmp1_reg_7_ ( .D(N1052), .CK(clk), .RN(rstn), .Q(x6_tmp1[7]) );
  DFFRHQX1 x6_tmp1_reg_6_ ( .D(N1051), .CK(clk), .RN(rstn), .Q(x6_tmp1[6]) );
  DFFRHQX1 x6_tmp1_reg_5_ ( .D(N1050), .CK(clk), .RN(rstn), .Q(x6_tmp1[5]) );
  DFFRHQX1 x6_tmp1_reg_4_ ( .D(N1049), .CK(clk), .RN(rstn), .Q(x6_tmp1[4]) );
  DFFRHQX1 x7_tmp1_reg_7_ ( .D(N1149), .CK(clk), .RN(rstn), .Q(x7_tmp1[7]) );
  DFFRHQX1 x7_tmp1_reg_6_ ( .D(N1148), .CK(clk), .RN(rstn), .Q(x7_tmp1[6]) );
  DFFRHQX1 x7_tmp1_reg_5_ ( .D(N1147), .CK(clk), .RN(rstn), .Q(x7_tmp1[5]) );
  DFFRHQX1 x7_tmp1_reg_4_ ( .D(N1146), .CK(clk), .RN(rstn), .Q(x7_tmp1[4]) );
  DFFRHQX1 x4_tmp1_reg_7_ ( .D(N767), .CK(clk), .RN(rstn), .Q(x4_tmp1[7]) );
  DFFRHQX1 x4_tmp1_reg_6_ ( .D(N766), .CK(clk), .RN(rstn), .Q(x4_tmp1[6]) );
  DFFRHQX1 x4_tmp1_reg_5_ ( .D(N765), .CK(clk), .RN(rstn), .Q(x4_tmp1[5]) );
  DFFRHQX1 x4_tmp1_reg_4_ ( .D(N764), .CK(clk), .RN(rstn), .Q(x4_tmp1[4]) );
  DFFRHQX1 x6_89_reg_0_ ( .D(N535), .CK(clk), .RN(rstn), .Q(x6_89[0]) );
  DFFRHQX1 x7_50_reg_6_ ( .D(N676), .CK(clk), .RN(rstn), .Q(x7_50[6]) );
  DFFRHQX1 x7_50_reg_5_ ( .D(N675), .CK(clk), .RN(rstn), .Q(x7_50[5]) );
  DFFRHQX1 x7_50_reg_4_ ( .D(N674), .CK(clk), .RN(rstn), .Q(x7_50[4]) );
  DFFRHQX1 x7_50_reg_3_ ( .D(N673), .CK(clk), .RN(rstn), .Q(x7_50[3]) );
  DFFRHQX1 x5_89_reg_6_ ( .D(N452), .CK(clk), .RN(rstn), .Q(x5_89[6]) );
  DFFRHQX1 x5_89_reg_5_ ( .D(N451), .CK(clk), .RN(rstn), .Q(x5_89[5]) );
  DFFRHQX1 x5_89_reg_4_ ( .D(N450), .CK(clk), .RN(rstn), .Q(x5_89[4]) );
  DFFRHQX1 x5_89_reg_3_ ( .D(N449), .CK(clk), .RN(rstn), .Q(x5_89[3]) );
  DFFRHQX1 x7_89_reg_6_ ( .D(N630), .CK(clk), .RN(rstn), .Q(x7_89[6]) );
  DFFRHQX1 x7_89_reg_5_ ( .D(N629), .CK(clk), .RN(rstn), .Q(x7_89[5]) );
  DFFRHQX1 x7_89_reg_4_ ( .D(N628), .CK(clk), .RN(rstn), .Q(x7_89[4]) );
  DFFRHQX1 x7_89_reg_3_ ( .D(N627), .CK(clk), .RN(rstn), .Q(x7_89[3]) );
  DFFRHQX1 x5_50_reg_6_ ( .D(N498), .CK(clk), .RN(rstn), .Q(x5_50[6]) );
  DFFRHQX1 x5_50_reg_5_ ( .D(N497), .CK(clk), .RN(rstn), .Q(x5_50[5]) );
  DFFRHQX1 x5_50_reg_4_ ( .D(N496), .CK(clk), .RN(rstn), .Q(x5_50[4]) );
  DFFRHQX1 x5_50_reg_3_ ( .D(N495), .CK(clk), .RN(rstn), .Q(x5_50[3]) );
  DFFRHQX1 y6_tmp_reg_12_ ( .D(N1536), .CK(clk), .RN(rstn), .Q(y6_tmp[12]) );
  DFFRHQX1 y7_tmp_reg_12_ ( .D(N1613), .CK(clk), .RN(rstn), .Q(y7_tmp[12]) );
  DFFRHQX1 y0_tmp_reg_14_ ( .D(N1229), .CK(clk), .RN(rstn), .Q(y0_tmp[14]) );
  DFFRHQX1 y0_tmp_reg_13_ ( .D(N1228), .CK(clk), .RN(rstn), .Q(y0_tmp[13]) );
  DFFRHQX1 y0_tmp_reg_12_ ( .D(N1227), .CK(clk), .RN(rstn), .Q(y0_tmp[12]) );
  DFFRHQX1 y1_tmp_reg_14_ ( .D(N1255), .CK(clk), .RN(rstn), .Q(y1_tmp[14]) );
  DFFRHQX1 y1_tmp_reg_13_ ( .D(N1254), .CK(clk), .RN(rstn), .Q(y1_tmp[13]) );
  DFFRHQX1 y1_tmp_reg_12_ ( .D(N1253), .CK(clk), .RN(rstn), .Q(y1_tmp[12]) );
  DFFRHQX1 y2_tmp_reg_14_ ( .D(N1281), .CK(clk), .RN(rstn), .Q(y2_tmp[14]) );
  DFFRHQX1 y2_tmp_reg_13_ ( .D(N1280), .CK(clk), .RN(rstn), .Q(y2_tmp[13]) );
  DFFRHQX1 y2_tmp_reg_12_ ( .D(N1279), .CK(clk), .RN(rstn), .Q(y2_tmp[12]) );
  DFFRHQX1 y3_tmp_reg_14_ ( .D(N1307), .CK(clk), .RN(rstn), .Q(y3_tmp[14]) );
  DFFRHQX1 y3_tmp_reg_13_ ( .D(N1306), .CK(clk), .RN(rstn), .Q(y3_tmp[13]) );
  DFFRHQX1 y3_tmp_reg_12_ ( .D(N1305), .CK(clk), .RN(rstn), .Q(y3_tmp[12]) );
  DFFRHQX1 y4_tmp_reg_12_ ( .D(N1382), .CK(clk), .RN(rstn), .Q(y4_tmp[12]) );
  DFFRHQX1 y5_tmp_reg_12_ ( .D(N1459), .CK(clk), .RN(rstn), .Q(y5_tmp[12]) );
  DFFRHQX1 x6_89_tmp2_reg_5_ ( .D(N215), .CK(clk), .RN(rstn), .Q(x6_89_tmp2[5]) );
  DFFRHQX1 x6_89_tmp2_reg_4_ ( .D(N214), .CK(clk), .RN(rstn), .Q(x6_89_tmp2[4]) );
  DFFRHQX1 x6_89_tmp2_reg_3_ ( .D(x6[0]), .CK(clk), .RN(rstn), .Q(
        x6_89_tmp2[3]) );
  DFFRHQX1 x5_89_tmp2_reg_5_ ( .D(N130), .CK(clk), .RN(rstn), .Q(x5_89_tmp2[5]) );
  DFFRHQX1 x5_89_tmp2_reg_4_ ( .D(N129), .CK(clk), .RN(rstn), .Q(x5_89_tmp2[4]) );
  DFFRHQX1 x5_89_tmp2_reg_3_ ( .D(x5[0]), .CK(clk), .RN(rstn), .Q(
        x5_89_tmp2[3]) );
  DFFRHQX1 x4_89_tmp2_reg_5_ ( .D(N45), .CK(clk), .RN(rstn), .Q(x4_89_tmp2[5])
         );
  DFFRHQX1 x4_89_tmp2_reg_4_ ( .D(N44), .CK(clk), .RN(rstn), .Q(x4_89_tmp2[4])
         );
  DFFRHQX1 x4_89_tmp2_reg_3_ ( .D(x4[0]), .CK(clk), .RN(rstn), .Q(
        x4_89_tmp2[3]) );
  DFFRHQX1 x7_89_tmp2_reg_5_ ( .D(N300), .CK(clk), .RN(rstn), .Q(x7_89_tmp2[5]) );
  DFFRHQX1 x7_89_tmp2_reg_4_ ( .D(N299), .CK(clk), .RN(rstn), .Q(x7_89_tmp2[4]) );
  DFFRHQX1 x7_89_tmp2_reg_3_ ( .D(x7[0]), .CK(clk), .RN(rstn), .Q(
        x7_89_tmp2[3]) );
  DFFRHQX1 x4_75_tmp2_reg_5_ ( .D(N66), .CK(clk), .RN(rstn), .Q(x4_75_tmp2[5])
         );
  DFFRHQX1 x4_75_tmp2_reg_4_ ( .D(N65), .CK(clk), .RN(rstn), .Q(x4_75_tmp2[4])
         );
  DFFRHQX1 x4_75_tmp2_reg_3_ ( .D(N64), .CK(clk), .RN(rstn), .Q(x4_75_tmp2[3])
         );
  DFFRHQX1 x4_75_tmp2_reg_2_ ( .D(x4[1]), .CK(clk), .RN(rstn), .Q(
        x4_75_tmp2[2]) );
  DFFRHQX1 x4_75_tmp2_reg_1_ ( .D(x4[0]), .CK(clk), .RN(rstn), .Q(
        x4_75_tmp2[1]) );
  DFFRHQX1 x5_75_tmp2_reg_5_ ( .D(N151), .CK(clk), .RN(rstn), .Q(x5_75_tmp2[5]) );
  DFFRHQX1 x5_75_tmp2_reg_4_ ( .D(N150), .CK(clk), .RN(rstn), .Q(x5_75_tmp2[4]) );
  DFFRHQX1 x5_75_tmp2_reg_3_ ( .D(N149), .CK(clk), .RN(rstn), .Q(x5_75_tmp2[3]) );
  DFFRHQX1 x5_75_tmp2_reg_2_ ( .D(x5[1]), .CK(clk), .RN(rstn), .Q(
        x5_75_tmp2[2]) );
  DFFRHQX1 x5_75_tmp2_reg_1_ ( .D(x5[0]), .CK(clk), .RN(rstn), .Q(
        x5_75_tmp2[1]) );
  DFFRHQX1 x6_75_tmp2_reg_5_ ( .D(N236), .CK(clk), .RN(rstn), .Q(x6_75_tmp2[5]) );
  DFFRHQX1 x6_75_tmp2_reg_4_ ( .D(N235), .CK(clk), .RN(rstn), .Q(x6_75_tmp2[4]) );
  DFFRHQX1 x6_75_tmp2_reg_3_ ( .D(N234), .CK(clk), .RN(rstn), .Q(x6_75_tmp2[3]) );
  DFFRHQX1 x6_75_tmp2_reg_2_ ( .D(x6[1]), .CK(clk), .RN(rstn), .Q(
        x6_75_tmp2[2]) );
  DFFRHQX1 x6_75_tmp2_reg_1_ ( .D(x6[0]), .CK(clk), .RN(rstn), .Q(
        x6_75_tmp2[1]) );
  DFFRHQX1 x7_75_tmp2_reg_5_ ( .D(N321), .CK(clk), .RN(rstn), .Q(x7_75_tmp2[5]) );
  DFFRHQX1 x7_75_tmp2_reg_4_ ( .D(N320), .CK(clk), .RN(rstn), .Q(x7_75_tmp2[4]) );
  DFFRHQX1 x7_75_tmp2_reg_3_ ( .D(N319), .CK(clk), .RN(rstn), .Q(x7_75_tmp2[3]) );
  DFFRHQX1 x7_75_tmp2_reg_2_ ( .D(x7[1]), .CK(clk), .RN(rstn), .Q(
        x7_75_tmp2[2]) );
  DFFRHQX1 x7_75_tmp2_reg_1_ ( .D(x7[0]), .CK(clk), .RN(rstn), .Q(
        x7_75_tmp2[1]) );
  DFFRHQX1 x6_50_reg_2_ ( .D(N583), .CK(clk), .RN(rstn), .Q(x6_50[2]) );
  DFFRHQX1 x6_50_reg_3_ ( .D(N584), .CK(clk), .RN(rstn), .Q(x6_50[3]) );
  DFFRHQX1 x6_50_reg_4_ ( .D(N585), .CK(clk), .RN(rstn), .Q(x6_50[4]) );
  DFFRHQX1 x6_50_reg_5_ ( .D(N586), .CK(clk), .RN(rstn), .Q(x6_50[5]) );
  DFFRHQX1 x6_50_reg_6_ ( .D(N587), .CK(clk), .RN(rstn), .Q(x6_50[6]) );
  DFFRHQX1 x7_18_reg_6_ ( .D(N698), .CK(clk), .RN(rstn), .Q(x7_18[6]) );
  DFFRHQX1 x7_18_reg_5_ ( .D(N697), .CK(clk), .RN(rstn), .Q(x7_18[5]) );
  DFFRHQX1 x7_18_reg_4_ ( .D(N696), .CK(clk), .RN(rstn), .Q(x7_18[4]) );
  DFFRHQX1 x7_18_reg_3_ ( .D(N695), .CK(clk), .RN(rstn), .Q(x7_18[3]) );
  DFFRHQX1 x7_18_reg_2_ ( .D(N694), .CK(clk), .RN(rstn), .Q(x7_18[2]) );
  DFFRHQX1 x6_89_reg_7_ ( .D(N542), .CK(clk), .RN(rstn), .Q(x6_89[7]) );
  DFFRHQX1 x6_89_reg_6_ ( .D(N541), .CK(clk), .RN(rstn), .Q(x6_89[6]) );
  DFFRHQX1 x6_89_reg_5_ ( .D(N540), .CK(clk), .RN(rstn), .Q(x6_89[5]) );
  DFFRHQX1 x6_89_reg_4_ ( .D(N539), .CK(clk), .RN(rstn), .Q(x6_89[4]) );
  DFFRHQX1 x7_75_reg_6_ ( .D(N653), .CK(clk), .RN(rstn), .Q(x7_75[6]) );
  DFFRHQX1 x7_75_reg_5_ ( .D(N652), .CK(clk), .RN(rstn), .Q(x7_75[5]) );
  DFFRHQX1 x7_75_reg_4_ ( .D(N651), .CK(clk), .RN(rstn), .Q(x7_75[4]) );
  DFFRHQX1 x7_75_reg_3_ ( .D(N650), .CK(clk), .RN(rstn), .Q(x7_75[3]) );
  DFFRHQX1 x7_75_reg_2_ ( .D(N649), .CK(clk), .RN(rstn), .Q(x7_75[2]) );
  DFFRHQX1 x4_tmp2_reg_7_ ( .D(N837), .CK(clk), .RN(rstn), .Q(x4_tmp2[7]) );
  DFFRHQX1 x4_tmp2_reg_6_ ( .D(N836), .CK(clk), .RN(rstn), .Q(x4_tmp2[6]) );
  DFFRHQX1 x4_tmp2_reg_5_ ( .D(N835), .CK(clk), .RN(rstn), .Q(x4_tmp2[5]) );
  DFFRHQX1 x4_tmp2_reg_4_ ( .D(N834), .CK(clk), .RN(rstn), .Q(x4_tmp2[4]) );
  DFFRHQX1 x4_tmp2_reg_3_ ( .D(N833), .CK(clk), .RN(rstn), .Q(x4_tmp2[3]) );
  DFFRHQX1 x5_tmp2_reg_7_ ( .D(N957), .CK(clk), .RN(rstn), .Q(x5_tmp2[7]) );
  DFFRHQX1 x5_tmp2_reg_6_ ( .D(N956), .CK(clk), .RN(rstn), .Q(x5_tmp2[6]) );
  DFFRHQX1 x5_tmp2_reg_5_ ( .D(N955), .CK(clk), .RN(rstn), .Q(x5_tmp2[5]) );
  DFFRHQX1 x5_tmp2_reg_4_ ( .D(N954), .CK(clk), .RN(rstn), .Q(x5_tmp2[4]) );
  DFFRHQX1 x5_tmp2_reg_3_ ( .D(N953), .CK(clk), .RN(rstn), .Q(x5_tmp2[3]) );
  DFFRHQX1 x6_tmp2_reg_7_ ( .D(N1100), .CK(clk), .RN(rstn), .Q(x6_tmp2[7]) );
  DFFRHQX1 x6_tmp2_reg_6_ ( .D(N1099), .CK(clk), .RN(rstn), .Q(x6_tmp2[6]) );
  DFFRHQX1 x6_tmp2_reg_5_ ( .D(N1098), .CK(clk), .RN(rstn), .Q(x6_tmp2[5]) );
  DFFRHQX1 x6_tmp2_reg_4_ ( .D(N1097), .CK(clk), .RN(rstn), .Q(x6_tmp2[4]) );
  DFFRHQX1 x6_tmp2_reg_3_ ( .D(N1096), .CK(clk), .RN(rstn), .Q(x6_tmp2[3]) );
  DFFRHQX1 x7_tmp2_reg_7_ ( .D(N1173), .CK(clk), .RN(rstn), .Q(x7_tmp2[7]) );
  DFFRHQX1 x7_tmp2_reg_6_ ( .D(N1172), .CK(clk), .RN(rstn), .Q(x7_tmp2[6]) );
  DFFRHQX1 x7_tmp2_reg_5_ ( .D(N1171), .CK(clk), .RN(rstn), .Q(x7_tmp2[5]) );
  DFFRHQX1 x7_tmp2_reg_4_ ( .D(N1170), .CK(clk), .RN(rstn), .Q(x7_tmp2[4]) );
  DFFRHQX1 x7_tmp2_reg_3_ ( .D(N1169), .CK(clk), .RN(rstn), .Q(x7_tmp2[3]) );
  DFFRHQX1 y6_tmp_reg_11_ ( .D(N1535), .CK(clk), .RN(rstn), .Q(y6_tmp[11]) );
  DFFRHQX1 y7_tmp_reg_11_ ( .D(N1612), .CK(clk), .RN(rstn), .Q(y7_tmp[11]) );
  DFFRHQX1 y0_tmp_reg_11_ ( .D(N1226), .CK(clk), .RN(rstn), .Q(y0_tmp[11]) );
  DFFRHQX1 y1_tmp_reg_11_ ( .D(N1252), .CK(clk), .RN(rstn), .Q(y1_tmp[11]) );
  DFFRHQX1 y2_tmp_reg_11_ ( .D(N1278), .CK(clk), .RN(rstn), .Q(y2_tmp[11]) );
  DFFRHQX1 y3_tmp_reg_11_ ( .D(N1304), .CK(clk), .RN(rstn), .Q(y3_tmp[11]) );
  DFFRHQX1 y4_tmp_reg_11_ ( .D(N1381), .CK(clk), .RN(rstn), .Q(y4_tmp[11]) );
  DFFRHQX1 y5_tmp_reg_11_ ( .D(N1458), .CK(clk), .RN(rstn), .Q(y5_tmp[11]) );
  DFFRHQX1 x7_tmp_reg_5_ ( .D(N1195), .CK(clk), .RN(rstn), .Q(x7_tmp[5]) );
  DFFRHQX1 x7_tmp_reg_6_ ( .D(N1196), .CK(clk), .RN(rstn), .Q(x7_tmp[6]) );
  DFFRHQX1 x7_tmp_reg_7_ ( .D(N1197), .CK(clk), .RN(rstn), .Q(x7_tmp[7]) );
  DFFRHQX1 x7_tmp_reg_8_ ( .D(N1198), .CK(clk), .RN(rstn), .Q(x7_tmp[8]) );
  DFFRHQX1 x7_tmp_reg_9_ ( .D(N1199), .CK(clk), .RN(rstn), .Q(x7_tmp[9]) );
  DFFRHQX1 x5_tmp_reg_9_ ( .D(N983), .CK(clk), .RN(rstn), .Q(x5_tmp[9]) );
  DFFRHQX1 x5_tmp_reg_8_ ( .D(N982), .CK(clk), .RN(rstn), .Q(x5_tmp[8]) );
  DFFRHQX1 x5_tmp_reg_7_ ( .D(N981), .CK(clk), .RN(rstn), .Q(x5_tmp[7]) );
  DFFRHQX1 x5_tmp_reg_6_ ( .D(N980), .CK(clk), .RN(rstn), .Q(x5_tmp[6]) );
  DFFRHQX1 x5_tmp_reg_5_ ( .D(N979), .CK(clk), .RN(rstn), .Q(x5_tmp[5]) );
  DFFRHQX1 x6_tmp_reg_9_ ( .D(N1126), .CK(clk), .RN(rstn), .Q(x6_tmp[9]) );
  DFFRHQX1 x6_tmp_reg_8_ ( .D(N1125), .CK(clk), .RN(rstn), .Q(x6_tmp[8]) );
  DFFRHQX1 x6_tmp_reg_7_ ( .D(N1124), .CK(clk), .RN(rstn), .Q(x6_tmp[7]) );
  DFFRHQX1 x6_tmp_reg_6_ ( .D(N1123), .CK(clk), .RN(rstn), .Q(x6_tmp[6]) );
  DFFRHQX1 x6_tmp_reg_5_ ( .D(N1122), .CK(clk), .RN(rstn), .Q(x6_tmp[5]) );
  DFFRHQX1 x4_tmp_reg_5_ ( .D(N859), .CK(clk), .RN(rstn), .Q(x4_tmp[5]) );
  DFFRHQX1 x4_tmp_reg_6_ ( .D(N860), .CK(clk), .RN(rstn), .Q(x4_tmp[6]) );
  DFFRHQX1 x4_tmp_reg_7_ ( .D(N861), .CK(clk), .RN(rstn), .Q(x4_tmp[7]) );
  DFFRHQX1 x4_tmp_reg_8_ ( .D(N862), .CK(clk), .RN(rstn), .Q(x4_tmp[8]) );
  DFFRHQX1 x4_tmp_reg_9_ ( .D(N863), .CK(clk), .RN(rstn), .Q(x4_tmp[9]) );
  DFFRHQX1 x7_89_tmp1_reg_1_ ( .D(x7[1]), .CK(clk), .RN(rstn), .Q(
        x7_89_tmp1[1]) );
  DFFRHQX1 x6_89_tmp1_reg_1_ ( .D(x6[1]), .CK(clk), .RN(rstn), .Q(
        x6_89_tmp1[1]) );
  DFFRHQX1 x5_89_tmp1_reg_1_ ( .D(x5[1]), .CK(clk), .RN(rstn), .Q(
        x5_89_tmp1[1]) );
  DFFRHQX1 x5_75_tmp1_reg_1_ ( .D(x5[1]), .CK(clk), .RN(rstn), .Q(
        x5_75_tmp1[1]) );
  DFFRHQX1 x4_75_tmp1_reg_1_ ( .D(x4[1]), .CK(clk), .RN(rstn), .Q(
        x4_75_tmp1[1]) );
  DFFRHQX1 x7_75_tmp1_reg_1_ ( .D(x7[1]), .CK(clk), .RN(rstn), .Q(
        x7_75_tmp1[1]) );
  DFFRHQX1 x6_75_tmp1_reg_1_ ( .D(x6[1]), .CK(clk), .RN(rstn), .Q(
        x6_75_tmp1[1]) );
  DFFRHQX1 x5_18_reg_3_ ( .D(N517), .CK(clk), .RN(rstn), .Q(x5_18[3]) );
  DFFRHQX1 x5_18_reg_2_ ( .D(N516), .CK(clk), .RN(rstn), .Q(x5_18[2]) );
  DFFRHQX1 x5_18_reg_1_ ( .D(N515), .CK(clk), .RN(rstn), .Q(x5_18[1]) );
  DFFRHQX1 x6_18_reg_2_ ( .D(N605), .CK(clk), .RN(rstn), .Q(x6_18[2]) );
  DFFRHQX1 x6_18_reg_1_ ( .D(N604), .CK(clk), .RN(rstn), .Q(x6_18[1]) );
  DFFRHQX1 x4_18_reg_2_ ( .D(N427), .CK(clk), .RN(rstn), .Q(x4_18[2]) );
  DFFRHQX1 x4_18_reg_1_ ( .D(N426), .CK(clk), .RN(rstn), .Q(x4_18[1]) );
  DFFRHQX1 x4_89_tmp1_reg_1_ ( .D(x4[1]), .CK(clk), .RN(rstn), .Q(
        x4_89_tmp1[1]) );
  DFFRHQX1 x4_89_reg_2_ ( .D(N359), .CK(clk), .RN(rstn), .Q(x4_89[2]) );
  DFFRHQX1 x4_89_reg_1_ ( .D(N358), .CK(clk), .RN(rstn), .Q(x4_89[1]) );
  DFFRHQX1 x4_75_reg_2_ ( .D(N382), .CK(clk), .RN(rstn), .Q(x4_75[2]) );
  DFFRHQX1 x4_75_reg_1_ ( .D(N381), .CK(clk), .RN(rstn), .Q(x4_75[1]) );
  DFFRHQX1 x5_75_reg_2_ ( .D(N471), .CK(clk), .RN(rstn), .Q(x5_75[2]) );
  DFFRHQX1 x5_75_reg_1_ ( .D(N470), .CK(clk), .RN(rstn), .Q(x5_75[1]) );
  DFFRHQX1 x6_75_reg_2_ ( .D(N560), .CK(clk), .RN(rstn), .Q(x6_75[2]) );
  DFFRHQX1 x6_75_reg_1_ ( .D(N559), .CK(clk), .RN(rstn), .Q(x6_75[1]) );
  DFFRHQX1 x4_50_reg_2_ ( .D(N405), .CK(clk), .RN(rstn), .Q(x4_50[2]) );
  DFFRHQX1 x4_50_reg_1_ ( .D(N404), .CK(clk), .RN(rstn), .Q(x4_50[1]) );
  DFFRHQX1 x5_tmp1_reg_3_ ( .D(N882), .CK(clk), .RN(rstn), .Q(x5_tmp1[3]) );
  DFFRHQX1 x5_tmp1_reg_2_ ( .D(N881), .CK(clk), .RN(rstn), .Q(x5_tmp1[2]) );
  DFFRHQX1 x5_tmp1_reg_1_ ( .D(N880), .CK(clk), .RN(rstn), .Q(x5_tmp1[1]) );
  DFFRHQX1 x6_tmp1_reg_3_ ( .D(N1048), .CK(clk), .RN(rstn), .Q(x6_tmp1[3]) );
  DFFRHQX1 x6_tmp1_reg_2_ ( .D(N1047), .CK(clk), .RN(rstn), .Q(x6_tmp1[2]) );
  DFFRHQX1 x6_tmp1_reg_1_ ( .D(N1046), .CK(clk), .RN(rstn), .Q(x6_tmp1[1]) );
  DFFRHQX1 x7_tmp1_reg_3_ ( .D(N1145), .CK(clk), .RN(rstn), .Q(x7_tmp1[3]) );
  DFFRHQX1 x7_tmp1_reg_2_ ( .D(N1144), .CK(clk), .RN(rstn), .Q(x7_tmp1[2]) );
  DFFRHQX1 x7_tmp1_reg_1_ ( .D(N1143), .CK(clk), .RN(rstn), .Q(x7_tmp1[1]) );
  DFFRHQX1 x4_tmp1_reg_3_ ( .D(N763), .CK(clk), .RN(rstn), .Q(x4_tmp1[3]) );
  DFFRHQX1 x4_tmp1_reg_2_ ( .D(N762), .CK(clk), .RN(rstn), .Q(x4_tmp1[2]) );
  DFFRHQX1 x4_tmp1_reg_1_ ( .D(N761), .CK(clk), .RN(rstn), .Q(x4_tmp1[1]) );
  DFFRHQX1 x7_50_reg_2_ ( .D(N672), .CK(clk), .RN(rstn), .Q(x7_50[2]) );
  DFFRHQX1 x7_50_reg_1_ ( .D(N671), .CK(clk), .RN(rstn), .Q(x7_50[1]) );
  DFFRHQX1 x7_50_reg_0_ ( .D(1'b0), .CK(clk), .RN(rstn), .Q(x7_50[0]) );
  DFFRHQX1 x5_89_reg_2_ ( .D(N448), .CK(clk), .RN(rstn), .Q(x5_89[2]) );
  DFFRHQX1 x5_89_reg_1_ ( .D(N447), .CK(clk), .RN(rstn), .Q(x5_89[1]) );
  DFFRHQX1 x5_89_reg_0_ ( .D(N446), .CK(clk), .RN(rstn), .Q(x5_89[0]) );
  DFFRHQX1 x7_89_reg_2_ ( .D(N626), .CK(clk), .RN(rstn), .Q(x7_89[2]) );
  DFFRHQX1 x7_89_reg_1_ ( .D(N625), .CK(clk), .RN(rstn), .Q(x7_89[1]) );
  DFFRHQX1 x7_89_reg_0_ ( .D(N624), .CK(clk), .RN(rstn), .Q(x7_89[0]) );
  DFFRHQX1 x5_50_reg_2_ ( .D(N494), .CK(clk), .RN(rstn), .Q(x5_50[2]) );
  DFFRHQX1 x5_50_reg_1_ ( .D(N493), .CK(clk), .RN(rstn), .Q(x5_50[1]) );
  DFFRHQX1 x5_50_reg_0_ ( .D(1'b0), .CK(clk), .RN(rstn), .Q(x5_50[0]) );
  DFFRHQX1 x6_50_reg_1_ ( .D(N582), .CK(clk), .RN(rstn), .Q(x6_50[1]) );
  DFFRHQX1 x7_18_reg_1_ ( .D(N693), .CK(clk), .RN(rstn), .Q(x7_18[1]) );
  DFFRHQX1 x6_89_reg_3_ ( .D(N538), .CK(clk), .RN(rstn), .Q(x6_89[3]) );
  DFFRHQX1 x6_89_reg_2_ ( .D(N537), .CK(clk), .RN(rstn), .Q(x6_89[2]) );
  DFFRHQX1 x6_89_reg_1_ ( .D(N536), .CK(clk), .RN(rstn), .Q(x6_89[1]) );
  DFFRHQX1 x7_75_reg_1_ ( .D(N648), .CK(clk), .RN(rstn), .Q(x7_75[1]) );
  DFFRHQX1 x4_tmp2_reg_2_ ( .D(N832), .CK(clk), .RN(rstn), .Q(x4_tmp2[2]) );
  DFFRHQX1 x4_tmp2_reg_1_ ( .D(N831), .CK(clk), .RN(rstn), .Q(x4_tmp2[1]) );
  DFFRHQX1 x5_tmp2_reg_2_ ( .D(N952), .CK(clk), .RN(rstn), .Q(x5_tmp2[2]) );
  DFFRHQX1 x5_tmp2_reg_1_ ( .D(N951), .CK(clk), .RN(rstn), .Q(x5_tmp2[1]) );
  DFFRHQX1 x6_tmp2_reg_2_ ( .D(N1095), .CK(clk), .RN(rstn), .Q(x6_tmp2[2]) );
  DFFRHQX1 x6_tmp2_reg_1_ ( .D(N1094), .CK(clk), .RN(rstn), .Q(x6_tmp2[1]) );
  DFFRHQX1 x7_tmp2_reg_2_ ( .D(N1168), .CK(clk), .RN(rstn), .Q(x7_tmp2[2]) );
  DFFRHQX1 x7_tmp2_reg_1_ ( .D(N1167), .CK(clk), .RN(rstn), .Q(x7_tmp2[1]) );
  DFFRHQX1 x6_50_reg_0_ ( .D(1'b0), .CK(clk), .RN(rstn), .Q(x6_50[0]) );
  DFFRHQX1 x7_75_reg_0_ ( .D(N647), .CK(clk), .RN(rstn), .Q(x7_75[0]) );
  DFFRHQX1 x4_tmp2_reg_0_ ( .D(N830), .CK(clk), .RN(rstn), .Q(x4_tmp2[0]) );
  DFFRHQX1 x5_tmp2_reg_0_ ( .D(N950), .CK(clk), .RN(rstn), .Q(x5_tmp2[0]) );
  DFFRHQX1 x6_tmp2_reg_0_ ( .D(N1093), .CK(clk), .RN(rstn), .Q(x6_tmp2[0]) );
  DFFRHQX1 x7_tmp2_reg_0_ ( .D(N1166), .CK(clk), .RN(rstn), .Q(x7_tmp2[0]) );
  DFFRHQX1 x5_75_reg_0_ ( .D(N469), .CK(clk), .RN(rstn), .Q(x5_75[0]) );
  DFFRHQX1 x4_50_reg_0_ ( .D(1'b0), .CK(clk), .RN(rstn), .Q(x4_50[0]) );
  DFFRHQX1 x5_tmp1_reg_0_ ( .D(N879), .CK(clk), .RN(rstn), .Q(x5_tmp1[0]) );
  DFFRHQX1 x6_tmp1_reg_0_ ( .D(N1045), .CK(clk), .RN(rstn), .Q(x6_tmp1[0]) );
  DFFRHQX1 x7_tmp1_reg_0_ ( .D(N1142), .CK(clk), .RN(rstn), .Q(x7_tmp1[0]) );
  DFFRHQX1 x4_tmp1_reg_0_ ( .D(N760), .CK(clk), .RN(rstn), .Q(x4_tmp1[0]) );
  DFFRHQX1 x7_tmp_reg_1_ ( .D(N1191), .CK(clk), .RN(rstn), .Q(x7_tmp[1]) );
  DFFRHQX1 x7_tmp_reg_2_ ( .D(N1192), .CK(clk), .RN(rstn), .Q(x7_tmp[2]) );
  DFFRHQX1 x7_tmp_reg_3_ ( .D(N1193), .CK(clk), .RN(rstn), .Q(x7_tmp[3]) );
  DFFRHQX1 x7_tmp_reg_4_ ( .D(N1194), .CK(clk), .RN(rstn), .Q(x7_tmp[4]) );
  DFFRHQX1 x5_tmp_reg_4_ ( .D(N978), .CK(clk), .RN(rstn), .Q(x5_tmp[4]) );
  DFFRHQX1 x5_tmp_reg_3_ ( .D(N977), .CK(clk), .RN(rstn), .Q(x5_tmp[3]) );
  DFFRHQX1 x5_tmp_reg_2_ ( .D(N976), .CK(clk), .RN(rstn), .Q(x5_tmp[2]) );
  DFFRHQX1 x5_tmp_reg_1_ ( .D(N975), .CK(clk), .RN(rstn), .Q(x5_tmp[1]) );
  DFFRHQX1 x6_tmp_reg_4_ ( .D(N1121), .CK(clk), .RN(rstn), .Q(x6_tmp[4]) );
  DFFRHQX1 x6_tmp_reg_3_ ( .D(N1120), .CK(clk), .RN(rstn), .Q(x6_tmp[3]) );
  DFFRHQX1 x6_tmp_reg_2_ ( .D(N1119), .CK(clk), .RN(rstn), .Q(x6_tmp[2]) );
  DFFRHQX1 x6_tmp_reg_1_ ( .D(N1118), .CK(clk), .RN(rstn), .Q(x6_tmp[1]) );
  DFFRHQX1 x4_tmp_reg_1_ ( .D(N855), .CK(clk), .RN(rstn), .Q(x4_tmp[1]) );
  DFFRHQX1 x4_tmp_reg_2_ ( .D(N856), .CK(clk), .RN(rstn), .Q(x4_tmp[2]) );
  DFFRHQX1 x4_tmp_reg_3_ ( .D(N857), .CK(clk), .RN(rstn), .Q(x4_tmp[3]) );
  DFFRHQX1 x4_tmp_reg_4_ ( .D(N858), .CK(clk), .RN(rstn), .Q(x4_tmp[4]) );
  DFFRHQX1 x4_75_reg_0_ ( .D(N380), .CK(clk), .RN(rstn), .Q(x4_75[0]) );
  DFFRHQX1 x6_75_reg_0_ ( .D(N558), .CK(clk), .RN(rstn), .Q(x6_75[0]) );
  DFFRHQX1 x7_tmp_reg_0_ ( .D(N1190), .CK(clk), .RN(rstn), .Q(x7_tmp[0]) );
  DFFRHQX1 x5_tmp_reg_0_ ( .D(N974), .CK(clk), .RN(rstn), .Q(x5_tmp[0]) );
  DFFRHQX1 x6_tmp_reg_0_ ( .D(N1117), .CK(clk), .RN(rstn), .Q(x6_tmp[0]) );
  DFFRHQX1 x4_tmp_reg_0_ ( .D(N854), .CK(clk), .RN(rstn), .Q(x4_tmp[0]) );
  DFFRHQX1 mode_delay1_reg_1_ ( .D(mode[1]), .CK(clk), .RN(rstn), .Q(
        mode_delay1[1]) );
  DFFRHQX1 mode_delay1_reg_0_ ( .D(mode[0]), .CK(clk), .RN(rstn), .Q(
        mode_delay1[0]) );
  AND2X2 U13 ( .A(y1_tmp[23]), .B(n92), .Y(y1[23]) );
  AND2X2 U14 ( .A(y1_tmp[24]), .B(n92), .Y(y1[24]) );
  AND2X2 U15 ( .A(y1_tmp[25]), .B(n92), .Y(y1[25]) );
  AND2X2 U16 ( .A(y2_tmp[17]), .B(n92), .Y(y2[17]) );
  AND2X2 U17 ( .A(y2_tmp[18]), .B(n92), .Y(y2[18]) );
  AND2X2 U18 ( .A(y2_tmp[19]), .B(n92), .Y(y2[19]) );
  AND2X2 U19 ( .A(y2_tmp[20]), .B(n92), .Y(y2[20]) );
  AND2X2 U47 ( .A(y2_tmp[21]), .B(n92), .Y(y2[21]) );
  AND2X2 U48 ( .A(y4_tmp[17]), .B(n92), .Y(y4[17]) );
  AND2X2 U49 ( .A(y4_tmp[19]), .B(n92), .Y(y4[19]) );
  AND2X2 U50 ( .A(y4_tmp[20]), .B(n92), .Y(y4[20]) );
  AND2X2 U51 ( .A(y4_tmp[21]), .B(n92), .Y(y4[21]) );
  AND2X2 U52 ( .A(y4_tmp[22]), .B(n92), .Y(y4[22]) );
  AND2X2 U53 ( .A(y4_tmp[23]), .B(n92), .Y(y4[23]) );
  AND2X2 U54 ( .A(y4_tmp[24]), .B(n92), .Y(y4[24]) );
  AND2X2 U55 ( .A(y4_tmp[25]), .B(n92), .Y(y4[25]) );
  AND2X2 U56 ( .A(y5_tmp[17]), .B(n92), .Y(y5[17]) );
  AND2X2 U57 ( .A(y5_tmp[18]), .B(n92), .Y(y5[18]) );
  AND2X2 U58 ( .A(y5_tmp[19]), .B(n92), .Y(y5[19]) );
  AND2X2 U59 ( .A(y5_tmp[20]), .B(n92), .Y(y5[20]) );
  AND2X2 U60 ( .A(y5_tmp[21]), .B(n92), .Y(y5[21]) );
  AND2X2 U61 ( .A(y5_tmp[23]), .B(n92), .Y(y5[23]) );
  AND2X2 U62 ( .A(y5_tmp[24]), .B(n92), .Y(y5[24]) );
  AND2X2 U94 ( .A(y0_tmp[20]), .B(n176), .Y(y0[20]) );
  AND2X2 U95 ( .A(y0_tmp[22]), .B(n171), .Y(y0[22]) );
  AND2X2 U96 ( .A(y0_tmp[23]), .B(n172), .Y(y0[23]) );
  AND2X2 U97 ( .A(y0_tmp[24]), .B(n174), .Y(y0[24]) );
  AND2X2 U98 ( .A(y0_tmp[25]), .B(n167), .Y(y0[25]) );
  AND2X2 U99 ( .A(y1_tmp[17]), .B(n176), .Y(y1[17]) );
  AND2X2 U100 ( .A(y1_tmp[18]), .B(n175), .Y(y1[18]) );
  AND2X2 U101 ( .A(y1_tmp[19]), .B(n171), .Y(y1[19]) );
  AND2X2 U102 ( .A(y1_tmp[20]), .B(n172), .Y(y1[20]) );
  AND2X2 U103 ( .A(y1_tmp[21]), .B(n174), .Y(y1[21]) );
  AND2X2 U104 ( .A(y1_tmp[22]), .B(n167), .Y(y1[22]) );
  AND2X2 U105 ( .A(y2_tmp[22]), .B(n176), .Y(y2[22]) );
  AND2X2 U106 ( .A(y2_tmp[23]), .B(n173), .Y(y2[23]) );
  AND2X2 U107 ( .A(y2_tmp[24]), .B(n166), .Y(y2[24]) );
  AND2X2 U108 ( .A(y2_tmp[25]), .B(n170), .Y(y2[25]) );
  AND2X2 U109 ( .A(y3_tmp[20]), .B(n168), .Y(y3[20]) );
  AND2X2 U110 ( .A(y3_tmp[21]), .B(n169), .Y(y3[21]) );
  AND2X2 U111 ( .A(y3_tmp[22]), .B(n175), .Y(y3[22]) );
  AND2X2 U112 ( .A(y3_tmp[23]), .B(n171), .Y(y3[23]) );
  AND2X2 U113 ( .A(y3_tmp[24]), .B(n172), .Y(y3[24]) );
  AND2X2 U114 ( .A(y3_tmp[25]), .B(n174), .Y(y3[25]) );
  AND2X2 U115 ( .A(y4_tmp[18]), .B(n167), .Y(y4[18]) );
  AND2X2 U116 ( .A(y5_tmp[22]), .B(n176), .Y(y5[22]) );
  AND2X2 U117 ( .A(y5_tmp[25]), .B(n173), .Y(y5[25]) );
  AND2X2 U118 ( .A(y6_tmp[17]), .B(n166), .Y(y6[17]) );
  AND2X2 U119 ( .A(y6_tmp[18]), .B(n170), .Y(y6[18]) );
  AND2X2 U120 ( .A(y6_tmp[19]), .B(n168), .Y(y6[19]) );
  AND2X2 U121 ( .A(y6_tmp[20]), .B(n169), .Y(y6[20]) );
  AND2X2 U122 ( .A(y6_tmp[22]), .B(n175), .Y(y6[22]) );
  AND2X2 U123 ( .A(y6_tmp[23]), .B(n171), .Y(y6[23]) );
  AND2X2 U124 ( .A(y6_tmp[24]), .B(n172), .Y(y6[24]) );
  AND2X2 U125 ( .A(y6_tmp[25]), .B(n174), .Y(y6[25]) );
  AND2X2 U126 ( .A(y0_tmp[17]), .B(n175), .Y(y0[17]) );
  AND2X2 U127 ( .A(y0_tmp[18]), .B(n166), .Y(y0[18]) );
  AND2X2 U128 ( .A(y0_tmp[19]), .B(n170), .Y(y0[19]) );
  AND2X2 U129 ( .A(y0_tmp[21]), .B(n168), .Y(y0[21]) );
  AND2X2 U130 ( .A(y3_tmp[17]), .B(n169), .Y(y3[17]) );
  AND2X2 U131 ( .A(y3_tmp[18]), .B(n173), .Y(y3[18]) );
  AND2X2 U132 ( .A(y3_tmp[19]), .B(n171), .Y(y3[19]) );
  AND2X2 U133 ( .A(y6_tmp[21]), .B(n172), .Y(y6[21]) );
  AND2X2 U134 ( .A(y7_tmp[17]), .B(n174), .Y(y7[17]) );
  AND2X2 U135 ( .A(y7_tmp[18]), .B(n176), .Y(y7[18]) );
  AND2X2 U136 ( .A(y7_tmp[19]), .B(n167), .Y(y7[19]) );
  AND2X2 U137 ( .A(y7_tmp[20]), .B(n175), .Y(y7[20]) );
  AND2X2 U138 ( .A(y7_tmp[21]), .B(n166), .Y(y7[21]) );
  AND2X2 U139 ( .A(y7_tmp[22]), .B(n170), .Y(y7[22]) );
  AND2X2 U140 ( .A(y7_tmp[23]), .B(n168), .Y(y7[23]) );
  AND2X2 U141 ( .A(y7_tmp[24]), .B(n169), .Y(y7[24]) );
  AND2X2 U142 ( .A(y7_tmp[25]), .B(n173), .Y(y7[25]) );
  INVX1 U143 ( .A(n158), .Y(n92) );
  INVX1 U144 ( .A(n157), .Y(n88) );
  INVX1 U145 ( .A(n158), .Y(n89) );
  INVX1 U146 ( .A(n158), .Y(n90) );
  INVX1 U147 ( .A(n158), .Y(n91) );
  INVX1 U148 ( .A(n157), .Y(n86) );
  INVX1 U149 ( .A(n157), .Y(n87) );
  INVX1 U150 ( .A(n156), .Y(n81) );
  INVX1 U151 ( .A(n157), .Y(n85) );
  INVX1 U152 ( .A(n156), .Y(n84) );
  INVX1 U153 ( .A(n156), .Y(n83) );
  INVX1 U154 ( .A(n156), .Y(n82) );
  INVX1 U155 ( .A(n159), .Y(n157) );
  INVX1 U156 ( .A(n454), .Y(n158) );
  INVX1 U157 ( .A(n162), .Y(n156) );
  INVX1 U158 ( .A(n159), .Y(n152) );
  INVX1 U159 ( .A(n160), .Y(n151) );
  INVX1 U160 ( .A(n160), .Y(n150) );
  INVX1 U161 ( .A(n160), .Y(n149) );
  INVX1 U162 ( .A(n163), .Y(n155) );
  INVX1 U163 ( .A(n159), .Y(n154) );
  INVX1 U164 ( .A(n159), .Y(n153) );
  INVX1 U165 ( .A(n161), .Y(n148) );
  INVX1 U166 ( .A(n160), .Y(n144) );
  INVX1 U167 ( .A(n162), .Y(n143) );
  INVX1 U168 ( .A(n162), .Y(n142) );
  INVX1 U169 ( .A(n162), .Y(n141) );
  INVX1 U170 ( .A(n161), .Y(n147) );
  INVX1 U171 ( .A(n161), .Y(n146) );
  INVX1 U172 ( .A(n161), .Y(n145) );
  INVX1 U173 ( .A(n163), .Y(n137) );
  INVX1 U174 ( .A(n163), .Y(n136) );
  INVX1 U175 ( .A(n164), .Y(n135) );
  INVX1 U176 ( .A(n164), .Y(n134) );
  INVX1 U177 ( .A(n162), .Y(n140) );
  INVX1 U178 ( .A(n163), .Y(n139) );
  INVX1 U179 ( .A(n163), .Y(n138) );
  INVX1 U180 ( .A(n164), .Y(n133) );
  INVX1 U181 ( .A(n165), .Y(n129) );
  INVX1 U182 ( .A(n163), .Y(n128) );
  INVX1 U183 ( .A(n164), .Y(n127) );
  INVX1 U184 ( .A(n165), .Y(n132) );
  INVX1 U185 ( .A(n165), .Y(n131) );
  INVX1 U186 ( .A(n165), .Y(n130) );
  INVX1 U187 ( .A(n167), .Y(n122) );
  INVX1 U188 ( .A(n167), .Y(n121) );
  INVX1 U189 ( .A(n167), .Y(n120) );
  INVX1 U190 ( .A(n168), .Y(n119) );
  INVX1 U191 ( .A(n170), .Y(n126) );
  INVX1 U192 ( .A(n166), .Y(n125) );
  INVX1 U193 ( .A(n166), .Y(n124) );
  INVX1 U194 ( .A(n166), .Y(n123) );
  INVX1 U195 ( .A(n168), .Y(n118) );
  INVX1 U196 ( .A(n169), .Y(n114) );
  INVX1 U197 ( .A(n170), .Y(n113) );
  INVX1 U198 ( .A(n170), .Y(n112) );
  INVX1 U199 ( .A(n170), .Y(n111) );
  INVX1 U200 ( .A(n171), .Y(n110) );
  INVX1 U201 ( .A(n168), .Y(n117) );
  INVX1 U202 ( .A(n169), .Y(n116) );
  INVX1 U203 ( .A(n169), .Y(n115) );
  INVX1 U204 ( .A(n172), .Y(n105) );
  INVX1 U205 ( .A(n173), .Y(n104) );
  INVX1 U206 ( .A(n173), .Y(n103) );
  INVX1 U207 ( .A(n173), .Y(n102) );
  INVX1 U208 ( .A(n171), .Y(n109) );
  INVX1 U209 ( .A(n171), .Y(n108) );
  INVX1 U210 ( .A(n172), .Y(n107) );
  INVX1 U211 ( .A(n172), .Y(n106) );
  INVX1 U212 ( .A(n174), .Y(n101) );
  INVX1 U213 ( .A(n175), .Y(n97) );
  INVX1 U214 ( .A(n175), .Y(n96) );
  INVX1 U215 ( .A(n176), .Y(n95) );
  INVX1 U216 ( .A(n176), .Y(n94) );
  INVX1 U217 ( .A(n176), .Y(n93) );
  INVX1 U218 ( .A(n174), .Y(n100) );
  INVX1 U219 ( .A(n174), .Y(n99) );
  INVX1 U220 ( .A(n175), .Y(n98) );
  ADDFX2 U221 ( .A(x7[15]), .B(x7[15]), .CI(N355), .CO(N356) );
  ADDFX2 U222 ( .A(x5[15]), .B(x5[15]), .CI(N185), .CO(N186) );
  ADDFX2 U223 ( .A(x6[15]), .B(x6[15]), .CI(N270), .CO(N271) );
  ADDFX2 U224 ( .A(x4[15]), .B(x4[15]), .CI(N100), .CO(N101) );
  ADDFX2 U225 ( .A(x7[15]), .B(x7[15]), .CI(N334), .CO(N335) );
  ADDFX2 U226 ( .A(x6[15]), .B(x6[15]), .CI(N249), .CO(N250) );
  ADDFX2 U227 ( .A(x5[15]), .B(x5[15]), .CI(N164), .CO(N165) );
  ADDFX2 U228 ( .A(x4[15]), .B(x4[15]), .CI(N79), .CO(N80) );
  ADDFX2 U229 ( .A(x7[15]), .B(x7[15]), .CI(N314), .CO(N315) );
  ADDFX2 U230 ( .A(x4[15]), .B(x4[15]), .CI(N59), .CO(N60) );
  ADDFX2 U231 ( .A(x5[15]), .B(x5[15]), .CI(N144), .CO(N145) );
  ADDFX2 U232 ( .A(x6[15]), .B(x6[15]), .CI(N229), .CO(N230) );
  INVX1 U233 ( .A(n177), .Y(n160) );
  INVX1 U234 ( .A(n181), .Y(n159) );
  INVX1 U235 ( .A(n182), .Y(n162) );
  INVX1 U236 ( .A(n178), .Y(n161) );
  INVX1 U237 ( .A(n182), .Y(n163) );
  INVX1 U238 ( .A(n181), .Y(n164) );
  INVX1 U239 ( .A(n181), .Y(n165) );
  INVX1 U240 ( .A(n180), .Y(n167) );
  INVX1 U241 ( .A(n180), .Y(n166) );
  INVX1 U242 ( .A(n179), .Y(n170) );
  INVX1 U243 ( .A(n179), .Y(n168) );
  INVX1 U244 ( .A(n179), .Y(n169) );
  INVX1 U245 ( .A(n178), .Y(n173) );
  INVX1 U246 ( .A(n178), .Y(n171) );
  INVX1 U247 ( .A(n178), .Y(n172) );
  INVX1 U248 ( .A(n177), .Y(n176) );
  INVX1 U249 ( .A(n177), .Y(n174) );
  INVX1 U250 ( .A(n177), .Y(n175) );
  ADDFX2 U251 ( .A(n41), .B(x7[15]), .CI(add_104_carry_18_), .CO(N355), .S(
        N354) );
  ADDFX2 U252 ( .A(n67), .B(x5[15]), .CI(add_86_carry_18_), .CO(N185), .S(N184) );
  ADDFX2 U253 ( .A(n54), .B(x6[15]), .CI(add_95_carry_18_), .CO(N270), .S(N269) );
  ADDFX2 U254 ( .A(n80), .B(x4[15]), .CI(add_77_carry_18_), .CO(N100), .S(N99)
         );
  ADDFX2 U255 ( .A(n41), .B(x7[15]), .CI(add_102_carry_17_), .CO(N334), .S(
        N333) );
  ADDFX2 U256 ( .A(n54), .B(x6[15]), .CI(add_93_carry_17_), .CO(N249), .S(N248) );
  ADDFX2 U257 ( .A(n67), .B(x5[15]), .CI(add_84_carry_17_), .CO(N164), .S(N163) );
  ADDFX2 U258 ( .A(n80), .B(x4[15]), .CI(add_75_carry_17_), .CO(N79), .S(N78)
         );
  ADDFX2 U259 ( .A(n41), .B(x7[15]), .CI(add_100_carry_18_), .CO(N314), .S(
        N313) );
  ADDFX2 U260 ( .A(n80), .B(x4[15]), .CI(add_73_carry_18_), .CO(N59), .S(N58)
         );
  ADDFX2 U261 ( .A(n67), .B(x5[15]), .CI(add_82_carry_18_), .CO(N144), .S(N143) );
  ADDFX2 U262 ( .A(n54), .B(x6[15]), .CI(add_91_carry_18_), .CO(N229), .S(N228) );
  ADDFX2 U263 ( .A(n80), .B(x4[15]), .CI(add_72_carry_20_), .CO(N38), .S(N37)
         );
  ADDFX2 U264 ( .A(n67), .B(x5[15]), .CI(add_81_carry_20_), .CO(N123), .S(N122) );
  ADDFX2 U265 ( .A(n54), .B(x6[15]), .CI(add_90_carry_20_), .CO(N208), .S(N207) );
  ADDFX2 U266 ( .A(n41), .B(x7[15]), .CI(add_99_carry_20_), .CO(N293), .S(N292) );
  ADDFX2 U267 ( .A(n2), .B(n5), .CI(add_104_carry_6_), .CO(add_104_carry_7_), 
        .S(N342) );
  ADDFX2 U268 ( .A(n3), .B(n6), .CI(add_104_carry_7_), .CO(add_104_carry_8_), 
        .S(N343) );
  ADDFX2 U269 ( .A(n4), .B(n7), .CI(add_104_carry_8_), .CO(add_104_carry_9_), 
        .S(N344) );
  ADDFX2 U270 ( .A(n5), .B(n8), .CI(add_104_carry_9_), .CO(add_104_carry_10_), 
        .S(N345) );
  ADDFX2 U271 ( .A(n6), .B(n36), .CI(add_104_carry_10_), .CO(add_104_carry_11_), .S(N346) );
  ADDFX2 U272 ( .A(n7), .B(n37), .CI(add_104_carry_11_), .CO(add_104_carry_12_), .S(N347) );
  ADDFX2 U273 ( .A(n8), .B(n38), .CI(add_104_carry_12_), .CO(add_104_carry_13_), .S(N348) );
  ADDFX2 U274 ( .A(n36), .B(n39), .CI(add_104_carry_13_), .CO(
        add_104_carry_14_), .S(N349) );
  ADDFX2 U275 ( .A(n37), .B(n40), .CI(add_104_carry_14_), .CO(
        add_104_carry_15_), .S(N350) );
  ADDFX2 U276 ( .A(n38), .B(n41), .CI(add_104_carry_15_), .CO(
        add_104_carry_16_), .S(N351) );
  ADDFX2 U277 ( .A(n39), .B(x7[15]), .CI(add_104_carry_16_), .CO(
        add_104_carry_17_), .S(N352) );
  ADDFX2 U278 ( .A(n40), .B(x7[15]), .CI(add_104_carry_17_), .CO(
        add_104_carry_18_), .S(N353) );
  ADDFX2 U279 ( .A(n55), .B(n58), .CI(add_86_carry_6_), .CO(add_86_carry_7_), 
        .S(N172) );
  ADDFX2 U280 ( .A(n56), .B(n59), .CI(add_86_carry_7_), .CO(add_86_carry_8_), 
        .S(N173) );
  ADDFX2 U281 ( .A(n57), .B(n60), .CI(add_86_carry_8_), .CO(add_86_carry_9_), 
        .S(N174) );
  ADDFX2 U282 ( .A(n58), .B(n61), .CI(add_86_carry_9_), .CO(add_86_carry_10_), 
        .S(N175) );
  ADDFX2 U283 ( .A(n59), .B(n62), .CI(add_86_carry_10_), .CO(add_86_carry_11_), 
        .S(N176) );
  ADDFX2 U284 ( .A(n60), .B(n63), .CI(add_86_carry_11_), .CO(add_86_carry_12_), 
        .S(N177) );
  ADDFX2 U285 ( .A(n61), .B(n64), .CI(add_86_carry_12_), .CO(add_86_carry_13_), 
        .S(N178) );
  ADDFX2 U286 ( .A(n62), .B(n65), .CI(add_86_carry_13_), .CO(add_86_carry_14_), 
        .S(N179) );
  ADDFX2 U287 ( .A(n63), .B(n66), .CI(add_86_carry_14_), .CO(add_86_carry_15_), 
        .S(N180) );
  ADDFX2 U288 ( .A(n64), .B(n67), .CI(add_86_carry_15_), .CO(add_86_carry_16_), 
        .S(N181) );
  ADDFX2 U289 ( .A(n65), .B(x5[15]), .CI(add_86_carry_16_), .CO(
        add_86_carry_17_), .S(N182) );
  ADDFX2 U290 ( .A(n66), .B(x5[15]), .CI(add_86_carry_17_), .CO(
        add_86_carry_18_), .S(N183) );
  ADDFX2 U291 ( .A(n42), .B(n45), .CI(add_95_carry_6_), .CO(add_95_carry_7_), 
        .S(N257) );
  ADDFX2 U292 ( .A(n43), .B(n46), .CI(add_95_carry_7_), .CO(add_95_carry_8_), 
        .S(N258) );
  ADDFX2 U293 ( .A(n44), .B(n47), .CI(add_95_carry_8_), .CO(add_95_carry_9_), 
        .S(N259) );
  ADDFX2 U294 ( .A(n45), .B(n48), .CI(add_95_carry_9_), .CO(add_95_carry_10_), 
        .S(N260) );
  ADDFX2 U295 ( .A(n46), .B(n49), .CI(add_95_carry_10_), .CO(add_95_carry_11_), 
        .S(N261) );
  ADDFX2 U296 ( .A(n47), .B(n50), .CI(add_95_carry_11_), .CO(add_95_carry_12_), 
        .S(N262) );
  ADDFX2 U297 ( .A(n48), .B(n51), .CI(add_95_carry_12_), .CO(add_95_carry_13_), 
        .S(N263) );
  ADDFX2 U298 ( .A(n49), .B(n52), .CI(add_95_carry_13_), .CO(add_95_carry_14_), 
        .S(N264) );
  ADDFX2 U299 ( .A(n50), .B(n53), .CI(add_95_carry_14_), .CO(add_95_carry_15_), 
        .S(N265) );
  ADDFX2 U300 ( .A(n51), .B(n54), .CI(add_95_carry_15_), .CO(add_95_carry_16_), 
        .S(N266) );
  ADDFX2 U301 ( .A(n52), .B(x6[15]), .CI(add_95_carry_16_), .CO(
        add_95_carry_17_), .S(N267) );
  ADDFX2 U302 ( .A(n53), .B(x6[15]), .CI(add_95_carry_17_), .CO(
        add_95_carry_18_), .S(N268) );
  ADDFX2 U303 ( .A(n68), .B(n71), .CI(add_77_carry_6_), .CO(add_77_carry_7_), 
        .S(N87) );
  ADDFX2 U304 ( .A(n69), .B(n72), .CI(add_77_carry_7_), .CO(add_77_carry_8_), 
        .S(N88) );
  ADDFX2 U305 ( .A(n70), .B(n73), .CI(add_77_carry_8_), .CO(add_77_carry_9_), 
        .S(N89) );
  ADDFX2 U306 ( .A(n71), .B(n74), .CI(add_77_carry_9_), .CO(add_77_carry_10_), 
        .S(N90) );
  ADDFX2 U307 ( .A(n72), .B(n75), .CI(add_77_carry_10_), .CO(add_77_carry_11_), 
        .S(N91) );
  ADDFX2 U308 ( .A(n73), .B(n76), .CI(add_77_carry_11_), .CO(add_77_carry_12_), 
        .S(N92) );
  ADDFX2 U309 ( .A(n74), .B(n77), .CI(add_77_carry_12_), .CO(add_77_carry_13_), 
        .S(N93) );
  ADDFX2 U310 ( .A(n75), .B(n78), .CI(add_77_carry_13_), .CO(add_77_carry_14_), 
        .S(N94) );
  ADDFX2 U311 ( .A(n76), .B(n79), .CI(add_77_carry_14_), .CO(add_77_carry_15_), 
        .S(N95) );
  ADDFX2 U312 ( .A(n77), .B(n80), .CI(add_77_carry_15_), .CO(add_77_carry_16_), 
        .S(N96) );
  ADDFX2 U313 ( .A(n78), .B(x4[15]), .CI(add_77_carry_16_), .CO(
        add_77_carry_17_), .S(N97) );
  ADDFX2 U314 ( .A(n79), .B(x4[15]), .CI(add_77_carry_17_), .CO(
        add_77_carry_18_), .S(N98) );
  ADDFX2 U315 ( .A(n2), .B(n4), .CI(add_102_carry_5_), .CO(add_102_carry_6_), 
        .S(N321) );
  ADDFX2 U316 ( .A(n3), .B(n5), .CI(add_102_carry_6_), .CO(add_102_carry_7_), 
        .S(N322) );
  ADDFX2 U317 ( .A(n4), .B(n6), .CI(add_102_carry_7_), .CO(add_102_carry_8_), 
        .S(N323) );
  ADDFX2 U318 ( .A(n5), .B(n7), .CI(add_102_carry_8_), .CO(add_102_carry_9_), 
        .S(N324) );
  ADDFX2 U319 ( .A(n6), .B(n8), .CI(add_102_carry_9_), .CO(add_102_carry_10_), 
        .S(N325) );
  ADDFX2 U320 ( .A(n7), .B(n36), .CI(add_102_carry_10_), .CO(add_102_carry_11_), .S(N326) );
  ADDFX2 U321 ( .A(n8), .B(n37), .CI(add_102_carry_11_), .CO(add_102_carry_12_), .S(N327) );
  ADDFX2 U322 ( .A(n36), .B(n38), .CI(add_102_carry_12_), .CO(
        add_102_carry_13_), .S(N328) );
  ADDFX2 U323 ( .A(n37), .B(n39), .CI(add_102_carry_13_), .CO(
        add_102_carry_14_), .S(N329) );
  ADDFX2 U324 ( .A(n38), .B(n40), .CI(add_102_carry_14_), .CO(
        add_102_carry_15_), .S(N330) );
  ADDFX2 U325 ( .A(n39), .B(n41), .CI(add_102_carry_15_), .CO(
        add_102_carry_16_), .S(N331) );
  ADDFX2 U326 ( .A(n40), .B(x7[15]), .CI(add_102_carry_16_), .CO(
        add_102_carry_17_), .S(N332) );
  ADDFX2 U327 ( .A(n42), .B(n44), .CI(add_93_carry_5_), .CO(add_93_carry_6_), 
        .S(N236) );
  ADDFX2 U328 ( .A(n43), .B(n45), .CI(add_93_carry_6_), .CO(add_93_carry_7_), 
        .S(N237) );
  ADDFX2 U329 ( .A(n44), .B(n46), .CI(add_93_carry_7_), .CO(add_93_carry_8_), 
        .S(N238) );
  ADDFX2 U330 ( .A(n45), .B(n47), .CI(add_93_carry_8_), .CO(add_93_carry_9_), 
        .S(N239) );
  ADDFX2 U331 ( .A(n46), .B(n48), .CI(add_93_carry_9_), .CO(add_93_carry_10_), 
        .S(N240) );
  ADDFX2 U332 ( .A(n47), .B(n49), .CI(add_93_carry_10_), .CO(add_93_carry_11_), 
        .S(N241) );
  ADDFX2 U333 ( .A(n48), .B(n50), .CI(add_93_carry_11_), .CO(add_93_carry_12_), 
        .S(N242) );
  ADDFX2 U334 ( .A(n49), .B(n51), .CI(add_93_carry_12_), .CO(add_93_carry_13_), 
        .S(N243) );
  ADDFX2 U335 ( .A(n50), .B(n52), .CI(add_93_carry_13_), .CO(add_93_carry_14_), 
        .S(N244) );
  ADDFX2 U336 ( .A(n51), .B(n53), .CI(add_93_carry_14_), .CO(add_93_carry_15_), 
        .S(N245) );
  ADDFX2 U337 ( .A(n52), .B(n54), .CI(add_93_carry_15_), .CO(add_93_carry_16_), 
        .S(N246) );
  ADDFX2 U338 ( .A(n53), .B(x6[15]), .CI(add_93_carry_16_), .CO(
        add_93_carry_17_), .S(N247) );
  ADDFX2 U339 ( .A(n55), .B(n57), .CI(add_84_carry_5_), .CO(add_84_carry_6_), 
        .S(N151) );
  ADDFX2 U340 ( .A(n56), .B(n58), .CI(add_84_carry_6_), .CO(add_84_carry_7_), 
        .S(N152) );
  ADDFX2 U341 ( .A(n57), .B(n59), .CI(add_84_carry_7_), .CO(add_84_carry_8_), 
        .S(N153) );
  ADDFX2 U342 ( .A(n58), .B(n60), .CI(add_84_carry_8_), .CO(add_84_carry_9_), 
        .S(N154) );
  ADDFX2 U343 ( .A(n59), .B(n61), .CI(add_84_carry_9_), .CO(add_84_carry_10_), 
        .S(N155) );
  ADDFX2 U344 ( .A(n60), .B(n62), .CI(add_84_carry_10_), .CO(add_84_carry_11_), 
        .S(N156) );
  ADDFX2 U345 ( .A(n61), .B(n63), .CI(add_84_carry_11_), .CO(add_84_carry_12_), 
        .S(N157) );
  ADDFX2 U346 ( .A(n62), .B(n64), .CI(add_84_carry_12_), .CO(add_84_carry_13_), 
        .S(N158) );
  ADDFX2 U347 ( .A(n63), .B(n65), .CI(add_84_carry_13_), .CO(add_84_carry_14_), 
        .S(N159) );
  ADDFX2 U348 ( .A(n64), .B(n66), .CI(add_84_carry_14_), .CO(add_84_carry_15_), 
        .S(N160) );
  ADDFX2 U349 ( .A(n65), .B(n67), .CI(add_84_carry_15_), .CO(add_84_carry_16_), 
        .S(N161) );
  ADDFX2 U350 ( .A(n66), .B(x5[15]), .CI(add_84_carry_16_), .CO(
        add_84_carry_17_), .S(N162) );
  ADDFX2 U351 ( .A(n68), .B(n70), .CI(add_75_carry_5_), .CO(add_75_carry_6_), 
        .S(N66) );
  ADDFX2 U352 ( .A(n69), .B(n71), .CI(add_75_carry_6_), .CO(add_75_carry_7_), 
        .S(N67) );
  ADDFX2 U353 ( .A(n70), .B(n72), .CI(add_75_carry_7_), .CO(add_75_carry_8_), 
        .S(N68) );
  ADDFX2 U354 ( .A(n71), .B(n73), .CI(add_75_carry_8_), .CO(add_75_carry_9_), 
        .S(N69) );
  ADDFX2 U355 ( .A(n72), .B(n74), .CI(add_75_carry_9_), .CO(add_75_carry_10_), 
        .S(N70) );
  ADDFX2 U356 ( .A(n73), .B(n75), .CI(add_75_carry_10_), .CO(add_75_carry_11_), 
        .S(N71) );
  ADDFX2 U357 ( .A(n74), .B(n76), .CI(add_75_carry_11_), .CO(add_75_carry_12_), 
        .S(N72) );
  ADDFX2 U358 ( .A(n75), .B(n77), .CI(add_75_carry_12_), .CO(add_75_carry_13_), 
        .S(N73) );
  ADDFX2 U359 ( .A(n76), .B(n78), .CI(add_75_carry_13_), .CO(add_75_carry_14_), 
        .S(N74) );
  ADDFX2 U360 ( .A(n77), .B(n79), .CI(add_75_carry_14_), .CO(add_75_carry_15_), 
        .S(N75) );
  ADDFX2 U361 ( .A(n78), .B(n80), .CI(add_75_carry_15_), .CO(add_75_carry_16_), 
        .S(N76) );
  ADDFX2 U362 ( .A(n79), .B(x4[15]), .CI(add_75_carry_16_), .CO(
        add_75_carry_17_), .S(N77) );
  ADDFX2 U363 ( .A(n2), .B(n3), .CI(add_100_carry_6_), .CO(add_100_carry_7_), 
        .S(N301) );
  ADDFX2 U364 ( .A(n3), .B(n4), .CI(add_100_carry_7_), .CO(add_100_carry_8_), 
        .S(N302) );
  ADDFX2 U365 ( .A(n4), .B(n5), .CI(add_100_carry_8_), .CO(add_100_carry_9_), 
        .S(N303) );
  ADDFX2 U366 ( .A(n5), .B(n6), .CI(add_100_carry_9_), .CO(add_100_carry_10_), 
        .S(N304) );
  ADDFX2 U367 ( .A(n6), .B(n7), .CI(add_100_carry_10_), .CO(add_100_carry_11_), 
        .S(N305) );
  ADDFX2 U368 ( .A(n7), .B(n8), .CI(add_100_carry_11_), .CO(add_100_carry_12_), 
        .S(N306) );
  ADDFX2 U369 ( .A(n8), .B(n36), .CI(add_100_carry_12_), .CO(add_100_carry_13_), .S(N307) );
  ADDFX2 U370 ( .A(n36), .B(n37), .CI(add_100_carry_13_), .CO(
        add_100_carry_14_), .S(N308) );
  ADDFX2 U371 ( .A(n37), .B(n38), .CI(add_100_carry_14_), .CO(
        add_100_carry_15_), .S(N309) );
  ADDFX2 U372 ( .A(n38), .B(n39), .CI(add_100_carry_15_), .CO(
        add_100_carry_16_), .S(N310) );
  ADDFX2 U373 ( .A(n39), .B(n40), .CI(add_100_carry_16_), .CO(
        add_100_carry_17_), .S(N311) );
  ADDFX2 U374 ( .A(n40), .B(n41), .CI(add_100_carry_17_), .CO(
        add_100_carry_18_), .S(N312) );
  ADDFX2 U375 ( .A(n68), .B(n74), .CI(add_72_carry_8_), .CO(add_72_carry_9_), 
        .S(N25) );
  ADDFX2 U376 ( .A(n69), .B(n75), .CI(add_72_carry_9_), .CO(add_72_carry_10_), 
        .S(N26) );
  ADDFX2 U377 ( .A(n70), .B(n76), .CI(add_72_carry_10_), .CO(add_72_carry_11_), 
        .S(N27) );
  ADDFX2 U378 ( .A(n71), .B(n77), .CI(add_72_carry_11_), .CO(add_72_carry_12_), 
        .S(N28) );
  ADDFX2 U379 ( .A(n72), .B(n78), .CI(add_72_carry_12_), .CO(add_72_carry_13_), 
        .S(N29) );
  ADDFX2 U380 ( .A(n73), .B(n79), .CI(add_72_carry_13_), .CO(add_72_carry_14_), 
        .S(N30) );
  ADDFX2 U381 ( .A(n74), .B(n80), .CI(add_72_carry_14_), .CO(add_72_carry_15_), 
        .S(N31) );
  ADDFX2 U382 ( .A(n75), .B(x4[15]), .CI(add_72_carry_15_), .CO(
        add_72_carry_16_), .S(N32) );
  ADDFX2 U383 ( .A(n76), .B(x4[15]), .CI(add_72_carry_16_), .CO(
        add_72_carry_17_), .S(N33) );
  ADDFX2 U384 ( .A(n77), .B(x4[15]), .CI(add_72_carry_17_), .CO(
        add_72_carry_18_), .S(N34) );
  ADDFX2 U385 ( .A(n78), .B(x4[15]), .CI(add_72_carry_18_), .CO(
        add_72_carry_19_), .S(N35) );
  ADDFX2 U386 ( .A(n79), .B(x4[15]), .CI(add_72_carry_19_), .CO(
        add_72_carry_20_), .S(N36) );
  ADDFX2 U387 ( .A(n68), .B(n69), .CI(add_73_carry_6_), .CO(add_73_carry_7_), 
        .S(N46) );
  ADDFX2 U388 ( .A(n69), .B(n70), .CI(add_73_carry_7_), .CO(add_73_carry_8_), 
        .S(N47) );
  ADDFX2 U389 ( .A(n70), .B(n71), .CI(add_73_carry_8_), .CO(add_73_carry_9_), 
        .S(N48) );
  ADDFX2 U390 ( .A(n71), .B(n72), .CI(add_73_carry_9_), .CO(add_73_carry_10_), 
        .S(N49) );
  ADDFX2 U391 ( .A(n72), .B(n73), .CI(add_73_carry_10_), .CO(add_73_carry_11_), 
        .S(N50) );
  ADDFX2 U392 ( .A(n73), .B(n74), .CI(add_73_carry_11_), .CO(add_73_carry_12_), 
        .S(N51) );
  ADDFX2 U393 ( .A(n74), .B(n75), .CI(add_73_carry_12_), .CO(add_73_carry_13_), 
        .S(N52) );
  ADDFX2 U394 ( .A(n75), .B(n76), .CI(add_73_carry_13_), .CO(add_73_carry_14_), 
        .S(N53) );
  ADDFX2 U395 ( .A(n76), .B(n77), .CI(add_73_carry_14_), .CO(add_73_carry_15_), 
        .S(N54) );
  ADDFX2 U396 ( .A(n77), .B(n78), .CI(add_73_carry_15_), .CO(add_73_carry_16_), 
        .S(N55) );
  ADDFX2 U397 ( .A(n78), .B(n79), .CI(add_73_carry_16_), .CO(add_73_carry_17_), 
        .S(N56) );
  ADDFX2 U398 ( .A(n79), .B(n80), .CI(add_73_carry_17_), .CO(add_73_carry_18_), 
        .S(N57) );
  ADDFX2 U399 ( .A(n55), .B(n56), .CI(add_82_carry_6_), .CO(add_82_carry_7_), 
        .S(N131) );
  ADDFX2 U400 ( .A(n56), .B(n57), .CI(add_82_carry_7_), .CO(add_82_carry_8_), 
        .S(N132) );
  ADDFX2 U401 ( .A(n57), .B(n58), .CI(add_82_carry_8_), .CO(add_82_carry_9_), 
        .S(N133) );
  ADDFX2 U402 ( .A(n58), .B(n59), .CI(add_82_carry_9_), .CO(add_82_carry_10_), 
        .S(N134) );
  ADDFX2 U403 ( .A(n59), .B(n60), .CI(add_82_carry_10_), .CO(add_82_carry_11_), 
        .S(N135) );
  ADDFX2 U404 ( .A(n60), .B(n61), .CI(add_82_carry_11_), .CO(add_82_carry_12_), 
        .S(N136) );
  ADDFX2 U405 ( .A(n61), .B(n62), .CI(add_82_carry_12_), .CO(add_82_carry_13_), 
        .S(N137) );
  ADDFX2 U406 ( .A(n62), .B(n63), .CI(add_82_carry_13_), .CO(add_82_carry_14_), 
        .S(N138) );
  ADDFX2 U407 ( .A(n63), .B(n64), .CI(add_82_carry_14_), .CO(add_82_carry_15_), 
        .S(N139) );
  ADDFX2 U408 ( .A(n64), .B(n65), .CI(add_82_carry_15_), .CO(add_82_carry_16_), 
        .S(N140) );
  ADDFX2 U409 ( .A(n65), .B(n66), .CI(add_82_carry_16_), .CO(add_82_carry_17_), 
        .S(N141) );
  ADDFX2 U410 ( .A(n66), .B(n67), .CI(add_82_carry_17_), .CO(add_82_carry_18_), 
        .S(N142) );
  ADDFX2 U411 ( .A(n42), .B(n43), .CI(add_91_carry_6_), .CO(add_91_carry_7_), 
        .S(N216) );
  ADDFX2 U412 ( .A(n43), .B(n44), .CI(add_91_carry_7_), .CO(add_91_carry_8_), 
        .S(N217) );
  ADDFX2 U413 ( .A(n44), .B(n45), .CI(add_91_carry_8_), .CO(add_91_carry_9_), 
        .S(N218) );
  ADDFX2 U414 ( .A(n45), .B(n46), .CI(add_91_carry_9_), .CO(add_91_carry_10_), 
        .S(N219) );
  ADDFX2 U415 ( .A(n46), .B(n47), .CI(add_91_carry_10_), .CO(add_91_carry_11_), 
        .S(N220) );
  ADDFX2 U416 ( .A(n47), .B(n48), .CI(add_91_carry_11_), .CO(add_91_carry_12_), 
        .S(N221) );
  ADDFX2 U417 ( .A(n48), .B(n49), .CI(add_91_carry_12_), .CO(add_91_carry_13_), 
        .S(N222) );
  ADDFX2 U418 ( .A(n49), .B(n50), .CI(add_91_carry_13_), .CO(add_91_carry_14_), 
        .S(N223) );
  ADDFX2 U419 ( .A(n50), .B(n51), .CI(add_91_carry_14_), .CO(add_91_carry_15_), 
        .S(N224) );
  ADDFX2 U420 ( .A(n51), .B(n52), .CI(add_91_carry_15_), .CO(add_91_carry_16_), 
        .S(N225) );
  ADDFX2 U421 ( .A(n52), .B(n53), .CI(add_91_carry_16_), .CO(add_91_carry_17_), 
        .S(N226) );
  ADDFX2 U422 ( .A(n53), .B(n54), .CI(add_91_carry_17_), .CO(add_91_carry_18_), 
        .S(N227) );
  ADDFX2 U423 ( .A(n55), .B(n61), .CI(add_81_carry_8_), .CO(add_81_carry_9_), 
        .S(N110) );
  ADDFX2 U424 ( .A(n56), .B(n62), .CI(add_81_carry_9_), .CO(add_81_carry_10_), 
        .S(N111) );
  ADDFX2 U425 ( .A(n57), .B(n63), .CI(add_81_carry_10_), .CO(add_81_carry_11_), 
        .S(N112) );
  ADDFX2 U426 ( .A(n58), .B(n64), .CI(add_81_carry_11_), .CO(add_81_carry_12_), 
        .S(N113) );
  ADDFX2 U427 ( .A(n59), .B(n65), .CI(add_81_carry_12_), .CO(add_81_carry_13_), 
        .S(N114) );
  ADDFX2 U428 ( .A(n60), .B(n66), .CI(add_81_carry_13_), .CO(add_81_carry_14_), 
        .S(N115) );
  ADDFX2 U429 ( .A(n61), .B(n67), .CI(add_81_carry_14_), .CO(add_81_carry_15_), 
        .S(N116) );
  ADDFX2 U430 ( .A(n62), .B(x5[15]), .CI(add_81_carry_15_), .CO(
        add_81_carry_16_), .S(N117) );
  ADDFX2 U431 ( .A(n63), .B(x5[15]), .CI(add_81_carry_16_), .CO(
        add_81_carry_17_), .S(N118) );
  ADDFX2 U432 ( .A(n64), .B(x5[15]), .CI(add_81_carry_17_), .CO(
        add_81_carry_18_), .S(N119) );
  ADDFX2 U433 ( .A(n65), .B(x5[15]), .CI(add_81_carry_18_), .CO(
        add_81_carry_19_), .S(N120) );
  ADDFX2 U434 ( .A(n66), .B(x5[15]), .CI(add_81_carry_19_), .CO(
        add_81_carry_20_), .S(N121) );
  ADDFX2 U435 ( .A(n42), .B(n48), .CI(add_90_carry_8_), .CO(add_90_carry_9_), 
        .S(N195) );
  ADDFX2 U436 ( .A(n43), .B(n49), .CI(add_90_carry_9_), .CO(add_90_carry_10_), 
        .S(N196) );
  ADDFX2 U437 ( .A(n44), .B(n50), .CI(add_90_carry_10_), .CO(add_90_carry_11_), 
        .S(N197) );
  ADDFX2 U438 ( .A(n45), .B(n51), .CI(add_90_carry_11_), .CO(add_90_carry_12_), 
        .S(N198) );
  ADDFX2 U439 ( .A(n46), .B(n52), .CI(add_90_carry_12_), .CO(add_90_carry_13_), 
        .S(N199) );
  ADDFX2 U440 ( .A(n47), .B(n53), .CI(add_90_carry_13_), .CO(add_90_carry_14_), 
        .S(N200) );
  ADDFX2 U441 ( .A(n48), .B(n54), .CI(add_90_carry_14_), .CO(add_90_carry_15_), 
        .S(N201) );
  ADDFX2 U442 ( .A(n49), .B(x6[15]), .CI(add_90_carry_15_), .CO(
        add_90_carry_16_), .S(N202) );
  ADDFX2 U443 ( .A(n50), .B(x6[15]), .CI(add_90_carry_16_), .CO(
        add_90_carry_17_), .S(N203) );
  ADDFX2 U444 ( .A(n51), .B(x6[15]), .CI(add_90_carry_17_), .CO(
        add_90_carry_18_), .S(N204) );
  ADDFX2 U445 ( .A(n52), .B(x6[15]), .CI(add_90_carry_18_), .CO(
        add_90_carry_19_), .S(N205) );
  ADDFX2 U446 ( .A(n53), .B(x6[15]), .CI(add_90_carry_19_), .CO(
        add_90_carry_20_), .S(N206) );
  ADDFX2 U447 ( .A(n2), .B(n8), .CI(add_99_carry_8_), .CO(add_99_carry_9_), 
        .S(N280) );
  ADDFX2 U448 ( .A(n3), .B(n36), .CI(add_99_carry_9_), .CO(add_99_carry_10_), 
        .S(N281) );
  ADDFX2 U449 ( .A(n4), .B(n37), .CI(add_99_carry_10_), .CO(add_99_carry_11_), 
        .S(N282) );
  ADDFX2 U450 ( .A(n5), .B(n38), .CI(add_99_carry_11_), .CO(add_99_carry_12_), 
        .S(N283) );
  ADDFX2 U451 ( .A(n6), .B(n39), .CI(add_99_carry_12_), .CO(add_99_carry_13_), 
        .S(N284) );
  ADDFX2 U452 ( .A(n7), .B(n40), .CI(add_99_carry_13_), .CO(add_99_carry_14_), 
        .S(N285) );
  ADDFX2 U453 ( .A(n8), .B(n41), .CI(add_99_carry_14_), .CO(add_99_carry_15_), 
        .S(N286) );
  ADDFX2 U454 ( .A(n36), .B(x7[15]), .CI(add_99_carry_15_), .CO(
        add_99_carry_16_), .S(N287) );
  ADDFX2 U455 ( .A(n37), .B(x7[15]), .CI(add_99_carry_16_), .CO(
        add_99_carry_17_), .S(N288) );
  ADDFX2 U456 ( .A(n38), .B(x7[15]), .CI(add_99_carry_17_), .CO(
        add_99_carry_18_), .S(N289) );
  ADDFX2 U457 ( .A(n39), .B(x7[15]), .CI(add_99_carry_18_), .CO(
        add_99_carry_19_), .S(N290) );
  ADDFX2 U458 ( .A(n40), .B(x7[15]), .CI(add_99_carry_19_), .CO(
        add_99_carry_20_), .S(N291) );
  INVX1 U459 ( .A(n454), .Y(n182) );
  INVX1 U460 ( .A(n454), .Y(n180) );
  INVX1 U461 ( .A(n454), .Y(n181) );
  INVX1 U462 ( .A(n454), .Y(n179) );
  INVX1 U463 ( .A(n454), .Y(n178) );
  INVX1 U464 ( .A(n454), .Y(n177) );
  INVX1 U465 ( .A(n582), .Y(y0[16]) );
  INVX1 U466 ( .A(n565), .Y(y1[16]) );
  INVX1 U467 ( .A(n548), .Y(y2[16]) );
  INVX1 U468 ( .A(n531), .Y(y3[16]) );
  INVX1 U469 ( .A(n514), .Y(y4[16]) );
  INVX1 U470 ( .A(n497), .Y(y5[16]) );
  INVX1 U471 ( .A(n480), .Y(y6[16]) );
  INVX1 U472 ( .A(n463), .Y(y7[16]) );
  INVX1 U473 ( .A(x5_tmp[2]), .Y(n323) );
  INVX1 U474 ( .A(x5_tmp[3]), .Y(n322) );
  INVX1 U475 ( .A(x5_tmp[4]), .Y(n321) );
  INVX1 U476 ( .A(x5_tmp[5]), .Y(n320) );
  INVX1 U477 ( .A(x5_tmp[6]), .Y(n319) );
  INVX1 U478 ( .A(x5_tmp[7]), .Y(n318) );
  INVX1 U479 ( .A(x5_tmp[8]), .Y(n317) );
  INVX1 U480 ( .A(x5_tmp[9]), .Y(n316) );
  INVX1 U481 ( .A(x5_tmp[10]), .Y(n315) );
  INVX1 U482 ( .A(x5_tmp[11]), .Y(n314) );
  INVX1 U483 ( .A(x5_tmp[12]), .Y(n313) );
  INVX1 U484 ( .A(x5_tmp[13]), .Y(n312) );
  INVX1 U485 ( .A(x5_tmp[14]), .Y(n311) );
  INVX1 U486 ( .A(x5_tmp[15]), .Y(n310) );
  INVX1 U487 ( .A(x5_tmp[16]), .Y(n309) );
  INVX1 U488 ( .A(x5_tmp[17]), .Y(n308) );
  INVX1 U489 ( .A(x5_tmp[18]), .Y(n307) );
  INVX1 U490 ( .A(x5_tmp[19]), .Y(n306) );
  INVX1 U491 ( .A(x5_tmp[20]), .Y(n305) );
  INVX1 U492 ( .A(x5_tmp[21]), .Y(n304) );
  INVX1 U493 ( .A(x5_tmp[22]), .Y(n303) );
  INVX1 U494 ( .A(x5_tmp[23]), .Y(n302) );
  INVX1 U495 ( .A(x4_tmp[2]), .Y(n353) );
  INVX1 U496 ( .A(x4_tmp[3]), .Y(n354) );
  INVX1 U497 ( .A(x4_tmp[4]), .Y(n355) );
  INVX1 U498 ( .A(x4_tmp[5]), .Y(n356) );
  INVX1 U499 ( .A(x4_tmp[6]), .Y(n357) );
  INVX1 U500 ( .A(x4_tmp[7]), .Y(n358) );
  INVX1 U501 ( .A(x4_tmp[8]), .Y(n359) );
  INVX1 U502 ( .A(x4_tmp[9]), .Y(n360) );
  INVX1 U503 ( .A(x4_tmp[10]), .Y(n361) );
  INVX1 U504 ( .A(x4_tmp[11]), .Y(n362) );
  INVX1 U505 ( .A(x4_tmp[12]), .Y(n363) );
  INVX1 U506 ( .A(x4_tmp[13]), .Y(n364) );
  INVX1 U507 ( .A(x4_tmp[14]), .Y(n365) );
  INVX1 U508 ( .A(x4_tmp[15]), .Y(n366) );
  INVX1 U509 ( .A(x4_tmp[16]), .Y(n367) );
  INVX1 U510 ( .A(x4_tmp[17]), .Y(n368) );
  INVX1 U511 ( .A(x4_tmp[18]), .Y(n369) );
  INVX1 U512 ( .A(x4_tmp[19]), .Y(n370) );
  INVX1 U513 ( .A(x4_tmp[20]), .Y(n371) );
  INVX1 U514 ( .A(x4_tmp[21]), .Y(n372) );
  INVX1 U515 ( .A(x4_tmp[22]), .Y(n373) );
  INVX1 U516 ( .A(x4_tmp[23]), .Y(n374) );
  INVX1 U517 ( .A(x7_tmp[2]), .Y(n278) );
  INVX1 U518 ( .A(x7_tmp[3]), .Y(n279) );
  INVX1 U519 ( .A(x7_tmp[4]), .Y(n280) );
  INVX1 U520 ( .A(x7_tmp[5]), .Y(n281) );
  INVX1 U521 ( .A(x7_tmp[6]), .Y(n282) );
  INVX1 U522 ( .A(x7_tmp[7]), .Y(n283) );
  INVX1 U523 ( .A(x7_tmp[8]), .Y(n284) );
  INVX1 U524 ( .A(x7_tmp[9]), .Y(n285) );
  INVX1 U525 ( .A(x7_tmp[10]), .Y(n286) );
  INVX1 U526 ( .A(x7_tmp[11]), .Y(n287) );
  INVX1 U527 ( .A(x7_tmp[12]), .Y(n288) );
  INVX1 U528 ( .A(x7_tmp[13]), .Y(n289) );
  INVX1 U529 ( .A(x7_tmp[14]), .Y(n290) );
  INVX1 U530 ( .A(x7_tmp[15]), .Y(n291) );
  INVX1 U531 ( .A(x7_tmp[16]), .Y(n292) );
  INVX1 U532 ( .A(x7_tmp[17]), .Y(n293) );
  INVX1 U533 ( .A(x7_tmp[18]), .Y(n294) );
  INVX1 U534 ( .A(x7_tmp[19]), .Y(n295) );
  INVX1 U535 ( .A(x7_tmp[20]), .Y(n296) );
  INVX1 U536 ( .A(x7_tmp[21]), .Y(n297) );
  INVX1 U537 ( .A(x7_tmp[22]), .Y(n298) );
  INVX1 U538 ( .A(x7_tmp[23]), .Y(n299) );
  INVX1 U539 ( .A(x6_tmp[2]), .Y(n348) );
  INVX1 U540 ( .A(x6_tmp[3]), .Y(n347) );
  INVX1 U541 ( .A(x6_tmp[4]), .Y(n346) );
  INVX1 U542 ( .A(x6_tmp[5]), .Y(n345) );
  INVX1 U543 ( .A(x6_tmp[6]), .Y(n344) );
  INVX1 U544 ( .A(x6_tmp[7]), .Y(n343) );
  INVX1 U545 ( .A(x6_tmp[8]), .Y(n342) );
  INVX1 U546 ( .A(x6_tmp[9]), .Y(n341) );
  INVX1 U547 ( .A(x6_tmp[10]), .Y(n340) );
  INVX1 U548 ( .A(x6_tmp[11]), .Y(n339) );
  INVX1 U549 ( .A(x6_tmp[12]), .Y(n338) );
  INVX1 U550 ( .A(x6_tmp[13]), .Y(n337) );
  INVX1 U551 ( .A(x6_tmp[14]), .Y(n336) );
  INVX1 U552 ( .A(x6_tmp[15]), .Y(n335) );
  INVX1 U553 ( .A(x6_tmp[16]), .Y(n334) );
  INVX1 U554 ( .A(x6_tmp[17]), .Y(n333) );
  INVX1 U555 ( .A(x6_tmp[18]), .Y(n332) );
  INVX1 U556 ( .A(x6_tmp[19]), .Y(n331) );
  INVX1 U557 ( .A(x6_tmp[20]), .Y(n330) );
  INVX1 U558 ( .A(x6_tmp[21]), .Y(n329) );
  INVX1 U559 ( .A(x6_tmp[22]), .Y(n328) );
  INVX1 U560 ( .A(x6_tmp[23]), .Y(n327) );
  INVX1 U561 ( .A(x5_tmp[1]), .Y(n324) );
  INVX1 U562 ( .A(x4_tmp[1]), .Y(n352) );
  INVX1 U563 ( .A(x7_tmp[1]), .Y(n277) );
  INVX1 U564 ( .A(x6_tmp[1]), .Y(n349) );
  INVX1 U565 ( .A(x5_tmp[0]), .Y(n325) );
  INVX1 U566 ( .A(x4_tmp[0]), .Y(n351) );
  INVX1 U567 ( .A(x7_tmp[0]), .Y(n276) );
  INVX1 U568 ( .A(x6_tmp[0]), .Y(n350) );
  INVX1 U569 ( .A(x7_89[0]), .Y(n253) );
  INVX1 U570 ( .A(x5_89[0]), .Y(n230) );
  INVX1 U571 ( .A(x7_50[0]), .Y(n207) );
  INVX1 U572 ( .A(x5_50[0]), .Y(n275) );
  INVX1 U573 ( .A(x7_89[2]), .Y(n251) );
  INVX1 U574 ( .A(x7_89[3]), .Y(n250) );
  INVX1 U575 ( .A(x7_89[4]), .Y(n249) );
  INVX1 U576 ( .A(x7_89[5]), .Y(n248) );
  INVX1 U577 ( .A(x7_89[6]), .Y(n247) );
  INVX1 U578 ( .A(x7_89[7]), .Y(n246) );
  INVX1 U579 ( .A(x7_89[8]), .Y(n245) );
  INVX1 U580 ( .A(x7_89[9]), .Y(n244) );
  INVX1 U581 ( .A(x7_89[10]), .Y(n243) );
  INVX1 U582 ( .A(x7_89[11]), .Y(n242) );
  INVX1 U583 ( .A(x7_89[12]), .Y(n241) );
  INVX1 U584 ( .A(x7_89[13]), .Y(n240) );
  INVX1 U585 ( .A(x7_89[14]), .Y(n239) );
  INVX1 U586 ( .A(x7_89[15]), .Y(n238) );
  INVX1 U587 ( .A(x7_89[16]), .Y(n237) );
  INVX1 U588 ( .A(x7_89[17]), .Y(n236) );
  INVX1 U589 ( .A(x7_89[18]), .Y(n235) );
  INVX1 U590 ( .A(x7_89[19]), .Y(n234) );
  INVX1 U591 ( .A(x7_89[20]), .Y(n233) );
  INVX1 U592 ( .A(x7_89[21]), .Y(n232) );
  INVX1 U593 ( .A(x5_89[2]), .Y(n228) );
  INVX1 U594 ( .A(x5_89[3]), .Y(n227) );
  INVX1 U595 ( .A(x5_89[4]), .Y(n226) );
  INVX1 U596 ( .A(x5_89[5]), .Y(n225) );
  INVX1 U597 ( .A(x5_89[6]), .Y(n224) );
  INVX1 U598 ( .A(x5_89[7]), .Y(n223) );
  INVX1 U599 ( .A(x5_89[8]), .Y(n222) );
  INVX1 U600 ( .A(x5_89[9]), .Y(n221) );
  INVX1 U601 ( .A(x5_89[10]), .Y(n220) );
  INVX1 U602 ( .A(x5_89[11]), .Y(n219) );
  INVX1 U603 ( .A(x5_89[12]), .Y(n218) );
  INVX1 U604 ( .A(x5_89[13]), .Y(n217) );
  INVX1 U605 ( .A(x5_89[14]), .Y(n216) );
  INVX1 U606 ( .A(x5_89[15]), .Y(n215) );
  INVX1 U607 ( .A(x5_89[16]), .Y(n214) );
  INVX1 U608 ( .A(x5_89[17]), .Y(n213) );
  INVX1 U609 ( .A(x5_89[18]), .Y(n212) );
  INVX1 U610 ( .A(x5_89[19]), .Y(n211) );
  INVX1 U611 ( .A(x5_89[20]), .Y(n210) );
  INVX1 U612 ( .A(x5_89[21]), .Y(n209) );
  INVX1 U613 ( .A(x7_50[2]), .Y(n205) );
  INVX1 U614 ( .A(x7_50[3]), .Y(n204) );
  INVX1 U615 ( .A(x7_50[4]), .Y(n203) );
  INVX1 U616 ( .A(x7_50[5]), .Y(n202) );
  INVX1 U617 ( .A(x7_50[6]), .Y(n201) );
  INVX1 U618 ( .A(x7_50[7]), .Y(n200) );
  INVX1 U619 ( .A(x7_50[8]), .Y(n199) );
  INVX1 U620 ( .A(x7_50[9]), .Y(n198) );
  INVX1 U621 ( .A(x7_50[10]), .Y(n197) );
  INVX1 U622 ( .A(x7_50[11]), .Y(n196) );
  INVX1 U623 ( .A(x7_50[12]), .Y(n195) );
  INVX1 U624 ( .A(x7_50[13]), .Y(n194) );
  INVX1 U625 ( .A(x7_50[14]), .Y(n193) );
  INVX1 U626 ( .A(x7_50[15]), .Y(n192) );
  INVX1 U627 ( .A(x7_50[16]), .Y(n191) );
  INVX1 U628 ( .A(x7_50[17]), .Y(n190) );
  INVX1 U629 ( .A(x7_50[18]), .Y(n189) );
  INVX1 U630 ( .A(x7_50[19]), .Y(n188) );
  INVX1 U631 ( .A(x7_50[20]), .Y(n187) );
  INVX1 U632 ( .A(x5_50[2]), .Y(n273) );
  INVX1 U633 ( .A(x5_50[3]), .Y(n272) );
  INVX1 U634 ( .A(x5_50[4]), .Y(n271) );
  INVX1 U635 ( .A(x5_50[5]), .Y(n270) );
  INVX1 U636 ( .A(x5_50[6]), .Y(n269) );
  INVX1 U637 ( .A(x5_50[7]), .Y(n268) );
  INVX1 U638 ( .A(x5_50[8]), .Y(n267) );
  INVX1 U639 ( .A(x5_50[9]), .Y(n266) );
  INVX1 U640 ( .A(x5_50[10]), .Y(n265) );
  INVX1 U641 ( .A(x5_50[11]), .Y(n264) );
  INVX1 U642 ( .A(x5_50[12]), .Y(n263) );
  INVX1 U643 ( .A(x5_50[13]), .Y(n262) );
  INVX1 U644 ( .A(x5_50[14]), .Y(n261) );
  INVX1 U645 ( .A(x5_50[15]), .Y(n260) );
  INVX1 U646 ( .A(x5_50[16]), .Y(n259) );
  INVX1 U647 ( .A(x5_50[17]), .Y(n258) );
  INVX1 U648 ( .A(x5_50[18]), .Y(n257) );
  INVX1 U649 ( .A(x5_50[19]), .Y(n256) );
  INVX1 U650 ( .A(x5_50[20]), .Y(n255) );
  INVX1 U651 ( .A(x7_50[1]), .Y(n206) );
  INVX1 U652 ( .A(x5_50[1]), .Y(n274) );
  INVX1 U653 ( .A(x7_89[1]), .Y(n252) );
  INVX1 U654 ( .A(x5_89[1]), .Y(n229) );
  AOI22X1 U655 ( .A0(N1710), .A1(n123), .B0(y4_tmp[15]), .B1(n86), .Y(n515) );
  AOI22X1 U656 ( .A0(N1727), .A1(n115), .B0(y5_tmp[15]), .B1(n84), .Y(n498) );
  AOI22X1 U657 ( .A0(N1744), .A1(n106), .B0(y6_tmp[15]), .B1(n83), .Y(n481) );
  AOI22X1 U658 ( .A0(N1761), .A1(n98), .B0(y7_tmp[15]), .B1(n81), .Y(n464) );
  INVX1 U659 ( .A(n584), .Y(y0[14]) );
  AOI22X1 U660 ( .A0(N1641), .A1(n154), .B0(y0_tmp[14]), .B1(n88), .Y(n584) );
  INVX1 U661 ( .A(n583), .Y(y0[15]) );
  AOI22X1 U662 ( .A0(N1642), .A1(n153), .B0(y0_tmp[15]), .B1(n88), .Y(n583) );
  INVX1 U663 ( .A(n567), .Y(y1[14]) );
  AOI22X1 U664 ( .A0(N1658), .A1(n145), .B0(y1_tmp[14]), .B1(n89), .Y(n567) );
  INVX1 U665 ( .A(n566), .Y(y1[15]) );
  AOI22X1 U666 ( .A0(N1659), .A1(n145), .B0(y1_tmp[15]), .B1(n89), .Y(n566) );
  INVX1 U667 ( .A(n550), .Y(y2[14]) );
  AOI22X1 U668 ( .A0(N1675), .A1(n139), .B0(y2_tmp[14]), .B1(n90), .Y(n550) );
  INVX1 U669 ( .A(n549), .Y(y2[15]) );
  AOI22X1 U670 ( .A0(N1676), .A1(n138), .B0(y2_tmp[15]), .B1(n91), .Y(n549) );
  INVX1 U671 ( .A(n533), .Y(y3[14]) );
  AOI22X1 U672 ( .A0(N1692), .A1(n130), .B0(y3_tmp[14]), .B1(n87), .Y(n533) );
  INVX1 U673 ( .A(n532), .Y(y3[15]) );
  AOI22X1 U674 ( .A0(N1693), .A1(n130), .B0(y3_tmp[15]), .B1(n87), .Y(n532) );
  INVX1 U675 ( .A(n515), .Y(y4[15]) );
  INVX1 U676 ( .A(n498), .Y(y5[15]) );
  INVX1 U677 ( .A(n481), .Y(y6[15]) );
  INVX1 U678 ( .A(n464), .Y(y7[15]) );
  INVX1 U679 ( .A(n585), .Y(y0[13]) );
  AOI22X1 U680 ( .A0(N1640), .A1(n154), .B0(y0_tmp[13]), .B1(n88), .Y(n585) );
  INVX1 U681 ( .A(n568), .Y(y1[13]) );
  AOI22X1 U682 ( .A0(N1657), .A1(n146), .B0(y1_tmp[13]), .B1(n89), .Y(n568) );
  INVX1 U683 ( .A(n551), .Y(y2[13]) );
  AOI22X1 U684 ( .A0(N1674), .A1(n139), .B0(y2_tmp[13]), .B1(n90), .Y(n551) );
  INVX1 U685 ( .A(n534), .Y(y3[13]) );
  AOI22X1 U686 ( .A0(N1691), .A1(n131), .B0(y3_tmp[13]), .B1(n87), .Y(n534) );
  AOI22X1 U687 ( .A0(N1708), .A1(n124), .B0(y4_tmp[13]), .B1(n86), .Y(n517) );
  AOI22X1 U688 ( .A0(N1709), .A1(n124), .B0(y4_tmp[14]), .B1(n86), .Y(n516) );
  AOI22X1 U689 ( .A0(N1725), .A1(n116), .B0(y5_tmp[13]), .B1(n84), .Y(n500) );
  AOI22X1 U690 ( .A0(N1726), .A1(n115), .B0(y5_tmp[14]), .B1(n84), .Y(n499) );
  AOI22X1 U691 ( .A0(N1742), .A1(n107), .B0(y6_tmp[13]), .B1(n83), .Y(n483) );
  AOI22X1 U692 ( .A0(N1743), .A1(n107), .B0(y6_tmp[14]), .B1(n83), .Y(n482) );
  AOI22X1 U693 ( .A0(N1759), .A1(n99), .B0(y7_tmp[13]), .B1(n82), .Y(n466) );
  AOI22X1 U694 ( .A0(N1760), .A1(n98), .B0(y7_tmp[14]), .B1(n81), .Y(n465) );
  AOI22X1 U695 ( .A0(N1705), .A1(n126), .B0(y4_tmp[10]), .B1(n86), .Y(n520) );
  AOI22X1 U696 ( .A0(N1722), .A1(n117), .B0(y5_tmp[10]), .B1(n85), .Y(n503) );
  AOI22X1 U697 ( .A0(N1739), .A1(n109), .B0(y6_tmp[10]), .B1(n83), .Y(n486) );
  AOI22X1 U698 ( .A0(N1756), .A1(n100), .B0(y7_tmp[10]), .B1(n82), .Y(n469) );
  AOI22X1 U699 ( .A0(N1706), .A1(n125), .B0(y4_tmp[11]), .B1(n86), .Y(n519) );
  AOI22X1 U700 ( .A0(N1707), .A1(n125), .B0(y4_tmp[12]), .B1(n86), .Y(n518) );
  AOI22X1 U701 ( .A0(N1723), .A1(n117), .B0(y5_tmp[11]), .B1(n85), .Y(n502) );
  AOI22X1 U702 ( .A0(N1724), .A1(n116), .B0(y5_tmp[12]), .B1(n84), .Y(n501) );
  AOI22X1 U703 ( .A0(N1740), .A1(n108), .B0(y6_tmp[11]), .B1(n83), .Y(n485) );
  AOI22X1 U704 ( .A0(N1741), .A1(n108), .B0(y6_tmp[12]), .B1(n83), .Y(n484) );
  AOI22X1 U705 ( .A0(N1757), .A1(n100), .B0(y7_tmp[11]), .B1(n82), .Y(n468) );
  AOI22X1 U706 ( .A0(N1758), .A1(n99), .B0(y7_tmp[12]), .B1(n82), .Y(n467) );
  INVX1 U707 ( .A(n574), .Y(y0[8]) );
  AOI22X1 U708 ( .A0(N1635), .A1(n149), .B0(y0_tmp[8]), .B1(n88), .Y(n574) );
  INVX1 U709 ( .A(n573), .Y(y0[9]) );
  AOI22X1 U710 ( .A0(N1636), .A1(n148), .B0(y0_tmp[9]), .B1(n89), .Y(n573) );
  INVX1 U711 ( .A(n557), .Y(y1[8]) );
  AOI22X1 U712 ( .A0(N1652), .A1(n141), .B0(y1_tmp[8]), .B1(n90), .Y(n557) );
  INVX1 U713 ( .A(n556), .Y(y1[9]) );
  AOI22X1 U714 ( .A0(N1653), .A1(n141), .B0(y1_tmp[9]), .B1(n90), .Y(n556) );
  INVX1 U715 ( .A(n540), .Y(y2[8]) );
  AOI22X1 U716 ( .A0(N1669), .A1(n134), .B0(y2_tmp[8]), .B1(n92), .Y(n540) );
  INVX1 U717 ( .A(n539), .Y(y2[9]) );
  AOI22X1 U718 ( .A0(N1670), .A1(n133), .B0(y2_tmp[9]), .B1(n92), .Y(n539) );
  INVX1 U719 ( .A(n466), .Y(y7[13]) );
  INVX1 U720 ( .A(n523), .Y(y3[8]) );
  AOI22X1 U721 ( .A0(N1686), .A1(n127), .B0(y3_tmp[8]), .B1(n86), .Y(n523) );
  INVX1 U722 ( .A(n522), .Y(y3[9]) );
  AOI22X1 U723 ( .A0(N1687), .A1(n127), .B0(y3_tmp[9]), .B1(n86), .Y(n522) );
  INVX1 U724 ( .A(n519), .Y(y4[11]) );
  INVX1 U725 ( .A(n518), .Y(y4[12]) );
  INVX1 U726 ( .A(n516), .Y(y4[14]) );
  INVX1 U727 ( .A(n502), .Y(y5[11]) );
  INVX1 U728 ( .A(n501), .Y(y5[12]) );
  INVX1 U729 ( .A(n499), .Y(y5[14]) );
  INVX1 U730 ( .A(n485), .Y(y6[11]) );
  INVX1 U731 ( .A(n484), .Y(y6[12]) );
  INVX1 U732 ( .A(n482), .Y(y6[14]) );
  ADDFX2 U733 ( .A(x4[1]), .B(n73), .CI(add_72_carry_7_), .CO(add_72_carry_8_), 
        .S(N24) );
  ADDFX2 U734 ( .A(x5[1]), .B(n60), .CI(add_81_carry_7_), .CO(add_81_carry_8_), 
        .S(N109) );
  ADDFX2 U735 ( .A(x6[1]), .B(n47), .CI(add_90_carry_7_), .CO(add_90_carry_8_), 
        .S(N194) );
  BUFX3 U736 ( .A(x5[7]), .Y(n60) );
  BUFX3 U737 ( .A(x5[8]), .Y(n61) );
  BUFX3 U738 ( .A(x6[7]), .Y(n47) );
  BUFX3 U739 ( .A(x6[8]), .Y(n48) );
  BUFX3 U740 ( .A(x4[7]), .Y(n73) );
  BUFX3 U741 ( .A(x4[8]), .Y(n74) );
  BUFX3 U742 ( .A(x7[7]), .Y(n7) );
  BUFX3 U743 ( .A(x7[8]), .Y(n8) );
  BUFX3 U744 ( .A(x4[4]), .Y(n70) );
  BUFX3 U745 ( .A(x4[5]), .Y(n71) );
  BUFX3 U746 ( .A(x5[4]), .Y(n57) );
  BUFX3 U747 ( .A(x5[5]), .Y(n58) );
  BUFX3 U748 ( .A(x6[4]), .Y(n44) );
  BUFX3 U749 ( .A(x6[5]), .Y(n45) );
  BUFX3 U750 ( .A(x5[6]), .Y(n59) );
  BUFX3 U751 ( .A(x6[6]), .Y(n46) );
  BUFX3 U752 ( .A(x4[6]), .Y(n72) );
  BUFX3 U753 ( .A(x7[4]), .Y(n4) );
  BUFX3 U754 ( .A(x7[5]), .Y(n5) );
  BUFX3 U755 ( .A(x7[6]), .Y(n6) );
  INVX1 U756 ( .A(n469), .Y(y7[10]) );
  INVX1 U757 ( .A(n468), .Y(y7[11]) );
  INVX1 U758 ( .A(n467), .Y(y7[12]) );
  INVX1 U759 ( .A(n465), .Y(y7[14]) );
  INVX1 U760 ( .A(n588), .Y(y0[10]) );
  AOI22X1 U761 ( .A0(N1637), .A1(n155), .B0(y0_tmp[10]), .B1(n91), .Y(n588) );
  INVX1 U762 ( .A(n587), .Y(y0[11]) );
  AOI22X1 U763 ( .A0(N1638), .A1(n155), .B0(y0_tmp[11]), .B1(n87), .Y(n587) );
  INVX1 U764 ( .A(n586), .Y(y0[12]) );
  AOI22X1 U765 ( .A0(N1639), .A1(n155), .B0(y0_tmp[12]), .B1(n87), .Y(n586) );
  INVX1 U766 ( .A(n571), .Y(y1[10]) );
  AOI22X1 U767 ( .A0(N1654), .A1(n147), .B0(y1_tmp[10]), .B1(n89), .Y(n571) );
  INVX1 U768 ( .A(n570), .Y(y1[11]) );
  AOI22X1 U769 ( .A0(N1655), .A1(n147), .B0(y1_tmp[11]), .B1(n89), .Y(n570) );
  INVX1 U770 ( .A(n569), .Y(y1[12]) );
  AOI22X1 U771 ( .A0(N1656), .A1(n146), .B0(y1_tmp[12]), .B1(n89), .Y(n569) );
  INVX1 U772 ( .A(n554), .Y(y2[10]) );
  AOI22X1 U773 ( .A0(N1671), .A1(n140), .B0(y2_tmp[10]), .B1(n90), .Y(n554) );
  INVX1 U774 ( .A(n553), .Y(y2[11]) );
  AOI22X1 U775 ( .A0(N1672), .A1(n140), .B0(y2_tmp[11]), .B1(n90), .Y(n553) );
  INVX1 U776 ( .A(n552), .Y(y2[12]) );
  AOI22X1 U777 ( .A0(N1673), .A1(n140), .B0(y2_tmp[12]), .B1(n90), .Y(n552) );
  INVX1 U778 ( .A(n537), .Y(y3[10]) );
  AOI22X1 U779 ( .A0(N1688), .A1(n132), .B0(y3_tmp[10]), .B1(n92), .Y(n537) );
  INVX1 U780 ( .A(n536), .Y(y3[11]) );
  AOI22X1 U781 ( .A0(N1689), .A1(n132), .B0(y3_tmp[11]), .B1(n92), .Y(n536) );
  INVX1 U782 ( .A(n535), .Y(y3[12]) );
  AOI22X1 U783 ( .A0(N1690), .A1(n131), .B0(y3_tmp[12]), .B1(n91), .Y(n535) );
  BUFX3 U784 ( .A(x4[3]), .Y(n69) );
  BUFX3 U785 ( .A(x5[3]), .Y(n56) );
  BUFX3 U786 ( .A(x6[3]), .Y(n43) );
  BUFX3 U787 ( .A(x7[3]), .Y(n3) );
  BUFX3 U788 ( .A(x4[2]), .Y(n68) );
  BUFX3 U789 ( .A(x5[2]), .Y(n55) );
  BUFX3 U790 ( .A(x6[2]), .Y(n42) );
  INVX1 U791 ( .A(n520), .Y(y4[10]) );
  INVX1 U792 ( .A(n517), .Y(y4[13]) );
  INVX1 U793 ( .A(n503), .Y(y5[10]) );
  INVX1 U794 ( .A(n500), .Y(y5[13]) );
  INVX1 U795 ( .A(n486), .Y(y6[10]) );
  INVX1 U796 ( .A(n483), .Y(y6[13]) );
  ADDFX2 U797 ( .A(x4[1]), .B(n68), .CI(add_73_carry_5_), .CO(add_73_carry_6_), 
        .S(N45) );
  ADDFX2 U798 ( .A(x5[1]), .B(n55), .CI(add_82_carry_5_), .CO(add_82_carry_6_), 
        .S(N130) );
  ADDFX2 U799 ( .A(x6[1]), .B(n42), .CI(add_91_carry_5_), .CO(add_91_carry_6_), 
        .S(N215) );
  ADDFX2 U800 ( .A(x7[1]), .B(n4), .CI(add_104_carry_5_), .CO(add_104_carry_6_), .S(N341) );
  ADDFX2 U801 ( .A(x5[1]), .B(n57), .CI(add_86_carry_5_), .CO(add_86_carry_6_), 
        .S(N171) );
  ADDFX2 U802 ( .A(x6[1]), .B(n44), .CI(add_95_carry_5_), .CO(add_95_carry_6_), 
        .S(N256) );
  ADDFX2 U803 ( .A(x4[1]), .B(n70), .CI(add_77_carry_5_), .CO(add_77_carry_6_), 
        .S(N86) );
  ADDFX2 U804 ( .A(x7[1]), .B(n3), .CI(add_102_carry_4_), .CO(add_102_carry_5_), .S(N320) );
  ADDFX2 U805 ( .A(x6[1]), .B(n43), .CI(add_93_carry_4_), .CO(add_93_carry_5_), 
        .S(N235) );
  ADDFX2 U806 ( .A(x5[1]), .B(n56), .CI(add_84_carry_4_), .CO(add_84_carry_5_), 
        .S(N150) );
  ADDFX2 U807 ( .A(x4[1]), .B(n69), .CI(add_75_carry_4_), .CO(add_75_carry_5_), 
        .S(N65) );
  ADDFX2 U808 ( .A(x7[1]), .B(n2), .CI(add_100_carry_5_), .CO(add_100_carry_6_), .S(N300) );
  ADDFX2 U809 ( .A(x7[1]), .B(n7), .CI(add_99_carry_7_), .CO(add_99_carry_8_), 
        .S(N279) );
  BUFX3 U810 ( .A(x7[2]), .Y(n2) );
  NAND2BX1 U811 ( .AN(mode_delay2[1]), .B(mode_delay2[0]), .Y(n454) );
  AOI22X1 U812 ( .A0(N1735), .A1(n103), .B0(y6_tmp[6]), .B1(n82), .Y(n474) );
  AOI22X1 U813 ( .A0(N1738), .A1(n101), .B0(y6_tmp[9]), .B1(n82), .Y(n471) );
  AOI22X1 U814 ( .A0(N1752), .A1(n94), .B0(y7_tmp[6]), .B1(n81), .Y(n457) );
  AOI22X1 U815 ( .A0(N1755), .A1(n93), .B0(y7_tmp[9]), .B1(n87), .Y(n453) );
  AOI22X1 U816 ( .A0(N1701), .A1(n120), .B0(y4_tmp[6]), .B1(n85), .Y(n508) );
  AOI22X1 U817 ( .A0(N1702), .A1(n119), .B0(y4_tmp[7]), .B1(n85), .Y(n507) );
  AOI22X1 U818 ( .A0(N1703), .A1(n119), .B0(y4_tmp[8]), .B1(n85), .Y(n506) );
  AOI22X1 U819 ( .A0(N1704), .A1(n118), .B0(y4_tmp[9]), .B1(n85), .Y(n505) );
  AOI22X1 U820 ( .A0(N1718), .A1(n111), .B0(y5_tmp[6]), .B1(n84), .Y(n491) );
  AOI22X1 U821 ( .A0(N1719), .A1(n111), .B0(y5_tmp[7]), .B1(n84), .Y(n490) );
  AOI22X1 U822 ( .A0(N1720), .A1(n110), .B0(y5_tmp[8]), .B1(n83), .Y(n489) );
  AOI22X1 U823 ( .A0(N1721), .A1(n110), .B0(y5_tmp[9]), .B1(n83), .Y(n488) );
  AOI22X1 U824 ( .A0(N1736), .A1(n102), .B0(y6_tmp[7]), .B1(n82), .Y(n473) );
  AOI22X1 U825 ( .A0(N1737), .A1(n102), .B0(y6_tmp[8]), .B1(n82), .Y(n472) );
  AOI22X1 U826 ( .A0(N1753), .A1(n94), .B0(y7_tmp[7]), .B1(n81), .Y(n456) );
  AOI22X1 U827 ( .A0(N1754), .A1(n93), .B0(y7_tmp[8]), .B1(n81), .Y(n455) );
  INVX1 U828 ( .A(n581), .Y(y0[1]) );
  AOI22X1 U829 ( .A0(N1628), .A1(n152), .B0(y0_tmp[1]), .B1(n88), .Y(n581) );
  INVX1 U830 ( .A(n580), .Y(y0[2]) );
  AOI22X1 U831 ( .A0(N1629), .A1(n152), .B0(y0_tmp[2]), .B1(n88), .Y(n580) );
  INVX1 U832 ( .A(n579), .Y(y0[3]) );
  AOI22X1 U833 ( .A0(N1630), .A1(n151), .B0(y0_tmp[3]), .B1(n88), .Y(n579) );
  INVX1 U834 ( .A(n577), .Y(y0[5]) );
  AOI22X1 U835 ( .A0(N1632), .A1(n150), .B0(y0_tmp[5]), .B1(n88), .Y(n577) );
  INVX1 U836 ( .A(n564), .Y(y1[1]) );
  AOI22X1 U837 ( .A0(N1645), .A1(n145), .B0(y1_tmp[1]), .B1(n89), .Y(n564) );
  INVX1 U838 ( .A(n563), .Y(y1[2]) );
  AOI22X1 U839 ( .A0(N1646), .A1(n144), .B0(y1_tmp[2]), .B1(n89), .Y(n563) );
  INVX1 U840 ( .A(n562), .Y(y1[3]) );
  AOI22X1 U841 ( .A0(N1647), .A1(n144), .B0(y1_tmp[3]), .B1(n89), .Y(n562) );
  INVX1 U842 ( .A(n560), .Y(y1[5]) );
  AOI22X1 U843 ( .A0(N1649), .A1(n143), .B0(y1_tmp[5]), .B1(n90), .Y(n560) );
  INVX1 U844 ( .A(n547), .Y(y2[1]) );
  AOI22X1 U845 ( .A0(N1662), .A1(n137), .B0(y2_tmp[1]), .B1(n91), .Y(n547) );
  INVX1 U846 ( .A(n546), .Y(y2[2]) );
  AOI22X1 U847 ( .A0(N1663), .A1(n137), .B0(y2_tmp[2]), .B1(n91), .Y(n546) );
  INVX1 U848 ( .A(n545), .Y(y2[3]) );
  AOI22X1 U849 ( .A0(N1664), .A1(n136), .B0(y2_tmp[3]), .B1(n91), .Y(n545) );
  INVX1 U850 ( .A(n543), .Y(y2[5]) );
  AOI22X1 U851 ( .A0(N1666), .A1(n135), .B0(y2_tmp[5]), .B1(n91), .Y(n543) );
  INVX1 U852 ( .A(n530), .Y(y3[1]) );
  AOI22X1 U853 ( .A0(N1679), .A1(n129), .B0(y3_tmp[1]), .B1(n87), .Y(n530) );
  INVX1 U854 ( .A(n529), .Y(y3[2]) );
  AOI22X1 U855 ( .A0(N1680), .A1(n129), .B0(y3_tmp[2]), .B1(n87), .Y(n529) );
  INVX1 U856 ( .A(n528), .Y(y3[3]) );
  AOI22X1 U857 ( .A0(N1681), .A1(n129), .B0(y3_tmp[3]), .B1(n87), .Y(n528) );
  INVX1 U858 ( .A(n526), .Y(y3[5]) );
  AOI22X1 U859 ( .A0(N1683), .A1(n128), .B0(y3_tmp[5]), .B1(n87), .Y(n526) );
  INVX1 U860 ( .A(n524), .Y(y3[7]) );
  AOI22X1 U861 ( .A0(N1685), .A1(n127), .B0(y3_tmp[7]), .B1(n86), .Y(n524) );
  BUFX3 U862 ( .A(x5[9]), .Y(n62) );
  BUFX3 U863 ( .A(x5[10]), .Y(n63) );
  BUFX3 U864 ( .A(x5[11]), .Y(n64) );
  BUFX3 U865 ( .A(x5[12]), .Y(n65) );
  BUFX3 U866 ( .A(x6[9]), .Y(n49) );
  BUFX3 U867 ( .A(x6[10]), .Y(n50) );
  BUFX3 U868 ( .A(x6[11]), .Y(n51) );
  BUFX3 U869 ( .A(x6[12]), .Y(n52) );
  BUFX3 U870 ( .A(x4[9]), .Y(n75) );
  BUFX3 U871 ( .A(x4[10]), .Y(n76) );
  BUFX3 U872 ( .A(x4[11]), .Y(n77) );
  BUFX3 U873 ( .A(x4[12]), .Y(n78) );
  BUFX3 U874 ( .A(x7[9]), .Y(n36) );
  BUFX3 U875 ( .A(x7[10]), .Y(n37) );
  BUFX3 U876 ( .A(x7[11]), .Y(n38) );
  BUFX3 U877 ( .A(x7[12]), .Y(n39) );
  INVX1 U878 ( .A(n589), .Y(y0[0]) );
  AOI22X1 U879 ( .A0(N1627), .A1(n155), .B0(y0_tmp[0]), .B1(n81), .Y(n589) );
  INVX1 U880 ( .A(n578), .Y(y0[4]) );
  AOI22X1 U881 ( .A0(N1631), .A1(n151), .B0(y0_tmp[4]), .B1(n88), .Y(n578) );
  INVX1 U882 ( .A(n576), .Y(y0[6]) );
  AOI22X1 U883 ( .A0(N1633), .A1(n150), .B0(y0_tmp[6]), .B1(n88), .Y(n576) );
  INVX1 U884 ( .A(n575), .Y(y0[7]) );
  AOI22X1 U885 ( .A0(N1634), .A1(n149), .B0(y0_tmp[7]), .B1(n88), .Y(n575) );
  INVX1 U886 ( .A(n572), .Y(y1[0]) );
  AOI22X1 U887 ( .A0(N1644), .A1(n148), .B0(y1_tmp[0]), .B1(n89), .Y(n572) );
  INVX1 U888 ( .A(n561), .Y(y1[4]) );
  AOI22X1 U889 ( .A0(N1648), .A1(n143), .B0(y1_tmp[4]), .B1(n90), .Y(n561) );
  INVX1 U890 ( .A(n559), .Y(y1[6]) );
  AOI22X1 U891 ( .A0(N1650), .A1(n142), .B0(y1_tmp[6]), .B1(n90), .Y(n559) );
  INVX1 U892 ( .A(n558), .Y(y1[7]) );
  AOI22X1 U893 ( .A0(N1651), .A1(n142), .B0(y1_tmp[7]), .B1(n90), .Y(n558) );
  INVX1 U894 ( .A(n555), .Y(y2[0]) );
  AOI22X1 U895 ( .A0(N1661), .A1(n139), .B0(y2_tmp[0]), .B1(n90), .Y(n555) );
  INVX1 U896 ( .A(n544), .Y(y2[4]) );
  AOI22X1 U897 ( .A0(N1665), .A1(n136), .B0(y2_tmp[4]), .B1(n91), .Y(n544) );
  INVX1 U898 ( .A(n542), .Y(y2[6]) );
  AOI22X1 U899 ( .A0(N1667), .A1(n135), .B0(y2_tmp[6]), .B1(n91), .Y(n542) );
  INVX1 U900 ( .A(n541), .Y(y2[7]) );
  AOI22X1 U901 ( .A0(N1668), .A1(n134), .B0(y2_tmp[7]), .B1(n91), .Y(n541) );
  INVX1 U902 ( .A(n538), .Y(y3[0]) );
  AOI22X1 U903 ( .A0(N1678), .A1(n133), .B0(y3_tmp[0]), .B1(n91), .Y(n538) );
  INVX1 U904 ( .A(n527), .Y(y3[4]) );
  AOI22X1 U905 ( .A0(N1682), .A1(n128), .B0(y3_tmp[4]), .B1(n87), .Y(n527) );
  INVX1 U906 ( .A(n525), .Y(y3[6]) );
  AOI22X1 U907 ( .A0(N1684), .A1(n180), .B0(y3_tmp[6]), .B1(n86), .Y(n525) );
  INVX1 U908 ( .A(n510), .Y(y4[4]) );
  INVX1 U909 ( .A(n509), .Y(y4[5]) );
  INVX1 U910 ( .A(n508), .Y(y4[6]) );
  INVX1 U911 ( .A(n507), .Y(y4[7]) );
  INVX1 U912 ( .A(n506), .Y(y4[8]) );
  INVX1 U913 ( .A(n505), .Y(y4[9]) );
  INVX1 U914 ( .A(n504), .Y(y5[0]) );
  INVX1 U915 ( .A(n496), .Y(y5[1]) );
  INVX1 U916 ( .A(n495), .Y(y5[2]) );
  INVX1 U917 ( .A(n494), .Y(y5[3]) );
  INVX1 U918 ( .A(n493), .Y(y5[4]) );
  INVX1 U919 ( .A(n492), .Y(y5[5]) );
  INVX1 U920 ( .A(n491), .Y(y5[6]) );
  INVX1 U921 ( .A(n490), .Y(y5[7]) );
  INVX1 U922 ( .A(n489), .Y(y5[8]) );
  INVX1 U923 ( .A(n488), .Y(y5[9]) );
  INVX1 U924 ( .A(n487), .Y(y6[0]) );
  INVX1 U925 ( .A(n479), .Y(y6[1]) );
  INVX1 U926 ( .A(n478), .Y(y6[2]) );
  INVX1 U927 ( .A(n477), .Y(y6[3]) );
  INVX1 U928 ( .A(n476), .Y(y6[4]) );
  INVX1 U929 ( .A(n475), .Y(y6[5]) );
  INVX1 U930 ( .A(n474), .Y(y6[6]) );
  INVX1 U931 ( .A(n473), .Y(y6[7]) );
  INVX1 U932 ( .A(n472), .Y(y6[8]) );
  INVX1 U933 ( .A(n471), .Y(y6[9]) );
  INVX1 U934 ( .A(n521), .Y(y4[0]) );
  INVX1 U935 ( .A(n513), .Y(y4[1]) );
  INVX1 U936 ( .A(n512), .Y(y4[2]) );
  INVX1 U937 ( .A(n511), .Y(y4[3]) );
  INVX1 U938 ( .A(n470), .Y(y7[0]) );
  INVX1 U939 ( .A(n462), .Y(y7[1]) );
  INVX1 U940 ( .A(n461), .Y(y7[2]) );
  INVX1 U941 ( .A(n460), .Y(y7[3]) );
  INVX1 U942 ( .A(n459), .Y(y7[4]) );
  INVX1 U943 ( .A(n458), .Y(y7[5]) );
  INVX1 U944 ( .A(n457), .Y(y7[6]) );
  INVX1 U945 ( .A(n456), .Y(y7[7]) );
  INVX1 U946 ( .A(n455), .Y(y7[8]) );
  INVX1 U947 ( .A(n453), .Y(y7[9]) );
  AOI22X1 U948 ( .A0(N1695), .A1(n126), .B0(y4_tmp[0]), .B1(n86), .Y(n521) );
  AOI22X1 U949 ( .A0(N1696), .A1(n122), .B0(y4_tmp[1]), .B1(n85), .Y(n513) );
  AOI22X1 U950 ( .A0(N1697), .A1(n122), .B0(y4_tmp[2]), .B1(n85), .Y(n512) );
  AOI22X1 U951 ( .A0(N1698), .A1(n121), .B0(y4_tmp[3]), .B1(n85), .Y(n511) );
  AOI22X1 U952 ( .A0(N1699), .A1(n121), .B0(y4_tmp[4]), .B1(n85), .Y(n510) );
  AOI22X1 U953 ( .A0(N1700), .A1(n120), .B0(y4_tmp[5]), .B1(n85), .Y(n509) );
  AOI22X1 U954 ( .A0(N1712), .A1(n118), .B0(y5_tmp[0]), .B1(n85), .Y(n504) );
  AOI22X1 U955 ( .A0(N1713), .A1(n114), .B0(y5_tmp[1]), .B1(n84), .Y(n496) );
  AOI22X1 U956 ( .A0(N1714), .A1(n113), .B0(y5_tmp[2]), .B1(n84), .Y(n495) );
  AOI22X1 U957 ( .A0(N1715), .A1(n113), .B0(y5_tmp[3]), .B1(n84), .Y(n494) );
  AOI22X1 U958 ( .A0(N1716), .A1(n112), .B0(y5_tmp[4]), .B1(n84), .Y(n493) );
  AOI22X1 U959 ( .A0(N1717), .A1(n112), .B0(y5_tmp[5]), .B1(n84), .Y(n492) );
  AOI22X1 U960 ( .A0(N1729), .A1(n109), .B0(y6_tmp[0]), .B1(n83), .Y(n487) );
  AOI22X1 U961 ( .A0(N1730), .A1(n105), .B0(y6_tmp[1]), .B1(n83), .Y(n479) );
  AOI22X1 U962 ( .A0(N1731), .A1(n105), .B0(y6_tmp[2]), .B1(n83), .Y(n478) );
  AOI22X1 U963 ( .A0(N1732), .A1(n104), .B0(y6_tmp[3]), .B1(n82), .Y(n477) );
  AOI22X1 U964 ( .A0(N1733), .A1(n104), .B0(y6_tmp[4]), .B1(n82), .Y(n476) );
  AOI22X1 U965 ( .A0(N1734), .A1(n103), .B0(y6_tmp[5]), .B1(n82), .Y(n475) );
  AOI22X1 U966 ( .A0(N1746), .A1(n101), .B0(y7_tmp[0]), .B1(n82), .Y(n470) );
  AOI22X1 U967 ( .A0(N1747), .A1(n97), .B0(y7_tmp[1]), .B1(n81), .Y(n462) );
  AOI22X1 U968 ( .A0(N1748), .A1(n96), .B0(y7_tmp[2]), .B1(n81), .Y(n461) );
  AOI22X1 U969 ( .A0(N1749), .A1(n96), .B0(y7_tmp[3]), .B1(n81), .Y(n460) );
  AOI22X1 U970 ( .A0(N1750), .A1(n95), .B0(y7_tmp[4]), .B1(n81), .Y(n459) );
  AOI22X1 U971 ( .A0(N1751), .A1(n95), .B0(y7_tmp[5]), .B1(n81), .Y(n458) );
  BUFX3 U972 ( .A(x5[13]), .Y(n66) );
  BUFX3 U973 ( .A(x5[14]), .Y(n67) );
  BUFX3 U974 ( .A(x6[13]), .Y(n53) );
  BUFX3 U975 ( .A(x6[14]), .Y(n54) );
  BUFX3 U976 ( .A(x4[13]), .Y(n79) );
  BUFX3 U977 ( .A(x4[14]), .Y(n80) );
  BUFX3 U978 ( .A(x7[13]), .Y(n40) );
  BUFX3 U979 ( .A(x7[14]), .Y(n41) );
  INVX1 U980 ( .A(x7_50[21]), .Y(n186) );
  INVX1 U981 ( .A(x5_50[21]), .Y(n254) );
  INVX1 U982 ( .A(x5_tmp[24]), .Y(n301) );
  INVX1 U983 ( .A(x4_tmp[24]), .Y(n375) );
  INVX1 U984 ( .A(x7_tmp[24]), .Y(n300) );
  INVX1 U985 ( .A(x6_tmp[24]), .Y(n326) );
  INVX1 U986 ( .A(x7_89[22]), .Y(n231) );
  INVX1 U987 ( .A(x5_89[22]), .Y(n208) );
  AOI22X1 U988 ( .A0(N1643), .A1(n153), .B0(y0_tmp[16]), .B1(n88), .Y(n582) );
  AOI22X1 U989 ( .A0(N1660), .A1(n126), .B0(y1_tmp[16]), .B1(n89), .Y(n565) );
  AOI22X1 U990 ( .A0(N1677), .A1(n138), .B0(y2_tmp[16]), .B1(n91), .Y(n548) );
  AOI22X1 U991 ( .A0(N1694), .A1(n119), .B0(y3_tmp[16]), .B1(n87), .Y(n531) );
  AOI22X1 U992 ( .A0(N1711), .A1(n123), .B0(y4_tmp[16]), .B1(n86), .Y(n514) );
  AOI22X1 U993 ( .A0(N1728), .A1(n114), .B0(y5_tmp[16]), .B1(n84), .Y(n497) );
  AOI22X1 U994 ( .A0(N1745), .A1(n106), .B0(y6_tmp[16]), .B1(n83), .Y(n480) );
  AOI22X1 U995 ( .A0(N1762), .A1(n97), .B0(y7_tmp[16]), .B1(n81), .Y(n463) );
  AND2X1 U1020 ( .A(add_184_carry_27_), .B(y4_tmp[25]), .Y(N1711) );
  XOR2X1 U1021 ( .A(y4_tmp[25]), .B(add_184_carry_27_), .Y(N1710) );
  AND2X1 U1022 ( .A(add_184_carry_26_), .B(y4_tmp[25]), .Y(add_184_carry_27_)
         );
  XOR2X1 U1023 ( .A(y4_tmp[25]), .B(add_184_carry_26_), .Y(N1709) );
  AND2X1 U1024 ( .A(add_184_carry_25_), .B(y4_tmp[25]), .Y(add_184_carry_26_)
         );
  XOR2X1 U1025 ( .A(y4_tmp[25]), .B(add_184_carry_25_), .Y(N1708) );
  AND2X1 U1026 ( .A(add_184_carry_24_), .B(y4_tmp[24]), .Y(add_184_carry_25_)
         );
  XOR2X1 U1027 ( .A(y4_tmp[24]), .B(add_184_carry_24_), .Y(N1707) );
  AND2X1 U1028 ( .A(add_184_carry_23_), .B(y4_tmp[23]), .Y(add_184_carry_24_)
         );
  XOR2X1 U1029 ( .A(y4_tmp[23]), .B(add_184_carry_23_), .Y(N1706) );
  AND2X1 U1030 ( .A(add_184_carry_22_), .B(y4_tmp[22]), .Y(add_184_carry_23_)
         );
  XOR2X1 U1031 ( .A(y4_tmp[22]), .B(add_184_carry_22_), .Y(N1705) );
  AND2X1 U1032 ( .A(add_184_carry_21_), .B(y4_tmp[21]), .Y(add_184_carry_22_)
         );
  XOR2X1 U1033 ( .A(y4_tmp[21]), .B(add_184_carry_21_), .Y(N1704) );
  AND2X1 U1034 ( .A(add_184_carry_20_), .B(y4_tmp[20]), .Y(add_184_carry_21_)
         );
  XOR2X1 U1035 ( .A(y4_tmp[20]), .B(add_184_carry_20_), .Y(N1703) );
  AND2X1 U1036 ( .A(add_184_carry_19_), .B(y4_tmp[19]), .Y(add_184_carry_20_)
         );
  XOR2X1 U1037 ( .A(y4_tmp[19]), .B(add_184_carry_19_), .Y(N1702) );
  AND2X1 U1038 ( .A(add_184_carry_18_), .B(y4_tmp[18]), .Y(add_184_carry_19_)
         );
  XOR2X1 U1039 ( .A(y4_tmp[18]), .B(add_184_carry_18_), .Y(N1701) );
  AND2X1 U1040 ( .A(add_184_carry_17_), .B(y4_tmp[17]), .Y(add_184_carry_18_)
         );
  XOR2X1 U1041 ( .A(y4_tmp[17]), .B(add_184_carry_17_), .Y(N1700) );
  AND2X1 U1042 ( .A(add_184_carry_16_), .B(y4_tmp[16]), .Y(add_184_carry_17_)
         );
  XOR2X1 U1043 ( .A(y4_tmp[16]), .B(add_184_carry_16_), .Y(N1699) );
  AND2X1 U1044 ( .A(add_184_carry_15_), .B(y4_tmp[15]), .Y(add_184_carry_16_)
         );
  XOR2X1 U1045 ( .A(y4_tmp[15]), .B(add_184_carry_15_), .Y(N1698) );
  AND2X1 U1046 ( .A(add_184_carry_14_), .B(y4_tmp[14]), .Y(add_184_carry_15_)
         );
  XOR2X1 U1047 ( .A(y4_tmp[14]), .B(add_184_carry_14_), .Y(N1697) );
  AND2X1 U1048 ( .A(add_184_carry_13_), .B(y4_tmp[13]), .Y(add_184_carry_14_)
         );
  XOR2X1 U1049 ( .A(y4_tmp[13]), .B(add_184_carry_13_), .Y(N1696) );
  AND2X1 U1050 ( .A(y4_tmp[11]), .B(y4_tmp[12]), .Y(add_184_carry_13_) );
  XOR2X1 U1051 ( .A(y4_tmp[12]), .B(y4_tmp[11]), .Y(N1695) );
  AND2X1 U1052 ( .A(add_185_carry_27_), .B(y5_tmp[25]), .Y(N1728) );
  XOR2X1 U1053 ( .A(y5_tmp[25]), .B(add_185_carry_27_), .Y(N1727) );
  AND2X1 U1054 ( .A(add_185_carry_26_), .B(y5_tmp[25]), .Y(add_185_carry_27_)
         );
  XOR2X1 U1055 ( .A(y5_tmp[25]), .B(add_185_carry_26_), .Y(N1726) );
  AND2X1 U1056 ( .A(add_185_carry_25_), .B(y5_tmp[25]), .Y(add_185_carry_26_)
         );
  XOR2X1 U1057 ( .A(y5_tmp[25]), .B(add_185_carry_25_), .Y(N1725) );
  AND2X1 U1058 ( .A(add_185_carry_24_), .B(y5_tmp[24]), .Y(add_185_carry_25_)
         );
  XOR2X1 U1059 ( .A(y5_tmp[24]), .B(add_185_carry_24_), .Y(N1724) );
  AND2X1 U1060 ( .A(add_185_carry_23_), .B(y5_tmp[23]), .Y(add_185_carry_24_)
         );
  XOR2X1 U1061 ( .A(y5_tmp[23]), .B(add_185_carry_23_), .Y(N1723) );
  AND2X1 U1062 ( .A(add_185_carry_22_), .B(y5_tmp[22]), .Y(add_185_carry_23_)
         );
  XOR2X1 U1063 ( .A(y5_tmp[22]), .B(add_185_carry_22_), .Y(N1722) );
  AND2X1 U1064 ( .A(add_185_carry_21_), .B(y5_tmp[21]), .Y(add_185_carry_22_)
         );
  XOR2X1 U1065 ( .A(y5_tmp[21]), .B(add_185_carry_21_), .Y(N1721) );
  AND2X1 U1066 ( .A(add_185_carry_20_), .B(y5_tmp[20]), .Y(add_185_carry_21_)
         );
  XOR2X1 U1067 ( .A(y5_tmp[20]), .B(add_185_carry_20_), .Y(N1720) );
  AND2X1 U1068 ( .A(add_185_carry_19_), .B(y5_tmp[19]), .Y(add_185_carry_20_)
         );
  XOR2X1 U1069 ( .A(y5_tmp[19]), .B(add_185_carry_19_), .Y(N1719) );
  AND2X1 U1070 ( .A(add_185_carry_18_), .B(y5_tmp[18]), .Y(add_185_carry_19_)
         );
  XOR2X1 U1071 ( .A(y5_tmp[18]), .B(add_185_carry_18_), .Y(N1718) );
  AND2X1 U1072 ( .A(add_185_carry_17_), .B(y5_tmp[17]), .Y(add_185_carry_18_)
         );
  XOR2X1 U1073 ( .A(y5_tmp[17]), .B(add_185_carry_17_), .Y(N1717) );
  AND2X1 U1074 ( .A(add_185_carry_16_), .B(y5_tmp[16]), .Y(add_185_carry_17_)
         );
  XOR2X1 U1075 ( .A(y5_tmp[16]), .B(add_185_carry_16_), .Y(N1716) );
  AND2X1 U1076 ( .A(add_185_carry_15_), .B(y5_tmp[15]), .Y(add_185_carry_16_)
         );
  XOR2X1 U1077 ( .A(y5_tmp[15]), .B(add_185_carry_15_), .Y(N1715) );
  AND2X1 U1078 ( .A(add_185_carry_14_), .B(y5_tmp[14]), .Y(add_185_carry_15_)
         );
  XOR2X1 U1079 ( .A(y5_tmp[14]), .B(add_185_carry_14_), .Y(N1714) );
  AND2X1 U1080 ( .A(add_185_carry_13_), .B(y5_tmp[13]), .Y(add_185_carry_14_)
         );
  XOR2X1 U1081 ( .A(y5_tmp[13]), .B(add_185_carry_13_), .Y(N1713) );
  AND2X1 U1082 ( .A(y5_tmp[11]), .B(y5_tmp[12]), .Y(add_185_carry_13_) );
  XOR2X1 U1083 ( .A(y5_tmp[12]), .B(y5_tmp[11]), .Y(N1712) );
  AND2X1 U1084 ( .A(add_186_carry_27_), .B(y6_tmp[25]), .Y(N1745) );
  XOR2X1 U1085 ( .A(y6_tmp[25]), .B(add_186_carry_27_), .Y(N1744) );
  AND2X1 U1086 ( .A(add_186_carry_26_), .B(y6_tmp[25]), .Y(add_186_carry_27_)
         );
  XOR2X1 U1087 ( .A(y6_tmp[25]), .B(add_186_carry_26_), .Y(N1743) );
  AND2X1 U1088 ( .A(add_186_carry_25_), .B(y6_tmp[25]), .Y(add_186_carry_26_)
         );
  XOR2X1 U1089 ( .A(y6_tmp[25]), .B(add_186_carry_25_), .Y(N1742) );
  AND2X1 U1090 ( .A(add_186_carry_24_), .B(y6_tmp[24]), .Y(add_186_carry_25_)
         );
  XOR2X1 U1091 ( .A(y6_tmp[24]), .B(add_186_carry_24_), .Y(N1741) );
  AND2X1 U1092 ( .A(add_186_carry_23_), .B(y6_tmp[23]), .Y(add_186_carry_24_)
         );
  XOR2X1 U1093 ( .A(y6_tmp[23]), .B(add_186_carry_23_), .Y(N1740) );
  AND2X1 U1094 ( .A(add_186_carry_22_), .B(y6_tmp[22]), .Y(add_186_carry_23_)
         );
  XOR2X1 U1095 ( .A(y6_tmp[22]), .B(add_186_carry_22_), .Y(N1739) );
  AND2X1 U1096 ( .A(add_186_carry_21_), .B(y6_tmp[21]), .Y(add_186_carry_22_)
         );
  XOR2X1 U1097 ( .A(y6_tmp[21]), .B(add_186_carry_21_), .Y(N1738) );
  AND2X1 U1098 ( .A(add_186_carry_20_), .B(y6_tmp[20]), .Y(add_186_carry_21_)
         );
  XOR2X1 U1099 ( .A(y6_tmp[20]), .B(add_186_carry_20_), .Y(N1737) );
  AND2X1 U1100 ( .A(add_186_carry_19_), .B(y6_tmp[19]), .Y(add_186_carry_20_)
         );
  XOR2X1 U1101 ( .A(y6_tmp[19]), .B(add_186_carry_19_), .Y(N1736) );
  AND2X1 U1102 ( .A(add_186_carry_18_), .B(y6_tmp[18]), .Y(add_186_carry_19_)
         );
  XOR2X1 U1103 ( .A(y6_tmp[18]), .B(add_186_carry_18_), .Y(N1735) );
  AND2X1 U1104 ( .A(add_186_carry_17_), .B(y6_tmp[17]), .Y(add_186_carry_18_)
         );
  XOR2X1 U1105 ( .A(y6_tmp[17]), .B(add_186_carry_17_), .Y(N1734) );
  AND2X1 U1106 ( .A(add_186_carry_16_), .B(y6_tmp[16]), .Y(add_186_carry_17_)
         );
  XOR2X1 U1107 ( .A(y6_tmp[16]), .B(add_186_carry_16_), .Y(N1733) );
  AND2X1 U1108 ( .A(add_186_carry_15_), .B(y6_tmp[15]), .Y(add_186_carry_16_)
         );
  XOR2X1 U1109 ( .A(y6_tmp[15]), .B(add_186_carry_15_), .Y(N1732) );
  AND2X1 U1110 ( .A(add_186_carry_14_), .B(y6_tmp[14]), .Y(add_186_carry_15_)
         );
  XOR2X1 U1111 ( .A(y6_tmp[14]), .B(add_186_carry_14_), .Y(N1731) );
  AND2X1 U1112 ( .A(add_186_carry_13_), .B(y6_tmp[13]), .Y(add_186_carry_14_)
         );
  XOR2X1 U1113 ( .A(y6_tmp[13]), .B(add_186_carry_13_), .Y(N1730) );
  AND2X1 U1114 ( .A(y6_tmp[11]), .B(y6_tmp[12]), .Y(add_186_carry_13_) );
  XOR2X1 U1115 ( .A(y6_tmp[12]), .B(y6_tmp[11]), .Y(N1729) );
  AND2X1 U1116 ( .A(add_187_carry_27_), .B(y7_tmp[25]), .Y(N1762) );
  XOR2X1 U1117 ( .A(y7_tmp[25]), .B(add_187_carry_27_), .Y(N1761) );
  AND2X1 U1118 ( .A(add_187_carry_26_), .B(y7_tmp[25]), .Y(add_187_carry_27_)
         );
  XOR2X1 U1119 ( .A(y7_tmp[25]), .B(add_187_carry_26_), .Y(N1760) );
  AND2X1 U1120 ( .A(add_187_carry_25_), .B(y7_tmp[25]), .Y(add_187_carry_26_)
         );
  XOR2X1 U1121 ( .A(y7_tmp[25]), .B(add_187_carry_25_), .Y(N1759) );
  AND2X1 U1122 ( .A(add_187_carry_24_), .B(y7_tmp[24]), .Y(add_187_carry_25_)
         );
  XOR2X1 U1123 ( .A(y7_tmp[24]), .B(add_187_carry_24_), .Y(N1758) );
  AND2X1 U1124 ( .A(add_187_carry_23_), .B(y7_tmp[23]), .Y(add_187_carry_24_)
         );
  XOR2X1 U1125 ( .A(y7_tmp[23]), .B(add_187_carry_23_), .Y(N1757) );
  AND2X1 U1126 ( .A(add_187_carry_22_), .B(y7_tmp[22]), .Y(add_187_carry_23_)
         );
  XOR2X1 U1127 ( .A(y7_tmp[22]), .B(add_187_carry_22_), .Y(N1756) );
  AND2X1 U1128 ( .A(add_187_carry_21_), .B(y7_tmp[21]), .Y(add_187_carry_22_)
         );
  XOR2X1 U1129 ( .A(y7_tmp[21]), .B(add_187_carry_21_), .Y(N1755) );
  AND2X1 U1130 ( .A(add_187_carry_20_), .B(y7_tmp[20]), .Y(add_187_carry_21_)
         );
  XOR2X1 U1131 ( .A(y7_tmp[20]), .B(add_187_carry_20_), .Y(N1754) );
  AND2X1 U1132 ( .A(add_187_carry_19_), .B(y7_tmp[19]), .Y(add_187_carry_20_)
         );
  XOR2X1 U1133 ( .A(y7_tmp[19]), .B(add_187_carry_19_), .Y(N1753) );
  AND2X1 U1134 ( .A(add_187_carry_18_), .B(y7_tmp[18]), .Y(add_187_carry_19_)
         );
  XOR2X1 U1135 ( .A(y7_tmp[18]), .B(add_187_carry_18_), .Y(N1752) );
  AND2X1 U1136 ( .A(add_187_carry_17_), .B(y7_tmp[17]), .Y(add_187_carry_18_)
         );
  XOR2X1 U1137 ( .A(y7_tmp[17]), .B(add_187_carry_17_), .Y(N1751) );
  AND2X1 U1138 ( .A(add_187_carry_16_), .B(y7_tmp[16]), .Y(add_187_carry_17_)
         );
  XOR2X1 U1139 ( .A(y7_tmp[16]), .B(add_187_carry_16_), .Y(N1750) );
  AND2X1 U1140 ( .A(add_187_carry_15_), .B(y7_tmp[15]), .Y(add_187_carry_16_)
         );
  XOR2X1 U1141 ( .A(y7_tmp[15]), .B(add_187_carry_15_), .Y(N1749) );
  AND2X1 U1142 ( .A(add_187_carry_14_), .B(y7_tmp[14]), .Y(add_187_carry_15_)
         );
  XOR2X1 U1143 ( .A(y7_tmp[14]), .B(add_187_carry_14_), .Y(N1748) );
  AND2X1 U1144 ( .A(add_187_carry_13_), .B(y7_tmp[13]), .Y(add_187_carry_14_)
         );
  XOR2X1 U1145 ( .A(y7_tmp[13]), .B(add_187_carry_13_), .Y(N1747) );
  AND2X1 U1146 ( .A(y7_tmp[11]), .B(y7_tmp[12]), .Y(add_187_carry_13_) );
  XOR2X1 U1147 ( .A(y7_tmp[12]), .B(y7_tmp[11]), .Y(N1746) );
  AND2X1 U1148 ( .A(add_180_carry_27_), .B(y0_tmp[25]), .Y(N1643) );
  XOR2X1 U1149 ( .A(y0_tmp[25]), .B(add_180_carry_27_), .Y(N1642) );
  AND2X1 U1150 ( .A(add_180_carry_26_), .B(y0_tmp[25]), .Y(add_180_carry_27_)
         );
  XOR2X1 U1151 ( .A(y0_tmp[25]), .B(add_180_carry_26_), .Y(N1641) );
  AND2X1 U1152 ( .A(add_180_carry_25_), .B(y0_tmp[25]), .Y(add_180_carry_26_)
         );
  XOR2X1 U1153 ( .A(y0_tmp[25]), .B(add_180_carry_25_), .Y(N1640) );
  AND2X1 U1154 ( .A(add_180_carry_24_), .B(y0_tmp[24]), .Y(add_180_carry_25_)
         );
  XOR2X1 U1155 ( .A(y0_tmp[24]), .B(add_180_carry_24_), .Y(N1639) );
  AND2X1 U1156 ( .A(add_180_carry_23_), .B(y0_tmp[23]), .Y(add_180_carry_24_)
         );
  XOR2X1 U1157 ( .A(y0_tmp[23]), .B(add_180_carry_23_), .Y(N1638) );
  AND2X1 U1158 ( .A(add_180_carry_22_), .B(y0_tmp[22]), .Y(add_180_carry_23_)
         );
  XOR2X1 U1159 ( .A(y0_tmp[22]), .B(add_180_carry_22_), .Y(N1637) );
  AND2X1 U1160 ( .A(add_180_carry_21_), .B(y0_tmp[21]), .Y(add_180_carry_22_)
         );
  XOR2X1 U1161 ( .A(y0_tmp[21]), .B(add_180_carry_21_), .Y(N1636) );
  AND2X1 U1162 ( .A(add_180_carry_20_), .B(y0_tmp[20]), .Y(add_180_carry_21_)
         );
  XOR2X1 U1163 ( .A(y0_tmp[20]), .B(add_180_carry_20_), .Y(N1635) );
  AND2X1 U1164 ( .A(add_180_carry_19_), .B(y0_tmp[19]), .Y(add_180_carry_20_)
         );
  XOR2X1 U1165 ( .A(y0_tmp[19]), .B(add_180_carry_19_), .Y(N1634) );
  AND2X1 U1166 ( .A(add_180_carry_18_), .B(y0_tmp[18]), .Y(add_180_carry_19_)
         );
  XOR2X1 U1167 ( .A(y0_tmp[18]), .B(add_180_carry_18_), .Y(N1633) );
  AND2X1 U1168 ( .A(add_180_carry_17_), .B(y0_tmp[17]), .Y(add_180_carry_18_)
         );
  XOR2X1 U1169 ( .A(y0_tmp[17]), .B(add_180_carry_17_), .Y(N1632) );
  AND2X1 U1170 ( .A(add_180_carry_16_), .B(y0_tmp[16]), .Y(add_180_carry_17_)
         );
  XOR2X1 U1171 ( .A(y0_tmp[16]), .B(add_180_carry_16_), .Y(N1631) );
  AND2X1 U1172 ( .A(add_180_carry_15_), .B(y0_tmp[15]), .Y(add_180_carry_16_)
         );
  XOR2X1 U1173 ( .A(y0_tmp[15]), .B(add_180_carry_15_), .Y(N1630) );
  AND2X1 U1174 ( .A(add_180_carry_14_), .B(y0_tmp[14]), .Y(add_180_carry_15_)
         );
  XOR2X1 U1175 ( .A(y0_tmp[14]), .B(add_180_carry_14_), .Y(N1629) );
  AND2X1 U1176 ( .A(add_180_carry_13_), .B(y0_tmp[13]), .Y(add_180_carry_14_)
         );
  XOR2X1 U1177 ( .A(y0_tmp[13]), .B(add_180_carry_13_), .Y(N1628) );
  AND2X1 U1178 ( .A(y0_tmp[11]), .B(y0_tmp[12]), .Y(add_180_carry_13_) );
  XOR2X1 U1179 ( .A(y0_tmp[12]), .B(y0_tmp[11]), .Y(N1627) );
  AND2X1 U1180 ( .A(add_181_carry_27_), .B(y1_tmp[25]), .Y(N1660) );
  XOR2X1 U1181 ( .A(y1_tmp[25]), .B(add_181_carry_27_), .Y(N1659) );
  AND2X1 U1182 ( .A(add_181_carry_26_), .B(y1_tmp[25]), .Y(add_181_carry_27_)
         );
  XOR2X1 U1183 ( .A(y1_tmp[25]), .B(add_181_carry_26_), .Y(N1658) );
  AND2X1 U1184 ( .A(add_181_carry_25_), .B(y1_tmp[25]), .Y(add_181_carry_26_)
         );
  XOR2X1 U1185 ( .A(y1_tmp[25]), .B(add_181_carry_25_), .Y(N1657) );
  AND2X1 U1186 ( .A(add_181_carry_24_), .B(y1_tmp[24]), .Y(add_181_carry_25_)
         );
  XOR2X1 U1187 ( .A(y1_tmp[24]), .B(add_181_carry_24_), .Y(N1656) );
  AND2X1 U1188 ( .A(add_181_carry_23_), .B(y1_tmp[23]), .Y(add_181_carry_24_)
         );
  XOR2X1 U1189 ( .A(y1_tmp[23]), .B(add_181_carry_23_), .Y(N1655) );
  AND2X1 U1190 ( .A(add_181_carry_22_), .B(y1_tmp[22]), .Y(add_181_carry_23_)
         );
  XOR2X1 U1191 ( .A(y1_tmp[22]), .B(add_181_carry_22_), .Y(N1654) );
  AND2X1 U1192 ( .A(add_181_carry_21_), .B(y1_tmp[21]), .Y(add_181_carry_22_)
         );
  XOR2X1 U1193 ( .A(y1_tmp[21]), .B(add_181_carry_21_), .Y(N1653) );
  AND2X1 U1194 ( .A(add_181_carry_20_), .B(y1_tmp[20]), .Y(add_181_carry_21_)
         );
  XOR2X1 U1195 ( .A(y1_tmp[20]), .B(add_181_carry_20_), .Y(N1652) );
  AND2X1 U1196 ( .A(add_181_carry_19_), .B(y1_tmp[19]), .Y(add_181_carry_20_)
         );
  XOR2X1 U1197 ( .A(y1_tmp[19]), .B(add_181_carry_19_), .Y(N1651) );
  AND2X1 U1198 ( .A(add_181_carry_18_), .B(y1_tmp[18]), .Y(add_181_carry_19_)
         );
  XOR2X1 U1199 ( .A(y1_tmp[18]), .B(add_181_carry_18_), .Y(N1650) );
  AND2X1 U1200 ( .A(add_181_carry_17_), .B(y1_tmp[17]), .Y(add_181_carry_18_)
         );
  XOR2X1 U1201 ( .A(y1_tmp[17]), .B(add_181_carry_17_), .Y(N1649) );
  AND2X1 U1202 ( .A(add_181_carry_16_), .B(y1_tmp[16]), .Y(add_181_carry_17_)
         );
  XOR2X1 U1203 ( .A(y1_tmp[16]), .B(add_181_carry_16_), .Y(N1648) );
  AND2X1 U1204 ( .A(add_181_carry_15_), .B(y1_tmp[15]), .Y(add_181_carry_16_)
         );
  XOR2X1 U1205 ( .A(y1_tmp[15]), .B(add_181_carry_15_), .Y(N1647) );
  AND2X1 U1206 ( .A(add_181_carry_14_), .B(y1_tmp[14]), .Y(add_181_carry_15_)
         );
  XOR2X1 U1207 ( .A(y1_tmp[14]), .B(add_181_carry_14_), .Y(N1646) );
  AND2X1 U1208 ( .A(add_181_carry_13_), .B(y1_tmp[13]), .Y(add_181_carry_14_)
         );
  XOR2X1 U1209 ( .A(y1_tmp[13]), .B(add_181_carry_13_), .Y(N1645) );
  AND2X1 U1210 ( .A(y1_tmp[11]), .B(y1_tmp[12]), .Y(add_181_carry_13_) );
  XOR2X1 U1211 ( .A(y1_tmp[12]), .B(y1_tmp[11]), .Y(N1644) );
  AND2X1 U1212 ( .A(add_182_carry_27_), .B(y2_tmp[25]), .Y(N1677) );
  XOR2X1 U1213 ( .A(y2_tmp[25]), .B(add_182_carry_27_), .Y(N1676) );
  AND2X1 U1214 ( .A(add_182_carry_26_), .B(y2_tmp[25]), .Y(add_182_carry_27_)
         );
  XOR2X1 U1215 ( .A(y2_tmp[25]), .B(add_182_carry_26_), .Y(N1675) );
  AND2X1 U1216 ( .A(add_182_carry_25_), .B(y2_tmp[25]), .Y(add_182_carry_26_)
         );
  XOR2X1 U1217 ( .A(y2_tmp[25]), .B(add_182_carry_25_), .Y(N1674) );
  AND2X1 U1218 ( .A(add_182_carry_24_), .B(y2_tmp[24]), .Y(add_182_carry_25_)
         );
  XOR2X1 U1219 ( .A(y2_tmp[24]), .B(add_182_carry_24_), .Y(N1673) );
  AND2X1 U1220 ( .A(add_182_carry_23_), .B(y2_tmp[23]), .Y(add_182_carry_24_)
         );
  XOR2X1 U1221 ( .A(y2_tmp[23]), .B(add_182_carry_23_), .Y(N1672) );
  AND2X1 U1222 ( .A(add_182_carry_22_), .B(y2_tmp[22]), .Y(add_182_carry_23_)
         );
  XOR2X1 U1223 ( .A(y2_tmp[22]), .B(add_182_carry_22_), .Y(N1671) );
  AND2X1 U1224 ( .A(add_182_carry_21_), .B(y2_tmp[21]), .Y(add_182_carry_22_)
         );
  XOR2X1 U1225 ( .A(y2_tmp[21]), .B(add_182_carry_21_), .Y(N1670) );
  AND2X1 U1226 ( .A(add_182_carry_20_), .B(y2_tmp[20]), .Y(add_182_carry_21_)
         );
  XOR2X1 U1227 ( .A(y2_tmp[20]), .B(add_182_carry_20_), .Y(N1669) );
  AND2X1 U1228 ( .A(add_182_carry_19_), .B(y2_tmp[19]), .Y(add_182_carry_20_)
         );
  XOR2X1 U1229 ( .A(y2_tmp[19]), .B(add_182_carry_19_), .Y(N1668) );
  AND2X1 U1230 ( .A(add_182_carry_18_), .B(y2_tmp[18]), .Y(add_182_carry_19_)
         );
  XOR2X1 U1231 ( .A(y2_tmp[18]), .B(add_182_carry_18_), .Y(N1667) );
  AND2X1 U1232 ( .A(add_182_carry_17_), .B(y2_tmp[17]), .Y(add_182_carry_18_)
         );
  XOR2X1 U1233 ( .A(y2_tmp[17]), .B(add_182_carry_17_), .Y(N1666) );
  AND2X1 U1234 ( .A(add_182_carry_16_), .B(y2_tmp[16]), .Y(add_182_carry_17_)
         );
  XOR2X1 U1235 ( .A(y2_tmp[16]), .B(add_182_carry_16_), .Y(N1665) );
  AND2X1 U1236 ( .A(add_182_carry_15_), .B(y2_tmp[15]), .Y(add_182_carry_16_)
         );
  XOR2X1 U1237 ( .A(y2_tmp[15]), .B(add_182_carry_15_), .Y(N1664) );
  AND2X1 U1238 ( .A(add_182_carry_14_), .B(y2_tmp[14]), .Y(add_182_carry_15_)
         );
  XOR2X1 U1239 ( .A(y2_tmp[14]), .B(add_182_carry_14_), .Y(N1663) );
  AND2X1 U1240 ( .A(add_182_carry_13_), .B(y2_tmp[13]), .Y(add_182_carry_14_)
         );
  XOR2X1 U1241 ( .A(y2_tmp[13]), .B(add_182_carry_13_), .Y(N1662) );
  AND2X1 U1242 ( .A(y2_tmp[11]), .B(y2_tmp[12]), .Y(add_182_carry_13_) );
  XOR2X1 U1243 ( .A(y2_tmp[12]), .B(y2_tmp[11]), .Y(N1661) );
  AND2X1 U1244 ( .A(add_183_carry_27_), .B(y3_tmp[25]), .Y(N1694) );
  XOR2X1 U1245 ( .A(y3_tmp[25]), .B(add_183_carry_27_), .Y(N1693) );
  AND2X1 U1246 ( .A(add_183_carry_26_), .B(y3_tmp[25]), .Y(add_183_carry_27_)
         );
  XOR2X1 U1247 ( .A(y3_tmp[25]), .B(add_183_carry_26_), .Y(N1692) );
  AND2X1 U1248 ( .A(add_183_carry_25_), .B(y3_tmp[25]), .Y(add_183_carry_26_)
         );
  XOR2X1 U1249 ( .A(y3_tmp[25]), .B(add_183_carry_25_), .Y(N1691) );
  AND2X1 U1250 ( .A(add_183_carry_24_), .B(y3_tmp[24]), .Y(add_183_carry_25_)
         );
  XOR2X1 U1251 ( .A(y3_tmp[24]), .B(add_183_carry_24_), .Y(N1690) );
  AND2X1 U1252 ( .A(add_183_carry_23_), .B(y3_tmp[23]), .Y(add_183_carry_24_)
         );
  XOR2X1 U1253 ( .A(y3_tmp[23]), .B(add_183_carry_23_), .Y(N1689) );
  AND2X1 U1254 ( .A(add_183_carry_22_), .B(y3_tmp[22]), .Y(add_183_carry_23_)
         );
  XOR2X1 U1255 ( .A(y3_tmp[22]), .B(add_183_carry_22_), .Y(N1688) );
  AND2X1 U1256 ( .A(add_183_carry_21_), .B(y3_tmp[21]), .Y(add_183_carry_22_)
         );
  XOR2X1 U1257 ( .A(y3_tmp[21]), .B(add_183_carry_21_), .Y(N1687) );
  AND2X1 U1258 ( .A(add_183_carry_20_), .B(y3_tmp[20]), .Y(add_183_carry_21_)
         );
  XOR2X1 U1259 ( .A(y3_tmp[20]), .B(add_183_carry_20_), .Y(N1686) );
  AND2X1 U1260 ( .A(add_183_carry_19_), .B(y3_tmp[19]), .Y(add_183_carry_20_)
         );
  XOR2X1 U1261 ( .A(y3_tmp[19]), .B(add_183_carry_19_), .Y(N1685) );
  AND2X1 U1262 ( .A(add_183_carry_18_), .B(y3_tmp[18]), .Y(add_183_carry_19_)
         );
  XOR2X1 U1263 ( .A(y3_tmp[18]), .B(add_183_carry_18_), .Y(N1684) );
  AND2X1 U1264 ( .A(add_183_carry_17_), .B(y3_tmp[17]), .Y(add_183_carry_18_)
         );
  XOR2X1 U1265 ( .A(y3_tmp[17]), .B(add_183_carry_17_), .Y(N1683) );
  AND2X1 U1266 ( .A(add_183_carry_16_), .B(y3_tmp[16]), .Y(add_183_carry_17_)
         );
  XOR2X1 U1267 ( .A(y3_tmp[16]), .B(add_183_carry_16_), .Y(N1682) );
  AND2X1 U1268 ( .A(add_183_carry_15_), .B(y3_tmp[15]), .Y(add_183_carry_16_)
         );
  XOR2X1 U1269 ( .A(y3_tmp[15]), .B(add_183_carry_15_), .Y(N1681) );
  AND2X1 U1270 ( .A(add_183_carry_14_), .B(y3_tmp[14]), .Y(add_183_carry_15_)
         );
  XOR2X1 U1271 ( .A(y3_tmp[14]), .B(add_183_carry_14_), .Y(N1680) );
  AND2X1 U1272 ( .A(add_183_carry_13_), .B(y3_tmp[13]), .Y(add_183_carry_14_)
         );
  XOR2X1 U1273 ( .A(y3_tmp[13]), .B(add_183_carry_13_), .Y(N1679) );
  AND2X1 U1274 ( .A(y3_tmp[11]), .B(y3_tmp[12]), .Y(add_183_carry_13_) );
  XOR2X1 U1275 ( .A(y3_tmp[12]), .B(y3_tmp[11]), .Y(N1678) );
  AND2X1 U1276 ( .A(x7[0]), .B(n3), .Y(add_104_carry_5_) );
  XOR2X1 U1277 ( .A(n3), .B(x7[0]), .Y(N340) );
  AND2X1 U1278 ( .A(x5[0]), .B(n56), .Y(add_86_carry_5_) );
  XOR2X1 U1279 ( .A(n56), .B(x5[0]), .Y(N170) );
  AND2X1 U1280 ( .A(x6[0]), .B(n43), .Y(add_95_carry_5_) );
  XOR2X1 U1281 ( .A(n43), .B(x6[0]), .Y(N255) );
  AND2X1 U1282 ( .A(x4[0]), .B(n69), .Y(add_77_carry_5_) );
  XOR2X1 U1283 ( .A(n69), .B(x4[0]), .Y(N85) );
  AND2X1 U1284 ( .A(x7[0]), .B(n2), .Y(add_102_carry_4_) );
  XOR2X1 U1285 ( .A(n2), .B(x7[0]), .Y(N319) );
  AND2X1 U1286 ( .A(x6[0]), .B(n42), .Y(add_93_carry_4_) );
  XOR2X1 U1287 ( .A(n42), .B(x6[0]), .Y(N234) );
  AND2X1 U1288 ( .A(x5[0]), .B(n55), .Y(add_84_carry_4_) );
  XOR2X1 U1289 ( .A(n55), .B(x5[0]), .Y(N149) );
  AND2X1 U1290 ( .A(x4[0]), .B(n68), .Y(add_75_carry_4_) );
  XOR2X1 U1291 ( .A(n68), .B(x4[0]), .Y(N64) );
  AND2X1 U1292 ( .A(x7[0]), .B(x7[1]), .Y(add_100_carry_5_) );
  XOR2X1 U1293 ( .A(x7[1]), .B(x7[0]), .Y(N299) );
  AND2X1 U1294 ( .A(x4[0]), .B(n72), .Y(add_72_carry_7_) );
  XOR2X1 U1295 ( .A(n72), .B(x4[0]), .Y(N23) );
  AND2X1 U1296 ( .A(x4[0]), .B(x4[1]), .Y(add_73_carry_5_) );
  XOR2X1 U1297 ( .A(x4[1]), .B(x4[0]), .Y(N44) );
  AND2X1 U1298 ( .A(x5[0]), .B(x5[1]), .Y(add_82_carry_5_) );
  XOR2X1 U1299 ( .A(x5[1]), .B(x5[0]), .Y(N129) );
  AND2X1 U1300 ( .A(x6[0]), .B(x6[1]), .Y(add_91_carry_5_) );
  XOR2X1 U1301 ( .A(x6[1]), .B(x6[0]), .Y(N214) );
  AND2X1 U1302 ( .A(x5[0]), .B(n59), .Y(add_81_carry_7_) );
  XOR2X1 U1303 ( .A(n59), .B(x5[0]), .Y(N108) );
  AND2X1 U1304 ( .A(x6[0]), .B(n46), .Y(add_90_carry_7_) );
  XOR2X1 U1305 ( .A(n46), .B(x6[0]), .Y(N193) );
  AND2X1 U1306 ( .A(x7[0]), .B(n6), .Y(add_99_carry_7_) );
  XOR2X1 U1307 ( .A(n6), .B(x7[0]), .Y(N278) );
endmodule


module idct_cal_shift12_add2048 ( clk, rstn, mode, start, x0, x1, x2, x3, x4, 
        x5, x6, x7, y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, 
        y14, y15, idct_ready, mode_out );
  input [1:0] mode;
  input [15:0] x0;
  input [15:0] x1;
  input [15:0] x2;
  input [15:0] x3;
  input [15:0] x4;
  input [15:0] x5;
  input [15:0] x6;
  input [15:0] x7;
  output [15:0] y0;
  output [15:0] y1;
  output [15:0] y2;
  output [15:0] y3;
  output [15:0] y4;
  output [15:0] y5;
  output [15:0] y6;
  output [15:0] y7;
  output [15:0] y8;
  output [15:0] y9;
  output [15:0] y10;
  output [15:0] y11;
  output [15:0] y12;
  output [15:0] y13;
  output [15:0] y14;
  output [15:0] y15;
  output [1:0] mode_out;
  input clk, rstn, start;
  output idct_ready;
  wire   idct4_ready, idct8_ready, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n325, n326, n327, n328, n329, n330, n331, n332;
  wire   [1:0] mode_delay2;
  wire   [1:0] mode_delay1;
  wire   [24:0] y0_idct4;
  wire   [24:0] y1_idct4;
  wire   [24:0] y2_idct4;
  wire   [24:0] y3_idct4;
  wire   [15:0] y0_idct8;
  wire   [15:0] y1_idct8;
  wire   [15:0] y2_idct8;
  wire   [15:0] y3_idct8;
  wire   [15:0] y4_idct8;
  wire   [15:0] y5_idct8;
  wire   [15:0] y6_idct8;
  wire   [15:0] y7_idct8;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75, 
        SYNOPSYS_UNCONNECTED__76, SYNOPSYS_UNCONNECTED__77, 
        SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79;

  CLKINVX8 U3 ( .A(n2), .Y(mode_out[0]) );
  AOI22X4 U4 ( .A0(idct_ready), .A1(mode_delay2[0]), .B0(n3), .B1(mode_out[0]), 
        .Y(n2) );
  NOR2BX4 U5 ( .AN(mode_out[1]), .B(idct_ready), .Y(mode_out[1]) );
  idct4_shift12_add2048 idct4_cal ( .clk(clk), .rstn(rstn), .mode(mode), 
        .start(start), .x0(x0), .x1(x1), .x2(x2), .x3(x3), .y0(y0_idct4), .y1(
        y1_idct4), .y2(y2_idct4), .y3(y3_idct4), .idct4_ready(idct4_ready) );
  idct8_shift12_add2048 idct8_cal ( .clk(clk), .rstn(rstn), .mode(mode), 
        .start(idct4_ready), .x0(y0_idct4), .x1(y1_idct4), .x2(y2_idct4), .x3(
        y3_idct4), .x4(x4), .x5(x5), .x6(x6), .x7(x7), .y0({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, y0_idct8}), .y1({
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, y1_idct8}), .y2({
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, y2_idct8}), .y3({
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, y3_idct8}), .y4({
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, y4_idct8}), .y5({
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, y5_idct8}), .y6({
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, y6_idct8}), .y7({
        SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75, 
        SYNOPSYS_UNCONNECTED__76, SYNOPSYS_UNCONNECTED__77, 
        SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79, y7_idct8}), 
        .idct8_ready(idct8_ready) );
  DFFRHQX1 mode_delay2_reg_1_ ( .D(mode_delay1[1]), .CK(clk), .RN(rstn), .Q(
        mode_delay2[1]) );
  DFFRHQX1 mode_delay2_reg_0_ ( .D(mode_delay1[0]), .CK(clk), .RN(rstn), .Q(
        mode_delay2[0]) );
  DFFRHQX1 mode_delay1_reg_1_ ( .D(mode[1]), .CK(clk), .RN(rstn), .Q(
        mode_delay1[1]) );
  DFFRHQX1 mode_delay1_reg_0_ ( .D(mode[0]), .CK(clk), .RN(rstn), .Q(
        mode_delay1[0]) );
  INVX1 U6 ( .A(1'b1), .Y(y15[0]) );
  INVX1 U8 ( .A(1'b1), .Y(y15[1]) );
  INVX1 U10 ( .A(1'b1), .Y(y15[2]) );
  INVX1 U12 ( .A(1'b1), .Y(y15[3]) );
  INVX1 U14 ( .A(1'b1), .Y(y15[4]) );
  INVX1 U16 ( .A(1'b1), .Y(y15[5]) );
  INVX1 U18 ( .A(1'b1), .Y(y15[6]) );
  INVX1 U20 ( .A(1'b1), .Y(y15[7]) );
  INVX1 U22 ( .A(1'b1), .Y(y15[8]) );
  INVX1 U24 ( .A(1'b1), .Y(y15[9]) );
  INVX1 U26 ( .A(1'b1), .Y(y15[10]) );
  INVX1 U28 ( .A(1'b1), .Y(y15[11]) );
  INVX1 U30 ( .A(1'b1), .Y(y15[12]) );
  INVX1 U32 ( .A(1'b1), .Y(y15[13]) );
  INVX1 U34 ( .A(1'b1), .Y(y15[14]) );
  INVX1 U36 ( .A(1'b1), .Y(y15[15]) );
  INVX1 U38 ( .A(1'b1), .Y(y14[0]) );
  INVX1 U40 ( .A(1'b1), .Y(y14[1]) );
  INVX1 U42 ( .A(1'b1), .Y(y14[2]) );
  INVX1 U44 ( .A(1'b1), .Y(y14[3]) );
  INVX1 U46 ( .A(1'b1), .Y(y14[4]) );
  INVX1 U48 ( .A(1'b1), .Y(y14[5]) );
  INVX1 U50 ( .A(1'b1), .Y(y14[6]) );
  INVX1 U52 ( .A(1'b1), .Y(y14[7]) );
  INVX1 U54 ( .A(1'b1), .Y(y14[8]) );
  INVX1 U56 ( .A(1'b1), .Y(y14[9]) );
  INVX1 U58 ( .A(1'b1), .Y(y14[10]) );
  INVX1 U60 ( .A(1'b1), .Y(y14[11]) );
  INVX1 U62 ( .A(1'b1), .Y(y14[12]) );
  INVX1 U64 ( .A(1'b1), .Y(y14[13]) );
  INVX1 U66 ( .A(1'b1), .Y(y14[14]) );
  INVX1 U68 ( .A(1'b1), .Y(y14[15]) );
  INVX1 U70 ( .A(1'b1), .Y(y13[0]) );
  INVX1 U72 ( .A(1'b1), .Y(y13[1]) );
  INVX1 U74 ( .A(1'b1), .Y(y13[2]) );
  INVX1 U76 ( .A(1'b1), .Y(y13[3]) );
  INVX1 U78 ( .A(1'b1), .Y(y13[4]) );
  INVX1 U80 ( .A(1'b1), .Y(y13[5]) );
  INVX1 U82 ( .A(1'b1), .Y(y13[6]) );
  INVX1 U84 ( .A(1'b1), .Y(y13[7]) );
  INVX1 U86 ( .A(1'b1), .Y(y13[8]) );
  INVX1 U88 ( .A(1'b1), .Y(y13[9]) );
  INVX1 U90 ( .A(1'b1), .Y(y13[10]) );
  INVX1 U92 ( .A(1'b1), .Y(y13[11]) );
  INVX1 U94 ( .A(1'b1), .Y(y13[12]) );
  INVX1 U96 ( .A(1'b1), .Y(y13[13]) );
  INVX1 U98 ( .A(1'b1), .Y(y13[14]) );
  INVX1 U100 ( .A(1'b1), .Y(y13[15]) );
  INVX1 U102 ( .A(1'b1), .Y(y12[0]) );
  INVX1 U104 ( .A(1'b1), .Y(y12[1]) );
  INVX1 U106 ( .A(1'b1), .Y(y12[2]) );
  INVX1 U108 ( .A(1'b1), .Y(y12[3]) );
  INVX1 U110 ( .A(1'b1), .Y(y12[4]) );
  INVX1 U112 ( .A(1'b1), .Y(y12[5]) );
  INVX1 U114 ( .A(1'b1), .Y(y12[6]) );
  INVX1 U116 ( .A(1'b1), .Y(y12[7]) );
  INVX1 U118 ( .A(1'b1), .Y(y12[8]) );
  INVX1 U120 ( .A(1'b1), .Y(y12[9]) );
  INVX1 U122 ( .A(1'b1), .Y(y12[10]) );
  INVX1 U124 ( .A(1'b1), .Y(y12[11]) );
  INVX1 U126 ( .A(1'b1), .Y(y12[12]) );
  INVX1 U128 ( .A(1'b1), .Y(y12[13]) );
  INVX1 U130 ( .A(1'b1), .Y(y12[14]) );
  INVX1 U132 ( .A(1'b1), .Y(y12[15]) );
  INVX1 U134 ( .A(1'b1), .Y(y11[0]) );
  INVX1 U136 ( .A(1'b1), .Y(y11[1]) );
  INVX1 U138 ( .A(1'b1), .Y(y11[2]) );
  INVX1 U140 ( .A(1'b1), .Y(y11[3]) );
  INVX1 U142 ( .A(1'b1), .Y(y11[4]) );
  INVX1 U144 ( .A(1'b1), .Y(y11[5]) );
  INVX1 U146 ( .A(1'b1), .Y(y11[6]) );
  INVX1 U148 ( .A(1'b1), .Y(y11[7]) );
  INVX1 U150 ( .A(1'b1), .Y(y11[8]) );
  INVX1 U152 ( .A(1'b1), .Y(y11[9]) );
  INVX1 U154 ( .A(1'b1), .Y(y11[10]) );
  INVX1 U156 ( .A(1'b1), .Y(y11[11]) );
  INVX1 U158 ( .A(1'b1), .Y(y11[12]) );
  INVX1 U160 ( .A(1'b1), .Y(y11[13]) );
  INVX1 U162 ( .A(1'b1), .Y(y11[14]) );
  INVX1 U164 ( .A(1'b1), .Y(y11[15]) );
  INVX1 U166 ( .A(1'b1), .Y(y10[0]) );
  INVX1 U168 ( .A(1'b1), .Y(y10[1]) );
  INVX1 U170 ( .A(1'b1), .Y(y10[2]) );
  INVX1 U172 ( .A(1'b1), .Y(y10[3]) );
  INVX1 U174 ( .A(1'b1), .Y(y10[4]) );
  INVX1 U176 ( .A(1'b1), .Y(y10[5]) );
  INVX1 U178 ( .A(1'b1), .Y(y10[6]) );
  INVX1 U180 ( .A(1'b1), .Y(y10[7]) );
  INVX1 U182 ( .A(1'b1), .Y(y10[8]) );
  INVX1 U184 ( .A(1'b1), .Y(y10[9]) );
  INVX1 U186 ( .A(1'b1), .Y(y10[10]) );
  INVX1 U188 ( .A(1'b1), .Y(y10[11]) );
  INVX1 U190 ( .A(1'b1), .Y(y10[12]) );
  INVX1 U192 ( .A(1'b1), .Y(y10[13]) );
  INVX1 U194 ( .A(1'b1), .Y(y10[14]) );
  INVX1 U196 ( .A(1'b1), .Y(y10[15]) );
  INVX1 U198 ( .A(1'b1), .Y(y9[0]) );
  INVX1 U200 ( .A(1'b1), .Y(y9[1]) );
  INVX1 U202 ( .A(1'b1), .Y(y9[2]) );
  INVX1 U204 ( .A(1'b1), .Y(y9[3]) );
  INVX1 U206 ( .A(1'b1), .Y(y9[4]) );
  INVX1 U208 ( .A(1'b1), .Y(y9[5]) );
  INVX1 U210 ( .A(1'b1), .Y(y9[6]) );
  INVX1 U212 ( .A(1'b1), .Y(y9[7]) );
  INVX1 U214 ( .A(1'b1), .Y(y9[8]) );
  INVX1 U216 ( .A(1'b1), .Y(y9[9]) );
  INVX1 U218 ( .A(1'b1), .Y(y9[10]) );
  INVX1 U220 ( .A(1'b1), .Y(y9[11]) );
  INVX1 U222 ( .A(1'b1), .Y(y9[12]) );
  INVX1 U224 ( .A(1'b1), .Y(y9[13]) );
  INVX1 U226 ( .A(1'b1), .Y(y9[14]) );
  INVX1 U228 ( .A(1'b1), .Y(y9[15]) );
  INVX1 U230 ( .A(1'b1), .Y(y8[0]) );
  INVX1 U232 ( .A(1'b1), .Y(y8[1]) );
  INVX1 U234 ( .A(1'b1), .Y(y8[2]) );
  INVX1 U236 ( .A(1'b1), .Y(y8[3]) );
  INVX1 U238 ( .A(1'b1), .Y(y8[4]) );
  INVX1 U240 ( .A(1'b1), .Y(y8[5]) );
  INVX1 U242 ( .A(1'b1), .Y(y8[6]) );
  INVX1 U244 ( .A(1'b1), .Y(y8[7]) );
  INVX1 U246 ( .A(1'b1), .Y(y8[8]) );
  INVX1 U248 ( .A(1'b1), .Y(y8[9]) );
  INVX1 U250 ( .A(1'b1), .Y(y8[10]) );
  INVX1 U252 ( .A(1'b1), .Y(y8[11]) );
  INVX1 U254 ( .A(1'b1), .Y(y8[12]) );
  INVX1 U256 ( .A(1'b1), .Y(y8[13]) );
  INVX1 U258 ( .A(1'b1), .Y(y8[14]) );
  INVX1 U260 ( .A(1'b1), .Y(y8[15]) );
  INVX1 U262 ( .A(n327), .Y(n325) );
  INVX1 U263 ( .A(n332), .Y(n329) );
  INVX1 U264 ( .A(n332), .Y(n330) );
  INVX1 U265 ( .A(n327), .Y(n326) );
  INVX1 U266 ( .A(n332), .Y(n331) );
  INVX1 U267 ( .A(n3), .Y(idct_ready) );
  INVX1 U268 ( .A(n6), .Y(n327) );
  INVX1 U269 ( .A(n332), .Y(n328) );
  INVX1 U270 ( .A(n4), .Y(n332) );
  INVX1 U271 ( .A(n64), .Y(y0[14]) );
  AOI22X1 U272 ( .A0(y0_idct8[14]), .A1(n328), .B0(y0_idct4[14]), .B1(n325), 
        .Y(n64) );
  INVX1 U273 ( .A(n63), .Y(y0[15]) );
  AOI22X1 U274 ( .A0(y0_idct8[15]), .A1(n328), .B0(y0_idct4[15]), .B1(n325), 
        .Y(n63) );
  INVX1 U275 ( .A(n48), .Y(y1[14]) );
  AOI22X1 U276 ( .A0(y1_idct8[14]), .A1(n329), .B0(y1_idct4[14]), .B1(n326), 
        .Y(n48) );
  INVX1 U277 ( .A(n47), .Y(y1[15]) );
  AOI22X1 U278 ( .A0(y1_idct8[15]), .A1(n330), .B0(y1_idct4[15]), .B1(n326), 
        .Y(n47) );
  INVX1 U279 ( .A(n32), .Y(y2[14]) );
  AOI22X1 U280 ( .A0(y2_idct8[14]), .A1(n329), .B0(y2_idct4[14]), .B1(n326), 
        .Y(n32) );
  INVX1 U281 ( .A(n31), .Y(y2[15]) );
  AOI22X1 U282 ( .A0(y2_idct8[15]), .A1(n329), .B0(y2_idct4[15]), .B1(n326), 
        .Y(n31) );
  INVX1 U283 ( .A(n16), .Y(y3[14]) );
  AOI22X1 U284 ( .A0(y3_idct8[14]), .A1(n330), .B0(y3_idct4[14]), .B1(n326), 
        .Y(n16) );
  INVX1 U285 ( .A(n15), .Y(y3[15]) );
  AOI22X1 U286 ( .A0(y3_idct8[15]), .A1(n330), .B0(y3_idct4[15]), .B1(n6), .Y(
        n15) );
  AND2X2 U287 ( .A(y4_idct8[15]), .B(n331), .Y(y4[15]) );
  AND2X2 U288 ( .A(y5_idct8[15]), .B(n331), .Y(y5[15]) );
  AND2X2 U289 ( .A(y6_idct8[15]), .B(n329), .Y(y6[15]) );
  AND2X2 U290 ( .A(y7_idct8[15]), .B(n4), .Y(y7[15]) );
  INVX1 U291 ( .A(n65), .Y(y0[13]) );
  AOI22X1 U292 ( .A0(y0_idct8[13]), .A1(n328), .B0(y0_idct4[13]), .B1(n325), 
        .Y(n65) );
  INVX1 U293 ( .A(n49), .Y(y1[13]) );
  AOI22X1 U294 ( .A0(y1_idct8[13]), .A1(n329), .B0(y1_idct4[13]), .B1(n326), 
        .Y(n49) );
  INVX1 U295 ( .A(n33), .Y(y2[13]) );
  AOI22X1 U296 ( .A0(y2_idct8[13]), .A1(n330), .B0(y2_idct4[13]), .B1(n326), 
        .Y(n33) );
  INVX1 U297 ( .A(n17), .Y(y3[13]) );
  AOI22X1 U298 ( .A0(y3_idct8[13]), .A1(n330), .B0(y3_idct4[13]), .B1(n326), 
        .Y(n17) );
  AOI22X1 U299 ( .A0(idct8_ready), .A1(n328), .B0(idct4_ready), .B1(n325), .Y(
        n3) );
  INVX1 U300 ( .A(n55), .Y(y0[8]) );
  AOI22X1 U301 ( .A0(y0_idct8[8]), .A1(n330), .B0(y0_idct4[8]), .B1(n326), .Y(
        n55) );
  INVX1 U302 ( .A(n54), .Y(y0[9]) );
  AOI22X1 U303 ( .A0(y0_idct8[9]), .A1(n329), .B0(y0_idct4[9]), .B1(n326), .Y(
        n54) );
  INVX1 U304 ( .A(n39), .Y(y1[8]) );
  AOI22X1 U305 ( .A0(y1_idct8[8]), .A1(n330), .B0(y1_idct4[8]), .B1(n6), .Y(
        n39) );
  INVX1 U306 ( .A(n38), .Y(y1[9]) );
  AOI22X1 U307 ( .A0(y1_idct8[9]), .A1(n330), .B0(y1_idct4[9]), .B1(n6), .Y(
        n38) );
  INVX1 U308 ( .A(n23), .Y(y2[8]) );
  AOI22X1 U309 ( .A0(y2_idct8[8]), .A1(n329), .B0(y2_idct4[8]), .B1(n326), .Y(
        n23) );
  INVX1 U310 ( .A(n22), .Y(y2[9]) );
  AOI22X1 U311 ( .A0(y2_idct8[9]), .A1(n329), .B0(y2_idct4[9]), .B1(n326), .Y(
        n22) );
  AND2X2 U312 ( .A(y7_idct8[13]), .B(n4), .Y(y7[13]) );
  INVX1 U313 ( .A(n7), .Y(y3[8]) );
  AOI22X1 U314 ( .A0(y3_idct8[8]), .A1(n330), .B0(y3_idct4[8]), .B1(n6), .Y(n7) );
  INVX1 U315 ( .A(n5), .Y(y3[9]) );
  AOI22X1 U316 ( .A0(y3_idct8[9]), .A1(n330), .B0(y3_idct4[9]), .B1(n6), .Y(n5) );
  NOR2BX1 U317 ( .AN(mode_delay2[0]), .B(mode_delay2[1]), .Y(n4) );
  AND2X2 U318 ( .A(y4_idct8[11]), .B(n331), .Y(y4[11]) );
  AND2X2 U319 ( .A(y4_idct8[12]), .B(n331), .Y(y4[12]) );
  AND2X2 U320 ( .A(y4_idct8[14]), .B(n331), .Y(y4[14]) );
  AND2X2 U321 ( .A(y5_idct8[11]), .B(n331), .Y(y5[11]) );
  AND2X2 U322 ( .A(y5_idct8[12]), .B(n331), .Y(y5[12]) );
  AND2X2 U323 ( .A(y5_idct8[14]), .B(n331), .Y(y5[14]) );
  AND2X2 U324 ( .A(y6_idct8[11]), .B(n330), .Y(y6[11]) );
  AND2X2 U325 ( .A(y6_idct8[12]), .B(n330), .Y(y6[12]) );
  AND2X2 U326 ( .A(y6_idct8[14]), .B(n330), .Y(y6[14]) );
  NOR2X1 U327 ( .A(mode_delay2[0]), .B(mode_delay2[1]), .Y(n6) );
  AND2X2 U328 ( .A(y7_idct8[10]), .B(n4), .Y(y7[10]) );
  AND2X2 U329 ( .A(y7_idct8[11]), .B(n4), .Y(y7[11]) );
  AND2X2 U330 ( .A(y7_idct8[12]), .B(n4), .Y(y7[12]) );
  AND2X2 U331 ( .A(y7_idct8[14]), .B(n4), .Y(y7[14]) );
  INVX1 U332 ( .A(n68), .Y(y0[10]) );
  AOI22X1 U333 ( .A0(y0_idct8[10]), .A1(n328), .B0(y0_idct4[10]), .B1(n325), 
        .Y(n68) );
  INVX1 U334 ( .A(n67), .Y(y0[11]) );
  AOI22X1 U335 ( .A0(y0_idct8[11]), .A1(n328), .B0(y0_idct4[11]), .B1(n325), 
        .Y(n67) );
  INVX1 U336 ( .A(n66), .Y(y0[12]) );
  AOI22X1 U337 ( .A0(y0_idct8[12]), .A1(n328), .B0(y0_idct4[12]), .B1(n325), 
        .Y(n66) );
  INVX1 U338 ( .A(n52), .Y(y1[10]) );
  AOI22X1 U339 ( .A0(y1_idct8[10]), .A1(n330), .B0(y1_idct4[10]), .B1(n326), 
        .Y(n52) );
  INVX1 U340 ( .A(n51), .Y(y1[11]) );
  AOI22X1 U341 ( .A0(y1_idct8[11]), .A1(n329), .B0(y1_idct4[11]), .B1(n326), 
        .Y(n51) );
  INVX1 U342 ( .A(n50), .Y(y1[12]) );
  AOI22X1 U343 ( .A0(y1_idct8[12]), .A1(n330), .B0(y1_idct4[12]), .B1(n326), 
        .Y(n50) );
  INVX1 U344 ( .A(n36), .Y(y2[10]) );
  AOI22X1 U345 ( .A0(y2_idct8[10]), .A1(n329), .B0(y2_idct4[10]), .B1(n6), .Y(
        n36) );
  INVX1 U346 ( .A(n35), .Y(y2[11]) );
  AOI22X1 U347 ( .A0(y2_idct8[11]), .A1(n329), .B0(y2_idct4[11]), .B1(n6), .Y(
        n35) );
  INVX1 U348 ( .A(n34), .Y(y2[12]) );
  AOI22X1 U349 ( .A0(y2_idct8[12]), .A1(n330), .B0(y2_idct4[12]), .B1(n326), 
        .Y(n34) );
  INVX1 U350 ( .A(n20), .Y(y3[10]) );
  AOI22X1 U351 ( .A0(y3_idct8[10]), .A1(n329), .B0(y3_idct4[10]), .B1(n326), 
        .Y(n20) );
  INVX1 U352 ( .A(n19), .Y(y3[11]) );
  AOI22X1 U353 ( .A0(y3_idct8[11]), .A1(n329), .B0(y3_idct4[11]), .B1(n6), .Y(
        n19) );
  INVX1 U354 ( .A(n18), .Y(y3[12]) );
  AOI22X1 U355 ( .A0(y3_idct8[12]), .A1(n330), .B0(y3_idct4[12]), .B1(n6), .Y(
        n18) );
  AND2X2 U356 ( .A(y4_idct8[10]), .B(n331), .Y(y4[10]) );
  AND2X2 U357 ( .A(y4_idct8[13]), .B(n331), .Y(y4[13]) );
  AND2X2 U358 ( .A(y5_idct8[10]), .B(n331), .Y(y5[10]) );
  AND2X2 U359 ( .A(y5_idct8[13]), .B(n331), .Y(y5[13]) );
  AND2X2 U360 ( .A(y6_idct8[10]), .B(n329), .Y(y6[10]) );
  AND2X2 U361 ( .A(y6_idct8[13]), .B(n329), .Y(y6[13]) );
  INVX1 U362 ( .A(n62), .Y(y0[1]) );
  AOI22X1 U363 ( .A0(y0_idct8[1]), .A1(n328), .B0(y0_idct4[1]), .B1(n325), .Y(
        n62) );
  INVX1 U364 ( .A(n61), .Y(y0[2]) );
  AOI22X1 U365 ( .A0(y0_idct8[2]), .A1(n328), .B0(y0_idct4[2]), .B1(n325), .Y(
        n61) );
  INVX1 U366 ( .A(n60), .Y(y0[3]) );
  AOI22X1 U367 ( .A0(y0_idct8[3]), .A1(n328), .B0(y0_idct4[3]), .B1(n325), .Y(
        n60) );
  INVX1 U368 ( .A(n58), .Y(y0[5]) );
  AOI22X1 U369 ( .A0(y0_idct8[5]), .A1(n328), .B0(y0_idct4[5]), .B1(n326), .Y(
        n58) );
  INVX1 U370 ( .A(n46), .Y(y1[1]) );
  AOI22X1 U371 ( .A0(y1_idct8[1]), .A1(n329), .B0(y1_idct4[1]), .B1(n6), .Y(
        n46) );
  INVX1 U372 ( .A(n45), .Y(y1[2]) );
  AOI22X1 U373 ( .A0(y1_idct8[2]), .A1(n330), .B0(y1_idct4[2]), .B1(n6), .Y(
        n45) );
  INVX1 U374 ( .A(n44), .Y(y1[3]) );
  AOI22X1 U375 ( .A0(y1_idct8[3]), .A1(n329), .B0(y1_idct4[3]), .B1(n6), .Y(
        n44) );
  INVX1 U376 ( .A(n42), .Y(y1[5]) );
  AOI22X1 U377 ( .A0(y1_idct8[5]), .A1(n330), .B0(y1_idct4[5]), .B1(n6), .Y(
        n42) );
  INVX1 U378 ( .A(n30), .Y(y2[1]) );
  AOI22X1 U379 ( .A0(y2_idct8[1]), .A1(n329), .B0(y2_idct4[1]), .B1(n326), .Y(
        n30) );
  INVX1 U380 ( .A(n29), .Y(y2[2]) );
  AOI22X1 U381 ( .A0(y2_idct8[2]), .A1(n329), .B0(y2_idct4[2]), .B1(n326), .Y(
        n29) );
  INVX1 U382 ( .A(n28), .Y(y2[3]) );
  AOI22X1 U383 ( .A0(y2_idct8[3]), .A1(n329), .B0(y2_idct4[3]), .B1(n326), .Y(
        n28) );
  INVX1 U384 ( .A(n26), .Y(y2[5]) );
  AOI22X1 U385 ( .A0(y2_idct8[5]), .A1(n329), .B0(y2_idct4[5]), .B1(n326), .Y(
        n26) );
  INVX1 U386 ( .A(n14), .Y(y3[1]) );
  AOI22X1 U387 ( .A0(y3_idct8[1]), .A1(n330), .B0(y3_idct4[1]), .B1(n326), .Y(
        n14) );
  INVX1 U388 ( .A(n13), .Y(y3[2]) );
  AOI22X1 U389 ( .A0(y3_idct8[2]), .A1(n330), .B0(y3_idct4[2]), .B1(n6), .Y(
        n13) );
  INVX1 U390 ( .A(n12), .Y(y3[3]) );
  AOI22X1 U391 ( .A0(y3_idct8[3]), .A1(n330), .B0(y3_idct4[3]), .B1(n326), .Y(
        n12) );
  INVX1 U392 ( .A(n10), .Y(y3[5]) );
  AOI22X1 U393 ( .A0(y3_idct8[5]), .A1(n330), .B0(y3_idct4[5]), .B1(n326), .Y(
        n10) );
  INVX1 U394 ( .A(n8), .Y(y3[7]) );
  AOI22X1 U395 ( .A0(y3_idct8[7]), .A1(n330), .B0(y3_idct4[7]), .B1(n6), .Y(n8) );
  INVX1 U396 ( .A(n69), .Y(y0[0]) );
  AOI22X1 U397 ( .A0(y0_idct8[0]), .A1(n328), .B0(y0_idct4[0]), .B1(n325), .Y(
        n69) );
  INVX1 U398 ( .A(n59), .Y(y0[4]) );
  AOI22X1 U399 ( .A0(y0_idct8[4]), .A1(n328), .B0(y0_idct4[4]), .B1(n325), .Y(
        n59) );
  INVX1 U400 ( .A(n57), .Y(y0[6]) );
  AOI22X1 U401 ( .A0(y0_idct8[6]), .A1(n330), .B0(y0_idct4[6]), .B1(n326), .Y(
        n57) );
  INVX1 U402 ( .A(n56), .Y(y0[7]) );
  AOI22X1 U403 ( .A0(y0_idct8[7]), .A1(n329), .B0(y0_idct4[7]), .B1(n326), .Y(
        n56) );
  INVX1 U404 ( .A(n53), .Y(y1[0]) );
  AOI22X1 U405 ( .A0(y1_idct8[0]), .A1(n329), .B0(y1_idct4[0]), .B1(n326), .Y(
        n53) );
  INVX1 U406 ( .A(n43), .Y(y1[4]) );
  AOI22X1 U407 ( .A0(y1_idct8[4]), .A1(n330), .B0(y1_idct4[4]), .B1(n6), .Y(
        n43) );
  INVX1 U408 ( .A(n41), .Y(y1[6]) );
  AOI22X1 U409 ( .A0(y1_idct8[6]), .A1(n329), .B0(y1_idct4[6]), .B1(n6), .Y(
        n41) );
  INVX1 U410 ( .A(n40), .Y(y1[7]) );
  AOI22X1 U411 ( .A0(y1_idct8[7]), .A1(n329), .B0(y1_idct4[7]), .B1(n6), .Y(
        n40) );
  INVX1 U412 ( .A(n37), .Y(y2[0]) );
  AOI22X1 U413 ( .A0(y2_idct8[0]), .A1(n330), .B0(y2_idct4[0]), .B1(n6), .Y(
        n37) );
  INVX1 U414 ( .A(n27), .Y(y2[4]) );
  AOI22X1 U415 ( .A0(y2_idct8[4]), .A1(n329), .B0(y2_idct4[4]), .B1(n326), .Y(
        n27) );
  INVX1 U416 ( .A(n25), .Y(y2[6]) );
  AOI22X1 U417 ( .A0(y2_idct8[6]), .A1(n329), .B0(y2_idct4[6]), .B1(n326), .Y(
        n25) );
  INVX1 U418 ( .A(n24), .Y(y2[7]) );
  AOI22X1 U419 ( .A0(y2_idct8[7]), .A1(n329), .B0(y2_idct4[7]), .B1(n325), .Y(
        n24) );
  INVX1 U420 ( .A(n21), .Y(y3[0]) );
  AOI22X1 U421 ( .A0(y3_idct8[0]), .A1(n329), .B0(y3_idct4[0]), .B1(n326), .Y(
        n21) );
  INVX1 U422 ( .A(n11), .Y(y3[4]) );
  AOI22X1 U423 ( .A0(y3_idct8[4]), .A1(n330), .B0(y3_idct4[4]), .B1(n6), .Y(
        n11) );
  INVX1 U424 ( .A(n9), .Y(y3[6]) );
  AOI22X1 U425 ( .A0(y3_idct8[6]), .A1(n330), .B0(y3_idct4[6]), .B1(n326), .Y(
        n9) );
  AND2X2 U426 ( .A(y4_idct8[4]), .B(n331), .Y(y4[4]) );
  AND2X2 U427 ( .A(y4_idct8[5]), .B(n331), .Y(y4[5]) );
  AND2X2 U428 ( .A(y4_idct8[6]), .B(n331), .Y(y4[6]) );
  AND2X2 U429 ( .A(y4_idct8[7]), .B(n331), .Y(y4[7]) );
  AND2X2 U430 ( .A(y4_idct8[8]), .B(n331), .Y(y4[8]) );
  AND2X2 U431 ( .A(y4_idct8[9]), .B(n331), .Y(y4[9]) );
  AND2X2 U432 ( .A(y5_idct8[0]), .B(n331), .Y(y5[0]) );
  AND2X2 U433 ( .A(y5_idct8[1]), .B(n331), .Y(y5[1]) );
  AND2X2 U434 ( .A(y5_idct8[2]), .B(n331), .Y(y5[2]) );
  AND2X2 U435 ( .A(y5_idct8[3]), .B(n331), .Y(y5[3]) );
  AND2X2 U436 ( .A(y5_idct8[4]), .B(n331), .Y(y5[4]) );
  AND2X2 U437 ( .A(y5_idct8[5]), .B(n331), .Y(y5[5]) );
  AND2X2 U438 ( .A(y5_idct8[6]), .B(n331), .Y(y5[6]) );
  AND2X2 U439 ( .A(y5_idct8[7]), .B(n331), .Y(y5[7]) );
  AND2X2 U440 ( .A(y5_idct8[8]), .B(n331), .Y(y5[8]) );
  AND2X2 U441 ( .A(y5_idct8[9]), .B(n331), .Y(y5[9]) );
  AND2X2 U442 ( .A(y6_idct8[0]), .B(n330), .Y(y6[0]) );
  AND2X2 U443 ( .A(y6_idct8[1]), .B(n330), .Y(y6[1]) );
  AND2X2 U444 ( .A(y6_idct8[2]), .B(n329), .Y(y6[2]) );
  AND2X2 U445 ( .A(y6_idct8[3]), .B(n329), .Y(y6[3]) );
  AND2X2 U446 ( .A(y6_idct8[4]), .B(n329), .Y(y6[4]) );
  AND2X2 U447 ( .A(y6_idct8[5]), .B(n328), .Y(y6[5]) );
  AND2X2 U448 ( .A(y6_idct8[6]), .B(n4), .Y(y6[6]) );
  AND2X2 U449 ( .A(y6_idct8[7]), .B(n4), .Y(y6[7]) );
  AND2X2 U450 ( .A(y6_idct8[8]), .B(n330), .Y(y6[8]) );
  AND2X2 U451 ( .A(y6_idct8[9]), .B(n4), .Y(y6[9]) );
  AND2X2 U452 ( .A(y4_idct8[0]), .B(n331), .Y(y4[0]) );
  AND2X2 U453 ( .A(y4_idct8[1]), .B(n331), .Y(y4[1]) );
  AND2X2 U454 ( .A(y4_idct8[2]), .B(n331), .Y(y4[2]) );
  AND2X2 U455 ( .A(y4_idct8[3]), .B(n331), .Y(y4[3]) );
  AND2X2 U456 ( .A(y7_idct8[0]), .B(n4), .Y(y7[0]) );
  AND2X2 U457 ( .A(y7_idct8[1]), .B(n4), .Y(y7[1]) );
  AND2X2 U458 ( .A(y7_idct8[2]), .B(n4), .Y(y7[2]) );
  AND2X2 U459 ( .A(y7_idct8[3]), .B(n4), .Y(y7[3]) );
  AND2X2 U460 ( .A(y7_idct8[4]), .B(n4), .Y(y7[4]) );
  AND2X2 U461 ( .A(y7_idct8[5]), .B(n4), .Y(y7[5]) );
  AND2X2 U462 ( .A(y7_idct8[6]), .B(n4), .Y(y7[6]) );
  AND2X2 U463 ( .A(y7_idct8[7]), .B(n4), .Y(y7[7]) );
  AND2X2 U464 ( .A(y7_idct8[8]), .B(n4), .Y(y7[8]) );
  AND2X2 U465 ( .A(y7_idct8[9]), .B(n4), .Y(y7[9]) );
endmodule


module p2s_1 ( clk, rstn, start, mode, cal_result, dout, p2s_ready, mode_out
 );
  input [1:0] mode;
  input [127:0] cal_result;
  output [15:0] dout;
  output [1:0] mode_out;
  input clk, rstn, start;
  output p2s_ready;
  wire   ready8, mode_reg_0_, shift4_flag, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n209, n210, n211, n212, n213, n214, n216, n217, n218, n219, n220,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n287, n307,
         n314, n447, n448, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
         n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
         n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
         n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
         n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
         n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
         n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
         n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
         n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
         n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
         n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
         n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
         n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
         n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
         n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
         n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
         n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
         n1266, n1267, n1268, n1269;
  wire   [5:0] start_reg4;
  wire   [143:0] result_reg4;
  wire   [127:0] result_reg8;

  AND2X4 U4 ( .A(mode_out[1]), .B(n1123), .Y(mode_out[1]) );
  OAI2BB1X4 U5 ( .A0N(n679), .A1N(mode_out[0]), .B0(n673), .Y(mode_out[0]) );
  DFFRHQX1 result_reg8_reg_111_ ( .D(n881), .CK(clk), .RN(rstn), .Q(
        result_reg8[111]) );
  DFFRHQX1 result_reg8_reg_110_ ( .D(n880), .CK(clk), .RN(rstn), .Q(
        result_reg8[110]) );
  DFFRHQX1 result_reg8_reg_109_ ( .D(n879), .CK(clk), .RN(rstn), .Q(
        result_reg8[109]) );
  DFFRHQX1 result_reg8_reg_108_ ( .D(n878), .CK(clk), .RN(rstn), .Q(
        result_reg8[108]) );
  DFFRHQX1 result_reg8_reg_107_ ( .D(n877), .CK(clk), .RN(rstn), .Q(
        result_reg8[107]) );
  DFFRHQX1 result_reg8_reg_106_ ( .D(n876), .CK(clk), .RN(rstn), .Q(
        result_reg8[106]) );
  DFFRHQX1 result_reg8_reg_105_ ( .D(n875), .CK(clk), .RN(rstn), .Q(
        result_reg8[105]) );
  DFFRHQX1 result_reg8_reg_104_ ( .D(n874), .CK(clk), .RN(rstn), .Q(
        result_reg8[104]) );
  DFFRHQX1 result_reg8_reg_103_ ( .D(n873), .CK(clk), .RN(rstn), .Q(
        result_reg8[103]) );
  DFFRHQX1 result_reg8_reg_102_ ( .D(n872), .CK(clk), .RN(rstn), .Q(
        result_reg8[102]) );
  DFFRHQX1 result_reg8_reg_101_ ( .D(n871), .CK(clk), .RN(rstn), .Q(
        result_reg8[101]) );
  DFFRHQX1 result_reg8_reg_100_ ( .D(n870), .CK(clk), .RN(rstn), .Q(
        result_reg8[100]) );
  DFFRHQX1 result_reg8_reg_99_ ( .D(n869), .CK(clk), .RN(rstn), .Q(
        result_reg8[99]) );
  DFFRHQX1 result_reg8_reg_98_ ( .D(n868), .CK(clk), .RN(rstn), .Q(
        result_reg8[98]) );
  DFFRHQX1 result_reg8_reg_97_ ( .D(n867), .CK(clk), .RN(rstn), .Q(
        result_reg8[97]) );
  DFFRHQX1 result_reg8_reg_96_ ( .D(n866), .CK(clk), .RN(rstn), .Q(
        result_reg8[96]) );
  DFFRHQX1 result_reg8_reg_95_ ( .D(n865), .CK(clk), .RN(rstn), .Q(
        result_reg8[95]) );
  DFFRHQX1 result_reg8_reg_94_ ( .D(n864), .CK(clk), .RN(rstn), .Q(
        result_reg8[94]) );
  DFFRHQX1 result_reg8_reg_93_ ( .D(n863), .CK(clk), .RN(rstn), .Q(
        result_reg8[93]) );
  DFFRHQX1 result_reg8_reg_92_ ( .D(n862), .CK(clk), .RN(rstn), .Q(
        result_reg8[92]) );
  DFFRHQX1 result_reg8_reg_91_ ( .D(n861), .CK(clk), .RN(rstn), .Q(
        result_reg8[91]) );
  DFFRHQX1 result_reg8_reg_90_ ( .D(n860), .CK(clk), .RN(rstn), .Q(
        result_reg8[90]) );
  DFFRHQX1 result_reg8_reg_89_ ( .D(n859), .CK(clk), .RN(rstn), .Q(
        result_reg8[89]) );
  DFFRHQX1 result_reg8_reg_88_ ( .D(n858), .CK(clk), .RN(rstn), .Q(
        result_reg8[88]) );
  DFFRHQX1 result_reg8_reg_87_ ( .D(n857), .CK(clk), .RN(rstn), .Q(
        result_reg8[87]) );
  DFFRHQX1 result_reg8_reg_86_ ( .D(n856), .CK(clk), .RN(rstn), .Q(
        result_reg8[86]) );
  DFFRHQX1 result_reg8_reg_85_ ( .D(n855), .CK(clk), .RN(rstn), .Q(
        result_reg8[85]) );
  DFFRHQX1 result_reg8_reg_84_ ( .D(n854), .CK(clk), .RN(rstn), .Q(
        result_reg8[84]) );
  DFFRHQX1 result_reg8_reg_83_ ( .D(n853), .CK(clk), .RN(rstn), .Q(
        result_reg8[83]) );
  DFFRHQX1 result_reg8_reg_82_ ( .D(n852), .CK(clk), .RN(rstn), .Q(
        result_reg8[82]) );
  DFFRHQX1 result_reg8_reg_81_ ( .D(n851), .CK(clk), .RN(rstn), .Q(
        result_reg8[81]) );
  DFFRHQX1 result_reg8_reg_80_ ( .D(n850), .CK(clk), .RN(rstn), .Q(
        result_reg8[80]) );
  DFFRHQX1 start_reg4_reg_5_ ( .D(n747), .CK(clk), .RN(rstn), .Q(start_reg4[5]) );
  DFFRHQX1 start_reg4_reg_4_ ( .D(n748), .CK(clk), .RN(rstn), .Q(start_reg4[4]) );
  DFFRHQX1 start_reg4_reg_3_ ( .D(n749), .CK(clk), .RN(rstn), .Q(start_reg4[3]) );
  DFFRHQX1 start_reg4_reg_2_ ( .D(n750), .CK(clk), .RN(rstn), .Q(start_reg4[2]) );
  DFFRHQX1 start_reg4_reg_1_ ( .D(n751), .CK(clk), .RN(rstn), .Q(start_reg4[1]) );
  DFFRHQX1 result_reg4_reg_95_ ( .D(n784), .CK(clk), .RN(rstn), .Q(
        result_reg4[95]) );
  DFFRHQX1 result_reg4_reg_94_ ( .D(n782), .CK(clk), .RN(rstn), .Q(
        result_reg4[94]) );
  DFFRHQX1 result_reg4_reg_93_ ( .D(n780), .CK(clk), .RN(rstn), .Q(
        result_reg4[93]) );
  DFFRHQX1 result_reg4_reg_92_ ( .D(n778), .CK(clk), .RN(rstn), .Q(
        result_reg4[92]) );
  DFFRHQX1 result_reg4_reg_91_ ( .D(n776), .CK(clk), .RN(rstn), .Q(
        result_reg4[91]) );
  DFFRHQX1 result_reg4_reg_90_ ( .D(n774), .CK(clk), .RN(rstn), .Q(
        result_reg4[90]) );
  DFFRHQX1 result_reg4_reg_89_ ( .D(n772), .CK(clk), .RN(rstn), .Q(
        result_reg4[89]) );
  DFFRHQX1 result_reg4_reg_88_ ( .D(n770), .CK(clk), .RN(rstn), .Q(
        result_reg4[88]) );
  DFFRHQX1 result_reg4_reg_87_ ( .D(n768), .CK(clk), .RN(rstn), .Q(
        result_reg4[87]) );
  DFFRHQX1 result_reg4_reg_86_ ( .D(n766), .CK(clk), .RN(rstn), .Q(
        result_reg4[86]) );
  DFFRHQX1 result_reg4_reg_85_ ( .D(n764), .CK(clk), .RN(rstn), .Q(
        result_reg4[85]) );
  DFFRHQX1 result_reg4_reg_84_ ( .D(n762), .CK(clk), .RN(rstn), .Q(
        result_reg4[84]) );
  DFFRHQX1 result_reg4_reg_83_ ( .D(n760), .CK(clk), .RN(rstn), .Q(
        result_reg4[83]) );
  DFFRHQX1 result_reg4_reg_82_ ( .D(n758), .CK(clk), .RN(rstn), .Q(
        result_reg4[82]) );
  DFFRHQX1 result_reg4_reg_81_ ( .D(n756), .CK(clk), .RN(rstn), .Q(
        result_reg4[81]) );
  DFFRHQX1 result_reg4_reg_80_ ( .D(n754), .CK(clk), .RN(rstn), .Q(
        result_reg4[80]) );
  DFFRHQX1 result_reg4_reg_79_ ( .D(n785), .CK(clk), .RN(rstn), .Q(
        result_reg4[79]) );
  DFFRHQX1 result_reg4_reg_78_ ( .D(n783), .CK(clk), .RN(rstn), .Q(
        result_reg4[78]) );
  DFFRHQX1 result_reg4_reg_77_ ( .D(n781), .CK(clk), .RN(rstn), .Q(
        result_reg4[77]) );
  DFFRHQX1 result_reg4_reg_76_ ( .D(n779), .CK(clk), .RN(rstn), .Q(
        result_reg4[76]) );
  DFFRHQX1 result_reg4_reg_75_ ( .D(n777), .CK(clk), .RN(rstn), .Q(
        result_reg4[75]) );
  DFFRHQX1 result_reg4_reg_74_ ( .D(n775), .CK(clk), .RN(rstn), .Q(
        result_reg4[74]) );
  DFFRHQX1 result_reg4_reg_73_ ( .D(n773), .CK(clk), .RN(rstn), .Q(
        result_reg4[73]) );
  DFFRHQX1 result_reg4_reg_72_ ( .D(n771), .CK(clk), .RN(rstn), .Q(
        result_reg4[72]) );
  DFFRHQX1 result_reg4_reg_71_ ( .D(n769), .CK(clk), .RN(rstn), .Q(
        result_reg4[71]) );
  DFFRHQX1 result_reg4_reg_70_ ( .D(n767), .CK(clk), .RN(rstn), .Q(
        result_reg4[70]) );
  DFFRHQX1 result_reg4_reg_69_ ( .D(n765), .CK(clk), .RN(rstn), .Q(
        result_reg4[69]) );
  DFFRHQX1 result_reg4_reg_68_ ( .D(n763), .CK(clk), .RN(rstn), .Q(
        result_reg4[68]) );
  DFFRHQX1 result_reg4_reg_67_ ( .D(n761), .CK(clk), .RN(rstn), .Q(
        result_reg4[67]) );
  DFFRHQX1 result_reg4_reg_66_ ( .D(n759), .CK(clk), .RN(rstn), .Q(
        result_reg4[66]) );
  DFFRHQX1 result_reg4_reg_65_ ( .D(n757), .CK(clk), .RN(rstn), .Q(
        result_reg4[65]) );
  DFFRHQX1 result_reg4_reg_64_ ( .D(n755), .CK(clk), .RN(rstn), .Q(
        result_reg4[64]) );
  DFFRHQX1 result_reg8_reg_63_ ( .D(n1253), .CK(clk), .RN(rstn), .Q(
        result_reg8[63]) );
  DFFRHQX1 result_reg8_reg_62_ ( .D(n1252), .CK(clk), .RN(rstn), .Q(
        result_reg8[62]) );
  DFFRHQX1 result_reg8_reg_61_ ( .D(n1251), .CK(clk), .RN(rstn), .Q(
        result_reg8[61]) );
  DFFRHQX1 result_reg8_reg_60_ ( .D(n1250), .CK(clk), .RN(rstn), .Q(
        result_reg8[60]) );
  DFFRHQX1 result_reg8_reg_59_ ( .D(n1249), .CK(clk), .RN(rstn), .Q(
        result_reg8[59]) );
  DFFRHQX1 result_reg8_reg_58_ ( .D(n1248), .CK(clk), .RN(rstn), .Q(
        result_reg8[58]) );
  DFFRHQX1 result_reg8_reg_57_ ( .D(n1247), .CK(clk), .RN(rstn), .Q(
        result_reg8[57]) );
  DFFRHQX1 result_reg8_reg_56_ ( .D(n1246), .CK(clk), .RN(rstn), .Q(
        result_reg8[56]) );
  DFFRHQX1 result_reg8_reg_55_ ( .D(n1245), .CK(clk), .RN(rstn), .Q(
        result_reg8[55]) );
  DFFRHQX1 result_reg8_reg_54_ ( .D(n1244), .CK(clk), .RN(rstn), .Q(
        result_reg8[54]) );
  DFFRHQX1 result_reg8_reg_53_ ( .D(n1243), .CK(clk), .RN(rstn), .Q(
        result_reg8[53]) );
  DFFRHQX1 result_reg8_reg_52_ ( .D(n1242), .CK(clk), .RN(rstn), .Q(
        result_reg8[52]) );
  DFFRHQX1 result_reg8_reg_51_ ( .D(n1241), .CK(clk), .RN(rstn), .Q(
        result_reg8[51]) );
  DFFRHQX1 result_reg8_reg_50_ ( .D(n1240), .CK(clk), .RN(rstn), .Q(
        result_reg8[50]) );
  DFFRHQX1 result_reg8_reg_49_ ( .D(n1239), .CK(clk), .RN(rstn), .Q(
        result_reg8[49]) );
  DFFRHQX1 result_reg8_reg_48_ ( .D(n1238), .CK(clk), .RN(rstn), .Q(
        result_reg8[48]) );
  DFFRHQX1 result_reg8_reg_47_ ( .D(n1237), .CK(clk), .RN(rstn), .Q(
        result_reg8[47]) );
  DFFRHQX1 result_reg8_reg_46_ ( .D(n1236), .CK(clk), .RN(rstn), .Q(
        result_reg8[46]) );
  DFFRHQX1 result_reg8_reg_45_ ( .D(n1235), .CK(clk), .RN(rstn), .Q(
        result_reg8[45]) );
  DFFRHQX1 result_reg8_reg_44_ ( .D(n1234), .CK(clk), .RN(rstn), .Q(
        result_reg8[44]) );
  DFFRHQX1 result_reg8_reg_43_ ( .D(n1233), .CK(clk), .RN(rstn), .Q(
        result_reg8[43]) );
  DFFRHQX1 result_reg8_reg_42_ ( .D(n1232), .CK(clk), .RN(rstn), .Q(
        result_reg8[42]) );
  DFFRHQX1 result_reg8_reg_41_ ( .D(n1231), .CK(clk), .RN(rstn), .Q(
        result_reg8[41]) );
  DFFRHQX1 result_reg8_reg_40_ ( .D(n1230), .CK(clk), .RN(rstn), .Q(
        result_reg8[40]) );
  DFFRHQX1 result_reg8_reg_39_ ( .D(n1229), .CK(clk), .RN(rstn), .Q(
        result_reg8[39]) );
  DFFRHQX1 result_reg8_reg_38_ ( .D(n1228), .CK(clk), .RN(rstn), .Q(
        result_reg8[38]) );
  DFFRHQX1 result_reg8_reg_37_ ( .D(n1227), .CK(clk), .RN(rstn), .Q(
        result_reg8[37]) );
  DFFRHQX1 result_reg8_reg_36_ ( .D(n1226), .CK(clk), .RN(rstn), .Q(
        result_reg8[36]) );
  DFFRHQX1 result_reg8_reg_35_ ( .D(n1225), .CK(clk), .RN(rstn), .Q(
        result_reg8[35]) );
  DFFRHQX1 result_reg8_reg_34_ ( .D(n1224), .CK(clk), .RN(rstn), .Q(
        result_reg8[34]) );
  DFFRHQX1 result_reg8_reg_33_ ( .D(n1223), .CK(clk), .RN(rstn), .Q(
        result_reg8[33]) );
  DFFRHQX1 result_reg8_reg_32_ ( .D(n1222), .CK(clk), .RN(rstn), .Q(
        result_reg8[32]) );
  DFFRHQX1 result_reg8_reg_31_ ( .D(n1221), .CK(clk), .RN(rstn), .Q(
        result_reg8[31]) );
  DFFRHQX1 result_reg8_reg_30_ ( .D(n1220), .CK(clk), .RN(rstn), .Q(
        result_reg8[30]) );
  DFFRHQX1 result_reg8_reg_29_ ( .D(n1219), .CK(clk), .RN(rstn), .Q(
        result_reg8[29]) );
  DFFRHQX1 result_reg8_reg_28_ ( .D(n1218), .CK(clk), .RN(rstn), .Q(
        result_reg8[28]) );
  DFFRHQX1 result_reg8_reg_27_ ( .D(n1217), .CK(clk), .RN(rstn), .Q(
        result_reg8[27]) );
  DFFRHQX1 result_reg8_reg_26_ ( .D(n1216), .CK(clk), .RN(rstn), .Q(
        result_reg8[26]) );
  DFFRHQX1 result_reg8_reg_25_ ( .D(n1215), .CK(clk), .RN(rstn), .Q(
        result_reg8[25]) );
  DFFRHQX1 result_reg8_reg_24_ ( .D(n1214), .CK(clk), .RN(rstn), .Q(
        result_reg8[24]) );
  DFFRHQX1 result_reg8_reg_23_ ( .D(n1213), .CK(clk), .RN(rstn), .Q(
        result_reg8[23]) );
  DFFRHQX1 result_reg8_reg_22_ ( .D(n1212), .CK(clk), .RN(rstn), .Q(
        result_reg8[22]) );
  DFFRHQX1 result_reg8_reg_21_ ( .D(n1211), .CK(clk), .RN(rstn), .Q(
        result_reg8[21]) );
  DFFRHQX1 result_reg8_reg_20_ ( .D(n1210), .CK(clk), .RN(rstn), .Q(
        result_reg8[20]) );
  DFFRHQX1 result_reg8_reg_19_ ( .D(n1209), .CK(clk), .RN(rstn), .Q(
        result_reg8[19]) );
  DFFRHQX1 result_reg8_reg_18_ ( .D(n1208), .CK(clk), .RN(rstn), .Q(
        result_reg8[18]) );
  DFFRHQX1 result_reg8_reg_17_ ( .D(n1207), .CK(clk), .RN(rstn), .Q(
        result_reg8[17]) );
  DFFRHQX1 result_reg8_reg_16_ ( .D(n1206), .CK(clk), .RN(rstn), .Q(
        result_reg8[16]) );
  DFFRHQX1 result_reg8_reg_79_ ( .D(n849), .CK(clk), .RN(rstn), .Q(
        result_reg8[79]) );
  DFFRHQX1 result_reg8_reg_78_ ( .D(n848), .CK(clk), .RN(rstn), .Q(
        result_reg8[78]) );
  DFFRHQX1 result_reg8_reg_77_ ( .D(n847), .CK(clk), .RN(rstn), .Q(
        result_reg8[77]) );
  DFFRHQX1 result_reg8_reg_76_ ( .D(n846), .CK(clk), .RN(rstn), .Q(
        result_reg8[76]) );
  DFFRHQX1 result_reg8_reg_75_ ( .D(n845), .CK(clk), .RN(rstn), .Q(
        result_reg8[75]) );
  DFFRHQX1 result_reg8_reg_74_ ( .D(n844), .CK(clk), .RN(rstn), .Q(
        result_reg8[74]) );
  DFFRHQX1 result_reg8_reg_73_ ( .D(n843), .CK(clk), .RN(rstn), .Q(
        result_reg8[73]) );
  DFFRHQX1 result_reg8_reg_72_ ( .D(n842), .CK(clk), .RN(rstn), .Q(
        result_reg8[72]) );
  DFFRHQX1 result_reg8_reg_71_ ( .D(n841), .CK(clk), .RN(rstn), .Q(
        result_reg8[71]) );
  DFFRHQX1 result_reg8_reg_70_ ( .D(n840), .CK(clk), .RN(rstn), .Q(
        result_reg8[70]) );
  DFFRHQX1 result_reg8_reg_69_ ( .D(n839), .CK(clk), .RN(rstn), .Q(
        result_reg8[69]) );
  DFFRHQX1 result_reg8_reg_68_ ( .D(n838), .CK(clk), .RN(rstn), .Q(
        result_reg8[68]) );
  DFFRHQX1 result_reg8_reg_67_ ( .D(n837), .CK(clk), .RN(rstn), .Q(
        result_reg8[67]) );
  DFFRHQX1 result_reg8_reg_66_ ( .D(n836), .CK(clk), .RN(rstn), .Q(
        result_reg8[66]) );
  DFFRHQX1 result_reg8_reg_65_ ( .D(n835), .CK(clk), .RN(rstn), .Q(
        result_reg8[65]) );
  DFFRHQX1 result_reg8_reg_64_ ( .D(n834), .CK(clk), .RN(rstn), .Q(
        result_reg8[64]) );
  DFFRHQX1 result_reg8_reg_15_ ( .D(n1205), .CK(clk), .RN(rstn), .Q(
        result_reg8[15]) );
  DFFRHQX1 result_reg8_reg_14_ ( .D(n1204), .CK(clk), .RN(rstn), .Q(
        result_reg8[14]) );
  DFFRHQX1 result_reg8_reg_13_ ( .D(n1203), .CK(clk), .RN(rstn), .Q(
        result_reg8[13]) );
  DFFRHQX1 result_reg8_reg_12_ ( .D(n1202), .CK(clk), .RN(rstn), .Q(
        result_reg8[12]) );
  DFFRHQX1 result_reg8_reg_11_ ( .D(n1201), .CK(clk), .RN(rstn), .Q(
        result_reg8[11]) );
  DFFRHQX1 result_reg8_reg_10_ ( .D(n1200), .CK(clk), .RN(rstn), .Q(
        result_reg8[10]) );
  DFFRHQX1 result_reg8_reg_9_ ( .D(n1199), .CK(clk), .RN(rstn), .Q(
        result_reg8[9]) );
  DFFRHQX1 result_reg8_reg_8_ ( .D(n1198), .CK(clk), .RN(rstn), .Q(
        result_reg8[8]) );
  DFFRHQX1 result_reg8_reg_7_ ( .D(n1197), .CK(clk), .RN(rstn), .Q(
        result_reg8[7]) );
  DFFRHQX1 result_reg8_reg_6_ ( .D(n1196), .CK(clk), .RN(rstn), .Q(
        result_reg8[6]) );
  DFFRHQX1 result_reg8_reg_5_ ( .D(n1195), .CK(clk), .RN(rstn), .Q(
        result_reg8[5]) );
  DFFRHQX1 result_reg8_reg_4_ ( .D(n1194), .CK(clk), .RN(rstn), .Q(
        result_reg8[4]) );
  DFFRHQX1 result_reg8_reg_3_ ( .D(n1193), .CK(clk), .RN(rstn), .Q(
        result_reg8[3]) );
  DFFRHQX1 result_reg8_reg_2_ ( .D(n1192), .CK(clk), .RN(rstn), .Q(
        result_reg8[2]) );
  DFFRHQX1 result_reg8_reg_1_ ( .D(n1191), .CK(clk), .RN(rstn), .Q(
        result_reg8[1]) );
  DFFRHQX1 result_reg8_reg_0_ ( .D(n1190), .CK(clk), .RN(rstn), .Q(
        result_reg8[0]) );
  DFFRHQX1 result_reg4_reg_143_ ( .D(n833), .CK(clk), .RN(rstn), .Q(
        result_reg4[143]) );
  DFFRHQX1 result_reg4_reg_142_ ( .D(n832), .CK(clk), .RN(rstn), .Q(
        result_reg4[142]) );
  DFFRHQX1 result_reg4_reg_141_ ( .D(n831), .CK(clk), .RN(rstn), .Q(
        result_reg4[141]) );
  DFFRHQX1 result_reg4_reg_140_ ( .D(n830), .CK(clk), .RN(rstn), .Q(
        result_reg4[140]) );
  DFFRHQX1 result_reg4_reg_139_ ( .D(n829), .CK(clk), .RN(rstn), .Q(
        result_reg4[139]) );
  DFFRHQX1 result_reg4_reg_138_ ( .D(n828), .CK(clk), .RN(rstn), .Q(
        result_reg4[138]) );
  DFFRHQX1 result_reg4_reg_137_ ( .D(n827), .CK(clk), .RN(rstn), .Q(
        result_reg4[137]) );
  DFFRHQX1 result_reg4_reg_136_ ( .D(n826), .CK(clk), .RN(rstn), .Q(
        result_reg4[136]) );
  DFFRHQX1 result_reg4_reg_135_ ( .D(n825), .CK(clk), .RN(rstn), .Q(
        result_reg4[135]) );
  DFFRHQX1 result_reg4_reg_134_ ( .D(n824), .CK(clk), .RN(rstn), .Q(
        result_reg4[134]) );
  DFFRHQX1 result_reg4_reg_133_ ( .D(n823), .CK(clk), .RN(rstn), .Q(
        result_reg4[133]) );
  DFFRHQX1 result_reg4_reg_132_ ( .D(n822), .CK(clk), .RN(rstn), .Q(
        result_reg4[132]) );
  DFFRHQX1 result_reg4_reg_131_ ( .D(n821), .CK(clk), .RN(rstn), .Q(
        result_reg4[131]) );
  DFFRHQX1 result_reg4_reg_130_ ( .D(n820), .CK(clk), .RN(rstn), .Q(
        result_reg4[130]) );
  DFFRHQX1 result_reg4_reg_129_ ( .D(n819), .CK(clk), .RN(rstn), .Q(
        result_reg4[129]) );
  DFFRHQX1 result_reg4_reg_128_ ( .D(n818), .CK(clk), .RN(rstn), .Q(
        result_reg4[128]) );
  DFFRHQX1 result_reg4_reg_127_ ( .D(n817), .CK(clk), .RN(rstn), .Q(
        result_reg4[127]) );
  DFFRHQX1 result_reg4_reg_126_ ( .D(n816), .CK(clk), .RN(rstn), .Q(
        result_reg4[126]) );
  DFFRHQX1 result_reg4_reg_125_ ( .D(n815), .CK(clk), .RN(rstn), .Q(
        result_reg4[125]) );
  DFFRHQX1 result_reg4_reg_124_ ( .D(n814), .CK(clk), .RN(rstn), .Q(
        result_reg4[124]) );
  DFFRHQX1 result_reg4_reg_123_ ( .D(n813), .CK(clk), .RN(rstn), .Q(
        result_reg4[123]) );
  DFFRHQX1 result_reg4_reg_122_ ( .D(n812), .CK(clk), .RN(rstn), .Q(
        result_reg4[122]) );
  DFFRHQX1 result_reg4_reg_121_ ( .D(n811), .CK(clk), .RN(rstn), .Q(
        result_reg4[121]) );
  DFFRHQX1 result_reg4_reg_120_ ( .D(n810), .CK(clk), .RN(rstn), .Q(
        result_reg4[120]) );
  DFFRHQX1 result_reg4_reg_119_ ( .D(n809), .CK(clk), .RN(rstn), .Q(
        result_reg4[119]) );
  DFFRHQX1 result_reg4_reg_118_ ( .D(n808), .CK(clk), .RN(rstn), .Q(
        result_reg4[118]) );
  DFFRHQX1 result_reg4_reg_117_ ( .D(n807), .CK(clk), .RN(rstn), .Q(
        result_reg4[117]) );
  DFFRHQX1 result_reg4_reg_116_ ( .D(n806), .CK(clk), .RN(rstn), .Q(
        result_reg4[116]) );
  DFFRHQX1 result_reg4_reg_115_ ( .D(n805), .CK(clk), .RN(rstn), .Q(
        result_reg4[115]) );
  DFFRHQX1 result_reg4_reg_114_ ( .D(n804), .CK(clk), .RN(rstn), .Q(
        result_reg4[114]) );
  DFFRHQX1 result_reg4_reg_113_ ( .D(n803), .CK(clk), .RN(rstn), .Q(
        result_reg4[113]) );
  DFFRHQX1 result_reg4_reg_112_ ( .D(n802), .CK(clk), .RN(rstn), .Q(
        result_reg4[112]) );
  DFFRHQX1 result_reg4_reg_111_ ( .D(n801), .CK(clk), .RN(rstn), .Q(
        result_reg4[111]) );
  DFFRHQX1 result_reg4_reg_110_ ( .D(n800), .CK(clk), .RN(rstn), .Q(
        result_reg4[110]) );
  DFFRHQX1 result_reg4_reg_109_ ( .D(n799), .CK(clk), .RN(rstn), .Q(
        result_reg4[109]) );
  DFFRHQX1 result_reg4_reg_108_ ( .D(n798), .CK(clk), .RN(rstn), .Q(
        result_reg4[108]) );
  DFFRHQX1 result_reg4_reg_107_ ( .D(n797), .CK(clk), .RN(rstn), .Q(
        result_reg4[107]) );
  DFFRHQX1 result_reg4_reg_106_ ( .D(n796), .CK(clk), .RN(rstn), .Q(
        result_reg4[106]) );
  DFFRHQX1 result_reg4_reg_105_ ( .D(n795), .CK(clk), .RN(rstn), .Q(
        result_reg4[105]) );
  DFFRHQX1 result_reg4_reg_104_ ( .D(n794), .CK(clk), .RN(rstn), .Q(
        result_reg4[104]) );
  DFFRHQX1 result_reg4_reg_103_ ( .D(n793), .CK(clk), .RN(rstn), .Q(
        result_reg4[103]) );
  DFFRHQX1 result_reg4_reg_102_ ( .D(n792), .CK(clk), .RN(rstn), .Q(
        result_reg4[102]) );
  DFFRHQX1 result_reg4_reg_101_ ( .D(n791), .CK(clk), .RN(rstn), .Q(
        result_reg4[101]) );
  DFFRHQX1 result_reg4_reg_100_ ( .D(n790), .CK(clk), .RN(rstn), .Q(
        result_reg4[100]) );
  DFFRHQX1 result_reg4_reg_99_ ( .D(n789), .CK(clk), .RN(rstn), .Q(
        result_reg4[99]) );
  DFFRHQX1 result_reg4_reg_98_ ( .D(n788), .CK(clk), .RN(rstn), .Q(
        result_reg4[98]) );
  DFFRHQX1 result_reg4_reg_97_ ( .D(n787), .CK(clk), .RN(rstn), .Q(
        result_reg4[97]) );
  DFFRHQX1 result_reg4_reg_96_ ( .D(n786), .CK(clk), .RN(rstn), .Q(
        result_reg4[96]) );
  DFFRHQX1 result_reg4_reg_15_ ( .D(n1141), .CK(clk), .RN(rstn), .Q(
        result_reg4[15]) );
  DFFRHQX1 result_reg4_reg_14_ ( .D(n1140), .CK(clk), .RN(rstn), .Q(
        result_reg4[14]) );
  DFFRHQX1 result_reg4_reg_13_ ( .D(n1139), .CK(clk), .RN(rstn), .Q(
        result_reg4[13]) );
  DFFRHQX1 result_reg4_reg_12_ ( .D(n1138), .CK(clk), .RN(rstn), .Q(
        result_reg4[12]) );
  DFFRHQX1 result_reg4_reg_11_ ( .D(n1137), .CK(clk), .RN(rstn), .Q(
        result_reg4[11]) );
  DFFRHQX1 result_reg4_reg_10_ ( .D(n1136), .CK(clk), .RN(rstn), .Q(
        result_reg4[10]) );
  DFFRHQX1 result_reg4_reg_9_ ( .D(n1135), .CK(clk), .RN(rstn), .Q(
        result_reg4[9]) );
  DFFRHQX1 result_reg4_reg_8_ ( .D(n1134), .CK(clk), .RN(rstn), .Q(
        result_reg4[8]) );
  DFFRHQX1 result_reg4_reg_7_ ( .D(n1133), .CK(clk), .RN(rstn), .Q(
        result_reg4[7]) );
  DFFRHQX1 result_reg4_reg_6_ ( .D(n1132), .CK(clk), .RN(rstn), .Q(
        result_reg4[6]) );
  DFFRHQX1 result_reg4_reg_5_ ( .D(n1131), .CK(clk), .RN(rstn), .Q(
        result_reg4[5]) );
  DFFRHQX1 result_reg4_reg_4_ ( .D(n1130), .CK(clk), .RN(rstn), .Q(
        result_reg4[4]) );
  DFFRHQX1 result_reg4_reg_3_ ( .D(n1129), .CK(clk), .RN(rstn), .Q(
        result_reg4[3]) );
  DFFRHQX1 result_reg4_reg_2_ ( .D(n1128), .CK(clk), .RN(rstn), .Q(
        result_reg4[2]) );
  DFFRHQX1 result_reg4_reg_1_ ( .D(n1127), .CK(clk), .RN(rstn), .Q(
        result_reg4[1]) );
  DFFRHQX1 result_reg4_reg_0_ ( .D(n1126), .CK(clk), .RN(rstn), .Q(
        result_reg4[0]) );
  DFFRHQX1 result_reg4_reg_63_ ( .D(n1189), .CK(clk), .RN(rstn), .Q(
        result_reg4[63]) );
  DFFRHQX1 result_reg4_reg_47_ ( .D(n1173), .CK(clk), .RN(rstn), .Q(
        result_reg4[47]) );
  DFFRHQX1 result_reg4_reg_31_ ( .D(n1157), .CK(clk), .RN(rstn), .Q(
        result_reg4[31]) );
  DFFRHQX1 result_reg4_reg_62_ ( .D(n1188), .CK(clk), .RN(rstn), .Q(
        result_reg4[62]) );
  DFFRHQX1 result_reg4_reg_46_ ( .D(n1172), .CK(clk), .RN(rstn), .Q(
        result_reg4[46]) );
  DFFRHQX1 result_reg4_reg_30_ ( .D(n1156), .CK(clk), .RN(rstn), .Q(
        result_reg4[30]) );
  DFFRHQX1 result_reg4_reg_61_ ( .D(n1187), .CK(clk), .RN(rstn), .Q(
        result_reg4[61]) );
  DFFRHQX1 result_reg4_reg_45_ ( .D(n1171), .CK(clk), .RN(rstn), .Q(
        result_reg4[45]) );
  DFFRHQX1 result_reg4_reg_29_ ( .D(n1155), .CK(clk), .RN(rstn), .Q(
        result_reg4[29]) );
  DFFRHQX1 result_reg4_reg_60_ ( .D(n1186), .CK(clk), .RN(rstn), .Q(
        result_reg4[60]) );
  DFFRHQX1 result_reg4_reg_44_ ( .D(n1170), .CK(clk), .RN(rstn), .Q(
        result_reg4[44]) );
  DFFRHQX1 result_reg4_reg_28_ ( .D(n1154), .CK(clk), .RN(rstn), .Q(
        result_reg4[28]) );
  DFFRHQX1 result_reg4_reg_59_ ( .D(n1185), .CK(clk), .RN(rstn), .Q(
        result_reg4[59]) );
  DFFRHQX1 result_reg4_reg_43_ ( .D(n1169), .CK(clk), .RN(rstn), .Q(
        result_reg4[43]) );
  DFFRHQX1 result_reg4_reg_27_ ( .D(n1153), .CK(clk), .RN(rstn), .Q(
        result_reg4[27]) );
  DFFRHQX1 result_reg4_reg_58_ ( .D(n1184), .CK(clk), .RN(rstn), .Q(
        result_reg4[58]) );
  DFFRHQX1 result_reg4_reg_42_ ( .D(n1168), .CK(clk), .RN(rstn), .Q(
        result_reg4[42]) );
  DFFRHQX1 result_reg4_reg_26_ ( .D(n1152), .CK(clk), .RN(rstn), .Q(
        result_reg4[26]) );
  DFFRHQX1 result_reg4_reg_57_ ( .D(n1183), .CK(clk), .RN(rstn), .Q(
        result_reg4[57]) );
  DFFRHQX1 result_reg4_reg_41_ ( .D(n1167), .CK(clk), .RN(rstn), .Q(
        result_reg4[41]) );
  DFFRHQX1 result_reg4_reg_25_ ( .D(n1151), .CK(clk), .RN(rstn), .Q(
        result_reg4[25]) );
  DFFRHQX1 result_reg4_reg_56_ ( .D(n1182), .CK(clk), .RN(rstn), .Q(
        result_reg4[56]) );
  DFFRHQX1 result_reg4_reg_40_ ( .D(n1166), .CK(clk), .RN(rstn), .Q(
        result_reg4[40]) );
  DFFRHQX1 result_reg4_reg_24_ ( .D(n1150), .CK(clk), .RN(rstn), .Q(
        result_reg4[24]) );
  DFFRHQX1 result_reg4_reg_55_ ( .D(n1181), .CK(clk), .RN(rstn), .Q(
        result_reg4[55]) );
  DFFRHQX1 result_reg4_reg_39_ ( .D(n1165), .CK(clk), .RN(rstn), .Q(
        result_reg4[39]) );
  DFFRHQX1 result_reg4_reg_23_ ( .D(n1149), .CK(clk), .RN(rstn), .Q(
        result_reg4[23]) );
  DFFRHQX1 result_reg4_reg_54_ ( .D(n1180), .CK(clk), .RN(rstn), .Q(
        result_reg4[54]) );
  DFFRHQX1 result_reg4_reg_38_ ( .D(n1164), .CK(clk), .RN(rstn), .Q(
        result_reg4[38]) );
  DFFRHQX1 result_reg4_reg_22_ ( .D(n1148), .CK(clk), .RN(rstn), .Q(
        result_reg4[22]) );
  DFFRHQX1 result_reg4_reg_53_ ( .D(n1179), .CK(clk), .RN(rstn), .Q(
        result_reg4[53]) );
  DFFRHQX1 result_reg4_reg_37_ ( .D(n1163), .CK(clk), .RN(rstn), .Q(
        result_reg4[37]) );
  DFFRHQX1 result_reg4_reg_21_ ( .D(n1147), .CK(clk), .RN(rstn), .Q(
        result_reg4[21]) );
  DFFRHQX1 result_reg4_reg_52_ ( .D(n1178), .CK(clk), .RN(rstn), .Q(
        result_reg4[52]) );
  DFFRHQX1 result_reg4_reg_36_ ( .D(n1162), .CK(clk), .RN(rstn), .Q(
        result_reg4[36]) );
  DFFRHQX1 result_reg4_reg_20_ ( .D(n1146), .CK(clk), .RN(rstn), .Q(
        result_reg4[20]) );
  DFFRHQX1 result_reg4_reg_51_ ( .D(n1177), .CK(clk), .RN(rstn), .Q(
        result_reg4[51]) );
  DFFRHQX1 result_reg4_reg_35_ ( .D(n1161), .CK(clk), .RN(rstn), .Q(
        result_reg4[35]) );
  DFFRHQX1 result_reg4_reg_19_ ( .D(n1145), .CK(clk), .RN(rstn), .Q(
        result_reg4[19]) );
  DFFRHQX1 result_reg4_reg_50_ ( .D(n1176), .CK(clk), .RN(rstn), .Q(
        result_reg4[50]) );
  DFFRHQX1 result_reg4_reg_34_ ( .D(n1160), .CK(clk), .RN(rstn), .Q(
        result_reg4[34]) );
  DFFRHQX1 result_reg4_reg_18_ ( .D(n1144), .CK(clk), .RN(rstn), .Q(
        result_reg4[18]) );
  DFFRHQX1 result_reg4_reg_49_ ( .D(n1175), .CK(clk), .RN(rstn), .Q(
        result_reg4[49]) );
  DFFRHQX1 result_reg4_reg_33_ ( .D(n1159), .CK(clk), .RN(rstn), .Q(
        result_reg4[33]) );
  DFFRHQX1 result_reg4_reg_17_ ( .D(n1143), .CK(clk), .RN(rstn), .Q(
        result_reg4[17]) );
  DFFRHQX1 result_reg4_reg_48_ ( .D(n1174), .CK(clk), .RN(rstn), .Q(
        result_reg4[48]) );
  DFFRHQX1 result_reg4_reg_32_ ( .D(n1158), .CK(clk), .RN(rstn), .Q(
        result_reg4[32]) );
  DFFRHQX1 result_reg4_reg_16_ ( .D(n1142), .CK(clk), .RN(rstn), .Q(
        result_reg4[16]) );
  DFFRHQX1 result_reg8_reg_127_ ( .D(n1269), .CK(clk), .RN(rstn), .Q(
        result_reg8[127]) );
  DFFRHQX1 result_reg8_reg_126_ ( .D(n1268), .CK(clk), .RN(rstn), .Q(
        result_reg8[126]) );
  DFFRHQX1 result_reg8_reg_125_ ( .D(n1267), .CK(clk), .RN(rstn), .Q(
        result_reg8[125]) );
  DFFRHQX1 result_reg8_reg_124_ ( .D(n1266), .CK(clk), .RN(rstn), .Q(
        result_reg8[124]) );
  DFFRHQX1 result_reg8_reg_123_ ( .D(n1265), .CK(clk), .RN(rstn), .Q(
        result_reg8[123]) );
  DFFRHQX1 result_reg8_reg_122_ ( .D(n1264), .CK(clk), .RN(rstn), .Q(
        result_reg8[122]) );
  DFFRHQX1 result_reg8_reg_121_ ( .D(n1263), .CK(clk), .RN(rstn), .Q(
        result_reg8[121]) );
  DFFRHQX1 result_reg8_reg_120_ ( .D(n1262), .CK(clk), .RN(rstn), .Q(
        result_reg8[120]) );
  DFFRHQX1 result_reg8_reg_119_ ( .D(n1261), .CK(clk), .RN(rstn), .Q(
        result_reg8[119]) );
  DFFRHQX1 result_reg8_reg_118_ ( .D(n1260), .CK(clk), .RN(rstn), .Q(
        result_reg8[118]) );
  DFFRHQX1 result_reg8_reg_117_ ( .D(n1259), .CK(clk), .RN(rstn), .Q(
        result_reg8[117]) );
  DFFRHQX1 result_reg8_reg_116_ ( .D(n1258), .CK(clk), .RN(rstn), .Q(
        result_reg8[116]) );
  DFFRHQX1 result_reg8_reg_115_ ( .D(n1257), .CK(clk), .RN(rstn), .Q(
        result_reg8[115]) );
  DFFRHQX1 result_reg8_reg_114_ ( .D(n1256), .CK(clk), .RN(rstn), .Q(
        result_reg8[114]) );
  DFFRHQX1 result_reg8_reg_113_ ( .D(n1255), .CK(clk), .RN(rstn), .Q(
        result_reg8[113]) );
  DFFRHQX1 result_reg8_reg_112_ ( .D(n1254), .CK(clk), .RN(rstn), .Q(
        result_reg8[112]) );
  DFFRHQX1 mode_reg_reg_0_ ( .D(n882), .CK(clk), .RN(rstn), .Q(mode_reg_0_) );
  DFFRHQX1 dout_reg_15_ ( .D(n883), .CK(clk), .RN(rstn), .Q(dout[15]) );
  DFFRHQX1 dout_reg_14_ ( .D(n884), .CK(clk), .RN(rstn), .Q(dout[14]) );
  DFFRHQX1 dout_reg_13_ ( .D(n885), .CK(clk), .RN(rstn), .Q(dout[13]) );
  DFFRHQX1 dout_reg_12_ ( .D(n886), .CK(clk), .RN(rstn), .Q(dout[12]) );
  DFFRHQX1 dout_reg_11_ ( .D(n887), .CK(clk), .RN(rstn), .Q(dout[11]) );
  DFFRHQX1 dout_reg_10_ ( .D(n888), .CK(clk), .RN(rstn), .Q(dout[10]) );
  DFFRHQX1 dout_reg_9_ ( .D(n889), .CK(clk), .RN(rstn), .Q(dout[9]) );
  DFFRHQX1 dout_reg_8_ ( .D(n890), .CK(clk), .RN(rstn), .Q(dout[8]) );
  DFFRHQX1 dout_reg_7_ ( .D(n891), .CK(clk), .RN(rstn), .Q(dout[7]) );
  DFFRHQX1 dout_reg_6_ ( .D(n892), .CK(clk), .RN(rstn), .Q(dout[6]) );
  DFFRHQX1 dout_reg_5_ ( .D(n893), .CK(clk), .RN(rstn), .Q(dout[5]) );
  DFFRHQX1 dout_reg_4_ ( .D(n894), .CK(clk), .RN(rstn), .Q(dout[4]) );
  DFFRHQX1 dout_reg_3_ ( .D(n895), .CK(clk), .RN(rstn), .Q(dout[3]) );
  DFFRHQX1 dout_reg_2_ ( .D(n896), .CK(clk), .RN(rstn), .Q(dout[2]) );
  DFFRHQX1 dout_reg_1_ ( .D(n897), .CK(clk), .RN(rstn), .Q(dout[1]) );
  DFFRHQX1 dout_reg_0_ ( .D(n898), .CK(clk), .RN(rstn), .Q(dout[0]) );
  DFFRHQX1 shift4_flag_reg ( .D(n753), .CK(clk), .RN(rstn), .Q(shift4_flag) );
  DFFRHQX1 start_reg4_reg_0_ ( .D(n752), .CK(clk), .RN(rstn), .Q(start_reg4[0]) );
  DFFRHQX1 ready8_reg ( .D(n746), .CK(clk), .RN(rstn), .Q(ready8) );
  OR3XL U3 ( .A(n1124), .B(n225), .C(n745), .Y(n81) );
  AND2X2 U6 ( .A(n1102), .B(n225), .Y(n82) );
  AND2X2 U7 ( .A(start), .B(n97), .Y(n83) );
  INVX1 U8 ( .A(n133), .Y(n92) );
  INVX1 U9 ( .A(n133), .Y(n93) );
  INVX1 U10 ( .A(n134), .Y(n94) );
  INVX1 U11 ( .A(n134), .Y(n95) );
  INVX1 U12 ( .A(n134), .Y(n96) );
  INVX1 U13 ( .A(n135), .Y(n98) );
  INVX1 U14 ( .A(n134), .Y(n97) );
  INVX1 U15 ( .A(n133), .Y(n91) );
  INVX1 U16 ( .A(n133), .Y(n99) );
  INVX1 U17 ( .A(n138), .Y(n134) );
  INVX1 U18 ( .A(n138), .Y(n133) );
  INVX1 U19 ( .A(n138), .Y(n135) );
  INVX1 U20 ( .A(n139), .Y(n112) );
  INVX1 U21 ( .A(n144), .Y(n108) );
  INVX1 U22 ( .A(n144), .Y(n110) );
  INVX1 U23 ( .A(n144), .Y(n109) );
  INVX1 U24 ( .A(n139), .Y(n111) );
  INVX1 U25 ( .A(n141), .Y(n122) );
  INVX1 U26 ( .A(n139), .Y(n129) );
  INVX1 U27 ( .A(n139), .Y(n130) );
  INVX1 U28 ( .A(n141), .Y(n123) );
  INVX1 U29 ( .A(n139), .Y(n131) );
  INVX1 U30 ( .A(n140), .Y(n125) );
  INVX1 U31 ( .A(n139), .Y(n132) );
  INVX1 U32 ( .A(n141), .Y(n124) );
  INVX1 U33 ( .A(n139), .Y(n128) );
  INVX1 U34 ( .A(n140), .Y(n127) );
  INVX1 U35 ( .A(n140), .Y(n126) );
  INVX1 U36 ( .A(n141), .Y(n120) );
  INVX1 U37 ( .A(n143), .Y(n116) );
  INVX1 U38 ( .A(n142), .Y(n113) );
  INVX1 U39 ( .A(n140), .Y(n121) );
  INVX1 U40 ( .A(n143), .Y(n115) );
  INVX1 U41 ( .A(n142), .Y(n117) );
  INVX1 U42 ( .A(n142), .Y(n118) );
  INVX1 U43 ( .A(n143), .Y(n114) );
  INVX1 U44 ( .A(n142), .Y(n119) );
  INVX1 U45 ( .A(n144), .Y(n107) );
  INVX1 U46 ( .A(n210), .Y(n103) );
  INVX1 U47 ( .A(n210), .Y(n101) );
  INVX1 U48 ( .A(n210), .Y(n102) );
  INVX1 U49 ( .A(n209), .Y(n105) );
  INVX1 U50 ( .A(n209), .Y(n106) );
  INVX1 U51 ( .A(n209), .Y(n104) );
  INVX1 U52 ( .A(n83), .Y(n89) );
  INVX1 U53 ( .A(n83), .Y(n90) );
  INVX1 U54 ( .A(n211), .Y(n136) );
  INVX1 U55 ( .A(n211), .Y(n137) );
  INVX1 U56 ( .A(n214), .Y(n138) );
  INVX1 U57 ( .A(n214), .Y(n139) );
  INVX1 U58 ( .A(n213), .Y(n141) );
  INVX1 U59 ( .A(n212), .Y(n140) );
  INVX1 U60 ( .A(n212), .Y(n144) );
  INVX1 U61 ( .A(n213), .Y(n142) );
  INVX1 U62 ( .A(n213), .Y(n143) );
  INVX1 U63 ( .A(n211), .Y(n100) );
  INVX1 U64 ( .A(n212), .Y(n211) );
  INVX1 U65 ( .A(n212), .Y(n210) );
  INVX1 U66 ( .A(n212), .Y(n209) );
  INVX1 U67 ( .A(n229), .Y(n225) );
  INVX1 U68 ( .A(n81), .Y(n223) );
  INVX1 U69 ( .A(n81), .Y(n224) );
  INVX1 U70 ( .A(n219), .Y(n217) );
  INVX1 U71 ( .A(n219), .Y(n218) );
  INVX1 U72 ( .A(n966), .Y(n214) );
  INVX1 U73 ( .A(n966), .Y(n213) );
  INVX1 U74 ( .A(n219), .Y(n216) );
  INVX1 U75 ( .A(n81), .Y(n222) );
  INVX1 U76 ( .A(n81), .Y(n220) );
  INVX1 U77 ( .A(n229), .Y(n226) );
  INVX1 U78 ( .A(n229), .Y(n227) );
  INVX1 U79 ( .A(n229), .Y(n228) );
  INVX1 U80 ( .A(n966), .Y(n212) );
  NAND2X1 U81 ( .A(n901), .B(n87), .Y(n966) );
  INVX1 U82 ( .A(start), .Y(n745) );
  INVX1 U83 ( .A(n84), .Y(n87) );
  INVX1 U84 ( .A(n1081), .Y(n219) );
  INVX1 U85 ( .A(n900), .Y(n1125) );
  INVX1 U86 ( .A(n84), .Y(n88) );
  INVX1 U87 ( .A(n1100), .Y(n229) );
  OAI222XL U88 ( .A0(n232), .A1(n89), .B0(n87), .B1(n712), .C0(n98), .C1(n728), 
        .Y(n784) );
  INVX1 U89 ( .A(cal_result[15]), .Y(n232) );
  OAI222XL U90 ( .A0(n248), .A1(n90), .B0(n88), .B1(n696), .C0(n97), .C1(n712), 
        .Y(n801) );
  INVX1 U91 ( .A(cal_result[31]), .Y(n248) );
  OAI222XL U92 ( .A0(n264), .A1(n89), .B0(n88), .B1(n680), .C0(n98), .C1(n696), 
        .Y(n817) );
  INVX1 U93 ( .A(cal_result[47]), .Y(n264) );
  OAI22X1 U94 ( .A0(n91), .A1(n680), .B0(n280), .B1(n90), .Y(n833) );
  INVX1 U95 ( .A(cal_result[63]), .Y(n280) );
  OAI222XL U96 ( .A0(n245), .A1(n90), .B0(n87), .B1(n727), .C0(n99), .C1(n743), 
        .Y(n754) );
  INVX1 U97 ( .A(cal_result[0]), .Y(n245) );
  OAI222XL U98 ( .A0(n244), .A1(n90), .B0(n87), .B1(n726), .C0(n99), .C1(n742), 
        .Y(n756) );
  INVX1 U99 ( .A(cal_result[1]), .Y(n244) );
  OAI222XL U100 ( .A0(n243), .A1(n90), .B0(n87), .B1(n725), .C0(n99), .C1(n741), .Y(n758) );
  INVX1 U101 ( .A(cal_result[2]), .Y(n243) );
  OAI222XL U102 ( .A0(n242), .A1(n90), .B0(n87), .B1(n724), .C0(n99), .C1(n740), .Y(n760) );
  INVX1 U103 ( .A(cal_result[3]), .Y(n242) );
  OAI222XL U104 ( .A0(n241), .A1(n90), .B0(n87), .B1(n723), .C0(n99), .C1(n739), .Y(n762) );
  INVX1 U105 ( .A(cal_result[4]), .Y(n241) );
  OAI222XL U106 ( .A0(n240), .A1(n90), .B0(n87), .B1(n722), .C0(n99), .C1(n738), .Y(n764) );
  INVX1 U107 ( .A(cal_result[5]), .Y(n240) );
  OAI222XL U108 ( .A0(n239), .A1(n90), .B0(n87), .B1(n721), .C0(n99), .C1(n737), .Y(n766) );
  INVX1 U109 ( .A(cal_result[6]), .Y(n239) );
  OAI222XL U110 ( .A0(n238), .A1(n90), .B0(n87), .B1(n720), .C0(n99), .C1(n736), .Y(n768) );
  INVX1 U111 ( .A(cal_result[7]), .Y(n238) );
  OAI222XL U112 ( .A0(n237), .A1(n90), .B0(n87), .B1(n719), .C0(n99), .C1(n735), .Y(n770) );
  INVX1 U113 ( .A(cal_result[8]), .Y(n237) );
  OAI222XL U114 ( .A0(n236), .A1(n89), .B0(n87), .B1(n718), .C0(n98), .C1(n734), .Y(n772) );
  INVX1 U115 ( .A(cal_result[9]), .Y(n236) );
  OAI222XL U116 ( .A0(n235), .A1(n89), .B0(n87), .B1(n717), .C0(n98), .C1(n733), .Y(n774) );
  INVX1 U117 ( .A(cal_result[10]), .Y(n235) );
  OAI222XL U118 ( .A0(n234), .A1(n89), .B0(n87), .B1(n716), .C0(n98), .C1(n732), .Y(n776) );
  INVX1 U119 ( .A(cal_result[11]), .Y(n234) );
  OAI222XL U120 ( .A0(n233), .A1(n89), .B0(n87), .B1(n715), .C0(n98), .C1(n731), .Y(n778) );
  INVX1 U121 ( .A(cal_result[12]), .Y(n233) );
  OAI222XL U122 ( .A0(n230), .A1(n89), .B0(n87), .B1(n714), .C0(n98), .C1(n730), .Y(n780) );
  INVX1 U123 ( .A(cal_result[13]), .Y(n230) );
  OAI222XL U124 ( .A0(n231), .A1(n89), .B0(n87), .B1(n713), .C0(n98), .C1(n729), .Y(n782) );
  INVX1 U125 ( .A(cal_result[14]), .Y(n231) );
  OAI222XL U126 ( .A0(n261), .A1(n89), .B0(n87), .B1(n711), .C0(n97), .C1(n727), .Y(n786) );
  INVX1 U127 ( .A(cal_result[16]), .Y(n261) );
  OAI222XL U128 ( .A0(n260), .A1(n89), .B0(n87), .B1(n710), .C0(n97), .C1(n726), .Y(n787) );
  INVX1 U129 ( .A(cal_result[17]), .Y(n260) );
  OAI222XL U130 ( .A0(n259), .A1(n89), .B0(n88), .B1(n709), .C0(n97), .C1(n725), .Y(n788) );
  INVX1 U131 ( .A(cal_result[18]), .Y(n259) );
  OAI222XL U132 ( .A0(n258), .A1(n89), .B0(n88), .B1(n708), .C0(n97), .C1(n724), .Y(n789) );
  INVX1 U133 ( .A(cal_result[19]), .Y(n258) );
  OAI222XL U134 ( .A0(n257), .A1(n89), .B0(n88), .B1(n707), .C0(n97), .C1(n723), .Y(n790) );
  INVX1 U135 ( .A(cal_result[20]), .Y(n257) );
  OAI222XL U136 ( .A0(n256), .A1(n89), .B0(n88), .B1(n706), .C0(n97), .C1(n722), .Y(n791) );
  INVX1 U137 ( .A(cal_result[21]), .Y(n256) );
  OAI222XL U138 ( .A0(n255), .A1(n89), .B0(n88), .B1(n705), .C0(n97), .C1(n721), .Y(n792) );
  INVX1 U139 ( .A(cal_result[22]), .Y(n255) );
  OAI222XL U140 ( .A0(n254), .A1(n89), .B0(n88), .B1(n704), .C0(n97), .C1(n720), .Y(n793) );
  INVX1 U141 ( .A(cal_result[23]), .Y(n254) );
  OAI222XL U142 ( .A0(n253), .A1(n89), .B0(n88), .B1(n703), .C0(n97), .C1(n719), .Y(n794) );
  INVX1 U143 ( .A(cal_result[24]), .Y(n253) );
  OAI222XL U144 ( .A0(n252), .A1(n89), .B0(n88), .B1(n702), .C0(n97), .C1(n718), .Y(n795) );
  INVX1 U145 ( .A(cal_result[25]), .Y(n252) );
  OAI222XL U146 ( .A0(n251), .A1(n89), .B0(n88), .B1(n701), .C0(n97), .C1(n717), .Y(n796) );
  INVX1 U147 ( .A(cal_result[26]), .Y(n251) );
  OAI222XL U148 ( .A0(n250), .A1(n89), .B0(n88), .B1(n700), .C0(n97), .C1(n716), .Y(n797) );
  INVX1 U149 ( .A(cal_result[27]), .Y(n250) );
  OAI222XL U150 ( .A0(n249), .A1(n89), .B0(n88), .B1(n699), .C0(n97), .C1(n715), .Y(n798) );
  INVX1 U151 ( .A(cal_result[28]), .Y(n249) );
  OAI222XL U152 ( .A0(n246), .A1(n89), .B0(n88), .B1(n698), .C0(n97), .C1(n714), .Y(n799) );
  INVX1 U153 ( .A(cal_result[29]), .Y(n246) );
  OAI222XL U154 ( .A0(n247), .A1(n89), .B0(n88), .B1(n697), .C0(n97), .C1(n713), .Y(n800) );
  INVX1 U155 ( .A(cal_result[30]), .Y(n247) );
  OAI222XL U156 ( .A0(n277), .A1(n89), .B0(n88), .B1(n695), .C0(n98), .C1(n711), .Y(n802) );
  INVX1 U157 ( .A(cal_result[32]), .Y(n277) );
  OAI222XL U158 ( .A0(n276), .A1(n90), .B0(n88), .B1(n694), .C0(n98), .C1(n710), .Y(n803) );
  INVX1 U159 ( .A(cal_result[33]), .Y(n276) );
  OAI222XL U160 ( .A0(n275), .A1(n89), .B0(n88), .B1(n693), .C0(n98), .C1(n709), .Y(n804) );
  INVX1 U161 ( .A(cal_result[34]), .Y(n275) );
  OAI222XL U162 ( .A0(n274), .A1(n90), .B0(n88), .B1(n692), .C0(n98), .C1(n708), .Y(n805) );
  INVX1 U163 ( .A(cal_result[35]), .Y(n274) );
  OAI222XL U164 ( .A0(n273), .A1(n89), .B0(n88), .B1(n691), .C0(n98), .C1(n707), .Y(n806) );
  INVX1 U165 ( .A(cal_result[36]), .Y(n273) );
  OAI222XL U166 ( .A0(n272), .A1(n90), .B0(n88), .B1(n690), .C0(n98), .C1(n706), .Y(n807) );
  INVX1 U167 ( .A(cal_result[37]), .Y(n272) );
  OAI222XL U168 ( .A0(n271), .A1(n89), .B0(n88), .B1(n689), .C0(n98), .C1(n705), .Y(n808) );
  INVX1 U169 ( .A(cal_result[38]), .Y(n271) );
  OAI222XL U170 ( .A0(n270), .A1(n90), .B0(n88), .B1(n688), .C0(n98), .C1(n704), .Y(n809) );
  INVX1 U171 ( .A(cal_result[39]), .Y(n270) );
  OAI222XL U172 ( .A0(n269), .A1(n89), .B0(n88), .B1(n687), .C0(n98), .C1(n703), .Y(n810) );
  INVX1 U173 ( .A(cal_result[40]), .Y(n269) );
  OAI222XL U174 ( .A0(n268), .A1(n90), .B0(n88), .B1(n686), .C0(n98), .C1(n702), .Y(n811) );
  INVX1 U175 ( .A(cal_result[41]), .Y(n268) );
  OAI222XL U176 ( .A0(n267), .A1(n89), .B0(n88), .B1(n685), .C0(n98), .C1(n701), .Y(n812) );
  INVX1 U177 ( .A(cal_result[42]), .Y(n267) );
  OAI222XL U178 ( .A0(n266), .A1(n90), .B0(n88), .B1(n684), .C0(n98), .C1(n700), .Y(n813) );
  INVX1 U179 ( .A(cal_result[43]), .Y(n266) );
  OAI222XL U180 ( .A0(n265), .A1(n89), .B0(n88), .B1(n683), .C0(n98), .C1(n699), .Y(n814) );
  INVX1 U181 ( .A(cal_result[44]), .Y(n265) );
  OAI222XL U182 ( .A0(n262), .A1(n90), .B0(n88), .B1(n682), .C0(n98), .C1(n698), .Y(n815) );
  INVX1 U183 ( .A(cal_result[45]), .Y(n262) );
  OAI222XL U184 ( .A0(n263), .A1(n89), .B0(n88), .B1(n681), .C0(n98), .C1(n697), .Y(n816) );
  INVX1 U185 ( .A(cal_result[46]), .Y(n263) );
  OAI22X1 U186 ( .A0(n91), .A1(n695), .B0(n671), .B1(n90), .Y(n818) );
  INVX1 U187 ( .A(cal_result[48]), .Y(n671) );
  OAI22X1 U188 ( .A0(n92), .A1(n694), .B0(n670), .B1(n90), .Y(n819) );
  INVX1 U189 ( .A(cal_result[49]), .Y(n670) );
  OAI22X1 U190 ( .A0(n91), .A1(n693), .B0(n669), .B1(n90), .Y(n820) );
  INVX1 U191 ( .A(cal_result[50]), .Y(n669) );
  OAI22X1 U192 ( .A0(n92), .A1(n692), .B0(n448), .B1(n90), .Y(n821) );
  INVX1 U193 ( .A(cal_result[51]), .Y(n448) );
  OAI22X1 U194 ( .A0(n91), .A1(n691), .B0(n447), .B1(n90), .Y(n822) );
  INVX1 U195 ( .A(cal_result[52]), .Y(n447) );
  OAI22X1 U196 ( .A0(n92), .A1(n690), .B0(n314), .B1(n90), .Y(n823) );
  INVX1 U197 ( .A(cal_result[53]), .Y(n314) );
  OAI22X1 U198 ( .A0(n91), .A1(n689), .B0(n307), .B1(n90), .Y(n824) );
  INVX1 U199 ( .A(cal_result[54]), .Y(n307) );
  OAI22X1 U200 ( .A0(n92), .A1(n688), .B0(n287), .B1(n90), .Y(n825) );
  INVX1 U201 ( .A(cal_result[55]), .Y(n287) );
  OAI22X1 U202 ( .A0(n91), .A1(n687), .B0(n285), .B1(n90), .Y(n826) );
  INVX1 U203 ( .A(cal_result[56]), .Y(n285) );
  OAI22X1 U204 ( .A0(n91), .A1(n686), .B0(n284), .B1(n90), .Y(n827) );
  INVX1 U205 ( .A(cal_result[57]), .Y(n284) );
  OAI22X1 U206 ( .A0(n91), .A1(n685), .B0(n283), .B1(n90), .Y(n828) );
  INVX1 U207 ( .A(cal_result[58]), .Y(n283) );
  OAI22X1 U208 ( .A0(n91), .A1(n684), .B0(n282), .B1(n90), .Y(n829) );
  INVX1 U209 ( .A(cal_result[59]), .Y(n282) );
  OAI22X1 U210 ( .A0(n91), .A1(n683), .B0(n281), .B1(n90), .Y(n830) );
  INVX1 U211 ( .A(cal_result[60]), .Y(n281) );
  OAI22X1 U212 ( .A0(n91), .A1(n682), .B0(n278), .B1(n90), .Y(n831) );
  INVX1 U213 ( .A(cal_result[61]), .Y(n278) );
  OAI22X1 U214 ( .A0(n91), .A1(n681), .B0(n279), .B1(n89), .Y(n832) );
  INVX1 U215 ( .A(cal_result[62]), .Y(n279) );
  NAND2X1 U216 ( .A(n968), .B(n1124), .Y(n901) );
  NOR2X1 U217 ( .A(n969), .B(n968), .Y(n1100) );
  AOI2BB1X1 U218 ( .A0N(n1124), .A1N(n969), .B0(n225), .Y(n1081) );
  NAND2X1 U219 ( .A(n1103), .B(n1101), .Y(n969) );
  NAND3X1 U220 ( .A(n672), .B(n745), .C(n1123), .Y(n967) );
  AND2X2 U221 ( .A(n1099), .B(n967), .Y(n1103) );
  NAND3X1 U222 ( .A(n1101), .B(n1102), .C(n967), .Y(n84) );
  NAND3X1 U223 ( .A(n1101), .B(n1102), .C(n901), .Y(n900) );
  OAI22X1 U224 ( .A0(n1125), .A1(n677), .B0(n900), .B1(n678), .Y(n751) );
  OAI22X1 U225 ( .A0(n1125), .A1(n676), .B0(n900), .B1(n677), .Y(n750) );
  OAI22X1 U226 ( .A0(n1125), .A1(n675), .B0(n900), .B1(n676), .Y(n749) );
  OAI22X1 U227 ( .A0(n1125), .A1(n674), .B0(n900), .B1(n675), .Y(n748) );
  OAI22X1 U228 ( .A0(n1125), .A1(n745), .B0(n900), .B1(n674), .Y(n747) );
  OAI22X1 U229 ( .A0(n1125), .A1(n678), .B0(n679), .B1(n900), .Y(n752) );
  AND2X2 U230 ( .A(n1101), .B(n745), .Y(n1104) );
  OAI21XL U231 ( .A0(n968), .A1(n672), .B0(n901), .Y(n753) );
  INVX1 U232 ( .A(n1123), .Y(p2s_ready) );
  OAI2BB1X1 U233 ( .A0N(n226), .A1N(result_reg8[79]), .B0(n1049), .Y(n849) );
  AOI22X1 U234 ( .A0(result_reg8[95]), .A1(n216), .B0(cal_result[79]), .B1(
        n222), .Y(n1049) );
  OAI2BB1X1 U235 ( .A0N(n225), .A1N(result_reg8[95]), .B0(n1065), .Y(n865) );
  AOI22X1 U236 ( .A0(result_reg8[111]), .A1(n216), .B0(cal_result[95]), .B1(
        n222), .Y(n1065) );
  OAI2BB1X1 U237 ( .A0N(n225), .A1N(result_reg8[111]), .B0(n1082), .Y(n881) );
  AOI22X1 U238 ( .A0(n1081), .A1(result_reg8[127]), .B0(cal_result[111]), .B1(
        n220), .Y(n1082) );
  INVX1 U239 ( .A(n1098), .Y(n1269) );
  AOI22X1 U240 ( .A0(n228), .A1(result_reg8[127]), .B0(cal_result[127]), .B1(
        n222), .Y(n1098) );
  INVX1 U241 ( .A(n983), .Y(n1203) );
  AOI222X1 U242 ( .A0(n224), .A1(cal_result[13]), .B0(n218), .B1(
        result_reg8[29]), .C0(n228), .C1(result_reg8[13]), .Y(n983) );
  INVX1 U243 ( .A(n984), .Y(n1204) );
  AOI222X1 U244 ( .A0(n224), .A1(cal_result[14]), .B0(n218), .B1(
        result_reg8[30]), .C0(n228), .C1(result_reg8[14]), .Y(n984) );
  INVX1 U245 ( .A(n985), .Y(n1205) );
  AOI222X1 U246 ( .A0(n224), .A1(cal_result[15]), .B0(n218), .B1(
        result_reg8[31]), .C0(n228), .C1(result_reg8[15]), .Y(n985) );
  INVX1 U247 ( .A(n999), .Y(n1219) );
  AOI222X1 U248 ( .A0(n224), .A1(cal_result[29]), .B0(n217), .B1(
        result_reg8[45]), .C0(n228), .C1(result_reg8[29]), .Y(n999) );
  INVX1 U249 ( .A(n1000), .Y(n1220) );
  AOI222X1 U250 ( .A0(n224), .A1(cal_result[30]), .B0(n217), .B1(
        result_reg8[46]), .C0(n226), .C1(result_reg8[30]), .Y(n1000) );
  INVX1 U251 ( .A(n1001), .Y(n1221) );
  AOI222X1 U252 ( .A0(n224), .A1(cal_result[31]), .B0(n217), .B1(
        result_reg8[47]), .C0(n227), .C1(result_reg8[31]), .Y(n1001) );
  INVX1 U253 ( .A(n1015), .Y(n1235) );
  AOI222X1 U254 ( .A0(n223), .A1(cal_result[45]), .B0(n217), .B1(
        result_reg8[61]), .C0(n227), .C1(result_reg8[45]), .Y(n1015) );
  INVX1 U255 ( .A(n1016), .Y(n1236) );
  AOI222X1 U256 ( .A0(n223), .A1(cal_result[46]), .B0(n217), .B1(
        result_reg8[62]), .C0(n227), .C1(result_reg8[46]), .Y(n1016) );
  INVX1 U257 ( .A(n1017), .Y(n1237) );
  AOI222X1 U258 ( .A0(n223), .A1(cal_result[47]), .B0(n217), .B1(
        result_reg8[63]), .C0(n227), .C1(result_reg8[47]), .Y(n1017) );
  INVX1 U259 ( .A(n1031), .Y(n1251) );
  AOI222X1 U260 ( .A0(n223), .A1(cal_result[61]), .B0(n218), .B1(
        result_reg8[77]), .C0(n227), .C1(result_reg8[61]), .Y(n1031) );
  INVX1 U261 ( .A(n1032), .Y(n1252) );
  AOI222X1 U262 ( .A0(n223), .A1(cal_result[62]), .B0(n218), .B1(
        result_reg8[78]), .C0(n227), .C1(result_reg8[62]), .Y(n1032) );
  INVX1 U263 ( .A(n1033), .Y(n1253) );
  AOI222X1 U264 ( .A0(n223), .A1(cal_result[63]), .B0(n218), .B1(
        result_reg8[79]), .C0(n226), .C1(result_reg8[63]), .Y(n1033) );
  NOR2X1 U265 ( .A(mode[1]), .B(n745), .Y(n968) );
  NAND3X1 U266 ( .A(n673), .B(n745), .C(start_reg4[0]), .Y(n1102) );
  NAND3X1 U267 ( .A(n1123), .B(n745), .C(shift4_flag), .Y(n1101) );
  INVX1 U268 ( .A(n1096), .Y(n1267) );
  AOI22X1 U269 ( .A0(n228), .A1(result_reg8[125]), .B0(cal_result[125]), .B1(
        n220), .Y(n1096) );
  OAI2BB1X1 U270 ( .A0N(n226), .A1N(result_reg8[75]), .B0(n1045), .Y(n845) );
  AOI22X1 U271 ( .A0(result_reg8[91]), .A1(n216), .B0(cal_result[75]), .B1(
        n220), .Y(n1045) );
  OAI2BB1X1 U272 ( .A0N(n226), .A1N(result_reg8[76]), .B0(n1046), .Y(n846) );
  AOI22X1 U273 ( .A0(result_reg8[92]), .A1(n216), .B0(cal_result[76]), .B1(
        n222), .Y(n1046) );
  OAI2BB1X1 U274 ( .A0N(n226), .A1N(result_reg8[78]), .B0(n1048), .Y(n848) );
  AOI22X1 U275 ( .A0(result_reg8[94]), .A1(n216), .B0(cal_result[78]), .B1(
        n220), .Y(n1048) );
  OAI2BB1X1 U276 ( .A0N(n226), .A1N(result_reg8[91]), .B0(n1061), .Y(n861) );
  AOI22X1 U277 ( .A0(result_reg8[107]), .A1(n216), .B0(cal_result[91]), .B1(
        n220), .Y(n1061) );
  OAI2BB1X1 U278 ( .A0N(n226), .A1N(result_reg8[92]), .B0(n1062), .Y(n862) );
  AOI22X1 U279 ( .A0(result_reg8[108]), .A1(n216), .B0(cal_result[92]), .B1(
        n222), .Y(n1062) );
  OAI2BB1X1 U280 ( .A0N(n225), .A1N(result_reg8[94]), .B0(n1064), .Y(n864) );
  AOI22X1 U281 ( .A0(result_reg8[110]), .A1(n216), .B0(cal_result[94]), .B1(
        n222), .Y(n1064) );
  OAI2BB1X1 U282 ( .A0N(n225), .A1N(result_reg8[107]), .B0(n1077), .Y(n877) );
  AOI22X1 U283 ( .A0(n1081), .A1(result_reg8[123]), .B0(cal_result[107]), .B1(
        n220), .Y(n1077) );
  OAI2BB1X1 U284 ( .A0N(n225), .A1N(result_reg8[108]), .B0(n1078), .Y(n878) );
  AOI22X1 U285 ( .A0(n218), .A1(result_reg8[124]), .B0(cal_result[108]), .B1(
        n220), .Y(n1078) );
  OAI2BB1X1 U286 ( .A0N(n225), .A1N(result_reg8[110]), .B0(n1080), .Y(n880) );
  AOI22X1 U287 ( .A0(n216), .A1(result_reg8[126]), .B0(cal_result[110]), .B1(
        n220), .Y(n1080) );
  NAND2X1 U288 ( .A(ready8), .B(n745), .Y(n1099) );
  OAI2BB2X1 U289 ( .B0(n106), .B1(n743), .A0N(n135), .A1N(result_reg4[64]), 
        .Y(n755) );
  OAI2BB2X1 U290 ( .B0(n105), .B1(n742), .A0N(n136), .A1N(result_reg4[65]), 
        .Y(n757) );
  OAI2BB2X1 U291 ( .B0(n103), .B1(n741), .A0N(n136), .A1N(result_reg4[66]), 
        .Y(n759) );
  OAI2BB2X1 U292 ( .B0(n100), .B1(n740), .A0N(n136), .A1N(result_reg4[67]), 
        .Y(n761) );
  OAI2BB2X1 U293 ( .B0(n107), .B1(n739), .A0N(n136), .A1N(result_reg4[68]), 
        .Y(n763) );
  OAI2BB2X1 U294 ( .B0(n100), .B1(n738), .A0N(n137), .A1N(result_reg4[69]), 
        .Y(n765) );
  OAI2BB2X1 U295 ( .B0(n101), .B1(n737), .A0N(n135), .A1N(result_reg4[70]), 
        .Y(n767) );
  OAI2BB2X1 U296 ( .B0(n104), .B1(n736), .A0N(n135), .A1N(result_reg4[71]), 
        .Y(n769) );
  OAI2BB2X1 U297 ( .B0(n107), .B1(n735), .A0N(n136), .A1N(result_reg4[72]), 
        .Y(n771) );
  OAI2BB2X1 U298 ( .B0(n103), .B1(n734), .A0N(n135), .A1N(result_reg4[73]), 
        .Y(n773) );
  OAI2BB2X1 U299 ( .B0(n102), .B1(n733), .A0N(n137), .A1N(result_reg4[74]), 
        .Y(n775) );
  OAI2BB2X1 U300 ( .B0(n101), .B1(n732), .A0N(n136), .A1N(result_reg4[75]), 
        .Y(n777) );
  OAI2BB2X1 U301 ( .B0(n102), .B1(n731), .A0N(n137), .A1N(result_reg4[76]), 
        .Y(n779) );
  OAI2BB2X1 U302 ( .B0(n105), .B1(n730), .A0N(n137), .A1N(result_reg4[77]), 
        .Y(n781) );
  OAI2BB2X1 U303 ( .B0(n106), .B1(n729), .A0N(n137), .A1N(result_reg4[78]), 
        .Y(n783) );
  OAI2BB2X1 U304 ( .B0(n104), .B1(n728), .A0N(n137), .A1N(result_reg4[79]), 
        .Y(n785) );
  INVX1 U305 ( .A(mode[0]), .Y(n1124) );
  INVX1 U306 ( .A(n1093), .Y(n1264) );
  AOI22X1 U307 ( .A0(n228), .A1(result_reg8[122]), .B0(cal_result[122]), .B1(
        n222), .Y(n1093) );
  INVX1 U308 ( .A(n1094), .Y(n1265) );
  AOI22X1 U309 ( .A0(n225), .A1(result_reg8[123]), .B0(cal_result[123]), .B1(
        n220), .Y(n1094) );
  INVX1 U310 ( .A(n1095), .Y(n1266) );
  AOI22X1 U311 ( .A0(n1100), .A1(result_reg8[124]), .B0(cal_result[124]), .B1(
        n220), .Y(n1095) );
  INVX1 U312 ( .A(n1097), .Y(n1268) );
  AOI22X1 U313 ( .A0(n1100), .A1(result_reg8[126]), .B0(cal_result[126]), .B1(
        n222), .Y(n1097) );
  OAI2BB1X1 U314 ( .A0N(n226), .A1N(result_reg8[74]), .B0(n1044), .Y(n844) );
  AOI22X1 U315 ( .A0(result_reg8[90]), .A1(n216), .B0(cal_result[74]), .B1(
        n222), .Y(n1044) );
  OAI2BB1X1 U316 ( .A0N(n226), .A1N(result_reg8[77]), .B0(n1047), .Y(n847) );
  AOI22X1 U317 ( .A0(result_reg8[93]), .A1(n218), .B0(cal_result[77]), .B1(
        n222), .Y(n1047) );
  OAI2BB1X1 U318 ( .A0N(n225), .A1N(result_reg8[90]), .B0(n1060), .Y(n860) );
  AOI22X1 U319 ( .A0(result_reg8[106]), .A1(n216), .B0(cal_result[90]), .B1(
        n222), .Y(n1060) );
  OAI2BB1X1 U320 ( .A0N(n226), .A1N(result_reg8[93]), .B0(n1063), .Y(n863) );
  AOI22X1 U321 ( .A0(result_reg8[109]), .A1(n216), .B0(cal_result[93]), .B1(
        n222), .Y(n1063) );
  OAI2BB1X1 U322 ( .A0N(n225), .A1N(result_reg8[106]), .B0(n1076), .Y(n876) );
  AOI22X1 U323 ( .A0(n216), .A1(result_reg8[122]), .B0(cal_result[106]), .B1(
        n220), .Y(n1076) );
  OAI2BB1X1 U324 ( .A0N(n225), .A1N(result_reg8[109]), .B0(n1079), .Y(n879) );
  AOI22X1 U325 ( .A0(n1081), .A1(result_reg8[125]), .B0(cal_result[109]), .B1(
        n220), .Y(n1079) );
  INVX1 U326 ( .A(n904), .Y(n1142) );
  AOI22X1 U327 ( .A0(n92), .A1(result_reg4[32]), .B0(n121), .B1(
        result_reg4[16]), .Y(n904) );
  INVX1 U328 ( .A(n903), .Y(n1158) );
  AOI22X1 U329 ( .A0(n92), .A1(result_reg4[48]), .B0(n116), .B1(
        result_reg4[32]), .Y(n903) );
  INVX1 U330 ( .A(n902), .Y(n1174) );
  AOI22X1 U331 ( .A0(n92), .A1(result_reg4[64]), .B0(n114), .B1(
        result_reg4[48]), .Y(n902) );
  INVX1 U332 ( .A(n908), .Y(n1143) );
  AOI22X1 U333 ( .A0(n93), .A1(result_reg4[33]), .B0(n122), .B1(
        result_reg4[17]), .Y(n908) );
  INVX1 U334 ( .A(n907), .Y(n1159) );
  AOI22X1 U335 ( .A0(n92), .A1(result_reg4[49]), .B0(n122), .B1(
        result_reg4[33]), .Y(n907) );
  INVX1 U336 ( .A(n906), .Y(n1175) );
  AOI22X1 U337 ( .A0(n93), .A1(result_reg4[65]), .B0(n131), .B1(
        result_reg4[49]), .Y(n906) );
  INVX1 U338 ( .A(n912), .Y(n1144) );
  AOI22X1 U339 ( .A0(n92), .A1(result_reg4[34]), .B0(n127), .B1(
        result_reg4[18]), .Y(n912) );
  INVX1 U340 ( .A(n911), .Y(n1160) );
  AOI22X1 U341 ( .A0(n93), .A1(result_reg4[50]), .B0(n118), .B1(
        result_reg4[34]), .Y(n911) );
  INVX1 U342 ( .A(n910), .Y(n1176) );
  AOI22X1 U343 ( .A0(n92), .A1(result_reg4[66]), .B0(n119), .B1(
        result_reg4[50]), .Y(n910) );
  INVX1 U344 ( .A(n916), .Y(n1145) );
  AOI22X1 U345 ( .A0(n94), .A1(result_reg4[35]), .B0(n126), .B1(
        result_reg4[19]), .Y(n916) );
  INVX1 U346 ( .A(n915), .Y(n1161) );
  AOI22X1 U347 ( .A0(n92), .A1(result_reg4[51]), .B0(n129), .B1(
        result_reg4[35]), .Y(n915) );
  INVX1 U348 ( .A(n914), .Y(n1177) );
  AOI22X1 U349 ( .A0(n93), .A1(result_reg4[67]), .B0(n124), .B1(
        result_reg4[51]), .Y(n914) );
  INVX1 U350 ( .A(n920), .Y(n1146) );
  AOI22X1 U351 ( .A0(n93), .A1(result_reg4[36]), .B0(n129), .B1(
        result_reg4[20]), .Y(n920) );
  INVX1 U352 ( .A(n919), .Y(n1162) );
  AOI22X1 U353 ( .A0(n93), .A1(result_reg4[52]), .B0(n131), .B1(
        result_reg4[36]), .Y(n919) );
  INVX1 U354 ( .A(n918), .Y(n1178) );
  AOI22X1 U355 ( .A0(n93), .A1(result_reg4[68]), .B0(n132), .B1(
        result_reg4[52]), .Y(n918) );
  INVX1 U356 ( .A(n924), .Y(n1147) );
  AOI22X1 U357 ( .A0(n94), .A1(result_reg4[37]), .B0(n130), .B1(
        result_reg4[21]), .Y(n924) );
  INVX1 U358 ( .A(n923), .Y(n1163) );
  AOI22X1 U359 ( .A0(n93), .A1(result_reg4[53]), .B0(n123), .B1(
        result_reg4[37]), .Y(n923) );
  INVX1 U360 ( .A(n922), .Y(n1179) );
  AOI22X1 U361 ( .A0(n93), .A1(result_reg4[69]), .B0(n130), .B1(
        result_reg4[53]), .Y(n922) );
  INVX1 U362 ( .A(n928), .Y(n1148) );
  AOI22X1 U363 ( .A0(n94), .A1(result_reg4[38]), .B0(n123), .B1(
        result_reg4[22]), .Y(n928) );
  INVX1 U364 ( .A(n927), .Y(n1164) );
  AOI22X1 U365 ( .A0(n94), .A1(result_reg4[54]), .B0(n125), .B1(
        result_reg4[38]), .Y(n927) );
  INVX1 U366 ( .A(n926), .Y(n1180) );
  AOI22X1 U367 ( .A0(n93), .A1(result_reg4[70]), .B0(n131), .B1(
        result_reg4[54]), .Y(n926) );
  INVX1 U368 ( .A(n932), .Y(n1149) );
  AOI22X1 U369 ( .A0(n94), .A1(result_reg4[39]), .B0(n125), .B1(
        result_reg4[23]), .Y(n932) );
  INVX1 U370 ( .A(n931), .Y(n1165) );
  AOI22X1 U371 ( .A0(n94), .A1(result_reg4[55]), .B0(n132), .B1(
        result_reg4[39]), .Y(n931) );
  INVX1 U372 ( .A(n930), .Y(n1181) );
  AOI22X1 U373 ( .A0(n94), .A1(result_reg4[71]), .B0(n124), .B1(
        result_reg4[55]), .Y(n930) );
  INVX1 U374 ( .A(n936), .Y(n1150) );
  AOI22X1 U375 ( .A0(n94), .A1(result_reg4[40]), .B0(n128), .B1(
        result_reg4[24]), .Y(n936) );
  INVX1 U376 ( .A(n935), .Y(n1166) );
  AOI22X1 U377 ( .A0(n95), .A1(result_reg4[56]), .B0(n128), .B1(
        result_reg4[40]), .Y(n935) );
  INVX1 U378 ( .A(n934), .Y(n1182) );
  AOI22X1 U379 ( .A0(n94), .A1(result_reg4[72]), .B0(n127), .B1(
        result_reg4[56]), .Y(n934) );
  INVX1 U380 ( .A(n940), .Y(n1151) );
  AOI22X1 U381 ( .A0(n95), .A1(result_reg4[41]), .B0(n115), .B1(
        result_reg4[25]), .Y(n940) );
  INVX1 U382 ( .A(n939), .Y(n1167) );
  AOI22X1 U383 ( .A0(n94), .A1(result_reg4[57]), .B0(n117), .B1(
        result_reg4[41]), .Y(n939) );
  INVX1 U384 ( .A(n938), .Y(n1183) );
  AOI22X1 U385 ( .A0(n95), .A1(result_reg4[73]), .B0(n126), .B1(
        result_reg4[57]), .Y(n938) );
  INVX1 U386 ( .A(n944), .Y(n1152) );
  AOI22X1 U387 ( .A0(n95), .A1(result_reg4[42]), .B0(n120), .B1(
        result_reg4[26]), .Y(n944) );
  INVX1 U388 ( .A(n943), .Y(n1168) );
  AOI22X1 U389 ( .A0(n95), .A1(result_reg4[58]), .B0(n120), .B1(
        result_reg4[42]), .Y(n943) );
  INVX1 U390 ( .A(n942), .Y(n1184) );
  AOI22X1 U391 ( .A0(n95), .A1(result_reg4[74]), .B0(n116), .B1(
        result_reg4[58]), .Y(n942) );
  INVX1 U392 ( .A(n948), .Y(n1153) );
  AOI22X1 U393 ( .A0(n95), .A1(result_reg4[43]), .B0(n129), .B1(
        result_reg4[27]), .Y(n948) );
  INVX1 U394 ( .A(n947), .Y(n1169) );
  AOI22X1 U395 ( .A0(n95), .A1(result_reg4[59]), .B0(n128), .B1(
        result_reg4[43]), .Y(n947) );
  INVX1 U396 ( .A(n946), .Y(n1185) );
  AOI22X1 U397 ( .A0(n95), .A1(result_reg4[75]), .B0(n120), .B1(
        result_reg4[59]), .Y(n946) );
  INVX1 U398 ( .A(n952), .Y(n1154) );
  AOI22X1 U399 ( .A0(n96), .A1(result_reg4[44]), .B0(n113), .B1(
        result_reg4[28]), .Y(n952) );
  INVX1 U400 ( .A(n951), .Y(n1170) );
  AOI22X1 U401 ( .A0(n96), .A1(result_reg4[60]), .B0(n116), .B1(
        result_reg4[44]), .Y(n951) );
  INVX1 U402 ( .A(n950), .Y(n1186) );
  AOI22X1 U403 ( .A0(n95), .A1(result_reg4[76]), .B0(n113), .B1(
        result_reg4[60]), .Y(n950) );
  INVX1 U404 ( .A(n956), .Y(n1155) );
  AOI22X1 U405 ( .A0(n96), .A1(result_reg4[45]), .B0(n121), .B1(
        result_reg4[29]), .Y(n956) );
  INVX1 U406 ( .A(n955), .Y(n1171) );
  AOI22X1 U407 ( .A0(n96), .A1(result_reg4[61]), .B0(n115), .B1(
        result_reg4[45]), .Y(n955) );
  INVX1 U408 ( .A(n954), .Y(n1187) );
  AOI22X1 U409 ( .A0(n96), .A1(result_reg4[77]), .B0(n121), .B1(
        result_reg4[61]), .Y(n954) );
  INVX1 U410 ( .A(n960), .Y(n1156) );
  AOI22X1 U411 ( .A0(n96), .A1(result_reg4[46]), .B0(n117), .B1(
        result_reg4[30]), .Y(n960) );
  INVX1 U412 ( .A(n959), .Y(n1172) );
  AOI22X1 U413 ( .A0(n96), .A1(result_reg4[62]), .B0(n118), .B1(
        result_reg4[46]), .Y(n959) );
  INVX1 U414 ( .A(n958), .Y(n1188) );
  AOI22X1 U415 ( .A0(n96), .A1(result_reg4[78]), .B0(n114), .B1(
        result_reg4[62]), .Y(n958) );
  INVX1 U416 ( .A(n964), .Y(n1157) );
  AOI22X1 U417 ( .A0(n97), .A1(result_reg4[47]), .B0(n119), .B1(
        result_reg4[31]), .Y(n964) );
  INVX1 U418 ( .A(n963), .Y(n1173) );
  AOI22X1 U419 ( .A0(n97), .A1(result_reg4[63]), .B0(n114), .B1(
        result_reg4[47]), .Y(n963) );
  INVX1 U420 ( .A(n962), .Y(n1189) );
  AOI22X1 U421 ( .A0(n97), .A1(result_reg4[79]), .B0(n130), .B1(
        result_reg4[63]), .Y(n962) );
  INVX1 U422 ( .A(n905), .Y(n1126) );
  AOI22X1 U423 ( .A0(n92), .A1(result_reg4[16]), .B0(result_reg4[0]), .B1(n112), .Y(n905) );
  INVX1 U424 ( .A(n909), .Y(n1127) );
  AOI22X1 U425 ( .A0(n92), .A1(result_reg4[17]), .B0(result_reg4[1]), .B1(n111), .Y(n909) );
  INVX1 U426 ( .A(n913), .Y(n1128) );
  AOI22X1 U427 ( .A0(n93), .A1(result_reg4[18]), .B0(result_reg4[2]), .B1(n112), .Y(n913) );
  INVX1 U428 ( .A(n917), .Y(n1129) );
  AOI22X1 U429 ( .A0(n93), .A1(result_reg4[19]), .B0(result_reg4[3]), .B1(n132), .Y(n917) );
  INVX1 U430 ( .A(n921), .Y(n1130) );
  AOI22X1 U431 ( .A0(n94), .A1(result_reg4[20]), .B0(result_reg4[4]), .B1(n110), .Y(n921) );
  INVX1 U432 ( .A(n925), .Y(n1131) );
  AOI22X1 U433 ( .A0(n93), .A1(result_reg4[21]), .B0(result_reg4[5]), .B1(n108), .Y(n925) );
  INVX1 U434 ( .A(n929), .Y(n1132) );
  AOI22X1 U435 ( .A0(n94), .A1(result_reg4[22]), .B0(result_reg4[6]), .B1(n109), .Y(n929) );
  INVX1 U436 ( .A(n933), .Y(n1133) );
  AOI22X1 U437 ( .A0(n94), .A1(result_reg4[23]), .B0(result_reg4[7]), .B1(n112), .Y(n933) );
  INVX1 U438 ( .A(n937), .Y(n1134) );
  AOI22X1 U439 ( .A0(n95), .A1(result_reg4[24]), .B0(result_reg4[8]), .B1(n110), .Y(n937) );
  INVX1 U440 ( .A(n941), .Y(n1135) );
  AOI22X1 U441 ( .A0(n95), .A1(result_reg4[25]), .B0(result_reg4[9]), .B1(n108), .Y(n941) );
  INVX1 U442 ( .A(n945), .Y(n1136) );
  AOI22X1 U443 ( .A0(n96), .A1(result_reg4[26]), .B0(result_reg4[10]), .B1(
        n111), .Y(n945) );
  INVX1 U444 ( .A(n949), .Y(n1137) );
  AOI22X1 U445 ( .A0(n95), .A1(result_reg4[27]), .B0(result_reg4[11]), .B1(
        n110), .Y(n949) );
  INVX1 U446 ( .A(n953), .Y(n1138) );
  AOI22X1 U447 ( .A0(n96), .A1(result_reg4[28]), .B0(result_reg4[12]), .B1(
        n109), .Y(n953) );
  INVX1 U448 ( .A(n957), .Y(n1139) );
  AOI22X1 U449 ( .A0(n96), .A1(result_reg4[29]), .B0(result_reg4[13]), .B1(
        n112), .Y(n957) );
  INVX1 U450 ( .A(n961), .Y(n1140) );
  AOI22X1 U451 ( .A0(n96), .A1(result_reg4[30]), .B0(result_reg4[14]), .B1(
        n111), .Y(n961) );
  INVX1 U452 ( .A(n965), .Y(n1141) );
  AOI22X1 U453 ( .A0(n96), .A1(result_reg4[31]), .B0(result_reg4[15]), .B1(
        n111), .Y(n965) );
  INVX1 U454 ( .A(n970), .Y(n1190) );
  AOI222X1 U455 ( .A0(n220), .A1(cal_result[0]), .B0(n1081), .B1(
        result_reg8[16]), .C0(n226), .C1(result_reg8[0]), .Y(n970) );
  INVX1 U456 ( .A(n971), .Y(n1191) );
  AOI222X1 U457 ( .A0(n220), .A1(cal_result[1]), .B0(n1081), .B1(
        result_reg8[17]), .C0(n228), .C1(result_reg8[1]), .Y(n971) );
  INVX1 U458 ( .A(n972), .Y(n1192) );
  AOI222X1 U459 ( .A0(n222), .A1(cal_result[2]), .B0(n218), .B1(
        result_reg8[18]), .C0(n228), .C1(result_reg8[2]), .Y(n972) );
  INVX1 U460 ( .A(n973), .Y(n1193) );
  AOI222X1 U461 ( .A0(n220), .A1(cal_result[3]), .B0(n218), .B1(
        result_reg8[19]), .C0(n228), .C1(result_reg8[3]), .Y(n973) );
  INVX1 U462 ( .A(n974), .Y(n1194) );
  AOI222X1 U463 ( .A0(n224), .A1(cal_result[4]), .B0(n218), .B1(
        result_reg8[20]), .C0(n228), .C1(result_reg8[4]), .Y(n974) );
  INVX1 U464 ( .A(n975), .Y(n1195) );
  AOI222X1 U465 ( .A0(n224), .A1(cal_result[5]), .B0(n218), .B1(
        result_reg8[21]), .C0(n228), .C1(result_reg8[5]), .Y(n975) );
  INVX1 U466 ( .A(n976), .Y(n1196) );
  AOI222X1 U467 ( .A0(n224), .A1(cal_result[6]), .B0(n218), .B1(
        result_reg8[22]), .C0(n228), .C1(result_reg8[6]), .Y(n976) );
  INVX1 U468 ( .A(n977), .Y(n1197) );
  AOI222X1 U469 ( .A0(n224), .A1(cal_result[7]), .B0(n218), .B1(
        result_reg8[23]), .C0(n228), .C1(result_reg8[7]), .Y(n977) );
  INVX1 U470 ( .A(n978), .Y(n1198) );
  AOI222X1 U471 ( .A0(n224), .A1(cal_result[8]), .B0(n218), .B1(
        result_reg8[24]), .C0(n228), .C1(result_reg8[8]), .Y(n978) );
  INVX1 U472 ( .A(n979), .Y(n1199) );
  AOI222X1 U473 ( .A0(n224), .A1(cal_result[9]), .B0(n218), .B1(
        result_reg8[25]), .C0(n228), .C1(result_reg8[9]), .Y(n979) );
  INVX1 U474 ( .A(n980), .Y(n1200) );
  AOI222X1 U475 ( .A0(n224), .A1(cal_result[10]), .B0(n218), .B1(
        result_reg8[26]), .C0(n228), .C1(result_reg8[10]), .Y(n980) );
  INVX1 U476 ( .A(n981), .Y(n1201) );
  AOI222X1 U477 ( .A0(n224), .A1(cal_result[11]), .B0(n218), .B1(
        result_reg8[27]), .C0(n228), .C1(result_reg8[11]), .Y(n981) );
  INVX1 U478 ( .A(n982), .Y(n1202) );
  AOI222X1 U479 ( .A0(n224), .A1(cal_result[12]), .B0(n218), .B1(
        result_reg8[28]), .C0(n228), .C1(result_reg8[12]), .Y(n982) );
  INVX1 U480 ( .A(n986), .Y(n1206) );
  AOI222X1 U481 ( .A0(n224), .A1(cal_result[16]), .B0(n217), .B1(
        result_reg8[32]), .C0(n228), .C1(result_reg8[16]), .Y(n986) );
  INVX1 U482 ( .A(n987), .Y(n1207) );
  AOI222X1 U483 ( .A0(n224), .A1(cal_result[17]), .B0(n217), .B1(
        result_reg8[33]), .C0(n228), .C1(result_reg8[17]), .Y(n987) );
  INVX1 U484 ( .A(n988), .Y(n1208) );
  AOI222X1 U485 ( .A0(n224), .A1(cal_result[18]), .B0(n217), .B1(
        result_reg8[34]), .C0(n228), .C1(result_reg8[18]), .Y(n988) );
  INVX1 U486 ( .A(n989), .Y(n1209) );
  AOI222X1 U487 ( .A0(n224), .A1(cal_result[19]), .B0(n217), .B1(
        result_reg8[35]), .C0(n228), .C1(result_reg8[19]), .Y(n989) );
  INVX1 U488 ( .A(n990), .Y(n1210) );
  AOI222X1 U489 ( .A0(n224), .A1(cal_result[20]), .B0(n217), .B1(
        result_reg8[36]), .C0(n228), .C1(result_reg8[20]), .Y(n990) );
  INVX1 U490 ( .A(n991), .Y(n1211) );
  AOI222X1 U491 ( .A0(n224), .A1(cal_result[21]), .B0(n217), .B1(
        result_reg8[37]), .C0(n228), .C1(result_reg8[21]), .Y(n991) );
  INVX1 U492 ( .A(n992), .Y(n1212) );
  AOI222X1 U493 ( .A0(n224), .A1(cal_result[22]), .B0(n217), .B1(
        result_reg8[38]), .C0(n228), .C1(result_reg8[22]), .Y(n992) );
  INVX1 U494 ( .A(n993), .Y(n1213) );
  AOI222X1 U495 ( .A0(n224), .A1(cal_result[23]), .B0(n217), .B1(
        result_reg8[39]), .C0(n228), .C1(result_reg8[23]), .Y(n993) );
  INVX1 U496 ( .A(n994), .Y(n1214) );
  AOI222X1 U497 ( .A0(n224), .A1(cal_result[24]), .B0(n217), .B1(
        result_reg8[40]), .C0(n228), .C1(result_reg8[24]), .Y(n994) );
  INVX1 U498 ( .A(n995), .Y(n1215) );
  AOI222X1 U499 ( .A0(n224), .A1(cal_result[25]), .B0(n217), .B1(
        result_reg8[41]), .C0(n228), .C1(result_reg8[25]), .Y(n995) );
  INVX1 U500 ( .A(n996), .Y(n1216) );
  AOI222X1 U501 ( .A0(n224), .A1(cal_result[26]), .B0(n217), .B1(
        result_reg8[42]), .C0(n228), .C1(result_reg8[26]), .Y(n996) );
  INVX1 U502 ( .A(n997), .Y(n1217) );
  AOI222X1 U503 ( .A0(n224), .A1(cal_result[27]), .B0(n217), .B1(
        result_reg8[43]), .C0(n228), .C1(result_reg8[27]), .Y(n997) );
  INVX1 U504 ( .A(n998), .Y(n1218) );
  AOI222X1 U505 ( .A0(n224), .A1(cal_result[28]), .B0(n217), .B1(
        result_reg8[44]), .C0(n228), .C1(result_reg8[28]), .Y(n998) );
  INVX1 U506 ( .A(n1002), .Y(n1222) );
  AOI222X1 U507 ( .A0(n224), .A1(cal_result[32]), .B0(n217), .B1(
        result_reg8[48]), .C0(n227), .C1(result_reg8[32]), .Y(n1002) );
  INVX1 U508 ( .A(n1003), .Y(n1223) );
  AOI222X1 U509 ( .A0(n224), .A1(cal_result[33]), .B0(n217), .B1(
        result_reg8[49]), .C0(n227), .C1(result_reg8[33]), .Y(n1003) );
  INVX1 U510 ( .A(n1004), .Y(n1224) );
  AOI222X1 U511 ( .A0(n224), .A1(cal_result[34]), .B0(n217), .B1(
        result_reg8[50]), .C0(n227), .C1(result_reg8[34]), .Y(n1004) );
  INVX1 U512 ( .A(n1005), .Y(n1225) );
  AOI222X1 U513 ( .A0(n224), .A1(cal_result[35]), .B0(n217), .B1(
        result_reg8[51]), .C0(n227), .C1(result_reg8[35]), .Y(n1005) );
  INVX1 U514 ( .A(n1006), .Y(n1226) );
  AOI222X1 U515 ( .A0(n223), .A1(cal_result[36]), .B0(n217), .B1(
        result_reg8[52]), .C0(n227), .C1(result_reg8[36]), .Y(n1006) );
  INVX1 U516 ( .A(n1007), .Y(n1227) );
  AOI222X1 U517 ( .A0(n223), .A1(cal_result[37]), .B0(n217), .B1(
        result_reg8[53]), .C0(n227), .C1(result_reg8[37]), .Y(n1007) );
  INVX1 U518 ( .A(n1008), .Y(n1228) );
  AOI222X1 U519 ( .A0(n223), .A1(cal_result[38]), .B0(n217), .B1(
        result_reg8[54]), .C0(n227), .C1(result_reg8[38]), .Y(n1008) );
  INVX1 U520 ( .A(n1009), .Y(n1229) );
  AOI222X1 U521 ( .A0(n223), .A1(cal_result[39]), .B0(n217), .B1(
        result_reg8[55]), .C0(n227), .C1(result_reg8[39]), .Y(n1009) );
  INVX1 U522 ( .A(n1010), .Y(n1230) );
  AOI222X1 U523 ( .A0(n223), .A1(cal_result[40]), .B0(n217), .B1(
        result_reg8[56]), .C0(n227), .C1(result_reg8[40]), .Y(n1010) );
  INVX1 U524 ( .A(n1011), .Y(n1231) );
  AOI222X1 U525 ( .A0(n223), .A1(cal_result[41]), .B0(n217), .B1(
        result_reg8[57]), .C0(n227), .C1(result_reg8[41]), .Y(n1011) );
  INVX1 U526 ( .A(n1012), .Y(n1232) );
  AOI222X1 U527 ( .A0(n223), .A1(cal_result[42]), .B0(n217), .B1(
        result_reg8[58]), .C0(n227), .C1(result_reg8[42]), .Y(n1012) );
  INVX1 U528 ( .A(n1013), .Y(n1233) );
  AOI222X1 U529 ( .A0(n223), .A1(cal_result[43]), .B0(n217), .B1(
        result_reg8[59]), .C0(n227), .C1(result_reg8[43]), .Y(n1013) );
  INVX1 U530 ( .A(n1014), .Y(n1234) );
  AOI222X1 U531 ( .A0(n223), .A1(cal_result[44]), .B0(n217), .B1(
        result_reg8[60]), .C0(n227), .C1(result_reg8[44]), .Y(n1014) );
  INVX1 U532 ( .A(n1018), .Y(n1238) );
  AOI222X1 U533 ( .A0(n223), .A1(cal_result[48]), .B0(n216), .B1(
        result_reg8[64]), .C0(n227), .C1(result_reg8[48]), .Y(n1018) );
  INVX1 U534 ( .A(n1019), .Y(n1239) );
  AOI222X1 U535 ( .A0(n223), .A1(cal_result[49]), .B0(n218), .B1(
        result_reg8[65]), .C0(n227), .C1(result_reg8[49]), .Y(n1019) );
  INVX1 U536 ( .A(n1020), .Y(n1240) );
  AOI222X1 U537 ( .A0(n223), .A1(cal_result[50]), .B0(n216), .B1(
        result_reg8[66]), .C0(n227), .C1(result_reg8[50]), .Y(n1020) );
  INVX1 U538 ( .A(n1021), .Y(n1241) );
  AOI222X1 U539 ( .A0(n223), .A1(cal_result[51]), .B0(n218), .B1(
        result_reg8[67]), .C0(n227), .C1(result_reg8[51]), .Y(n1021) );
  INVX1 U540 ( .A(n1022), .Y(n1242) );
  AOI222X1 U541 ( .A0(n223), .A1(cal_result[52]), .B0(n216), .B1(
        result_reg8[68]), .C0(n227), .C1(result_reg8[52]), .Y(n1022) );
  INVX1 U542 ( .A(n1023), .Y(n1243) );
  AOI222X1 U543 ( .A0(n223), .A1(cal_result[53]), .B0(n218), .B1(
        result_reg8[69]), .C0(n227), .C1(result_reg8[53]), .Y(n1023) );
  INVX1 U544 ( .A(n1024), .Y(n1244) );
  AOI222X1 U545 ( .A0(n223), .A1(cal_result[54]), .B0(n216), .B1(
        result_reg8[70]), .C0(n227), .C1(result_reg8[54]), .Y(n1024) );
  INVX1 U546 ( .A(n1025), .Y(n1245) );
  AOI222X1 U547 ( .A0(n223), .A1(cal_result[55]), .B0(n218), .B1(
        result_reg8[71]), .C0(n227), .C1(result_reg8[55]), .Y(n1025) );
  INVX1 U548 ( .A(n1026), .Y(n1246) );
  AOI222X1 U549 ( .A0(n223), .A1(cal_result[56]), .B0(n1081), .B1(
        result_reg8[72]), .C0(n227), .C1(result_reg8[56]), .Y(n1026) );
  INVX1 U550 ( .A(n1027), .Y(n1247) );
  AOI222X1 U551 ( .A0(n223), .A1(cal_result[57]), .B0(n1081), .B1(
        result_reg8[73]), .C0(n227), .C1(result_reg8[57]), .Y(n1027) );
  INVX1 U552 ( .A(n1028), .Y(n1248) );
  AOI222X1 U553 ( .A0(n223), .A1(cal_result[58]), .B0(n1081), .B1(
        result_reg8[74]), .C0(n227), .C1(result_reg8[58]), .Y(n1028) );
  INVX1 U554 ( .A(n1029), .Y(n1249) );
  AOI222X1 U555 ( .A0(n223), .A1(cal_result[59]), .B0(n1081), .B1(
        result_reg8[75]), .C0(n227), .C1(result_reg8[59]), .Y(n1029) );
  INVX1 U556 ( .A(n1030), .Y(n1250) );
  AOI222X1 U557 ( .A0(n223), .A1(cal_result[60]), .B0(n1081), .B1(
        result_reg8[76]), .C0(n227), .C1(result_reg8[60]), .Y(n1030) );
  NOR2X1 U558 ( .A(start_reg4[0]), .B(ready8), .Y(n1123) );
  BUFX3 U559 ( .A(n1121), .Y(n86) );
  OAI21XL U560 ( .A0(n1104), .A1(mode_reg_0_), .B0(n1102), .Y(n1121) );
  OAI2BB2X1 U561 ( .B0(n82), .B1(n1122), .A0N(dout[0]), .A1N(n82), .Y(n898) );
  AOI22X1 U562 ( .A0(result_reg4[0]), .A1(n86), .B0(result_reg8[0]), .B1(n85), 
        .Y(n1122) );
  OAI2BB2X1 U563 ( .B0(n82), .B1(n1119), .A0N(dout[1]), .A1N(n82), .Y(n897) );
  AOI22X1 U564 ( .A0(result_reg4[1]), .A1(n86), .B0(result_reg8[1]), .B1(n85), 
        .Y(n1119) );
  OAI2BB2X1 U565 ( .B0(n82), .B1(n1118), .A0N(dout[2]), .A1N(n82), .Y(n896) );
  AOI22X1 U566 ( .A0(result_reg4[2]), .A1(n86), .B0(result_reg8[2]), .B1(n85), 
        .Y(n1118) );
  OAI2BB2X1 U567 ( .B0(n82), .B1(n1117), .A0N(dout[3]), .A1N(n82), .Y(n895) );
  AOI22X1 U568 ( .A0(result_reg4[3]), .A1(n86), .B0(result_reg8[3]), .B1(n85), 
        .Y(n1117) );
  OAI2BB2X1 U569 ( .B0(n82), .B1(n1116), .A0N(dout[4]), .A1N(n82), .Y(n894) );
  AOI22X1 U570 ( .A0(result_reg4[4]), .A1(n86), .B0(result_reg8[4]), .B1(n85), 
        .Y(n1116) );
  OAI2BB2X1 U571 ( .B0(n82), .B1(n1115), .A0N(dout[5]), .A1N(n82), .Y(n893) );
  AOI22X1 U572 ( .A0(result_reg4[5]), .A1(n86), .B0(result_reg8[5]), .B1(n85), 
        .Y(n1115) );
  OAI2BB2X1 U573 ( .B0(n82), .B1(n1114), .A0N(dout[6]), .A1N(n82), .Y(n892) );
  AOI22X1 U574 ( .A0(result_reg4[6]), .A1(n86), .B0(result_reg8[6]), .B1(n85), 
        .Y(n1114) );
  OAI2BB2X1 U575 ( .B0(n82), .B1(n1113), .A0N(dout[7]), .A1N(n82), .Y(n891) );
  AOI22X1 U576 ( .A0(result_reg4[7]), .A1(n86), .B0(result_reg8[7]), .B1(n85), 
        .Y(n1113) );
  OAI2BB2X1 U577 ( .B0(n82), .B1(n1112), .A0N(dout[8]), .A1N(n82), .Y(n890) );
  AOI22X1 U578 ( .A0(result_reg4[8]), .A1(n86), .B0(result_reg8[8]), .B1(n85), 
        .Y(n1112) );
  OAI2BB2X1 U579 ( .B0(n82), .B1(n1111), .A0N(dout[9]), .A1N(n82), .Y(n889) );
  AOI22X1 U580 ( .A0(result_reg4[9]), .A1(n86), .B0(result_reg8[9]), .B1(n85), 
        .Y(n1111) );
  OAI2BB2X1 U581 ( .B0(n82), .B1(n1110), .A0N(dout[10]), .A1N(n82), .Y(n888)
         );
  AOI22X1 U582 ( .A0(result_reg4[10]), .A1(n86), .B0(result_reg8[10]), .B1(n85), .Y(n1110) );
  OAI2BB2X1 U583 ( .B0(n82), .B1(n1109), .A0N(dout[11]), .A1N(n82), .Y(n887)
         );
  AOI22X1 U584 ( .A0(result_reg4[11]), .A1(n86), .B0(result_reg8[11]), .B1(n85), .Y(n1109) );
  OAI2BB2X1 U585 ( .B0(n82), .B1(n1108), .A0N(dout[12]), .A1N(n82), .Y(n886)
         );
  AOI22X1 U586 ( .A0(result_reg4[12]), .A1(n86), .B0(result_reg8[12]), .B1(n85), .Y(n1108) );
  OAI2BB2X1 U587 ( .B0(n82), .B1(n1107), .A0N(dout[13]), .A1N(n82), .Y(n885)
         );
  AOI22X1 U588 ( .A0(result_reg4[13]), .A1(n86), .B0(result_reg8[13]), .B1(n85), .Y(n1107) );
  OAI2BB2X1 U589 ( .B0(n82), .B1(n1106), .A0N(dout[14]), .A1N(n82), .Y(n884)
         );
  AOI22X1 U590 ( .A0(result_reg4[14]), .A1(n86), .B0(result_reg8[14]), .B1(n85), .Y(n1106) );
  OAI2BB2X1 U591 ( .B0(n82), .B1(n1105), .A0N(dout[15]), .A1N(n82), .Y(n883)
         );
  AOI22X1 U592 ( .A0(result_reg4[15]), .A1(n86), .B0(result_reg8[15]), .B1(n85), .Y(n1105) );
  BUFX3 U593 ( .A(n1120), .Y(n85) );
  OAI21XL U594 ( .A0(n1104), .A1(n744), .B0(n1103), .Y(n1120) );
  INVX1 U595 ( .A(mode_reg_0_), .Y(n744) );
  INVX1 U596 ( .A(ready8), .Y(n673) );
  INVX1 U597 ( .A(shift4_flag), .Y(n672) );
  INVX1 U598 ( .A(start_reg4[0]), .Y(n679) );
  OAI2BB1X1 U599 ( .A0N(n226), .A1N(result_reg8[68]), .B0(n1038), .Y(n838) );
  AOI22X1 U600 ( .A0(result_reg8[84]), .A1(n216), .B0(cal_result[68]), .B1(
        n220), .Y(n1038) );
  OAI2BB1X1 U601 ( .A0N(n226), .A1N(result_reg8[69]), .B0(n1039), .Y(n839) );
  AOI22X1 U602 ( .A0(result_reg8[85]), .A1(n218), .B0(cal_result[69]), .B1(
        n220), .Y(n1039) );
  OAI2BB1X1 U603 ( .A0N(n226), .A1N(result_reg8[70]), .B0(n1040), .Y(n840) );
  AOI22X1 U604 ( .A0(result_reg8[86]), .A1(n218), .B0(cal_result[70]), .B1(
        n222), .Y(n1040) );
  OAI2BB1X1 U605 ( .A0N(n226), .A1N(result_reg8[71]), .B0(n1041), .Y(n841) );
  AOI22X1 U606 ( .A0(result_reg8[87]), .A1(n216), .B0(cal_result[71]), .B1(
        n222), .Y(n1041) );
  OAI2BB1X1 U607 ( .A0N(n226), .A1N(result_reg8[72]), .B0(n1042), .Y(n842) );
  AOI22X1 U608 ( .A0(result_reg8[88]), .A1(n216), .B0(cal_result[72]), .B1(
        n220), .Y(n1042) );
  OAI2BB1X1 U609 ( .A0N(n226), .A1N(result_reg8[73]), .B0(n1043), .Y(n843) );
  AOI22X1 U610 ( .A0(result_reg8[89]), .A1(n218), .B0(cal_result[73]), .B1(
        n220), .Y(n1043) );
  OAI2BB1X1 U611 ( .A0N(n226), .A1N(result_reg8[80]), .B0(n1050), .Y(n850) );
  AOI22X1 U612 ( .A0(result_reg8[96]), .A1(n216), .B0(cal_result[80]), .B1(
        n220), .Y(n1050) );
  OAI2BB1X1 U613 ( .A0N(n226), .A1N(result_reg8[81]), .B0(n1051), .Y(n851) );
  AOI22X1 U614 ( .A0(result_reg8[97]), .A1(n218), .B0(cal_result[81]), .B1(
        n220), .Y(n1051) );
  OAI2BB1X1 U615 ( .A0N(n226), .A1N(result_reg8[82]), .B0(n1052), .Y(n852) );
  AOI22X1 U616 ( .A0(result_reg8[98]), .A1(n216), .B0(cal_result[82]), .B1(
        n222), .Y(n1052) );
  OAI2BB1X1 U617 ( .A0N(n226), .A1N(result_reg8[83]), .B0(n1053), .Y(n853) );
  AOI22X1 U618 ( .A0(result_reg8[99]), .A1(n216), .B0(cal_result[83]), .B1(
        n222), .Y(n1053) );
  OAI2BB1X1 U619 ( .A0N(n226), .A1N(result_reg8[84]), .B0(n1054), .Y(n854) );
  AOI22X1 U620 ( .A0(result_reg8[100]), .A1(n216), .B0(cal_result[84]), .B1(
        n222), .Y(n1054) );
  OAI2BB1X1 U621 ( .A0N(n226), .A1N(result_reg8[85]), .B0(n1055), .Y(n855) );
  AOI22X1 U622 ( .A0(result_reg8[101]), .A1(n216), .B0(cal_result[85]), .B1(
        n220), .Y(n1055) );
  OAI2BB1X1 U623 ( .A0N(n226), .A1N(result_reg8[86]), .B0(n1056), .Y(n856) );
  AOI22X1 U624 ( .A0(result_reg8[102]), .A1(n218), .B0(cal_result[86]), .B1(
        n222), .Y(n1056) );
  OAI2BB1X1 U625 ( .A0N(n226), .A1N(result_reg8[87]), .B0(n1057), .Y(n857) );
  AOI22X1 U626 ( .A0(result_reg8[103]), .A1(n216), .B0(cal_result[87]), .B1(
        n222), .Y(n1057) );
  OAI2BB1X1 U627 ( .A0N(n226), .A1N(result_reg8[88]), .B0(n1058), .Y(n858) );
  AOI22X1 U628 ( .A0(result_reg8[104]), .A1(n216), .B0(cal_result[88]), .B1(
        n222), .Y(n1058) );
  OAI2BB1X1 U629 ( .A0N(n226), .A1N(result_reg8[89]), .B0(n1059), .Y(n859) );
  AOI22X1 U630 ( .A0(result_reg8[105]), .A1(n216), .B0(cal_result[89]), .B1(
        n220), .Y(n1059) );
  OAI2BB1X1 U631 ( .A0N(n225), .A1N(result_reg8[96]), .B0(n1066), .Y(n866) );
  AOI22X1 U632 ( .A0(n216), .A1(result_reg8[112]), .B0(cal_result[96]), .B1(
        n222), .Y(n1066) );
  OAI2BB1X1 U633 ( .A0N(n225), .A1N(result_reg8[97]), .B0(n1067), .Y(n867) );
  AOI22X1 U634 ( .A0(n1081), .A1(result_reg8[113]), .B0(cal_result[97]), .B1(
        n222), .Y(n1067) );
  OAI2BB1X1 U635 ( .A0N(n225), .A1N(result_reg8[98]), .B0(n1068), .Y(n868) );
  AOI22X1 U636 ( .A0(n218), .A1(result_reg8[114]), .B0(cal_result[98]), .B1(
        n222), .Y(n1068) );
  OAI2BB1X1 U637 ( .A0N(n225), .A1N(result_reg8[99]), .B0(n1069), .Y(n869) );
  AOI22X1 U638 ( .A0(n1081), .A1(result_reg8[115]), .B0(cal_result[99]), .B1(
        n222), .Y(n1069) );
  OAI2BB1X1 U639 ( .A0N(n225), .A1N(result_reg8[100]), .B0(n1070), .Y(n870) );
  AOI22X1 U640 ( .A0(n216), .A1(result_reg8[116]), .B0(cal_result[100]), .B1(
        n222), .Y(n1070) );
  OAI2BB1X1 U641 ( .A0N(n225), .A1N(result_reg8[101]), .B0(n1071), .Y(n871) );
  AOI22X1 U642 ( .A0(n1081), .A1(result_reg8[117]), .B0(cal_result[101]), .B1(
        n222), .Y(n1071) );
  OAI2BB1X1 U643 ( .A0N(n225), .A1N(result_reg8[102]), .B0(n1072), .Y(n872) );
  AOI22X1 U644 ( .A0(n1081), .A1(result_reg8[118]), .B0(cal_result[102]), .B1(
        n222), .Y(n1072) );
  OAI2BB1X1 U645 ( .A0N(n225), .A1N(result_reg8[103]), .B0(n1073), .Y(n873) );
  AOI22X1 U646 ( .A0(n1081), .A1(result_reg8[119]), .B0(cal_result[103]), .B1(
        n222), .Y(n1073) );
  OAI2BB1X1 U647 ( .A0N(n225), .A1N(result_reg8[104]), .B0(n1074), .Y(n874) );
  AOI22X1 U648 ( .A0(n216), .A1(result_reg8[120]), .B0(cal_result[104]), .B1(
        n220), .Y(n1074) );
  OAI2BB1X1 U649 ( .A0N(n225), .A1N(result_reg8[105]), .B0(n1075), .Y(n875) );
  AOI22X1 U650 ( .A0(n1081), .A1(result_reg8[121]), .B0(cal_result[105]), .B1(
        n220), .Y(n1075) );
  OAI2BB1X1 U651 ( .A0N(n226), .A1N(result_reg8[64]), .B0(n1034), .Y(n834) );
  AOI22X1 U652 ( .A0(result_reg8[80]), .A1(n216), .B0(cal_result[64]), .B1(
        n223), .Y(n1034) );
  OAI2BB1X1 U653 ( .A0N(n226), .A1N(result_reg8[65]), .B0(n1035), .Y(n835) );
  AOI22X1 U654 ( .A0(result_reg8[81]), .A1(n218), .B0(cal_result[65]), .B1(
        n223), .Y(n1035) );
  OAI2BB1X1 U655 ( .A0N(n226), .A1N(result_reg8[66]), .B0(n1036), .Y(n836) );
  AOI22X1 U656 ( .A0(result_reg8[82]), .A1(n218), .B0(cal_result[66]), .B1(
        n223), .Y(n1036) );
  OAI2BB1X1 U657 ( .A0N(n226), .A1N(result_reg8[67]), .B0(n1037), .Y(n837) );
  AOI22X1 U658 ( .A0(result_reg8[83]), .A1(n218), .B0(cal_result[67]), .B1(
        n223), .Y(n1037) );
  INVX1 U659 ( .A(n1083), .Y(n1254) );
  AOI22X1 U660 ( .A0(n225), .A1(result_reg8[112]), .B0(cal_result[112]), .B1(
        n220), .Y(n1083) );
  INVX1 U661 ( .A(n1084), .Y(n1255) );
  AOI22X1 U662 ( .A0(n225), .A1(result_reg8[113]), .B0(cal_result[113]), .B1(
        n220), .Y(n1084) );
  INVX1 U663 ( .A(n1085), .Y(n1256) );
  AOI22X1 U664 ( .A0(n225), .A1(result_reg8[114]), .B0(cal_result[114]), .B1(
        n220), .Y(n1085) );
  INVX1 U665 ( .A(n1086), .Y(n1257) );
  AOI22X1 U666 ( .A0(n1100), .A1(result_reg8[115]), .B0(cal_result[115]), .B1(
        n220), .Y(n1086) );
  INVX1 U667 ( .A(n1087), .Y(n1258) );
  AOI22X1 U668 ( .A0(n225), .A1(result_reg8[116]), .B0(cal_result[116]), .B1(
        n222), .Y(n1087) );
  INVX1 U669 ( .A(n1088), .Y(n1259) );
  AOI22X1 U670 ( .A0(n1100), .A1(result_reg8[117]), .B0(cal_result[117]), .B1(
        n220), .Y(n1088) );
  INVX1 U671 ( .A(n1089), .Y(n1260) );
  AOI22X1 U672 ( .A0(n1100), .A1(result_reg8[118]), .B0(cal_result[118]), .B1(
        n222), .Y(n1089) );
  INVX1 U673 ( .A(n1090), .Y(n1261) );
  AOI22X1 U674 ( .A0(n1100), .A1(result_reg8[119]), .B0(cal_result[119]), .B1(
        n220), .Y(n1090) );
  INVX1 U675 ( .A(n1091), .Y(n1262) );
  AOI22X1 U676 ( .A0(n1100), .A1(result_reg8[120]), .B0(cal_result[120]), .B1(
        n220), .Y(n1091) );
  INVX1 U677 ( .A(n1092), .Y(n1263) );
  AOI22X1 U678 ( .A0(n1100), .A1(result_reg8[121]), .B0(cal_result[121]), .B1(
        n222), .Y(n1092) );
  OAI2BB2X1 U679 ( .B0(n673), .B1(n899), .A0N(n899), .A1N(start), .Y(n746) );
  OAI2BB1X1 U680 ( .A0N(mode[0]), .A1N(n968), .B0(n1099), .Y(n899) );
  OAI2BB1X1 U681 ( .A0N(n1102), .A1N(mode_reg_0_), .B0(n1099), .Y(n882) );
  INVX1 U682 ( .A(result_reg4[128]), .Y(n695) );
  INVX1 U683 ( .A(result_reg4[129]), .Y(n694) );
  INVX1 U684 ( .A(result_reg4[130]), .Y(n693) );
  INVX1 U685 ( .A(result_reg4[131]), .Y(n692) );
  INVX1 U686 ( .A(result_reg4[132]), .Y(n691) );
  INVX1 U687 ( .A(result_reg4[133]), .Y(n690) );
  INVX1 U688 ( .A(result_reg4[134]), .Y(n689) );
  INVX1 U689 ( .A(result_reg4[135]), .Y(n688) );
  INVX1 U690 ( .A(result_reg4[136]), .Y(n687) );
  INVX1 U691 ( .A(result_reg4[137]), .Y(n686) );
  INVX1 U692 ( .A(result_reg4[138]), .Y(n685) );
  INVX1 U693 ( .A(result_reg4[139]), .Y(n684) );
  INVX1 U694 ( .A(result_reg4[140]), .Y(n683) );
  INVX1 U695 ( .A(result_reg4[141]), .Y(n682) );
  INVX1 U696 ( .A(result_reg4[142]), .Y(n681) );
  INVX1 U697 ( .A(result_reg4[143]), .Y(n680) );
  INVX1 U698 ( .A(result_reg4[96]), .Y(n727) );
  INVX1 U699 ( .A(result_reg4[97]), .Y(n726) );
  INVX1 U700 ( .A(result_reg4[98]), .Y(n725) );
  INVX1 U701 ( .A(result_reg4[99]), .Y(n724) );
  INVX1 U702 ( .A(result_reg4[100]), .Y(n723) );
  INVX1 U703 ( .A(result_reg4[101]), .Y(n722) );
  INVX1 U704 ( .A(result_reg4[102]), .Y(n721) );
  INVX1 U705 ( .A(result_reg4[103]), .Y(n720) );
  INVX1 U706 ( .A(result_reg4[104]), .Y(n719) );
  INVX1 U707 ( .A(result_reg4[105]), .Y(n718) );
  INVX1 U708 ( .A(result_reg4[106]), .Y(n717) );
  INVX1 U709 ( .A(result_reg4[107]), .Y(n716) );
  INVX1 U710 ( .A(result_reg4[108]), .Y(n715) );
  INVX1 U711 ( .A(result_reg4[109]), .Y(n714) );
  INVX1 U712 ( .A(result_reg4[110]), .Y(n713) );
  INVX1 U713 ( .A(result_reg4[111]), .Y(n712) );
  INVX1 U714 ( .A(result_reg4[112]), .Y(n711) );
  INVX1 U715 ( .A(result_reg4[113]), .Y(n710) );
  INVX1 U716 ( .A(result_reg4[114]), .Y(n709) );
  INVX1 U717 ( .A(result_reg4[115]), .Y(n708) );
  INVX1 U718 ( .A(result_reg4[116]), .Y(n707) );
  INVX1 U719 ( .A(result_reg4[117]), .Y(n706) );
  INVX1 U720 ( .A(result_reg4[118]), .Y(n705) );
  INVX1 U721 ( .A(result_reg4[119]), .Y(n704) );
  INVX1 U722 ( .A(result_reg4[120]), .Y(n703) );
  INVX1 U723 ( .A(result_reg4[121]), .Y(n702) );
  INVX1 U724 ( .A(result_reg4[122]), .Y(n701) );
  INVX1 U725 ( .A(result_reg4[123]), .Y(n700) );
  INVX1 U726 ( .A(result_reg4[124]), .Y(n699) );
  INVX1 U727 ( .A(result_reg4[125]), .Y(n698) );
  INVX1 U728 ( .A(result_reg4[126]), .Y(n697) );
  INVX1 U729 ( .A(result_reg4[127]), .Y(n696) );
  INVX1 U730 ( .A(start_reg4[1]), .Y(n678) );
  INVX1 U731 ( .A(start_reg4[2]), .Y(n677) );
  INVX1 U732 ( .A(start_reg4[3]), .Y(n676) );
  INVX1 U733 ( .A(start_reg4[4]), .Y(n675) );
  INVX1 U734 ( .A(start_reg4[5]), .Y(n674) );
  INVX1 U735 ( .A(result_reg4[80]), .Y(n743) );
  INVX1 U736 ( .A(result_reg4[81]), .Y(n742) );
  INVX1 U737 ( .A(result_reg4[82]), .Y(n741) );
  INVX1 U738 ( .A(result_reg4[83]), .Y(n740) );
  INVX1 U739 ( .A(result_reg4[84]), .Y(n739) );
  INVX1 U740 ( .A(result_reg4[85]), .Y(n738) );
  INVX1 U741 ( .A(result_reg4[86]), .Y(n737) );
  INVX1 U742 ( .A(result_reg4[87]), .Y(n736) );
  INVX1 U743 ( .A(result_reg4[88]), .Y(n735) );
  INVX1 U744 ( .A(result_reg4[89]), .Y(n734) );
  INVX1 U745 ( .A(result_reg4[90]), .Y(n733) );
  INVX1 U746 ( .A(result_reg4[91]), .Y(n732) );
  INVX1 U747 ( .A(result_reg4[92]), .Y(n731) );
  INVX1 U748 ( .A(result_reg4[93]), .Y(n730) );
  INVX1 U749 ( .A(result_reg4[94]), .Y(n729) );
  INVX1 U750 ( .A(result_reg4[95]), .Y(n728) );
endmodule


module idct ( clk, rstn, mode, start, din, dout, dout_mode );
  input [1:0] mode;
  input [15:0] din;
  output [15:0] dout;
  output [1:0] dout_mode;
  input clk, rstn, start;
  wire   s2p_ready_col, even_odd_ready_col, idct_ready_col, p2s_ready_mem,
         en_ram8x8_1, wr_rd_ram8x8_1, en_ram8x8_2, wr_rd_ram8x8_2, en_ram4x4_1,
         wr_rd_ram4x4_1, en_ram4x4_2, wr_rd_ram4x4_2, en_ram4x4_3,
         wr_rd_ram4x4_3, en_ram4x4_4, wr_rd_ram4x4_4, ram8x8_1_ready,
         ram8x8_2_ready, ram4x4_1_ready, ram4x4_2_ready, ram4x4_3_ready,
         ram4x4_4_ready, mem_ctrl_tran_ready, s2p_ready_row,
         even_odd_ready_row, idct_ready_row, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n1, n2;
  wire   [255:0] idct_in_col;
  wire   [1:0] s2p1_mode;
  wire   [255:0] idct_in_col_tran;
  wire   [1:0] even_odd_col_mode;
  wire   [127:0] idct_out_col;
  wire   [1:0] idct_cal_col_mode;
  wire   [15:0] mem_in;
  wire   [1:0] p2s1_mode;
  wire   [5:0] addr_ram8x8_1;
  wire   [5:0] addr_ram8x8_2;
  wire   [3:0] addr_ram4x4_1;
  wire   [3:0] addr_ram4x4_2;
  wire   [3:0] addr_ram4x4_3;
  wire   [3:0] addr_ram4x4_4;
  wire   [1:0] mem_ctrl_tran_mode;
  wire   [15:0] dout8x8_1;
  wire   [15:0] dout8x8_2;
  wire   [15:0] dout4x4_1;
  wire   [15:0] dout4x4_2;
  wire   [15:0] dout4x4_3;
  wire   [15:0] dout4x4_4;
  wire   [15:0] ram_out_wire;
  wire   [255:0] idct_in_row;
  wire   [1:0] s2p2_mode;
  wire   [255:0] idct_in_row_tran;
  wire   [1:0] even_odd_row_mode;
  wire   [127:0] idct_out_row;
  wire   [1:0] idct_cal_row_mode;

  s2p_0 inst_s2p1 ( .clk(clk), .rstn(rstn), .start(start), .mode(mode), .din(
        din), .dout(idct_in_col), .s2p_ready(s2p_ready_col), .mode_out(
        s2p1_mode) );
  even_odd_0 even_odd_col ( .clk(clk), .rstn(rstn), .mode(s2p1_mode), .start(
        s2p_ready_col), .din(idct_in_col), .dout(idct_in_col_tran), 
        .even_odd_ready(even_odd_ready_col), .mode_out(even_odd_col_mode) );
  idct_cal_shift7_add64 idct_cal_col ( .clk(clk), .rstn(rstn), .mode(
        even_odd_col_mode), .start(even_odd_ready_col), .x0(
        idct_in_col_tran[255:240]), .x1(idct_in_col_tran[239:224]), .x2(
        idct_in_col_tran[223:208]), .x3(idct_in_col_tran[207:192]), .x4(
        idct_in_col_tran[191:176]), .x5(idct_in_col_tran[175:160]), .x6(
        idct_in_col_tran[159:144]), .x7(idct_in_col_tran[143:128]), .y0(
        idct_out_col[15:0]), .y1(idct_out_col[31:16]), .y2(idct_out_col[47:32]), .y3(idct_out_col[63:48]), .y4(idct_out_col[79:64]), .y5(idct_out_col[95:80]), 
        .y6(idct_out_col[111:96]), .y7(idct_out_col[127:112]), .idct_ready(
        idct_ready_col), .mode_out(idct_cal_col_mode) );
  p2s_0 inst_p2s1 ( .clk(clk), .rstn(rstn), .start(idct_ready_col), .mode(
        idct_cal_col_mode), .cal_result(idct_out_col), .dout(mem_in), 
        .p2s_ready(p2s_ready_mem), .mode_out(p2s1_mode) );
  mem_ctrl_tran inst_mem_ctrl_tran ( .clk(clk), .rstn(rstn), .start(
        p2s_ready_mem), .mode(p2s1_mode), .en_ram8x8_1(en_ram8x8_1), 
        .wr_rd_ram8x8_1(wr_rd_ram8x8_1), .addr_ram8x8_1(addr_ram8x8_1), 
        .en_ram8x8_2(en_ram8x8_2), .wr_rd_ram8x8_2(wr_rd_ram8x8_2), 
        .addr_ram8x8_2(addr_ram8x8_2), .en_ram4x4_1(en_ram4x4_1), 
        .wr_rd_ram4x4_1(wr_rd_ram4x4_1), .addr_ram4x4_1(addr_ram4x4_1), 
        .en_ram4x4_2(en_ram4x4_2), .wr_rd_ram4x4_2(wr_rd_ram4x4_2), 
        .addr_ram4x4_2(addr_ram4x4_2), .en_ram4x4_3(en_ram4x4_3), 
        .wr_rd_ram4x4_3(wr_rd_ram4x4_3), .addr_ram4x4_3(addr_ram4x4_3), 
        .en_ram4x4_4(en_ram4x4_4), .wr_rd_ram4x4_4(wr_rd_ram4x4_4), 
        .addr_ram4x4_4(addr_ram4x4_4), .ram8x8_1_ready(ram8x8_1_ready), 
        .ram8x8_2_ready(ram8x8_2_ready), .ram4x4_1_ready(ram4x4_1_ready), 
        .ram4x4_2_ready(ram4x4_2_ready), .ram4x4_3_ready(ram4x4_3_ready), 
        .ram4x4_4_ready(ram4x4_4_ready), .mode_out(mem_ctrl_tran_mode) );
  mem8x8_0 ram8x8_1 ( .clk(clk), .rstn(rstn), .en(en_ram8x8_1), .wr_rd(
        wr_rd_ram8x8_1), .addr(addr_ram8x8_1), .din(mem_in), .dout(dout8x8_1)
         );
  mem8x8_1 ram8x8_2 ( .clk(clk), .rstn(rstn), .en(en_ram8x8_2), .wr_rd(
        wr_rd_ram8x8_2), .addr(addr_ram8x8_2), .din(mem_in), .dout(dout8x8_2)
         );
  mem4x4_0 ram4x4_1 ( .clk(clk), .rstn(rstn), .en(en_ram4x4_1), .wr_rd(
        wr_rd_ram4x4_1), .addr(addr_ram4x4_1), .din(mem_in), .dout(dout4x4_1)
         );
  mem4x4_3 ram4x4_2 ( .clk(clk), .rstn(rstn), .en(en_ram4x4_2), .wr_rd(
        wr_rd_ram4x4_2), .addr(addr_ram4x4_2), .din(mem_in), .dout(dout4x4_2)
         );
  mem4x4_2 ram4x4_3 ( .clk(clk), .rstn(rstn), .en(en_ram4x4_3), .wr_rd(
        wr_rd_ram4x4_3), .addr(addr_ram4x4_3), .din(mem_in), .dout(dout4x4_3)
         );
  mem4x4_1 ram4x4_4 ( .clk(clk), .rstn(rstn), .en(en_ram4x4_4), .wr_rd(
        wr_rd_ram4x4_4), .addr(addr_ram4x4_4), .din(mem_in), .dout(dout4x4_4)
         );
  s2p_1 inst_s2p2 ( .clk(clk), .rstn(rstn), .start(mem_ctrl_tran_ready), 
        .mode(mem_ctrl_tran_mode), .din(ram_out_wire), .dout(idct_in_row), 
        .s2p_ready(s2p_ready_row), .mode_out(s2p2_mode) );
  even_odd_1 even_odd_row ( .clk(clk), .rstn(rstn), .mode(s2p2_mode), .start(
        s2p_ready_row), .din(idct_in_row), .dout(idct_in_row_tran), 
        .even_odd_ready(even_odd_ready_row), .mode_out(even_odd_row_mode) );
  idct_cal_shift12_add2048 idct_cal_row ( .clk(clk), .rstn(rstn), .mode(
        even_odd_row_mode), .start(even_odd_ready_row), .x0(
        idct_in_row_tran[255:240]), .x1(idct_in_row_tran[239:224]), .x2(
        idct_in_row_tran[223:208]), .x3(idct_in_row_tran[207:192]), .x4(
        idct_in_row_tran[191:176]), .x5(idct_in_row_tran[175:160]), .x6(
        idct_in_row_tran[159:144]), .x7(idct_in_row_tran[143:128]), .y0(
        idct_out_row[15:0]), .y1(idct_out_row[31:16]), .y2(idct_out_row[47:32]), .y3(idct_out_row[63:48]), .y4(idct_out_row[79:64]), .y5(idct_out_row[95:80]), 
        .y6(idct_out_row[111:96]), .y7(idct_out_row[127:112]), .idct_ready(
        idct_ready_row), .mode_out(idct_cal_row_mode) );
  p2s_1 inst_p2s2 ( .clk(clk), .rstn(rstn), .start(idct_ready_row), .mode(
        idct_cal_row_mode), .cal_result(idct_out_row), .dout(dout), .mode_out(
        dout_mode) );
  NAND2X1 U1 ( .A(n25), .B(n26), .Y(ram_out_wire[1]) );
  AOI222X1 U2 ( .A0(dout8x8_2[1]), .A1(n8), .B0(dout4x4_2[1]), .B1(n9), .C0(
        dout4x4_1[1]), .C1(n10), .Y(n25) );
  AOI222X1 U3 ( .A0(dout4x4_3[1]), .A1(n5), .B0(dout8x8_1[1]), .B1(n6), .C0(
        dout4x4_4[1]), .C1(n7), .Y(n26) );
  NAND2X1 U4 ( .A(n23), .B(n24), .Y(ram_out_wire[2]) );
  AOI222X1 U5 ( .A0(dout8x8_2[2]), .A1(n8), .B0(dout4x4_2[2]), .B1(n9), .C0(
        dout4x4_1[2]), .C1(n10), .Y(n23) );
  AOI222X1 U6 ( .A0(dout4x4_3[2]), .A1(n5), .B0(dout8x8_1[2]), .B1(n6), .C0(
        dout4x4_4[2]), .C1(n7), .Y(n24) );
  NAND2X1 U7 ( .A(n21), .B(n22), .Y(ram_out_wire[3]) );
  AOI222X1 U8 ( .A0(dout8x8_2[3]), .A1(n8), .B0(dout4x4_2[3]), .B1(n9), .C0(
        dout4x4_1[3]), .C1(n10), .Y(n21) );
  AOI222X1 U9 ( .A0(dout4x4_3[3]), .A1(n5), .B0(dout8x8_1[3]), .B1(n6), .C0(
        dout4x4_4[3]), .C1(n7), .Y(n22) );
  NAND2X1 U10 ( .A(n19), .B(n20), .Y(ram_out_wire[4]) );
  AOI222X1 U11 ( .A0(dout8x8_2[4]), .A1(n8), .B0(dout4x4_2[4]), .B1(n9), .C0(
        dout4x4_1[4]), .C1(n10), .Y(n19) );
  AOI222X1 U12 ( .A0(dout4x4_3[4]), .A1(n5), .B0(dout8x8_1[4]), .B1(n6), .C0(
        dout4x4_4[4]), .C1(n7), .Y(n20) );
  NAND2X1 U13 ( .A(n17), .B(n18), .Y(ram_out_wire[5]) );
  AOI222X1 U14 ( .A0(dout8x8_2[5]), .A1(n8), .B0(dout4x4_2[5]), .B1(n9), .C0(
        dout4x4_1[5]), .C1(n10), .Y(n17) );
  AOI222X1 U15 ( .A0(dout4x4_3[5]), .A1(n5), .B0(dout8x8_1[5]), .B1(n6), .C0(
        dout4x4_4[5]), .C1(n7), .Y(n18) );
  NAND2X1 U16 ( .A(n15), .B(n16), .Y(ram_out_wire[6]) );
  AOI222X1 U17 ( .A0(dout8x8_2[6]), .A1(n8), .B0(dout4x4_2[6]), .B1(n9), .C0(
        dout4x4_1[6]), .C1(n10), .Y(n15) );
  AOI222X1 U18 ( .A0(dout4x4_3[6]), .A1(n5), .B0(dout8x8_1[6]), .B1(n6), .C0(
        dout4x4_4[6]), .C1(n7), .Y(n16) );
  NAND2X1 U19 ( .A(n13), .B(n14), .Y(ram_out_wire[7]) );
  AOI222X1 U20 ( .A0(dout8x8_2[7]), .A1(n8), .B0(dout4x4_2[7]), .B1(n9), .C0(
        dout4x4_1[7]), .C1(n10), .Y(n13) );
  AOI222X1 U21 ( .A0(dout4x4_3[7]), .A1(n5), .B0(dout8x8_1[7]), .B1(n6), .C0(
        dout4x4_4[7]), .C1(n7), .Y(n14) );
  NAND2X1 U22 ( .A(n11), .B(n12), .Y(ram_out_wire[8]) );
  AOI222X1 U23 ( .A0(dout8x8_2[8]), .A1(n8), .B0(dout4x4_2[8]), .B1(n9), .C0(
        dout4x4_1[8]), .C1(n10), .Y(n11) );
  AOI222X1 U24 ( .A0(dout4x4_3[8]), .A1(n5), .B0(dout8x8_1[8]), .B1(n6), .C0(
        dout4x4_4[8]), .C1(n7), .Y(n12) );
  NAND2X1 U25 ( .A(n3), .B(n4), .Y(ram_out_wire[9]) );
  AOI222X1 U26 ( .A0(dout8x8_2[9]), .A1(n8), .B0(dout4x4_2[9]), .B1(n9), .C0(
        dout4x4_1[9]), .C1(n10), .Y(n3) );
  AOI222X1 U27 ( .A0(dout4x4_3[9]), .A1(n5), .B0(dout8x8_1[9]), .B1(n6), .C0(
        dout4x4_4[9]), .C1(n7), .Y(n4) );
  NAND2X1 U28 ( .A(n37), .B(n38), .Y(ram_out_wire[10]) );
  AOI222X1 U29 ( .A0(dout8x8_2[10]), .A1(n8), .B0(dout4x4_2[10]), .B1(n9), 
        .C0(dout4x4_1[10]), .C1(n10), .Y(n37) );
  AOI222X1 U30 ( .A0(dout4x4_3[10]), .A1(n5), .B0(dout8x8_1[10]), .B1(n6), 
        .C0(dout4x4_4[10]), .C1(n7), .Y(n38) );
  NAND2X1 U31 ( .A(n35), .B(n36), .Y(ram_out_wire[11]) );
  AOI222X1 U32 ( .A0(dout8x8_2[11]), .A1(n8), .B0(dout4x4_2[11]), .B1(n9), 
        .C0(dout4x4_1[11]), .C1(n10), .Y(n35) );
  AOI222X1 U33 ( .A0(dout4x4_3[11]), .A1(n5), .B0(dout8x8_1[11]), .B1(n6), 
        .C0(dout4x4_4[11]), .C1(n7), .Y(n36) );
  NAND2X1 U34 ( .A(n33), .B(n34), .Y(ram_out_wire[12]) );
  AOI222X1 U35 ( .A0(dout8x8_2[12]), .A1(n8), .B0(dout4x4_2[12]), .B1(n9), 
        .C0(dout4x4_1[12]), .C1(n10), .Y(n33) );
  AOI222X1 U36 ( .A0(dout4x4_3[12]), .A1(n5), .B0(dout8x8_1[12]), .B1(n6), 
        .C0(dout4x4_4[12]), .C1(n7), .Y(n34) );
  NAND2X1 U37 ( .A(n39), .B(n40), .Y(ram_out_wire[0]) );
  AOI222X1 U38 ( .A0(dout8x8_2[0]), .A1(n8), .B0(dout4x4_2[0]), .B1(n9), .C0(
        dout4x4_1[0]), .C1(n10), .Y(n39) );
  AOI222X1 U39 ( .A0(dout4x4_3[0]), .A1(n5), .B0(dout8x8_1[0]), .B1(n6), .C0(
        dout4x4_4[0]), .C1(n7), .Y(n40) );
  NAND2X1 U40 ( .A(n31), .B(n32), .Y(ram_out_wire[13]) );
  AOI222X1 U41 ( .A0(dout8x8_2[13]), .A1(n8), .B0(dout4x4_2[13]), .B1(n9), 
        .C0(dout4x4_1[13]), .C1(n10), .Y(n31) );
  AOI222X1 U42 ( .A0(dout4x4_3[13]), .A1(n5), .B0(dout8x8_1[13]), .B1(n6), 
        .C0(dout4x4_4[13]), .C1(n7), .Y(n32) );
  NAND2X1 U43 ( .A(n29), .B(n30), .Y(ram_out_wire[14]) );
  AOI222X1 U44 ( .A0(dout8x8_2[14]), .A1(n8), .B0(dout4x4_2[14]), .B1(n9), 
        .C0(dout4x4_1[14]), .C1(n10), .Y(n29) );
  AOI222X1 U45 ( .A0(dout4x4_3[14]), .A1(n5), .B0(dout8x8_1[14]), .B1(n6), 
        .C0(dout4x4_4[14]), .C1(n7), .Y(n30) );
  NAND2X1 U46 ( .A(n27), .B(n28), .Y(ram_out_wire[15]) );
  AOI222X1 U47 ( .A0(dout8x8_2[15]), .A1(n8), .B0(dout4x4_2[15]), .B1(n9), 
        .C0(dout4x4_1[15]), .C1(n10), .Y(n27) );
  AOI222X1 U48 ( .A0(dout4x4_3[15]), .A1(n5), .B0(dout8x8_1[15]), .B1(n6), 
        .C0(dout4x4_4[15]), .C1(n7), .Y(n28) );
  NOR4BX1 U49 ( .AN(n41), .B(n10), .C(n8), .D(n9), .Y(n6) );
  NOR2X1 U50 ( .A(n5), .B(n7), .Y(n41) );
  NAND2X1 U51 ( .A(n43), .B(n42), .Y(mem_ctrl_tran_ready) );
  NOR4BBX1 U52 ( .AN(n42), .BN(ram8x8_2_ready), .C(ram8x8_1_ready), .D(
        ram4x4_4_ready), .Y(n8) );
  NOR4BX1 U53 ( .AN(n43), .B(n1), .C(ram4x4_1_ready), .D(ram4x4_2_ready), .Y(
        n5) );
  NOR4BX1 U54 ( .AN(n43), .B(n2), .C(ram4x4_1_ready), .D(ram4x4_3_ready), .Y(
        n9) );
  NOR4BBX1 U55 ( .AN(n42), .BN(ram4x4_4_ready), .C(ram8x8_1_ready), .D(
        ram8x8_2_ready), .Y(n7) );
  NOR3X1 U56 ( .A(ram8x8_1_ready), .B(ram8x8_2_ready), .C(ram4x4_4_ready), .Y(
        n43) );
  AND4X2 U57 ( .A(ram4x4_1_ready), .B(n43), .C(n2), .D(n1), .Y(n10) );
  NOR3X1 U58 ( .A(ram4x4_2_ready), .B(ram4x4_3_ready), .C(ram4x4_1_ready), .Y(
        n42) );
  INVX1 U59 ( .A(ram4x4_3_ready), .Y(n1) );
  INVX1 U60 ( .A(ram4x4_2_ready), .Y(n2) );
endmodule


module idct_chip ( clk, rstn, mode, start, din, dout, dout_mode );
  input [1:0] mode;
  input [15:0] din;
  output [15:0] dout;
  output [1:0] dout_mode;
  input clk, rstn, start;
  wire   net_clk, net_rstn, net_start;
  wire   [1:0] net_mode;
  wire   [15:0] net_din;
  wire   [15:0] net_dout;
  wire   [1:0] net_dout_mode;

  PIW PIW_clk ( .PAD(clk), .C(net_clk) );
  PIW PIW_rstn ( .PAD(rstn), .C(net_rstn) );
  PIW PIW_start ( .PAD(start), .C(net_start) );
  PIW PIW_mode0 ( .PAD(mode[0]), .C(net_mode[0]) );
  PIW PIW_mode1 ( .PAD(mode[1]), .C(net_mode[1]) );
  PIW PIW_din0 ( .PAD(din[0]), .C(net_din[0]) );
  PIW PIW_din1 ( .PAD(din[1]), .C(net_din[1]) );
  PIW PIW_din2 ( .PAD(din[2]), .C(net_din[2]) );
  PIW PIW_din3 ( .PAD(din[3]), .C(net_din[3]) );
  PIW PIW_din4 ( .PAD(din[4]), .C(net_din[4]) );
  PIW PIW_din5 ( .PAD(din[5]), .C(net_din[5]) );
  PIW PIW_din6 ( .PAD(din[6]), .C(net_din[6]) );
  PIW PIW_din7 ( .PAD(din[7]), .C(net_din[7]) );
  PIW PIW_din8 ( .PAD(din[8]), .C(net_din[8]) );
  PIW PIW_din9 ( .PAD(din[9]), .C(net_din[9]) );
  PIW PIW_din10 ( .PAD(din[10]), .C(net_din[10]) );
  PIW PIW_din11 ( .PAD(din[11]), .C(net_din[11]) );
  PIW PIW_din12 ( .PAD(din[12]), .C(net_din[12]) );
  PIW PIW_din13 ( .PAD(din[13]), .C(net_din[13]) );
  PIW PIW_din14 ( .PAD(din[14]), .C(net_din[14]) );
  PIW PIW_din15 ( .PAD(din[15]), .C(net_din[15]) );
  PO8W PO8W_dout0 ( .I(net_dout[0]), .PAD(dout[0]) );
  PO8W PO8W_dout1 ( .I(net_dout[1]), .PAD(dout[1]) );
  PO8W PO8W_dout2 ( .I(net_dout[2]), .PAD(dout[2]) );
  PO8W PO8W_dout3 ( .I(net_dout[3]), .PAD(dout[3]) );
  PO8W PO8W_dout4 ( .I(net_dout[4]), .PAD(dout[4]) );
  PO8W PO8W_dout5 ( .I(net_dout[5]), .PAD(dout[5]) );
  PO8W PO8W_dout6 ( .I(net_dout[6]), .PAD(dout[6]) );
  PO8W PO8W_dout7 ( .I(net_dout[7]), .PAD(dout[7]) );
  PO8W PO8W_dout8 ( .I(net_dout[8]), .PAD(dout[8]) );
  PO8W PO8W_dout9 ( .I(net_dout[9]), .PAD(dout[9]) );
  PO8W PO8W_dout10 ( .I(net_dout[10]), .PAD(dout[10]) );
  PO8W PO8W_dout11 ( .I(net_dout[11]), .PAD(dout[11]) );
  PO8W PO8W_dout12 ( .I(net_dout[12]), .PAD(dout[12]) );
  PO8W PO8W_dout13 ( .I(net_dout[13]), .PAD(dout[13]) );
  PO8W PO8W_dout14 ( .I(net_dout[14]), .PAD(dout[14]) );
  PO8W PO8W_dout15 ( .I(net_dout[15]), .PAD(dout[15]) );
  PO8W PO8W_dout_mode0 ( .I(net_dout_mode[0]), .PAD(dout_mode[0]) );
  PO8W PO8W_dout_mode1 ( .I(net_dout_mode[1]), .PAD(dout_mode[1]) );
  idct inst_idct ( .clk(net_clk), .rstn(net_rstn), .mode(net_mode), .start(
        net_start), .din(net_din), .dout(net_dout), .dout_mode(net_dout_mode)
         );
endmodule

